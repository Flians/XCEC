//
// Conformal-LEC Version 20.10-d213 (02-Sep-2020)
//
module top(RIae76b68_57,RIae76be0_58,RIae78a58_123,RIae78ad0_124,RIae76028_33,RIae760a0_34,RIae76118_35,RIae76190_36,RIae762f8_39,
        RIae76370_40,RIae76208_37,RIae76280_38,RIae763e8_41,RIae76460_42,RIae764d8_43,RIae76550_44,RIae76730_48,RIae766b8_47,RIae76640_46,
        RIae765c8_45,RIae76988_53,RIae76a00_54,RIae76a78_55,RIae76af0_56,RIae767a8_49,RIae76820_50,RIae76898_51,RIae76910_52,RIae77798_83,
        RIae77810_84,RIae77888_85,RIae77900_86,RIae77a68_89,RIae77ae0_90,RIae77978_87,RIae779f0_88,RIae77108_69,RIae77180_70,RIae77018_67,
        RIae77090_68,RIae772e8_73,RIae77360_74,RIae771f8_71,RIae77270_72,RIae76c58_59,RIae76cd0_60,RIae76d48_61,RIae76dc0_62,RIae76f28_65,
        RIae76fa0_66,RIae76e38_63,RIae76eb0_64,RIae780f8_103,RIae78170_104,RIae782d8_107,RIae78350_108,RIae77f18_99,RIae77f90_100,RIae78008_101,
        RIae78080_102,RIae77e28_97,RIae77ea0_98,RIae78698_115,RIae78710_116,RIae78968_121,RIae789e0_122,RIae78878_119,RIae788f0_120,RIae78788_117,
        RIae78800_118,RIae77b58_91,RIae77bd0_92,RIae77c48_93,RIae77cc0_94,RIae77d38_95,RIae77db0_96,RIae785a8_113,RIae78620_114,RIae781e8_105,
        RIae78260_106,RIae784b8_111,RIae78530_112,RIae783c8_109,RIae78440_110,RIae774c8_77,RIae77540_78,RIae776a8_81,RIae77720_82,RIae77450_76,
        RIae773d8_75,RIae775b8_79,RIae77630_80,RIae755d8_11,RIae75650_12,RIae754e8_9,RIae75560_10,RIae75830_16,RIae757b8_15,RIae756c8_13,
        RIae75740_14,RIae75380_6,RIae75308_5,RIae75218_3,RIae75290_4,RIae75128_1,RIae751a0_2,RIae753f8_7,RIae75470_8,RIae75998_19,
        RIae75a10_20,RIae758a8_17,RIae75920_18,RIae75b78_23,RIae75bf0_24,RIae75a88_21,RIae75b00_22,RIae75e48_29,RIae75ec0_30,RIae75f38_31,
        RIae75fb0_32,RIae75c68_25,RIae75ce0_26,RIae75d58_27,RIae75dd0_28,RIae78cb0_128,RIae78d28_129,RIae78f80_134,RIae79070_136,RIae790e8_137,
        RIae78da0_130,RIae78e18_131,RIae78b48_125,RIae78bc0_126,RIae78c38_127,RIae78e90_132,RIae78ff8_135,RIae79160_138,RIae791d8_139,RIae79250_140,
        RIae792c8_141,RIae78f08_133,RIae79340_142,RIae793b8_143,RIae79ac0_158,RIae79b38_159,RIae79688_149,RIae799d0_156,RIae79610_148,RIae798e0_154,
        RIae79958_155,RIae794a8_145,RIae79700_150,RIae797f0_152,RIae79778_151,RIae79598_147,RIae79430_144,RIae79520_146,RIae79a48_157,RIae79868_153,
        RIae79ca0_162,RIae79d18_163,RIae79c28_161,RIae79bb0_160,RIae79d90_164,RIae79e08_165,RIae79e80_166,RIae79ef8_167,RIae79fe8_169,RIae79f70_168,
        RIae7a6f0_184,RIae7a858_187,RIae7a8d0_188,RIae7a2b8_175,RIae7a678_183,RIae7a768_185,RIae7a7e0_186,RIae7a510_180,RIae7a600_182,RIae7a3a8_177,
        RIae7a240_174,RIae7a330_176,RIae7a948_189,RIae7a060_170,RIae7a150_172,RIae7a0d8_171,RIae7a1c8_173,RIae7a9c0_190,RIae7aa38_191,RIae7a588_181,
        RIae7a498_179,RIae7a420_178,RIae7aab0_192,RIae7aee8_201,RIae7af60_202,RIae7afd8_203,RIae7b050_204,RIae7b0c8_205,RIae7b140_206,RIae7b230_208,
        RIae7b1b8_207,RIae7ab28_193,RIae7aba0_194,RIae7ac90_196,RIae7ac18_195,RIae7ad08_197,RIae7ad80_198,RIae7adf8_199,RIae7ae70_200,RIae7ba28_225,
        RIae7baa0_226,RIae7bb18_227,RIae7bb90_228,RIae7bed8_235,RIae7bf50_236,RIae7bde8_233,RIae7be60_234,RIae7b848_221,RIae7b8c0_222,RIae7b9b0_224,
        RIae7b938_223,RIae7b668_217,RIae7b6e0_218,RIae7b758_219,RIae7b7d0_220,RIae7bfc8_237,RIae7c040_238,RIae7c0b8_239,RIae7c130_240,RIae7c658_251,
        RIae7c6d0_252,RIae7bc08_229,RIae7bc80_230,RIae7c748_253,RIae7c7c0_254,RIae7c8b0_256,RIae7c838_255,RIae7bcf8_231,RIae7bd70_232,RIae7c568_249,
        RIae7c5e0_250,RIae7c388_245,RIae7c400_246,RIae7c478_247,RIae7c4f0_248,RIae7c1a8_241,RIae7c220_242,RIae7c298_243,RIae7c310_244,RIae7b488_213,
        RIae7b500_214,RIae7b5f0_216,RIae7b578_215,RIae7b398_211,RIae7b410_212,RIae7b2a8_209,RIae7b320_210,R_101_77c8620,R_102_af8fd30,R_103_af901c8,
        R_104_af9a140,R_105_af99768,R_106_af8be30,R_107_77c1150,R_108_af8ddb0,R_109_af8f010,R_10a_af996c0,R_10b_77c34c0,R_10c_77c28f0,R_10d_af8d090,
        R_10e_77ca5a0,R_10f_77ce4a0,R_110_77cd780,R_111_af8f2b0,R_112_77c6550,R_113_af98ee0,R_114_77c2068,R_115_af99ea0,R_116_77c0eb0,R_117_77cc280,
        R_118_77bf860,R_119_77c9f10,R_11a_af8bf80,R_11b_77bf320,R_11c_77c4fa8,R_11d_af99ab0,R_11e_77ca258,R_11f_af92880,R_120_af91c08,R_121_af92298,
        R_122_af99ca8,R_123_af990d8,R_124_77c5638,R_125_af8e6e0,R_126_77c3aa8,R_127_77c8d58,R_128_77c1fc0,R_129_77c6748,R_12a_77c3370,R_12b_af99d50,
        R_12c_77c5248,R_12d_77ca840,R_12e_af8eec0,R_12f_77c1498,R_130_77c5398,R_131_77c0820,R_132_af8d480,R_133_77ce890,R_134_af97c80,R_135_77c65f8,
        R_136_af8d678,R_137_77c3e98,R_138_af8e0f8,R_139_af99378,R_13a_77c7078,R_13b_77ce740,R_13c_af97fc8,R_13d_77c62b0,R_13e_77c27a0,R_13f_af979e0,
        R_140_77c25a8,R_141_af921f0,R_142_af8b7a0,R_143_77bfcf8,R_144_af92148,R_145_77c1c78,R_146_77cb560,R_147_af99960,R_148_af92490,R_149_77c9298,
        R_14a_77cb170,R_14b_af98268,R_14c_77bf9b0,R_14d_af91b60,R_14e_af8f208,R_14f_77c7a50,R_150_af99030,R_151_77c67f0,R_152_af8c370,R_153_77c8818,
        R_154_77c6d30,R_155_af98c40,R_156_77c9538,R_157_af96f60,R_158_af96d68,R_159_af8d870,R_15a_af8e830,R_15b_77ccbb0,R_15c_af8c610,R_15d_77c6898,
        R_15e_af8cb50,R_15f_af92538,R_160_af975f0,R_161_77c71c8,R_162_af8d720,R_163_77cb608,R_164_af8b650,R_165_af988f8,R_166_77c41e0,R_167_af8e398,
        R_168_af974a0,R_169_af8d330,R_16a_af8c0d0,R_16b_77cc520,R_16c_77cb8a8,R_16d_77ccda8,R_16e_af973f8,R_16f_77cd6d8,R_170_af99ff0,R_171_77c54e8,
        R_172_77c3808,R_173_77c0580,R_174_af99618,R_175_77cd198,R_176_77c0628,R_177_af97698);
input RIae76b68_57,RIae76be0_58,RIae78a58_123,RIae78ad0_124,RIae76028_33,RIae760a0_34,RIae76118_35,RIae76190_36,RIae762f8_39,
        RIae76370_40,RIae76208_37,RIae76280_38,RIae763e8_41,RIae76460_42,RIae764d8_43,RIae76550_44,RIae76730_48,RIae766b8_47,RIae76640_46,
        RIae765c8_45,RIae76988_53,RIae76a00_54,RIae76a78_55,RIae76af0_56,RIae767a8_49,RIae76820_50,RIae76898_51,RIae76910_52,RIae77798_83,
        RIae77810_84,RIae77888_85,RIae77900_86,RIae77a68_89,RIae77ae0_90,RIae77978_87,RIae779f0_88,RIae77108_69,RIae77180_70,RIae77018_67,
        RIae77090_68,RIae772e8_73,RIae77360_74,RIae771f8_71,RIae77270_72,RIae76c58_59,RIae76cd0_60,RIae76d48_61,RIae76dc0_62,RIae76f28_65,
        RIae76fa0_66,RIae76e38_63,RIae76eb0_64,RIae780f8_103,RIae78170_104,RIae782d8_107,RIae78350_108,RIae77f18_99,RIae77f90_100,RIae78008_101,
        RIae78080_102,RIae77e28_97,RIae77ea0_98,RIae78698_115,RIae78710_116,RIae78968_121,RIae789e0_122,RIae78878_119,RIae788f0_120,RIae78788_117,
        RIae78800_118,RIae77b58_91,RIae77bd0_92,RIae77c48_93,RIae77cc0_94,RIae77d38_95,RIae77db0_96,RIae785a8_113,RIae78620_114,RIae781e8_105,
        RIae78260_106,RIae784b8_111,RIae78530_112,RIae783c8_109,RIae78440_110,RIae774c8_77,RIae77540_78,RIae776a8_81,RIae77720_82,RIae77450_76,
        RIae773d8_75,RIae775b8_79,RIae77630_80,RIae755d8_11,RIae75650_12,RIae754e8_9,RIae75560_10,RIae75830_16,RIae757b8_15,RIae756c8_13,
        RIae75740_14,RIae75380_6,RIae75308_5,RIae75218_3,RIae75290_4,RIae75128_1,RIae751a0_2,RIae753f8_7,RIae75470_8,RIae75998_19,
        RIae75a10_20,RIae758a8_17,RIae75920_18,RIae75b78_23,RIae75bf0_24,RIae75a88_21,RIae75b00_22,RIae75e48_29,RIae75ec0_30,RIae75f38_31,
        RIae75fb0_32,RIae75c68_25,RIae75ce0_26,RIae75d58_27,RIae75dd0_28,RIae78cb0_128,RIae78d28_129,RIae78f80_134,RIae79070_136,RIae790e8_137,
        RIae78da0_130,RIae78e18_131,RIae78b48_125,RIae78bc0_126,RIae78c38_127,RIae78e90_132,RIae78ff8_135,RIae79160_138,RIae791d8_139,RIae79250_140,
        RIae792c8_141,RIae78f08_133,RIae79340_142,RIae793b8_143,RIae79ac0_158,RIae79b38_159,RIae79688_149,RIae799d0_156,RIae79610_148,RIae798e0_154,
        RIae79958_155,RIae794a8_145,RIae79700_150,RIae797f0_152,RIae79778_151,RIae79598_147,RIae79430_144,RIae79520_146,RIae79a48_157,RIae79868_153,
        RIae79ca0_162,RIae79d18_163,RIae79c28_161,RIae79bb0_160,RIae79d90_164,RIae79e08_165,RIae79e80_166,RIae79ef8_167,RIae79fe8_169,RIae79f70_168,
        RIae7a6f0_184,RIae7a858_187,RIae7a8d0_188,RIae7a2b8_175,RIae7a678_183,RIae7a768_185,RIae7a7e0_186,RIae7a510_180,RIae7a600_182,RIae7a3a8_177,
        RIae7a240_174,RIae7a330_176,RIae7a948_189,RIae7a060_170,RIae7a150_172,RIae7a0d8_171,RIae7a1c8_173,RIae7a9c0_190,RIae7aa38_191,RIae7a588_181,
        RIae7a498_179,RIae7a420_178,RIae7aab0_192,RIae7aee8_201,RIae7af60_202,RIae7afd8_203,RIae7b050_204,RIae7b0c8_205,RIae7b140_206,RIae7b230_208,
        RIae7b1b8_207,RIae7ab28_193,RIae7aba0_194,RIae7ac90_196,RIae7ac18_195,RIae7ad08_197,RIae7ad80_198,RIae7adf8_199,RIae7ae70_200,RIae7ba28_225,
        RIae7baa0_226,RIae7bb18_227,RIae7bb90_228,RIae7bed8_235,RIae7bf50_236,RIae7bde8_233,RIae7be60_234,RIae7b848_221,RIae7b8c0_222,RIae7b9b0_224,
        RIae7b938_223,RIae7b668_217,RIae7b6e0_218,RIae7b758_219,RIae7b7d0_220,RIae7bfc8_237,RIae7c040_238,RIae7c0b8_239,RIae7c130_240,RIae7c658_251,
        RIae7c6d0_252,RIae7bc08_229,RIae7bc80_230,RIae7c748_253,RIae7c7c0_254,RIae7c8b0_256,RIae7c838_255,RIae7bcf8_231,RIae7bd70_232,RIae7c568_249,
        RIae7c5e0_250,RIae7c388_245,RIae7c400_246,RIae7c478_247,RIae7c4f0_248,RIae7c1a8_241,RIae7c220_242,RIae7c298_243,RIae7c310_244,RIae7b488_213,
        RIae7b500_214,RIae7b5f0_216,RIae7b578_215,RIae7b398_211,RIae7b410_212,RIae7b2a8_209,RIae7b320_210;
output R_101_77c8620,R_102_af8fd30,R_103_af901c8,R_104_af9a140,R_105_af99768,R_106_af8be30,R_107_77c1150,R_108_af8ddb0,R_109_af8f010,
        R_10a_af996c0,R_10b_77c34c0,R_10c_77c28f0,R_10d_af8d090,R_10e_77ca5a0,R_10f_77ce4a0,R_110_77cd780,R_111_af8f2b0,R_112_77c6550,R_113_af98ee0,
        R_114_77c2068,R_115_af99ea0,R_116_77c0eb0,R_117_77cc280,R_118_77bf860,R_119_77c9f10,R_11a_af8bf80,R_11b_77bf320,R_11c_77c4fa8,R_11d_af99ab0,
        R_11e_77ca258,R_11f_af92880,R_120_af91c08,R_121_af92298,R_122_af99ca8,R_123_af990d8,R_124_77c5638,R_125_af8e6e0,R_126_77c3aa8,R_127_77c8d58,
        R_128_77c1fc0,R_129_77c6748,R_12a_77c3370,R_12b_af99d50,R_12c_77c5248,R_12d_77ca840,R_12e_af8eec0,R_12f_77c1498,R_130_77c5398,R_131_77c0820,
        R_132_af8d480,R_133_77ce890,R_134_af97c80,R_135_77c65f8,R_136_af8d678,R_137_77c3e98,R_138_af8e0f8,R_139_af99378,R_13a_77c7078,R_13b_77ce740,
        R_13c_af97fc8,R_13d_77c62b0,R_13e_77c27a0,R_13f_af979e0,R_140_77c25a8,R_141_af921f0,R_142_af8b7a0,R_143_77bfcf8,R_144_af92148,R_145_77c1c78,
        R_146_77cb560,R_147_af99960,R_148_af92490,R_149_77c9298,R_14a_77cb170,R_14b_af98268,R_14c_77bf9b0,R_14d_af91b60,R_14e_af8f208,R_14f_77c7a50,
        R_150_af99030,R_151_77c67f0,R_152_af8c370,R_153_77c8818,R_154_77c6d30,R_155_af98c40,R_156_77c9538,R_157_af96f60,R_158_af96d68,R_159_af8d870,
        R_15a_af8e830,R_15b_77ccbb0,R_15c_af8c610,R_15d_77c6898,R_15e_af8cb50,R_15f_af92538,R_160_af975f0,R_161_77c71c8,R_162_af8d720,R_163_77cb608,
        R_164_af8b650,R_165_af988f8,R_166_77c41e0,R_167_af8e398,R_168_af974a0,R_169_af8d330,R_16a_af8c0d0,R_16b_77cc520,R_16c_77cb8a8,R_16d_77ccda8,
        R_16e_af973f8,R_16f_77cd6d8,R_170_af99ff0,R_171_77c54e8,R_172_77c3808,R_173_77c0580,R_174_af99618,R_175_77cd198,R_176_77c0628,R_177_af97698;

wire \376_ZERO , \377_ONE , \378 , \379 , \380 , \381 , \382 , \383 , \384 ,
         \385 , \386 , \387 , \388 , \389 , \390 , \391 , \392 , \393 , \394 ,
         \395 , \396 , \397 , \398 , \399 , \400 , \401 , \402 , \403 , \404 ,
         \405 , \406 , \407 , \408 , \409 , \410 , \411 , \412 , \413 , \414 ,
         \415 , \416 , \417 , \418 , \419 , \420 , \421 , \422 , \423 , \424 ,
         \425 , \426 , \427 , \428 , \429 , \430 , \431 , \432 , \433 , \434 ,
         \435 , \436 , \437 , \438 , \439 , \440 , \441 , \442 , \443 , \444 ,
         \445 , \446 , \447 , \448 , \449 , \450 , \451 , \452 , \453 , \454 ,
         \455 , \456 , \457 , \458 , \459 , \460 , \461 , \462 , \463 , \464 ,
         \465 , \466 , \467 , \468 , \469 , \470 , \471 , \472 , \473 , \474 ,
         \475 , \476 , \477 , \478 , \479 , \480 , \481 , \482 , \483 , \484 ,
         \485 , \486 , \487 , \488 , \489 , \490 , \491 , \492 , \493 , \494 ,
         \495 , \496 , \497 , \498 , \499 , \500 , \501 , \502 , \503 , \504 ,
         \505 , \506 , \507 , \508 , \509 , \510 , \511 , \512 , \513 , \514 ,
         \515 , \516 , \517 , \518 , \519 , \520 , \521 , \522 , \523 , \524 ,
         \525 , \526 , \527 , \528 , \529 , \530 , \531 , \532 , \533 , \534 ,
         \535 , \536 , \537 , \538 , \539 , \540 , \541 , \542 , \543 , \544 ,
         \545 , \546 , \547 , \548 , \549 , \550 , \551 , \552 , \553 , \554 ,
         \555 , \556 , \557 , \558 , \559 , \560 , \561 , \562 , \563 , \564 ,
         \565 , \566 , \567 , \568 , \569 , \570 , \571 , \572 , \573 , \574 ,
         \575 , \576 , \577 , \578 , \579 , \580 , \581 , \582 , \583 , \584 ,
         \585 , \586 , \587 , \588 , \589 , \590 , \591 , \592 , \593 , \594 ,
         \595 , \596 , \597 , \598 , \599 , \600 , \601 , \602 , \603 , \604 ,
         \605 , \606 , \607 , \608 , \609 , \610 , \611 , \612 , \613 , \614 ,
         \615 , \616 , \617 , \618 , \619 , \620 , \621 , \622 , \623 , \624 ,
         \625 , \626 , \627 , \628 , \629 , \630 , \631 , \632 , \633 , \634 ,
         \635 , \636 , \637 , \638 , \639 , \640 , \641 , \642 , \643 , \644 ,
         \645 , \646 , \647 , \648 , \649 , \650 , \651 , \652 , \653 , \654 ,
         \655 , \656 , \657 , \658 , \659 , \660 , \661 , \662 , \663 , \664 ,
         \665 , \666 , \667 , \668 , \669 , \670 , \671 , \672 , \673 , \674 ,
         \675 , \676 , \677 , \678 , \679 , \680 , \681 , \682 , \683 , \684 ,
         \685 , \686 , \687 , \688 , \689 , \690 , \691 , \692 , \693 , \694 ,
         \695 , \696 , \697 , \698 , \699 , \700 , \701 , \702 , \703 , \704 ,
         \705 , \706 , \707 , \708 , \709 , \710 , \711 , \712 , \713 , \714 ,
         \715 , \716 , \717 , \718 , \719 , \720 , \721 , \722 , \723 , \724 ,
         \725 , \726 , \727 , \728 , \729 , \730 , \731 , \732 , \733 , \734 ,
         \735 , \736 , \737 , \738 , \739 , \740 , \741 , \742 , \743 , \744 ,
         \745 , \746 , \747 , \748 , \749 , \750 , \751 , \752 , \753 , \754 ,
         \755 , \756 , \757 , \758 , \759 , \760 , \761 , \762 , \763 , \764 ,
         \765 , \766 , \767 , \768 , \769 , \770 , \771 , \772 , \773 , \774 ,
         \775 , \776 , \777 , \778 , \779 , \780 , \781 , \782 , \783 , \784 ,
         \785 , \786 , \787 , \788 , \789 , \790 , \791 , \792 , \793 , \794 ,
         \795 , \796 , \797 , \798 , \799 , \800 , \801 , \802 , \803 , \804 ,
         \805 , \806 , \807 , \808 , \809 , \810 , \811 , \812 , \813 , \814 ,
         \815 , \816 , \817 , \818 , \819 , \820 , \821 , \822 , \823 , \824 ,
         \825 , \826 , \827 , \828 , \829 , \830 , \831 , \832 , \833 , \834 ,
         \835 , \836 , \837 , \838 , \839 , \840 , \841 , \842 , \843 , \844 ,
         \845 , \846 , \847 , \848 , \849 , \850 , \851 , \852 , \853 , \854 ,
         \855 , \856 , \857 , \858 , \859 , \860 , \861 , \862 , \863 , \864 ,
         \865 , \866 , \867 , \868 , \869 , \870 , \871 , \872 , \873 , \874 ,
         \875 , \876 , \877 , \878 , \879 , \880 , \881 , \882 , \883 , \884 ,
         \885 , \886 , \887 , \888 , \889 , \890 , \891 , \892 , \893 , \894 ,
         \895 , \896 , \897 , \898 , \899 , \900 , \901 , \902 , \903 , \904 ,
         \905 , \906 , \907 , \908 , \909 , \910 , \911 , \912 , \913 , \914 ,
         \915 , \916 , \917 , \918 , \919 , \920 , \921 , \922 , \923 , \924 ,
         \925 , \926 , \927 , \928 , \929 , \930 , \931 , \932 , \933 , \934 ,
         \935 , \936 , \937 , \938 , \939 , \940 , \941 , \942 , \943 , \944 ,
         \945 , \946 , \947 , \948 , \949 , \950 , \951 , \952 , \953 , \954 ,
         \955 , \956 , \957 , \958 , \959 , \960 , \961 , \962 , \963 , \964 ,
         \965 , \966 , \967 , \968 , \969 , \970 , \971 , \972 , \973 , \974 ,
         \975 , \976 , \977 , \978 , \979 , \980 , \981 , \982 , \983 , \984 ,
         \985 , \986 , \987 , \988 , \989 , \990 , \991 , \992 , \993 , \994 ,
         \995 , \996 , \997 , \998 , \999 , \1000 , \1001 , \1002 , \1003 , \1004 ,
         \1005 , \1006 , \1007 , \1008 , \1009 , \1010 , \1011 , \1012 , \1013 , \1014 ,
         \1015 , \1016 , \1017 , \1018 , \1019 , \1020 , \1021 , \1022 , \1023 , \1024 ,
         \1025 , \1026 , \1027 , \1028 , \1029 , \1030 , \1031 , \1032 , \1033 , \1034 ,
         \1035 , \1036 , \1037 , \1038 , \1039 , \1040 , \1041 , \1042 , \1043 , \1044 ,
         \1045 , \1046 , \1047 , \1048 , \1049 , \1050 , \1051 , \1052 , \1053 , \1054 ,
         \1055 , \1056 , \1057 , \1058 , \1059 , \1060 , \1061 , \1062 , \1063 , \1064 ,
         \1065 , \1066 , \1067 , \1068 , \1069 , \1070 , \1071 , \1072 , \1073 , \1074 ,
         \1075 , \1076 , \1077 , \1078 , \1079 , \1080 , \1081 , \1082 , \1083 , \1084 ,
         \1085 , \1086 , \1087 , \1088 , \1089 , \1090 , \1091 , \1092 , \1093 , \1094 ,
         \1095 , \1096 , \1097 , \1098 , \1099 , \1100 , \1101 , \1102 , \1103 , \1104 ,
         \1105 , \1106 , \1107 , \1108 , \1109 , \1110 , \1111 , \1112 , \1113 , \1114 ,
         \1115 , \1116 , \1117 , \1118 , \1119 , \1120 , \1121 , \1122 , \1123 , \1124 ,
         \1125 , \1126 , \1127 , \1128 , \1129 , \1130 , \1131 , \1132 , \1133 , \1134 ,
         \1135 , \1136 , \1137 , \1138 , \1139 , \1140 , \1141 , \1142 , \1143 , \1144 ,
         \1145 , \1146 , \1147 , \1148 , \1149 , \1150 , \1151 , \1152 , \1153 , \1154 ,
         \1155 , \1156 , \1157 , \1158 , \1159 , \1160 , \1161 , \1162 , \1163 , \1164 ,
         \1165 , \1166 , \1167 , \1168 , \1169 , \1170 , \1171 , \1172 , \1173 , \1174 ,
         \1175 , \1176 , \1177 , \1178 , \1179 , \1180 , \1181 , \1182 , \1183 , \1184 ,
         \1185 , \1186 , \1187 , \1188 , \1189 , \1190 , \1191 , \1192 , \1193 , \1194 ,
         \1195 , \1196 , \1197 , \1198 , \1199 , \1200 , \1201 , \1202 , \1203 , \1204 ,
         \1205 , \1206 , \1207 , \1208 , \1209 , \1210 , \1211 , \1212 , \1213 , \1214 ,
         \1215 , \1216 , \1217 , \1218 , \1219 , \1220 , \1221 , \1222 , \1223 , \1224 ,
         \1225 , \1226 , \1227 , \1228 , \1229 , \1230 , \1231 , \1232 , \1233 , \1234 ,
         \1235 , \1236 , \1237 , \1238 , \1239 , \1240 , \1241 , \1242 , \1243 , \1244 ,
         \1245 , \1246 , \1247 , \1248 , \1249 , \1250 , \1251 , \1252 , \1253 , \1254 ,
         \1255 , \1256 , \1257 , \1258 , \1259 , \1260 , \1261 , \1262 , \1263 , \1264 ,
         \1265 , \1266 , \1267 , \1268 , \1269 , \1270 , \1271 , \1272 , \1273 , \1274 ,
         \1275 , \1276 , \1277 , \1278 , \1279 , \1280 , \1281 , \1282 , \1283 , \1284 ,
         \1285 , \1286 , \1287 , \1288 , \1289 , \1290 , \1291 , \1292 , \1293 , \1294 ,
         \1295 , \1296 , \1297 , \1298 , \1299 , \1300 , \1301 , \1302 , \1303 , \1304 ,
         \1305 , \1306 , \1307 , \1308 , \1309 , \1310 , \1311 , \1312 , \1313 , \1314 ,
         \1315 , \1316 , \1317 , \1318 , \1319 , \1320 , \1321 , \1322 , \1323 , \1324 ,
         \1325 , \1326 , \1327 , \1328 , \1329 , \1330 , \1331 , \1332 , \1333 , \1334 ,
         \1335 , \1336 , \1337 , \1338 , \1339 , \1340 , \1341 , \1342 , \1343 , \1344 ,
         \1345 , \1346 , \1347 , \1348 , \1349 , \1350 , \1351 , \1352 , \1353 , \1354 ,
         \1355 , \1356 , \1357 , \1358 , \1359 , \1360 , \1361 , \1362 , \1363 , \1364 ,
         \1365 , \1366 , \1367 , \1368 , \1369 , \1370 , \1371 , \1372 , \1373 , \1374 ,
         \1375 , \1376 , \1377 , \1378 , \1379 , \1380 , \1381 , \1382 , \1383 , \1384 ,
         \1385 , \1386 , \1387 , \1388 , \1389 , \1390 , \1391 , \1392 , \1393 , \1394 ,
         \1395 , \1396 , \1397 , \1398 , \1399 , \1400 , \1401 , \1402 , \1403 , \1404 ,
         \1405 , \1406 , \1407 , \1408 , \1409 , \1410 , \1411 , \1412 , \1413 , \1414 ,
         \1415 , \1416 , \1417 , \1418 , \1419 , \1420 , \1421 , \1422 , \1423 , \1424 ,
         \1425 , \1426 , \1427 , \1428 , \1429 , \1430 , \1431 , \1432 , \1433 , \1434 ,
         \1435 , \1436 , \1437 , \1438 , \1439 , \1440 , \1441 , \1442 , \1443 , \1444 ,
         \1445 , \1446 , \1447 , \1448 , \1449 , \1450 , \1451 , \1452 , \1453 , \1454 ,
         \1455 , \1456 , \1457 , \1458 , \1459 , \1460 , \1461 , \1462 , \1463 , \1464 ,
         \1465 , \1466 , \1467 , \1468 , \1469 , \1470 , \1471 , \1472 , \1473 , \1474 ,
         \1475 , \1476 , \1477 , \1478 , \1479 , \1480 , \1481 , \1482 , \1483 , \1484 ,
         \1485 , \1486 , \1487 , \1488 , \1489 , \1490 , \1491 , \1492 , \1493 , \1494 ,
         \1495 , \1496 , \1497 , \1498 , \1499 , \1500 , \1501 , \1502 , \1503 , \1504 ,
         \1505 , \1506 , \1507 , \1508 , \1509 , \1510 , \1511 , \1512 , \1513 , \1514 ,
         \1515 , \1516 , \1517 , \1518 , \1519 , \1520 , \1521 , \1522 , \1523 , \1524 ,
         \1525 , \1526 , \1527 , \1528 , \1529 , \1530 , \1531 , \1532 , \1533 , \1534 ,
         \1535 , \1536 , \1537 , \1538 , \1539 , \1540 , \1541 , \1542 , \1543 , \1544 ,
         \1545 , \1546 , \1547 , \1548 , \1549 , \1550 , \1551 , \1552 , \1553 , \1554 ,
         \1555 , \1556 , \1557 , \1558 , \1559 , \1560 , \1561 , \1562 , \1563 , \1564 ,
         \1565 , \1566 , \1567 , \1568 , \1569 , \1570 , \1571 , \1572 , \1573 , \1574 ,
         \1575 , \1576 , \1577 , \1578 , \1579 , \1580 , \1581 , \1582 , \1583 , \1584 ,
         \1585 , \1586 , \1587 , \1588 , \1589 , \1590 , \1591 , \1592 , \1593 , \1594 ,
         \1595 , \1596 , \1597 , \1598 , \1599 , \1600 , \1601 , \1602 , \1603 , \1604 ,
         \1605 , \1606 , \1607 , \1608 , \1609 , \1610 , \1611 , \1612 , \1613 , \1614 ,
         \1615 , \1616 , \1617 , \1618 , \1619 , \1620 , \1621 , \1622 , \1623 , \1624 ,
         \1625 , \1626 , \1627 , \1628 , \1629 , \1630 , \1631 , \1632 , \1633 , \1634 ,
         \1635 , \1636 , \1637 , \1638 , \1639 , \1640 , \1641 , \1642 , \1643 , \1644 ,
         \1645 , \1646 , \1647 , \1648 , \1649 , \1650 , \1651 , \1652 , \1653 , \1654 ,
         \1655 , \1656 , \1657 , \1658 , \1659 , \1660 , \1661 , \1662 , \1663 , \1664 ,
         \1665 , \1666 , \1667 , \1668 , \1669 , \1670 , \1671 , \1672 , \1673 , \1674 ,
         \1675 , \1676 , \1677 , \1678 , \1679 , \1680 , \1681 , \1682 , \1683 , \1684 ,
         \1685 , \1686 , \1687 , \1688 , \1689 , \1690 , \1691 , \1692 , \1693 , \1694 ,
         \1695 , \1696 , \1697 , \1698 , \1699 , \1700 , \1701 , \1702 , \1703 , \1704 ,
         \1705 , \1706 , \1707 , \1708 , \1709 , \1710 , \1711 , \1712 , \1713 , \1714 ,
         \1715 , \1716 , \1717 , \1718 , \1719 , \1720 , \1721 , \1722 , \1723 , \1724 ,
         \1725 , \1726 , \1727 , \1728 , \1729 , \1730 , \1731 , \1732 , \1733 , \1734 ,
         \1735 , \1736 , \1737 , \1738 , \1739 , \1740 , \1741 , \1742 , \1743 , \1744 ,
         \1745 , \1746 , \1747 , \1748 , \1749 , \1750 , \1751 , \1752 , \1753 , \1754 ,
         \1755 , \1756 , \1757 , \1758 , \1759 , \1760 , \1761 , \1762 , \1763 , \1764 ,
         \1765 , \1766 , \1767 , \1768 , \1769 , \1770 , \1771 , \1772 , \1773 , \1774 ,
         \1775 , \1776 , \1777 , \1778 , \1779 , \1780 , \1781 , \1782 , \1783 , \1784 ,
         \1785 , \1786 , \1787 , \1788 , \1789 , \1790 , \1791 , \1792 , \1793 , \1794 ,
         \1795 , \1796 , \1797 , \1798 , \1799 , \1800 , \1801 , \1802 , \1803 , \1804 ,
         \1805 , \1806 , \1807 , \1808 , \1809 , \1810 , \1811 , \1812 , \1813 , \1814 ,
         \1815 , \1816 , \1817 , \1818 , \1819 , \1820 , \1821 , \1822 , \1823 , \1824 ,
         \1825 , \1826 , \1827 , \1828 , \1829 , \1830 , \1831 , \1832 , \1833 , \1834 ,
         \1835 , \1836 , \1837 , \1838 , \1839 , \1840 , \1841 , \1842 , \1843 , \1844 ,
         \1845 , \1846 , \1847 , \1848 , \1849 , \1850 , \1851 , \1852 , \1853 , \1854 ,
         \1855 , \1856 , \1857 , \1858 , \1859 , \1860 , \1861 , \1862 , \1863 , \1864 ,
         \1865 , \1866 , \1867 , \1868 , \1869 , \1870 , \1871 , \1872 , \1873 , \1874 ,
         \1875 , \1876 , \1877 , \1878 , \1879 , \1880 , \1881 , \1882 , \1883 , \1884 ,
         \1885 , \1886 , \1887 , \1888 , \1889 , \1890 , \1891 , \1892 , \1893 , \1894 ,
         \1895 , \1896 , \1897 , \1898 , \1899 , \1900 , \1901 , \1902 , \1903 , \1904 ,
         \1905 , \1906 , \1907 , \1908 , \1909 , \1910 , \1911 , \1912 , \1913 , \1914 ,
         \1915 , \1916 , \1917 , \1918 , \1919 , \1920 , \1921 , \1922 , \1923 , \1924 ,
         \1925 , \1926 , \1927 , \1928 , \1929 , \1930 , \1931 , \1932 , \1933 , \1934 ,
         \1935 , \1936 , \1937 , \1938 , \1939 , \1940 , \1941 , \1942 , \1943 , \1944 ,
         \1945 , \1946 , \1947 , \1948 , \1949 , \1950 , \1951 , \1952 , \1953 , \1954 ,
         \1955 , \1956 , \1957 , \1958 , \1959 , \1960 , \1961 , \1962 , \1963 , \1964 ,
         \1965 , \1966 , \1967 , \1968 , \1969 , \1970 , \1971 , \1972 , \1973 , \1974 ,
         \1975 , \1976 , \1977 , \1978 , \1979 , \1980 , \1981 , \1982 , \1983 , \1984 ,
         \1985 , \1986 , \1987 , \1988 , \1989 , \1990 , \1991 , \1992 , \1993 , \1994 ,
         \1995 , \1996 , \1997 , \1998 , \1999 , \2000 , \2001 , \2002 , \2003 , \2004 ,
         \2005 , \2006 , \2007 , \2008 , \2009 , \2010 , \2011 , \2012 , \2013 , \2014 ,
         \2015 , \2016 , \2017 , \2018 , \2019 , \2020 , \2021 , \2022 , \2023 , \2024 ,
         \2025 , \2026 , \2027 , \2028 , \2029 , \2030 , \2031 , \2032 , \2033 , \2034 ,
         \2035 , \2036 , \2037 , \2038 , \2039 , \2040 , \2041 , \2042 , \2043 , \2044 ,
         \2045 , \2046 , \2047 , \2048 , \2049 , \2050 , \2051 , \2052 , \2053 , \2054 ,
         \2055 , \2056 , \2057 , \2058 , \2059 , \2060 , \2061 , \2062 , \2063 , \2064 ,
         \2065 , \2066 , \2067 , \2068 , \2069 , \2070 , \2071 , \2072 , \2073 , \2074 ,
         \2075 , \2076 , \2077 , \2078 , \2079 , \2080 , \2081 , \2082 , \2083 , \2084 ,
         \2085 , \2086 , \2087 , \2088 , \2089 , \2090 , \2091 , \2092 , \2093 , \2094 ,
         \2095 , \2096 , \2097 , \2098 , \2099 , \2100 , \2101 , \2102 , \2103 , \2104 ,
         \2105 , \2106 , \2107 , \2108 , \2109 , \2110 , \2111 , \2112 , \2113 , \2114 ,
         \2115 , \2116 , \2117 , \2118 , \2119 , \2120 , \2121 , \2122 , \2123 , \2124 ,
         \2125 , \2126 , \2127 , \2128 , \2129 , \2130 , \2131 , \2132 , \2133 , \2134 ,
         \2135 , \2136 , \2137 , \2138 , \2139 , \2140 , \2141 , \2142 , \2143 , \2144 ,
         \2145 , \2146 , \2147 , \2148 , \2149 , \2150 , \2151 , \2152 , \2153 , \2154 ,
         \2155 , \2156 , \2157 , \2158 , \2159 , \2160 , \2161 , \2162 , \2163 , \2164 ,
         \2165 , \2166 , \2167 , \2168 , \2169 , \2170 , \2171 , \2172 , \2173 , \2174 ,
         \2175 , \2176 , \2177 , \2178 , \2179 , \2180 , \2181 , \2182 , \2183 , \2184 ,
         \2185 , \2186 , \2187 , \2188 , \2189 , \2190 , \2191 , \2192 , \2193 , \2194 ,
         \2195 , \2196 , \2197 , \2198 , \2199 , \2200 , \2201 , \2202 , \2203 , \2204 ,
         \2205 , \2206 , \2207 , \2208 , \2209 , \2210 , \2211 , \2212 , \2213 , \2214 ,
         \2215 , \2216 , \2217 , \2218 , \2219 , \2220 , \2221 , \2222 , \2223 , \2224 ,
         \2225 , \2226 , \2227 , \2228 , \2229 , \2230 , \2231 , \2232 , \2233 , \2234 ,
         \2235 , \2236 , \2237 , \2238 , \2239 , \2240 , \2241 , \2242 , \2243 , \2244 ,
         \2245 , \2246 , \2247 , \2248 , \2249 , \2250 , \2251 , \2252 , \2253 , \2254 ,
         \2255 , \2256 , \2257 , \2258 , \2259 , \2260 , \2261 , \2262 , \2263 , \2264 ,
         \2265 , \2266 , \2267 , \2268 , \2269 , \2270 , \2271 , \2272 , \2273 , \2274 ,
         \2275 , \2276 , \2277 , \2278 , \2279 , \2280 , \2281 , \2282 , \2283 , \2284 ,
         \2285 , \2286 , \2287 , \2288 , \2289 , \2290 , \2291 , \2292 , \2293 , \2294 ,
         \2295 , \2296 , \2297 , \2298 , \2299 , \2300 , \2301 , \2302 , \2303 , \2304 ,
         \2305 , \2306 , \2307 , \2308 , \2309 , \2310 , \2311 , \2312 , \2313 , \2314 ,
         \2315 , \2316 , \2317 , \2318 , \2319 , \2320 , \2321 , \2322 , \2323 , \2324 ,
         \2325 , \2326 , \2327 , \2328 , \2329 , \2330 , \2331 , \2332 , \2333 , \2334 ,
         \2335 , \2336 , \2337 , \2338 , \2339 , \2340 , \2341 , \2342 , \2343 , \2344 ,
         \2345 , \2346 , \2347 , \2348 , \2349 , \2350 , \2351 , \2352 , \2353 , \2354 ,
         \2355 , \2356 , \2357 , \2358 , \2359 , \2360 , \2361 , \2362 , \2363 , \2364 ,
         \2365 , \2366 , \2367 , \2368 , \2369 , \2370 , \2371 , \2372 , \2373 , \2374 ,
         \2375 , \2376 , \2377 , \2378 , \2379 , \2380 , \2381 , \2382 , \2383 , \2384 ,
         \2385 , \2386 , \2387 , \2388 , \2389 , \2390 , \2391 , \2392 , \2393 , \2394 ,
         \2395 , \2396 , \2397 , \2398 , \2399 , \2400 , \2401 , \2402 , \2403 , \2404 ,
         \2405 , \2406 , \2407 , \2408 , \2409 , \2410 , \2411 , \2412 , \2413 , \2414 ,
         \2415 , \2416 , \2417 , \2418 , \2419 , \2420 , \2421 , \2422 , \2423 , \2424 ,
         \2425 , \2426 , \2427 , \2428 , \2429 , \2430 , \2431 , \2432 , \2433 , \2434 ,
         \2435 , \2436 , \2437 , \2438 , \2439 , \2440 , \2441 , \2442 , \2443 , \2444 ,
         \2445 , \2446 , \2447 , \2448 , \2449 , \2450 , \2451 , \2452 , \2453 , \2454 ,
         \2455 , \2456 , \2457 , \2458 , \2459 , \2460 , \2461 , \2462 , \2463 , \2464 ,
         \2465 , \2466 , \2467 , \2468 , \2469 , \2470 , \2471 , \2472 , \2473 , \2474 ,
         \2475 , \2476 , \2477 , \2478 , \2479 , \2480 , \2481 , \2482 , \2483 , \2484 ,
         \2485 , \2486 , \2487 , \2488 , \2489 , \2490 , \2491 , \2492 , \2493 , \2494 ,
         \2495 , \2496 , \2497 , \2498 , \2499 , \2500 , \2501 , \2502 , \2503 , \2504 ,
         \2505 , \2506 , \2507 , \2508 , \2509 , \2510 , \2511 , \2512 , \2513 , \2514 ,
         \2515 , \2516 , \2517 , \2518 , \2519 , \2520 , \2521 , \2522 , \2523 , \2524 ,
         \2525 , \2526 , \2527 , \2528 , \2529 , \2530 , \2531 , \2532 , \2533 , \2534 ,
         \2535 , \2536 , \2537 , \2538 , \2539 , \2540 , \2541 , \2542 , \2543 , \2544 ,
         \2545 , \2546 , \2547 , \2548 , \2549 , \2550 , \2551 , \2552 , \2553 , \2554 ,
         \2555 , \2556 , \2557 , \2558 , \2559 , \2560 , \2561 , \2562 , \2563 , \2564 ,
         \2565 , \2566 , \2567 , \2568 , \2569 , \2570 , \2571 , \2572 , \2573 , \2574 ,
         \2575 , \2576 , \2577 , \2578 , \2579 , \2580 , \2581 , \2582 , \2583 , \2584 ,
         \2585 , \2586 , \2587 , \2588 , \2589 , \2590 , \2591 , \2592 , \2593 , \2594 ,
         \2595 , \2596 , \2597 , \2598 , \2599 , \2600 , \2601 , \2602 , \2603 , \2604 ,
         \2605 , \2606 , \2607 , \2608 , \2609 , \2610 , \2611 , \2612 , \2613 , \2614 ,
         \2615 , \2616 , \2617 , \2618 , \2619 , \2620 , \2621 , \2622 , \2623 , \2624 ,
         \2625 , \2626 , \2627 , \2628 , \2629 , \2630 , \2631 , \2632 , \2633 , \2634 ,
         \2635 , \2636 , \2637 , \2638 , \2639 , \2640 , \2641 , \2642 , \2643 , \2644 ,
         \2645 , \2646 , \2647 , \2648 , \2649 , \2650 , \2651 , \2652 , \2653 , \2654 ,
         \2655 , \2656 , \2657 , \2658 , \2659 , \2660 , \2661 , \2662 , \2663 , \2664 ,
         \2665 , \2666 , \2667 , \2668 , \2669 , \2670 , \2671 , \2672 , \2673 , \2674 ,
         \2675 , \2676 , \2677 , \2678 , \2679 , \2680 , \2681 , \2682 , \2683 , \2684 ,
         \2685 , \2686 , \2687 , \2688 , \2689 , \2690 , \2691 , \2692 , \2693 , \2694 ,
         \2695 , \2696 , \2697 , \2698 , \2699 , \2700 , \2701 , \2702 , \2703 , \2704 ,
         \2705 , \2706 , \2707 , \2708 , \2709 , \2710 , \2711 , \2712 , \2713 , \2714 ,
         \2715 , \2716 , \2717 , \2718 , \2719 , \2720 , \2721 , \2722 , \2723 , \2724 ,
         \2725 , \2726 , \2727 , \2728 , \2729 , \2730 , \2731 , \2732 , \2733 , \2734 ,
         \2735 , \2736 , \2737 , \2738 , \2739 , \2740 , \2741 , \2742 , \2743 , \2744 ,
         \2745 , \2746 , \2747 , \2748 , \2749 , \2750 , \2751 , \2752 , \2753 , \2754 ,
         \2755 , \2756 , \2757 , \2758 , \2759 , \2760 , \2761 , \2762 , \2763 , \2764 ,
         \2765 , \2766 , \2767 , \2768 , \2769 , \2770 , \2771 , \2772 , \2773 , \2774 ,
         \2775 , \2776 , \2777 , \2778 , \2779 , \2780 , \2781 , \2782 , \2783 , \2784 ,
         \2785 , \2786 , \2787 , \2788 , \2789 , \2790 , \2791 , \2792 , \2793 , \2794 ,
         \2795 , \2796 , \2797 , \2798 , \2799 , \2800 , \2801 , \2802 , \2803 , \2804 ,
         \2805 , \2806 , \2807 , \2808 , \2809 , \2810 , \2811 , \2812 , \2813 , \2814 ,
         \2815 , \2816 , \2817 , \2818 , \2819 , \2820 , \2821 , \2822 , \2823 , \2824 ,
         \2825 , \2826 , \2827 , \2828 , \2829 , \2830 , \2831 , \2832 , \2833 , \2834 ,
         \2835 , \2836 , \2837 , \2838 , \2839 , \2840 , \2841 , \2842 , \2843 , \2844 ,
         \2845 , \2846 , \2847 , \2848 , \2849 , \2850 , \2851 , \2852 , \2853 , \2854 ,
         \2855 , \2856 , \2857 , \2858 , \2859 , \2860 , \2861 , \2862 , \2863 , \2864 ,
         \2865 , \2866 , \2867 , \2868 , \2869 , \2870 , \2871 , \2872 , \2873 , \2874 ,
         \2875 , \2876 , \2877 , \2878 , \2879 , \2880 , \2881 , \2882 , \2883 , \2884 ,
         \2885 , \2886 , \2887 , \2888 , \2889 , \2890 , \2891 , \2892 , \2893 , \2894 ,
         \2895 , \2896 , \2897 , \2898 , \2899 , \2900 , \2901 , \2902 , \2903 , \2904 ,
         \2905 , \2906 , \2907 , \2908 , \2909 , \2910 , \2911 , \2912 , \2913 , \2914 ,
         \2915 , \2916 , \2917 , \2918 , \2919 , \2920 , \2921 , \2922 , \2923 , \2924 ,
         \2925 , \2926 , \2927 , \2928 , \2929 , \2930 , \2931 , \2932 , \2933 , \2934 ,
         \2935 , \2936 , \2937 , \2938 , \2939 , \2940 , \2941 , \2942 , \2943 , \2944 ,
         \2945 , \2946 , \2947 , \2948 , \2949 , \2950 , \2951 , \2952 , \2953 , \2954 ,
         \2955 , \2956 , \2957 , \2958 , \2959 , \2960 , \2961 , \2962 , \2963 , \2964 ,
         \2965 , \2966 , \2967 , \2968 , \2969 , \2970 , \2971 , \2972 , \2973 , \2974 ,
         \2975 , \2976 , \2977 , \2978 , \2979 , \2980 , \2981 , \2982 , \2983 , \2984 ,
         \2985 , \2986 , \2987 , \2988 , \2989 , \2990 , \2991 , \2992 , \2993 , \2994 ,
         \2995 , \2996 , \2997 , \2998 , \2999 , \3000 , \3001 , \3002 , \3003 , \3004 ,
         \3005 , \3006 , \3007 , \3008 , \3009 , \3010 , \3011 , \3012 , \3013 , \3014 ,
         \3015 , \3016 , \3017 , \3018 , \3019 , \3020 , \3021 , \3022 , \3023 , \3024 ,
         \3025 , \3026 , \3027 , \3028 , \3029 , \3030 , \3031 , \3032 , \3033 , \3034 ,
         \3035 , \3036 , \3037 , \3038 , \3039 , \3040 , \3041 , \3042 , \3043 , \3044 ,
         \3045 , \3046 , \3047 , \3048 , \3049 , \3050 , \3051 , \3052 , \3053 , \3054 ,
         \3055 , \3056 , \3057 , \3058 , \3059 , \3060 , \3061 , \3062 , \3063 , \3064 ,
         \3065 , \3066 , \3067 , \3068 , \3069 , \3070 , \3071 , \3072 , \3073 , \3074 ,
         \3075 , \3076 , \3077 , \3078 , \3079 , \3080 , \3081 , \3082 , \3083 , \3084 ,
         \3085 , \3086 , \3087 , \3088 , \3089 , \3090 , \3091 , \3092 , \3093 , \3094 ,
         \3095 , \3096 , \3097 , \3098 , \3099 , \3100 , \3101 , \3102 , \3103 , \3104 ,
         \3105 , \3106 , \3107 , \3108 , \3109 , \3110 , \3111 , \3112 , \3113 , \3114 ,
         \3115 , \3116 , \3117 , \3118 , \3119 , \3120 , \3121 , \3122 , \3123 , \3124 ,
         \3125 , \3126 , \3127 , \3128 , \3129 , \3130 , \3131 , \3132 , \3133 , \3134 ,
         \3135 , \3136 , \3137 , \3138 , \3139 , \3140 , \3141 , \3142 , \3143 , \3144 ,
         \3145 , \3146 , \3147 , \3148 , \3149 , \3150 , \3151 , \3152 , \3153 , \3154 ,
         \3155 , \3156 , \3157 , \3158 , \3159 , \3160 , \3161 , \3162 , \3163 , \3164 ,
         \3165 , \3166 , \3167 , \3168 , \3169 , \3170 , \3171 , \3172 , \3173 , \3174 ,
         \3175 , \3176 , \3177 , \3178 , \3179 , \3180 , \3181 , \3182 , \3183 , \3184 ,
         \3185 , \3186 , \3187 , \3188 , \3189 , \3190 , \3191 , \3192 , \3193 , \3194 ,
         \3195 , \3196 , \3197 , \3198 , \3199 , \3200 , \3201 , \3202 , \3203 , \3204 ,
         \3205 , \3206 , \3207 , \3208 , \3209 , \3210 , \3211 , \3212 , \3213 , \3214 ,
         \3215 , \3216 , \3217 , \3218 , \3219 , \3220 , \3221 , \3222 , \3223 , \3224 ,
         \3225 , \3226 , \3227 , \3228 , \3229 , \3230 , \3231 , \3232 , \3233 , \3234 ,
         \3235 , \3236 , \3237 , \3238 , \3239 , \3240 , \3241 , \3242 , \3243 , \3244 ,
         \3245 , \3246 , \3247 , \3248 , \3249 , \3250 , \3251 , \3252 , \3253 , \3254 ,
         \3255 , \3256 , \3257 , \3258 , \3259 , \3260 , \3261 , \3262 , \3263 , \3264 ,
         \3265 , \3266 , \3267 , \3268 , \3269 , \3270 , \3271 , \3272 , \3273 , \3274 ,
         \3275 , \3276 , \3277 , \3278 , \3279 , \3280 , \3281 , \3282 , \3283 , \3284 ,
         \3285 , \3286 , \3287 , \3288 , \3289 , \3290 , \3291 , \3292 , \3293 , \3294 ,
         \3295 , \3296 , \3297 , \3298 , \3299 , \3300 , \3301 , \3302 , \3303 , \3304 ,
         \3305 , \3306 , \3307 , \3308 , \3309 , \3310 , \3311 , \3312 , \3313 , \3314 ,
         \3315 , \3316 , \3317 , \3318 , \3319 , \3320 , \3321 , \3322 , \3323 , \3324 ,
         \3325 , \3326 , \3327 , \3328 , \3329 , \3330 , \3331 , \3332 , \3333 , \3334 ,
         \3335 , \3336 , \3337 , \3338 , \3339 , \3340 , \3341 , \3342 , \3343 , \3344 ,
         \3345 , \3346 , \3347 , \3348 , \3349 , \3350 , \3351 , \3352 , \3353 , \3354 ,
         \3355 , \3356 , \3357 , \3358 , \3359 , \3360 , \3361 , \3362 , \3363 , \3364 ,
         \3365 , \3366 , \3367 , \3368 , \3369 , \3370 , \3371 , \3372 , \3373 , \3374 ,
         \3375 , \3376 , \3377 , \3378 , \3379 , \3380 , \3381 , \3382 , \3383 , \3384 ,
         \3385 , \3386 , \3387 , \3388 , \3389 , \3390 , \3391 , \3392 , \3393 , \3394 ,
         \3395 , \3396 , \3397 , \3398 , \3399 , \3400 , \3401 , \3402 , \3403 , \3404 ,
         \3405 , \3406 , \3407 , \3408 , \3409 , \3410 , \3411 , \3412 , \3413 , \3414 ,
         \3415 , \3416 , \3417 , \3418 , \3419 , \3420 , \3421 , \3422 , \3423 , \3424 ,
         \3425 , \3426 , \3427 , \3428 , \3429 , \3430 , \3431 , \3432 , \3433 , \3434 ,
         \3435 , \3436 , \3437 , \3438 , \3439 , \3440 , \3441 , \3442 , \3443 , \3444 ,
         \3445 , \3446 , \3447 , \3448 , \3449 , \3450 , \3451 , \3452 , \3453 , \3454 ,
         \3455 , \3456 , \3457 , \3458 , \3459 , \3460 , \3461 , \3462 , \3463 , \3464 ,
         \3465 , \3466 , \3467 , \3468 , \3469 , \3470 , \3471 , \3472 , \3473 , \3474 ,
         \3475 , \3476 , \3477 , \3478 , \3479 , \3480 , \3481 , \3482 , \3483 , \3484 ,
         \3485 , \3486 , \3487 , \3488 , \3489 , \3490 , \3491 , \3492 , \3493 , \3494 ,
         \3495 , \3496 , \3497 , \3498 , \3499 , \3500 , \3501 , \3502 , \3503 , \3504 ,
         \3505 , \3506 , \3507 , \3508 , \3509 , \3510 , \3511 , \3512 , \3513 , \3514 ,
         \3515 , \3516 , \3517 , \3518 , \3519 , \3520 , \3521 , \3522 , \3523 , \3524 ,
         \3525 , \3526 , \3527 , \3528 , \3529 , \3530 , \3531 , \3532 , \3533 , \3534 ,
         \3535 , \3536 , \3537 , \3538 , \3539 , \3540 , \3541 , \3542 , \3543 , \3544 ,
         \3545 , \3546 , \3547 , \3548 , \3549 , \3550 , \3551 , \3552 , \3553 , \3554 ,
         \3555 , \3556 , \3557 , \3558 , \3559 , \3560 , \3561 , \3562 , \3563 , \3564 ,
         \3565 , \3566 , \3567 , \3568 , \3569 , \3570 , \3571 , \3572 , \3573 , \3574 ,
         \3575 , \3576 , \3577 , \3578 , \3579 , \3580 , \3581 , \3582 , \3583 , \3584 ,
         \3585 , \3586 , \3587 , \3588 , \3589 , \3590 , \3591 , \3592 , \3593 , \3594 ,
         \3595 , \3596 , \3597 , \3598 , \3599 , \3600 , \3601 , \3602 , \3603 , \3604 ,
         \3605 , \3606 , \3607 , \3608 , \3609 , \3610 , \3611 , \3612 , \3613 , \3614 ,
         \3615 , \3616 , \3617 , \3618 , \3619 , \3620 , \3621 , \3622 , \3623 , \3624 ,
         \3625 , \3626 , \3627 , \3628 , \3629 , \3630 , \3631 , \3632 , \3633 , \3634 ,
         \3635 , \3636 , \3637 , \3638 , \3639 , \3640 , \3641 , \3642 , \3643 , \3644 ,
         \3645 , \3646 , \3647 , \3648 , \3649 , \3650 , \3651 , \3652 , \3653 , \3654 ,
         \3655 , \3656 , \3657 , \3658 , \3659 , \3660 , \3661 , \3662 , \3663 , \3664 ,
         \3665 , \3666 , \3667 , \3668 , \3669 , \3670 , \3671 , \3672 , \3673 , \3674 ,
         \3675 , \3676 , \3677 , \3678 , \3679 , \3680 , \3681 , \3682 , \3683 , \3684 ,
         \3685 , \3686 , \3687 , \3688 , \3689 , \3690 , \3691 , \3692 , \3693 , \3694 ,
         \3695 , \3696 , \3697 , \3698 , \3699 , \3700 , \3701 , \3702 , \3703 , \3704 ,
         \3705 , \3706 , \3707 , \3708 , \3709 , \3710 , \3711 , \3712 , \3713 , \3714 ,
         \3715 , \3716 , \3717 , \3718 , \3719 , \3720 , \3721 , \3722 , \3723 , \3724 ,
         \3725 , \3726 , \3727 , \3728 , \3729 , \3730 , \3731 , \3732 , \3733 , \3734 ,
         \3735 , \3736 , \3737 , \3738 , \3739 , \3740 , \3741 , \3742 , \3743 , \3744 ,
         \3745 , \3746 , \3747 , \3748 , \3749 , \3750 , \3751 , \3752 , \3753 , \3754 ,
         \3755 , \3756 , \3757 , \3758 , \3759 , \3760 , \3761 , \3762 , \3763 , \3764 ,
         \3765 , \3766 , \3767 , \3768 , \3769 , \3770 , \3771 , \3772 , \3773 , \3774 ,
         \3775 , \3776 , \3777 , \3778 , \3779 , \3780 , \3781 , \3782 , \3783 , \3784 ,
         \3785 , \3786 , \3787 , \3788 , \3789 , \3790 , \3791 , \3792 , \3793 , \3794 ,
         \3795 , \3796 , \3797 , \3798 , \3799 , \3800 , \3801 , \3802 , \3803 , \3804 ,
         \3805 , \3806 , \3807 , \3808 , \3809 , \3810 , \3811 , \3812 , \3813 , \3814 ,
         \3815 , \3816 , \3817 , \3818 , \3819 , \3820 , \3821 , \3822 , \3823 , \3824 ,
         \3825 , \3826 , \3827 , \3828 , \3829 , \3830 , \3831 , \3832 , \3833 , \3834 ,
         \3835 , \3836 , \3837 , \3838 , \3839 , \3840 , \3841 , \3842 , \3843 , \3844 ,
         \3845 , \3846 , \3847 , \3848 , \3849 , \3850 , \3851 , \3852 , \3853 , \3854 ,
         \3855 , \3856 , \3857 , \3858 , \3859 , \3860 , \3861 , \3862 , \3863 , \3864 ,
         \3865 , \3866 , \3867 , \3868 , \3869 , \3870 , \3871 , \3872 , \3873 , \3874 ,
         \3875 , \3876 , \3877 , \3878 , \3879 , \3880 , \3881 , \3882 , \3883 , \3884 ,
         \3885 , \3886 , \3887 , \3888 , \3889 , \3890 , \3891 , \3892 , \3893 , \3894 ,
         \3895 , \3896 , \3897 , \3898 , \3899 , \3900 , \3901 , \3902 , \3903 , \3904 ,
         \3905 , \3906 , \3907 , \3908 , \3909 , \3910 , \3911 , \3912 , \3913 , \3914 ,
         \3915 , \3916 , \3917 , \3918 , \3919 , \3920 , \3921 , \3922 , \3923 , \3924 ,
         \3925 , \3926 , \3927 , \3928 , \3929 , \3930 , \3931 , \3932 , \3933 , \3934 ,
         \3935 , \3936 , \3937 , \3938 , \3939 , \3940 , \3941 , \3942 , \3943 , \3944 ,
         \3945 , \3946 , \3947 , \3948 , \3949 , \3950 , \3951 , \3952 , \3953 , \3954 ,
         \3955 , \3956 , \3957 , \3958 , \3959 , \3960 , \3961 , \3962 , \3963 , \3964 ,
         \3965 , \3966 , \3967 , \3968 , \3969 , \3970 , \3971 , \3972 , \3973 , \3974 ,
         \3975 , \3976 , \3977 , \3978 , \3979 , \3980 , \3981 , \3982 , \3983 , \3984 ,
         \3985 , \3986 , \3987 , \3988 , \3989 , \3990 , \3991 , \3992 , \3993 , \3994 ,
         \3995 , \3996 , \3997 , \3998 , \3999 , \4000 , \4001 , \4002 , \4003 , \4004 ,
         \4005 , \4006 , \4007 , \4008 , \4009 , \4010 , \4011 , \4012 , \4013 , \4014 ,
         \4015 , \4016 , \4017 , \4018 , \4019 , \4020 , \4021 , \4022 , \4023 , \4024 ,
         \4025 , \4026 , \4027 , \4028 , \4029 , \4030 , \4031 , \4032 , \4033 , \4034 ,
         \4035 , \4036 , \4037 , \4038 , \4039 , \4040 , \4041 , \4042 , \4043 , \4044 ,
         \4045 , \4046 , \4047 , \4048 , \4049 , \4050 , \4051 , \4052 , \4053 , \4054 ,
         \4055 , \4056 , \4057 , \4058 , \4059 , \4060 , \4061 , \4062 , \4063 , \4064 ,
         \4065 , \4066 , \4067 , \4068 , \4069 , \4070 , \4071 , \4072 , \4073 , \4074 ,
         \4075 , \4076 , \4077 , \4078 , \4079 , \4080 , \4081 , \4082 , \4083 , \4084 ,
         \4085 , \4086 , \4087 , \4088 , \4089 , \4090 , \4091 , \4092 , \4093 , \4094 ,
         \4095 , \4096 , \4097 , \4098 , \4099 , \4100 , \4101 , \4102 , \4103 , \4104 ,
         \4105 , \4106 , \4107 , \4108 , \4109 , \4110 , \4111 , \4112 , \4113 , \4114 ,
         \4115 , \4116 , \4117 , \4118 , \4119 , \4120 , \4121 , \4122 , \4123 , \4124 ,
         \4125 , \4126 , \4127 , \4128 , \4129 , \4130 , \4131 , \4132 , \4133 , \4134 ,
         \4135 , \4136 , \4137 , \4138 , \4139 , \4140 , \4141 , \4142 , \4143 , \4144 ,
         \4145 , \4146 , \4147 , \4148 , \4149 , \4150 , \4151 , \4152 , \4153 , \4154 ,
         \4155 , \4156 , \4157 , \4158 , \4159 , \4160 , \4161 , \4162 , \4163 , \4164 ,
         \4165 , \4166 , \4167 , \4168 , \4169 , \4170 , \4171 , \4172 , \4173 , \4174 ,
         \4175 , \4176 , \4177 , \4178 , \4179 , \4180 , \4181 , \4182 , \4183 , \4184 ,
         \4185 , \4186 , \4187 , \4188 , \4189 , \4190 , \4191 , \4192 , \4193 , \4194 ,
         \4195 , \4196 , \4197 , \4198 , \4199 , \4200 , \4201 , \4202 , \4203 , \4204 ,
         \4205 , \4206 , \4207 , \4208 , \4209 , \4210 , \4211 , \4212 , \4213 , \4214 ,
         \4215 , \4216 , \4217 , \4218 , \4219 , \4220 , \4221 , \4222 , \4223 , \4224 ,
         \4225 , \4226 , \4227 , \4228 , \4229 , \4230 , \4231 , \4232 , \4233 , \4234 ,
         \4235 , \4236 , \4237 , \4238 , \4239 , \4240 , \4241 , \4242 , \4243 , \4244 ,
         \4245 , \4246 , \4247 , \4248 , \4249 , \4250 , \4251 , \4252 , \4253 , \4254 ,
         \4255 , \4256 , \4257 , \4258 , \4259 , \4260 , \4261 , \4262 , \4263 , \4264 ,
         \4265 , \4266 , \4267 , \4268 , \4269 , \4270 , \4271 , \4272 , \4273 , \4274 ,
         \4275 , \4276 , \4277 , \4278 , \4279 , \4280 , \4281 , \4282 , \4283 , \4284 ,
         \4285 , \4286 , \4287 , \4288 , \4289 , \4290 , \4291 , \4292 , \4293 , \4294 ,
         \4295 , \4296 , \4297 , \4298 , \4299 , \4300 , \4301 , \4302 , \4303 , \4304 ,
         \4305 , \4306 , \4307 , \4308 , \4309 , \4310 , \4311 , \4312 , \4313 , \4314 ,
         \4315 , \4316 , \4317 , \4318 , \4319 , \4320 , \4321 , \4322 , \4323 , \4324 ,
         \4325 , \4326 , \4327 , \4328 , \4329 , \4330 , \4331 , \4332 , \4333 , \4334 ,
         \4335 , \4336 , \4337 , \4338 , \4339 , \4340 , \4341 , \4342 , \4343 , \4344 ,
         \4345 , \4346 , \4347 , \4348 , \4349 , \4350 , \4351 , \4352 , \4353 , \4354 ,
         \4355 , \4356 , \4357 , \4358 , \4359 , \4360 , \4361 , \4362 , \4363 , \4364 ,
         \4365 , \4366 , \4367 , \4368 , \4369 , \4370 , \4371 , \4372 , \4373 , \4374 ,
         \4375 , \4376 , \4377 , \4378 , \4379 , \4380 , \4381 , \4382 , \4383 , \4384 ,
         \4385 , \4386 , \4387 , \4388 , \4389 , \4390 , \4391 , \4392 , \4393 , \4394 ,
         \4395 , \4396 , \4397 , \4398 , \4399 , \4400 , \4401 , \4402 , \4403 , \4404 ,
         \4405 , \4406 , \4407 , \4408 , \4409 , \4410 , \4411 , \4412 , \4413 , \4414 ,
         \4415 , \4416 , \4417 , \4418 , \4419 , \4420 , \4421 , \4422 , \4423 , \4424 ,
         \4425 , \4426 , \4427 , \4428 , \4429 , \4430 , \4431 , \4432 , \4433 , \4434 ,
         \4435 , \4436 , \4437 , \4438 , \4439 , \4440 , \4441 , \4442 , \4443 , \4444 ,
         \4445 , \4446 , \4447 , \4448 , \4449 , \4450 , \4451 , \4452 , \4453 , \4454 ,
         \4455 , \4456 , \4457 , \4458 , \4459 , \4460 , \4461 , \4462 , \4463 , \4464 ,
         \4465 , \4466 , \4467 , \4468 , \4469 , \4470 , \4471 , \4472 , \4473 , \4474 ,
         \4475 , \4476 , \4477 , \4478 , \4479 , \4480 , \4481 , \4482 , \4483 , \4484 ,
         \4485 , \4486 , \4487 , \4488 , \4489 , \4490 , \4491 , \4492 , \4493 , \4494 ,
         \4495 , \4496 , \4497 , \4498 , \4499 , \4500 , \4501 , \4502 , \4503 , \4504 ,
         \4505 , \4506 , \4507 , \4508 , \4509 , \4510 , \4511 , \4512 , \4513 , \4514 ,
         \4515 , \4516 , \4517 , \4518 , \4519 , \4520 , \4521 , \4522 , \4523 , \4524 ,
         \4525 , \4526 , \4527 , \4528 , \4529 , \4530 , \4531 , \4532 , \4533 , \4534 ,
         \4535 , \4536 , \4537 , \4538 , \4539 , \4540 , \4541 , \4542 , \4543 , \4544 ,
         \4545 , \4546 , \4547 , \4548 , \4549 , \4550 , \4551 , \4552 , \4553 , \4554 ,
         \4555 , \4556 , \4557 , \4558 , \4559 , \4560 , \4561 , \4562 , \4563 , \4564 ,
         \4565 , \4566 , \4567 , \4568 , \4569 , \4570 , \4571 , \4572 , \4573 , \4574 ,
         \4575 , \4576 , \4577 , \4578 , \4579 , \4580 , \4581 , \4582 , \4583 , \4584 ,
         \4585 , \4586 , \4587 , \4588 , \4589 , \4590 , \4591 , \4592 , \4593 , \4594 ,
         \4595 , \4596 , \4597 , \4598 , \4599 , \4600 , \4601 , \4602 , \4603 , \4604 ,
         \4605 , \4606 , \4607 , \4608 , \4609 , \4610 , \4611 , \4612 , \4613 , \4614 ,
         \4615 , \4616 , \4617 , \4618 , \4619 , \4620 , \4621 , \4622 , \4623 , \4624 ,
         \4625 , \4626 , \4627 , \4628 , \4629 , \4630 , \4631 , \4632 , \4633 , \4634 ,
         \4635 , \4636 , \4637 , \4638 , \4639 , \4640 , \4641 , \4642 , \4643 , \4644 ,
         \4645 , \4646 , \4647 , \4648 , \4649 , \4650 , \4651 , \4652 , \4653 , \4654 ,
         \4655 , \4656 , \4657 , \4658 , \4659 , \4660 , \4661 , \4662 , \4663 , \4664 ,
         \4665 , \4666 , \4667 , \4668 , \4669 , \4670 , \4671 , \4672 , \4673 , \4674 ,
         \4675 , \4676 , \4677 , \4678 , \4679 , \4680 , \4681 , \4682 , \4683 , \4684 ,
         \4685 , \4686 , \4687 , \4688 , \4689 , \4690 , \4691 , \4692 , \4693 , \4694 ,
         \4695 , \4696 , \4697 , \4698 , \4699 , \4700 , \4701 , \4702 , \4703 , \4704 ,
         \4705 , \4706 , \4707 , \4708 , \4709 , \4710 , \4711 , \4712 , \4713 , \4714 ,
         \4715 , \4716 , \4717 , \4718 , \4719 , \4720 , \4721 , \4722 , \4723 , \4724 ,
         \4725 , \4726 , \4727 , \4728 , \4729 , \4730 , \4731 , \4732 , \4733 , \4734 ,
         \4735 , \4736 , \4737 , \4738 , \4739 , \4740 , \4741 , \4742 , \4743 , \4744 ,
         \4745 , \4746 , \4747 , \4748 , \4749 , \4750 , \4751 , \4752 , \4753 , \4754 ,
         \4755 , \4756 , \4757 , \4758 , \4759 , \4760 , \4761 , \4762 , \4763 , \4764 ,
         \4765 , \4766 , \4767 , \4768 , \4769 , \4770 , \4771 , \4772 , \4773 , \4774 ,
         \4775 , \4776 , \4777 , \4778 , \4779 , \4780 , \4781 , \4782 , \4783 , \4784 ,
         \4785 , \4786 , \4787 , \4788 , \4789 , \4790 , \4791 , \4792 , \4793 , \4794 ,
         \4795 , \4796 , \4797 , \4798 , \4799 , \4800 , \4801 , \4802 , \4803 , \4804 ,
         \4805 , \4806 , \4807 , \4808 , \4809 , \4810 , \4811 , \4812 , \4813 , \4814 ,
         \4815 , \4816 , \4817 , \4818 , \4819 , \4820 , \4821 , \4822 , \4823 , \4824 ,
         \4825 , \4826 , \4827 , \4828 , \4829 , \4830 , \4831 , \4832 , \4833 , \4834 ,
         \4835 , \4836 , \4837 , \4838 , \4839 , \4840 , \4841 , \4842 , \4843 , \4844 ,
         \4845 , \4846 , \4847 , \4848 , \4849 , \4850 , \4851 , \4852 , \4853 , \4854 ,
         \4855 , \4856 , \4857 , \4858 , \4859 , \4860 , \4861 , \4862 , \4863 , \4864 ,
         \4865 , \4866 , \4867 , \4868 , \4869 , \4870 , \4871 , \4872 , \4873 , \4874 ,
         \4875 , \4876 , \4877 , \4878 , \4879 , \4880 , \4881 , \4882 , \4883 , \4884 ,
         \4885 , \4886 , \4887 , \4888 , \4889 , \4890 , \4891 , \4892 , \4893 , \4894 ,
         \4895 , \4896 , \4897 , \4898 , \4899 , \4900 , \4901 , \4902 , \4903 , \4904 ,
         \4905 , \4906 , \4907 , \4908 , \4909 , \4910 , \4911 , \4912 , \4913 , \4914 ,
         \4915 , \4916 , \4917 , \4918 , \4919 , \4920 , \4921 , \4922 , \4923 , \4924 ,
         \4925 , \4926 , \4927 , \4928 , \4929 , \4930 , \4931 , \4932 , \4933 , \4934 ,
         \4935 , \4936 , \4937 , \4938 , \4939 , \4940 , \4941 , \4942 , \4943 , \4944 ,
         \4945 , \4946 , \4947 , \4948 , \4949 , \4950 , \4951 , \4952 , \4953 , \4954 ,
         \4955 , \4956 , \4957 , \4958 , \4959 , \4960 , \4961 , \4962 , \4963 , \4964 ,
         \4965 , \4966 , \4967 , \4968 , \4969 , \4970 , \4971 , \4972 , \4973 , \4974 ,
         \4975 , \4976 , \4977 , \4978 , \4979 , \4980 , \4981 , \4982 , \4983 , \4984 ,
         \4985 , \4986 , \4987 , \4988 , \4989 , \4990 , \4991 , \4992 , \4993 , \4994 ,
         \4995 , \4996 , \4997 , \4998 , \4999 , \5000 , \5001 , \5002 , \5003 , \5004 ,
         \5005 , \5006 , \5007 , \5008 , \5009 , \5010 , \5011 , \5012 , \5013 , \5014 ,
         \5015 , \5016 , \5017 , \5018 , \5019 , \5020 , \5021 , \5022 , \5023 , \5024 ,
         \5025 , \5026 , \5027 , \5028 , \5029 , \5030 , \5031 , \5032 , \5033 , \5034 ,
         \5035 , \5036 , \5037 , \5038 , \5039 , \5040 , \5041 , \5042 , \5043 , \5044 ,
         \5045 , \5046 , \5047 , \5048 , \5049 , \5050 , \5051 , \5052 , \5053 , \5054 ,
         \5055 , \5056 , \5057 , \5058 , \5059 , \5060 , \5061 , \5062 , \5063 , \5064 ,
         \5065 , \5066 , \5067 , \5068 , \5069 , \5070 , \5071 , \5072 , \5073 , \5074 ,
         \5075 , \5076 , \5077 , \5078 , \5079 , \5080 , \5081 , \5082 , \5083 , \5084 ,
         \5085 , \5086 , \5087 , \5088 , \5089 , \5090 , \5091 , \5092 , \5093 , \5094 ,
         \5095 , \5096 , \5097 , \5098 , \5099 , \5100 , \5101 , \5102 , \5103 , \5104 ,
         \5105 , \5106 , \5107 , \5108 , \5109 , \5110 , \5111 , \5112 , \5113 , \5114 ,
         \5115 , \5116 , \5117 , \5118 , \5119 , \5120 , \5121 , \5122 , \5123 , \5124 ,
         \5125 , \5126 , \5127 , \5128 , \5129 , \5130 , \5131 , \5132 , \5133 , \5134 ,
         \5135 , \5136 , \5137 , \5138 , \5139 , \5140 , \5141 , \5142 , \5143 , \5144 ,
         \5145 , \5146 , \5147 , \5148 , \5149 , \5150 , \5151 , \5152 , \5153 , \5154 ,
         \5155 , \5156 , \5157 , \5158 , \5159 , \5160 , \5161 , \5162 , \5163 , \5164 ,
         \5165 , \5166 , \5167 , \5168 , \5169 , \5170 , \5171 , \5172 , \5173 , \5174 ,
         \5175 , \5176 , \5177 , \5178 , \5179 , \5180 , \5181 , \5182 , \5183 , \5184 ,
         \5185 , \5186 , \5187 , \5188 , \5189 , \5190 , \5191 , \5192 , \5193 , \5194 ,
         \5195 , \5196 , \5197 , \5198 , \5199 , \5200 , \5201 , \5202 , \5203 , \5204 ,
         \5205 , \5206 , \5207 , \5208 , \5209 , \5210 , \5211 , \5212 , \5213 , \5214 ,
         \5215 , \5216 , \5217 , \5218 , \5219 , \5220 , \5221 , \5222 , \5223 , \5224 ,
         \5225 , \5226 , \5227 , \5228 , \5229 , \5230 , \5231 , \5232 , \5233 , \5234 ,
         \5235 , \5236 , \5237 , \5238 , \5239 , \5240 , \5241 , \5242 , \5243 , \5244 ,
         \5245 , \5246 , \5247 , \5248 , \5249 , \5250 , \5251 , \5252 , \5253 , \5254 ,
         \5255 , \5256 , \5257 , \5258 , \5259 , \5260 , \5261 , \5262 , \5263 , \5264 ,
         \5265 , \5266 , \5267 , \5268 , \5269 , \5270 , \5271 , \5272 , \5273 , \5274 ,
         \5275 , \5276 , \5277 , \5278 , \5279 , \5280 , \5281 , \5282 , \5283 , \5284 ,
         \5285 , \5286 , \5287 , \5288 , \5289 , \5290 , \5291 , \5292 , \5293 , \5294 ,
         \5295 , \5296 , \5297 , \5298 , \5299 , \5300 , \5301 , \5302 , \5303 , \5304 ,
         \5305 , \5306 , \5307 , \5308 , \5309 , \5310 , \5311 , \5312 , \5313 , \5314 ,
         \5315 , \5316 , \5317 , \5318 , \5319 , \5320 , \5321 , \5322 , \5323 , \5324 ,
         \5325 , \5326 , \5327 , \5328 , \5329 , \5330 , \5331 , \5332 , \5333 , \5334 ,
         \5335 , \5336 , \5337 , \5338 , \5339 , \5340 , \5341 , \5342 , \5343 , \5344 ,
         \5345 , \5346 , \5347 , \5348 , \5349 , \5350 , \5351 , \5352 , \5353 , \5354 ,
         \5355 , \5356 , \5357 , \5358 , \5359 , \5360 , \5361 , \5362 , \5363 , \5364 ,
         \5365 , \5366 , \5367 , \5368 , \5369 , \5370 , \5371 , \5372 , \5373 , \5374 ,
         \5375 , \5376 , \5377 , \5378 , \5379 , \5380 , \5381 , \5382 , \5383 , \5384 ,
         \5385 , \5386 , \5387 , \5388 , \5389 , \5390 , \5391 , \5392 , \5393 , \5394 ,
         \5395 , \5396 , \5397 , \5398 , \5399 , \5400 , \5401 , \5402 , \5403 , \5404 ,
         \5405 , \5406 , \5407 , \5408 , \5409 , \5410 , \5411 , \5412 , \5413 , \5414 ,
         \5415 , \5416 , \5417 , \5418 , \5419 , \5420 , \5421 , \5422 , \5423 , \5424 ,
         \5425 , \5426 , \5427 , \5428 , \5429 , \5430 , \5431 , \5432 , \5433 , \5434 ,
         \5435 , \5436 , \5437 , \5438 , \5439 , \5440 , \5441 , \5442 , \5443 , \5444 ,
         \5445 , \5446 , \5447 , \5448 , \5449 , \5450 , \5451 , \5452 , \5453 , \5454 ,
         \5455 , \5456 , \5457 , \5458 , \5459 , \5460 , \5461 , \5462 , \5463 , \5464 ,
         \5465 , \5466 , \5467 , \5468 , \5469 , \5470 , \5471 , \5472 , \5473 , \5474 ,
         \5475 , \5476 , \5477 , \5478 , \5479 , \5480 , \5481 , \5482 , \5483 , \5484 ,
         \5485 , \5486 , \5487 , \5488 , \5489 , \5490 , \5491 , \5492 , \5493 , \5494 ,
         \5495 , \5496 , \5497 , \5498 , \5499 , \5500 , \5501 , \5502 , \5503 , \5504 ,
         \5505 , \5506 , \5507 , \5508 , \5509 , \5510 , \5511 , \5512 , \5513 , \5514 ,
         \5515 , \5516 , \5517 , \5518 , \5519 , \5520 , \5521 , \5522 , \5523 , \5524 ,
         \5525 , \5526 , \5527 , \5528 , \5529 , \5530 , \5531 , \5532 , \5533 , \5534 ,
         \5535 , \5536 , \5537 , \5538 , \5539 , \5540 , \5541 , \5542 , \5543 , \5544 ,
         \5545 , \5546 , \5547 , \5548 , \5549 , \5550 , \5551 , \5552 , \5553 , \5554 ,
         \5555 , \5556 , \5557 , \5558 , \5559 , \5560 , \5561 , \5562 , \5563 , \5564 ,
         \5565 , \5566 , \5567 , \5568 , \5569 , \5570 , \5571 , \5572 , \5573 , \5574 ,
         \5575 , \5576 , \5577 , \5578 , \5579 , \5580 , \5581 , \5582 , \5583 , \5584 ,
         \5585 , \5586 , \5587 , \5588 , \5589 , \5590 , \5591 , \5592 , \5593 , \5594 ,
         \5595 , \5596 , \5597 , \5598 , \5599 , \5600 , \5601 , \5602 , \5603 , \5604 ,
         \5605 , \5606 , \5607 , \5608 , \5609 , \5610 , \5611 , \5612 , \5613 , \5614 ,
         \5615 , \5616 , \5617 , \5618 , \5619 , \5620 , \5621 , \5622 , \5623 , \5624 ,
         \5625 , \5626 , \5627 , \5628 , \5629 , \5630 , \5631 , \5632 , \5633 , \5634 ,
         \5635 , \5636 , \5637 , \5638 , \5639 , \5640 , \5641 , \5642 , \5643 , \5644 ,
         \5645 , \5646 , \5647 , \5648 , \5649 , \5650 , \5651 , \5652 , \5653 , \5654 ,
         \5655 , \5656 , \5657 , \5658 , \5659 , \5660 , \5661 , \5662 , \5663 , \5664 ,
         \5665 , \5666 , \5667 , \5668 , \5669 , \5670 , \5671 , \5672 , \5673 , \5674 ,
         \5675 , \5676 , \5677 , \5678 , \5679 , \5680 , \5681 , \5682 , \5683 , \5684 ,
         \5685 , \5686 , \5687 , \5688 , \5689 , \5690 , \5691 , \5692 , \5693 , \5694 ,
         \5695 , \5696 , \5697 , \5698 , \5699 , \5700 , \5701 , \5702 , \5703 , \5704 ,
         \5705 , \5706 , \5707 , \5708 , \5709 , \5710 , \5711 , \5712 , \5713 , \5714 ,
         \5715 , \5716 , \5717 , \5718 , \5719 , \5720 , \5721 , \5722 , \5723 , \5724 ,
         \5725 , \5726 , \5727 , \5728 , \5729 , \5730 , \5731 , \5732 , \5733 , \5734 ,
         \5735 , \5736 , \5737 , \5738 , \5739 , \5740 , \5741 , \5742 , \5743 , \5744 ,
         \5745 , \5746 , \5747 , \5748 , \5749 , \5750 , \5751 , \5752 , \5753 , \5754 ,
         \5755 , \5756 , \5757 , \5758 , \5759 , \5760 , \5761 , \5762 , \5763 , \5764 ,
         \5765 , \5766 , \5767 , \5768 , \5769 , \5770 , \5771 , \5772 , \5773 , \5774 ,
         \5775 , \5776 , \5777 , \5778 , \5779 , \5780 , \5781 , \5782 , \5783 , \5784 ,
         \5785 , \5786 , \5787 , \5788 , \5789 , \5790 , \5791 , \5792 , \5793 , \5794 ,
         \5795 , \5796 , \5797 , \5798 , \5799 , \5800 , \5801 , \5802 , \5803 , \5804 ,
         \5805 , \5806 , \5807 , \5808 , \5809 , \5810 , \5811 , \5812 , \5813 , \5814 ,
         \5815 , \5816 , \5817 , \5818 , \5819 , \5820 , \5821 , \5822 , \5823 , \5824 ,
         \5825 , \5826 , \5827 , \5828 , \5829 , \5830 , \5831 , \5832 , \5833 , \5834 ,
         \5835 , \5836 , \5837 , \5838 , \5839 , \5840 , \5841 , \5842 , \5843 , \5844 ,
         \5845 , \5846 , \5847 , \5848 , \5849 , \5850 , \5851 , \5852 , \5853 , \5854 ,
         \5855 , \5856 , \5857 , \5858 , \5859 , \5860 , \5861 , \5862 , \5863 , \5864 ,
         \5865 , \5866 , \5867 , \5868 , \5869 , \5870 , \5871 , \5872 , \5873 , \5874 ,
         \5875 , \5876 , \5877 , \5878 , \5879 , \5880 , \5881 , \5882 , \5883 , \5884 ,
         \5885 , \5886 , \5887 , \5888 , \5889 , \5890 , \5891 , \5892 , \5893 , \5894 ,
         \5895 , \5896 , \5897 , \5898 , \5899 , \5900 , \5901 , \5902 , \5903 , \5904 ,
         \5905 , \5906 , \5907 , \5908 , \5909 , \5910 , \5911 , \5912 , \5913 , \5914 ,
         \5915 , \5916 , \5917 , \5918 , \5919 , \5920 , \5921 , \5922 , \5923 , \5924 ,
         \5925 , \5926 , \5927 , \5928 , \5929 , \5930 , \5931 , \5932 , \5933 , \5934 ,
         \5935 , \5936 , \5937 , \5938 , \5939 , \5940 , \5941 , \5942 , \5943 , \5944 ,
         \5945 , \5946 , \5947 , \5948 , \5949 , \5950 , \5951 , \5952 , \5953 , \5954 ,
         \5955 , \5956 , \5957 , \5958 , \5959 , \5960 , \5961 , \5962 , \5963 , \5964 ,
         \5965 , \5966 , \5967 , \5968 , \5969 , \5970 , \5971 , \5972 , \5973 , \5974 ,
         \5975 , \5976 , \5977 , \5978 , \5979 , \5980 , \5981 , \5982 , \5983 , \5984 ,
         \5985 , \5986 , \5987 , \5988 , \5989 , \5990 , \5991 , \5992 , \5993 , \5994 ,
         \5995 , \5996 , \5997 , \5998 , \5999 , \6000 , \6001 , \6002 , \6003 , \6004 ,
         \6005 , \6006 , \6007 , \6008 , \6009 , \6010 , \6011 , \6012 , \6013 , \6014 ,
         \6015 , \6016 , \6017 , \6018 , \6019 , \6020 , \6021 , \6022 , \6023 , \6024 ,
         \6025 , \6026 , \6027 , \6028 , \6029 , \6030 , \6031 , \6032 , \6033 , \6034 ,
         \6035 , \6036 , \6037 , \6038 , \6039 , \6040 , \6041 , \6042 , \6043 , \6044 ,
         \6045 , \6046 , \6047 , \6048 , \6049 , \6050 , \6051 , \6052 , \6053 , \6054 ,
         \6055 , \6056 , \6057 , \6058 , \6059 , \6060 , \6061 , \6062 , \6063 , \6064 ,
         \6065 , \6066 , \6067 , \6068 , \6069 , \6070 , \6071 , \6072 , \6073 , \6074 ,
         \6075 , \6076 , \6077 , \6078 , \6079 , \6080 , \6081 , \6082 , \6083 , \6084 ,
         \6085 , \6086 , \6087 , \6088 , \6089 , \6090 , \6091 , \6092 , \6093 , \6094 ,
         \6095 , \6096 , \6097 , \6098 , \6099 , \6100 , \6101 , \6102 , \6103 , \6104 ,
         \6105 , \6106 , \6107 , \6108 , \6109 , \6110 , \6111 , \6112 , \6113 , \6114 ,
         \6115 , \6116 , \6117 , \6118 , \6119 , \6120 , \6121 , \6122 , \6123 , \6124 ,
         \6125 , \6126 , \6127 , \6128 , \6129 , \6130 , \6131 , \6132 , \6133 , \6134 ,
         \6135 , \6136 , \6137 , \6138 , \6139 , \6140 , \6141 , \6142 , \6143 , \6144 ,
         \6145 , \6146 , \6147 , \6148 , \6149 , \6150 , \6151 , \6152 , \6153 , \6154 ,
         \6155 , \6156 , \6157 , \6158 , \6159 , \6160 , \6161 , \6162 , \6163 , \6164 ,
         \6165 , \6166 , \6167 , \6168 , \6169 , \6170 , \6171 , \6172 , \6173 , \6174 ,
         \6175 , \6176 , \6177 , \6178 , \6179 , \6180 , \6181 , \6182 , \6183 , \6184 ,
         \6185 , \6186 , \6187 , \6188 , \6189 , \6190 , \6191 , \6192 , \6193 , \6194 ,
         \6195 , \6196 , \6197 , \6198 , \6199 , \6200 , \6201 , \6202 , \6203 , \6204 ,
         \6205 , \6206 , \6207 , \6208 , \6209 , \6210 , \6211 , \6212 , \6213 , \6214 ,
         \6215 , \6216 , \6217 , \6218 , \6219 , \6220 , \6221 , \6222 , \6223 , \6224 ,
         \6225 , \6226 , \6227 , \6228 , \6229 , \6230 , \6231 , \6232 , \6233 , \6234 ,
         \6235 , \6236 , \6237 , \6238 , \6239 , \6240 , \6241 , \6242 , \6243 , \6244 ,
         \6245 , \6246 , \6247 , \6248 , \6249 , \6250 , \6251 , \6252 , \6253 , \6254 ,
         \6255 , \6256 , \6257 , \6258 , \6259 , \6260 , \6261 , \6262 , \6263 , \6264 ,
         \6265 , \6266 , \6267 , \6268 , \6269 , \6270 , \6271 , \6272 , \6273 , \6274 ,
         \6275 , \6276 , \6277 , \6278 , \6279 , \6280 , \6281 , \6282 , \6283 , \6284 ,
         \6285 , \6286 , \6287 , \6288 , \6289 , \6290 , \6291 , \6292 , \6293 , \6294 ,
         \6295 , \6296 , \6297 , \6298 , \6299 , \6300 , \6301 , \6302 , \6303 , \6304 ,
         \6305 , \6306 , \6307 , \6308 , \6309 , \6310 , \6311 , \6312 , \6313 , \6314 ,
         \6315 , \6316 , \6317 , \6318 , \6319 , \6320 , \6321 , \6322 , \6323 , \6324 ,
         \6325 , \6326 , \6327 , \6328 , \6329 , \6330 , \6331 , \6332 , \6333 , \6334 ,
         \6335 , \6336 , \6337 , \6338 , \6339 , \6340 , \6341 , \6342 , \6343 , \6344 ,
         \6345 , \6346 , \6347 , \6348 , \6349 , \6350 , \6351 , \6352 , \6353 , \6354 ,
         \6355 , \6356 , \6357 , \6358 , \6359 , \6360 , \6361 , \6362 , \6363 , \6364 ,
         \6365 , \6366 , \6367 , \6368 , \6369 , \6370 , \6371 , \6372 , \6373 , \6374 ,
         \6375 , \6376 , \6377 , \6378 , \6379 , \6380 , \6381 , \6382 , \6383 , \6384 ,
         \6385 , \6386 , \6387 , \6388 , \6389 , \6390 , \6391 , \6392 , \6393 , \6394 ,
         \6395 , \6396 , \6397 , \6398 , \6399 , \6400 , \6401 , \6402 , \6403 , \6404 ,
         \6405 , \6406 , \6407 , \6408 , \6409 , \6410 , \6411 , \6412 , \6413 , \6414 ,
         \6415 , \6416 , \6417 , \6418 , \6419 , \6420 , \6421 , \6422 , \6423 , \6424 ,
         \6425 , \6426 , \6427 , \6428 , \6429 , \6430 , \6431 , \6432 , \6433 , \6434 ,
         \6435 , \6436 , \6437 , \6438 , \6439 , \6440 , \6441 , \6442 , \6443 , \6444 ,
         \6445 , \6446 , \6447 , \6448 , \6449 , \6450 , \6451 , \6452 , \6453 , \6454 ,
         \6455 , \6456 , \6457 , \6458 , \6459 , \6460 , \6461 , \6462 , \6463 , \6464 ,
         \6465 , \6466 , \6467 , \6468 , \6469 , \6470 , \6471 , \6472 , \6473 , \6474 ,
         \6475 , \6476 , \6477 , \6478 , \6479 , \6480 , \6481 , \6482 , \6483 , \6484 ,
         \6485 , \6486 , \6487 , \6488 , \6489 , \6490 , \6491 , \6492 , \6493 , \6494 ,
         \6495 , \6496 , \6497 , \6498 , \6499 , \6500 , \6501 , \6502 , \6503 , \6504 ,
         \6505 , \6506 , \6507 , \6508 , \6509 , \6510 , \6511 , \6512 , \6513 , \6514 ,
         \6515 , \6516 , \6517 , \6518 , \6519 , \6520 , \6521 , \6522 , \6523 , \6524 ,
         \6525 , \6526 , \6527 , \6528 , \6529 , \6530 , \6531 , \6532 , \6533 , \6534 ,
         \6535 , \6536 , \6537 , \6538 , \6539 , \6540 , \6541 , \6542 , \6543 , \6544 ,
         \6545 , \6546 , \6547 , \6548 , \6549 , \6550 , \6551 , \6552 , \6553 , \6554 ,
         \6555 , \6556 , \6557 , \6558 , \6559 , \6560 , \6561 , \6562 , \6563 , \6564 ,
         \6565 , \6566 , \6567 , \6568 , \6569 , \6570 , \6571 , \6572 , \6573 , \6574 ,
         \6575 , \6576 , \6577 , \6578 , \6579 , \6580 , \6581 , \6582 , \6583 , \6584 ,
         \6585 , \6586 , \6587 , \6588 , \6589 , \6590 , \6591 , \6592 , \6593 , \6594 ,
         \6595 , \6596 , \6597 , \6598 , \6599 , \6600 , \6601 , \6602 , \6603 , \6604 ,
         \6605 , \6606 , \6607 , \6608 , \6609 , \6610 , \6611 , \6612 , \6613 , \6614 ,
         \6615 , \6616 , \6617 , \6618 , \6619 , \6620 , \6621 , \6622 , \6623 , \6624 ,
         \6625 , \6626 , \6627 , \6628 , \6629 , \6630 , \6631 , \6632 , \6633 , \6634 ,
         \6635 , \6636 , \6637 , \6638 , \6639 , \6640 , \6641 , \6642 , \6643 , \6644 ,
         \6645 , \6646 , \6647 , \6648 , \6649 , \6650 , \6651 , \6652 , \6653 , \6654 ,
         \6655 , \6656 , \6657 , \6658 , \6659 , \6660 , \6661 , \6662 , \6663 , \6664 ,
         \6665 , \6666 , \6667 , \6668 , \6669 , \6670 , \6671 , \6672 , \6673 , \6674 ,
         \6675 , \6676 , \6677 , \6678 , \6679 , \6680 , \6681 , \6682 , \6683 , \6684 ,
         \6685 , \6686 , \6687 , \6688 , \6689 , \6690 , \6691 , \6692 , \6693 , \6694 ,
         \6695 , \6696 , \6697 , \6698 , \6699 , \6700 , \6701 , \6702 , \6703 , \6704 ,
         \6705 , \6706 , \6707 , \6708 , \6709 , \6710 , \6711 , \6712 , \6713 , \6714 ,
         \6715 , \6716 , \6717 , \6718 , \6719 , \6720 , \6721 , \6722 , \6723 , \6724 ,
         \6725 , \6726 , \6727 , \6728 , \6729 , \6730 , \6731 , \6732 , \6733 , \6734 ,
         \6735 , \6736 , \6737 , \6738 , \6739 , \6740 , \6741 , \6742 , \6743 , \6744 ,
         \6745 , \6746 , \6747 , \6748 , \6749 , \6750 , \6751 , \6752 , \6753 , \6754 ,
         \6755 , \6756 , \6757 , \6758 , \6759 , \6760 , \6761 , \6762 , \6763 , \6764 ,
         \6765 , \6766 , \6767 , \6768 , \6769 , \6770 , \6771 , \6772 , \6773 , \6774 ,
         \6775 , \6776 , \6777 , \6778 , \6779 , \6780 , \6781 , \6782 , \6783 , \6784 ,
         \6785 , \6786 , \6787 , \6788 , \6789 , \6790 , \6791 , \6792 , \6793 , \6794 ,
         \6795 , \6796 , \6797 , \6798 , \6799 , \6800 , \6801 , \6802 , \6803 , \6804 ,
         \6805 , \6806 , \6807 , \6808 , \6809 , \6810 , \6811 , \6812 , \6813 , \6814 ,
         \6815 , \6816 , \6817 , \6818 , \6819 , \6820 , \6821 , \6822 , \6823 , \6824 ,
         \6825 , \6826 , \6827 , \6828 , \6829 , \6830 , \6831 , \6832 , \6833 , \6834 ,
         \6835 , \6836 , \6837 , \6838 , \6839 , \6840 , \6841 , \6842 , \6843 , \6844 ,
         \6845 , \6846 , \6847 , \6848 , \6849 , \6850 , \6851 , \6852 , \6853 , \6854 ,
         \6855 , \6856 , \6857 , \6858 , \6859 , \6860 , \6861 , \6862 , \6863 , \6864 ,
         \6865 , \6866 , \6867 , \6868 , \6869 , \6870 , \6871 , \6872 , \6873 , \6874 ,
         \6875 , \6876 , \6877 , \6878 , \6879 , \6880 , \6881 , \6882 , \6883 , \6884 ,
         \6885 , \6886 , \6887 , \6888 , \6889 , \6890 , \6891 , \6892 , \6893 , \6894 ,
         \6895 , \6896 , \6897 , \6898 , \6899 , \6900 , \6901 , \6902 , \6903 , \6904 ,
         \6905 , \6906 , \6907 , \6908 , \6909 , \6910 , \6911 , \6912 , \6913 , \6914 ,
         \6915 , \6916 , \6917 , \6918 , \6919 , \6920 , \6921 , \6922 , \6923 , \6924 ,
         \6925 , \6926 , \6927 , \6928 , \6929 , \6930 , \6931 , \6932 , \6933 , \6934 ,
         \6935 , \6936 , \6937 , \6938 , \6939 , \6940 , \6941 , \6942 , \6943 , \6944 ,
         \6945 , \6946 , \6947 , \6948 , \6949 , \6950 , \6951 , \6952 , \6953 , \6954 ,
         \6955 , \6956 , \6957 , \6958 , \6959 , \6960 , \6961 , \6962 , \6963 , \6964 ,
         \6965 , \6966 , \6967 , \6968 , \6969 , \6970 , \6971 , \6972 , \6973 , \6974 ,
         \6975 , \6976 , \6977 , \6978 , \6979 , \6980 , \6981 , \6982 , \6983 , \6984 ,
         \6985 , \6986 , \6987 , \6988 , \6989 , \6990 , \6991 , \6992 , \6993 , \6994 ,
         \6995 , \6996 , \6997 , \6998 , \6999 , \7000 , \7001 , \7002 , \7003 , \7004 ,
         \7005 , \7006 , \7007 , \7008 , \7009 , \7010 , \7011 , \7012 , \7013 , \7014 ,
         \7015 , \7016 , \7017 , \7018 , \7019 , \7020 , \7021 , \7022 , \7023 , \7024 ,
         \7025 , \7026 , \7027 , \7028 , \7029 , \7030 , \7031 , \7032 , \7033 , \7034 ,
         \7035 , \7036 , \7037 , \7038 , \7039 , \7040 , \7041 , \7042 , \7043 , \7044 ,
         \7045 , \7046 , \7047 , \7048 , \7049 , \7050 , \7051 , \7052 , \7053 , \7054 ,
         \7055 , \7056 , \7057 , \7058 , \7059 , \7060 , \7061 , \7062 , \7063 , \7064 ,
         \7065 , \7066 , \7067 , \7068 , \7069 , \7070 , \7071 , \7072 , \7073 , \7074 ,
         \7075 , \7076 , \7077 , \7078 , \7079 , \7080 , \7081 , \7082 , \7083 , \7084 ,
         \7085 , \7086 , \7087 , \7088 , \7089 , \7090 , \7091 , \7092 , \7093 , \7094 ,
         \7095 , \7096 , \7097 , \7098 , \7099 , \7100 , \7101 , \7102 , \7103 , \7104 ,
         \7105 , \7106 , \7107 , \7108 , \7109 , \7110 , \7111 , \7112 , \7113 , \7114 ,
         \7115 , \7116 , \7117 , \7118 , \7119 , \7120 , \7121 , \7122 , \7123 , \7124 ,
         \7125 , \7126 , \7127 , \7128 , \7129 , \7130 , \7131 , \7132 , \7133 , \7134 ,
         \7135 , \7136 , \7137 , \7138 , \7139 , \7140 , \7141 , \7142 , \7143 , \7144 ,
         \7145 , \7146 , \7147 , \7148 , \7149 , \7150 , \7151 , \7152 , \7153 , \7154 ,
         \7155 , \7156 , \7157 , \7158 , \7159 , \7160 , \7161 , \7162 , \7163 , \7164 ,
         \7165 , \7166 , \7167 , \7168 , \7169 , \7170 , \7171 , \7172 , \7173 , \7174 ,
         \7175 , \7176 , \7177 , \7178 , \7179 , \7180 , \7181 , \7182 , \7183 , \7184 ,
         \7185 , \7186 , \7187 , \7188 , \7189 , \7190 , \7191 , \7192 , \7193 , \7194 ,
         \7195 , \7196 , \7197 , \7198 , \7199 , \7200 , \7201 , \7202 , \7203 , \7204 ,
         \7205 , \7206 , \7207 , \7208 , \7209 , \7210 , \7211 , \7212 , \7213 , \7214 ,
         \7215 , \7216 , \7217 , \7218 , \7219 , \7220 , \7221 , \7222 , \7223 , \7224 ,
         \7225 , \7226 , \7227 , \7228 , \7229 , \7230 , \7231 , \7232 , \7233 , \7234 ,
         \7235 , \7236 , \7237 , \7238 , \7239 , \7240 , \7241 , \7242 , \7243 , \7244 ,
         \7245 , \7246 , \7247 , \7248 , \7249 , \7250 , \7251 , \7252 , \7253 , \7254 ,
         \7255 , \7256 , \7257 , \7258 , \7259 , \7260 , \7261 , \7262 , \7263 , \7264 ,
         \7265 , \7266 , \7267 , \7268 , \7269 , \7270 , \7271 , \7272 , \7273 , \7274 ,
         \7275 , \7276 , \7277 , \7278 , \7279 , \7280 , \7281 , \7282 , \7283 , \7284 ,
         \7285 , \7286 , \7287 , \7288 , \7289 , \7290 , \7291 , \7292 , \7293 , \7294 ,
         \7295 , \7296 , \7297 , \7298 , \7299 , \7300 , \7301 , \7302 , \7303 , \7304 ,
         \7305 , \7306 , \7307 , \7308 , \7309 , \7310 , \7311 , \7312 , \7313 , \7314 ,
         \7315 , \7316 , \7317 , \7318 , \7319 , \7320 , \7321 , \7322 , \7323 , \7324 ,
         \7325 , \7326 , \7327 , \7328 , \7329 , \7330 , \7331 , \7332 , \7333 , \7334 ,
         \7335 , \7336 , \7337 , \7338 , \7339 , \7340 , \7341 , \7342 , \7343 , \7344 ,
         \7345 , \7346 , \7347 , \7348 , \7349 , \7350 , \7351 , \7352 , \7353 , \7354 ,
         \7355 , \7356 , \7357 , \7358 , \7359 , \7360 , \7361 , \7362 , \7363 , \7364 ,
         \7365 , \7366 , \7367 , \7368 , \7369 , \7370 , \7371 , \7372 , \7373 , \7374 ,
         \7375 , \7376 , \7377 , \7378 , \7379 , \7380 , \7381 , \7382 , \7383 , \7384 ,
         \7385 , \7386 , \7387 , \7388 , \7389 , \7390 , \7391 , \7392 , \7393 , \7394 ,
         \7395 , \7396 , \7397 , \7398 , \7399 , \7400 , \7401 , \7402 , \7403 , \7404 ,
         \7405 , \7406 , \7407 , \7408 , \7409 , \7410 , \7411 , \7412 , \7413 , \7414 ,
         \7415 , \7416 , \7417 , \7418 , \7419 , \7420 , \7421 , \7422 , \7423 , \7424 ,
         \7425 , \7426 , \7427 , \7428 , \7429 , \7430 , \7431 , \7432 , \7433 , \7434 ,
         \7435 , \7436 , \7437 , \7438 , \7439 , \7440 , \7441 , \7442 , \7443 , \7444 ,
         \7445 , \7446 , \7447 , \7448 , \7449 , \7450 , \7451 , \7452 , \7453 , \7454 ,
         \7455 , \7456 , \7457 , \7458 , \7459 , \7460 , \7461 , \7462 , \7463 , \7464 ,
         \7465 , \7466 , \7467 , \7468 , \7469 , \7470 , \7471 , \7472 , \7473 , \7474 ,
         \7475 , \7476 , \7477 , \7478 , \7479 , \7480 , \7481 , \7482 , \7483 , \7484 ,
         \7485 , \7486 , \7487 , \7488 , \7489 , \7490 , \7491 , \7492 , \7493 , \7494 ,
         \7495 , \7496 , \7497 , \7498 , \7499 , \7500 , \7501 , \7502 , \7503 , \7504 ,
         \7505 , \7506 , \7507 , \7508 , \7509 , \7510 , \7511 , \7512 , \7513 , \7514 ,
         \7515 , \7516 , \7517 , \7518 , \7519 , \7520 , \7521 , \7522 , \7523 , \7524 ,
         \7525 , \7526 , \7527 , \7528 , \7529 , \7530 , \7531 , \7532 , \7533 , \7534 ,
         \7535 , \7536 , \7537 , \7538 , \7539 , \7540 , \7541 , \7542 , \7543 , \7544 ,
         \7545 , \7546 , \7547 , \7548 , \7549 , \7550 , \7551 , \7552 , \7553 , \7554 ,
         \7555 , \7556 , \7557 , \7558 , \7559 , \7560 , \7561 , \7562 , \7563 , \7564 ,
         \7565 , \7566 , \7567 , \7568 , \7569 , \7570 , \7571 , \7572 , \7573 , \7574 ,
         \7575 , \7576 , \7577 , \7578 , \7579 , \7580 , \7581 , \7582 , \7583 , \7584 ,
         \7585 , \7586 , \7587 , \7588 , \7589 , \7590 , \7591 , \7592 , \7593 , \7594 ,
         \7595 , \7596 , \7597 , \7598 , \7599 , \7600 , \7601 , \7602 , \7603 , \7604 ,
         \7605 , \7606 , \7607 , \7608 , \7609 , \7610 , \7611 , \7612 , \7613 , \7614 ,
         \7615 , \7616 , \7617 , \7618 , \7619 , \7620 , \7621 , \7622 , \7623 , \7624 ,
         \7625 , \7626 , \7627 , \7628 , \7629 , \7630 , \7631 , \7632 , \7633 , \7634 ,
         \7635 , \7636 , \7637 , \7638 , \7639 , \7640 , \7641 , \7642 , \7643 , \7644 ,
         \7645 , \7646 , \7647 , \7648 , \7649 , \7650 , \7651 , \7652 , \7653 , \7654 ,
         \7655 , \7656 , \7657 , \7658 , \7659 , \7660 , \7661 , \7662 , \7663 , \7664 ,
         \7665 , \7666 , \7667 , \7668 , \7669 , \7670 , \7671 , \7672 , \7673 , \7674 ,
         \7675 , \7676 , \7677 , \7678 , \7679 , \7680 , \7681 , \7682 , \7683 , \7684 ,
         \7685 , \7686 , \7687 , \7688 , \7689 , \7690 , \7691 , \7692 , \7693 , \7694 ,
         \7695 , \7696 , \7697 , \7698 , \7699 , \7700 , \7701 , \7702 , \7703 , \7704 ,
         \7705 , \7706 , \7707 , \7708 , \7709 , \7710 , \7711 , \7712 , \7713 , \7714 ,
         \7715 , \7716 , \7717 , \7718 , \7719 , \7720 , \7721 , \7722 , \7723 , \7724 ,
         \7725 , \7726 , \7727 , \7728 , \7729 , \7730 , \7731 , \7732 , \7733 , \7734 ,
         \7735 , \7736 , \7737 , \7738 , \7739 , \7740 , \7741 , \7742 , \7743 , \7744 ,
         \7745 , \7746 , \7747 , \7748 , \7749 , \7750 , \7751 , \7752 , \7753 , \7754 ,
         \7755 , \7756 , \7757 , \7758 , \7759 , \7760 , \7761 , \7762 , \7763 , \7764 ,
         \7765 , \7766 , \7767 , \7768 , \7769 , \7770 , \7771 , \7772 , \7773 , \7774 ,
         \7775 , \7776 , \7777 , \7778 , \7779 , \7780 , \7781 , \7782 , \7783 , \7784 ,
         \7785 , \7786 , \7787 , \7788 , \7789 , \7790 , \7791 , \7792 , \7793 , \7794 ,
         \7795 , \7796 , \7797 , \7798 , \7799 , \7800 , \7801 , \7802 , \7803 , \7804 ,
         \7805 , \7806 , \7807 , \7808 , \7809 , \7810 , \7811 , \7812 , \7813 , \7814 ,
         \7815 , \7816 , \7817 , \7818 , \7819 , \7820 , \7821 , \7822 , \7823 , \7824 ,
         \7825 , \7826 , \7827 , \7828 , \7829 , \7830 , \7831 , \7832 , \7833 , \7834 ,
         \7835 , \7836 , \7837 , \7838 , \7839 , \7840 , \7841 , \7842 , \7843 , \7844 ,
         \7845 , \7846 , \7847 , \7848 , \7849 , \7850 , \7851 , \7852 , \7853 , \7854 ,
         \7855 , \7856 , \7857 , \7858 , \7859 , \7860 , \7861 , \7862 , \7863 , \7864 ,
         \7865 , \7866 , \7867 , \7868 , \7869 , \7870 , \7871 , \7872 , \7873 , \7874 ,
         \7875 , \7876 , \7877 , \7878 , \7879 , \7880 , \7881 , \7882 , \7883 , \7884 ,
         \7885 , \7886 , \7887 , \7888 , \7889 , \7890 , \7891 , \7892 , \7893 , \7894 ,
         \7895 , \7896 , \7897 , \7898 , \7899 , \7900 , \7901 , \7902 , \7903 , \7904 ,
         \7905 , \7906 , \7907 , \7908 , \7909 , \7910 , \7911 , \7912 , \7913 , \7914 ,
         \7915 , \7916 , \7917 , \7918 , \7919 , \7920 , \7921 , \7922 , \7923 , \7924 ,
         \7925 , \7926 , \7927 , \7928 , \7929 , \7930 , \7931 , \7932 , \7933 , \7934 ,
         \7935 , \7936 , \7937 , \7938 , \7939 , \7940 , \7941 , \7942 , \7943 , \7944 ,
         \7945 , \7946 , \7947 , \7948 , \7949 , \7950 , \7951 , \7952 , \7953 , \7954 ,
         \7955 , \7956 , \7957 , \7958 , \7959 , \7960 , \7961 , \7962 , \7963 , \7964 ,
         \7965 , \7966 , \7967 , \7968 , \7969 , \7970 , \7971 , \7972 , \7973 , \7974 ,
         \7975 , \7976 , \7977 , \7978 , \7979 , \7980 , \7981 , \7982 , \7983 , \7984 ,
         \7985 , \7986 , \7987 , \7988 , \7989 , \7990 , \7991 , \7992 , \7993 , \7994 ,
         \7995 , \7996 , \7997 , \7998 , \7999 , \8000 , \8001 , \8002 , \8003 , \8004 ,
         \8005 , \8006 , \8007 , \8008 , \8009 , \8010 , \8011 , \8012 , \8013 , \8014 ,
         \8015 , \8016 , \8017 , \8018 , \8019 , \8020 , \8021 , \8022 , \8023 , \8024 ,
         \8025 , \8026 , \8027 , \8028 , \8029 , \8030 , \8031 , \8032 , \8033 , \8034 ,
         \8035 , \8036 , \8037 , \8038 , \8039 , \8040 , \8041 , \8042 , \8043 , \8044 ,
         \8045 , \8046 , \8047 , \8048 , \8049 , \8050 , \8051 , \8052 , \8053 , \8054 ,
         \8055 , \8056 , \8057 , \8058 , \8059 , \8060 , \8061 , \8062 , \8063 , \8064 ,
         \8065 , \8066 , \8067 , \8068 , \8069 , \8070 , \8071 , \8072 , \8073 , \8074 ,
         \8075 , \8076 , \8077 , \8078 , \8079 , \8080 , \8081 , \8082 , \8083 , \8084 ,
         \8085 , \8086 , \8087 , \8088 , \8089 , \8090 , \8091 , \8092 , \8093 , \8094 ,
         \8095 , \8096 , \8097 , \8098 , \8099 , \8100 , \8101 , \8102 , \8103 , \8104 ,
         \8105 , \8106 , \8107 , \8108 , \8109 , \8110 , \8111 , \8112 , \8113 , \8114 ,
         \8115 , \8116 , \8117 , \8118 , \8119 , \8120 , \8121 , \8122 , \8123 , \8124 ,
         \8125 , \8126 , \8127 , \8128 , \8129 , \8130 , \8131 , \8132 , \8133 , \8134 ,
         \8135 , \8136 , \8137 , \8138 , \8139 , \8140 , \8141 , \8142 , \8143 , \8144 ,
         \8145 , \8146 , \8147 , \8148 , \8149 , \8150 , \8151 , \8152 , \8153 , \8154 ,
         \8155 , \8156 , \8157 , \8158 , \8159 , \8160 , \8161 , \8162 , \8163 , \8164 ,
         \8165 , \8166 , \8167 , \8168 , \8169 , \8170 , \8171 , \8172 , \8173 , \8174 ,
         \8175 , \8176 , \8177 , \8178 , \8179 , \8180 , \8181 , \8182 , \8183 , \8184 ,
         \8185 , \8186 , \8187 , \8188 , \8189 , \8190 , \8191 , \8192 , \8193 , \8194 ,
         \8195 , \8196 , \8197 , \8198 , \8199 , \8200 , \8201 , \8202 , \8203 , \8204 ,
         \8205 , \8206 , \8207 , \8208 , \8209 , \8210 , \8211 , \8212 , \8213 , \8214 ,
         \8215 , \8216 , \8217 , \8218 , \8219 , \8220 , \8221 , \8222 , \8223 , \8224 ,
         \8225 , \8226 , \8227 , \8228 , \8229 , \8230 , \8231 , \8232 , \8233 , \8234 ,
         \8235 , \8236 , \8237 , \8238 , \8239 , \8240 , \8241 , \8242 , \8243 , \8244 ,
         \8245 , \8246 , \8247 , \8248 , \8249 , \8250 , \8251 , \8252 , \8253 , \8254 ,
         \8255 , \8256 , \8257 , \8258 , \8259 , \8260 , \8261 , \8262 , \8263 , \8264 ,
         \8265 , \8266 , \8267 , \8268 , \8269 , \8270 , \8271 , \8272 , \8273 , \8274 ,
         \8275 , \8276 , \8277 , \8278 , \8279 , \8280 , \8281 , \8282 , \8283 , \8284 ,
         \8285 , \8286 , \8287 , \8288 , \8289 , \8290 , \8291 , \8292 , \8293 , \8294 ,
         \8295 , \8296 , \8297 , \8298 , \8299 , \8300 , \8301 , \8302 , \8303 , \8304 ,
         \8305 , \8306 , \8307 , \8308 , \8309 , \8310 , \8311 , \8312 , \8313 , \8314 ,
         \8315 , \8316 , \8317 , \8318 , \8319 , \8320 , \8321 , \8322 , \8323 , \8324 ,
         \8325 , \8326 , \8327 , \8328 , \8329 , \8330 , \8331 , \8332 , \8333 , \8334 ,
         \8335 , \8336 , \8337 , \8338 , \8339 , \8340 , \8341 , \8342 , \8343 , \8344 ,
         \8345 , \8346 , \8347 , \8348 , \8349 , \8350 , \8351 , \8352 , \8353 , \8354 ,
         \8355 , \8356 , \8357 , \8358 , \8359 , \8360 , \8361 , \8362 , \8363 , \8364 ,
         \8365 , \8366 , \8367 , \8368 , \8369 , \8370 , \8371 , \8372 , \8373 , \8374 ,
         \8375 , \8376 , \8377 , \8378 , \8379 , \8380 , \8381 , \8382 , \8383 , \8384 ,
         \8385 , \8386 , \8387 , \8388 , \8389 , \8390 , \8391 , \8392 , \8393 , \8394 ,
         \8395 , \8396 , \8397 , \8398 , \8399 , \8400 , \8401 , \8402 , \8403 , \8404 ,
         \8405 , \8406 , \8407 , \8408 , \8409 , \8410 , \8411 , \8412 , \8413 , \8414 ,
         \8415 , \8416 , \8417 , \8418 , \8419 , \8420 , \8421 , \8422 , \8423 , \8424 ,
         \8425 , \8426 , \8427 , \8428 , \8429 , \8430 , \8431 , \8432 , \8433 , \8434 ,
         \8435 , \8436 , \8437 , \8438 , \8439 , \8440 , \8441 , \8442 , \8443 , \8444 ,
         \8445 , \8446 , \8447 , \8448 , \8449 , \8450 , \8451 , \8452 , \8453 , \8454 ,
         \8455 , \8456 , \8457 , \8458 , \8459 , \8460 , \8461 , \8462 , \8463 , \8464 ,
         \8465 , \8466 , \8467 , \8468 , \8469 , \8470 , \8471 , \8472 , \8473 , \8474 ,
         \8475 , \8476 , \8477 , \8478 , \8479 , \8480 , \8481 , \8482 , \8483 , \8484 ,
         \8485 , \8486 , \8487 , \8488 , \8489 , \8490 , \8491 , \8492 , \8493 , \8494 ,
         \8495 , \8496 , \8497 , \8498 , \8499 , \8500 , \8501 , \8502 , \8503 , \8504 ,
         \8505 , \8506 , \8507 , \8508 , \8509 , \8510 , \8511 , \8512 , \8513 , \8514 ,
         \8515 , \8516 , \8517 , \8518 , \8519 , \8520 , \8521 , \8522 , \8523 , \8524 ,
         \8525 , \8526 , \8527 , \8528 , \8529 , \8530 , \8531 , \8532 , \8533 , \8534 ,
         \8535 , \8536 , \8537 , \8538 , \8539 , \8540 , \8541 , \8542 , \8543 , \8544 ,
         \8545 , \8546 , \8547 , \8548 , \8549 , \8550 , \8551 , \8552 , \8553 , \8554 ,
         \8555 , \8556 , \8557 , \8558 , \8559 , \8560 , \8561 , \8562 , \8563 , \8564 ,
         \8565 , \8566 , \8567 , \8568 , \8569 , \8570 , \8571 , \8572 , \8573 , \8574 ,
         \8575 , \8576 , \8577 , \8578 , \8579 , \8580 , \8581 , \8582 , \8583 , \8584 ,
         \8585 , \8586 , \8587 , \8588 , \8589 , \8590 , \8591 , \8592 , \8593 , \8594 ,
         \8595 , \8596 , \8597 , \8598 , \8599 , \8600 , \8601 , \8602 , \8603 , \8604 ,
         \8605 , \8606 , \8607 , \8608 , \8609 , \8610 , \8611 , \8612 , \8613 , \8614 ,
         \8615 , \8616 , \8617 , \8618 , \8619 , \8620 , \8621 , \8622 , \8623 , \8624 ,
         \8625 , \8626 , \8627 , \8628 , \8629 , \8630 , \8631 , \8632 , \8633 , \8634 ,
         \8635 , \8636 , \8637 , \8638 , \8639 , \8640 , \8641 , \8642 , \8643 , \8644 ,
         \8645 , \8646 , \8647 , \8648 , \8649 , \8650 , \8651 , \8652 , \8653 , \8654 ,
         \8655 , \8656 , \8657 , \8658 , \8659 , \8660 , \8661 , \8662 , \8663 , \8664 ,
         \8665 , \8666 , \8667 , \8668 , \8669 , \8670 , \8671 , \8672 , \8673 , \8674 ,
         \8675 , \8676 , \8677 , \8678 , \8679 , \8680 , \8681 , \8682 , \8683 , \8684 ,
         \8685 , \8686 , \8687 , \8688 , \8689 , \8690 , \8691 , \8692 , \8693 , \8694 ,
         \8695 , \8696 , \8697 , \8698 , \8699 , \8700 , \8701 , \8702 , \8703 , \8704 ,
         \8705 , \8706 , \8707 , \8708 , \8709 , \8710 , \8711 , \8712 , \8713 , \8714 ,
         \8715 , \8716 , \8717 , \8718 , \8719 , \8720 , \8721 , \8722 , \8723 , \8724 ,
         \8725 , \8726 , \8727 , \8728 , \8729 , \8730 , \8731 , \8732 , \8733 , \8734 ,
         \8735 , \8736 , \8737 , \8738 , \8739 , \8740 , \8741 , \8742 , \8743 , \8744 ,
         \8745 , \8746 , \8747 , \8748 , \8749 , \8750 , \8751 , \8752 , \8753 , \8754 ,
         \8755 , \8756 , \8757 , \8758 , \8759 , \8760 , \8761 , \8762 , \8763 , \8764 ,
         \8765 , \8766 , \8767 , \8768 , \8769 , \8770 , \8771 , \8772 , \8773 , \8774 ,
         \8775 , \8776 , \8777 , \8778 , \8779 , \8780 , \8781 , \8782 , \8783 , \8784 ,
         \8785 , \8786 , \8787 , \8788 , \8789 , \8790 , \8791 , \8792 , \8793 , \8794 ,
         \8795 , \8796 , \8797 , \8798 , \8799 , \8800 , \8801 , \8802 , \8803 , \8804 ,
         \8805 , \8806 , \8807 , \8808 , \8809 , \8810 , \8811 , \8812 , \8813 , \8814 ,
         \8815 , \8816 , \8817 , \8818 , \8819 , \8820 , \8821 , \8822 , \8823 , \8824 ,
         \8825 , \8826 , \8827 , \8828 , \8829 , \8830 , \8831 , \8832 , \8833 , \8834 ,
         \8835 , \8836 , \8837 , \8838 , \8839 , \8840 , \8841 , \8842 , \8843 , \8844 ,
         \8845 , \8846 , \8847 , \8848 , \8849 , \8850 , \8851 , \8852 , \8853 , \8854 ,
         \8855 , \8856 , \8857 , \8858 , \8859 , \8860 , \8861 , \8862 , \8863 , \8864 ,
         \8865 , \8866 , \8867 , \8868 , \8869 , \8870 , \8871 , \8872 , \8873 , \8874 ,
         \8875 , \8876 , \8877 , \8878 , \8879 , \8880 , \8881 , \8882 , \8883 , \8884 ,
         \8885 , \8886 , \8887 , \8888 , \8889 , \8890 , \8891 , \8892 , \8893 , \8894 ,
         \8895 , \8896 , \8897 , \8898 , \8899 , \8900 , \8901 , \8902 , \8903 , \8904 ,
         \8905 , \8906 , \8907 , \8908 , \8909 , \8910 , \8911 , \8912 , \8913 , \8914 ,
         \8915 , \8916 , \8917 , \8918 , \8919 , \8920 , \8921 , \8922 , \8923 , \8924 ,
         \8925 , \8926 , \8927 , \8928 , \8929 , \8930 , \8931 , \8932 , \8933 , \8934 ,
         \8935 , \8936 , \8937 , \8938 , \8939 , \8940 , \8941 , \8942 , \8943 , \8944 ,
         \8945 , \8946 , \8947 , \8948 , \8949 , \8950 , \8951 , \8952 , \8953 , \8954 ,
         \8955 , \8956 , \8957 , \8958 , \8959 , \8960 , \8961 , \8962 , \8963 , \8964 ,
         \8965 , \8966 , \8967 , \8968 , \8969 , \8970 , \8971 , \8972 , \8973 , \8974 ,
         \8975 , \8976 , \8977 , \8978 , \8979 , \8980 , \8981 , \8982 , \8983 , \8984 ,
         \8985 , \8986 , \8987 , \8988 , \8989 , \8990 , \8991 , \8992 , \8993 , \8994 ,
         \8995 , \8996 , \8997 , \8998 , \8999 , \9000 , \9001 , \9002 , \9003 , \9004 ,
         \9005 , \9006 , \9007 , \9008 , \9009 , \9010 , \9011 , \9012 , \9013 , \9014 ,
         \9015 , \9016 , \9017 , \9018 , \9019 , \9020 , \9021 , \9022 , \9023 , \9024 ,
         \9025 , \9026 , \9027 , \9028 , \9029 , \9030 , \9031 , \9032 , \9033 , \9034 ,
         \9035 , \9036 , \9037 , \9038 , \9039 , \9040 , \9041 , \9042 , \9043 , \9044 ,
         \9045 , \9046 , \9047 , \9048 , \9049 , \9050 , \9051 , \9052 , \9053 , \9054 ,
         \9055 , \9056 , \9057 , \9058 , \9059 , \9060 , \9061 , \9062 , \9063 , \9064 ,
         \9065 , \9066 , \9067 , \9068 , \9069 , \9070 , \9071 , \9072 , \9073 , \9074 ,
         \9075 , \9076 , \9077 , \9078 , \9079 , \9080 , \9081 , \9082 , \9083 , \9084 ,
         \9085 , \9086 , \9087 , \9088 , \9089 , \9090 , \9091 , \9092 , \9093 , \9094 ,
         \9095 , \9096 , \9097 , \9098 , \9099 , \9100 , \9101 , \9102 , \9103 , \9104 ,
         \9105 , \9106 , \9107 , \9108 , \9109 , \9110 , \9111 , \9112 , \9113 , \9114 ,
         \9115 , \9116 , \9117 , \9118 , \9119 , \9120 , \9121 , \9122 , \9123 , \9124 ,
         \9125 , \9126 , \9127 , \9128 , \9129 , \9130 , \9131 , \9132 , \9133 , \9134 ,
         \9135 , \9136 , \9137 , \9138 , \9139 , \9140 , \9141 , \9142 , \9143 , \9144 ,
         \9145 , \9146 , \9147 , \9148 , \9149 , \9150 , \9151 , \9152 , \9153 , \9154 ,
         \9155 , \9156 , \9157 , \9158 , \9159 , \9160 , \9161 , \9162 , \9163 , \9164 ,
         \9165 , \9166 , \9167 , \9168 , \9169 , \9170 , \9171 , \9172 , \9173 , \9174 ,
         \9175 , \9176 , \9177 , \9178 , \9179 , \9180 , \9181 , \9182 , \9183 , \9184 ,
         \9185 , \9186 , \9187 , \9188 , \9189 , \9190 , \9191 , \9192 , \9193 , \9194 ,
         \9195 , \9196 , \9197 , \9198 , \9199 , \9200 , \9201 , \9202 , \9203 , \9204 ,
         \9205 , \9206 , \9207 , \9208 , \9209 , \9210 , \9211 , \9212 , \9213 , \9214 ,
         \9215 , \9216 , \9217 , \9218 , \9219 , \9220 , \9221 , \9222 , \9223 , \9224 ,
         \9225 , \9226 , \9227 , \9228 , \9229 , \9230 , \9231 , \9232 , \9233 , \9234 ,
         \9235 , \9236 , \9237 , \9238 , \9239 , \9240 , \9241 , \9242 , \9243 , \9244 ,
         \9245 , \9246 , \9247 , \9248 , \9249 , \9250 , \9251 , \9252 , \9253 , \9254 ,
         \9255 , \9256 , \9257 , \9258 , \9259 , \9260 , \9261 , \9262 , \9263 , \9264 ,
         \9265 , \9266 , \9267 , \9268 , \9269 , \9270 , \9271 , \9272 , \9273 , \9274 ,
         \9275 , \9276 , \9277 , \9278 , \9279 , \9280 , \9281 , \9282 , \9283 , \9284 ,
         \9285 , \9286 , \9287 , \9288 , \9289 , \9290 , \9291 , \9292 , \9293 , \9294 ,
         \9295 , \9296 , \9297 , \9298 , \9299 , \9300 , \9301 , \9302 , \9303 , \9304 ,
         \9305 , \9306 , \9307 , \9308 , \9309 , \9310 , \9311 , \9312 , \9313 , \9314 ,
         \9315 , \9316 , \9317 , \9318 , \9319 , \9320 , \9321 , \9322 , \9323 , \9324 ,
         \9325 , \9326 , \9327 , \9328 , \9329 , \9330 , \9331 , \9332 , \9333 , \9334 ,
         \9335 , \9336 , \9337 , \9338 , \9339 , \9340 , \9341 , \9342 , \9343 , \9344 ,
         \9345 , \9346 , \9347 , \9348 , \9349 , \9350 , \9351 , \9352 , \9353 , \9354 ,
         \9355 , \9356 , \9357 , \9358 , \9359 , \9360 , \9361 , \9362 , \9363 , \9364 ,
         \9365 , \9366 , \9367 , \9368 , \9369 , \9370 , \9371 , \9372 , \9373 , \9374 ,
         \9375 , \9376 , \9377 , \9378 , \9379 , \9380 , \9381 , \9382 , \9383 , \9384 ,
         \9385 , \9386 , \9387 , \9388 , \9389 , \9390 , \9391 , \9392 , \9393 , \9394 ,
         \9395 , \9396 , \9397 , \9398 , \9399 , \9400 , \9401 , \9402 , \9403 , \9404 ,
         \9405 , \9406 , \9407 , \9408 , \9409 , \9410 , \9411 , \9412 , \9413 , \9414 ,
         \9415 , \9416 , \9417 , \9418 , \9419 , \9420 , \9421 , \9422 , \9423 , \9424 ,
         \9425 , \9426 , \9427 , \9428 , \9429 , \9430 , \9431 , \9432 , \9433 , \9434 ,
         \9435 , \9436 , \9437 , \9438 , \9439 , \9440 , \9441 , \9442 , \9443 , \9444 ,
         \9445 , \9446 , \9447 , \9448 , \9449 , \9450 , \9451 , \9452 , \9453 , \9454 ,
         \9455 , \9456 , \9457 , \9458 , \9459 , \9460 , \9461 , \9462 , \9463 , \9464 ,
         \9465 , \9466 , \9467 , \9468 , \9469 , \9470 , \9471 , \9472 , \9473 , \9474 ,
         \9475 , \9476 , \9477 , \9478 , \9479 , \9480 , \9481 , \9482 , \9483 , \9484 ,
         \9485 , \9486 , \9487 , \9488 , \9489 , \9490 , \9491 , \9492 , \9493 , \9494 ,
         \9495 , \9496 , \9497 , \9498 , \9499 , \9500 , \9501 , \9502 , \9503 , \9504 ,
         \9505 , \9506 , \9507 , \9508 , \9509 , \9510 , \9511 , \9512 , \9513 , \9514 ,
         \9515 , \9516 , \9517 , \9518 , \9519 , \9520 , \9521 , \9522 , \9523 , \9524 ,
         \9525 , \9526 , \9527 , \9528 , \9529 , \9530 , \9531 , \9532 , \9533 , \9534 ,
         \9535 , \9536 , \9537 , \9538 , \9539 , \9540 , \9541 , \9542 , \9543 , \9544 ,
         \9545 , \9546 , \9547 , \9548 , \9549 , \9550 , \9551 , \9552 , \9553 , \9554 ,
         \9555 , \9556 , \9557 , \9558 , \9559 , \9560 , \9561 , \9562 , \9563 , \9564 ,
         \9565 , \9566 , \9567 , \9568 , \9569 , \9570 , \9571 , \9572 , \9573 , \9574 ,
         \9575 , \9576 , \9577 , \9578 , \9579 , \9580 , \9581 , \9582 , \9583 , \9584 ,
         \9585 , \9586 , \9587 , \9588 , \9589 , \9590 , \9591 , \9592 , \9593 , \9594 ,
         \9595 , \9596 , \9597 , \9598 , \9599 , \9600 , \9601 , \9602 , \9603 , \9604 ,
         \9605 , \9606 , \9607 , \9608 , \9609 , \9610 , \9611 , \9612 , \9613 , \9614 ,
         \9615 , \9616 , \9617 , \9618 , \9619 , \9620 , \9621 , \9622 , \9623 , \9624 ,
         \9625 , \9626 , \9627 , \9628 , \9629 , \9630 , \9631 , \9632 , \9633 , \9634 ,
         \9635 , \9636 , \9637 , \9638 , \9639 , \9640 , \9641 , \9642 , \9643 , \9644 ,
         \9645 , \9646 , \9647 , \9648 , \9649 , \9650 , \9651 , \9652 , \9653 , \9654 ,
         \9655 , \9656 , \9657 , \9658 , \9659 , \9660 , \9661 , \9662 , \9663 , \9664 ,
         \9665 , \9666 , \9667 , \9668 , \9669 , \9670 , \9671 , \9672 , \9673 , \9674 ,
         \9675 , \9676 , \9677 , \9678 , \9679 , \9680 , \9681 , \9682 , \9683 , \9684 ,
         \9685 , \9686 , \9687 , \9688 , \9689 , \9690 , \9691 , \9692 , \9693 , \9694 ,
         \9695 , \9696 , \9697 , \9698 , \9699 , \9700 , \9701 , \9702 , \9703 , \9704 ,
         \9705 , \9706 , \9707 , \9708 , \9709 , \9710 , \9711 , \9712 , \9713 , \9714 ,
         \9715 , \9716 , \9717 , \9718 , \9719 , \9720 , \9721 , \9722 , \9723 , \9724 ,
         \9725 , \9726 , \9727 , \9728 , \9729 , \9730 , \9731 , \9732 , \9733 , \9734 ,
         \9735 , \9736 , \9737 , \9738 , \9739 , \9740 , \9741 , \9742 , \9743 , \9744 ,
         \9745 , \9746 , \9747 , \9748 , \9749 , \9750 , \9751 , \9752 , \9753 , \9754 ,
         \9755 , \9756 , \9757 , \9758 , \9759 , \9760 , \9761 , \9762 , \9763 , \9764 ,
         \9765 , \9766 , \9767 , \9768 , \9769 , \9770 , \9771 , \9772 , \9773 , \9774 ,
         \9775 , \9776 , \9777 , \9778 , \9779 , \9780 , \9781 , \9782 , \9783 , \9784 ,
         \9785 , \9786 , \9787 , \9788 , \9789 , \9790 , \9791 , \9792 , \9793 , \9794 ,
         \9795 , \9796 , \9797 , \9798 , \9799 , \9800 , \9801 , \9802 , \9803 , \9804 ,
         \9805 , \9806 , \9807 , \9808 , \9809 , \9810 , \9811 , \9812 , \9813 , \9814 ,
         \9815 , \9816 , \9817 , \9818 , \9819 , \9820 , \9821 , \9822 , \9823 , \9824 ,
         \9825 , \9826 , \9827 , \9828 , \9829 , \9830 , \9831 , \9832 , \9833 , \9834 ,
         \9835 , \9836 , \9837 , \9838 , \9839 , \9840 , \9841 , \9842 , \9843 , \9844 ,
         \9845 , \9846 , \9847 , \9848 , \9849 , \9850 , \9851 , \9852 , \9853 , \9854 ,
         \9855 , \9856 , \9857 , \9858 , \9859 , \9860 , \9861 , \9862 , \9863 , \9864 ,
         \9865 , \9866 , \9867 , \9868 , \9869 , \9870 , \9871 , \9872 , \9873 , \9874 ,
         \9875 , \9876 , \9877 , \9878 , \9879 , \9880 , \9881 , \9882 , \9883 , \9884 ,
         \9885 , \9886 , \9887 , \9888 , \9889 , \9890 , \9891 , \9892 , \9893 , \9894 ,
         \9895 , \9896 , \9897 , \9898 , \9899 , \9900 , \9901 , \9902 , \9903 , \9904 ,
         \9905 , \9906 , \9907 , \9908 , \9909 , \9910 , \9911 , \9912 , \9913 , \9914 ,
         \9915 , \9916 , \9917 , \9918 , \9919 , \9920 , \9921 , \9922 , \9923 , \9924 ,
         \9925 , \9926 , \9927 , \9928 , \9929 , \9930 , \9931 , \9932 , \9933 , \9934 ,
         \9935 , \9936 , \9937 , \9938 , \9939 , \9940 , \9941 , \9942 , \9943 , \9944 ,
         \9945 , \9946 , \9947 , \9948 , \9949 , \9950 , \9951 , \9952 , \9953 , \9954 ,
         \9955 , \9956 , \9957 , \9958 , \9959 , \9960 , \9961 , \9962 , \9963 , \9964 ,
         \9965 , \9966 , \9967 , \9968 , \9969 , \9970 , \9971 , \9972 , \9973 , \9974 ,
         \9975 , \9976 , \9977 , \9978 , \9979 , \9980 , \9981 , \9982 , \9983 , \9984 ,
         \9985 , \9986 , \9987 , \9988 , \9989 , \9990 , \9991 , \9992 , \9993 , \9994 ,
         \9995 , \9996 , \9997 , \9998 , \9999 , \10000 , \10001 , \10002 , \10003 , \10004 ,
         \10005 , \10006 , \10007 , \10008 , \10009 , \10010 , \10011 , \10012 , \10013 , \10014 ,
         \10015 , \10016 , \10017 , \10018 , \10019 , \10020 , \10021 , \10022 , \10023 , \10024 ,
         \10025 , \10026 , \10027 , \10028 , \10029 , \10030 , \10031 , \10032 , \10033 , \10034 ,
         \10035 , \10036 , \10037 , \10038 , \10039 , \10040 , \10041 , \10042 , \10043 , \10044 ,
         \10045 , \10046 , \10047 , \10048 , \10049 , \10050 , \10051 , \10052 , \10053 , \10054 ,
         \10055 , \10056 , \10057 , \10058 , \10059 , \10060 , \10061 , \10062 , \10063 , \10064 ,
         \10065 , \10066 , \10067 , \10068 , \10069 , \10070 , \10071 , \10072 , \10073 , \10074 ,
         \10075 , \10076 , \10077 , \10078 , \10079 , \10080 , \10081 , \10082 , \10083 , \10084 ,
         \10085 , \10086 , \10087 , \10088 , \10089 , \10090 , \10091 , \10092 , \10093 , \10094 ,
         \10095 , \10096 , \10097 , \10098 , \10099 , \10100 , \10101 , \10102 , \10103 , \10104 ,
         \10105 , \10106 , \10107 , \10108 , \10109 , \10110 , \10111 , \10112 , \10113 , \10114 ,
         \10115 , \10116 , \10117 , \10118 , \10119 , \10120 , \10121 , \10122 , \10123 , \10124 ,
         \10125 , \10126 , \10127 , \10128 , \10129 , \10130 , \10131 , \10132 , \10133 , \10134 ,
         \10135 , \10136 , \10137 , \10138 , \10139 , \10140 , \10141 , \10142 , \10143 , \10144 ,
         \10145 , \10146 , \10147 , \10148 , \10149 , \10150 , \10151 , \10152 , \10153 , \10154 ,
         \10155 , \10156 , \10157 , \10158 , \10159 , \10160 , \10161 , \10162 , \10163 , \10164 ,
         \10165 , \10166 , \10167 , \10168 , \10169 , \10170 , \10171 , \10172 , \10173 , \10174 ,
         \10175 , \10176 , \10177 , \10178 , \10179 , \10180 , \10181 , \10182 , \10183 , \10184 ,
         \10185 , \10186 , \10187 , \10188 , \10189 , \10190 , \10191 , \10192 , \10193 , \10194 ,
         \10195 , \10196 , \10197 , \10198 , \10199 , \10200 , \10201 , \10202 , \10203 , \10204 ,
         \10205 , \10206 , \10207 , \10208 , \10209 , \10210 , \10211 , \10212 , \10213 , \10214 ,
         \10215 , \10216 , \10217 , \10218 , \10219 , \10220 , \10221 , \10222 , \10223 , \10224 ,
         \10225 , \10226 , \10227 , \10228 , \10229 , \10230 , \10231 , \10232 , \10233 , \10234 ,
         \10235 , \10236 , \10237 , \10238 , \10239 , \10240 , \10241 , \10242 , \10243 , \10244 ,
         \10245 , \10246 , \10247 , \10248 , \10249 , \10250 , \10251 , \10252 , \10253 , \10254 ,
         \10255 , \10256 , \10257 , \10258 , \10259 , \10260 , \10261 , \10262 , \10263 , \10264 ,
         \10265 , \10266 , \10267 , \10268 , \10269 , \10270 , \10271 , \10272 , \10273 , \10274 ,
         \10275 , \10276 , \10277 , \10278 , \10279 , \10280 , \10281 , \10282 , \10283 , \10284 ,
         \10285 , \10286 , \10287 , \10288 , \10289 , \10290 , \10291 , \10292 , \10293 , \10294 ,
         \10295 , \10296 , \10297 , \10298 , \10299 , \10300 , \10301 , \10302 , \10303 , \10304 ,
         \10305 , \10306 , \10307 , \10308 , \10309 , \10310 , \10311 , \10312 , \10313 , \10314 ,
         \10315 , \10316 , \10317 , \10318 , \10319 , \10320 , \10321 , \10322 , \10323 , \10324 ,
         \10325 , \10326 , \10327 , \10328 , \10329 , \10330 , \10331 , \10332 , \10333 , \10334 ,
         \10335 , \10336 , \10337 , \10338 , \10339 , \10340 , \10341 , \10342 , \10343 , \10344 ,
         \10345 , \10346 , \10347 , \10348 , \10349 , \10350 , \10351 , \10352 , \10353 , \10354 ,
         \10355 , \10356 , \10357 , \10358 , \10359 , \10360 , \10361 , \10362 , \10363 , \10364 ,
         \10365 , \10366 , \10367 , \10368 , \10369 , \10370 , \10371 , \10372 , \10373 , \10374 ,
         \10375 , \10376 , \10377 , \10378 , \10379 , \10380 , \10381 , \10382 , \10383 , \10384 ,
         \10385 , \10386 , \10387 , \10388 , \10389 , \10390 , \10391 , \10392 , \10393 , \10394 ,
         \10395 , \10396 , \10397 , \10398 , \10399 , \10400 , \10401 , \10402 , \10403 , \10404 ,
         \10405 , \10406 , \10407 , \10408 , \10409 , \10410 , \10411 , \10412 , \10413 , \10414 ,
         \10415 , \10416 , \10417 , \10418 , \10419 , \10420 , \10421 , \10422 , \10423 , \10424 ,
         \10425 , \10426 , \10427 , \10428 , \10429 , \10430 , \10431 , \10432 , \10433 , \10434 ,
         \10435 , \10436 , \10437 , \10438 , \10439 , \10440 , \10441 , \10442 , \10443 , \10444 ,
         \10445 , \10446 , \10447 , \10448 , \10449 , \10450 , \10451 , \10452 , \10453 , \10454 ,
         \10455 , \10456 , \10457 , \10458 , \10459 , \10460 , \10461 , \10462 , \10463 , \10464 ,
         \10465 , \10466 , \10467 , \10468 , \10469 , \10470 , \10471 , \10472 , \10473 , \10474 ,
         \10475 , \10476 , \10477 , \10478 , \10479 , \10480 , \10481 , \10482 , \10483 , \10484 ,
         \10485 , \10486 , \10487 , \10488 , \10489 , \10490 , \10491 , \10492 , \10493 , \10494 ,
         \10495 , \10496 , \10497 , \10498 , \10499 , \10500 , \10501 , \10502 , \10503 , \10504 ,
         \10505 , \10506 , \10507 , \10508 , \10509 , \10510 , \10511 , \10512 , \10513 , \10514 ,
         \10515 , \10516 , \10517 , \10518 , \10519 , \10520 , \10521 , \10522 , \10523 , \10524 ,
         \10525 , \10526 , \10527 , \10528 , \10529 , \10530 , \10531 , \10532 , \10533 , \10534 ,
         \10535 , \10536 , \10537 , \10538 , \10539 , \10540 , \10541 , \10542 , \10543 , \10544 ,
         \10545 , \10546 , \10547 , \10548 , \10549 , \10550 , \10551 , \10552 , \10553 , \10554 ,
         \10555 , \10556 , \10557 , \10558 , \10559 , \10560 , \10561 , \10562 , \10563 , \10564 ,
         \10565 , \10566 , \10567 , \10568 , \10569 , \10570 , \10571 , \10572 , \10573 , \10574 ,
         \10575 , \10576 , \10577 , \10578 , \10579 , \10580 , \10581 , \10582 , \10583 , \10584 ,
         \10585 , \10586 , \10587 , \10588 , \10589 , \10590 , \10591 , \10592 , \10593 , \10594 ,
         \10595 , \10596 , \10597 , \10598 , \10599 , \10600 , \10601 , \10602 , \10603 , \10604 ,
         \10605 , \10606 , \10607 , \10608 , \10609 , \10610 , \10611 , \10612 , \10613 , \10614 ,
         \10615 , \10616 , \10617 , \10618 , \10619 , \10620 , \10621 , \10622 , \10623 , \10624 ,
         \10625 , \10626 , \10627 , \10628 , \10629 , \10630 , \10631 , \10632 , \10633 , \10634 ,
         \10635 , \10636 , \10637 , \10638 , \10639 , \10640 , \10641 , \10642 , \10643 , \10644 ,
         \10645 , \10646 , \10647 , \10648 , \10649 , \10650 , \10651 , \10652 , \10653 , \10654 ,
         \10655 , \10656 , \10657 , \10658 , \10659 , \10660 , \10661 , \10662 , \10663 , \10664 ,
         \10665 , \10666 , \10667 , \10668 , \10669 , \10670 , \10671 , \10672 , \10673 , \10674 ,
         \10675 , \10676 , \10677 , \10678 , \10679 , \10680 , \10681 , \10682 , \10683 , \10684 ,
         \10685 , \10686 , \10687 , \10688 , \10689 , \10690 , \10691 , \10692 , \10693 , \10694 ,
         \10695 , \10696 , \10697 , \10698 , \10699 , \10700 , \10701 , \10702 , \10703 , \10704 ,
         \10705 , \10706 , \10707 , \10708 , \10709 , \10710 , \10711 , \10712 , \10713 , \10714 ,
         \10715 , \10716 , \10717 , \10718 , \10719 , \10720 , \10721 , \10722 , \10723 , \10724 ,
         \10725 , \10726 , \10727 , \10728 , \10729 , \10730 , \10731 , \10732 , \10733 , \10734 ,
         \10735 , \10736 , \10737 , \10738 , \10739 , \10740 , \10741 , \10742 , \10743 , \10744 ,
         \10745 , \10746 , \10747 , \10748 , \10749 , \10750 , \10751 , \10752 , \10753 , \10754 ,
         \10755 , \10756 , \10757 , \10758 , \10759 , \10760 , \10761 , \10762 , \10763 , \10764 ,
         \10765 , \10766 , \10767 , \10768 , \10769 , \10770 , \10771 , \10772 , \10773 , \10774 ,
         \10775 , \10776 , \10777 , \10778 , \10779 , \10780 , \10781 , \10782 , \10783 , \10784 ,
         \10785 , \10786 , \10787 , \10788 , \10789 , \10790 , \10791 , \10792 , \10793 , \10794 ,
         \10795 , \10796 , \10797 , \10798 , \10799 , \10800 , \10801 , \10802 , \10803 , \10804 ,
         \10805 , \10806 , \10807 , \10808 , \10809 , \10810 , \10811 , \10812 , \10813 , \10814 ,
         \10815 , \10816 , \10817 , \10818 , \10819 , \10820 , \10821 , \10822 , \10823 , \10824 ,
         \10825 , \10826 , \10827 , \10828 , \10829 , \10830 , \10831 , \10832 , \10833 , \10834 ,
         \10835 , \10836 , \10837 , \10838 , \10839 , \10840 , \10841 , \10842 , \10843 , \10844 ,
         \10845 , \10846 , \10847 , \10848 , \10849 , \10850 , \10851 , \10852 , \10853 , \10854 ,
         \10855 , \10856 , \10857 , \10858 , \10859 , \10860 , \10861 , \10862 , \10863 , \10864 ,
         \10865 , \10866 , \10867 , \10868 , \10869 , \10870 , \10871 , \10872 , \10873 , \10874 ,
         \10875 , \10876 , \10877 , \10878 , \10879 , \10880 , \10881 , \10882 , \10883 , \10884 ,
         \10885 , \10886 , \10887 , \10888 , \10889 , \10890 , \10891 , \10892 , \10893 , \10894 ,
         \10895 , \10896 , \10897 , \10898 , \10899 , \10900 , \10901 , \10902 , \10903 , \10904 ,
         \10905 , \10906 , \10907 , \10908 , \10909 , \10910 , \10911 , \10912 , \10913 , \10914 ,
         \10915 , \10916 , \10917 , \10918 , \10919 , \10920 , \10921 , \10922 , \10923 , \10924 ,
         \10925 , \10926 , \10927 , \10928 , \10929 , \10930 , \10931 , \10932 , \10933 , \10934 ,
         \10935 , \10936 , \10937 , \10938 , \10939 , \10940 , \10941 , \10942 , \10943 , \10944 ,
         \10945 , \10946 , \10947 , \10948 , \10949 , \10950 , \10951 , \10952 , \10953 , \10954 ,
         \10955 , \10956 , \10957 , \10958 , \10959 , \10960 , \10961 , \10962 , \10963 , \10964 ,
         \10965 , \10966 , \10967 , \10968 , \10969 , \10970 , \10971 , \10972 , \10973 , \10974 ,
         \10975 , \10976 , \10977 , \10978 , \10979 , \10980 , \10981 , \10982 , \10983 , \10984 ,
         \10985 , \10986 , \10987 , \10988 , \10989 , \10990 , \10991 , \10992 , \10993 , \10994 ,
         \10995 , \10996 , \10997 , \10998 , \10999 , \11000 , \11001 , \11002 , \11003 , \11004 ,
         \11005 , \11006 , \11007 , \11008 , \11009 , \11010 , \11011 , \11012 , \11013 , \11014 ,
         \11015 , \11016 , \11017 , \11018 , \11019 , \11020 , \11021 , \11022 , \11023 , \11024 ,
         \11025 , \11026 , \11027 , \11028 , \11029 , \11030 , \11031 , \11032 , \11033 , \11034 ,
         \11035 , \11036 , \11037 , \11038 , \11039 , \11040 , \11041 , \11042 , \11043 , \11044 ,
         \11045 , \11046 , \11047 , \11048 , \11049 , \11050 , \11051 , \11052 , \11053 , \11054 ,
         \11055 , \11056 , \11057 , \11058 , \11059 , \11060 , \11061 , \11062 , \11063 , \11064 ,
         \11065 , \11066 , \11067 , \11068 , \11069 , \11070 , \11071 , \11072 , \11073 , \11074 ,
         \11075 , \11076 , \11077 , \11078 , \11079 , \11080 , \11081 , \11082 , \11083 , \11084 ,
         \11085 , \11086 , \11087 , \11088 , \11089 , \11090 , \11091 , \11092 , \11093 , \11094 ,
         \11095 , \11096 , \11097 , \11098 , \11099 , \11100 , \11101 , \11102 , \11103 , \11104 ,
         \11105 , \11106 , \11107 , \11108 , \11109 , \11110 , \11111 , \11112 , \11113 , \11114 ,
         \11115 , \11116 , \11117 , \11118 , \11119 , \11120 , \11121 , \11122 , \11123 , \11124 ,
         \11125 , \11126 , \11127 , \11128 , \11129 , \11130 , \11131 , \11132 , \11133 , \11134 ,
         \11135 , \11136 , \11137 , \11138 , \11139 , \11140 , \11141 , \11142 , \11143 , \11144 ,
         \11145 , \11146 , \11147 , \11148 , \11149 , \11150 , \11151 , \11152 , \11153 , \11154 ,
         \11155 , \11156 , \11157 , \11158 , \11159 , \11160 , \11161 , \11162 , \11163 , \11164 ,
         \11165 , \11166 , \11167 , \11168 , \11169 , \11170 , \11171 , \11172 , \11173 , \11174 ,
         \11175 , \11176 , \11177 , \11178 , \11179 , \11180 , \11181 , \11182 , \11183 , \11184 ,
         \11185 , \11186 , \11187 , \11188 , \11189 , \11190 , \11191 , \11192 , \11193 , \11194 ,
         \11195 , \11196 , \11197 , \11198 , \11199 , \11200 , \11201 , \11202 , \11203 , \11204 ,
         \11205 , \11206 , \11207 , \11208 , \11209 , \11210 , \11211 , \11212 , \11213 , \11214 ,
         \11215 , \11216 , \11217 , \11218 , \11219 , \11220 , \11221 , \11222 , \11223 , \11224 ,
         \11225 , \11226 , \11227 , \11228 , \11229 , \11230 , \11231 , \11232 , \11233 , \11234 ,
         \11235 , \11236 , \11237 , \11238 , \11239 , \11240 , \11241 , \11242 , \11243 , \11244 ,
         \11245 , \11246 , \11247 , \11248 , \11249 , \11250 , \11251 , \11252 , \11253 , \11254 ,
         \11255 , \11256 , \11257 , \11258 , \11259 , \11260 , \11261 , \11262 , \11263 , \11264 ,
         \11265 , \11266 , \11267 , \11268 , \11269 , \11270 , \11271 , \11272 , \11273 , \11274 ,
         \11275 , \11276 , \11277 , \11278 , \11279 , \11280 , \11281 , \11282 , \11283 , \11284 ,
         \11285 , \11286 , \11287 , \11288 , \11289 , \11290 , \11291 , \11292 , \11293 , \11294 ,
         \11295 , \11296 , \11297 , \11298 , \11299 , \11300 , \11301 , \11302 , \11303 , \11304 ,
         \11305 , \11306 , \11307 , \11308 , \11309 , \11310 , \11311 , \11312 , \11313 , \11314 ,
         \11315 , \11316 , \11317 , \11318 , \11319 , \11320 , \11321 , \11322 , \11323 , \11324 ,
         \11325 , \11326 , \11327 , \11328 , \11329 , \11330 , \11331 , \11332 , \11333 , \11334 ,
         \11335 , \11336 , \11337 , \11338 , \11339 , \11340 , \11341 , \11342 , \11343 , \11344 ,
         \11345 , \11346 , \11347 , \11348 , \11349 , \11350 , \11351 , \11352 , \11353 , \11354 ,
         \11355 , \11356 , \11357 , \11358 , \11359 , \11360 , \11361 , \11362 , \11363 , \11364 ,
         \11365 , \11366 , \11367 , \11368 , \11369 , \11370 , \11371 , \11372 , \11373 , \11374 ,
         \11375 , \11376 , \11377 , \11378 , \11379 , \11380 , \11381 , \11382 , \11383 , \11384 ,
         \11385 , \11386 , \11387 , \11388 , \11389 , \11390 , \11391 , \11392 , \11393 , \11394 ,
         \11395 , \11396 , \11397 , \11398 , \11399 , \11400 , \11401 , \11402 , \11403 , \11404 ,
         \11405 , \11406 , \11407 , \11408 , \11409 , \11410 , \11411 , \11412 , \11413 , \11414 ,
         \11415 , \11416 , \11417 , \11418 , \11419 , \11420 , \11421 , \11422 , \11423 , \11424 ,
         \11425 , \11426 , \11427 , \11428 , \11429 , \11430 , \11431 , \11432 , \11433 , \11434 ,
         \11435 , \11436 , \11437 , \11438 , \11439 , \11440 , \11441 , \11442 , \11443 , \11444 ,
         \11445 , \11446 , \11447 , \11448 , \11449 , \11450 , \11451 , \11452 , \11453 , \11454 ,
         \11455 , \11456 , \11457 , \11458 , \11459 , \11460 , \11461 , \11462 , \11463 , \11464 ,
         \11465 , \11466 , \11467 , \11468 , \11469 , \11470 , \11471 , \11472 , \11473 , \11474 ,
         \11475 , \11476 , \11477 , \11478 , \11479 , \11480 , \11481 , \11482 , \11483 , \11484 ,
         \11485 , \11486 , \11487 , \11488 , \11489 , \11490 , \11491 , \11492 , \11493 , \11494 ,
         \11495 , \11496 , \11497 , \11498 , \11499 , \11500 , \11501 , \11502 , \11503 , \11504 ,
         \11505 , \11506 , \11507 , \11508 , \11509 , \11510 , \11511 , \11512 , \11513 , \11514 ,
         \11515 , \11516 , \11517 , \11518 , \11519 , \11520 , \11521 , \11522 , \11523 , \11524 ,
         \11525 , \11526 , \11527 , \11528 , \11529 , \11530 , \11531 , \11532 , \11533 , \11534 ,
         \11535 , \11536 , \11537 , \11538 , \11539 , \11540 , \11541 , \11542 , \11543 , \11544 ,
         \11545 , \11546 , \11547 , \11548 , \11549 , \11550 , \11551 , \11552 , \11553 , \11554 ,
         \11555 , \11556 , \11557 , \11558 , \11559 , \11560 , \11561 , \11562 , \11563 , \11564 ,
         \11565 , \11566 , \11567 , \11568 , \11569 , \11570 , \11571 , \11572 , \11573 , \11574 ,
         \11575 , \11576 , \11577 , \11578 , \11579 , \11580 , \11581 , \11582 , \11583 , \11584 ,
         \11585 , \11586 , \11587 , \11588 , \11589 , \11590 , \11591 , \11592 , \11593 , \11594 ,
         \11595 , \11596 , \11597 , \11598 , \11599 , \11600 , \11601 , \11602 , \11603 , \11604 ,
         \11605 , \11606 , \11607 , \11608 , \11609 , \11610 , \11611 , \11612 , \11613 , \11614 ,
         \11615 , \11616 , \11617 , \11618 , \11619 , \11620 , \11621 , \11622 , \11623 , \11624 ,
         \11625 , \11626 , \11627 , \11628 , \11629 , \11630 , \11631 , \11632 , \11633 , \11634 ,
         \11635 , \11636 , \11637 , \11638 , \11639 , \11640 , \11641 , \11642 , \11643 , \11644 ,
         \11645 , \11646 , \11647 , \11648 , \11649 , \11650 , \11651 , \11652 , \11653 , \11654 ,
         \11655 , \11656 , \11657 , \11658 , \11659 , \11660 , \11661 , \11662 , \11663 , \11664 ,
         \11665 , \11666 , \11667 , \11668 , \11669 , \11670 , \11671 , \11672 , \11673 , \11674 ,
         \11675 , \11676 , \11677 , \11678 , \11679 , \11680 , \11681 , \11682 , \11683 , \11684 ,
         \11685 , \11686 , \11687 , \11688 , \11689 , \11690 , \11691 , \11692 , \11693 , \11694 ,
         \11695 , \11696 , \11697 , \11698 , \11699 , \11700 , \11701 , \11702 , \11703 , \11704 ,
         \11705 , \11706 , \11707 , \11708 , \11709 , \11710 , \11711 , \11712 , \11713 , \11714 ,
         \11715 , \11716 , \11717 , \11718 , \11719 , \11720 , \11721 , \11722 , \11723 , \11724 ,
         \11725 , \11726 , \11727 , \11728 , \11729 , \11730 , \11731 , \11732 , \11733 , \11734 ,
         \11735 , \11736 , \11737 , \11738 , \11739 , \11740 , \11741 , \11742 , \11743 , \11744 ,
         \11745 , \11746 , \11747 , \11748 , \11749 , \11750 , \11751 , \11752 , \11753 , \11754 ,
         \11755 , \11756 , \11757 , \11758 , \11759 , \11760 , \11761 , \11762 , \11763 , \11764 ,
         \11765 , \11766 , \11767 , \11768 , \11769 , \11770 , \11771 , \11772 , \11773 , \11774 ,
         \11775 , \11776 , \11777 , \11778 , \11779 , \11780 , \11781 , \11782 , \11783 , \11784 ,
         \11785 , \11786 , \11787 , \11788 , \11789 , \11790 , \11791 , \11792 , \11793 , \11794 ,
         \11795 , \11796 , \11797 , \11798 , \11799 , \11800 , \11801 , \11802 , \11803 , \11804 ,
         \11805 , \11806 , \11807 , \11808 , \11809 , \11810 , \11811 , \11812 , \11813 , \11814 ,
         \11815 , \11816 , \11817 , \11818 , \11819 , \11820 , \11821 , \11822 , \11823 , \11824 ,
         \11825 , \11826 , \11827 , \11828 , \11829 , \11830 , \11831 , \11832 , \11833 , \11834 ,
         \11835 , \11836 , \11837 , \11838 , \11839 , \11840 , \11841 , \11842 , \11843 , \11844 ,
         \11845 , \11846 , \11847 , \11848 , \11849 , \11850 , \11851 , \11852 , \11853 , \11854 ,
         \11855 , \11856 , \11857 , \11858 , \11859 , \11860 , \11861 , \11862 , \11863 , \11864 ,
         \11865 , \11866 , \11867 , \11868 , \11869 , \11870 , \11871 , \11872 , \11873 , \11874 ,
         \11875 , \11876 , \11877 , \11878 , \11879 , \11880 , \11881 , \11882 , \11883 , \11884 ,
         \11885 , \11886 , \11887 , \11888 , \11889 , \11890 , \11891 , \11892 , \11893 , \11894 ,
         \11895 , \11896 , \11897 , \11898 , \11899 , \11900 , \11901 , \11902 , \11903 , \11904 ,
         \11905 , \11906 , \11907 , \11908 , \11909 , \11910 , \11911 , \11912 , \11913 , \11914 ,
         \11915 , \11916 , \11917 , \11918 , \11919 , \11920 , \11921 , \11922 , \11923 , \11924 ,
         \11925 , \11926 , \11927 , \11928 , \11929 , \11930 , \11931 , \11932 , \11933 , \11934 ,
         \11935 , \11936 , \11937 , \11938 , \11939 , \11940 , \11941 , \11942 , \11943 , \11944 ,
         \11945 , \11946 , \11947 , \11948 , \11949 , \11950 , \11951 , \11952 , \11953 , \11954 ,
         \11955 , \11956 , \11957 , \11958 , \11959 , \11960 , \11961 , \11962 , \11963 , \11964 ,
         \11965 , \11966 , \11967 , \11968 , \11969 , \11970 , \11971 , \11972 , \11973 , \11974 ,
         \11975 , \11976 , \11977 , \11978 , \11979 , \11980 , \11981 , \11982 , \11983 , \11984 ,
         \11985 , \11986 , \11987 , \11988 , \11989 , \11990 , \11991 , \11992 , \11993 , \11994 ,
         \11995 , \11996 , \11997 , \11998 , \11999 , \12000 , \12001 , \12002 , \12003 , \12004 ,
         \12005 , \12006 , \12007 , \12008 , \12009 , \12010 , \12011 , \12012 , \12013 , \12014 ,
         \12015 , \12016 , \12017 , \12018 , \12019 , \12020 , \12021 , \12022 , \12023 , \12024 ,
         \12025 , \12026 , \12027 , \12028 , \12029 , \12030 , \12031 , \12032 , \12033 , \12034 ,
         \12035 , \12036 , \12037 , \12038 , \12039 , \12040 , \12041 , \12042 , \12043 , \12044 ,
         \12045 , \12046 , \12047 , \12048 , \12049 , \12050 , \12051 , \12052 , \12053 , \12054 ,
         \12055 , \12056 , \12057 , \12058 , \12059 , \12060 , \12061 , \12062 , \12063 , \12064 ,
         \12065 , \12066 , \12067 , \12068 , \12069 , \12070 , \12071 , \12072 , \12073 , \12074 ,
         \12075 , \12076 , \12077 , \12078 , \12079 , \12080 , \12081 , \12082 , \12083 , \12084 ,
         \12085 , \12086 , \12087 , \12088 , \12089 , \12090 , \12091 , \12092 , \12093 , \12094 ,
         \12095 , \12096 , \12097 , \12098 , \12099 , \12100 , \12101 , \12102 , \12103 , \12104 ,
         \12105 , \12106 , \12107 , \12108 , \12109 , \12110 , \12111 , \12112 , \12113 , \12114 ,
         \12115 , \12116 , \12117 , \12118 , \12119 , \12120 , \12121 , \12122 , \12123 , \12124 ,
         \12125 , \12126 , \12127 , \12128 , \12129 , \12130 , \12131 , \12132 , \12133 , \12134 ,
         \12135 , \12136 , \12137 , \12138 , \12139 , \12140 , \12141 , \12142 , \12143 , \12144 ,
         \12145 , \12146 , \12147 , \12148 , \12149 , \12150 , \12151 , \12152 , \12153 , \12154 ,
         \12155 , \12156 , \12157 , \12158 , \12159 , \12160 , \12161 , \12162 , \12163 , \12164 ,
         \12165 , \12166 , \12167 , \12168 , \12169 , \12170 , \12171 , \12172 , \12173 , \12174 ,
         \12175 , \12176 , \12177 , \12178 , \12179 , \12180 , \12181 , \12182 , \12183 , \12184 ,
         \12185 , \12186 , \12187 , \12188 , \12189 , \12190 , \12191 , \12192 , \12193 , \12194 ,
         \12195 , \12196 , \12197 , \12198 , \12199 , \12200 , \12201 , \12202 , \12203 , \12204 ,
         \12205 , \12206 , \12207 , \12208 , \12209 , \12210 , \12211 , \12212 , \12213 , \12214 ,
         \12215 , \12216 , \12217 , \12218 , \12219 , \12220 , \12221 , \12222 , \12223 , \12224 ,
         \12225 , \12226 , \12227 , \12228 , \12229 , \12230 , \12231 , \12232 , \12233 , \12234 ,
         \12235 , \12236 , \12237 , \12238 , \12239 , \12240 , \12241 , \12242 , \12243 , \12244 ,
         \12245 , \12246 , \12247 , \12248 , \12249 , \12250 , \12251 , \12252 , \12253 , \12254 ,
         \12255 , \12256 , \12257 , \12258 , \12259 , \12260 , \12261 , \12262 , \12263 , \12264 ,
         \12265 , \12266 , \12267 , \12268 , \12269 , \12270 , \12271 , \12272 , \12273 , \12274 ,
         \12275 , \12276 , \12277 , \12278 , \12279 , \12280 , \12281 , \12282 , \12283 , \12284 ,
         \12285 , \12286 , \12287 , \12288 , \12289 , \12290 , \12291 , \12292 , \12293 , \12294 ,
         \12295 , \12296 , \12297 , \12298 , \12299 , \12300 , \12301 , \12302 , \12303 , \12304 ,
         \12305 , \12306 , \12307 , \12308 , \12309 , \12310 , \12311 , \12312 , \12313 , \12314 ,
         \12315 , \12316 , \12317 , \12318 , \12319 , \12320 , \12321 , \12322 , \12323 , \12324 ,
         \12325 , \12326 , \12327 , \12328 , \12329 , \12330 , \12331 , \12332 , \12333 , \12334 ,
         \12335 , \12336 , \12337 , \12338 , \12339 , \12340 , \12341 , \12342 , \12343 , \12344 ,
         \12345 , \12346 , \12347 , \12348 , \12349 , \12350 , \12351 , \12352 , \12353 , \12354 ,
         \12355 , \12356 , \12357 , \12358 , \12359 , \12360 , \12361 , \12362 , \12363 , \12364 ,
         \12365 , \12366 , \12367 , \12368 , \12369 , \12370 , \12371 , \12372 , \12373 , \12374 ,
         \12375 , \12376 , \12377 , \12378 , \12379 , \12380 , \12381 , \12382 , \12383 , \12384 ,
         \12385 , \12386 , \12387 , \12388 , \12389 , \12390 , \12391 , \12392 , \12393 , \12394 ,
         \12395 , \12396 , \12397 , \12398 , \12399 , \12400 , \12401 , \12402 , \12403 , \12404 ,
         \12405 , \12406 , \12407 , \12408 , \12409 , \12410 , \12411 , \12412 , \12413 , \12414 ,
         \12415 , \12416 , \12417 , \12418 , \12419 , \12420 , \12421 , \12422 , \12423 , \12424 ,
         \12425 , \12426 , \12427 , \12428 , \12429 , \12430 , \12431 , \12432 , \12433 , \12434 ,
         \12435 , \12436 , \12437 , \12438 , \12439 , \12440 , \12441 , \12442 , \12443 , \12444 ,
         \12445 , \12446 , \12447 , \12448 , \12449 , \12450 , \12451 , \12452 , \12453 , \12454 ,
         \12455 , \12456 , \12457 , \12458 , \12459 , \12460 , \12461 , \12462 , \12463 , \12464 ,
         \12465 , \12466 , \12467 , \12468 , \12469 , \12470 , \12471 , \12472 , \12473 , \12474 ,
         \12475 , \12476 , \12477 , \12478 , \12479 , \12480 , \12481 , \12482 , \12483 , \12484 ,
         \12485 , \12486 , \12487 , \12488 , \12489 , \12490 , \12491 , \12492 , \12493 , \12494 ,
         \12495 , \12496 , \12497 , \12498 , \12499 , \12500 , \12501 , \12502 , \12503 , \12504 ,
         \12505 , \12506 , \12507 , \12508 , \12509 , \12510 , \12511 , \12512 , \12513 , \12514 ,
         \12515 , \12516 , \12517 , \12518 , \12519 , \12520 , \12521 , \12522 , \12523 , \12524 ,
         \12525 , \12526 , \12527 , \12528 , \12529 , \12530 , \12531 , \12532 , \12533 , \12534 ,
         \12535 , \12536 , \12537 , \12538 , \12539 , \12540 , \12541 , \12542 , \12543 , \12544 ,
         \12545 , \12546 , \12547 , \12548 , \12549 , \12550 , \12551 , \12552 , \12553 , \12554 ,
         \12555 , \12556 , \12557 , \12558 , \12559 , \12560 , \12561 , \12562 , \12563 , \12564 ,
         \12565 , \12566 , \12567 , \12568 , \12569 , \12570 , \12571 , \12572 , \12573 , \12574 ,
         \12575 , \12576 , \12577 , \12578 , \12579 , \12580 , \12581 , \12582 , \12583 , \12584 ,
         \12585 , \12586 , \12587 , \12588 , \12589 , \12590 , \12591 , \12592 , \12593 , \12594 ,
         \12595 , \12596 , \12597 , \12598 , \12599 , \12600 , \12601 , \12602 , \12603 , \12604 ,
         \12605 , \12606 , \12607 , \12608 , \12609 , \12610 , \12611 , \12612 , \12613 , \12614 ,
         \12615 , \12616 , \12617 , \12618 , \12619 , \12620 , \12621 , \12622 , \12623 , \12624 ,
         \12625 , \12626 , \12627 , \12628 , \12629 , \12630 , \12631 , \12632 , \12633 , \12634 ,
         \12635 , \12636 , \12637 , \12638 , \12639 , \12640 , \12641 , \12642 , \12643 , \12644 ,
         \12645 , \12646 , \12647 , \12648 , \12649 , \12650 , \12651 , \12652 , \12653 , \12654 ,
         \12655 , \12656 , \12657 , \12658 , \12659 , \12660 , \12661 , \12662 , \12663 , \12664 ,
         \12665 , \12666 , \12667 , \12668 , \12669 , \12670 , \12671 , \12672 , \12673 , \12674 ,
         \12675 , \12676 , \12677 , \12678 , \12679 , \12680 , \12681 , \12682 , \12683 , \12684 ,
         \12685 , \12686 , \12687 , \12688 , \12689 , \12690 , \12691 , \12692 , \12693 , \12694 ,
         \12695 , \12696 , \12697 , \12698 , \12699 , \12700 , \12701 , \12702 , \12703 , \12704 ,
         \12705 , \12706 , \12707 , \12708 , \12709 , \12710 , \12711 , \12712 , \12713 , \12714 ,
         \12715 , \12716 , \12717 , \12718 , \12719 , \12720 , \12721 , \12722 , \12723 , \12724 ,
         \12725 , \12726 , \12727 , \12728 , \12729 , \12730 , \12731 , \12732 , \12733 , \12734 ,
         \12735 , \12736 , \12737 , \12738 , \12739 , \12740 , \12741 , \12742 , \12743 , \12744 ,
         \12745 , \12746 , \12747 , \12748 , \12749 , \12750 , \12751 , \12752 , \12753 , \12754 ,
         \12755 , \12756 , \12757 , \12758 , \12759 , \12760 , \12761 , \12762 , \12763 , \12764 ,
         \12765 , \12766 , \12767 , \12768 , \12769 , \12770 , \12771 , \12772 , \12773 , \12774 ,
         \12775 , \12776 , \12777 , \12778 , \12779 , \12780 , \12781 , \12782 , \12783 , \12784 ,
         \12785 , \12786 , \12787 , \12788 , \12789 , \12790 , \12791 , \12792 , \12793 , \12794 ,
         \12795 , \12796 , \12797 , \12798 , \12799 , \12800 , \12801 , \12802 , \12803 , \12804 ,
         \12805 , \12806 , \12807 , \12808 , \12809 , \12810 , \12811 , \12812 , \12813 , \12814 ,
         \12815 , \12816 , \12817 , \12818 , \12819 , \12820 , \12821 , \12822 , \12823 , \12824 ,
         \12825 , \12826 , \12827 , \12828 , \12829 , \12830 , \12831 , \12832 , \12833 , \12834 ,
         \12835 , \12836 , \12837 , \12838 , \12839 , \12840 , \12841 , \12842 , \12843 , \12844 ,
         \12845 , \12846 , \12847 , \12848 , \12849 , \12850 , \12851 , \12852 , \12853 , \12854 ,
         \12855 , \12856 , \12857 , \12858 , \12859 , \12860 , \12861 , \12862 , \12863 , \12864 ,
         \12865 , \12866 , \12867 , \12868 , \12869 , \12870 , \12871 , \12872 , \12873 , \12874 ,
         \12875 , \12876 , \12877 , \12878 , \12879 , \12880 , \12881 , \12882 , \12883 , \12884 ,
         \12885 , \12886 , \12887 , \12888 , \12889 , \12890 , \12891 , \12892 , \12893 , \12894 ,
         \12895 , \12896 , \12897 , \12898 , \12899 , \12900 , \12901 , \12902 , \12903 , \12904 ,
         \12905 , \12906 , \12907 , \12908 , \12909 , \12910 , \12911 , \12912 , \12913 , \12914 ,
         \12915 , \12916 , \12917 , \12918 , \12919 , \12920 , \12921 , \12922 , \12923 , \12924 ,
         \12925 , \12926 , \12927 , \12928 , \12929 , \12930 , \12931 , \12932 , \12933 , \12934 ,
         \12935 , \12936 , \12937 , \12938 , \12939 , \12940 , \12941 , \12942 , \12943 , \12944 ,
         \12945 , \12946 , \12947 , \12948 , \12949 , \12950 , \12951 , \12952 , \12953 , \12954 ,
         \12955 , \12956 , \12957 , \12958 , \12959 , \12960 , \12961 , \12962 , \12963 , \12964 ,
         \12965 , \12966 , \12967 , \12968 , \12969 , \12970 , \12971 , \12972 , \12973 , \12974 ,
         \12975 , \12976 , \12977 , \12978 , \12979 , \12980 , \12981 , \12982 , \12983 , \12984 ,
         \12985 , \12986 , \12987 , \12988 , \12989 , \12990 , \12991 , \12992 , \12993 , \12994 ,
         \12995 , \12996 , \12997 , \12998 , \12999 , \13000 , \13001 , \13002 , \13003 , \13004 ,
         \13005 , \13006 , \13007 , \13008 , \13009 , \13010 , \13011 , \13012 , \13013 , \13014 ,
         \13015 , \13016 , \13017 , \13018 , \13019 , \13020 , \13021 , \13022 , \13023 , \13024 ,
         \13025 , \13026 , \13027 , \13028 , \13029 , \13030 , \13031 , \13032 , \13033 , \13034 ,
         \13035 , \13036 , \13037 , \13038 , \13039 , \13040 , \13041 , \13042 , \13043 , \13044 ,
         \13045 , \13046 , \13047 , \13048 , \13049 , \13050 , \13051 , \13052 , \13053 , \13054 ,
         \13055 , \13056 , \13057 , \13058 , \13059 , \13060 , \13061 , \13062 , \13063 , \13064 ,
         \13065 , \13066 , \13067 , \13068 , \13069 , \13070 , \13071 , \13072 , \13073 , \13074 ,
         \13075 , \13076 , \13077 , \13078 , \13079 , \13080 , \13081 , \13082 , \13083 , \13084 ,
         \13085 , \13086 , \13087 , \13088 , \13089 , \13090 , \13091 , \13092 , \13093 , \13094 ,
         \13095 , \13096 , \13097 , \13098 , \13099 , \13100 , \13101 , \13102 , \13103 , \13104 ,
         \13105 , \13106 , \13107 , \13108 , \13109 , \13110 , \13111 , \13112 , \13113 , \13114 ,
         \13115 , \13116 , \13117 , \13118 , \13119 , \13120 , \13121 , \13122 , \13123 , \13124 ,
         \13125 , \13126 , \13127 , \13128 , \13129 , \13130 , \13131 , \13132 , \13133 , \13134 ,
         \13135 , \13136 , \13137 , \13138 , \13139 , \13140 , \13141 , \13142 , \13143 , \13144 ,
         \13145 , \13146 , \13147 , \13148 , \13149 , \13150 , \13151 , \13152 , \13153 , \13154 ,
         \13155 , \13156 , \13157 , \13158 , \13159 , \13160 , \13161 , \13162 , \13163 , \13164 ,
         \13165 , \13166 , \13167 , \13168 , \13169 , \13170 , \13171 , \13172 , \13173 , \13174 ,
         \13175 , \13176 , \13177 , \13178 , \13179 , \13180 , \13181 , \13182 , \13183 , \13184 ,
         \13185 , \13186 , \13187 , \13188 , \13189 , \13190 , \13191 , \13192 , \13193 , \13194 ,
         \13195 , \13196 , \13197 , \13198 , \13199 , \13200 , \13201 , \13202 , \13203 , \13204 ,
         \13205 , \13206 , \13207 , \13208 , \13209 , \13210 , \13211 , \13212 , \13213 , \13214 ,
         \13215 , \13216 , \13217 , \13218 , \13219 , \13220 , \13221 , \13222 , \13223 , \13224 ,
         \13225 , \13226 , \13227 , \13228 , \13229 , \13230 , \13231 , \13232 , \13233 , \13234 ,
         \13235 , \13236 , \13237 , \13238 , \13239 , \13240 , \13241 , \13242 , \13243 , \13244 ,
         \13245 , \13246 , \13247 , \13248 , \13249 , \13250 , \13251 , \13252 , \13253 , \13254 ,
         \13255 , \13256 , \13257 , \13258 , \13259 , \13260 , \13261 , \13262 , \13263 , \13264 ,
         \13265 , \13266 , \13267 , \13268 , \13269 , \13270 , \13271 , \13272 , \13273 , \13274 ,
         \13275 , \13276 , \13277 , \13278 , \13279 , \13280 , \13281 , \13282 , \13283 , \13284 ,
         \13285 , \13286 , \13287 , \13288 , \13289 , \13290 , \13291 , \13292 , \13293 , \13294 ,
         \13295 , \13296 , \13297 , \13298 , \13299 , \13300 , \13301 , \13302 , \13303 , \13304 ,
         \13305 , \13306 , \13307 , \13308 , \13309 , \13310 , \13311 , \13312 , \13313 , \13314 ,
         \13315 , \13316 , \13317 , \13318 , \13319 , \13320 , \13321 , \13322 , \13323 , \13324 ,
         \13325 , \13326 , \13327 , \13328 , \13329 , \13330 , \13331 , \13332 , \13333 , \13334 ,
         \13335 , \13336 , \13337 , \13338 , \13339 , \13340 , \13341 , \13342 , \13343 , \13344 ,
         \13345 , \13346 , \13347 , \13348 , \13349 , \13350 , \13351 , \13352 , \13353 , \13354 ,
         \13355 , \13356 , \13357 , \13358 , \13359 , \13360 , \13361 , \13362 , \13363 , \13364 ,
         \13365 , \13366 , \13367 , \13368 , \13369 , \13370 , \13371 , \13372 , \13373 , \13374 ,
         \13375 , \13376 , \13377 , \13378 , \13379 , \13380 , \13381 , \13382 , \13383 , \13384 ,
         \13385 , \13386 , \13387 , \13388 , \13389 , \13390 , \13391 , \13392 , \13393 , \13394 ,
         \13395 , \13396 , \13397 , \13398 , \13399 , \13400 , \13401 , \13402 , \13403 , \13404 ,
         \13405 , \13406 , \13407 , \13408 , \13409 , \13410 , \13411 , \13412 , \13413 , \13414 ,
         \13415 , \13416 , \13417 , \13418 , \13419 , \13420 , \13421 , \13422 , \13423 , \13424 ,
         \13425 , \13426 , \13427 , \13428 , \13429 , \13430 , \13431 , \13432 , \13433 , \13434 ,
         \13435 , \13436 , \13437 , \13438 , \13439 , \13440 , \13441 , \13442 , \13443 , \13444 ,
         \13445 , \13446 , \13447 , \13448 , \13449 , \13450 , \13451 , \13452 , \13453 , \13454 ,
         \13455 , \13456 , \13457 , \13458 , \13459 , \13460 , \13461 , \13462 , \13463 , \13464 ,
         \13465 , \13466 , \13467 , \13468 , \13469 , \13470 , \13471 , \13472 , \13473 , \13474 ,
         \13475 , \13476 , \13477 , \13478 , \13479 , \13480 , \13481 , \13482 , \13483 , \13484 ,
         \13485 , \13486 , \13487 , \13488 , \13489 , \13490 , \13491 , \13492 , \13493 , \13494 ,
         \13495 , \13496 , \13497 , \13498 , \13499 , \13500 , \13501 , \13502 , \13503 , \13504 ,
         \13505 , \13506 , \13507 , \13508 , \13509 , \13510 , \13511 , \13512 , \13513 , \13514 ,
         \13515 , \13516 , \13517 , \13518 , \13519 , \13520 , \13521 , \13522 , \13523 , \13524 ,
         \13525 , \13526 , \13527 , \13528 , \13529 , \13530 , \13531 , \13532 , \13533 , \13534 ,
         \13535 , \13536 , \13537 , \13538 , \13539 , \13540 , \13541 , \13542 , \13543 , \13544 ,
         \13545 , \13546 , \13547 , \13548 , \13549 , \13550 , \13551 , \13552 , \13553 , \13554 ,
         \13555 , \13556 , \13557 , \13558 , \13559 , \13560 , \13561 , \13562 , \13563 , \13564 ,
         \13565 , \13566 , \13567 , \13568 , \13569 , \13570 , \13571 , \13572 , \13573 , \13574 ,
         \13575 , \13576 , \13577 , \13578 , \13579 , \13580 , \13581 , \13582 , \13583 , \13584 ,
         \13585 , \13586 , \13587 , \13588 , \13589 , \13590 , \13591 , \13592 , \13593 , \13594 ,
         \13595 , \13596 , \13597 , \13598 , \13599 , \13600 , \13601 , \13602 , \13603 , \13604 ,
         \13605 , \13606 , \13607 , \13608 , \13609 , \13610 , \13611 , \13612 , \13613 , \13614 ,
         \13615 , \13616 , \13617 , \13618 , \13619 , \13620 , \13621 , \13622 , \13623 , \13624 ,
         \13625 , \13626 , \13627 , \13628 , \13629 , \13630 , \13631 , \13632 , \13633 , \13634 ,
         \13635 , \13636 , \13637 , \13638 , \13639 , \13640 , \13641 , \13642 , \13643 , \13644 ,
         \13645 , \13646 , \13647 , \13648 , \13649 , \13650 , \13651 , \13652 , \13653 , \13654 ,
         \13655 , \13656 , \13657 , \13658 , \13659 , \13660 , \13661 , \13662 , \13663 , \13664 ,
         \13665 , \13666 , \13667 , \13668 , \13669 , \13670 , \13671 , \13672 , \13673 , \13674 ,
         \13675 , \13676 , \13677 , \13678 , \13679 , \13680 , \13681 , \13682 , \13683 , \13684 ,
         \13685 , \13686 , \13687 , \13688 , \13689 , \13690 , \13691 , \13692 , \13693 , \13694 ,
         \13695 , \13696 , \13697 , \13698 , \13699 , \13700 , \13701 , \13702 , \13703 , \13704 ,
         \13705 , \13706 , \13707 , \13708 , \13709 , \13710 , \13711 , \13712 , \13713 , \13714 ,
         \13715 , \13716 , \13717 , \13718 , \13719 , \13720 , \13721 , \13722 , \13723 , \13724 ,
         \13725 , \13726 , \13727 , \13728 , \13729 , \13730 , \13731 , \13732 , \13733 , \13734 ,
         \13735 , \13736 , \13737 , \13738 , \13739 , \13740 , \13741 , \13742 , \13743 , \13744 ,
         \13745 , \13746 , \13747 , \13748 , \13749 , \13750 , \13751 , \13752 , \13753 , \13754 ,
         \13755 , \13756 , \13757 , \13758 , \13759 , \13760 , \13761 , \13762 , \13763 , \13764 ,
         \13765 , \13766 , \13767 , \13768 , \13769 , \13770 , \13771 , \13772 , \13773 , \13774 ,
         \13775 , \13776 , \13777 , \13778 , \13779 , \13780 , \13781 , \13782 , \13783 , \13784 ,
         \13785 , \13786 , \13787 , \13788 , \13789 , \13790 , \13791 , \13792 , \13793 , \13794 ,
         \13795 , \13796 , \13797 , \13798 , \13799 , \13800 , \13801 , \13802 , \13803 , \13804 ,
         \13805 , \13806 , \13807 , \13808 , \13809 , \13810 , \13811 , \13812 , \13813 , \13814 ,
         \13815 , \13816 , \13817 , \13818 , \13819 , \13820 , \13821 , \13822 , \13823 , \13824 ,
         \13825 , \13826 , \13827 , \13828 , \13829 , \13830 , \13831 , \13832 , \13833 , \13834 ,
         \13835 , \13836 , \13837 , \13838 , \13839 , \13840 , \13841 , \13842 , \13843 , \13844 ,
         \13845 , \13846 , \13847 , \13848 , \13849 , \13850 , \13851 , \13852 , \13853 , \13854 ,
         \13855 , \13856 , \13857 , \13858 , \13859 , \13860 , \13861 , \13862 , \13863 , \13864 ,
         \13865 , \13866 , \13867 , \13868 , \13869 , \13870 , \13871 , \13872 , \13873 , \13874 ,
         \13875 , \13876 , \13877 , \13878 , \13879 , \13880 , \13881 , \13882 , \13883 , \13884 ,
         \13885 , \13886 , \13887 , \13888 , \13889 , \13890 , \13891 , \13892 , \13893 , \13894 ,
         \13895 , \13896 , \13897 , \13898 , \13899 , \13900 , \13901 , \13902 , \13903 , \13904 ,
         \13905 , \13906 , \13907 , \13908 , \13909 , \13910 , \13911 , \13912 , \13913 , \13914 ,
         \13915 , \13916 , \13917 , \13918 , \13919 , \13920 , \13921 , \13922 , \13923 , \13924 ,
         \13925 , \13926 , \13927 , \13928 , \13929 , \13930 , \13931 , \13932 , \13933 , \13934 ,
         \13935 , \13936 , \13937 , \13938 , \13939 , \13940 , \13941 , \13942 , \13943 , \13944 ,
         \13945 , \13946 , \13947 , \13948 , \13949 , \13950 , \13951 , \13952 , \13953 , \13954 ,
         \13955 , \13956 , \13957 , \13958 , \13959 , \13960 , \13961 , \13962 , \13963 , \13964 ,
         \13965 , \13966 , \13967 , \13968 , \13969 , \13970 , \13971 , \13972 , \13973 , \13974 ,
         \13975 , \13976 , \13977 , \13978 , \13979 , \13980 , \13981 , \13982 , \13983 , \13984 ,
         \13985 , \13986 , \13987 , \13988 , \13989 , \13990 , \13991 , \13992 , \13993 , \13994 ,
         \13995 , \13996 , \13997 , \13998 , \13999 , \14000 , \14001 , \14002 , \14003 , \14004 ,
         \14005 , \14006 , \14007 , \14008 , \14009 , \14010 , \14011 , \14012 , \14013 , \14014 ,
         \14015 , \14016 , \14017 , \14018 , \14019 , \14020 , \14021 , \14022 , \14023 , \14024 ,
         \14025 , \14026 , \14027 , \14028 , \14029 , \14030 , \14031 , \14032 , \14033 , \14034 ,
         \14035 , \14036 , \14037 , \14038 , \14039 , \14040 , \14041 , \14042 , \14043 , \14044 ,
         \14045 , \14046 , \14047 , \14048 , \14049 , \14050 , \14051 , \14052 , \14053 , \14054 ,
         \14055 , \14056 , \14057 , \14058 , \14059 , \14060 , \14061 , \14062 , \14063 , \14064 ,
         \14065 , \14066 , \14067 , \14068 , \14069 , \14070 , \14071 , \14072 , \14073 , \14074 ,
         \14075 , \14076 , \14077 , \14078 , \14079 , \14080 , \14081 , \14082 , \14083 , \14084 ,
         \14085 , \14086 , \14087 , \14088 , \14089 , \14090 , \14091 , \14092 , \14093 , \14094 ,
         \14095 , \14096 , \14097 , \14098 , \14099 , \14100 , \14101 , \14102 , \14103 , \14104 ,
         \14105 , \14106 , \14107 , \14108 , \14109 , \14110 , \14111 , \14112 , \14113 , \14114 ,
         \14115 , \14116 , \14117 , \14118 , \14119 , \14120 , \14121 , \14122 , \14123 , \14124 ,
         \14125 , \14126 , \14127 , \14128 , \14129 , \14130 , \14131 , \14132 , \14133 , \14134 ,
         \14135 , \14136 , \14137 , \14138 , \14139 , \14140 , \14141 , \14142 , \14143 , \14144 ,
         \14145 , \14146 , \14147 , \14148 , \14149 , \14150 , \14151 , \14152 , \14153 , \14154 ,
         \14155 , \14156 , \14157 , \14158 , \14159 , \14160 , \14161 , \14162 , \14163 , \14164 ,
         \14165 , \14166 , \14167 , \14168 , \14169 , \14170 , \14171 , \14172 , \14173 , \14174 ,
         \14175 , \14176 , \14177 , \14178 , \14179 , \14180 , \14181 , \14182 , \14183 , \14184 ,
         \14185 , \14186 , \14187 , \14188 , \14189 , \14190 , \14191 , \14192 , \14193 , \14194 ,
         \14195 , \14196 , \14197 , \14198 , \14199 , \14200 , \14201 , \14202 , \14203 , \14204 ,
         \14205 , \14206 , \14207 , \14208 , \14209 , \14210 , \14211 , \14212 , \14213 , \14214 ,
         \14215 , \14216 , \14217 , \14218 , \14219 , \14220 , \14221 , \14222 , \14223 , \14224 ,
         \14225 , \14226 , \14227 , \14228 , \14229 , \14230 , \14231 , \14232 , \14233 , \14234 ,
         \14235 , \14236 , \14237 , \14238 , \14239 , \14240 , \14241 , \14242 , \14243 , \14244 ,
         \14245 , \14246 , \14247 , \14248 , \14249 , \14250 , \14251 , \14252 , \14253 , \14254 ,
         \14255 , \14256 , \14257 , \14258 , \14259 , \14260 , \14261 , \14262 , \14263 , \14264 ,
         \14265 , \14266 , \14267 , \14268 , \14269 , \14270 , \14271 , \14272 , \14273 , \14274 ,
         \14275 , \14276 , \14277 , \14278 , \14279 , \14280 , \14281 , \14282 , \14283 , \14284 ,
         \14285 , \14286 , \14287 , \14288 , \14289 , \14290 , \14291 , \14292 , \14293 , \14294 ,
         \14295 , \14296 , \14297 , \14298 , \14299 , \14300 , \14301 , \14302 , \14303 , \14304 ,
         \14305 , \14306 , \14307 , \14308 , \14309 , \14310 , \14311 , \14312 , \14313 , \14314 ,
         \14315 , \14316 , \14317 , \14318 , \14319 , \14320 , \14321 , \14322 , \14323 , \14324 ,
         \14325 , \14326 , \14327 , \14328 , \14329 , \14330 , \14331 , \14332 , \14333 , \14334 ,
         \14335 , \14336 , \14337 , \14338 , \14339 , \14340 , \14341 , \14342 , \14343 , \14344 ,
         \14345 , \14346 , \14347 , \14348 , \14349 , \14350 , \14351 , \14352 , \14353 , \14354 ,
         \14355 , \14356 , \14357 , \14358 , \14359 , \14360 , \14361 , \14362 , \14363 , \14364 ,
         \14365 , \14366 , \14367 , \14368 , \14369 , \14370 , \14371 , \14372 , \14373 , \14374 ,
         \14375 , \14376 , \14377 , \14378 , \14379 , \14380 , \14381 , \14382 , \14383 , \14384 ,
         \14385 , \14386 , \14387 , \14388 , \14389 , \14390 , \14391 , \14392 , \14393 , \14394 ,
         \14395 , \14396 , \14397 , \14398 , \14399 , \14400 , \14401 , \14402 , \14403 , \14404 ,
         \14405 , \14406 , \14407 , \14408 , \14409 , \14410 , \14411 , \14412 , \14413 , \14414 ,
         \14415 , \14416 , \14417 , \14418 , \14419 , \14420 , \14421 , \14422 , \14423 , \14424 ,
         \14425 , \14426 , \14427 , \14428 , \14429 , \14430 , \14431 , \14432 , \14433 , \14434 ,
         \14435 , \14436 , \14437 , \14438 , \14439 , \14440 , \14441 , \14442 , \14443 , \14444 ,
         \14445 , \14446 , \14447 , \14448 , \14449 , \14450 , \14451 , \14452 , \14453 , \14454 ,
         \14455 , \14456 , \14457 , \14458 , \14459 , \14460 , \14461 , \14462 , \14463 , \14464 ,
         \14465 , \14466 , \14467 , \14468 , \14469 , \14470 , \14471 , \14472 , \14473 , \14474 ,
         \14475 , \14476 , \14477 , \14478 , \14479 , \14480 , \14481 , \14482 , \14483 , \14484 ,
         \14485 , \14486 , \14487 , \14488 , \14489 , \14490 , \14491 , \14492 , \14493 , \14494 ,
         \14495 , \14496 , \14497 , \14498 , \14499 , \14500 , \14501 , \14502 , \14503 , \14504 ,
         \14505 , \14506 , \14507 , \14508 , \14509 , \14510 , \14511 , \14512 , \14513 , \14514 ,
         \14515 , \14516 , \14517 , \14518 , \14519 , \14520 , \14521 , \14522 , \14523 , \14524 ,
         \14525 , \14526 , \14527 , \14528 , \14529 , \14530 , \14531 , \14532 , \14533 , \14534 ,
         \14535 , \14536 , \14537 , \14538 , \14539 , \14540 , \14541 , \14542 , \14543 , \14544 ,
         \14545 , \14546 , \14547 , \14548 , \14549 , \14550 , \14551 , \14552 , \14553 , \14554 ,
         \14555 , \14556 , \14557 , \14558 , \14559 , \14560 , \14561 , \14562 , \14563 , \14564 ,
         \14565 , \14566 , \14567 , \14568 , \14569 , \14570 , \14571 , \14572 , \14573 , \14574 ,
         \14575 , \14576 , \14577 , \14578 , \14579 , \14580 , \14581 , \14582 , \14583 , \14584 ,
         \14585 , \14586 , \14587 , \14588 , \14589 , \14590 , \14591 , \14592 , \14593 , \14594 ,
         \14595 , \14596 , \14597 , \14598 , \14599 , \14600 , \14601 , \14602 , \14603 , \14604 ,
         \14605 , \14606 , \14607 , \14608 , \14609 , \14610 , \14611 , \14612 , \14613 , \14614 ,
         \14615 , \14616 , \14617 , \14618 , \14619 , \14620 , \14621 , \14622 , \14623 , \14624 ,
         \14625 , \14626 , \14627 , \14628 , \14629 , \14630 , \14631 , \14632 , \14633 , \14634 ,
         \14635 , \14636 , \14637 , \14638 , \14639 , \14640 , \14641 , \14642 , \14643 , \14644 ,
         \14645 , \14646 , \14647 , \14648 , \14649 , \14650 , \14651 , \14652 , \14653 , \14654 ,
         \14655 , \14656 , \14657 , \14658 , \14659 , \14660 , \14661 , \14662 , \14663 , \14664 ,
         \14665 , \14666 , \14667 , \14668 , \14669 , \14670 , \14671 , \14672 , \14673 , \14674 ,
         \14675 , \14676 , \14677 , \14678 , \14679 , \14680 , \14681 , \14682 , \14683 , \14684 ,
         \14685 , \14686 , \14687 , \14688 , \14689 , \14690 , \14691 , \14692 , \14693 , \14694 ,
         \14695 , \14696 , \14697 , \14698 , \14699 , \14700 , \14701 , \14702 , \14703 , \14704 ,
         \14705 , \14706 , \14707 , \14708 , \14709 , \14710 , \14711 , \14712 , \14713 , \14714 ,
         \14715 , \14716 , \14717 , \14718 , \14719 , \14720 , \14721 , \14722 , \14723 , \14724 ,
         \14725 , \14726 , \14727 , \14728 , \14729 , \14730 , \14731 , \14732 , \14733 , \14734 ,
         \14735 , \14736 , \14737 , \14738 , \14739 , \14740 , \14741 , \14742 , \14743 , \14744 ,
         \14745 , \14746 , \14747 , \14748 , \14749 , \14750 , \14751 , \14752 , \14753 , \14754 ,
         \14755 , \14756 , \14757 , \14758 , \14759 , \14760 , \14761 , \14762 , \14763 , \14764 ,
         \14765 , \14766 , \14767 , \14768 , \14769 , \14770 , \14771 , \14772 , \14773 , \14774 ,
         \14775 , \14776 , \14777 , \14778 , \14779 , \14780 , \14781 , \14782 , \14783 , \14784 ,
         \14785 , \14786 , \14787 , \14788 , \14789 , \14790 , \14791 , \14792 , \14793 , \14794 ,
         \14795 , \14796 , \14797 , \14798 , \14799 , \14800 , \14801 , \14802 , \14803 , \14804 ,
         \14805 , \14806 , \14807 , \14808 , \14809 , \14810 , \14811 , \14812 , \14813 , \14814 ,
         \14815 , \14816 , \14817 , \14818 , \14819 , \14820 , \14821 , \14822 , \14823 , \14824 ,
         \14825 , \14826 , \14827 , \14828 , \14829 , \14830 , \14831 , \14832 , \14833 , \14834 ,
         \14835 , \14836 , \14837 , \14838 , \14839 , \14840 , \14841 , \14842 , \14843 , \14844 ,
         \14845 , \14846 , \14847 , \14848 , \14849 , \14850 , \14851 , \14852 , \14853 , \14854 ,
         \14855 , \14856 , \14857 , \14858 , \14859 , \14860 , \14861 , \14862 , \14863 , \14864 ,
         \14865 , \14866 , \14867 , \14868 , \14869 , \14870 , \14871 , \14872 , \14873 , \14874 ,
         \14875 , \14876 , \14877 , \14878 , \14879 , \14880 , \14881 , \14882 , \14883 , \14884 ,
         \14885 , \14886 , \14887 , \14888 , \14889 , \14890 , \14891 , \14892 , \14893 , \14894 ,
         \14895 , \14896 , \14897 , \14898 , \14899 , \14900 , \14901 , \14902 , \14903 , \14904 ,
         \14905 , \14906 , \14907 , \14908 , \14909 , \14910 , \14911 , \14912 , \14913 , \14914 ,
         \14915 , \14916 , \14917 , \14918 , \14919 , \14920 , \14921 , \14922 , \14923 , \14924 ,
         \14925 , \14926 , \14927 , \14928 , \14929 , \14930 , \14931 , \14932 , \14933 , \14934 ,
         \14935 , \14936 , \14937 , \14938 , \14939 , \14940 , \14941 , \14942 , \14943 , \14944 ,
         \14945 , \14946 , \14947 , \14948 , \14949 , \14950 , \14951 , \14952 , \14953 , \14954 ,
         \14955 , \14956 , \14957 , \14958 , \14959 , \14960 , \14961 , \14962 , \14963 , \14964 ,
         \14965 , \14966 , \14967 , \14968 , \14969 , \14970 , \14971 , \14972 , \14973 , \14974 ,
         \14975 , \14976 , \14977 , \14978 , \14979 , \14980 , \14981 , \14982 , \14983 , \14984 ,
         \14985 , \14986 , \14987 , \14988 , \14989 , \14990 , \14991 , \14992 , \14993 , \14994 ,
         \14995 , \14996 , \14997 , \14998 , \14999 , \15000 , \15001 , \15002 , \15003 , \15004 ,
         \15005 , \15006 , \15007 , \15008 , \15009 , \15010 , \15011 , \15012 , \15013 , \15014 ,
         \15015 , \15016 , \15017 , \15018 , \15019 , \15020 , \15021 , \15022 , \15023 , \15024 ,
         \15025 , \15026 , \15027 , \15028 , \15029 , \15030 , \15031 , \15032 , \15033 , \15034 ,
         \15035 , \15036 , \15037 , \15038 , \15039 , \15040 , \15041 , \15042 , \15043 , \15044 ,
         \15045 , \15046 , \15047 , \15048 , \15049 , \15050 , \15051 , \15052 , \15053 , \15054 ,
         \15055 , \15056 , \15057 , \15058 , \15059 , \15060 , \15061 , \15062 , \15063 , \15064 ,
         \15065 , \15066 , \15067 , \15068 , \15069 , \15070 , \15071 , \15072 , \15073 , \15074 ,
         \15075 , \15076 , \15077 , \15078 , \15079 , \15080 , \15081 , \15082 , \15083 , \15084 ,
         \15085 , \15086 , \15087 , \15088 , \15089 , \15090 , \15091 , \15092 , \15093 , \15094 ,
         \15095 , \15096 , \15097 , \15098 , \15099 , \15100 , \15101 , \15102 , \15103 , \15104 ,
         \15105 , \15106 , \15107 , \15108 , \15109 , \15110 , \15111 , \15112 , \15113 , \15114 ,
         \15115 , \15116 , \15117 , \15118 , \15119 , \15120 , \15121 , \15122 , \15123 , \15124 ,
         \15125 , \15126 , \15127 , \15128 , \15129 , \15130 , \15131 , \15132 , \15133 , \15134 ,
         \15135 , \15136 , \15137 , \15138 , \15139 , \15140 , \15141 , \15142 , \15143 , \15144 ,
         \15145 , \15146 , \15147 , \15148 , \15149 , \15150 , \15151 , \15152 , \15153 , \15154 ,
         \15155 , \15156 , \15157 , \15158 , \15159 , \15160 , \15161 , \15162 , \15163 , \15164 ,
         \15165 , \15166 , \15167 , \15168 , \15169 , \15170 , \15171 , \15172 , \15173 , \15174 ,
         \15175 , \15176 , \15177 , \15178 , \15179 , \15180 , \15181 , \15182 , \15183 , \15184 ,
         \15185 , \15186 , \15187 , \15188 , \15189 , \15190 , \15191 , \15192 , \15193 , \15194 ,
         \15195 , \15196 , \15197 , \15198 , \15199 , \15200 , \15201 , \15202 , \15203 , \15204 ,
         \15205 , \15206 , \15207 , \15208 , \15209 , \15210 , \15211 , \15212 , \15213 , \15214 ,
         \15215 , \15216 , \15217 , \15218 , \15219 , \15220 , \15221 , \15222 , \15223 , \15224 ,
         \15225 , \15226 , \15227 , \15228 , \15229 , \15230 , \15231 , \15232 , \15233 , \15234 ,
         \15235 , \15236 , \15237 , \15238 , \15239 , \15240 , \15241 , \15242 , \15243 , \15244 ,
         \15245 , \15246 , \15247 , \15248 , \15249 , \15250 , \15251 , \15252 , \15253 , \15254 ,
         \15255 , \15256 , \15257 , \15258 , \15259 , \15260 , \15261 , \15262 , \15263 , \15264 ,
         \15265 , \15266 , \15267 , \15268 , \15269 , \15270 , \15271 , \15272 , \15273 , \15274 ,
         \15275 , \15276 , \15277 , \15278 , \15279 , \15280 , \15281 , \15282 , \15283 , \15284 ,
         \15285 , \15286 , \15287 , \15288 , \15289 , \15290 , \15291 , \15292 , \15293 , \15294 ,
         \15295 , \15296 , \15297 , \15298 , \15299 , \15300 , \15301 , \15302 , \15303 , \15304 ,
         \15305 , \15306 , \15307 , \15308 , \15309 , \15310 , \15311 , \15312 , \15313 , \15314 ,
         \15315 , \15316 , \15317 , \15318 , \15319 , \15320 , \15321 , \15322 , \15323 , \15324 ,
         \15325 , \15326 , \15327 , \15328 , \15329 , \15330 , \15331 , \15332 , \15333 , \15334 ,
         \15335 , \15336 , \15337 , \15338 , \15339 , \15340 , \15341 , \15342 , \15343 , \15344 ,
         \15345 , \15346 , \15347 , \15348 , \15349 , \15350 , \15351 , \15352 , \15353 , \15354 ,
         \15355 , \15356 , \15357 , \15358 , \15359 , \15360 , \15361 , \15362 , \15363 , \15364 ,
         \15365 , \15366 , \15367 , \15368 , \15369 , \15370 , \15371 , \15372 , \15373 , \15374 ,
         \15375 , \15376 , \15377 , \15378 , \15379 , \15380 , \15381 , \15382 , \15383 , \15384 ,
         \15385 , \15386 , \15387 , \15388 , \15389 , \15390 , \15391 , \15392 , \15393 , \15394 ,
         \15395 , \15396 , \15397 , \15398 , \15399 , \15400 , \15401 , \15402 , \15403 , \15404 ,
         \15405 , \15406 , \15407 , \15408 , \15409 , \15410 , \15411 , \15412 , \15413 , \15414 ,
         \15415 , \15416 , \15417 , \15418 , \15419 , \15420 , \15421 , \15422 , \15423 , \15424 ,
         \15425 , \15426 , \15427 , \15428 , \15429 , \15430 , \15431 , \15432 , \15433 , \15434 ,
         \15435 , \15436 , \15437 , \15438 , \15439 , \15440 , \15441 , \15442 , \15443 , \15444 ,
         \15445 , \15446 , \15447 , \15448 , \15449 , \15450 , \15451 , \15452 , \15453 , \15454 ,
         \15455 , \15456 , \15457 , \15458 , \15459 , \15460 , \15461 , \15462 , \15463 , \15464 ,
         \15465 , \15466 , \15467 , \15468 , \15469 , \15470 , \15471 , \15472 , \15473 , \15474 ,
         \15475 , \15476 , \15477 , \15478 , \15479 , \15480 , \15481 , \15482 , \15483 , \15484 ,
         \15485 , \15486 , \15487 , \15488 , \15489 , \15490 , \15491 , \15492 , \15493 , \15494 ,
         \15495 , \15496 , \15497 , \15498 , \15499 , \15500 , \15501 , \15502 , \15503 , \15504 ,
         \15505 , \15506 , \15507 , \15508 , \15509 , \15510 , \15511 , \15512 , \15513 , \15514 ,
         \15515 , \15516 , \15517 , \15518 , \15519 , \15520 , \15521 , \15522 , \15523 , \15524 ,
         \15525 , \15526 , \15527 , \15528 , \15529 , \15530 , \15531 , \15532 , \15533 , \15534 ,
         \15535 , \15536 , \15537 , \15538 , \15539 , \15540 , \15541 , \15542 , \15543 , \15544 ,
         \15545 , \15546 , \15547 , \15548 , \15549 , \15550 , \15551 , \15552 , \15553 , \15554 ,
         \15555 , \15556 , \15557 , \15558 , \15559 , \15560 , \15561 , \15562 , \15563 , \15564 ,
         \15565 , \15566 , \15567 , \15568 , \15569 , \15570 , \15571 , \15572 , \15573 , \15574 ,
         \15575 , \15576 , \15577 , \15578 , \15579 , \15580 , \15581 , \15582 , \15583 , \15584 ,
         \15585 , \15586 , \15587 , \15588 , \15589 , \15590 , \15591 , \15592 , \15593 , \15594 ,
         \15595 , \15596 , \15597 , \15598 , \15599 , \15600 , \15601 , \15602 , \15603 , \15604 ,
         \15605 , \15606 , \15607 , \15608 , \15609 , \15610 , \15611 , \15612 , \15613 , \15614 ,
         \15615 , \15616 , \15617 , \15618 , \15619 , \15620 , \15621 , \15622 , \15623 , \15624 ,
         \15625 , \15626 , \15627 , \15628 , \15629 , \15630 , \15631 , \15632 , \15633 , \15634 ,
         \15635 , \15636 , \15637 , \15638 , \15639 , \15640 , \15641 , \15642 , \15643 , \15644 ,
         \15645 , \15646 , \15647 , \15648 , \15649 , \15650 , \15651 , \15652 , \15653 , \15654 ,
         \15655 , \15656 , \15657 , \15658 , \15659 , \15660 , \15661 , \15662 , \15663 , \15664 ,
         \15665 , \15666 , \15667 , \15668 , \15669 , \15670 , \15671 , \15672 , \15673 , \15674 ,
         \15675 , \15676 , \15677 , \15678 , \15679 , \15680 , \15681 , \15682 , \15683 , \15684 ,
         \15685 , \15686 , \15687 , \15688 , \15689 , \15690 , \15691 , \15692 , \15693 , \15694 ,
         \15695 , \15696 , \15697 , \15698 , \15699 , \15700 , \15701 , \15702 , \15703 , \15704 ,
         \15705 , \15706 , \15707 , \15708 , \15709 , \15710 , \15711 , \15712 , \15713 , \15714 ,
         \15715 , \15716 , \15717 , \15718 , \15719 , \15720 , \15721 , \15722 , \15723 , \15724 ,
         \15725 , \15726 , \15727 , \15728 , \15729 , \15730 , \15731 , \15732 , \15733 , \15734 ,
         \15735 , \15736 , \15737 , \15738 , \15739 , \15740 , \15741 , \15742 , \15743 , \15744 ,
         \15745 , \15746 , \15747 , \15748 , \15749 , \15750 , \15751 , \15752 , \15753 , \15754 ,
         \15755 , \15756 , \15757 , \15758 , \15759 , \15760 , \15761 , \15762 , \15763 , \15764 ,
         \15765 , \15766 , \15767 , \15768 , \15769 , \15770 , \15771 , \15772 , \15773 , \15774 ,
         \15775 , \15776 , \15777 , \15778 , \15779 , \15780 , \15781 , \15782 , \15783 , \15784 ,
         \15785 , \15786 , \15787 , \15788 , \15789 , \15790 , \15791 , \15792 , \15793 , \15794 ,
         \15795 , \15796 , \15797 , \15798 , \15799 , \15800 , \15801 , \15802 , \15803 , \15804 ,
         \15805 , \15806 , \15807 , \15808 , \15809 , \15810 , \15811 , \15812 , \15813 , \15814 ,
         \15815 , \15816 , \15817 , \15818 , \15819 , \15820 , \15821 , \15822 , \15823 , \15824 ,
         \15825 , \15826 , \15827 , \15828 , \15829 , \15830 , \15831 , \15832 , \15833 , \15834 ,
         \15835 , \15836 , \15837 , \15838 , \15839 , \15840 , \15841 , \15842 , \15843 , \15844 ,
         \15845 , \15846 , \15847 , \15848 , \15849 , \15850 , \15851 , \15852 , \15853 , \15854 ,
         \15855 , \15856 , \15857 , \15858 , \15859 , \15860 , \15861 , \15862 , \15863 , \15864 ,
         \15865 , \15866 , \15867 , \15868 , \15869 , \15870 , \15871 , \15872 , \15873 , \15874 ,
         \15875 , \15876 , \15877 , \15878 , \15879 , \15880 , \15881 , \15882 , \15883 , \15884 ,
         \15885 , \15886 , \15887 , \15888 , \15889 , \15890 , \15891 , \15892 , \15893 , \15894 ,
         \15895 , \15896 , \15897 , \15898 , \15899 , \15900 , \15901 , \15902 , \15903 , \15904 ,
         \15905 , \15906 , \15907 , \15908 , \15909 , \15910 , \15911 , \15912 , \15913 , \15914 ,
         \15915 , \15916 , \15917 , \15918 , \15919 , \15920 , \15921 , \15922 , \15923 , \15924 ,
         \15925 , \15926 , \15927 , \15928 , \15929 , \15930 , \15931 , \15932 , \15933 , \15934 ,
         \15935 , \15936 , \15937 , \15938 , \15939 , \15940 , \15941 , \15942 , \15943 , \15944 ,
         \15945 , \15946 , \15947 , \15948 , \15949 , \15950 , \15951 , \15952 , \15953 , \15954 ,
         \15955 , \15956 , \15957 , \15958 , \15959 , \15960 , \15961 , \15962 , \15963 , \15964 ,
         \15965 , \15966 , \15967 , \15968 , \15969 , \15970 , \15971 , \15972 , \15973 , \15974 ,
         \15975 , \15976 , \15977 , \15978 , \15979 , \15980 , \15981 , \15982 , \15983 , \15984 ,
         \15985 , \15986 , \15987 , \15988 , \15989 , \15990 , \15991 , \15992 , \15993 , \15994 ,
         \15995 , \15996 , \15997 , \15998 , \15999 , \16000 , \16001 , \16002 , \16003 , \16004 ,
         \16005 , \16006 , \16007 , \16008 , \16009 , \16010 , \16011 , \16012 , \16013 , \16014 ,
         \16015 , \16016 , \16017 , \16018 , \16019 , \16020 , \16021 , \16022 , \16023 , \16024 ,
         \16025 , \16026 , \16027 , \16028 , \16029 , \16030 , \16031 , \16032 , \16033 , \16034 ,
         \16035 , \16036 , \16037 , \16038 , \16039 , \16040 , \16041 , \16042 , \16043 , \16044 ,
         \16045 , \16046 , \16047 , \16048 , \16049 , \16050 , \16051 , \16052 , \16053 , \16054 ,
         \16055 , \16056 , \16057 , \16058 , \16059 , \16060 , \16061 , \16062 , \16063 , \16064 ,
         \16065 , \16066 , \16067 , \16068 , \16069 , \16070 , \16071 , \16072 , \16073 , \16074 ,
         \16075 , \16076 , \16077 , \16078 , \16079 , \16080 , \16081 , \16082 , \16083 , \16084 ,
         \16085 , \16086 , \16087 , \16088 , \16089 , \16090 , \16091 , \16092 , \16093 , \16094 ,
         \16095 , \16096 , \16097 , \16098 , \16099 , \16100 , \16101 , \16102 , \16103 , \16104 ,
         \16105 , \16106 , \16107 , \16108 , \16109 , \16110 , \16111 , \16112 , \16113 , \16114 ,
         \16115 , \16116 , \16117 , \16118 , \16119 , \16120 , \16121 , \16122 , \16123 , \16124 ,
         \16125 , \16126 , \16127 , \16128 , \16129 , \16130 , \16131 , \16132 , \16133 , \16134 ,
         \16135 , \16136 , \16137 , \16138 , \16139 , \16140 , \16141 , \16142 , \16143 , \16144 ,
         \16145 , \16146 , \16147 , \16148 , \16149 , \16150 , \16151 , \16152 , \16153 , \16154 ,
         \16155 , \16156 , \16157 , \16158 , \16159 , \16160 , \16161 , \16162 , \16163 , \16164 ,
         \16165 , \16166 , \16167 , \16168 , \16169 , \16170 , \16171 , \16172 , \16173 , \16174 ,
         \16175 , \16176 , \16177 , \16178 , \16179 , \16180 , \16181 , \16182 , \16183 , \16184 ,
         \16185 , \16186 , \16187 , \16188 , \16189 , \16190 , \16191 , \16192 , \16193 , \16194 ,
         \16195 , \16196 , \16197 , \16198 , \16199 , \16200 , \16201 , \16202 , \16203 , \16204 ,
         \16205 , \16206 , \16207 , \16208 , \16209 , \16210 , \16211 , \16212 , \16213 , \16214 ,
         \16215 , \16216 , \16217 , \16218 , \16219 , \16220 , \16221 , \16222 , \16223 , \16224 ,
         \16225 , \16226 , \16227 , \16228 , \16229 , \16230 , \16231 , \16232 , \16233 , \16234 ,
         \16235 , \16236 , \16237 , \16238 , \16239 , \16240 , \16241 , \16242 , \16243 , \16244 ,
         \16245 , \16246 , \16247 , \16248 , \16249 , \16250 , \16251 , \16252 , \16253 , \16254 ,
         \16255 , \16256 , \16257 , \16258 , \16259 , \16260 , \16261 , \16262 , \16263 , \16264 ,
         \16265 , \16266 , \16267 , \16268 , \16269 , \16270 , \16271 , \16272 , \16273 , \16274 ,
         \16275 , \16276 , \16277 , \16278 , \16279 , \16280 , \16281 , \16282 , \16283 , \16284 ,
         \16285 , \16286 , \16287 , \16288 , \16289 , \16290 , \16291 , \16292 , \16293 , \16294 ,
         \16295 , \16296 , \16297 , \16298 , \16299 , \16300 , \16301 , \16302 , \16303 , \16304 ,
         \16305 , \16306 , \16307 , \16308 , \16309 , \16310 , \16311 , \16312 , \16313 , \16314 ,
         \16315 , \16316 , \16317 , \16318 , \16319 , \16320 , \16321 , \16322 , \16323 , \16324 ,
         \16325 , \16326 , \16327 , \16328 , \16329 , \16330 , \16331 , \16332 , \16333 , \16334 ,
         \16335 , \16336 , \16337 , \16338 , \16339 , \16340 , \16341 , \16342 , \16343 , \16344 ,
         \16345 , \16346 , \16347 , \16348 , \16349 , \16350 , \16351 , \16352 , \16353 , \16354 ,
         \16355 , \16356 , \16357 , \16358 , \16359 , \16360 , \16361 , \16362 , \16363 , \16364 ,
         \16365 , \16366 , \16367 , \16368 , \16369 , \16370 , \16371 , \16372 , \16373 , \16374 ,
         \16375 , \16376 , \16377 , \16378 , \16379 , \16380 , \16381 , \16382 , \16383 , \16384 ,
         \16385 , \16386 , \16387 , \16388 , \16389 , \16390 , \16391 , \16392 , \16393 , \16394 ,
         \16395 , \16396 , \16397 , \16398 , \16399 , \16400 , \16401 , \16402 , \16403 , \16404 ,
         \16405 , \16406 , \16407 , \16408 , \16409 , \16410 , \16411 , \16412 , \16413 , \16414 ,
         \16415 , \16416 , \16417 , \16418 , \16419 , \16420 , \16421 , \16422 , \16423 , \16424 ,
         \16425 , \16426 , \16427 , \16428 , \16429 , \16430 , \16431 , \16432 , \16433 , \16434 ,
         \16435 , \16436 , \16437 , \16438 , \16439 , \16440 , \16441 , \16442 , \16443 , \16444 ,
         \16445 , \16446 , \16447 , \16448 , \16449 , \16450 , \16451 , \16452 , \16453 , \16454 ,
         \16455 , \16456 , \16457 , \16458 , \16459 , \16460 , \16461 , \16462 , \16463 , \16464 ,
         \16465 , \16466 , \16467 , \16468 , \16469 , \16470 , \16471 , \16472 , \16473 , \16474 ,
         \16475 , \16476 , \16477 , \16478 , \16479 , \16480 , \16481 , \16482 , \16483 , \16484 ,
         \16485 , \16486 , \16487 , \16488 , \16489 , \16490 , \16491 , \16492 , \16493 , \16494 ,
         \16495 , \16496 , \16497 , \16498 , \16499 , \16500 , \16501 , \16502 , \16503 , \16504 ,
         \16505 , \16506 , \16507 , \16508 , \16509 , \16510 , \16511 , \16512 , \16513 , \16514 ,
         \16515 , \16516 , \16517 , \16518 , \16519 , \16520 , \16521 , \16522 , \16523 , \16524 ,
         \16525 , \16526 , \16527 , \16528 , \16529 , \16530 , \16531 , \16532 , \16533 , \16534 ,
         \16535 , \16536 , \16537 , \16538 , \16539 , \16540 , \16541 , \16542 , \16543 , \16544 ,
         \16545 , \16546 , \16547 , \16548 , \16549 , \16550 , \16551 , \16552 , \16553 , \16554 ,
         \16555 , \16556 , \16557 , \16558 , \16559 , \16560 , \16561 , \16562 , \16563 , \16564 ,
         \16565 , \16566 , \16567 , \16568 , \16569 , \16570 , \16571 , \16572 , \16573 , \16574 ,
         \16575 , \16576 , \16577 , \16578 , \16579 , \16580 , \16581 , \16582 , \16583 , \16584 ,
         \16585 , \16586 , \16587 , \16588 , \16589 , \16590 , \16591 , \16592 , \16593 , \16594 ,
         \16595 , \16596 , \16597 , \16598 , \16599 , \16600 , \16601 , \16602 , \16603 , \16604 ,
         \16605 , \16606 , \16607 , \16608 , \16609 , \16610 , \16611 , \16612 , \16613 , \16614 ,
         \16615 , \16616 , \16617 , \16618 , \16619 , \16620 , \16621 , \16622 , \16623 , \16624 ,
         \16625 , \16626 , \16627 , \16628 , \16629 , \16630 , \16631 , \16632 , \16633 , \16634 ,
         \16635 , \16636 , \16637 , \16638 , \16639 , \16640 , \16641 , \16642 , \16643 , \16644 ,
         \16645 , \16646 , \16647 , \16648 , \16649 , \16650 , \16651 , \16652 , \16653 , \16654 ,
         \16655 , \16656 , \16657 , \16658 , \16659 , \16660 , \16661 , \16662 , \16663 , \16664 ,
         \16665 , \16666 , \16667 , \16668 , \16669 , \16670 , \16671 , \16672 , \16673 , \16674 ,
         \16675 , \16676 , \16677 , \16678 , \16679 , \16680 , \16681 , \16682 , \16683 , \16684 ,
         \16685 , \16686 , \16687 , \16688 , \16689 , \16690 , \16691 , \16692 , \16693 , \16694 ,
         \16695 , \16696 , \16697 , \16698 , \16699 , \16700 , \16701 , \16702 , \16703 , \16704 ,
         \16705 , \16706 , \16707 , \16708 , \16709 , \16710 , \16711 , \16712 , \16713 , \16714 ,
         \16715 , \16716 , \16717 , \16718 , \16719 , \16720 , \16721 , \16722 , \16723 , \16724 ,
         \16725 , \16726 , \16727 , \16728 , \16729 , \16730 , \16731 , \16732 , \16733 , \16734 ,
         \16735 , \16736 , \16737 , \16738 , \16739 , \16740 , \16741 , \16742 , \16743 , \16744 ,
         \16745 , \16746 , \16747 , \16748 , \16749 , \16750 , \16751 , \16752 , \16753 , \16754 ,
         \16755 , \16756 , \16757 , \16758 , \16759 , \16760 , \16761 , \16762 , \16763 , \16764 ,
         \16765 , \16766 , \16767 , \16768 , \16769 , \16770 , \16771 , \16772 , \16773 , \16774 ,
         \16775 , \16776 , \16777 , \16778 , \16779 , \16780 , \16781 , \16782 , \16783 , \16784 ,
         \16785 , \16786 , \16787 , \16788 , \16789 , \16790 , \16791 , \16792 , \16793 , \16794 ,
         \16795 , \16796 , \16797 , \16798 , \16799 , \16800 , \16801 , \16802 , \16803 , \16804 ,
         \16805 , \16806 , \16807 , \16808 , \16809 , \16810 , \16811 , \16812 , \16813 , \16814 ,
         \16815 , \16816 , \16817 , \16818 , \16819 , \16820 , \16821 , \16822 , \16823 , \16824 ,
         \16825 , \16826 , \16827 , \16828 , \16829 , \16830 , \16831 , \16832 , \16833 , \16834 ,
         \16835 , \16836 , \16837 , \16838 , \16839 , \16840 , \16841 , \16842 , \16843 , \16844 ,
         \16845 , \16846 , \16847 , \16848 , \16849 , \16850 , \16851 , \16852 , \16853 , \16854 ,
         \16855 , \16856 , \16857 , \16858 , \16859 , \16860 , \16861 , \16862 , \16863 , \16864 ,
         \16865 , \16866 , \16867 , \16868 , \16869 , \16870 , \16871 , \16872 , \16873 , \16874 ,
         \16875 , \16876 , \16877 , \16878 , \16879 , \16880 , \16881 , \16882 , \16883 , \16884 ,
         \16885 , \16886 , \16887 , \16888 , \16889 , \16890 , \16891 , \16892 , \16893 , \16894 ,
         \16895 , \16896 , \16897 , \16898 , \16899 , \16900 , \16901 , \16902 , \16903 , \16904 ,
         \16905 , \16906 , \16907 , \16908 , \16909 , \16910 , \16911 , \16912 , \16913 , \16914 ,
         \16915 , \16916 , \16917 , \16918 , \16919 , \16920 , \16921 , \16922 , \16923 , \16924 ,
         \16925 , \16926 , \16927 , \16928 , \16929 , \16930 , \16931 , \16932 , \16933 , \16934 ,
         \16935 , \16936 , \16937 , \16938 , \16939 , \16940 , \16941 , \16942 , \16943 , \16944 ,
         \16945 , \16946 , \16947 , \16948 , \16949 , \16950 , \16951 , \16952 , \16953 , \16954 ,
         \16955 , \16956 , \16957 , \16958 , \16959 , \16960 , \16961 , \16962 , \16963 , \16964 ,
         \16965 , \16966 , \16967 , \16968 , \16969 , \16970 , \16971 , \16972 , \16973 , \16974 ,
         \16975 , \16976 , \16977 , \16978 , \16979 , \16980 , \16981 , \16982 , \16983 , \16984 ,
         \16985 , \16986 , \16987 , \16988 , \16989 , \16990 , \16991 , \16992 , \16993 , \16994 ,
         \16995 , \16996 , \16997 , \16998 , \16999 , \17000 , \17001 , \17002 , \17003 , \17004 ,
         \17005 , \17006 , \17007 , \17008 , \17009 , \17010 , \17011 , \17012 , \17013 , \17014 ,
         \17015 , \17016 , \17017 , \17018 , \17019 , \17020 , \17021 , \17022 , \17023 , \17024 ,
         \17025 , \17026 , \17027 , \17028 , \17029 , \17030 , \17031 , \17032 , \17033 , \17034 ,
         \17035 , \17036 , \17037 , \17038 , \17039 , \17040 , \17041 , \17042 , \17043 , \17044 ,
         \17045 , \17046 , \17047 , \17048 , \17049 , \17050 , \17051 , \17052 , \17053 , \17054 ,
         \17055 , \17056 , \17057 , \17058 , \17059 , \17060 , \17061 , \17062 , \17063 , \17064 ,
         \17065 , \17066 , \17067 , \17068 , \17069 , \17070 , \17071 , \17072 , \17073 , \17074 ,
         \17075 , \17076 , \17077 , \17078 , \17079 , \17080 , \17081 , \17082 , \17083 , \17084 ,
         \17085 , \17086 , \17087 , \17088 , \17089 , \17090 , \17091 , \17092 , \17093 , \17094 ,
         \17095 , \17096 , \17097 , \17098 , \17099 , \17100 , \17101 , \17102 , \17103 , \17104 ,
         \17105 , \17106 , \17107 , \17108 , \17109 , \17110 , \17111 , \17112 , \17113 , \17114 ,
         \17115 , \17116 , \17117 , \17118 , \17119 , \17120 , \17121 , \17122 , \17123 , \17124 ,
         \17125 , \17126 , \17127 , \17128 , \17129 , \17130 , \17131 , \17132 , \17133 , \17134 ,
         \17135 , \17136 , \17137 , \17138 , \17139 , \17140 , \17141 , \17142 , \17143 , \17144 ,
         \17145 , \17146 , \17147 , \17148 , \17149 , \17150 , \17151 , \17152 , \17153 , \17154 ,
         \17155 , \17156 , \17157 , \17158 , \17159 , \17160 , \17161 , \17162 , \17163 , \17164 ,
         \17165 , \17166 , \17167 , \17168 , \17169 , \17170 , \17171 , \17172 , \17173 , \17174 ,
         \17175 , \17176 , \17177 , \17178 , \17179 , \17180 , \17181 , \17182 , \17183 , \17184 ,
         \17185 , \17186 , \17187 , \17188 , \17189 , \17190 , \17191 , \17192 , \17193 , \17194 ,
         \17195 , \17196 , \17197 , \17198 , \17199 , \17200 , \17201 , \17202 , \17203 , \17204 ,
         \17205 , \17206 , \17207 , \17208 , \17209 , \17210 , \17211 , \17212 , \17213 , \17214 ,
         \17215 , \17216 , \17217 , \17218 , \17219 , \17220 , \17221 , \17222 , \17223 , \17224 ,
         \17225 , \17226 , \17227 , \17228 , \17229 , \17230 , \17231 , \17232 , \17233 , \17234 ,
         \17235 , \17236 , \17237 , \17238 , \17239 , \17240 , \17241 , \17242 , \17243 , \17244 ,
         \17245 , \17246 , \17247 , \17248 , \17249 , \17250 , \17251 , \17252 , \17253 , \17254 ,
         \17255 , \17256 , \17257 , \17258 , \17259 , \17260 , \17261 , \17262 , \17263 , \17264 ,
         \17265 , \17266 , \17267 , \17268 , \17269 , \17270 , \17271 , \17272 , \17273 , \17274 ,
         \17275 , \17276 , \17277 , \17278 , \17279 , \17280 , \17281 , \17282 , \17283 , \17284 ,
         \17285 , \17286 , \17287 , \17288 , \17289 , \17290 , \17291 , \17292 , \17293 , \17294 ,
         \17295 , \17296 , \17297 , \17298 , \17299 , \17300 , \17301 , \17302 , \17303 , \17304 ,
         \17305 , \17306 , \17307 , \17308 , \17309 , \17310 , \17311 , \17312 , \17313 , \17314 ,
         \17315 , \17316 , \17317 , \17318 , \17319 , \17320 , \17321 , \17322 , \17323 , \17324 ,
         \17325 , \17326 , \17327 , \17328 , \17329 , \17330 , \17331 , \17332 , \17333 , \17334 ,
         \17335 , \17336 , \17337 , \17338 , \17339 , \17340 , \17341 , \17342 , \17343 , \17344 ,
         \17345 , \17346 , \17347 , \17348 , \17349 , \17350 , \17351 , \17352 , \17353 , \17354 ,
         \17355 , \17356 , \17357 , \17358 , \17359 , \17360 , \17361 , \17362 , \17363 , \17364 ,
         \17365 , \17366 , \17367 , \17368 , \17369 , \17370 , \17371 , \17372 , \17373 , \17374 ,
         \17375 , \17376 , \17377 , \17378 , \17379 , \17380 , \17381 , \17382 , \17383 , \17384 ,
         \17385 , \17386 , \17387 , \17388 , \17389 , \17390 , \17391 , \17392 , \17393 , \17394 ,
         \17395 , \17396 , \17397 , \17398 , \17399 , \17400 , \17401 , \17402 , \17403 , \17404 ,
         \17405 , \17406 , \17407 , \17408 , \17409 , \17410 , \17411 , \17412 , \17413 , \17414 ,
         \17415 , \17416 , \17417 , \17418 , \17419 , \17420 , \17421 , \17422 , \17423 , \17424 ,
         \17425 , \17426 , \17427 , \17428 , \17429 , \17430 , \17431 , \17432 , \17433 , \17434 ,
         \17435 , \17436 , \17437 , \17438 , \17439 , \17440 , \17441 , \17442 , \17443 , \17444 ,
         \17445 , \17446 , \17447 , \17448 , \17449 , \17450 , \17451 , \17452 , \17453 , \17454 ,
         \17455 , \17456 , \17457 , \17458 , \17459 , \17460 , \17461 , \17462 , \17463 , \17464 ,
         \17465 , \17466 , \17467 , \17468 , \17469 , \17470 , \17471 , \17472 , \17473 , \17474 ,
         \17475 , \17476 , \17477 , \17478 , \17479 , \17480 , \17481 , \17482 , \17483 , \17484 ,
         \17485 , \17486 , \17487 , \17488 , \17489 , \17490 , \17491 , \17492 , \17493 , \17494 ,
         \17495 , \17496 , \17497 , \17498 , \17499 , \17500 , \17501 , \17502 , \17503 , \17504 ,
         \17505 , \17506 , \17507 , \17508 , \17509 , \17510 , \17511 , \17512 , \17513 , \17514 ,
         \17515 , \17516 , \17517 , \17518 , \17519 , \17520 , \17521 , \17522 , \17523 , \17524 ,
         \17525 , \17526 , \17527 , \17528 , \17529 , \17530 , \17531 , \17532 , \17533 , \17534 ,
         \17535 , \17536 , \17537 , \17538 , \17539 , \17540 , \17541 , \17542 , \17543 , \17544 ,
         \17545 , \17546 , \17547 , \17548 , \17549 , \17550 , \17551 , \17552 , \17553 , \17554 ,
         \17555 , \17556 , \17557 , \17558 , \17559 , \17560 , \17561 , \17562 , \17563 , \17564 ,
         \17565 , \17566 , \17567 , \17568 , \17569 , \17570 , \17571 , \17572 , \17573 , \17574 ,
         \17575 , \17576 , \17577 , \17578 , \17579 , \17580 , \17581 , \17582 , \17583 , \17584 ,
         \17585 , \17586 , \17587 , \17588 , \17589 , \17590 , \17591 , \17592 , \17593 , \17594 ,
         \17595 , \17596 , \17597 , \17598 , \17599 , \17600 , \17601 , \17602 , \17603 , \17604 ,
         \17605 , \17606 , \17607 , \17608 , \17609 , \17610 , \17611 , \17612 , \17613 , \17614 ,
         \17615 , \17616 , \17617 , \17618 , \17619 , \17620 , \17621 , \17622 , \17623 , \17624 ,
         \17625 , \17626 , \17627 , \17628 , \17629 , \17630 , \17631 , \17632 , \17633 , \17634 ,
         \17635 , \17636 , \17637 , \17638 , \17639 , \17640 , \17641 , \17642 , \17643 , \17644 ,
         \17645 , \17646 , \17647 , \17648 , \17649 , \17650 , \17651 , \17652 , \17653 , \17654 ,
         \17655 , \17656 , \17657 , \17658 , \17659 , \17660 , \17661 , \17662 , \17663 , \17664 ,
         \17665 , \17666 , \17667 , \17668 , \17669 , \17670 , \17671 , \17672 , \17673 , \17674 ,
         \17675 , \17676 , \17677 , \17678 , \17679 , \17680 , \17681 , \17682 , \17683 , \17684 ,
         \17685 , \17686 , \17687 , \17688 , \17689 , \17690 , \17691 , \17692 , \17693 , \17694 ,
         \17695 , \17696 , \17697 , \17698 , \17699 , \17700 , \17701 , \17702 , \17703 , \17704 ,
         \17705 , \17706 , \17707 , \17708 , \17709 , \17710 , \17711 , \17712 , \17713 , \17714 ,
         \17715 , \17716 , \17717 , \17718 , \17719 , \17720 , \17721 , \17722 , \17723 , \17724 ,
         \17725 , \17726 , \17727 , \17728 , \17729 , \17730 , \17731 , \17732 , \17733 , \17734 ,
         \17735 , \17736 , \17737 , \17738 , \17739 , \17740 , \17741 , \17742 , \17743 , \17744 ,
         \17745 , \17746 , \17747 , \17748 , \17749 , \17750 , \17751 , \17752 , \17753 , \17754 ,
         \17755 , \17756 , \17757 , \17758 , \17759 , \17760 , \17761 , \17762 , \17763 , \17764 ,
         \17765 , \17766 , \17767 , \17768 , \17769 , \17770 , \17771 , \17772 , \17773 , \17774 ,
         \17775 , \17776 , \17777 , \17778 , \17779 , \17780 , \17781 , \17782 , \17783 , \17784 ,
         \17785 , \17786 , \17787 , \17788 , \17789 , \17790 , \17791 , \17792 , \17793 , \17794 ,
         \17795 , \17796 , \17797 , \17798 , \17799 , \17800 , \17801 , \17802 , \17803 , \17804 ,
         \17805 , \17806 , \17807 , \17808 , \17809 , \17810 , \17811 , \17812 , \17813 , \17814 ,
         \17815 , \17816 , \17817 , \17818 , \17819 , \17820 , \17821 , \17822 , \17823 , \17824 ,
         \17825 , \17826 , \17827 , \17828 , \17829 , \17830 , \17831 , \17832 , \17833 , \17834 ,
         \17835 , \17836 , \17837 , \17838 , \17839 , \17840 , \17841 , \17842 , \17843 , \17844 ,
         \17845 , \17846 , \17847 , \17848 , \17849 , \17850 , \17851 , \17852 , \17853 , \17854 ,
         \17855 , \17856 , \17857 , \17858 , \17859 , \17860 , \17861 , \17862 , \17863 , \17864 ,
         \17865 , \17866 , \17867 , \17868 , \17869 , \17870 , \17871 , \17872 , \17873 , \17874 ,
         \17875 , \17876 , \17877 , \17878 , \17879 , \17880 , \17881 , \17882 , \17883 , \17884 ,
         \17885 , \17886 , \17887 , \17888 , \17889 , \17890 , \17891 , \17892 , \17893 , \17894 ,
         \17895 , \17896 , \17897 , \17898 , \17899 , \17900 , \17901 , \17902 , \17903 , \17904 ,
         \17905 , \17906 , \17907 , \17908 , \17909 , \17910 , \17911 , \17912 , \17913 , \17914 ,
         \17915 , \17916 , \17917 , \17918 , \17919 , \17920 , \17921 , \17922 , \17923 , \17924 ,
         \17925 , \17926 , \17927 , \17928 , \17929 , \17930 , \17931 , \17932 , \17933 , \17934 ,
         \17935 , \17936 , \17937 , \17938 , \17939 , \17940 , \17941 , \17942 , \17943 , \17944 ,
         \17945 , \17946 , \17947 , \17948 , \17949 , \17950 , \17951 , \17952 , \17953 , \17954 ,
         \17955 , \17956 , \17957 , \17958 , \17959 , \17960 , \17961 , \17962 , \17963 , \17964 ,
         \17965 , \17966 , \17967 , \17968 , \17969 , \17970 , \17971 , \17972 , \17973 , \17974 ,
         \17975 , \17976 , \17977 , \17978 , \17979 , \17980 , \17981 , \17982 , \17983 , \17984 ,
         \17985 , \17986 , \17987 , \17988 , \17989 , \17990 , \17991 , \17992 , \17993 , \17994 ,
         \17995 , \17996 , \17997 , \17998 , \17999 , \18000 , \18001 , \18002 , \18003 , \18004 ,
         \18005 , \18006 , \18007 , \18008 , \18009 , \18010 , \18011 , \18012 , \18013 , \18014 ,
         \18015 , \18016 , \18017 , \18018 , \18019 , \18020 , \18021 , \18022 , \18023 , \18024 ,
         \18025 , \18026 , \18027 , \18028 , \18029 , \18030 , \18031 , \18032 , \18033 , \18034 ,
         \18035 , \18036 , \18037 , \18038 , \18039 , \18040 , \18041 , \18042 , \18043 , \18044 ,
         \18045 , \18046 , \18047 , \18048 , \18049 , \18050 , \18051 , \18052 , \18053 , \18054 ,
         \18055 , \18056 , \18057 , \18058 , \18059 , \18060 , \18061 , \18062 , \18063 , \18064 ,
         \18065 , \18066 , \18067 , \18068 , \18069 , \18070 , \18071 , \18072 , \18073 , \18074 ,
         \18075 , \18076 , \18077 , \18078 , \18079 , \18080 , \18081 , \18082 , \18083 , \18084 ,
         \18085 , \18086 , \18087 , \18088 , \18089 , \18090 , \18091 , \18092 , \18093 , \18094 ,
         \18095 , \18096 , \18097 , \18098 , \18099 , \18100 , \18101 , \18102 , \18103 , \18104 ,
         \18105 , \18106 , \18107 , \18108 , \18109 , \18110 , \18111 , \18112 , \18113 , \18114 ,
         \18115 , \18116 , \18117 , \18118 , \18119 , \18120 , \18121 , \18122 , \18123 , \18124 ,
         \18125 , \18126 , \18127 , \18128 , \18129 , \18130 , \18131 , \18132 , \18133 , \18134 ,
         \18135 , \18136 , \18137 , \18138 , \18139 , \18140 , \18141 , \18142 , \18143 , \18144 ,
         \18145 , \18146 , \18147 , \18148 , \18149 , \18150 , \18151 , \18152 , \18153 , \18154 ,
         \18155 , \18156 , \18157 , \18158 , \18159 , \18160 , \18161 , \18162 , \18163 , \18164 ,
         \18165 , \18166 , \18167 , \18168 , \18169 , \18170 , \18171 , \18172 , \18173 , \18174 ,
         \18175 , \18176 , \18177 , \18178 , \18179 , \18180 , \18181 , \18182 , \18183 , \18184 ,
         \18185 , \18186 , \18187 , \18188 , \18189 , \18190 , \18191 , \18192 , \18193 , \18194 ,
         \18195 , \18196 , \18197 , \18198 , \18199 , \18200 , \18201 , \18202 , \18203 , \18204 ,
         \18205 , \18206 , \18207 , \18208 , \18209 , \18210 , \18211 , \18212 , \18213 , \18214 ,
         \18215 , \18216 , \18217 , \18218 , \18219 , \18220 , \18221 , \18222 , \18223 , \18224 ,
         \18225 , \18226 , \18227 , \18228 , \18229 , \18230 , \18231 , \18232 , \18233 , \18234 ,
         \18235 , \18236 , \18237 , \18238 , \18239 , \18240 , \18241 , \18242 , \18243 , \18244 ,
         \18245 , \18246 , \18247 , \18248 , \18249 , \18250 , \18251 , \18252 , \18253 , \18254 ,
         \18255 , \18256 , \18257 , \18258 , \18259 , \18260 , \18261 , \18262 , \18263 , \18264 ,
         \18265 , \18266 , \18267 , \18268 , \18269 , \18270 , \18271 , \18272 , \18273 , \18274 ,
         \18275 , \18276 , \18277 , \18278 , \18279 , \18280 , \18281 , \18282 , \18283 , \18284 ,
         \18285 , \18286 , \18287 , \18288 , \18289 , \18290 , \18291 , \18292 , \18293 , \18294 ,
         \18295 , \18296 , \18297 , \18298 , \18299 , \18300 , \18301 , \18302 , \18303 , \18304 ,
         \18305 , \18306 , \18307 , \18308 , \18309 , \18310 , \18311 , \18312 , \18313 , \18314 ,
         \18315 , \18316 , \18317 , \18318 , \18319 , \18320 , \18321 , \18322 , \18323 , \18324 ,
         \18325 , \18326 , \18327 , \18328 , \18329 , \18330 , \18331 , \18332 , \18333 , \18334 ,
         \18335 , \18336 , \18337 , \18338 , \18339 , \18340 , \18341 , \18342 , \18343 , \18344 ,
         \18345 , \18346 , \18347 , \18348 , \18349 , \18350 , \18351 , \18352 , \18353 , \18354 ,
         \18355 , \18356 , \18357 , \18358 , \18359 , \18360 , \18361 , \18362 , \18363 , \18364 ,
         \18365 , \18366 , \18367 , \18368 , \18369 , \18370 , \18371 , \18372 , \18373 , \18374 ,
         \18375 , \18376 , \18377 , \18378 , \18379 , \18380 , \18381 , \18382 , \18383 , \18384 ,
         \18385 , \18386 , \18387 , \18388 , \18389 , \18390 , \18391 , \18392 , \18393 , \18394 ,
         \18395 , \18396 , \18397 , \18398 , \18399 , \18400 , \18401 , \18402 , \18403 , \18404 ,
         \18405 , \18406 , \18407 , \18408 , \18409 , \18410 , \18411 , \18412 , \18413 , \18414 ,
         \18415 , \18416 , \18417 , \18418 , \18419 , \18420 , \18421 , \18422 , \18423 , \18424 ,
         \18425 , \18426 , \18427 , \18428 , \18429 , \18430 , \18431 , \18432 , \18433 , \18434 ,
         \18435 , \18436 , \18437 , \18438 , \18439 , \18440 , \18441 , \18442 , \18443 , \18444 ,
         \18445 , \18446 , \18447 , \18448 , \18449 , \18450 , \18451 , \18452 , \18453 , \18454 ,
         \18455 , \18456 , \18457 , \18458 , \18459 , \18460 , \18461 , \18462 , \18463 , \18464 ,
         \18465 , \18466 , \18467 , \18468 , \18469 , \18470 , \18471 , \18472 , \18473 , \18474 ,
         \18475 , \18476 , \18477 , \18478 , \18479 , \18480 , \18481 , \18482 , \18483 , \18484 ,
         \18485 , \18486 , \18487 , \18488 , \18489 , \18490 , \18491 , \18492 , \18493 , \18494 ,
         \18495 , \18496 , \18497 , \18498 , \18499 , \18500 , \18501 , \18502 , \18503 , \18504 ,
         \18505 , \18506 , \18507 , \18508 , \18509 , \18510 , \18511 , \18512 , \18513 , \18514 ,
         \18515 , \18516 , \18517 , \18518 , \18519 , \18520 , \18521 , \18522 , \18523 , \18524 ,
         \18525 , \18526 , \18527 , \18528 , \18529 , \18530 , \18531 , \18532 , \18533 , \18534 ,
         \18535 , \18536 , \18537 , \18538 , \18539 , \18540 , \18541 , \18542 , \18543 , \18544 ,
         \18545 , \18546 , \18547 , \18548 , \18549 , \18550 , \18551 , \18552 , \18553 , \18554 ,
         \18555 , \18556 , \18557 , \18558 , \18559 , \18560 , \18561 , \18562 , \18563 , \18564 ,
         \18565 , \18566 , \18567 , \18568 , \18569 , \18570 , \18571 , \18572 , \18573 , \18574 ,
         \18575 , \18576 , \18577 , \18578 , \18579 , \18580 , \18581 , \18582 , \18583 , \18584 ,
         \18585 , \18586 , \18587 , \18588 , \18589 , \18590 , \18591 , \18592 , \18593 , \18594 ,
         \18595 , \18596 , \18597 , \18598 , \18599 , \18600 , \18601 , \18602 , \18603 , \18604 ,
         \18605 , \18606 , \18607 , \18608 , \18609 , \18610 , \18611 , \18612 , \18613 , \18614 ,
         \18615 , \18616 , \18617 , \18618 , \18619 , \18620 , \18621 , \18622 , \18623 , \18624 ,
         \18625 , \18626 , \18627 , \18628 , \18629 , \18630 , \18631 , \18632 , \18633 , \18634 ,
         \18635 , \18636 , \18637 , \18638 , \18639 , \18640 , \18641 , \18642 , \18643 , \18644 ,
         \18645 , \18646 , \18647 , \18648 , \18649 , \18650 , \18651 , \18652 , \18653 , \18654 ,
         \18655 , \18656 , \18657 , \18658 , \18659 , \18660 , \18661 , \18662 , \18663 , \18664 ,
         \18665 , \18666 , \18667 , \18668 , \18669 , \18670 , \18671 , \18672 , \18673 , \18674 ,
         \18675 , \18676 , \18677 , \18678 , \18679 , \18680 , \18681 , \18682 , \18683 , \18684 ,
         \18685 , \18686 , \18687 , \18688 , \18689 , \18690 , \18691 , \18692 , \18693 , \18694 ,
         \18695 , \18696 , \18697 , \18698 , \18699 , \18700 , \18701 , \18702 , \18703 , \18704 ,
         \18705 , \18706 , \18707 , \18708 , \18709 , \18710 , \18711 , \18712 , \18713 , \18714 ,
         \18715 , \18716 , \18717 , \18718 , \18719 , \18720 , \18721 , \18722 , \18723 , \18724 ,
         \18725 , \18726 , \18727 , \18728 , \18729 , \18730 , \18731 , \18732 , \18733 , \18734 ,
         \18735 , \18736 , \18737 , \18738 , \18739 , \18740 , \18741 , \18742 , \18743 , \18744 ,
         \18745 , \18746 , \18747 , \18748 , \18749 , \18750 , \18751 , \18752 , \18753 , \18754 ,
         \18755 , \18756 , \18757 , \18758 , \18759 , \18760 , \18761 , \18762 , \18763 , \18764 ,
         \18765 , \18766 , \18767 , \18768 , \18769 , \18770 , \18771 , \18772 , \18773 , \18774 ,
         \18775 , \18776 , \18777 , \18778 , \18779 , \18780 , \18781 , \18782 , \18783 , \18784 ,
         \18785 , \18786 , \18787 , \18788 , \18789 , \18790 , \18791 , \18792 , \18793 , \18794 ,
         \18795 , \18796 , \18797 , \18798 , \18799 , \18800 , \18801 , \18802 , \18803 , \18804 ,
         \18805 , \18806 , \18807 , \18808 , \18809 , \18810 , \18811 , \18812 , \18813 , \18814 ,
         \18815 , \18816 , \18817 , \18818 , \18819 , \18820 , \18821 , \18822 , \18823 , \18824 ,
         \18825 , \18826 , \18827 , \18828 , \18829 , \18830 , \18831 , \18832 , \18833 , \18834 ,
         \18835 , \18836 , \18837 , \18838 , \18839 , \18840 , \18841 , \18842 , \18843 , \18844 ,
         \18845 , \18846 , \18847 , \18848 , \18849 , \18850 , \18851 , \18852 , \18853 , \18854 ,
         \18855 , \18856 , \18857 , \18858 , \18859 , \18860 , \18861 , \18862 , \18863 , \18864 ,
         \18865 , \18866 , \18867 , \18868 , \18869 , \18870 , \18871 , \18872 , \18873 , \18874 ,
         \18875 , \18876 , \18877 , \18878 , \18879 , \18880 , \18881 , \18882 , \18883 , \18884 ,
         \18885 , \18886 , \18887 , \18888 , \18889 , \18890 , \18891 , \18892 , \18893 , \18894 ,
         \18895 , \18896 , \18897 , \18898 , \18899 , \18900 , \18901 , \18902 , \18903 , \18904 ,
         \18905 , \18906 , \18907 , \18908 , \18909 , \18910 , \18911 , \18912 , \18913 , \18914 ,
         \18915 , \18916 , \18917 , \18918 , \18919 , \18920 , \18921 , \18922 , \18923 , \18924 ,
         \18925 , \18926 , \18927 , \18928 , \18929 , \18930 , \18931 , \18932 , \18933 , \18934 ,
         \18935 , \18936 , \18937 , \18938 , \18939 , \18940 , \18941 , \18942 , \18943 , \18944 ,
         \18945 , \18946 , \18947 , \18948 , \18949 , \18950 , \18951 , \18952 , \18953 , \18954 ,
         \18955 , \18956 , \18957 , \18958 , \18959 , \18960 , \18961 , \18962 , \18963 , \18964 ,
         \18965 , \18966 , \18967 , \18968 , \18969 , \18970 , \18971 , \18972 , \18973 , \18974 ,
         \18975 , \18976 , \18977 , \18978 , \18979 , \18980 , \18981 , \18982 , \18983 , \18984 ,
         \18985 , \18986 , \18987 , \18988 , \18989 , \18990 , \18991 , \18992 , \18993 , \18994 ,
         \18995 , \18996 , \18997 , \18998 , \18999 , \19000 , \19001 , \19002 , \19003 , \19004 ,
         \19005 , \19006 , \19007 , \19008 , \19009 , \19010 , \19011 , \19012 , \19013 , \19014 ,
         \19015 , \19016 , \19017 , \19018 , \19019 , \19020 , \19021 , \19022 , \19023 , \19024 ,
         \19025 , \19026 , \19027 , \19028 , \19029 , \19030 , \19031 , \19032 , \19033 , \19034 ,
         \19035 , \19036 , \19037 , \19038 , \19039 , \19040 , \19041 , \19042 , \19043 , \19044 ,
         \19045 , \19046 , \19047 , \19048 , \19049 , \19050 , \19051 , \19052 , \19053 , \19054 ,
         \19055 , \19056 , \19057 , \19058 , \19059 , \19060 , \19061 , \19062 , \19063 , \19064 ,
         \19065 , \19066 , \19067 , \19068 , \19069 , \19070 , \19071 , \19072 , \19073 , \19074 ,
         \19075 , \19076 , \19077 , \19078 , \19079 , \19080 , \19081 , \19082 , \19083 , \19084 ,
         \19085 , \19086 , \19087 , \19088 , \19089 , \19090 , \19091 , \19092 , \19093 , \19094 ,
         \19095 , \19096 , \19097 , \19098 , \19099 , \19100 , \19101 , \19102 , \19103 , \19104 ,
         \19105 , \19106 , \19107 , \19108 , \19109 , \19110 , \19111 , \19112 , \19113 , \19114 ,
         \19115 , \19116 , \19117 , \19118 , \19119 , \19120 , \19121 , \19122 , \19123 , \19124 ,
         \19125 , \19126 , \19127 , \19128 , \19129 , \19130 , \19131 , \19132 , \19133 , \19134 ,
         \19135 , \19136 , \19137 , \19138 , \19139 , \19140 , \19141 , \19142 , \19143 , \19144 ,
         \19145 , \19146 , \19147 , \19148 , \19149 , \19150 , \19151 , \19152 , \19153 , \19154 ,
         \19155 , \19156 , \19157 , \19158 , \19159 , \19160 , \19161 , \19162 , \19163 , \19164 ,
         \19165 , \19166 , \19167 , \19168 , \19169 , \19170 , \19171 , \19172 , \19173 , \19174 ,
         \19175 , \19176 , \19177 , \19178 , \19179 , \19180 , \19181 , \19182 , \19183 , \19184 ,
         \19185 , \19186 , \19187 , \19188 , \19189 , \19190 , \19191 , \19192 , \19193 , \19194 ,
         \19195 , \19196 , \19197 , \19198 , \19199 , \19200 , \19201 , \19202 , \19203 , \19204 ,
         \19205 , \19206 , \19207 , \19208 , \19209 , \19210 , \19211 , \19212 , \19213 , \19214 ,
         \19215 , \19216 , \19217 , \19218 , \19219 , \19220 , \19221 , \19222 , \19223 , \19224 ,
         \19225 , \19226 , \19227 , \19228 , \19229 , \19230 , \19231 , \19232 , \19233 , \19234 ,
         \19235 , \19236 , \19237 , \19238 , \19239 , \19240 , \19241 , \19242 , \19243 , \19244 ,
         \19245 , \19246 , \19247 , \19248 , \19249 , \19250 , \19251 , \19252 , \19253 , \19254 ,
         \19255 , \19256 , \19257 , \19258 , \19259 , \19260 , \19261 , \19262 , \19263 , \19264 ,
         \19265 , \19266 , \19267 , \19268 , \19269 , \19270 , \19271 , \19272 , \19273 , \19274 ,
         \19275 , \19276 , \19277 , \19278 , \19279 , \19280 , \19281 , \19282 , \19283 , \19284 ,
         \19285 , \19286 , \19287 , \19288 , \19289 , \19290 , \19291 , \19292 , \19293 , \19294 ,
         \19295 , \19296 , \19297 , \19298 , \19299 , \19300 , \19301 , \19302 , \19303 , \19304 ,
         \19305 , \19306 , \19307 , \19308 , \19309 , \19310 , \19311 , \19312 , \19313 , \19314 ,
         \19315 , \19316 , \19317 , \19318 , \19319 , \19320 , \19321 , \19322 , \19323 , \19324 ,
         \19325 , \19326 , \19327 , \19328 , \19329 , \19330 , \19331 , \19332 , \19333 , \19334 ,
         \19335 , \19336 , \19337 , \19338 , \19339 , \19340 , \19341 , \19342 , \19343 , \19344 ,
         \19345 , \19346 , \19347 , \19348 , \19349 , \19350 , \19351 , \19352 , \19353 , \19354 ,
         \19355 , \19356 , \19357 , \19358 , \19359 , \19360 , \19361 , \19362 , \19363 , \19364 ,
         \19365 , \19366 , \19367 , \19368 , \19369 , \19370 , \19371 , \19372 , \19373 , \19374 ,
         \19375 , \19376 , \19377 , \19378 , \19379 , \19380 , \19381 , \19382 , \19383 , \19384 ,
         \19385 , \19386 , \19387 , \19388 , \19389 , \19390 , \19391 , \19392 , \19393 , \19394 ,
         \19395 , \19396 , \19397 , \19398 , \19399 , \19400 , \19401 , \19402 , \19403 , \19404 ,
         \19405 , \19406 , \19407 , \19408 , \19409 , \19410 , \19411 , \19412 , \19413 , \19414 ,
         \19415 , \19416 , \19417 , \19418 , \19419 , \19420 , \19421 , \19422 , \19423 , \19424 ,
         \19425 , \19426 , \19427 , \19428 , \19429 , \19430 , \19431 , \19432 , \19433 , \19434 ,
         \19435 , \19436 , \19437 , \19438 , \19439 , \19440 , \19441 , \19442 , \19443 , \19444 ,
         \19445 , \19446 , \19447 , \19448 , \19449 , \19450 , \19451 , \19452 , \19453 , \19454 ,
         \19455 , \19456 , \19457 , \19458 , \19459 , \19460 , \19461 , \19462 , \19463 , \19464 ,
         \19465 , \19466 , \19467 , \19468 , \19469 , \19470 , \19471 , \19472 , \19473 , \19474 ,
         \19475 , \19476 , \19477 , \19478 , \19479 , \19480 , \19481 , \19482 , \19483 , \19484 ,
         \19485 , \19486 , \19487 , \19488 , \19489 , \19490 , \19491 , \19492 , \19493 , \19494 ,
         \19495 , \19496 , \19497 , \19498 , \19499 , \19500 , \19501 , \19502 , \19503 , \19504 ,
         \19505 , \19506 , \19507 , \19508 , \19509 , \19510 , \19511 , \19512 , \19513 , \19514 ,
         \19515 , \19516 , \19517 , \19518 , \19519 , \19520 , \19521 , \19522 , \19523 , \19524 ,
         \19525 , \19526 , \19527 , \19528 , \19529 , \19530 , \19531 , \19532 , \19533 , \19534 ,
         \19535 , \19536 , \19537 , \19538 , \19539 , \19540 , \19541 , \19542 , \19543 , \19544 ,
         \19545 , \19546 , \19547 , \19548 , \19549 , \19550 , \19551 , \19552 , \19553 , \19554 ,
         \19555 , \19556 , \19557 , \19558 , \19559 , \19560 , \19561 , \19562 , \19563 , \19564 ,
         \19565 , \19566 , \19567 , \19568 , \19569 , \19570 , \19571 , \19572 , \19573 , \19574 ,
         \19575 , \19576 , \19577 , \19578 , \19579 , \19580 , \19581 , \19582 , \19583 , \19584 ,
         \19585 , \19586 , \19587 , \19588 , \19589 , \19590 , \19591 , \19592 , \19593 , \19594 ,
         \19595 , \19596 , \19597 , \19598 , \19599 , \19600 , \19601 , \19602 , \19603 , \19604 ,
         \19605 , \19606 , \19607 , \19608 , \19609 , \19610 , \19611 , \19612 , \19613 , \19614 ,
         \19615 , \19616 , \19617 , \19618 , \19619 , \19620 , \19621 , \19622 , \19623 , \19624 ,
         \19625 , \19626 , \19627 , \19628 , \19629 , \19630 , \19631 , \19632 , \19633 , \19634 ,
         \19635 , \19636 , \19637 , \19638 , \19639 , \19640 , \19641 , \19642 , \19643 , \19644 ,
         \19645 , \19646 , \19647 , \19648 , \19649 , \19650 , \19651 , \19652 , \19653 , \19654 ,
         \19655 , \19656 , \19657 , \19658 , \19659 , \19660 , \19661 , \19662 , \19663 , \19664 ,
         \19665 , \19666 , \19667 , \19668 , \19669 , \19670 , \19671 , \19672 , \19673 , \19674 ,
         \19675 , \19676 , \19677 , \19678 , \19679 , \19680 , \19681 , \19682 , \19683 , \19684 ,
         \19685 , \19686 , \19687 , \19688 , \19689 , \19690 , \19691 , \19692 , \19693 , \19694 ,
         \19695 , \19696 , \19697 , \19698 , \19699 , \19700 , \19701 , \19702 , \19703 , \19704 ,
         \19705 , \19706 , \19707 , \19708 , \19709 , \19710 , \19711 , \19712 , \19713 , \19714 ,
         \19715 , \19716 , \19717 , \19718 , \19719 , \19720 , \19721 , \19722 , \19723 , \19724 ,
         \19725 , \19726 , \19727 , \19728 , \19729 , \19730 , \19731 , \19732 , \19733 , \19734 ,
         \19735 , \19736 , \19737 , \19738 , \19739 , \19740 , \19741 , \19742 , \19743 , \19744 ,
         \19745 , \19746 , \19747 , \19748 , \19749 , \19750 , \19751 , \19752 , \19753 , \19754 ,
         \19755 , \19756 , \19757 , \19758 , \19759 , \19760 , \19761 , \19762 , \19763 , \19764 ,
         \19765 , \19766 , \19767 , \19768 , \19769 , \19770 , \19771 , \19772 , \19773 , \19774 ,
         \19775 , \19776 , \19777 , \19778 , \19779 , \19780 , \19781 , \19782 , \19783 , \19784 ,
         \19785 , \19786 , \19787 , \19788 , \19789 , \19790 , \19791 , \19792 , \19793 , \19794 ,
         \19795 , \19796 , \19797 , \19798 , \19799 , \19800 , \19801 , \19802 , \19803 , \19804 ,
         \19805 , \19806 , \19807 , \19808 , \19809 , \19810 , \19811 , \19812 , \19813 , \19814 ,
         \19815 , \19816 , \19817 , \19818 , \19819 , \19820 , \19821 , \19822 , \19823 , \19824 ,
         \19825 , \19826 , \19827 , \19828 , \19829 , \19830 , \19831 , \19832 , \19833 , \19834 ,
         \19835 , \19836 , \19837 , \19838 , \19839 , \19840 , \19841 , \19842 , \19843 , \19844 ,
         \19845 , \19846 , \19847 , \19848 , \19849 , \19850 , \19851 , \19852 , \19853 , \19854 ,
         \19855 , \19856 , \19857 , \19858 , \19859 , \19860 , \19861 , \19862 , \19863 , \19864 ,
         \19865 , \19866 , \19867 , \19868 , \19869 , \19870 , \19871 , \19872 , \19873 , \19874 ,
         \19875 , \19876 , \19877 , \19878 , \19879 , \19880 , \19881 , \19882 , \19883 , \19884 ,
         \19885 , \19886 , \19887 , \19888 , \19889 , \19890 , \19891 , \19892 , \19893 , \19894 ,
         \19895 , \19896 , \19897 , \19898 , \19899 , \19900 , \19901 , \19902 , \19903 , \19904 ,
         \19905 , \19906 , \19907 , \19908 , \19909 , \19910 , \19911 , \19912 , \19913 , \19914 ,
         \19915 , \19916 , \19917 , \19918 , \19919 , \19920 , \19921 , \19922 , \19923 , \19924 ,
         \19925 , \19926 , \19927 , \19928 , \19929 , \19930 , \19931 , \19932 , \19933 , \19934 ,
         \19935 , \19936 , \19937 , \19938 , \19939 , \19940 , \19941 , \19942 , \19943 , \19944 ,
         \19945 , \19946 , \19947 , \19948 , \19949 , \19950 , \19951 , \19952 , \19953 , \19954 ,
         \19955 , \19956 , \19957 , \19958 , \19959 , \19960 , \19961 , \19962 , \19963 , \19964 ,
         \19965 , \19966 , \19967 , \19968 , \19969 , \19970 , \19971 , \19972 , \19973 , \19974 ,
         \19975 , \19976 , \19977 , \19978 , \19979 , \19980 , \19981 , \19982 , \19983 , \19984 ,
         \19985 , \19986 , \19987 , \19988 , \19989 , \19990 , \19991 , \19992 , \19993 , \19994 ,
         \19995 , \19996 , \19997 , \19998 , \19999 , \20000 , \20001 , \20002 , \20003 , \20004 ,
         \20005 , \20006 , \20007 , \20008 , \20009 , \20010 , \20011 , \20012 , \20013 , \20014 ,
         \20015 , \20016 , \20017 , \20018 , \20019 , \20020 , \20021 , \20022 , \20023 , \20024 ,
         \20025 , \20026 , \20027 , \20028 , \20029 , \20030 , \20031 , \20032 , \20033 , \20034 ,
         \20035 , \20036 , \20037 , \20038 , \20039 , \20040 , \20041 , \20042 , \20043 , \20044 ,
         \20045 , \20046 , \20047 , \20048 , \20049 , \20050 , \20051 , \20052 , \20053 , \20054 ,
         \20055 , \20056 , \20057 , \20058 , \20059 , \20060 , \20061 , \20062 , \20063 , \20064 ,
         \20065 , \20066 , \20067 , \20068 , \20069 , \20070 , \20071 , \20072 , \20073 , \20074 ,
         \20075 , \20076 , \20077 , \20078 , \20079 , \20080 , \20081 , \20082 , \20083 , \20084 ,
         \20085 , \20086 , \20087 , \20088 , \20089 , \20090 , \20091 , \20092 , \20093 , \20094 ,
         \20095 , \20096 , \20097 , \20098 , \20099 , \20100 , \20101 , \20102 , \20103 , \20104 ,
         \20105 , \20106 , \20107 , \20108 , \20109 , \20110 , \20111 , \20112 , \20113 , \20114 ,
         \20115 , \20116 , \20117 , \20118 , \20119 , \20120 , \20121 , \20122 , \20123 , \20124 ,
         \20125 , \20126 , \20127 , \20128 , \20129 , \20130 , \20131 , \20132 , \20133 , \20134 ,
         \20135 , \20136 , \20137 , \20138 , \20139 , \20140 , \20141 , \20142 , \20143 , \20144 ,
         \20145 , \20146 , \20147 , \20148 , \20149 , \20150 , \20151 , \20152 , \20153 , \20154 ,
         \20155 , \20156 , \20157 , \20158 , \20159 , \20160 , \20161 , \20162 , \20163 , \20164 ,
         \20165 , \20166 , \20167 , \20168 , \20169 , \20170 , \20171 , \20172 , \20173 , \20174 ,
         \20175 , \20176 , \20177 , \20178 , \20179 , \20180 , \20181 , \20182 , \20183 , \20184 ,
         \20185 , \20186 , \20187 , \20188 , \20189 , \20190 , \20191 , \20192 , \20193 , \20194 ,
         \20195 , \20196 , \20197 , \20198 , \20199 , \20200 , \20201 , \20202 , \20203 , \20204 ,
         \20205 , \20206 , \20207 , \20208 , \20209 , \20210 , \20211 , \20212 , \20213 , \20214 ,
         \20215 , \20216 , \20217 , \20218 , \20219 , \20220 , \20221 , \20222 , \20223 , \20224 ,
         \20225 , \20226 , \20227 , \20228 , \20229 , \20230 , \20231 , \20232 , \20233 , \20234 ,
         \20235 , \20236 , \20237 , \20238 , \20239 , \20240 , \20241 , \20242 , \20243 , \20244 ,
         \20245 , \20246 , \20247 , \20248 , \20249 , \20250 , \20251 , \20252 , \20253 , \20254 ,
         \20255 , \20256 , \20257 , \20258 , \20259 , \20260 , \20261 , \20262 , \20263 , \20264 ,
         \20265 , \20266 , \20267 , \20268 , \20269 , \20270 , \20271 , \20272 , \20273 , \20274 ,
         \20275 , \20276 , \20277 , \20278 , \20279 , \20280 , \20281 , \20282 , \20283 , \20284 ,
         \20285 , \20286 , \20287 , \20288 , \20289 , \20290 , \20291 , \20292 , \20293 , \20294 ,
         \20295 , \20296 , \20297 , \20298 , \20299 , \20300 , \20301 , \20302 , \20303 , \20304 ,
         \20305 , \20306 , \20307 , \20308 , \20309 , \20310 , \20311 , \20312 , \20313 , \20314 ,
         \20315 , \20316 , \20317 , \20318 , \20319 , \20320 , \20321 , \20322 , \20323 , \20324 ,
         \20325 , \20326 , \20327 , \20328 , \20329 , \20330 , \20331 , \20332 , \20333 , \20334 ,
         \20335 , \20336 , \20337 , \20338 , \20339 , \20340 , \20341 , \20342 , \20343 , \20344 ,
         \20345 , \20346 , \20347 , \20348 , \20349 , \20350 , \20351 , \20352 , \20353 , \20354 ,
         \20355 , \20356 , \20357 , \20358 , \20359 , \20360 , \20361 , \20362 , \20363 , \20364 ,
         \20365 , \20366 , \20367 , \20368 , \20369 , \20370 , \20371 , \20372 , \20373 , \20374 ,
         \20375 , \20376 , \20377 , \20378 , \20379 , \20380 , \20381 , \20382 , \20383 , \20384 ,
         \20385 , \20386 , \20387 , \20388 , \20389 , \20390 , \20391 , \20392 , \20393 , \20394 ,
         \20395 , \20396 , \20397 , \20398 , \20399 , \20400 , \20401 , \20402 , \20403 , \20404 ,
         \20405 , \20406 , \20407 , \20408 , \20409 , \20410 , \20411 , \20412 , \20413 , \20414 ,
         \20415 , \20416 , \20417 , \20418 , \20419 , \20420 , \20421 , \20422 , \20423 , \20424 ,
         \20425 , \20426 , \20427 , \20428 , \20429 , \20430 , \20431 , \20432 , \20433 , \20434 ,
         \20435 , \20436 , \20437 , \20438 , \20439 , \20440 , \20441 , \20442 , \20443 , \20444 ,
         \20445 , \20446 , \20447 , \20448 , \20449 , \20450 , \20451 , \20452 , \20453 , \20454 ,
         \20455 , \20456 , \20457 , \20458 , \20459 , \20460 , \20461 , \20462 , \20463 , \20464 ,
         \20465 , \20466 , \20467 , \20468 , \20469 , \20470 , \20471 , \20472 , \20473 , \20474 ,
         \20475 , \20476 , \20477 , \20478 , \20479 , \20480 , \20481 , \20482 , \20483 , \20484 ,
         \20485 , \20486 , \20487 , \20488 , \20489 , \20490 , \20491 , \20492 , \20493 , \20494 ,
         \20495 , \20496 , \20497 , \20498 , \20499 , \20500 , \20501 , \20502 , \20503 , \20504 ,
         \20505 , \20506 , \20507 , \20508 , \20509 , \20510 , \20511 , \20512 , \20513 , \20514 ,
         \20515 , \20516 , \20517 , \20518 , \20519 , \20520 , \20521 , \20522 , \20523 , \20524 ,
         \20525 , \20526 , \20527 , \20528 , \20529 , \20530 , \20531 , \20532 , \20533 , \20534 ,
         \20535 , \20536 , \20537 , \20538 , \20539 , \20540 , \20541 , \20542 , \20543 , \20544 ,
         \20545 , \20546 , \20547 , \20548 , \20549 , \20550 , \20551 , \20552 , \20553 , \20554 ,
         \20555 , \20556 , \20557 , \20558 , \20559 , \20560 , \20561 , \20562 , \20563 , \20564 ,
         \20565 , \20566 , \20567 , \20568 , \20569 , \20570 , \20571 , \20572 , \20573 , \20574 ,
         \20575 , \20576 , \20577 , \20578 , \20579 , \20580 , \20581 , \20582 , \20583 , \20584 ,
         \20585 , \20586 , \20587 , \20588 , \20589 , \20590 , \20591 , \20592 , \20593 , \20594 ,
         \20595 , \20596 , \20597 , \20598 , \20599 , \20600 , \20601 , \20602 , \20603 , \20604 ,
         \20605 , \20606 , \20607 , \20608 , \20609 , \20610 , \20611 , \20612 , \20613 , \20614 ,
         \20615 , \20616 , \20617 , \20618 , \20619 , \20620 , \20621 , \20622 , \20623 , \20624 ,
         \20625 , \20626 , \20627 , \20628 , \20629 , \20630 , \20631 , \20632 , \20633 , \20634 ,
         \20635 , \20636 , \20637 , \20638 , \20639 , \20640 , \20641 , \20642 , \20643 , \20644 ,
         \20645 , \20646 , \20647 , \20648 , \20649 , \20650 , \20651 , \20652 , \20653 , \20654 ,
         \20655 , \20656 , \20657 , \20658 , \20659 , \20660 , \20661 , \20662 , \20663 , \20664 ,
         \20665 , \20666 , \20667 , \20668 , \20669 , \20670 , \20671 , \20672 , \20673 , \20674 ,
         \20675 , \20676 , \20677 , \20678 , \20679 , \20680 , \20681 , \20682 , \20683 , \20684 ,
         \20685 , \20686 , \20687 , \20688 , \20689 , \20690 , \20691 , \20692 , \20693 , \20694 ,
         \20695 , \20696 , \20697 , \20698 , \20699 , \20700 , \20701 , \20702 , \20703 , \20704 ,
         \20705 , \20706 , \20707 , \20708 , \20709 , \20710 , \20711 , \20712 , \20713 , \20714 ,
         \20715 , \20716 , \20717 , \20718 , \20719 , \20720 , \20721 , \20722 , \20723 , \20724 ,
         \20725 , \20726 , \20727 , \20728 , \20729 , \20730 , \20731 , \20732 , \20733 , \20734 ,
         \20735 , \20736 , \20737 , \20738 , \20739 , \20740 , \20741 , \20742 , \20743 , \20744 ,
         \20745 , \20746 , \20747 , \20748 , \20749 , \20750 , \20751 , \20752 , \20753 , \20754 ,
         \20755 , \20756 , \20757 , \20758 , \20759 , \20760 , \20761 , \20762 , \20763 , \20764 ,
         \20765 , \20766 , \20767 , \20768 , \20769 , \20770 , \20771 , \20772 , \20773 , \20774 ,
         \20775 , \20776 , \20777 , \20778 , \20779 , \20780 , \20781 , \20782 , \20783 , \20784 ,
         \20785 , \20786 , \20787 , \20788 , \20789 , \20790 , \20791 , \20792 , \20793 , \20794 ,
         \20795 , \20796 , \20797 , \20798 , \20799 , \20800 , \20801 , \20802 , \20803 , \20804 ,
         \20805 , \20806 , \20807 , \20808 , \20809 , \20810 , \20811 , \20812 , \20813 , \20814 ,
         \20815 , \20816 , \20817 , \20818 , \20819 , \20820 , \20821 , \20822 , \20823 , \20824 ,
         \20825 , \20826 , \20827 , \20828 , \20829 , \20830 , \20831 , \20832 , \20833 , \20834 ,
         \20835 , \20836 , \20837 , \20838 , \20839 , \20840 , \20841 , \20842 , \20843 , \20844 ,
         \20845 , \20846 , \20847 , \20848 , \20849 , \20850 , \20851 , \20852 , \20853 , \20854 ,
         \20855 , \20856 , \20857 , \20858 , \20859 , \20860 , \20861 , \20862 , \20863 , \20864 ,
         \20865 , \20866 , \20867 , \20868 , \20869 , \20870 , \20871 , \20872 , \20873 , \20874 ,
         \20875 , \20876 , \20877 , \20878 , \20879 , \20880 , \20881 , \20882 , \20883 , \20884 ,
         \20885 , \20886 , \20887 , \20888 , \20889 , \20890 , \20891 , \20892 , \20893 , \20894 ,
         \20895 , \20896 , \20897 , \20898 , \20899 , \20900 , \20901 , \20902 , \20903 , \20904 ,
         \20905 , \20906 , \20907 , \20908 , \20909 , \20910 , \20911 , \20912 , \20913 , \20914 ,
         \20915 , \20916 , \20917 , \20918 , \20919 , \20920 , \20921 , \20922 , \20923 , \20924 ,
         \20925 , \20926 , \20927 , \20928 , \20929 , \20930 , \20931 , \20932 , \20933 , \20934 ,
         \20935 , \20936 , \20937 , \20938 , \20939 , \20940 , \20941 , \20942 , \20943 , \20944 ,
         \20945 , \20946 , \20947 , \20948 , \20949 , \20950 , \20951 , \20952 , \20953 , \20954 ,
         \20955 , \20956 , \20957 , \20958 , \20959 , \20960 , \20961 , \20962 , \20963 , \20964 ,
         \20965 , \20966 , \20967 , \20968 , \20969 , \20970 , \20971 , \20972 , \20973 , \20974 ,
         \20975 , \20976 , \20977 , \20978 , \20979 , \20980 , \20981 , \20982 , \20983 , \20984 ,
         \20985 , \20986 , \20987 , \20988 , \20989 , \20990 , \20991 , \20992 , \20993 , \20994 ,
         \20995 , \20996 , \20997 , \20998 , \20999 , \21000 , \21001 , \21002 , \21003 , \21004 ,
         \21005 , \21006 , \21007 , \21008 , \21009 , \21010 , \21011 , \21012 , \21013 , \21014 ,
         \21015 , \21016 , \21017 , \21018 , \21019 , \21020 , \21021 , \21022 , \21023 , \21024 ,
         \21025 , \21026 , \21027 , \21028 , \21029 , \21030 , \21031 , \21032 , \21033 , \21034 ,
         \21035 , \21036 , \21037 , \21038 , \21039 , \21040 , \21041 , \21042 , \21043 , \21044 ,
         \21045 , \21046 , \21047 , \21048 , \21049 , \21050 , \21051 , \21052 , \21053 , \21054 ,
         \21055 , \21056 , \21057 , \21058 , \21059 , \21060 , \21061 , \21062 , \21063 , \21064 ,
         \21065 , \21066 , \21067 , \21068 , \21069 , \21070 , \21071 , \21072 , \21073 , \21074 ,
         \21075 , \21076 , \21077 , \21078 , \21079 , \21080 , \21081 , \21082 , \21083 , \21084 ,
         \21085 , \21086 , \21087 , \21088 , \21089 , \21090 , \21091 , \21092 , \21093 , \21094 ,
         \21095 , \21096 , \21097 , \21098 , \21099 , \21100 , \21101 , \21102 , \21103 , \21104 ,
         \21105 , \21106 , \21107 , \21108 , \21109 , \21110 , \21111 , \21112 , \21113 , \21114 ,
         \21115 , \21116 , \21117 , \21118 , \21119 , \21120 , \21121 , \21122 , \21123 , \21124 ,
         \21125 , \21126 , \21127 , \21128 , \21129 , \21130 , \21131 , \21132 , \21133 , \21134 ,
         \21135 , \21136 , \21137 , \21138 , \21139 , \21140 , \21141 , \21142 , \21143 , \21144 ,
         \21145 , \21146 , \21147 , \21148 , \21149 , \21150 , \21151 , \21152 , \21153 , \21154 ,
         \21155 , \21156 , \21157 , \21158 , \21159 , \21160 , \21161 , \21162 , \21163 , \21164 ,
         \21165 , \21166 , \21167 , \21168 , \21169 , \21170 , \21171 , \21172 , \21173 , \21174 ,
         \21175 , \21176 , \21177 , \21178 , \21179 , \21180 , \21181 , \21182 , \21183 , \21184 ,
         \21185 , \21186 , \21187 , \21188 , \21189 , \21190 , \21191 , \21192 , \21193 , \21194 ,
         \21195 , \21196 , \21197 , \21198 , \21199 , \21200 , \21201 , \21202 , \21203 , \21204 ,
         \21205 , \21206 , \21207 , \21208 , \21209 , \21210 , \21211 , \21212 , \21213 , \21214 ,
         \21215 , \21216 , \21217 , \21218 , \21219 , \21220 , \21221 , \21222 , \21223 , \21224 ,
         \21225 , \21226 , \21227 , \21228 , \21229 , \21230 , \21231 , \21232 , \21233 , \21234 ,
         \21235 , \21236 , \21237 , \21238 , \21239 , \21240 , \21241 , \21242 , \21243 , \21244 ,
         \21245 , \21246 , \21247 , \21248 , \21249 , \21250 , \21251 , \21252 , \21253 , \21254 ,
         \21255 , \21256 , \21257 , \21258 , \21259 , \21260 , \21261 , \21262 , \21263 , \21264 ,
         \21265 , \21266 , \21267 , \21268 , \21269 , \21270 , \21271 , \21272 , \21273 , \21274 ,
         \21275 , \21276 , \21277 , \21278 , \21279 , \21280 , \21281 , \21282 , \21283 , \21284 ,
         \21285 , \21286 , \21287 , \21288 , \21289 , \21290 , \21291 , \21292 , \21293 , \21294 ,
         \21295 , \21296 , \21297 , \21298 , \21299 , \21300 , \21301 , \21302 , \21303 , \21304 ,
         \21305 , \21306 , \21307 , \21308 , \21309 , \21310 , \21311 , \21312 , \21313 , \21314 ,
         \21315 , \21316 , \21317 , \21318 , \21319 , \21320 , \21321 , \21322 , \21323 , \21324 ,
         \21325 , \21326 , \21327 , \21328 , \21329 , \21330 , \21331 , \21332 , \21333 , \21334 ,
         \21335 , \21336 , \21337 , \21338 , \21339 , \21340 , \21341 , \21342 , \21343 , \21344 ,
         \21345 , \21346 , \21347 , \21348 , \21349 , \21350 , \21351 , \21352 , \21353 , \21354 ,
         \21355 , \21356 , \21357 , \21358 , \21359 , \21360 , \21361 , \21362 , \21363 , \21364 ,
         \21365 , \21366 , \21367 , \21368 , \21369 , \21370 , \21371 , \21372 , \21373 , \21374 ,
         \21375 , \21376 , \21377 , \21378 , \21379 , \21380 , \21381 , \21382 , \21383 , \21384 ,
         \21385 , \21386 , \21387 , \21388 , \21389 , \21390 , \21391 , \21392 , \21393 , \21394 ,
         \21395 , \21396 , \21397 , \21398 , \21399 , \21400 , \21401 , \21402 , \21403 , \21404 ,
         \21405 , \21406 , \21407 , \21408 , \21409 , \21410 , \21411 , \21412 , \21413 , \21414 ,
         \21415 , \21416 , \21417 , \21418 , \21419 , \21420 , \21421 , \21422 , \21423 , \21424 ,
         \21425 , \21426 , \21427 , \21428 , \21429 , \21430 , \21431 , \21432 , \21433 , \21434 ,
         \21435 , \21436 , \21437 , \21438 , \21439 , \21440 , \21441 , \21442 , \21443 , \21444 ,
         \21445 , \21446 , \21447 , \21448 , \21449 , \21450 , \21451 , \21452 , \21453 , \21454 ,
         \21455 , \21456 , \21457 , \21458 , \21459 , \21460 , \21461 , \21462 , \21463 , \21464 ,
         \21465 , \21466 , \21467 , \21468 , \21469 , \21470 , \21471 , \21472 , \21473 , \21474 ,
         \21475 , \21476 , \21477 , \21478 , \21479 , \21480 , \21481 , \21482 , \21483 , \21484 ,
         \21485 , \21486 , \21487 , \21488 , \21489 , \21490 , \21491 , \21492 , \21493 , \21494 ,
         \21495 , \21496 , \21497 , \21498 , \21499 , \21500 , \21501 , \21502 , \21503 , \21504 ,
         \21505 , \21506 , \21507 , \21508 , \21509 , \21510 , \21511 , \21512 , \21513 , \21514 ,
         \21515 , \21516 , \21517 , \21518 , \21519 , \21520 , \21521 , \21522 , \21523 , \21524 ,
         \21525 , \21526 , \21527 , \21528 , \21529 , \21530 , \21531 , \21532 , \21533 , \21534 ,
         \21535 , \21536 , \21537 , \21538 , \21539 , \21540 , \21541 , \21542 , \21543 , \21544 ,
         \21545 , \21546 , \21547 , \21548 , \21549 , \21550 , \21551 , \21552 , \21553 , \21554 ,
         \21555 , \21556 , \21557 , \21558 , \21559 , \21560 , \21561 , \21562 , \21563 , \21564 ,
         \21565 , \21566 , \21567 , \21568 , \21569 , \21570 , \21571 , \21572 , \21573 , \21574 ,
         \21575 , \21576 , \21577 , \21578 , \21579 , \21580 , \21581 , \21582 , \21583 , \21584 ,
         \21585 , \21586 , \21587 , \21588 , \21589 , \21590 , \21591 , \21592 , \21593 , \21594 ,
         \21595 , \21596 , \21597 , \21598 , \21599 , \21600 , \21601 , \21602 , \21603 , \21604 ,
         \21605 , \21606 , \21607 , \21608 , \21609 , \21610 , \21611 , \21612 , \21613 , \21614 ,
         \21615 , \21616 , \21617 , \21618 , \21619 , \21620 , \21621 , \21622 , \21623 , \21624 ,
         \21625 , \21626 , \21627 , \21628 , \21629 , \21630 , \21631 , \21632 , \21633 , \21634 ,
         \21635 , \21636 , \21637 , \21638 , \21639 , \21640 , \21641 , \21642 , \21643 , \21644 ,
         \21645 , \21646 , \21647 , \21648 , \21649 , \21650 , \21651 , \21652 , \21653 , \21654 ,
         \21655 , \21656 , \21657 , \21658 , \21659 , \21660 , \21661 , \21662 , \21663 , \21664 ,
         \21665 , \21666 , \21667 , \21668 , \21669 , \21670 , \21671 , \21672 , \21673 , \21674 ,
         \21675 , \21676 , \21677 , \21678 , \21679 , \21680 , \21681 , \21682 , \21683 , \21684 ,
         \21685 , \21686 , \21687 , \21688 , \21689 , \21690 , \21691 , \21692 , \21693 , \21694 ,
         \21695 , \21696 , \21697 , \21698 , \21699 , \21700 , \21701 , \21702 , \21703 , \21704 ,
         \21705 , \21706 , \21707 , \21708 , \21709 , \21710 , \21711 , \21712 , \21713 , \21714 ,
         \21715 , \21716 , \21717 , \21718 , \21719 , \21720 , \21721 , \21722 , \21723 , \21724 ,
         \21725 , \21726 , \21727 , \21728 , \21729 , \21730 , \21731 , \21732 , \21733 , \21734 ,
         \21735 , \21736 , \21737 , \21738 , \21739 , \21740 , \21741 , \21742 , \21743 , \21744 ,
         \21745 , \21746 , \21747 , \21748 , \21749 , \21750 , \21751 , \21752 , \21753 , \21754 ,
         \21755 , \21756 , \21757 , \21758 , \21759 , \21760 , \21761 , \21762 , \21763 , \21764 ,
         \21765 , \21766 , \21767 , \21768 , \21769 , \21770 , \21771 , \21772 , \21773 , \21774 ,
         \21775 , \21776 , \21777 , \21778 , \21779 , \21780 , \21781 , \21782 , \21783 , \21784 ,
         \21785 , \21786 , \21787 , \21788 , \21789 , \21790 , \21791 , \21792 , \21793 , \21794 ,
         \21795 , \21796 , \21797 , \21798 , \21799 , \21800 , \21801 , \21802 , \21803 , \21804 ,
         \21805 , \21806 , \21807 , \21808 , \21809 , \21810 , \21811 , \21812 , \21813 , \21814 ,
         \21815 , \21816 , \21817 , \21818 , \21819 , \21820 , \21821 , \21822 , \21823 , \21824 ,
         \21825 , \21826 , \21827 , \21828 , \21829 , \21830 , \21831 , \21832 , \21833 , \21834 ,
         \21835 , \21836 , \21837 , \21838 , \21839 , \21840 , \21841 , \21842 , \21843 , \21844 ,
         \21845 , \21846 , \21847 , \21848 , \21849 , \21850 , \21851 , \21852 , \21853 , \21854 ,
         \21855 , \21856 , \21857 , \21858 , \21859 , \21860 , \21861 , \21862 , \21863 , \21864 ,
         \21865 , \21866 , \21867 , \21868 , \21869 , \21870 , \21871 , \21872 , \21873 , \21874 ,
         \21875 , \21876 , \21877 , \21878 , \21879 , \21880 , \21881 , \21882 , \21883 , \21884 ,
         \21885 , \21886 , \21887 , \21888 , \21889 , \21890 , \21891 , \21892 , \21893 , \21894 ,
         \21895 , \21896 , \21897 , \21898 , \21899 , \21900 , \21901 , \21902 , \21903 , \21904 ,
         \21905 , \21906 , \21907 , \21908 , \21909 , \21910 , \21911 , \21912 , \21913 , \21914 ,
         \21915 , \21916 , \21917 , \21918 , \21919 , \21920 , \21921 , \21922 , \21923 , \21924 ,
         \21925 , \21926 , \21927 , \21928 , \21929 , \21930 , \21931 , \21932 , \21933 , \21934 ,
         \21935 , \21936 , \21937 , \21938 , \21939 , \21940 , \21941 , \21942 , \21943 , \21944 ,
         \21945 , \21946 , \21947 , \21948 , \21949 , \21950 , \21951 , \21952 , \21953 , \21954 ,
         \21955 , \21956 , \21957 , \21958 , \21959 , \21960 , \21961 , \21962 , \21963 , \21964 ,
         \21965 , \21966 , \21967 , \21968 , \21969 , \21970 , \21971 , \21972 , \21973 , \21974 ,
         \21975 , \21976 , \21977 , \21978 , \21979 , \21980 , \21981 , \21982 , \21983 , \21984 ,
         \21985 , \21986 , \21987 , \21988 , \21989 , \21990 , \21991 , \21992 , \21993 , \21994 ,
         \21995 , \21996 , \21997 , \21998 , \21999 , \22000 , \22001 , \22002 , \22003 , \22004 ,
         \22005 , \22006 , \22007 , \22008 , \22009 , \22010 , \22011 , \22012 , \22013 , \22014 ,
         \22015 , \22016 , \22017 , \22018 , \22019 , \22020 , \22021 , \22022 , \22023 , \22024 ,
         \22025 , \22026 , \22027 , \22028 , \22029 , \22030 , \22031 , \22032 , \22033 , \22034 ,
         \22035 , \22036 , \22037 , \22038 , \22039 , \22040 , \22041 , \22042 , \22043 , \22044 ,
         \22045 , \22046 , \22047 , \22048 , \22049 , \22050 , \22051 , \22052 , \22053 , \22054 ,
         \22055 , \22056 , \22057 , \22058 , \22059 , \22060 , \22061 , \22062 , \22063 , \22064 ,
         \22065 , \22066 , \22067 , \22068 , \22069 , \22070 , \22071 , \22072 , \22073 , \22074 ,
         \22075 , \22076 , \22077 , \22078 , \22079 , \22080 , \22081 , \22082 , \22083 , \22084 ,
         \22085 , \22086 , \22087 , \22088 , \22089 , \22090 , \22091 , \22092 , \22093 , \22094 ,
         \22095 , \22096 , \22097 , \22098 , \22099 , \22100 , \22101 , \22102 , \22103 , \22104 ,
         \22105 , \22106 , \22107 , \22108 , \22109 , \22110 , \22111 , \22112 , \22113 , \22114 ,
         \22115 , \22116 , \22117 , \22118 , \22119 , \22120 , \22121 , \22122 , \22123 , \22124 ,
         \22125 , \22126 , \22127 , \22128 , \22129 , \22130 , \22131 , \22132 , \22133 , \22134 ,
         \22135 , \22136 , \22137 , \22138 , \22139 , \22140 , \22141 , \22142 , \22143 , \22144 ,
         \22145 , \22146 , \22147 , \22148 , \22149 , \22150 , \22151 , \22152 , \22153 , \22154 ,
         \22155 , \22156 , \22157 , \22158 , \22159 , \22160 , \22161 , \22162 , \22163 , \22164 ,
         \22165 , \22166 , \22167 , \22168 , \22169 , \22170 , \22171 , \22172 , \22173 , \22174 ,
         \22175 , \22176 , \22177 , \22178 , \22179 , \22180 , \22181 , \22182 , \22183 , \22184 ,
         \22185 , \22186 , \22187 , \22188 , \22189 , \22190 , \22191 , \22192 , \22193 , \22194 ,
         \22195 , \22196 , \22197 , \22198 , \22199 , \22200 , \22201 , \22202 , \22203 , \22204 ,
         \22205 , \22206 , \22207 , \22208 , \22209 , \22210 , \22211 , \22212 , \22213 , \22214 ,
         \22215 , \22216 , \22217 , \22218 , \22219 , \22220 , \22221 , \22222 , \22223 , \22224 ,
         \22225 , \22226 , \22227 , \22228 , \22229 , \22230 , \22231 , \22232 , \22233 , \22234 ,
         \22235 , \22236 , \22237 , \22238 , \22239 , \22240 , \22241 , \22242 , \22243 , \22244 ,
         \22245 , \22246 , \22247 , \22248 , \22249 , \22250 , \22251 , \22252 , \22253 , \22254 ,
         \22255 , \22256 , \22257 , \22258 , \22259 , \22260 , \22261 , \22262 , \22263 , \22264 ,
         \22265 , \22266 , \22267 , \22268 , \22269 , \22270 , \22271 , \22272 , \22273 , \22274 ,
         \22275 , \22276 , \22277 , \22278 , \22279 , \22280 , \22281 , \22282 , \22283 , \22284 ,
         \22285 , \22286 , \22287 , \22288 , \22289 , \22290 , \22291 , \22292 , \22293 , \22294 ,
         \22295 , \22296 , \22297 , \22298 , \22299 , \22300 , \22301 , \22302 , \22303 , \22304 ,
         \22305 , \22306 , \22307 , \22308 , \22309 , \22310 , \22311 , \22312 , \22313 , \22314 ,
         \22315 , \22316 , \22317 , \22318 , \22319 , \22320 , \22321 , \22322 , \22323 , \22324 ,
         \22325 , \22326 , \22327 , \22328 , \22329 , \22330 , \22331 , \22332 , \22333 , \22334 ,
         \22335 , \22336 , \22337 , \22338 , \22339 , \22340 , \22341 , \22342 , \22343 , \22344 ,
         \22345 , \22346 , \22347 , \22348 , \22349 , \22350 , \22351 , \22352 , \22353 , \22354 ,
         \22355 , \22356 , \22357 , \22358 , \22359 , \22360 , \22361 , \22362 , \22363 , \22364 ,
         \22365 , \22366 , \22367 , \22368 , \22369 , \22370 , \22371 , \22372 , \22373 , \22374 ,
         \22375 , \22376 , \22377 , \22378 , \22379 , \22380 , \22381 , \22382 , \22383 , \22384 ,
         \22385 , \22386 , \22387 , \22388 , \22389 , \22390 , \22391 , \22392 , \22393 , \22394 ,
         \22395 , \22396 , \22397 , \22398 , \22399 , \22400 , \22401 , \22402 , \22403 , \22404 ,
         \22405 , \22406 , \22407 , \22408 , \22409 , \22410 , \22411 , \22412 , \22413 , \22414 ,
         \22415 , \22416 , \22417 , \22418 , \22419 , \22420 , \22421 , \22422 , \22423 , \22424 ,
         \22425 , \22426 , \22427 , \22428 , \22429 , \22430 , \22431 , \22432 , \22433 , \22434 ,
         \22435 , \22436 , \22437 , \22438 , \22439 , \22440 , \22441 , \22442 , \22443 , \22444 ,
         \22445 , \22446 , \22447 , \22448 , \22449 , \22450 , \22451 , \22452 , \22453 , \22454 ,
         \22455 , \22456 , \22457 , \22458 , \22459 , \22460 , \22461 , \22462 , \22463 , \22464 ,
         \22465 , \22466 , \22467 , \22468 , \22469 , \22470 , \22471 , \22472 , \22473 , \22474 ,
         \22475 , \22476 , \22477 , \22478 , \22479 , \22480 , \22481 , \22482 , \22483 , \22484 ,
         \22485 , \22486 , \22487 , \22488 , \22489 , \22490 , \22491 , \22492 , \22493 , \22494 ,
         \22495 , \22496 , \22497 , \22498 , \22499 , \22500 , \22501 , \22502 , \22503 , \22504 ,
         \22505 , \22506 , \22507 , \22508 , \22509 , \22510 , \22511 , \22512 , \22513 , \22514 ,
         \22515 , \22516 , \22517 , \22518 , \22519 , \22520 , \22521 , \22522 , \22523 , \22524 ,
         \22525 , \22526 , \22527 , \22528 , \22529 , \22530 , \22531 , \22532 , \22533 , \22534 ,
         \22535 , \22536 , \22537 , \22538 , \22539 , \22540 , \22541 , \22542 , \22543 , \22544 ,
         \22545 , \22546 , \22547 , \22548 , \22549 , \22550 , \22551 , \22552 , \22553 , \22554 ,
         \22555 , \22556 , \22557 , \22558 , \22559 , \22560 , \22561 , \22562 , \22563 , \22564 ,
         \22565 , \22566 , \22567 , \22568 , \22569 , \22570 , \22571 , \22572 , \22573 , \22574 ,
         \22575 , \22576 , \22577 , \22578 , \22579 , \22580 , \22581 , \22582 , \22583 , \22584 ,
         \22585 , \22586 , \22587 , \22588 , \22589 , \22590 , \22591 , \22592 , \22593 , \22594 ,
         \22595 , \22596 , \22597 , \22598 , \22599 , \22600 , \22601 , \22602 , \22603 , \22604 ,
         \22605 , \22606 , \22607 , \22608 , \22609 , \22610 , \22611 , \22612 , \22613 , \22614 ,
         \22615 , \22616 , \22617 , \22618 , \22619 , \22620 , \22621 , \22622 , \22623 , \22624 ,
         \22625 , \22626 , \22627 , \22628 , \22629 , \22630 , \22631 , \22632 , \22633 , \22634 ,
         \22635 , \22636 , \22637 , \22638 , \22639 , \22640 , \22641 , \22642 , \22643 , \22644 ,
         \22645 , \22646 , \22647 , \22648 , \22649 , \22650 , \22651 , \22652 , \22653 , \22654 ,
         \22655 , \22656 , \22657 , \22658 , \22659 , \22660 , \22661 , \22662 , \22663 , \22664 ,
         \22665 , \22666 , \22667 , \22668 , \22669 , \22670 , \22671 , \22672 , \22673 , \22674 ,
         \22675 , \22676 , \22677 , \22678 , \22679 , \22680 , \22681 , \22682 , \22683 , \22684 ,
         \22685 , \22686 , \22687 , \22688 , \22689 , \22690 , \22691 , \22692 , \22693 , \22694 ,
         \22695 , \22696 , \22697 , \22698 , \22699 , \22700 , \22701 , \22702 , \22703 , \22704 ,
         \22705 , \22706 , \22707 , \22708 , \22709 , \22710 , \22711 , \22712 , \22713 , \22714 ,
         \22715 , \22716 , \22717 , \22718 , \22719 , \22720 , \22721 , \22722 , \22723 , \22724 ,
         \22725 , \22726 , \22727 , \22728 , \22729 , \22730 , \22731 , \22732 , \22733 , \22734 ,
         \22735 , \22736 , \22737 , \22738 , \22739 , \22740 , \22741 , \22742 , \22743 , \22744 ,
         \22745 , \22746 , \22747 , \22748 , \22749 , \22750 , \22751 , \22752 , \22753 , \22754 ,
         \22755 , \22756 , \22757 , \22758 , \22759 , \22760 , \22761 , \22762 , \22763 , \22764 ,
         \22765 , \22766 , \22767 , \22768 , \22769 , \22770 , \22771 , \22772 , \22773 , \22774 ,
         \22775 , \22776 , \22777 , \22778 , \22779 , \22780 , \22781 , \22782 , \22783 , \22784 ,
         \22785 , \22786 , \22787 , \22788 , \22789 , \22790 , \22791 , \22792 , \22793 , \22794 ,
         \22795 , \22796 , \22797 , \22798 , \22799 , \22800 , \22801 , \22802 , \22803 , \22804 ,
         \22805 , \22806 , \22807 , \22808 , \22809 , \22810 , \22811 , \22812 , \22813 , \22814 ,
         \22815 , \22816 , \22817 , \22818 , \22819 , \22820 , \22821 , \22822 , \22823 , \22824 ,
         \22825 , \22826 , \22827 , \22828 , \22829 , \22830 , \22831 , \22832 , \22833 , \22834 ,
         \22835 , \22836 , \22837 , \22838 , \22839 , \22840 , \22841 , \22842 , \22843 , \22844 ,
         \22845 , \22846 , \22847 , \22848 , \22849 , \22850 , \22851 , \22852 , \22853 , \22854 ,
         \22855 , \22856 , \22857 , \22858 , \22859 , \22860 , \22861 , \22862 , \22863 , \22864 ,
         \22865 , \22866 , \22867 , \22868 , \22869 , \22870 , \22871 , \22872 , \22873 , \22874 ,
         \22875 , \22876 , \22877 , \22878 , \22879 , \22880 , \22881 , \22882 , \22883 , \22884 ,
         \22885 , \22886 , \22887 , \22888 , \22889 , \22890 , \22891 , \22892 , \22893 , \22894 ,
         \22895 , \22896 , \22897 , \22898 , \22899 , \22900 , \22901 , \22902 , \22903 , \22904 ,
         \22905 , \22906 , \22907 , \22908 , \22909 , \22910 , \22911 , \22912 , \22913 , \22914 ,
         \22915 , \22916 , \22917 , \22918 , \22919 , \22920 , \22921 , \22922 , \22923 , \22924 ,
         \22925 , \22926 , \22927 , \22928 , \22929 , \22930 , \22931 , \22932 , \22933 , \22934 ,
         \22935 , \22936 , \22937 , \22938 , \22939 , \22940 , \22941 , \22942 , \22943 , \22944 ,
         \22945 , \22946 , \22947 , \22948 , \22949 , \22950 , \22951 , \22952 , \22953 , \22954 ,
         \22955 , \22956 , \22957 , \22958 , \22959 , \22960 , \22961 , \22962 , \22963 , \22964 ,
         \22965 , \22966 , \22967 , \22968 , \22969 , \22970 , \22971 , \22972 , \22973 , \22974 ,
         \22975 , \22976 , \22977 , \22978 , \22979 , \22980 , \22981 , \22982 , \22983 , \22984 ,
         \22985 , \22986 , \22987 , \22988 , \22989 , \22990 , \22991 , \22992 , \22993 , \22994 ,
         \22995 , \22996 , \22997 , \22998 , \22999 , \23000 , \23001 , \23002 , \23003 , \23004 ,
         \23005 , \23006 , \23007 , \23008 , \23009 , \23010 , \23011 , \23012 , \23013 , \23014 ,
         \23015 , \23016 , \23017 , \23018 , \23019 , \23020 , \23021 , \23022 , \23023 , \23024 ,
         \23025 , \23026 , \23027 , \23028 , \23029 , \23030 , \23031 , \23032 , \23033 , \23034 ,
         \23035 , \23036 , \23037 , \23038 , \23039 , \23040 , \23041 , \23042 , \23043 , \23044 ,
         \23045 , \23046 , \23047 , \23048 , \23049 , \23050 , \23051 , \23052 , \23053 , \23054 ,
         \23055 , \23056 , \23057 , \23058 , \23059 , \23060 , \23061 , \23062 , \23063 , \23064 ,
         \23065 , \23066 , \23067 , \23068 , \23069 , \23070 , \23071 , \23072 , \23073 , \23074 ,
         \23075 , \23076 , \23077 , \23078 , \23079 , \23080 , \23081 , \23082 , \23083 , \23084 ,
         \23085 , \23086 , \23087 , \23088 , \23089 , \23090 , \23091 , \23092 , \23093 , \23094 ,
         \23095 , \23096 , \23097 , \23098 , \23099 , \23100 , \23101 , \23102 , \23103 , \23104 ,
         \23105 , \23106 , \23107 , \23108 , \23109 , \23110 , \23111 , \23112 , \23113 , \23114 ,
         \23115 , \23116 , \23117 , \23118 , \23119 , \23120 , \23121 , \23122 , \23123 , \23124 ,
         \23125 , \23126 , \23127 , \23128 , \23129 , \23130 , \23131 , \23132 , \23133 , \23134 ,
         \23135 , \23136 , \23137 , \23138 , \23139 , \23140 , \23141 , \23142 , \23143 , \23144 ,
         \23145 , \23146 , \23147 , \23148 , \23149 , \23150 , \23151 , \23152 , \23153 , \23154 ,
         \23155 , \23156 , \23157 , \23158 , \23159 , \23160 , \23161 , \23162 , \23163 , \23164 ,
         \23165 , \23166 , \23167 , \23168 , \23169 , \23170 , \23171 , \23172 , \23173 , \23174 ,
         \23175 , \23176 , \23177 , \23178 , \23179 , \23180 , \23181 , \23182 , \23183 , \23184 ,
         \23185 , \23186 , \23187 , \23188 , \23189 , \23190 , \23191 , \23192 , \23193 , \23194 ,
         \23195 , \23196 , \23197 , \23198 , \23199 , \23200 , \23201 , \23202 , \23203 , \23204 ,
         \23205 , \23206 , \23207 , \23208 , \23209 , \23210 , \23211 , \23212 , \23213 , \23214 ,
         \23215 , \23216 , \23217 , \23218 , \23219 , \23220 , \23221 , \23222 , \23223 , \23224 ,
         \23225 , \23226 , \23227 , \23228 , \23229 , \23230 , \23231 , \23232 , \23233 , \23234 ,
         \23235 , \23236 , \23237 , \23238 , \23239 , \23240 , \23241 , \23242 , \23243 , \23244 ,
         \23245 , \23246 , \23247 , \23248 , \23249 , \23250 , \23251 , \23252 , \23253 , \23254 ,
         \23255 , \23256 , \23257 , \23258 , \23259 , \23260 , \23261 , \23262 , \23263 , \23264 ,
         \23265 , \23266 , \23267 , \23268 , \23269 , \23270 , \23271 , \23272 , \23273 , \23274 ,
         \23275 , \23276 , \23277 , \23278 , \23279 , \23280 , \23281 , \23282 , \23283 , \23284 ,
         \23285 , \23286 , \23287 , \23288 , \23289 , \23290 , \23291 , \23292 , \23293 , \23294 ,
         \23295 , \23296 , \23297 , \23298 , \23299 , \23300 , \23301 , \23302 , \23303 , \23304 ,
         \23305 , \23306 , \23307 , \23308 , \23309 , \23310 , \23311 , \23312 , \23313 , \23314 ,
         \23315 , \23316 , \23317 , \23318 , \23319 , \23320 , \23321 , \23322 , \23323 , \23324 ,
         \23325 , \23326 , \23327 , \23328 , \23329 , \23330 , \23331 , \23332 , \23333 , \23334 ,
         \23335 , \23336 , \23337 , \23338 , \23339 , \23340 , \23341 , \23342 , \23343 , \23344 ,
         \23345 , \23346 , \23347 , \23348 , \23349 , \23350 , \23351 , \23352 , \23353 , \23354 ,
         \23355 , \23356 , \23357 , \23358 , \23359 , \23360 , \23361 , \23362 , \23363 , \23364 ,
         \23365 , \23366 , \23367 , \23368 , \23369 , \23370 , \23371 , \23372 , \23373 , \23374 ,
         \23375 , \23376 , \23377 , \23378 , \23379 , \23380 , \23381 , \23382 , \23383 , \23384 ,
         \23385 , \23386 , \23387 , \23388 , \23389 , \23390 , \23391 , \23392 , \23393 , \23394 ,
         \23395 , \23396 , \23397 , \23398 , \23399 , \23400 , \23401 , \23402 , \23403 , \23404 ,
         \23405 , \23406 , \23407 , \23408 , \23409 , \23410 , \23411 , \23412 , \23413 , \23414 ,
         \23415 , \23416 , \23417 , \23418 , \23419 , \23420 , \23421 , \23422 , \23423 , \23424 ,
         \23425 , \23426 , \23427 , \23428 , \23429 , \23430 , \23431 , \23432 , \23433 , \23434 ,
         \23435 , \23436 , \23437 , \23438 , \23439 , \23440 , \23441 , \23442 , \23443 , \23444 ,
         \23445 , \23446 , \23447 , \23448 , \23449 , \23450 , \23451 , \23452 , \23453 , \23454 ,
         \23455 , \23456 , \23457 , \23458 , \23459 , \23460 , \23461 , \23462 , \23463 , \23464 ,
         \23465 , \23466 , \23467 , \23468 , \23469 , \23470 , \23471 , \23472 , \23473 , \23474 ,
         \23475 , \23476 , \23477 , \23478 , \23479 , \23480 , \23481 , \23482 , \23483 , \23484 ,
         \23485 , \23486 , \23487 , \23488 , \23489 , \23490 , \23491 , \23492 , \23493 , \23494 ,
         \23495 , \23496 , \23497 , \23498 , \23499 , \23500 , \23501 , \23502 , \23503 , \23504 ,
         \23505 , \23506 , \23507 , \23508 , \23509 , \23510 , \23511 , \23512 , \23513 , \23514 ,
         \23515 , \23516 , \23517 , \23518 , \23519 , \23520 , \23521 , \23522 , \23523 , \23524 ,
         \23525 , \23526 , \23527 , \23528 , \23529 , \23530 , \23531 , \23532 , \23533 , \23534 ,
         \23535 , \23536 , \23537 , \23538 , \23539 , \23540 , \23541 , \23542 , \23543 , \23544 ,
         \23545 , \23546 , \23547 , \23548 , \23549 , \23550 , \23551 , \23552 , \23553 , \23554 ,
         \23555 , \23556 , \23557 , \23558 , \23559 , \23560 , \23561 , \23562 , \23563 , \23564 ,
         \23565 , \23566 , \23567 , \23568 , \23569 , \23570 , \23571 , \23572 , \23573 , \23574 ,
         \23575 , \23576 , \23577 , \23578 , \23579 , \23580 , \23581 , \23582 , \23583 , \23584 ,
         \23585 , \23586 , \23587 , \23588 , \23589 , \23590 , \23591 , \23592 , \23593 , \23594 ,
         \23595 , \23596 , \23597 , \23598 , \23599 , \23600 , \23601 , \23602 , \23603 , \23604 ,
         \23605 , \23606 , \23607 , \23608 , \23609 , \23610 , \23611 , \23612 , \23613 , \23614 ,
         \23615 , \23616 , \23617 , \23618 , \23619 , \23620 , \23621 , \23622 , \23623 , \23624 ,
         \23625 , \23626 , \23627 , \23628 , \23629 , \23630 , \23631 , \23632 , \23633 , \23634 ,
         \23635 , \23636 , \23637 , \23638 , \23639 , \23640 , \23641 , \23642 , \23643 , \23644 ,
         \23645 , \23646 , \23647 , \23648 , \23649 , \23650 , \23651 , \23652 , \23653 , \23654 ,
         \23655 , \23656 , \23657 , \23658 , \23659 , \23660 , \23661 , \23662 , \23663 , \23664 ,
         \23665 , \23666 , \23667 , \23668 , \23669 , \23670 , \23671 , \23672 , \23673 , \23674 ,
         \23675 , \23676 , \23677 , \23678 , \23679 , \23680 , \23681 , \23682 , \23683 , \23684 ,
         \23685 , \23686 , \23687 , \23688 , \23689 , \23690 , \23691 , \23692 , \23693 , \23694 ,
         \23695 , \23696 , \23697 , \23698 , \23699 , \23700 , \23701 , \23702 , \23703 , \23704 ,
         \23705 , \23706 , \23707 , \23708 , \23709 , \23710 , \23711 , \23712 , \23713 , \23714 ,
         \23715 , \23716 , \23717 , \23718 , \23719 , \23720 , \23721 , \23722 , \23723 , \23724 ,
         \23725 , \23726 , \23727 , \23728 , \23729 , \23730 , \23731 , \23732 , \23733 , \23734 ,
         \23735 , \23736 , \23737 , \23738 , \23739 , \23740 , \23741 , \23742 , \23743 , \23744 ,
         \23745 , \23746 , \23747 , \23748 , \23749 , \23750 , \23751 , \23752 , \23753 , \23754 ,
         \23755 , \23756 , \23757 , \23758 , \23759 , \23760 , \23761 , \23762 , \23763 , \23764 ,
         \23765 , \23766 , \23767 , \23768 , \23769 , \23770 , \23771 , \23772 , \23773 , \23774 ,
         \23775 , \23776 , \23777 , \23778 , \23779 , \23780 , \23781 , \23782 , \23783 , \23784 ,
         \23785 , \23786 , \23787 , \23788 , \23789 , \23790 , \23791 , \23792 , \23793 , \23794 ,
         \23795 , \23796 , \23797 , \23798 , \23799 , \23800 , \23801 , \23802 , \23803 , \23804 ,
         \23805 , \23806 , \23807 , \23808 , \23809 , \23810 , \23811 , \23812 , \23813 , \23814 ,
         \23815 , \23816 , \23817 , \23818 , \23819 , \23820 , \23821 , \23822 , \23823 , \23824 ,
         \23825 , \23826 , \23827 , \23828 , \23829 , \23830 , \23831 , \23832 , \23833 , \23834 ,
         \23835 , \23836 , \23837 , \23838 , \23839 , \23840 , \23841 , \23842 , \23843 , \23844 ,
         \23845 , \23846 , \23847 , \23848 , \23849 , \23850 , \23851 , \23852 , \23853 , \23854 ,
         \23855 , \23856 , \23857 , \23858 , \23859 , \23860 , \23861 , \23862 , \23863 , \23864 ,
         \23865 , \23866 , \23867 , \23868 , \23869 , \23870 , \23871 , \23872 , \23873 , \23874 ,
         \23875 , \23876 , \23877 , \23878 , \23879 , \23880 , \23881 , \23882 , \23883 , \23884 ,
         \23885 , \23886 , \23887 , \23888 , \23889 , \23890 , \23891 , \23892 , \23893 , \23894 ,
         \23895 , \23896 , \23897 , \23898 , \23899 , \23900 , \23901 , \23902 , \23903 , \23904 ,
         \23905 , \23906 , \23907 , \23908 , \23909 , \23910 , \23911 , \23912 , \23913 , \23914 ,
         \23915 , \23916 , \23917 , \23918 , \23919 , \23920 , \23921 , \23922 , \23923 , \23924 ,
         \23925 , \23926 , \23927 , \23928 , \23929 , \23930 , \23931 , \23932 , \23933 , \23934 ,
         \23935 , \23936 , \23937 , \23938 , \23939 , \23940 , \23941 , \23942 , \23943 , \23944 ,
         \23945 , \23946 , \23947 , \23948 , \23949 , \23950 , \23951 , \23952 , \23953 , \23954 ,
         \23955 , \23956 , \23957 , \23958 , \23959 , \23960 , \23961 , \23962 , \23963 , \23964 ,
         \23965 , \23966 , \23967 , \23968 , \23969 , \23970 , \23971 , \23972 , \23973 , \23974 ,
         \23975 , \23976 , \23977 , \23978 , \23979 , \23980 , \23981 , \23982 , \23983 , \23984 ,
         \23985 , \23986 , \23987 , \23988 , \23989 , \23990 , \23991 , \23992 , \23993 , \23994 ,
         \23995 , \23996 , \23997 , \23998 , \23999 , \24000 , \24001 , \24002 , \24003 , \24004 ,
         \24005 , \24006 , \24007 , \24008 , \24009 , \24010 , \24011 , \24012 , \24013 , \24014 ,
         \24015 , \24016 , \24017 , \24018 , \24019 , \24020 , \24021 , \24022 , \24023 , \24024 ,
         \24025 , \24026 , \24027 , \24028 , \24029 , \24030 , \24031 , \24032 , \24033 , \24034 ,
         \24035 , \24036 , \24037 , \24038 , \24039 , \24040 , \24041 , \24042 , \24043 , \24044 ,
         \24045 , \24046 , \24047 , \24048 , \24049 , \24050 , \24051 , \24052 , \24053 , \24054 ,
         \24055 , \24056 , \24057 , \24058 , \24059 , \24060 , \24061 , \24062 , \24063 , \24064 ,
         \24065 , \24066 , \24067 , \24068 , \24069 , \24070 , \24071 , \24072 , \24073 , \24074 ,
         \24075 , \24076 , \24077 , \24078 , \24079 , \24080 , \24081 , \24082 , \24083 , \24084 ,
         \24085 , \24086 , \24087 , \24088 , \24089 , \24090 , \24091 , \24092 , \24093 , \24094 ,
         \24095 , \24096 , \24097 , \24098 , \24099 , \24100 , \24101 , \24102 , \24103 , \24104 ,
         \24105 , \24106 , \24107 , \24108 , \24109 , \24110 , \24111 , \24112 , \24113 , \24114 ,
         \24115 , \24116 , \24117 , \24118 , \24119 , \24120 , \24121 , \24122 , \24123 , \24124 ,
         \24125 , \24126 , \24127 , \24128 , \24129 , \24130 , \24131 , \24132 , \24133 , \24134 ,
         \24135 , \24136 , \24137 , \24138 , \24139 , \24140 , \24141 , \24142 , \24143 , \24144 ,
         \24145 , \24146 , \24147 , \24148 , \24149 , \24150 , \24151 , \24152 , \24153 , \24154 ,
         \24155 , \24156 , \24157 , \24158 , \24159 , \24160 , \24161 , \24162 , \24163 , \24164 ,
         \24165 , \24166 , \24167 , \24168 , \24169 , \24170 , \24171 , \24172 , \24173 , \24174 ,
         \24175 , \24176 , \24177 , \24178 , \24179 , \24180 , \24181 , \24182 , \24183 , \24184 ,
         \24185 , \24186 , \24187 , \24188 , \24189 , \24190 , \24191 , \24192 , \24193 , \24194 ,
         \24195 , \24196 , \24197 , \24198 , \24199 , \24200 , \24201 , \24202 , \24203 , \24204 ,
         \24205 , \24206 , \24207 , \24208 , \24209 , \24210 , \24211 , \24212 , \24213 , \24214 ,
         \24215 , \24216 , \24217 , \24218 , \24219 , \24220 , \24221 , \24222 , \24223 , \24224 ,
         \24225 , \24226 , \24227 , \24228 , \24229 , \24230 , \24231 , \24232 , \24233 , \24234 ,
         \24235 , \24236 , \24237 , \24238 , \24239 , \24240 , \24241 , \24242 , \24243 , \24244 ,
         \24245 , \24246 , \24247 , \24248 , \24249 , \24250 , \24251 , \24252 , \24253 , \24254 ,
         \24255 , \24256 , \24257 , \24258 , \24259 , \24260 , \24261 , \24262 , \24263 , \24264 ,
         \24265 , \24266 , \24267 , \24268 , \24269 , \24270 , \24271 , \24272 , \24273 , \24274 ,
         \24275 , \24276 , \24277 , \24278 , \24279 , \24280 , \24281 , \24282 , \24283 , \24284 ,
         \24285 , \24286 , \24287 , \24288 , \24289 , \24290 , \24291 , \24292 , \24293 , \24294 ,
         \24295 , \24296 , \24297 , \24298 , \24299 , \24300 , \24301 , \24302 , \24303 , \24304 ,
         \24305 , \24306 , \24307 , \24308 , \24309 , \24310 , \24311 , \24312 , \24313 , \24314 ,
         \24315 , \24316 , \24317 , \24318 , \24319 , \24320 , \24321 , \24322 , \24323 , \24324 ,
         \24325 , \24326 , \24327 , \24328 , \24329 , \24330 , \24331 , \24332 , \24333 , \24334 ,
         \24335 , \24336 , \24337 , \24338 , \24339 , \24340 , \24341 , \24342 , \24343 , \24344 ,
         \24345 , \24346 , \24347 , \24348 , \24349 , \24350 , \24351 , \24352 , \24353 , \24354 ,
         \24355 , \24356 , \24357 , \24358 , \24359 , \24360 , \24361 , \24362 , \24363 , \24364 ,
         \24365 , \24366 , \24367 , \24368 , \24369 , \24370 , \24371 , \24372 , \24373 , \24374 ,
         \24375 , \24376 , \24377 , \24378 , \24379 , \24380 , \24381 , \24382 , \24383 , \24384 ,
         \24385 , \24386 , \24387 , \24388 , \24389 , \24390 , \24391 , \24392 , \24393 , \24394 ,
         \24395 , \24396 , \24397 , \24398 , \24399 , \24400 , \24401 , \24402 , \24403 , \24404 ,
         \24405 , \24406 , \24407 , \24408 , \24409 , \24410 , \24411 , \24412 , \24413 , \24414 ,
         \24415 , \24416 , \24417 , \24418 , \24419 , \24420 , \24421 , \24422 , \24423 , \24424 ,
         \24425 , \24426 , \24427 , \24428 , \24429 , \24430 , \24431 , \24432 , \24433 , \24434 ,
         \24435 , \24436 , \24437 , \24438 , \24439 , \24440 , \24441 , \24442 , \24443 , \24444 ,
         \24445 , \24446 , \24447 , \24448 , \24449 , \24450 , \24451 , \24452 , \24453 , \24454 ,
         \24455 , \24456 , \24457 , \24458 , \24459 , \24460 , \24461 , \24462 , \24463 , \24464 ,
         \24465 , \24466 , \24467 , \24468 , \24469 , \24470 , \24471 , \24472 , \24473 , \24474 ,
         \24475 , \24476 , \24477 , \24478 , \24479 , \24480 , \24481 , \24482 , \24483 , \24484 ,
         \24485 , \24486 , \24487 , \24488 , \24489 , \24490 , \24491 , \24492 , \24493 , \24494 ,
         \24495 , \24496 , \24497 , \24498 , \24499 , \24500 , \24501 , \24502 , \24503 , \24504 ,
         \24505 , \24506 , \24507 , \24508 , \24509 , \24510 , \24511 , \24512 , \24513 , \24514 ,
         \24515 , \24516 , \24517 , \24518 , \24519 , \24520 , \24521 , \24522 , \24523 , \24524 ,
         \24525 , \24526 , \24527 , \24528 , \24529 , \24530 , \24531 , \24532 , \24533 , \24534 ,
         \24535 , \24536 , \24537 , \24538 , \24539 , \24540 , \24541 , \24542 , \24543 , \24544 ,
         \24545 , \24546 , \24547 , \24548 , \24549 , \24550 , \24551 , \24552 , \24553 , \24554 ,
         \24555 , \24556 , \24557 , \24558 , \24559 , \24560 , \24561 , \24562 , \24563 , \24564 ,
         \24565 , \24566 , \24567 , \24568 , \24569 , \24570 , \24571 , \24572 , \24573 , \24574 ,
         \24575 , \24576 , \24577 , \24578 , \24579 , \24580 , \24581 , \24582 , \24583 , \24584 ,
         \24585 , \24586 , \24587 , \24588 , \24589 , \24590 , \24591 , \24592 , \24593 , \24594 ,
         \24595 , \24596 , \24597 , \24598 , \24599 , \24600 , \24601 , \24602 , \24603 , \24604 ,
         \24605 , \24606 , \24607 , \24608 , \24609 , \24610 , \24611 , \24612 , \24613 , \24614 ,
         \24615 , \24616 , \24617 , \24618 , \24619 , \24620 , \24621 , \24622 , \24623 , \24624 ,
         \24625 , \24626 , \24627 , \24628 , \24629 , \24630 , \24631 , \24632 , \24633 , \24634 ,
         \24635 , \24636 , \24637 , \24638 , \24639 , \24640 , \24641 , \24642 , \24643 , \24644 ,
         \24645 , \24646 , \24647 , \24648 , \24649 , \24650 , \24651 , \24652 , \24653 , \24654 ,
         \24655 , \24656 , \24657 , \24658 , \24659 , \24660 , \24661 , \24662 , \24663 , \24664 ,
         \24665 , \24666 , \24667 , \24668 , \24669 , \24670 , \24671 , \24672 , \24673 , \24674 ,
         \24675 , \24676 , \24677 , \24678 , \24679 , \24680 , \24681 , \24682 , \24683 , \24684 ,
         \24685 , \24686 , \24687 , \24688 , \24689 , \24690 , \24691 , \24692 , \24693 , \24694 ,
         \24695 , \24696 , \24697 , \24698 , \24699 , \24700 , \24701 , \24702 , \24703 , \24704 ,
         \24705 , \24706 , \24707 , \24708 , \24709 , \24710 , \24711 , \24712 , \24713 , \24714 ,
         \24715 , \24716 , \24717 , \24718 , \24719 , \24720 , \24721 , \24722 , \24723 , \24724 ,
         \24725 , \24726 , \24727 , \24728 , \24729 , \24730 , \24731 , \24732 , \24733 , \24734 ,
         \24735 , \24736 , \24737 , \24738 , \24739 , \24740 , \24741 , \24742 , \24743 , \24744 ,
         \24745 , \24746 , \24747 , \24748 , \24749 , \24750 , \24751 , \24752 , \24753 , \24754 ,
         \24755 , \24756 , \24757 , \24758 , \24759 , \24760 , \24761 , \24762 , \24763 , \24764 ,
         \24765 , \24766 , \24767 , \24768 , \24769 , \24770 , \24771 , \24772 , \24773 , \24774 ,
         \24775 , \24776 , \24777 , \24778 , \24779 , \24780 , \24781 , \24782 , \24783 , \24784 ,
         \24785 , \24786 , \24787 , \24788 , \24789 , \24790 , \24791 , \24792 , \24793 , \24794 ,
         \24795 , \24796 , \24797 , \24798 , \24799 , \24800 , \24801 , \24802 , \24803 , \24804 ,
         \24805 , \24806 , \24807 , \24808 , \24809 , \24810 , \24811 , \24812 , \24813 , \24814 ,
         \24815 , \24816 , \24817 , \24818 , \24819 , \24820 , \24821 , \24822 , \24823 , \24824 ,
         \24825 , \24826 , \24827 , \24828 , \24829 , \24830 , \24831 , \24832 , \24833 , \24834 ,
         \24835 , \24836 , \24837 , \24838 , \24839 , \24840 , \24841 , \24842 , \24843 , \24844 ,
         \24845 , \24846 , \24847 , \24848 , \24849 , \24850 , \24851 , \24852 , \24853 , \24854 ,
         \24855 , \24856 , \24857 , \24858 , \24859 , \24860 , \24861 , \24862 , \24863 , \24864 ,
         \24865 , \24866 , \24867 , \24868 , \24869 , \24870 , \24871 , \24872 , \24873 , \24874 ,
         \24875 , \24876 , \24877 , \24878 , \24879 , \24880 , \24881 , \24882 , \24883 , \24884 ,
         \24885 , \24886 , \24887 , \24888 , \24889 , \24890 , \24891 , \24892 , \24893 , \24894 ,
         \24895 , \24896 , \24897 , \24898 , \24899 , \24900 , \24901 , \24902 , \24903 , \24904 ,
         \24905 , \24906 , \24907 , \24908 , \24909 , \24910 , \24911 , \24912 , \24913 , \24914 ,
         \24915 , \24916 , \24917 , \24918 , \24919 , \24920 , \24921 , \24922 , \24923 , \24924 ,
         \24925 , \24926 , \24927 , \24928 , \24929 , \24930 , \24931 , \24932 , \24933 , \24934 ,
         \24935 , \24936 , \24937 , \24938 , \24939 , \24940 , \24941 , \24942 , \24943 , \24944 ,
         \24945 , \24946 , \24947 , \24948 , \24949 , \24950 , \24951 , \24952 , \24953 , \24954 ,
         \24955 , \24956 , \24957 , \24958 , \24959 , \24960 , \24961 , \24962 , \24963 , \24964 ,
         \24965 , \24966 , \24967 , \24968 , \24969 , \24970 , \24971 , \24972 , \24973 , \24974 ,
         \24975 , \24976 , \24977 , \24978 , \24979 , \24980 , \24981 , \24982 , \24983 , \24984 ,
         \24985 , \24986 , \24987 , \24988 , \24989 , \24990 , \24991 , \24992 , \24993 , \24994 ,
         \24995 , \24996 , \24997 , \24998 , \24999 , \25000 , \25001 , \25002 , \25003 , \25004 ,
         \25005 , \25006 , \25007 , \25008 , \25009 , \25010 , \25011 , \25012 , \25013 , \25014 ,
         \25015 , \25016 , \25017 , \25018 , \25019 , \25020 , \25021 , \25022 , \25023 , \25024 ,
         \25025 , \25026 , \25027 , \25028 , \25029 , \25030 , \25031 , \25032 , \25033 , \25034 ,
         \25035 , \25036 , \25037 , \25038 , \25039 , \25040 , \25041 , \25042 , \25043 , \25044 ,
         \25045 , \25046 , \25047 , \25048 , \25049 , \25050 , \25051 , \25052 , \25053 , \25054 ,
         \25055 , \25056 , \25057 , \25058 , \25059 , \25060 , \25061 , \25062 , \25063 , \25064 ,
         \25065 , \25066 , \25067 , \25068 , \25069 , \25070 , \25071 , \25072 , \25073 , \25074 ,
         \25075 , \25076 , \25077 , \25078 , \25079 , \25080 , \25081 , \25082 , \25083 , \25084 ,
         \25085 , \25086 , \25087 , \25088 , \25089 , \25090 , \25091 , \25092 , \25093 , \25094 ,
         \25095 , \25096 , \25097 , \25098 , \25099 , \25100 , \25101 , \25102 , \25103 , \25104 ,
         \25105 , \25106 , \25107 , \25108 , \25109 , \25110 , \25111 , \25112 , \25113 , \25114 ,
         \25115 , \25116 , \25117 , \25118 , \25119 , \25120 , \25121 , \25122 , \25123 , \25124 ,
         \25125 , \25126 , \25127 , \25128 , \25129 , \25130 , \25131 , \25132 , \25133 , \25134 ,
         \25135 , \25136 , \25137 , \25138 , \25139 , \25140 , \25141 , \25142 , \25143 , \25144 ,
         \25145 , \25146 , \25147 , \25148 , \25149 , \25150 , \25151 , \25152 , \25153 , \25154 ,
         \25155 , \25156 , \25157 , \25158 , \25159 , \25160 , \25161 , \25162 , \25163 , \25164 ,
         \25165 , \25166 , \25167 , \25168 , \25169 , \25170 , \25171 , \25172 , \25173 , \25174 ,
         \25175 , \25176 , \25177 , \25178 , \25179 , \25180 , \25181 , \25182 , \25183 , \25184 ,
         \25185 , \25186 , \25187 , \25188 , \25189 , \25190 , \25191 , \25192 , \25193 , \25194 ,
         \25195 , \25196 , \25197 , \25198 , \25199 , \25200 , \25201 , \25202 , \25203 , \25204 ,
         \25205 , \25206 , \25207 , \25208 , \25209 , \25210 , \25211 , \25212 , \25213 , \25214 ,
         \25215 , \25216 , \25217 , \25218 , \25219 , \25220 , \25221 , \25222 , \25223 , \25224 ,
         \25225 , \25226 , \25227 , \25228 , \25229 , \25230 , \25231 , \25232 , \25233 , \25234 ,
         \25235 , \25236 , \25237 , \25238 , \25239 , \25240 , \25241 , \25242 , \25243 , \25244 ,
         \25245 , \25246 , \25247 , \25248 , \25249 , \25250 , \25251 , \25252 , \25253 , \25254 ,
         \25255 , \25256 , \25257 , \25258 , \25259 , \25260 , \25261 , \25262 , \25263 , \25264 ,
         \25265 , \25266 , \25267 , \25268 , \25269 , \25270 , \25271 , \25272 , \25273 , \25274 ,
         \25275 , \25276 , \25277 , \25278 , \25279 , \25280 , \25281 , \25282 , \25283 , \25284 ,
         \25285 , \25286 , \25287 , \25288 , \25289 , \25290 , \25291 , \25292 , \25293 , \25294 ,
         \25295 , \25296 , \25297 , \25298 , \25299 , \25300 , \25301 , \25302 , \25303 , \25304 ,
         \25305 , \25306 , \25307 , \25308 , \25309 , \25310 , \25311 , \25312 , \25313 , \25314 ,
         \25315 , \25316 , \25317 , \25318 , \25319 , \25320 , \25321 , \25322 , \25323 , \25324 ,
         \25325 , \25326 , \25327 , \25328 , \25329 , \25330 , \25331 , \25332 , \25333 , \25334 ,
         \25335 , \25336 , \25337 , \25338 , \25339 , \25340 , \25341 , \25342 , \25343 , \25344 ,
         \25345 , \25346 , \25347 , \25348 , \25349 , \25350 , \25351 , \25352 , \25353 , \25354 ,
         \25355 , \25356 , \25357 , \25358 , \25359 , \25360 , \25361 , \25362 , \25363 , \25364 ,
         \25365 , \25366 , \25367 , \25368 , \25369 , \25370 , \25371 , \25372 , \25373 , \25374 ,
         \25375 , \25376 , \25377 , \25378 , \25379 , \25380 , \25381 , \25382 , \25383 , \25384 ,
         \25385 , \25386 , \25387 , \25388 , \25389 , \25390 , \25391 , \25392 , \25393 , \25394 ,
         \25395 , \25396 , \25397 , \25398 , \25399 , \25400 , \25401 , \25402 , \25403 , \25404 ,
         \25405 , \25406 , \25407 , \25408 , \25409 , \25410 , \25411 , \25412 , \25413 , \25414 ,
         \25415 , \25416 , \25417 , \25418 , \25419 , \25420 , \25421 , \25422 , \25423 , \25424 ,
         \25425 , \25426 , \25427 , \25428 , \25429 , \25430 , \25431 , \25432 , \25433 , \25434 ,
         \25435 , \25436 , \25437 , \25438 , \25439 , \25440 , \25441 , \25442 , \25443 , \25444 ,
         \25445 , \25446 , \25447 , \25448 , \25449 , \25450 , \25451 , \25452 , \25453 , \25454 ,
         \25455 , \25456 , \25457 , \25458 , \25459 , \25460 , \25461 , \25462 , \25463 , \25464 ,
         \25465 , \25466 , \25467 , \25468 , \25469 , \25470 , \25471 , \25472 , \25473 , \25474 ,
         \25475 , \25476 , \25477 , \25478 , \25479 , \25480 , \25481 , \25482 , \25483 , \25484 ,
         \25485 , \25486 , \25487 , \25488 , \25489 , \25490 , \25491 , \25492 , \25493 , \25494 ,
         \25495 , \25496 , \25497 , \25498 , \25499 , \25500 , \25501 , \25502 , \25503 , \25504 ,
         \25505 , \25506 , \25507 , \25508 , \25509 , \25510 , \25511 , \25512 , \25513 , \25514 ,
         \25515 , \25516 , \25517 , \25518 , \25519 , \25520 , \25521 , \25522 , \25523 , \25524 ,
         \25525 , \25526 , \25527 , \25528 , \25529 , \25530 , \25531 , \25532 , \25533 , \25534 ,
         \25535 , \25536 , \25537 , \25538 , \25539 , \25540 , \25541 , \25542 , \25543 , \25544 ,
         \25545 , \25546 , \25547 , \25548 , \25549 , \25550 , \25551 , \25552 , \25553 , \25554 ,
         \25555 , \25556 , \25557 , \25558 , \25559 , \25560 , \25561 , \25562 , \25563 , \25564 ,
         \25565 , \25566 , \25567 , \25568 , \25569 , \25570 , \25571 , \25572 , \25573 , \25574 ,
         \25575 , \25576 , \25577 , \25578 , \25579 , \25580 , \25581 , \25582 , \25583 , \25584 ,
         \25585 , \25586 , \25587 , \25588 , \25589 , \25590 , \25591 , \25592 , \25593 , \25594 ,
         \25595 , \25596 , \25597 , \25598 , \25599 , \25600 , \25601 , \25602 , \25603 , \25604 ,
         \25605 , \25606 , \25607 , \25608 , \25609 , \25610 , \25611 , \25612 , \25613 , \25614 ,
         \25615 , \25616 , \25617 , \25618 , \25619 , \25620 , \25621 , \25622 , \25623 , \25624 ,
         \25625 , \25626 , \25627 , \25628 , \25629 , \25630 , \25631 , \25632 , \25633 , \25634 ,
         \25635 , \25636 , \25637 , \25638 , \25639 , \25640 , \25641 , \25642 , \25643 , \25644 ,
         \25645 , \25646 , \25647 , \25648 , \25649 , \25650 , \25651 , \25652 , \25653 , \25654 ,
         \25655 , \25656 , \25657 , \25658 , \25659 , \25660 , \25661 , \25662 , \25663 , \25664 ,
         \25665 , \25666 , \25667 , \25668 , \25669 , \25670 , \25671 , \25672 , \25673 , \25674 ,
         \25675 , \25676 , \25677 , \25678 , \25679 , \25680 , \25681 , \25682 , \25683 , \25684 ,
         \25685 , \25686 , \25687 , \25688 , \25689 , \25690 , \25691 , \25692 , \25693 , \25694 ,
         \25695 , \25696 , \25697 , \25698 , \25699 , \25700 , \25701 , \25702 , \25703 , \25704 ,
         \25705 , \25706 , \25707 , \25708 , \25709 , \25710 , \25711 , \25712 , \25713 , \25714 ,
         \25715 , \25716 , \25717 , \25718 , \25719 , \25720 , \25721 , \25722 , \25723 , \25724 ,
         \25725 , \25726 , \25727 , \25728 , \25729 , \25730 , \25731 , \25732 , \25733 , \25734 ,
         \25735 , \25736 , \25737 , \25738 , \25739 , \25740 , \25741 , \25742 , \25743 , \25744 ,
         \25745 , \25746 , \25747 , \25748 , \25749 , \25750 , \25751 , \25752 , \25753 , \25754 ,
         \25755 , \25756 , \25757 , \25758 , \25759 , \25760 , \25761 , \25762 , \25763 , \25764 ,
         \25765 , \25766 , \25767 , \25768 , \25769 , \25770 , \25771 , \25772 , \25773 , \25774 ,
         \25775 , \25776 , \25777 , \25778 , \25779 , \25780 , \25781 , \25782 , \25783 , \25784 ,
         \25785 , \25786 , \25787 , \25788 , \25789 , \25790 , \25791 , \25792 , \25793 , \25794 ,
         \25795 , \25796 , \25797 , \25798 , \25799 , \25800 , \25801 , \25802 , \25803 , \25804 ,
         \25805 , \25806 , \25807 , \25808 , \25809 , \25810 , \25811 , \25812 , \25813 , \25814 ,
         \25815 , \25816 , \25817 , \25818 , \25819 , \25820 , \25821 , \25822 , \25823 , \25824 ,
         \25825 , \25826 , \25827 , \25828 , \25829 , \25830 , \25831 , \25832 , \25833 , \25834 ,
         \25835 , \25836 , \25837 , \25838 , \25839 , \25840 , \25841 , \25842 , \25843 , \25844 ,
         \25845 , \25846 , \25847 , \25848 , \25849 , \25850 , \25851 , \25852 , \25853 , \25854 ,
         \25855 , \25856 , \25857 , \25858 , \25859 , \25860 , \25861 , \25862 , \25863 , \25864 ,
         \25865 , \25866 , \25867 , \25868 , \25869 , \25870 , \25871 , \25872 , \25873 , \25874 ,
         \25875 , \25876 , \25877 , \25878 , \25879 , \25880 , \25881 , \25882 , \25883 , \25884 ,
         \25885 , \25886 , \25887 , \25888 , \25889 , \25890 , \25891 , \25892 , \25893 , \25894 ,
         \25895 , \25896 , \25897 , \25898 , \25899 , \25900 , \25901 , \25902 , \25903 , \25904 ,
         \25905 , \25906 , \25907 , \25908 , \25909 , \25910 , \25911 , \25912 , \25913 , \25914 ,
         \25915 , \25916 , \25917 , \25918 , \25919 , \25920 , \25921 , \25922 , \25923 , \25924 ,
         \25925 , \25926 , \25927 , \25928 , \25929 , \25930 , \25931 , \25932 , \25933 , \25934 ,
         \25935 , \25936 , \25937 , \25938 , \25939 , \25940 , \25941 , \25942 , \25943 , \25944 ,
         \25945 , \25946 , \25947 , \25948 , \25949 , \25950 , \25951 , \25952 , \25953 , \25954 ,
         \25955 , \25956 , \25957 , \25958 , \25959 , \25960 , \25961 , \25962 , \25963 , \25964 ,
         \25965 , \25966 , \25967 , \25968 , \25969 , \25970 , \25971 , \25972 , \25973 , \25974 ,
         \25975 , \25976 , \25977 , \25978 , \25979 , \25980 , \25981 , \25982 , \25983 , \25984 ,
         \25985 , \25986 , \25987 , \25988 , \25989 , \25990 , \25991 , \25992 , \25993 , \25994 ,
         \25995 , \25996 , \25997 , \25998 , \25999 , \26000 , \26001 , \26002 , \26003 , \26004 ,
         \26005 , \26006 , \26007 , \26008 , \26009 , \26010 , \26011 , \26012 , \26013 , \26014 ,
         \26015 , \26016 , \26017 , \26018 , \26019 , \26020 , \26021 , \26022 , \26023 , \26024 ,
         \26025 , \26026 , \26027 , \26028 , \26029 , \26030 , \26031 , \26032 , \26033 , \26034 ,
         \26035 , \26036 , \26037 , \26038 , \26039 , \26040 , \26041 , \26042 , \26043 , \26044 ,
         \26045 , \26046 , \26047 , \26048 , \26049 , \26050 , \26051 , \26052 , \26053 , \26054 ,
         \26055 , \26056 , \26057 , \26058 , \26059 , \26060 , \26061 , \26062 , \26063 , \26064 ,
         \26065 , \26066 , \26067 , \26068 , \26069 , \26070 , \26071 , \26072 , \26073 , \26074 ,
         \26075 , \26076 , \26077 , \26078 , \26079 , \26080 , \26081 , \26082 , \26083 , \26084 ,
         \26085 , \26086 , \26087 , \26088 , \26089 , \26090 , \26091 , \26092 , \26093 , \26094 ,
         \26095 , \26096 , \26097 , \26098 , \26099 , \26100 , \26101 , \26102 , \26103 , \26104 ,
         \26105 , \26106 , \26107 , \26108 , \26109 , \26110 , \26111 , \26112 , \26113 , \26114 ,
         \26115 , \26116 , \26117 , \26118 , \26119 , \26120 , \26121 , \26122 , \26123 , \26124 ,
         \26125 , \26126 , \26127 , \26128 , \26129 , \26130 , \26131 , \26132 , \26133 , \26134 ,
         \26135 , \26136 , \26137 , \26138 , \26139 , \26140 , \26141 , \26142 , \26143 , \26144 ,
         \26145 , \26146 , \26147 , \26148 , \26149 , \26150 , \26151 , \26152 , \26153 , \26154 ,
         \26155 , \26156 , \26157 , \26158 , \26159 , \26160 , \26161 , \26162 , \26163 , \26164 ,
         \26165 , \26166 , \26167 , \26168 , \26169 , \26170 , \26171 , \26172 , \26173 , \26174 ,
         \26175 , \26176 , \26177 , \26178 , \26179 , \26180 , \26181 , \26182 , \26183 , \26184 ,
         \26185 , \26186 , \26187 , \26188 , \26189 , \26190 , \26191 , \26192 , \26193 , \26194 ,
         \26195 , \26196 , \26197 , \26198 , \26199 , \26200 , \26201 , \26202 , \26203 , \26204 ,
         \26205 , \26206 , \26207 , \26208 , \26209 , \26210 , \26211 , \26212 , \26213 , \26214 ,
         \26215 , \26216 , \26217 , \26218 , \26219 , \26220 , \26221 , \26222 , \26223 , \26224 ,
         \26225 , \26226 , \26227 , \26228 , \26229 , \26230 , \26231 , \26232 , \26233 , \26234 ,
         \26235 , \26236 , \26237 , \26238 , \26239 , \26240 , \26241 , \26242 , \26243 , \26244 ,
         \26245 , \26246 , \26247 , \26248 , \26249 , \26250 , \26251 , \26252 , \26253 , \26254 ,
         \26255 , \26256 , \26257 , \26258 , \26259 , \26260 , \26261 , \26262 , \26263 , \26264 ,
         \26265 , \26266 , \26267 , \26268 , \26269 , \26270 , \26271 , \26272 , \26273 , \26274 ,
         \26275 , \26276 , \26277 , \26278 , \26279 , \26280 , \26281 , \26282 , \26283 , \26284 ,
         \26285 , \26286 , \26287 , \26288 , \26289 , \26290 , \26291 , \26292 , \26293 , \26294 ,
         \26295 , \26296 , \26297 , \26298 , \26299 , \26300 , \26301 , \26302 , \26303 , \26304 ,
         \26305 , \26306 , \26307 , \26308 , \26309 , \26310 , \26311 , \26312 , \26313 , \26314 ,
         \26315 , \26316 , \26317 , \26318 , \26319 , \26320 , \26321 , \26322 , \26323 , \26324 ,
         \26325 , \26326 , \26327 , \26328 , \26329 , \26330 , \26331 , \26332 , \26333 , \26334 ,
         \26335 , \26336 , \26337 , \26338 , \26339 , \26340 , \26341 , \26342 , \26343 , \26344 ,
         \26345 , \26346 , \26347 , \26348 , \26349 , \26350 , \26351 , \26352 , \26353 , \26354 ,
         \26355 , \26356 , \26357 , \26358 , \26359 , \26360 , \26361 , \26362 , \26363 , \26364 ,
         \26365 , \26366 , \26367 , \26368 , \26369 , \26370 , \26371 , \26372 , \26373 , \26374 ,
         \26375 , \26376 , \26377 , \26378 , \26379 , \26380 , \26381 , \26382 , \26383 , \26384 ,
         \26385 , \26386 , \26387 , \26388 , \26389 , \26390 , \26391 , \26392 , \26393 , \26394 ,
         \26395 , \26396 , \26397 , \26398 , \26399 , \26400 , \26401 , \26402 , \26403 , \26404 ,
         \26405 , \26406 , \26407 , \26408 , \26409 , \26410 , \26411 , \26412 , \26413 , \26414 ,
         \26415 , \26416 , \26417 , \26418 , \26419 , \26420 , \26421 , \26422 , \26423 , \26424 ,
         \26425 , \26426 , \26427 , \26428 , \26429 , \26430 , \26431 , \26432 , \26433 , \26434 ,
         \26435 , \26436 , \26437 , \26438 , \26439 , \26440 , \26441 , \26442 , \26443 , \26444 ,
         \26445 , \26446 , \26447 , \26448 , \26449 , \26450 , \26451 , \26452 , \26453 , \26454 ,
         \26455 , \26456 , \26457 , \26458 , \26459 , \26460 , \26461 , \26462 , \26463 , \26464 ,
         \26465 , \26466 , \26467 , \26468 , \26469 , \26470 , \26471 , \26472 , \26473 , \26474 ,
         \26475 , \26476 , \26477 , \26478 , \26479 , \26480 , \26481 , \26482 , \26483 , \26484 ,
         \26485 , \26486 , \26487 , \26488 , \26489 , \26490 , \26491 , \26492 , \26493 , \26494 ,
         \26495 , \26496 , \26497 , \26498 , \26499 , \26500 , \26501 , \26502 , \26503 , \26504 ,
         \26505 , \26506 , \26507 , \26508 , \26509 , \26510 , \26511 , \26512 , \26513 , \26514 ,
         \26515 , \26516 , \26517 , \26518 , \26519 , \26520 , \26521 , \26522 , \26523 , \26524 ,
         \26525 , \26526 , \26527 , \26528 , \26529 , \26530 , \26531 , \26532 , \26533 , \26534 ,
         \26535 , \26536 , \26537 , \26538 , \26539 , \26540 , \26541 , \26542 , \26543 , \26544 ,
         \26545 , \26546 , \26547 , \26548 , \26549 , \26550 , \26551 , \26552 , \26553 , \26554 ,
         \26555 , \26556 , \26557 , \26558 , \26559 , \26560 , \26561 , \26562 , \26563 , \26564 ,
         \26565 , \26566 , \26567 , \26568 , \26569 , \26570 , \26571 , \26572 , \26573 , \26574 ,
         \26575 , \26576 , \26577 , \26578 , \26579 , \26580 , \26581 , \26582 , \26583 , \26584 ,
         \26585 , \26586 , \26587 , \26588 , \26589 , \26590 , \26591 , \26592 , \26593 , \26594 ,
         \26595 , \26596 , \26597 , \26598 , \26599 , \26600 , \26601 , \26602 , \26603 , \26604 ,
         \26605 , \26606 , \26607 , \26608 , \26609 , \26610 , \26611 , \26612 , \26613 , \26614 ,
         \26615 , \26616 , \26617 , \26618 , \26619 , \26620 , \26621 , \26622 , \26623 , \26624 ,
         \26625 , \26626 , \26627 , \26628 , \26629 , \26630 , \26631 , \26632 , \26633 , \26634 ,
         \26635 , \26636 , \26637 , \26638 , \26639 , \26640 , \26641 , \26642 , \26643 , \26644 ,
         \26645 , \26646 , \26647 , \26648 , \26649 , \26650 , \26651 , \26652 , \26653 , \26654 ,
         \26655 , \26656 , \26657 , \26658 , \26659 , \26660 , \26661 , \26662 , \26663 , \26664 ,
         \26665 , \26666 , \26667 , \26668 , \26669 , \26670 , \26671 , \26672 , \26673 , \26674 ,
         \26675 , \26676 , \26677 , \26678 , \26679 , \26680 , \26681 , \26682 , \26683 , \26684 ,
         \26685 , \26686 , \26687 , \26688 , \26689 , \26690 , \26691 , \26692 , \26693 , \26694 ,
         \26695 , \26696 , \26697 , \26698 , \26699 , \26700 , \26701 , \26702 , \26703 , \26704 ,
         \26705 , \26706 , \26707 , \26708 , \26709 , \26710 , \26711 , \26712 , \26713 , \26714 ,
         \26715 , \26716 , \26717 , \26718 , \26719 , \26720 , \26721 , \26722 , \26723 , \26724 ,
         \26725 , \26726 , \26727 , \26728 , \26729 , \26730 , \26731 , \26732 , \26733 , \26734 ,
         \26735 , \26736 , \26737 , \26738 , \26739 , \26740 , \26741 , \26742 , \26743 , \26744 ,
         \26745 , \26746 , \26747 , \26748 , \26749 , \26750 , \26751 , \26752 , \26753 , \26754 ,
         \26755 , \26756 , \26757 , \26758 , \26759 , \26760 , \26761 , \26762 , \26763 , \26764 ,
         \26765 , \26766 , \26767 , \26768 , \26769 , \26770 , \26771 , \26772 , \26773 , \26774 ,
         \26775 , \26776 , \26777 , \26778 , \26779 , \26780 , \26781 , \26782 , \26783 , \26784 ,
         \26785 , \26786 , \26787 , \26788 , \26789 , \26790 , \26791 , \26792 , \26793 , \26794 ,
         \26795 , \26796 , \26797 , \26798 , \26799 , \26800 , \26801 , \26802 , \26803 , \26804 ,
         \26805 , \26806 , \26807 , \26808 , \26809 , \26810 , \26811 , \26812 , \26813 , \26814 ,
         \26815 , \26816 , \26817 , \26818 , \26819 , \26820 , \26821 , \26822 , \26823 , \26824 ,
         \26825 , \26826 , \26827 , \26828 , \26829 , \26830 , \26831 , \26832 , \26833 , \26834 ,
         \26835 , \26836 , \26837 , \26838 , \26839 , \26840 , \26841 , \26842 , \26843 , \26844 ,
         \26845 , \26846 , \26847 , \26848 , \26849 , \26850 , \26851 , \26852 , \26853 , \26854 ,
         \26855 , \26856 , \26857 , \26858 , \26859 , \26860 , \26861 , \26862 , \26863 , \26864 ,
         \26865 , \26866 , \26867 , \26868 , \26869 , \26870 , \26871 , \26872 , \26873 , \26874 ,
         \26875 , \26876 , \26877 , \26878 , \26879 , \26880 , \26881 , \26882 , \26883 , \26884 ,
         \26885 , \26886 , \26887 , \26888 , \26889 , \26890 , \26891 , \26892 , \26893 , \26894 ,
         \26895 , \26896 , \26897 , \26898 , \26899 , \26900 , \26901 , \26902 , \26903 , \26904 ,
         \26905 , \26906 , \26907 , \26908 , \26909 , \26910 , \26911 , \26912 , \26913 , \26914 ,
         \26915 , \26916 , \26917 , \26918 , \26919 , \26920 , \26921 , \26922 , \26923 , \26924 ,
         \26925 , \26926 , \26927 , \26928 , \26929 , \26930 , \26931 , \26932 , \26933 , \26934 ,
         \26935 , \26936 , \26937 , \26938 , \26939 , \26940 , \26941 , \26942 , \26943 , \26944 ,
         \26945 , \26946 , \26947 , \26948 , \26949 , \26950 , \26951 , \26952 , \26953 , \26954 ,
         \26955 , \26956 , \26957 , \26958 , \26959 , \26960 , \26961 , \26962 , \26963 , \26964 ,
         \26965 , \26966 , \26967 , \26968 , \26969 , \26970 , \26971 , \26972 , \26973 , \26974 ,
         \26975 , \26976 , \26977 , \26978 , \26979 , \26980 , \26981 , \26982 , \26983 , \26984 ,
         \26985 , \26986 , \26987 , \26988 , \26989 , \26990 , \26991 , \26992 , \26993 , \26994 ,
         \26995 , \26996 , \26997 , \26998 , \26999 , \27000 , \27001 , \27002 , \27003 , \27004 ,
         \27005 , \27006 , \27007 , \27008 , \27009 , \27010 , \27011 , \27012 , \27013 , \27014 ,
         \27015 , \27016 , \27017 , \27018 , \27019 , \27020 , \27021 , \27022 , \27023 , \27024 ,
         \27025 , \27026 , \27027 , \27028 , \27029 , \27030 , \27031 , \27032 , \27033 , \27034 ,
         \27035 , \27036 , \27037 , \27038 , \27039 , \27040 , \27041 , \27042 , \27043 , \27044 ,
         \27045 , \27046 , \27047 , \27048 , \27049 , \27050 , \27051 , \27052 , \27053 , \27054 ,
         \27055 , \27056 , \27057 , \27058 , \27059 , \27060 , \27061 , \27062 , \27063 , \27064 ,
         \27065 , \27066 , \27067 , \27068 , \27069 , \27070 , \27071 , \27072 , \27073 , \27074 ,
         \27075 , \27076 , \27077 , \27078 , \27079 , \27080 , \27081 , \27082 , \27083 , \27084 ,
         \27085 , \27086 , \27087 , \27088 , \27089 , \27090 , \27091 , \27092 , \27093 , \27094 ,
         \27095 , \27096 , \27097 , \27098 , \27099 , \27100 , \27101 , \27102 , \27103 , \27104 ,
         \27105 , \27106 , \27107 , \27108 , \27109 , \27110 , \27111 , \27112 , \27113 , \27114 ,
         \27115 , \27116 , \27117 , \27118 , \27119 , \27120 , \27121 , \27122 , \27123 , \27124 ,
         \27125 , \27126 , \27127 , \27128 , \27129 , \27130 , \27131 , \27132 , \27133 , \27134 ,
         \27135 , \27136 , \27137 , \27138 , \27139 , \27140 , \27141 , \27142 , \27143 , \27144 ,
         \27145 , \27146 , \27147 , \27148 , \27149 , \27150 , \27151 , \27152 , \27153 , \27154 ,
         \27155 , \27156 , \27157 , \27158 , \27159 , \27160 , \27161 , \27162 , \27163 , \27164 ,
         \27165 , \27166 , \27167 , \27168 , \27169 , \27170 , \27171 , \27172 , \27173 , \27174 ,
         \27175 , \27176 , \27177 , \27178 , \27179 , \27180 , \27181 , \27182 , \27183 , \27184 ,
         \27185 , \27186 , \27187 , \27188 , \27189 , \27190 , \27191 , \27192 , \27193 , \27194 ,
         \27195 , \27196 , \27197 , \27198 , \27199 , \27200 , \27201 , \27202 , \27203 , \27204 ,
         \27205 , \27206 , \27207 , \27208 , \27209 , \27210 , \27211 , \27212 , \27213 , \27214 ,
         \27215 , \27216 , \27217 , \27218 , \27219 , \27220 , \27221 , \27222 , \27223 , \27224 ,
         \27225 , \27226 , \27227 , \27228 , \27229 , \27230 , \27231 , \27232 , \27233 , \27234 ,
         \27235 , \27236 , \27237 , \27238 , \27239 , \27240 , \27241 , \27242 , \27243 , \27244 ,
         \27245 , \27246 , \27247 , \27248 , \27249 , \27250 , \27251 , \27252 , \27253 , \27254 ,
         \27255 , \27256 , \27257 , \27258 , \27259 , \27260 , \27261 , \27262 , \27263 , \27264 ,
         \27265 , \27266 , \27267 , \27268 , \27269 , \27270 , \27271 , \27272 , \27273 , \27274 ,
         \27275 , \27276 , \27277 , \27278 , \27279 , \27280 , \27281 , \27282 , \27283 , \27284 ,
         \27285 , \27286 , \27287 , \27288 , \27289 , \27290 , \27291 , \27292 , \27293 , \27294 ,
         \27295 , \27296 , \27297 , \27298 , \27299 , \27300 , \27301 , \27302 , \27303 , \27304 ,
         \27305 , \27306 , \27307 , \27308 , \27309 , \27310 , \27311 , \27312 , \27313 , \27314 ,
         \27315 , \27316 , \27317 , \27318 , \27319 , \27320 , \27321 , \27322 , \27323 , \27324 ,
         \27325 , \27326 , \27327 , \27328 , \27329 , \27330 , \27331 , \27332 , \27333 , \27334 ,
         \27335 , \27336 , \27337 , \27338 , \27339 , \27340 , \27341 , \27342 , \27343 , \27344 ,
         \27345 , \27346 , \27347 , \27348 , \27349 , \27350 , \27351 , \27352 , \27353 , \27354 ,
         \27355 , \27356 , \27357 , \27358 , \27359 , \27360 , \27361 , \27362 , \27363 , \27364 ,
         \27365 , \27366 , \27367 , \27368 , \27369 , \27370 , \27371 , \27372 , \27373 , \27374 ,
         \27375 , \27376 , \27377 , \27378 , \27379 , \27380 , \27381 , \27382 , \27383 , \27384 ,
         \27385 , \27386 , \27387 , \27388 , \27389 , \27390 , \27391 , \27392 , \27393 , \27394 ,
         \27395 , \27396 , \27397 , \27398 , \27399 , \27400 , \27401 , \27402 , \27403 , \27404 ,
         \27405 , \27406 , \27407 , \27408 , \27409 , \27410 , \27411 , \27412 , \27413 , \27414 ,
         \27415 , \27416 , \27417 , \27418 , \27419 , \27420 , \27421 , \27422 , \27423 , \27424 ,
         \27425 , \27426 , \27427 , \27428 , \27429 , \27430 , \27431 , \27432 , \27433 , \27434 ,
         \27435 , \27436 , \27437 , \27438 , \27439 , \27440 , \27441 , \27442 , \27443 , \27444 ,
         \27445 , \27446 , \27447 , \27448 , \27449 , \27450 , \27451 , \27452 , \27453 , \27454 ,
         \27455 , \27456 , \27457 , \27458 , \27459 , \27460 , \27461 , \27462 , \27463 , \27464 ,
         \27465 , \27466 , \27467 , \27468 , \27469 , \27470 , \27471 , \27472 , \27473 , \27474 ,
         \27475 , \27476 , \27477 , \27478 , \27479 , \27480 , \27481 , \27482 , \27483 , \27484 ,
         \27485 , \27486 , \27487 , \27488 , \27489 , \27490 , \27491 , \27492 , \27493 , \27494 ,
         \27495 , \27496 , \27497 , \27498 , \27499 , \27500 , \27501 , \27502 , \27503 , \27504 ,
         \27505 , \27506 , \27507 , \27508 , \27509 , \27510 , \27511 , \27512 , \27513 , \27514 ,
         \27515 , \27516 , \27517 , \27518 , \27519 , \27520 , \27521 , \27522 , \27523 , \27524 ,
         \27525 , \27526 , \27527 , \27528 , \27529 , \27530 , \27531 , \27532 , \27533 , \27534 ,
         \27535 , \27536 , \27537 , \27538 , \27539 , \27540 , \27541 , \27542 , \27543 , \27544 ,
         \27545 , \27546 , \27547 , \27548 , \27549 , \27550 , \27551 , \27552 , \27553 , \27554 ,
         \27555 , \27556 , \27557 , \27558 , \27559 , \27560 , \27561 , \27562 , \27563 , \27564 ,
         \27565 , \27566 , \27567 , \27568 , \27569 , \27570 , \27571 , \27572 , \27573 , \27574 ,
         \27575 , \27576 , \27577 , \27578 , \27579 , \27580 , \27581 , \27582 , \27583 , \27584 ,
         \27585 , \27586 , \27587 , \27588 , \27589 , \27590 , \27591 , \27592 , \27593 , \27594 ,
         \27595 , \27596 , \27597 , \27598 , \27599 , \27600 , \27601 , \27602 , \27603 , \27604 ,
         \27605 , \27606 , \27607 , \27608 , \27609 , \27610 , \27611 , \27612 , \27613 , \27614 ,
         \27615 , \27616 , \27617 , \27618 , \27619 , \27620 , \27621 , \27622 , \27623 , \27624 ,
         \27625 , \27626 , \27627 , \27628 , \27629 , \27630 , \27631 , \27632 , \27633 , \27634 ,
         \27635 , \27636 , \27637 , \27638 , \27639 , \27640 , \27641 , \27642 , \27643 , \27644 ,
         \27645 , \27646 , \27647 , \27648 , \27649 , \27650 , \27651 , \27652 , \27653 , \27654 ,
         \27655 , \27656 , \27657 , \27658 , \27659 , \27660 , \27661 , \27662 , \27663 , \27664 ,
         \27665 , \27666 , \27667 , \27668 , \27669 , \27670 , \27671 , \27672 , \27673 , \27674 ,
         \27675 , \27676 , \27677 , \27678 , \27679 , \27680 , \27681 , \27682 , \27683 , \27684 ,
         \27685 , \27686 , \27687 , \27688 , \27689 , \27690 , \27691 , \27692 , \27693 , \27694 ,
         \27695 , \27696 , \27697 , \27698 , \27699 , \27700 , \27701 , \27702 , \27703 , \27704 ,
         \27705 , \27706 , \27707 , \27708 , \27709 , \27710 , \27711 , \27712 , \27713 , \27714 ,
         \27715 , \27716 , \27717 , \27718 , \27719 , \27720 , \27721 , \27722 , \27723 , \27724 ,
         \27725 , \27726 , \27727 , \27728 , \27729 , \27730 , \27731 , \27732 , \27733 , \27734 ,
         \27735 , \27736 , \27737 , \27738 , \27739 , \27740 , \27741 , \27742 , \27743 , \27744 ,
         \27745 , \27746 , \27747 , \27748 , \27749 , \27750 , \27751 , \27752 , \27753 , \27754 ,
         \27755 , \27756 , \27757 , \27758 , \27759 , \27760 , \27761 , \27762 , \27763 , \27764 ,
         \27765 , \27766 , \27767 , \27768 , \27769 , \27770 , \27771 , \27772 , \27773 , \27774 ,
         \27775 , \27776 , \27777 , \27778 , \27779 , \27780 , \27781 , \27782 , \27783 , \27784 ,
         \27785 , \27786 , \27787 , \27788 , \27789 , \27790 , \27791 , \27792 , \27793 , \27794 ,
         \27795 , \27796 , \27797 , \27798 , \27799 , \27800 , \27801 , \27802 , \27803 , \27804 ,
         \27805 , \27806 , \27807 , \27808 , \27809 , \27810 , \27811 , \27812 , \27813 , \27814 ,
         \27815 , \27816 , \27817 , \27818 , \27819 , \27820 , \27821 , \27822 , \27823 , \27824 ,
         \27825 , \27826 , \27827 , \27828 , \27829 , \27830 , \27831 , \27832 , \27833 , \27834 ,
         \27835 , \27836 , \27837 , \27838 , \27839 , \27840 , \27841 , \27842 , \27843 , \27844 ,
         \27845 , \27846 , \27847 , \27848 , \27849 , \27850 , \27851 , \27852 , \27853 , \27854 ,
         \27855 , \27856 , \27857 , \27858 , \27859 , \27860 , \27861 , \27862 , \27863 , \27864 ,
         \27865 , \27866 , \27867 , \27868 , \27869 , \27870 , \27871 , \27872 , \27873 , \27874 ,
         \27875 , \27876 , \27877 , \27878 , \27879 , \27880 , \27881 , \27882 , \27883 , \27884 ,
         \27885 , \27886 , \27887 , \27888 , \27889 , \27890 , \27891 , \27892 , \27893 , \27894 ,
         \27895 , \27896 , \27897 , \27898 , \27899 , \27900 , \27901 , \27902 , \27903 , \27904 ,
         \27905 , \27906 , \27907 , \27908 , \27909 , \27910 , \27911 , \27912 , \27913 , \27914 ,
         \27915 , \27916 , \27917 , \27918 , \27919 , \27920 , \27921 , \27922 , \27923 , \27924 ,
         \27925 , \27926 , \27927 , \27928 , \27929 , \27930 , \27931 , \27932 , \27933 , \27934 ,
         \27935 , \27936 , \27937 , \27938 , \27939 , \27940 , \27941 , \27942 , \27943 , \27944 ,
         \27945 , \27946 , \27947 , \27948 , \27949 , \27950 , \27951 , \27952 , \27953 , \27954 ,
         \27955 , \27956 , \27957 , \27958 , \27959 , \27960 , \27961 , \27962 , \27963 , \27964 ,
         \27965 , \27966 , \27967 , \27968 , \27969 , \27970 , \27971 , \27972 , \27973 , \27974 ,
         \27975 , \27976 , \27977 , \27978 , \27979 , \27980 , \27981 , \27982 , \27983 , \27984 ,
         \27985 , \27986 , \27987 , \27988 , \27989 , \27990 , \27991 , \27992 , \27993 , \27994 ,
         \27995 , \27996 , \27997 , \27998 , \27999 , \28000 , \28001 , \28002 , \28003 , \28004 ,
         \28005 , \28006 , \28007 , \28008 , \28009 , \28010 , \28011 , \28012 , \28013 , \28014 ,
         \28015 , \28016 , \28017 , \28018 , \28019 , \28020 , \28021 , \28022 , \28023 , \28024 ,
         \28025 , \28026 , \28027 , \28028 , \28029 , \28030 , \28031 , \28032 , \28033 , \28034 ,
         \28035 , \28036 , \28037 , \28038 , \28039 , \28040 , \28041 , \28042 , \28043 , \28044 ,
         \28045 , \28046 , \28047 , \28048 , \28049 , \28050 , \28051 , \28052 , \28053 , \28054 ,
         \28055 , \28056 , \28057 , \28058 , \28059 , \28060 , \28061 , \28062 , \28063 , \28064 ,
         \28065 , \28066 , \28067 , \28068 , \28069 , \28070 , \28071 , \28072 , \28073 , \28074 ,
         \28075 , \28076 , \28077 , \28078 , \28079 , \28080 , \28081 , \28082 , \28083 , \28084 ,
         \28085 , \28086 , \28087 , \28088 , \28089 , \28090 , \28091 , \28092 , \28093 , \28094 ,
         \28095 , \28096 , \28097 , \28098 , \28099 , \28100 , \28101 , \28102 , \28103 , \28104 ,
         \28105 , \28106 , \28107 , \28108 , \28109 , \28110 , \28111 , \28112 , \28113 , \28114 ,
         \28115 , \28116 , \28117 , \28118 , \28119 , \28120 , \28121 , \28122 , \28123 , \28124 ,
         \28125 , \28126 , \28127 , \28128 , \28129 , \28130 , \28131 , \28132 , \28133 , \28134 ,
         \28135 , \28136 , \28137 , \28138 , \28139 , \28140 , \28141 , \28142 , \28143 , \28144 ,
         \28145 , \28146 , \28147 , \28148 , \28149 , \28150 , \28151 , \28152 , \28153 , \28154 ,
         \28155 , \28156 , \28157 , \28158 , \28159 , \28160 , \28161 , \28162 , \28163 , \28164 ,
         \28165 , \28166 , \28167 , \28168 , \28169 , \28170 , \28171 , \28172 , \28173 , \28174 ,
         \28175 , \28176 , \28177 , \28178 , \28179 , \28180 , \28181 , \28182 , \28183 , \28184 ,
         \28185 , \28186 , \28187 , \28188 , \28189 , \28190 , \28191 , \28192 , \28193 , \28194 ,
         \28195 , \28196 , \28197 , \28198 , \28199 , \28200 , \28201 , \28202 , \28203 , \28204 ,
         \28205 , \28206 , \28207 , \28208 , \28209 , \28210 , \28211 , \28212 , \28213 , \28214 ,
         \28215 , \28216 , \28217 , \28218 , \28219 , \28220 , \28221 , \28222 , \28223 , \28224 ,
         \28225 , \28226 , \28227 , \28228 , \28229 , \28230 , \28231 , \28232 , \28233 , \28234 ,
         \28235 , \28236 , \28237 , \28238 , \28239 , \28240 , \28241 , \28242 , \28243 , \28244 ,
         \28245 , \28246 , \28247 , \28248 , \28249 , \28250 , \28251 , \28252 , \28253 , \28254 ,
         \28255 , \28256 , \28257 , \28258 , \28259 , \28260 , \28261 , \28262 , \28263 , \28264 ,
         \28265 , \28266 , \28267 , \28268 , \28269 , \28270 , \28271 , \28272 , \28273 , \28274 ,
         \28275 , \28276 , \28277 , \28278 , \28279 , \28280 , \28281 , \28282 , \28283 , \28284 ,
         \28285 , \28286 , \28287 , \28288 , \28289 , \28290 , \28291 , \28292 , \28293 , \28294 ,
         \28295 , \28296 , \28297 , \28298 , \28299 , \28300 , \28301 , \28302 , \28303 , \28304 ,
         \28305 , \28306 , \28307 , \28308 , \28309 , \28310 , \28311 , \28312 , \28313 , \28314 ,
         \28315 , \28316 , \28317 , \28318 , \28319 , \28320 , \28321 , \28322 , \28323 , \28324 ,
         \28325 , \28326 , \28327 , \28328 , \28329 , \28330 , \28331 , \28332 , \28333 , \28334 ,
         \28335 , \28336 , \28337 , \28338 , \28339 , \28340 , \28341 , \28342 , \28343 , \28344 ,
         \28345 , \28346 , \28347 , \28348 , \28349 , \28350 , \28351 , \28352 , \28353 , \28354 ,
         \28355 , \28356 , \28357 , \28358 , \28359 , \28360 , \28361 , \28362 , \28363 , \28364 ,
         \28365 , \28366 , \28367 , \28368 , \28369 , \28370 , \28371 , \28372 , \28373 , \28374 ,
         \28375 , \28376 , \28377 , \28378 , \28379 , \28380 , \28381 , \28382 , \28383 , \28384 ,
         \28385 , \28386 , \28387 , \28388 , \28389 , \28390 , \28391 , \28392 , \28393 , \28394 ,
         \28395 , \28396 , \28397 , \28398 , \28399 , \28400 , \28401 , \28402 , \28403 , \28404 ,
         \28405 , \28406 , \28407 , \28408 , \28409 , \28410 , \28411 , \28412 , \28413 , \28414 ,
         \28415 , \28416 , \28417 , \28418 , \28419 , \28420 , \28421 , \28422 , \28423 , \28424 ,
         \28425 , \28426 , \28427 , \28428 , \28429 , \28430 , \28431 , \28432 , \28433 , \28434 ,
         \28435 , \28436 , \28437 , \28438 , \28439 , \28440 , \28441 , \28442 , \28443 , \28444 ,
         \28445 , \28446 , \28447 , \28448 , \28449 , \28450 , \28451 , \28452 , \28453 , \28454 ,
         \28455 , \28456 , \28457 , \28458 , \28459 , \28460 , \28461 , \28462 , \28463 , \28464 ,
         \28465 , \28466 , \28467 , \28468 , \28469 , \28470 , \28471 , \28472 , \28473 , \28474 ,
         \28475 , \28476 , \28477 , \28478 , \28479 , \28480 , \28481 , \28482 , \28483 , \28484 ,
         \28485 , \28486 , \28487 , \28488 , \28489 , \28490 , \28491 , \28492 , \28493 , \28494 ,
         \28495 , \28496 , \28497 , \28498 , \28499 , \28500 , \28501 , \28502 , \28503 , \28504 ,
         \28505 , \28506 , \28507 , \28508 , \28509 , \28510 , \28511 , \28512 , \28513 , \28514 ,
         \28515 , \28516 , \28517 , \28518 , \28519 , \28520 , \28521 , \28522 , \28523 , \28524 ,
         \28525 , \28526 , \28527 , \28528 , \28529 , \28530 , \28531 , \28532 , \28533 , \28534 ,
         \28535 , \28536 , \28537 , \28538 , \28539 , \28540 , \28541 , \28542 , \28543 , \28544 ,
         \28545 , \28546 , \28547 , \28548 , \28549 , \28550 , \28551 , \28552 , \28553 , \28554 ,
         \28555 , \28556 , \28557 , \28558 , \28559 , \28560 , \28561 , \28562 , \28563 , \28564 ,
         \28565 , \28566 , \28567 , \28568 , \28569 , \28570 , \28571 , \28572 , \28573 , \28574 ,
         \28575 , \28576 , \28577 , \28578 , \28579 , \28580 , \28581 , \28582 , \28583 , \28584 ,
         \28585 , \28586 , \28587 , \28588 , \28589 , \28590 , \28591 , \28592 , \28593 , \28594 ,
         \28595 , \28596 , \28597 , \28598 , \28599 , \28600 , \28601 , \28602 , \28603 , \28604 ,
         \28605 , \28606 , \28607 , \28608 , \28609 , \28610 , \28611 , \28612 , \28613 , \28614 ,
         \28615 , \28616 , \28617 , \28618 , \28619 , \28620 , \28621 , \28622 , \28623 , \28624 ,
         \28625 , \28626 , \28627 , \28628 , \28629 , \28630 , \28631 , \28632 , \28633 , \28634 ,
         \28635 , \28636 , \28637 , \28638 , \28639 , \28640 , \28641 , \28642 , \28643 , \28644 ,
         \28645 , \28646 , \28647 , \28648 , \28649 , \28650 , \28651 , \28652 , \28653 , \28654 ,
         \28655 , \28656 , \28657 , \28658 , \28659 , \28660 , \28661 , \28662 , \28663 , \28664 ,
         \28665 , \28666 , \28667 , \28668 , \28669 , \28670 , \28671 , \28672 , \28673 , \28674 ,
         \28675 , \28676 , \28677 , \28678 , \28679 , \28680 , \28681 , \28682 , \28683 , \28684 ,
         \28685 , \28686 , \28687 , \28688 , \28689 , \28690 , \28691 , \28692 , \28693 , \28694 ,
         \28695 , \28696 , \28697 , \28698 , \28699 , \28700 , \28701 , \28702 , \28703 , \28704 ,
         \28705 , \28706 , \28707 , \28708 , \28709 , \28710 , \28711 , \28712 , \28713 , \28714 ,
         \28715 , \28716 , \28717 , \28718 , \28719 , \28720 , \28721 , \28722 , \28723 , \28724 ,
         \28725 , \28726 , \28727 , \28728 , \28729 , \28730 , \28731 , \28732 , \28733 , \28734 ,
         \28735 , \28736 , \28737 , \28738 , \28739 , \28740 , \28741 , \28742 , \28743 , \28744 ,
         \28745 , \28746 , \28747 , \28748 , \28749 , \28750 , \28751 , \28752 , \28753 , \28754 ,
         \28755 , \28756 , \28757 , \28758 , \28759 , \28760 , \28761 , \28762 , \28763 , \28764 ,
         \28765 , \28766 , \28767 , \28768 , \28769 , \28770 , \28771 , \28772 , \28773 , \28774 ,
         \28775 , \28776 , \28777 , \28778 , \28779 , \28780 , \28781 , \28782 , \28783 , \28784 ,
         \28785 , \28786 , \28787 , \28788 , \28789 , \28790 , \28791 , \28792 , \28793 , \28794 ,
         \28795 , \28796 , \28797 , \28798 , \28799 , \28800 , \28801 , \28802 , \28803 , \28804 ,
         \28805 , \28806 , \28807 , \28808 , \28809 , \28810 , \28811 , \28812 , \28813 , \28814 ,
         \28815 , \28816 , \28817 , \28818 , \28819 , \28820 , \28821 , \28822 , \28823 , \28824 ,
         \28825 , \28826 , \28827 , \28828 , \28829 , \28830 , \28831 , \28832 , \28833 , \28834 ,
         \28835 , \28836 , \28837 , \28838 , \28839 , \28840 , \28841 , \28842 , \28843 , \28844 ,
         \28845 , \28846 , \28847 , \28848 , \28849 , \28850 , \28851 , \28852 , \28853 , \28854 ,
         \28855 , \28856 , \28857 , \28858 , \28859 , \28860 , \28861 , \28862 , \28863 , \28864 ,
         \28865 , \28866 , \28867 , \28868 , \28869 , \28870 , \28871 , \28872 , \28873 , \28874 ,
         \28875 , \28876 , \28877 , \28878 , \28879 , \28880 , \28881 , \28882 , \28883 , \28884 ,
         \28885 , \28886 , \28887 , \28888 , \28889 , \28890 , \28891 , \28892 , \28893 , \28894 ,
         \28895 , \28896 , \28897 , \28898 , \28899 , \28900 , \28901 , \28902 , \28903 , \28904 ,
         \28905 , \28906 , \28907 , \28908 , \28909 , \28910 , \28911 , \28912 , \28913 , \28914 ,
         \28915 , \28916 , \28917 , \28918 , \28919 , \28920 , \28921 , \28922 , \28923 , \28924 ,
         \28925 , \28926 , \28927 , \28928 , \28929 , \28930 , \28931 , \28932 , \28933 , \28934 ,
         \28935 , \28936 , \28937 , \28938 , \28939 , \28940 , \28941 , \28942 , \28943 , \28944 ,
         \28945 , \28946 , \28947 , \28948 , \28949 , \28950 , \28951 , \28952 , \28953 , \28954 ,
         \28955 , \28956 , \28957 , \28958 , \28959 , \28960 , \28961 , \28962 , \28963 , \28964 ,
         \28965 , \28966 , \28967 , \28968 , \28969 , \28970 , \28971 , \28972 , \28973 , \28974 ,
         \28975 , \28976 , \28977 , \28978 , \28979 , \28980 , \28981 , \28982 , \28983 , \28984 ,
         \28985 , \28986 , \28987 , \28988 , \28989 , \28990 , \28991 , \28992 , \28993 , \28994 ,
         \28995 , \28996 , \28997 , \28998 , \28999 , \29000 , \29001 , \29002 , \29003 , \29004 ,
         \29005 , \29006 , \29007 , \29008 , \29009 , \29010 , \29011 , \29012 , \29013 , \29014 ,
         \29015 , \29016 , \29017 , \29018 , \29019 , \29020 , \29021 , \29022 , \29023 , \29024 ,
         \29025 , \29026 , \29027 , \29028 , \29029 , \29030 , \29031 , \29032 , \29033 , \29034 ,
         \29035 , \29036 , \29037 , \29038 , \29039 , \29040 , \29041 , \29042 , \29043 , \29044 ,
         \29045 , \29046 , \29047 , \29048 , \29049 , \29050 , \29051 , \29052 , \29053 , \29054 ,
         \29055 , \29056 , \29057 , \29058 , \29059 , \29060 , \29061 , \29062 , \29063 , \29064 ,
         \29065 , \29066 , \29067 , \29068 , \29069 , \29070 , \29071 , \29072 , \29073 , \29074 ,
         \29075 , \29076 , \29077 , \29078 , \29079 , \29080 , \29081 , \29082 , \29083 , \29084 ,
         \29085 , \29086 , \29087 , \29088 , \29089 , \29090 , \29091 , \29092 , \29093 , \29094 ,
         \29095 , \29096 , \29097 , \29098 , \29099 , \29100 , \29101 , \29102 , \29103 , \29104 ,
         \29105 , \29106 , \29107 , \29108 , \29109 , \29110 , \29111 , \29112 , \29113 , \29114 ,
         \29115 , \29116 , \29117 , \29118 , \29119 , \29120 , \29121 , \29122 , \29123 , \29124 ,
         \29125 , \29126 , \29127 , \29128 , \29129 , \29130 , \29131 , \29132 , \29133 , \29134 ,
         \29135 , \29136 , \29137 , \29138 , \29139 , \29140 , \29141 , \29142 , \29143 , \29144 ,
         \29145 , \29146 , \29147 , \29148 , \29149 , \29150 , \29151 , \29152 , \29153 , \29154 ,
         \29155 , \29156 , \29157 , \29158 , \29159 , \29160 , \29161 , \29162 , \29163 , \29164 ,
         \29165 , \29166 , \29167 , \29168 , \29169 , \29170 , \29171 , \29172 , \29173 , \29174 ,
         \29175 , \29176 , \29177 , \29178 , \29179 , \29180 , \29181 , \29182 , \29183 , \29184 ,
         \29185 , \29186 , \29187 , \29188 , \29189 , \29190 , \29191 , \29192 , \29193 , \29194 ,
         \29195 , \29196 , \29197 , \29198 , \29199 , \29200 , \29201 , \29202 , \29203 , \29204 ,
         \29205 , \29206 , \29207 , \29208 , \29209 , \29210 , \29211 , \29212 , \29213 , \29214 ,
         \29215 , \29216 , \29217 , \29218 , \29219 , \29220 , \29221 , \29222 , \29223 , \29224 ,
         \29225 , \29226 , \29227 , \29228 , \29229 , \29230 , \29231 , \29232 , \29233 , \29234 ,
         \29235 , \29236 , \29237 , \29238 , \29239 , \29240 , \29241 , \29242 , \29243 , \29244 ,
         \29245 , \29246 , \29247 , \29248 , \29249 , \29250 , \29251 , \29252 , \29253 , \29254 ,
         \29255 , \29256 , \29257 , \29258 , \29259 , \29260 , \29261 , \29262 , \29263 , \29264 ,
         \29265 , \29266 , \29267 , \29268 , \29269 , \29270 , \29271 , \29272 , \29273 , \29274 ,
         \29275 , \29276 , \29277 , \29278 , \29279 , \29280 , \29281 , \29282 , \29283 , \29284 ,
         \29285 , \29286 , \29287 , \29288 , \29289 , \29290 , \29291 , \29292 , \29293 , \29294 ,
         \29295 , \29296 , \29297 , \29298 , \29299 , \29300 , \29301 , \29302 , \29303 , \29304 ,
         \29305 , \29306 , \29307 , \29308 , \29309 , \29310 , \29311 , \29312 , \29313 , \29314 ,
         \29315 , \29316 , \29317 , \29318 , \29319 , \29320 , \29321 , \29322 , \29323 , \29324 ,
         \29325 , \29326 , \29327 , \29328 , \29329 , \29330 , \29331 , \29332 , \29333 , \29334 ,
         \29335 , \29336 , \29337 , \29338 , \29339 , \29340 , \29341 , \29342 , \29343 , \29344 ,
         \29345 , \29346 , \29347 , \29348 , \29349 , \29350 , \29351 , \29352 , \29353 , \29354 ,
         \29355 , \29356 , \29357 , \29358 , \29359 , \29360 , \29361 , \29362 , \29363 , \29364 ,
         \29365 , \29366 , \29367 , \29368 , \29369 , \29370 , \29371 , \29372 , \29373 , \29374 ,
         \29375 , \29376 , \29377 , \29378 , \29379 , \29380 , \29381 , \29382 , \29383 , \29384 ,
         \29385 , \29386 , \29387 , \29388 , \29389 , \29390 , \29391 , \29392 , \29393 , \29394 ,
         \29395 , \29396 , \29397 , \29398 , \29399 , \29400 , \29401 , \29402 , \29403 , \29404 ,
         \29405 , \29406 , \29407 , \29408 , \29409 , \29410 , \29411 , \29412 , \29413 , \29414 ,
         \29415 , \29416 , \29417 , \29418 , \29419 , \29420 , \29421 , \29422 , \29423 , \29424 ,
         \29425 , \29426 , \29427 , \29428 , \29429 , \29430 , \29431 , \29432 , \29433 , \29434 ,
         \29435 , \29436 , \29437 , \29438 , \29439 , \29440 , \29441 , \29442 , \29443 , \29444 ,
         \29445 , \29446 , \29447 , \29448 , \29449 , \29450 , \29451 , \29452 , \29453 , \29454 ,
         \29455 , \29456 , \29457 , \29458 , \29459 , \29460 , \29461 , \29462 , \29463 , \29464 ,
         \29465 , \29466 , \29467 , \29468 , \29469 , \29470 , \29471 , \29472 , \29473 , \29474 ,
         \29475 , \29476 , \29477 , \29478 , \29479 , \29480 , \29481 , \29482 , \29483 , \29484 ,
         \29485 , \29486 , \29487 , \29488 , \29489 , \29490 , \29491 , \29492 , \29493 , \29494 ,
         \29495 , \29496 , \29497 , \29498 , \29499 , \29500 , \29501 , \29502 , \29503 , \29504 ,
         \29505 , \29506 , \29507 , \29508 , \29509 , \29510 , \29511 , \29512 , \29513 , \29514 ,
         \29515 , \29516 , \29517 , \29518 , \29519 , \29520 , \29521 , \29522 , \29523 , \29524 ,
         \29525 , \29526 , \29527 , \29528 , \29529 , \29530 , \29531 , \29532 , \29533 , \29534 ,
         \29535 , \29536 , \29537 , \29538 , \29539 , \29540 , \29541 , \29542 , \29543 , \29544 ,
         \29545 , \29546 , \29547 , \29548 , \29549 , \29550 , \29551 , \29552 , \29553 , \29554 ,
         \29555 , \29556 , \29557 , \29558 , \29559 , \29560 , \29561 , \29562 , \29563 , \29564 ,
         \29565 , \29566 , \29567 , \29568 , \29569 , \29570 , \29571 , \29572 , \29573 , \29574 ,
         \29575 , \29576 , \29577 , \29578 , \29579 , \29580 , \29581 , \29582 , \29583 , \29584 ,
         \29585 , \29586 , \29587 , \29588 , \29589 , \29590 , \29591 , \29592 , \29593 , \29594 ,
         \29595 , \29596 , \29597 , \29598 , \29599 , \29600 , \29601 , \29602 , \29603 , \29604 ,
         \29605 , \29606 , \29607 , \29608 , \29609 , \29610 , \29611 , \29612 , \29613 , \29614 ,
         \29615 , \29616 , \29617 , \29618 , \29619 , \29620 , \29621 , \29622 , \29623 , \29624 ,
         \29625 , \29626 , \29627 , \29628 , \29629 , \29630 , \29631 , \29632 , \29633 , \29634 ,
         \29635 , \29636 , \29637 , \29638 , \29639 , \29640 , \29641 , \29642 , \29643 , \29644 ,
         \29645 , \29646 , \29647 , \29648 , \29649 , \29650 , \29651 , \29652 , \29653 , \29654 ,
         \29655 , \29656 , \29657 , \29658 , \29659 , \29660 , \29661 , \29662 , \29663 , \29664 ,
         \29665 , \29666 , \29667 , \29668 , \29669 , \29670 , \29671 , \29672 , \29673 , \29674 ,
         \29675 , \29676 , \29677 , \29678 , \29679 , \29680 , \29681 , \29682 , \29683 , \29684 ,
         \29685 , \29686 , \29687 , \29688 , \29689 , \29690 , \29691 , \29692 , \29693 , \29694 ,
         \29695 , \29696 , \29697 , \29698 , \29699 , \29700 , \29701 , \29702 , \29703 , \29704 ,
         \29705 , \29706 , \29707 , \29708 , \29709 , \29710 , \29711 , \29712 , \29713 , \29714 ,
         \29715 , \29716 , \29717 , \29718 , \29719 , \29720 , \29721 , \29722 , \29723 , \29724 ,
         \29725 , \29726 , \29727 , \29728 , \29729 , \29730 , \29731 , \29732 , \29733 , \29734 ,
         \29735 , \29736 , \29737 , \29738 , \29739 , \29740 , \29741 , \29742 , \29743 , \29744 ,
         \29745 , \29746 , \29747 , \29748 , \29749 , \29750 , \29751 , \29752 , \29753 , \29754 ,
         \29755 , \29756 , \29757 , \29758 , \29759 , \29760 , \29761 , \29762 , \29763 , \29764 ,
         \29765 , \29766 , \29767 , \29768 , \29769 , \29770 , \29771 , \29772 , \29773 , \29774 ,
         \29775 , \29776 , \29777 , \29778 , \29779 , \29780 , \29781 , \29782 , \29783 , \29784 ,
         \29785 , \29786 , \29787 , \29788 , \29789 , \29790 , \29791 , \29792 , \29793 , \29794 ,
         \29795 , \29796 , \29797 , \29798 , \29799 , \29800 , \29801 , \29802 , \29803 , \29804 ,
         \29805 , \29806 , \29807 , \29808 , \29809 , \29810 , \29811 , \29812 , \29813 , \29814 ,
         \29815 , \29816 , \29817 , \29818 , \29819 , \29820 , \29821 , \29822 , \29823 , \29824 ,
         \29825 , \29826 , \29827 , \29828 , \29829 , \29830 , \29831 , \29832 , \29833 , \29834 ,
         \29835 , \29836 , \29837 , \29838 , \29839 , \29840 , \29841 , \29842 , \29843 , \29844 ,
         \29845 , \29846 , \29847 , \29848 , \29849 , \29850 , \29851 , \29852 , \29853 , \29854 ,
         \29855 , \29856 , \29857 , \29858 , \29859 , \29860 , \29861 , \29862 , \29863 , \29864 ,
         \29865 , \29866 , \29867 , \29868 , \29869 , \29870 , \29871 , \29872 , \29873 , \29874 ,
         \29875 , \29876 , \29877 , \29878 , \29879 , \29880 , \29881 , \29882 , \29883 , \29884 ,
         \29885 , \29886 , \29887 , \29888 , \29889 , \29890 , \29891 , \29892 , \29893 , \29894 ,
         \29895 , \29896 , \29897 , \29898 , \29899 , \29900 , \29901 , \29902 , \29903 , \29904 ,
         \29905 , \29906 , \29907 , \29908 , \29909 , \29910 , \29911 , \29912 , \29913 , \29914 ,
         \29915 , \29916 , \29917 , \29918 , \29919 , \29920 , \29921 , \29922 , \29923 , \29924 ,
         \29925 , \29926 , \29927 , \29928 , \29929 , \29930 , \29931 , \29932 , \29933 , \29934 ,
         \29935 , \29936 , \29937 , \29938 , \29939 , \29940 , \29941 , \29942 , \29943 , \29944 ,
         \29945 , \29946 , \29947 , \29948 , \29949 , \29950 , \29951 , \29952 , \29953 , \29954 ,
         \29955 , \29956 , \29957 , \29958 , \29959 , \29960 , \29961 , \29962 , \29963 , \29964 ,
         \29965 , \29966 , \29967 , \29968 , \29969 , \29970 , \29971 , \29972 , \29973 , \29974 ,
         \29975 , \29976 , \29977 , \29978 , \29979 , \29980 , \29981 , \29982 , \29983 , \29984 ,
         \29985 , \29986 , \29987 , \29988 , \29989 , \29990 , \29991 , \29992 , \29993 , \29994 ,
         \29995 , \29996 , \29997 , \29998 , \29999 , \30000 , \30001 , \30002 , \30003 , \30004 ,
         \30005 , \30006 , \30007 , \30008 , \30009 , \30010 , \30011 , \30012 , \30013 , \30014 ,
         \30015 , \30016 , \30017 , \30018 , \30019 , \30020 , \30021 , \30022 , \30023 , \30024 ,
         \30025 , \30026 , \30027 , \30028 , \30029 , \30030 , \30031 , \30032 , \30033 , \30034 ,
         \30035 , \30036 , \30037 , \30038 , \30039 , \30040 , \30041 , \30042 , \30043 , \30044 ,
         \30045 , \30046 , \30047 , \30048 , \30049 , \30050 , \30051 , \30052 , \30053 , \30054 ,
         \30055 , \30056 , \30057 , \30058 , \30059 , \30060 , \30061 , \30062 , \30063 , \30064 ,
         \30065 , \30066 , \30067 , \30068 , \30069 , \30070 , \30071 , \30072 , \30073 , \30074 ,
         \30075 , \30076 , \30077 , \30078 , \30079 , \30080 , \30081 , \30082 , \30083 , \30084 ,
         \30085 , \30086 , \30087 , \30088 , \30089 , \30090 , \30091 , \30092 , \30093 , \30094 ,
         \30095 , \30096 , \30097 , \30098 , \30099 , \30100 , \30101 , \30102 , \30103 , \30104 ,
         \30105 , \30106 , \30107 , \30108 , \30109 , \30110 , \30111 , \30112 , \30113 , \30114 ,
         \30115 , \30116 , \30117 , \30118 , \30119 , \30120 , \30121 , \30122 , \30123 , \30124 ,
         \30125 , \30126 , \30127 , \30128 , \30129 , \30130 , \30131 , \30132 , \30133 , \30134 ,
         \30135 , \30136 , \30137 , \30138 , \30139 , \30140 , \30141 , \30142 , \30143 , \30144 ,
         \30145 , \30146 , \30147 , \30148 , \30149 , \30150 , \30151 , \30152 , \30153 , \30154 ,
         \30155 , \30156 , \30157 , \30158 , \30159 , \30160 , \30161 , \30162 , \30163 , \30164 ,
         \30165 , \30166 , \30167 , \30168 , \30169 , \30170 , \30171 , \30172 , \30173 , \30174 ,
         \30175 , \30176 , \30177 , \30178 , \30179 , \30180 , \30181 , \30182 , \30183 , \30184 ,
         \30185 , \30186 , \30187 , \30188 , \30189 , \30190 , \30191 , \30192 , \30193 , \30194 ,
         \30195 , \30196 , \30197 , \30198 , \30199 , \30200 , \30201 , \30202 , \30203 , \30204 ,
         \30205 , \30206 , \30207 , \30208 , \30209 , \30210 , \30211 , \30212 , \30213 , \30214 ,
         \30215 , \30216 , \30217 , \30218 , \30219 , \30220 , \30221 , \30222 , \30223 , \30224 ,
         \30225 , \30226 , \30227 , \30228 , \30229 , \30230 , \30231 , \30232 , \30233 , \30234 ,
         \30235 , \30236 , \30237 , \30238 , \30239 , \30240 , \30241 , \30242 , \30243 , \30244 ,
         \30245 , \30246 , \30247 , \30248 , \30249 , \30250 , \30251 , \30252 , \30253 , \30254 ,
         \30255 , \30256 , \30257 , \30258 , \30259 , \30260 , \30261 , \30262 , \30263 , \30264 ,
         \30265 , \30266 , \30267 , \30268 , \30269 , \30270 , \30271 , \30272 , \30273 , \30274 ,
         \30275 , \30276 , \30277 , \30278 , \30279 , \30280 , \30281 , \30282 , \30283 , \30284 ,
         \30285 , \30286 , \30287 , \30288 , \30289 , \30290 , \30291 , \30292 , \30293 , \30294 ,
         \30295 , \30296 , \30297 , \30298 , \30299 , \30300 , \30301 , \30302 , \30303 , \30304 ,
         \30305 , \30306 , \30307 , \30308 , \30309 , \30310 , \30311 , \30312 , \30313 , \30314 ,
         \30315 , \30316 , \30317 , \30318 , \30319 , \30320 , \30321 , \30322 , \30323 , \30324 ,
         \30325 , \30326 , \30327 , \30328 , \30329 , \30330 , \30331 , \30332 , \30333 , \30334 ,
         \30335 , \30336 , \30337 , \30338 , \30339 , \30340 , \30341 , \30342 , \30343 , \30344 ,
         \30345 , \30346 , \30347 , \30348 , \30349 , \30350 , \30351 , \30352 , \30353 , \30354 ,
         \30355 , \30356 , \30357 , \30358 , \30359 , \30360 , \30361 , \30362 , \30363 , \30364 ,
         \30365 , \30366 , \30367 , \30368 , \30369 , \30370 , \30371 , \30372 , \30373 , \30374 ,
         \30375 , \30376 , \30377 , \30378 , \30379 , \30380 , \30381 , \30382 , \30383 , \30384 ,
         \30385 , \30386 , \30387 , \30388 , \30389 , \30390 , \30391 , \30392 , \30393 , \30394 ,
         \30395 , \30396 , \30397 , \30398 , \30399 , \30400 , \30401 , \30402 , \30403 , \30404 ,
         \30405 , \30406 , \30407 , \30408 , \30409 , \30410 , \30411 , \30412 , \30413 , \30414 ,
         \30415 , \30416 , \30417 , \30418 , \30419 , \30420 , \30421 , \30422 , \30423 , \30424 ,
         \30425 , \30426 , \30427 , \30428 , \30429 , \30430 , \30431 , \30432 , \30433 , \30434 ,
         \30435 , \30436 , \30437 , \30438 , \30439 , \30440 , \30441 , \30442 , \30443 , \30444 ,
         \30445 , \30446 , \30447 , \30448 , \30449 , \30450 , \30451 , \30452 , \30453 , \30454 ,
         \30455 , \30456 , \30457 , \30458 , \30459 , \30460 , \30461 , \30462 , \30463 , \30464 ,
         \30465 , \30466 , \30467 , \30468 , \30469 , \30470 , \30471 , \30472 , \30473 , \30474 ,
         \30475 , \30476 , \30477 , \30478 , \30479 , \30480 , \30481 , \30482 , \30483 , \30484 ,
         \30485 , \30486 , \30487 , \30488 , \30489 , \30490 , \30491 , \30492 , \30493 , \30494 ,
         \30495 , \30496 , \30497 , \30498 , \30499 , \30500 , \30501 , \30502 , \30503 , \30504 ,
         \30505 , \30506 , \30507 , \30508 , \30509 , \30510 , \30511 , \30512 , \30513 , \30514 ,
         \30515 , \30516 , \30517 , \30518 , \30519 , \30520 , \30521 , \30522 , \30523 , \30524 ,
         \30525 , \30526 , \30527 , \30528 , \30529 , \30530 , \30531 , \30532 , \30533 , \30534 ,
         \30535 , \30536 , \30537 , \30538 , \30539 , \30540 , \30541 , \30542 , \30543 , \30544 ,
         \30545 , \30546 , \30547 , \30548 , \30549 , \30550 , \30551 , \30552 , \30553 , \30554 ,
         \30555 , \30556 , \30557 , \30558 , \30559 , \30560 , \30561 , \30562 , \30563 , \30564 ,
         \30565 , \30566 , \30567 , \30568 , \30569 , \30570 , \30571 , \30572 , \30573 , \30574 ,
         \30575 , \30576 , \30577 , \30578 , \30579 , \30580 , \30581 , \30582 , \30583 , \30584 ,
         \30585 , \30586 , \30587 , \30588 , \30589 , \30590 , \30591 , \30592 , \30593 , \30594 ,
         \30595 , \30596 , \30597 , \30598 , \30599 , \30600 , \30601 , \30602 , \30603 , \30604 ,
         \30605 , \30606 , \30607 , \30608 , \30609 , \30610 , \30611 , \30612 , \30613 , \30614 ,
         \30615 , \30616 , \30617 , \30618 , \30619 , \30620 , \30621 , \30622 , \30623 , \30624 ,
         \30625 , \30626 , \30627 , \30628 , \30629 , \30630 , \30631 , \30632 , \30633 , \30634 ,
         \30635 , \30636 , \30637 , \30638 , \30639 , \30640 , \30641 , \30642 , \30643 , \30644 ,
         \30645 , \30646 , \30647 , \30648 , \30649 , \30650 , \30651 , \30652 , \30653 , \30654 ,
         \30655 , \30656 , \30657 , \30658 , \30659 , \30660 , \30661 , \30662 , \30663 , \30664 ,
         \30665 , \30666 , \30667 , \30668 , \30669 , \30670 , \30671 , \30672 , \30673 , \30674 ,
         \30675 , \30676 , \30677 , \30678 , \30679 , \30680 , \30681 , \30682 , \30683 , \30684 ,
         \30685 , \30686 , \30687 , \30688 , \30689 , \30690 , \30691 , \30692 , \30693 , \30694 ,
         \30695 , \30696 , \30697 , \30698 , \30699 , \30700 , \30701 , \30702 , \30703 , \30704 ,
         \30705 , \30706 , \30707 , \30708 , \30709 , \30710 , \30711 , \30712 , \30713 , \30714 ,
         \30715 , \30716 , \30717 , \30718 , \30719 , \30720 , \30721 , \30722 , \30723 , \30724 ,
         \30725 , \30726 , \30727 , \30728 , \30729 , \30730 , \30731 , \30732 , \30733 , \30734 ,
         \30735 , \30736 , \30737 , \30738 , \30739 , \30740 , \30741 , \30742 , \30743 , \30744 ,
         \30745 , \30746 , \30747 , \30748 , \30749 , \30750 , \30751 , \30752 , \30753 , \30754 ,
         \30755 , \30756 , \30757 , \30758 , \30759 , \30760 , \30761 , \30762 , \30763 , \30764 ,
         \30765 , \30766 , \30767 , \30768 , \30769 , \30770 , \30771 , \30772 , \30773 , \30774 ,
         \30775 , \30776 , \30777 , \30778 , \30779 , \30780 , \30781 , \30782 , \30783 , \30784 ,
         \30785 , \30786 , \30787 , \30788 , \30789 , \30790 , \30791 , \30792 , \30793 , \30794 ,
         \30795 , \30796 , \30797 , \30798 , \30799 , \30800 , \30801 , \30802 , \30803 , \30804 ,
         \30805 , \30806 , \30807 , \30808 , \30809 , \30810 , \30811 , \30812 , \30813 , \30814 ,
         \30815 , \30816 , \30817 , \30818 , \30819 , \30820 , \30821 , \30822 , \30823 , \30824 ,
         \30825 , \30826 , \30827 , \30828 , \30829 , \30830 , \30831 , \30832 , \30833 , \30834 ,
         \30835 , \30836 , \30837 , \30838 , \30839 , \30840 , \30841 , \30842 , \30843 , \30844 ,
         \30845 , \30846 , \30847 , \30848 , \30849 , \30850 , \30851 , \30852 , \30853 , \30854 ,
         \30855 , \30856 , \30857 , \30858 , \30859 , \30860 , \30861 , \30862 , \30863 , \30864 ,
         \30865 , \30866 , \30867 , \30868 , \30869 , \30870 , \30871 , \30872 , \30873 , \30874 ,
         \30875 , \30876 , \30877 , \30878 , \30879 , \30880 , \30881 , \30882 , \30883 , \30884 ,
         \30885 , \30886 , \30887 , \30888 , \30889 , \30890 , \30891 , \30892 , \30893 , \30894 ,
         \30895 , \30896 , \30897 , \30898 , \30899 , \30900 , \30901 , \30902 , \30903 , \30904 ,
         \30905 , \30906 , \30907 , \30908 , \30909 , \30910 , \30911 , \30912 , \30913 , \30914 ,
         \30915 , \30916 , \30917 , \30918 , \30919 , \30920 , \30921 , \30922 , \30923 , \30924 ,
         \30925 , \30926 , \30927 , \30928 , \30929 , \30930 , \30931 , \30932 , \30933 , \30934 ,
         \30935 , \30936 , \30937 , \30938 , \30939 , \30940 , \30941 , \30942 , \30943 , \30944 ,
         \30945 , \30946 , \30947 , \30948 , \30949 , \30950 , \30951 , \30952 , \30953 , \30954 ,
         \30955 , \30956 , \30957 , \30958 , \30959 , \30960 , \30961 , \30962 , \30963 , \30964 ,
         \30965 , \30966 , \30967 , \30968 , \30969 , \30970 , \30971 , \30972 , \30973 , \30974 ,
         \30975 , \30976 , \30977 , \30978 , \30979 , \30980 , \30981 , \30982 , \30983 , \30984 ,
         \30985 , \30986 , \30987 , \30988 , \30989 , \30990 , \30991 , \30992 , \30993 , \30994 ,
         \30995 , \30996 , \30997 , \30998 , \30999 , \31000 , \31001 , \31002 , \31003 , \31004 ,
         \31005 , \31006 , \31007 , \31008 , \31009 , \31010 , \31011 , \31012 , \31013 , \31014 ,
         \31015 , \31016 , \31017 , \31018 , \31019 , \31020 , \31021 , \31022 , \31023 , \31024 ,
         \31025 , \31026 , \31027 , \31028 , \31029 , \31030 , \31031 , \31032 , \31033 , \31034 ,
         \31035 , \31036 , \31037 , \31038 , \31039 , \31040 , \31041 , \31042 , \31043 , \31044 ,
         \31045 , \31046 , \31047 , \31048 , \31049 , \31050 , \31051 , \31052 , \31053 , \31054 ,
         \31055 , \31056 , \31057 , \31058 , \31059 , \31060 , \31061 , \31062 , \31063 , \31064 ,
         \31065 , \31066 , \31067 , \31068 , \31069 , \31070 , \31071 , \31072 , \31073 , \31074 ,
         \31075 , \31076 , \31077 , \31078 , \31079 , \31080 , \31081 , \31082 , \31083 , \31084 ,
         \31085 , \31086 , \31087 , \31088 , \31089 , \31090 , \31091 , \31092 , \31093 , \31094 ,
         \31095 , \31096 , \31097 , \31098 , \31099 , \31100 , \31101 , \31102 , \31103 , \31104 ,
         \31105 , \31106 , \31107 , \31108 , \31109 , \31110 , \31111 , \31112 , \31113 , \31114 ,
         \31115 , \31116 , \31117 , \31118 , \31119 , \31120 , \31121 , \31122 , \31123 , \31124 ,
         \31125 , \31126 , \31127 , \31128 , \31129 , \31130 , \31131 , \31132 , \31133 , \31134 ,
         \31135 , \31136 , \31137 , \31138 , \31139 , \31140 , \31141 , \31142 , \31143 , \31144 ,
         \31145 , \31146 , \31147 , \31148 , \31149 , \31150 , \31151 , \31152 , \31153 , \31154 ,
         \31155 , \31156 , \31157 , \31158 , \31159 , \31160 , \31161 , \31162 , \31163 , \31164 ,
         \31165 , \31166 , \31167 , \31168 , \31169 , \31170 , \31171 , \31172 , \31173 , \31174 ,
         \31175 , \31176 , \31177 , \31178 , \31179 , \31180 , \31181 , \31182 , \31183 , \31184 ,
         \31185 , \31186 , \31187 , \31188 , \31189 , \31190 , \31191 , \31192 , \31193 , \31194 ,
         \31195 , \31196 , \31197 , \31198 , \31199 , \31200 , \31201 , \31202 , \31203 , \31204 ,
         \31205 , \31206 , \31207 , \31208 , \31209 , \31210 , \31211 , \31212 , \31213 , \31214 ,
         \31215 , \31216 , \31217 , \31218 , \31219 , \31220 , \31221 , \31222 , \31223 , \31224 ,
         \31225 , \31226 , \31227 , \31228 , \31229 , \31230 , \31231 , \31232 , \31233 , \31234 ,
         \31235 , \31236 , \31237 , \31238 , \31239 , \31240 , \31241 , \31242 , \31243 , \31244 ,
         \31245 , \31246 , \31247 , \31248 , \31249 , \31250 , \31251 , \31252 , \31253 , \31254 ,
         \31255 , \31256 , \31257 , \31258 , \31259 , \31260 , \31261 , \31262 , \31263 , \31264 ,
         \31265 , \31266 , \31267 , \31268 , \31269 , \31270 , \31271 , \31272 , \31273 , \31274 ,
         \31275 , \31276 , \31277 , \31278 , \31279 , \31280 , \31281 , \31282 , \31283 , \31284 ,
         \31285 , \31286 , \31287 , \31288 , \31289 , \31290 , \31291 , \31292 , \31293 , \31294 ,
         \31295 , \31296 , \31297 , \31298 , \31299 , \31300 , \31301 , \31302 , \31303 , \31304 ,
         \31305 , \31306 , \31307 , \31308 , \31309 , \31310 , \31311 , \31312 , \31313 , \31314 ,
         \31315 , \31316 , \31317 , \31318 , \31319 , \31320 , \31321 , \31322 , \31323 , \31324 ,
         \31325 , \31326 , \31327 , \31328 , \31329 , \31330 , \31331 , \31332 , \31333 , \31334 ,
         \31335 , \31336 , \31337 , \31338 , \31339 , \31340 , \31341 , \31342 , \31343 , \31344 ,
         \31345 , \31346 , \31347 , \31348 , \31349 , \31350 , \31351 , \31352 , \31353 , \31354 ,
         \31355 , \31356 , \31357 , \31358 , \31359 , \31360 , \31361 , \31362 , \31363 , \31364 ,
         \31365 , \31366 , \31367 , \31368 , \31369 , \31370 , \31371 , \31372 , \31373 , \31374 ,
         \31375 , \31376 , \31377 , \31378 , \31379 , \31380 , \31381 , \31382 , \31383 , \31384 ,
         \31385 , \31386 , \31387 , \31388 , \31389 , \31390 , \31391 , \31392 , \31393 , \31394 ,
         \31395 , \31396 , \31397 , \31398 , \31399 , \31400 , \31401 , \31402 , \31403 , \31404 ,
         \31405 , \31406 , \31407 , \31408 , \31409 , \31410 , \31411 , \31412 , \31413 , \31414 ,
         \31415 , \31416 , \31417 , \31418 , \31419 , \31420 , \31421 , \31422 , \31423 , \31424 ,
         \31425 , \31426 , \31427 , \31428 , \31429 , \31430 , \31431 , \31432 , \31433 , \31434 ,
         \31435 , \31436 , \31437 , \31438 , \31439 , \31440 , \31441 , \31442 , \31443 , \31444 ,
         \31445 , \31446 , \31447 , \31448 , \31449 , \31450 , \31451 , \31452 , \31453 , \31454 ,
         \31455 , \31456 , \31457 , \31458 , \31459 , \31460 , \31461 , \31462 , \31463 , \31464 ,
         \31465 , \31466 , \31467 , \31468 , \31469 , \31470 , \31471 , \31472 , \31473 , \31474 ,
         \31475 , \31476 , \31477 , \31478 , \31479 , \31480 , \31481 , \31482 , \31483 , \31484 ,
         \31485 , \31486 , \31487 , \31488 , \31489 , \31490 , \31491 , \31492 , \31493 , \31494 ,
         \31495 , \31496 , \31497 , \31498 , \31499 , \31500 , \31501 , \31502 , \31503 , \31504 ,
         \31505 , \31506 , \31507 , \31508 , \31509 , \31510 , \31511 , \31512 , \31513 , \31514 ,
         \31515 , \31516 , \31517 , \31518 , \31519 , \31520 , \31521 , \31522 , \31523 , \31524 ,
         \31525 , \31526 , \31527 , \31528 , \31529 , \31530 , \31531 , \31532 , \31533 , \31534 ,
         \31535 , \31536 , \31537 , \31538 , \31539 , \31540 , \31541 , \31542 , \31543 , \31544 ,
         \31545 , \31546 , \31547 , \31548 , \31549 , \31550 , \31551 , \31552 , \31553 , \31554 ,
         \31555 , \31556 , \31557 , \31558 , \31559 , \31560 , \31561 , \31562 , \31563 , \31564 ,
         \31565 , \31566 , \31567 , \31568 , \31569 , \31570 , \31571 , \31572 , \31573 , \31574 ,
         \31575 , \31576 , \31577 , \31578 , \31579 , \31580 , \31581 , \31582 , \31583 , \31584 ,
         \31585 , \31586 , \31587 , \31588 , \31589 , \31590 , \31591 , \31592 , \31593 , \31594 ,
         \31595 , \31596 , \31597 , \31598 , \31599 , \31600 , \31601 , \31602 , \31603 , \31604 ,
         \31605 , \31606 , \31607 , \31608 , \31609 , \31610 , \31611 , \31612 , \31613 , \31614 ,
         \31615 , \31616 , \31617 , \31618 , \31619 , \31620 , \31621 , \31622 , \31623 , \31624 ,
         \31625 , \31626 , \31627 , \31628 , \31629 , \31630 , \31631 , \31632 , \31633 , \31634 ,
         \31635 , \31636 , \31637 , \31638 , \31639 , \31640 , \31641 , \31642 , \31643 , \31644 ,
         \31645 , \31646 , \31647 , \31648 , \31649 , \31650 , \31651 , \31652 , \31653 , \31654 ,
         \31655 , \31656 , \31657 , \31658 , \31659 , \31660 , \31661 , \31662 , \31663 , \31664 ,
         \31665 , \31666 , \31667 , \31668 , \31669 , \31670 , \31671 , \31672 , \31673 , \31674 ,
         \31675 , \31676 , \31677 , \31678 , \31679 , \31680 , \31681 , \31682 , \31683 , \31684 ,
         \31685 , \31686 , \31687 , \31688 , \31689 , \31690 , \31691 , \31692 , \31693 , \31694 ,
         \31695 , \31696 , \31697 , \31698 , \31699 , \31700 , \31701 , \31702 , \31703 , \31704 ,
         \31705 , \31706 , \31707 , \31708 , \31709 , \31710 , \31711 , \31712 , \31713 , \31714 ,
         \31715 , \31716 , \31717 , \31718 , \31719 , \31720 , \31721 , \31722 , \31723 , \31724 ,
         \31725 , \31726 , \31727 , \31728 , \31729 , \31730 , \31731 , \31732 , \31733 , \31734 ,
         \31735 , \31736 , \31737 , \31738 , \31739 , \31740 , \31741 , \31742 , \31743 , \31744 ,
         \31745 , \31746 , \31747 , \31748 , \31749 , \31750 , \31751 , \31752 , \31753 , \31754 ,
         \31755 , \31756 , \31757 , \31758 , \31759 , \31760 , \31761 , \31762 , \31763 , \31764 ,
         \31765 , \31766 , \31767 , \31768 , \31769 , \31770 , \31771 , \31772 , \31773 , \31774 ,
         \31775 , \31776 , \31777 , \31778 , \31779 , \31780 , \31781 , \31782 , \31783 , \31784 ,
         \31785 , \31786 , \31787 , \31788 , \31789 , \31790 , \31791 , \31792 , \31793 , \31794 ,
         \31795 , \31796 , \31797 , \31798 , \31799 , \31800 , \31801 , \31802 , \31803 , \31804 ,
         \31805 , \31806 , \31807 , \31808 , \31809 , \31810 , \31811 , \31812 , \31813 , \31814 ,
         \31815 , \31816 , \31817 , \31818 , \31819 , \31820 , \31821 , \31822 , \31823 , \31824 ,
         \31825 , \31826 , \31827 , \31828 , \31829 , \31830 , \31831 , \31832 , \31833 , \31834 ,
         \31835 , \31836 , \31837 , \31838 , \31839 , \31840 , \31841 , \31842 , \31843 , \31844 ,
         \31845 , \31846 , \31847 , \31848 , \31849 , \31850 , \31851 , \31852 , \31853 , \31854 ,
         \31855 , \31856 , \31857 , \31858 , \31859 , \31860 , \31861 , \31862 , \31863 , \31864 ,
         \31865 , \31866 , \31867 , \31868 , \31869 , \31870 , \31871 , \31872 , \31873 , \31874 ,
         \31875 , \31876 , \31877 , \31878 , \31879 , \31880 , \31881 , \31882 , \31883 , \31884 ,
         \31885 , \31886 , \31887 , \31888 , \31889 , \31890 , \31891 , \31892 , \31893 , \31894 ,
         \31895 , \31896 , \31897 , \31898 , \31899 , \31900 , \31901 , \31902 , \31903 , \31904 ,
         \31905 , \31906 , \31907 , \31908 , \31909 , \31910 , \31911 , \31912 , \31913 , \31914 ,
         \31915 , \31916 , \31917 , \31918 , \31919 , \31920 , \31921 , \31922 , \31923 , \31924 ,
         \31925 , \31926 , \31927 , \31928 , \31929 , \31930 , \31931 , \31932 , \31933 , \31934 ,
         \31935 , \31936 , \31937 , \31938 , \31939 , \31940 , \31941 , \31942 , \31943 , \31944 ,
         \31945 , \31946 , \31947 , \31948 , \31949 , \31950 , \31951 , \31952 , \31953 , \31954 ,
         \31955 , \31956 , \31957 , \31958 , \31959 , \31960 , \31961 , \31962 , \31963 , \31964 ,
         \31965 , \31966 , \31967 , \31968 , \31969 , \31970 , \31971 , \31972 , \31973 , \31974 ,
         \31975 , \31976 , \31977 , \31978 , \31979 , \31980 , \31981 , \31982 , \31983 , \31984 ,
         \31985 , \31986 , \31987 , \31988 , \31989 , \31990 , \31991 , \31992 , \31993 , \31994 ,
         \31995 , \31996 , \31997 , \31998 , \31999 , \32000 , \32001 , \32002 , \32003 , \32004 ,
         \32005 , \32006 , \32007 , \32008 , \32009 , \32010 , \32011 , \32012 , \32013 , \32014 ,
         \32015 , \32016 , \32017 , \32018 , \32019 , \32020 , \32021 , \32022 , \32023 , \32024 ,
         \32025 , \32026 , \32027 , \32028 , \32029 , \32030 , \32031 , \32032 , \32033 , \32034 ,
         \32035 , \32036 , \32037 , \32038 , \32039 , \32040 , \32041 , \32042 , \32043 , \32044 ,
         \32045 , \32046 , \32047 , \32048 , \32049 , \32050 , \32051 , \32052 , \32053 , \32054 ,
         \32055 , \32056 , \32057 , \32058 , \32059 , \32060 , \32061 , \32062 , \32063 , \32064 ,
         \32065 , \32066 , \32067 , \32068 , \32069 , \32070 , \32071 , \32072 , \32073 , \32074 ,
         \32075 , \32076 , \32077 , \32078 , \32079 , \32080 , \32081 , \32082 , \32083 , \32084 ,
         \32085 , \32086 , \32087 , \32088 , \32089 , \32090 , \32091 , \32092 , \32093 , \32094 ,
         \32095 , \32096 , \32097 , \32098 , \32099 , \32100 , \32101 , \32102 , \32103 , \32104 ,
         \32105 , \32106 , \32107 , \32108 , \32109 , \32110 , \32111 , \32112 , \32113 , \32114 ,
         \32115 , \32116 , \32117 , \32118 , \32119 , \32120 , \32121 , \32122 , \32123 , \32124 ,
         \32125 , \32126 , \32127 , \32128 , \32129 , \32130 , \32131 , \32132 , \32133 , \32134 ,
         \32135 , \32136 , \32137 , \32138 , \32139 , \32140 , \32141 , \32142 , \32143 , \32144 ,
         \32145 , \32146 , \32147 , \32148 , \32149 , \32150 , \32151 , \32152 , \32153 , \32154 ,
         \32155 , \32156 , \32157 , \32158 , \32159 , \32160 , \32161 , \32162 , \32163 , \32164 ,
         \32165 , \32166 , \32167 , \32168 , \32169 , \32170 , \32171 , \32172 , \32173 , \32174 ,
         \32175 , \32176 , \32177 , \32178 , \32179 , \32180 , \32181 , \32182 , \32183 , \32184 ,
         \32185 , \32186 , \32187 , \32188 , \32189 , \32190 , \32191 , \32192 , \32193 , \32194 ,
         \32195 , \32196 , \32197 , \32198 , \32199 , \32200 , \32201 , \32202 , \32203 , \32204 ,
         \32205 , \32206 , \32207 , \32208 , \32209 , \32210 , \32211 , \32212 , \32213 , \32214 ,
         \32215 , \32216 , \32217 , \32218 , \32219 , \32220 , \32221 , \32222 , \32223 , \32224 ,
         \32225 , \32226 , \32227 , \32228 , \32229 , \32230 , \32231 , \32232 , \32233 , \32234 ,
         \32235 , \32236 , \32237 , \32238 , \32239 , \32240 , \32241 , \32242 , \32243 , \32244 ,
         \32245 , \32246 , \32247 , \32248 , \32249 , \32250 , \32251 , \32252 , \32253 , \32254 ,
         \32255 , \32256 , \32257 , \32258 , \32259 , \32260 , \32261 , \32262 , \32263 , \32264 ,
         \32265 , \32266 , \32267 , \32268 , \32269 , \32270 , \32271 , \32272 , \32273 , \32274 ,
         \32275 , \32276 , \32277 , \32278 , \32279 , \32280 , \32281 , \32282 , \32283 , \32284 ,
         \32285 , \32286 , \32287 , \32288 , \32289 , \32290 , \32291 , \32292 , \32293 , \32294 ,
         \32295 , \32296 , \32297 , \32298 , \32299 , \32300 , \32301 , \32302 , \32303 , \32304 ,
         \32305 , \32306 , \32307 , \32308 , \32309 , \32310 , \32311 , \32312 , \32313 , \32314 ,
         \32315 , \32316 , \32317 , \32318 , \32319 , \32320 , \32321 , \32322 , \32323 , \32324 ,
         \32325 , \32326 , \32327 , \32328 , \32329 , \32330 , \32331 , \32332 , \32333 , \32334 ,
         \32335 , \32336 , \32337 , \32338 , \32339 , \32340 , \32341 , \32342 , \32343 , \32344 ,
         \32345 , \32346 , \32347 , \32348 , \32349 , \32350 , \32351 , \32352 , \32353 , \32354 ,
         \32355 , \32356 , \32357 , \32358 , \32359 , \32360 , \32361 , \32362 , \32363 , \32364 ,
         \32365 , \32366 , \32367 , \32368 , \32369 , \32370 , \32371 , \32372 , \32373 , \32374 ,
         \32375 , \32376 , \32377 , \32378 , \32379 , \32380 , \32381 , \32382 , \32383 , \32384 ,
         \32385 , \32386 , \32387 , \32388 , \32389 , \32390 , \32391 , \32392 , \32393 , \32394 ,
         \32395 , \32396 , \32397 , \32398 , \32399 , \32400 , \32401 , \32402 , \32403 , \32404 ,
         \32405 , \32406 , \32407 , \32408 , \32409 , \32410 , \32411 , \32412 , \32413 , \32414 ,
         \32415 , \32416 , \32417 , \32418 , \32419 , \32420 , \32421 , \32422 , \32423 , \32424 ,
         \32425 , \32426 , \32427 , \32428 , \32429 , \32430 , \32431 , \32432 , \32433 , \32434 ,
         \32435 , \32436 , \32437 , \32438 , \32439 , \32440 , \32441 , \32442 , \32443 , \32444 ,
         \32445 , \32446 , \32447 , \32448 , \32449 , \32450 , \32451 , \32452 , \32453 , \32454 ,
         \32455 , \32456 , \32457 , \32458 , \32459 , \32460 , \32461 , \32462 , \32463 , \32464 ,
         \32465 , \32466 , \32467 , \32468 , \32469 , \32470 , \32471 , \32472 , \32473 , \32474 ,
         \32475 , \32476 , \32477 , \32478 , \32479 , \32480 , \32481 , \32482 , \32483 , \32484 ,
         \32485 , \32486 , \32487 , \32488 , \32489 , \32490 , \32491 , \32492 , \32493 , \32494 ,
         \32495 , \32496 , \32497 , \32498 , \32499 , \32500 , \32501 , \32502 , \32503 , \32504 ,
         \32505 , \32506 , \32507 , \32508 , \32509 , \32510 , \32511 , \32512 , \32513 , \32514 ,
         \32515 , \32516 , \32517 , \32518 , \32519 , \32520 , \32521 , \32522 , \32523 , \32524 ,
         \32525 , \32526 , \32527 , \32528 , \32529 , \32530 , \32531 , \32532 , \32533 , \32534 ,
         \32535 , \32536 , \32537 , \32538 , \32539 , \32540 , \32541 , \32542 , \32543 , \32544 ,
         \32545 , \32546 , \32547 , \32548 , \32549 , \32550 , \32551 , \32552 , \32553 , \32554 ,
         \32555 , \32556 , \32557 , \32558 , \32559 , \32560 , \32561 , \32562 , \32563 , \32564 ,
         \32565 , \32566 , \32567 , \32568 , \32569 , \32570 , \32571 , \32572 , \32573 , \32574 ,
         \32575 , \32576 , \32577 , \32578 , \32579 , \32580 , \32581 , \32582 , \32583 , \32584 ,
         \32585 , \32586 , \32587 , \32588 , \32589 , \32590 , \32591 , \32592 , \32593 , \32594 ,
         \32595 , \32596 , \32597 , \32598 , \32599 , \32600 , \32601 , \32602 , \32603 , \32604 ,
         \32605 , \32606 , \32607 , \32608 , \32609 , \32610 , \32611 , \32612 , \32613 , \32614 ,
         \32615 , \32616 , \32617 , \32618 , \32619 , \32620 , \32621 , \32622 , \32623 , \32624 ,
         \32625 , \32626 , \32627 , \32628 , \32629 , \32630 , \32631 , \32632 , \32633 , \32634 ,
         \32635 , \32636 , \32637 , \32638 , \32639 , \32640 , \32641 , \32642 , \32643 , \32644 ,
         \32645 , \32646 , \32647 , \32648 , \32649 , \32650 , \32651 , \32652 , \32653 , \32654 ,
         \32655 , \32656 , \32657 , \32658 , \32659 , \32660 , \32661 , \32662 , \32663 , \32664 ,
         \32665 , \32666 , \32667 , \32668 , \32669 , \32670 , \32671 , \32672 , \32673 , \32674 ,
         \32675 , \32676 , \32677 , \32678 , \32679 , \32680 , \32681 , \32682 , \32683 , \32684 ,
         \32685 , \32686 , \32687 , \32688 , \32689 , \32690 , \32691 , \32692 , \32693 , \32694 ,
         \32695 , \32696 , \32697 , \32698 , \32699 , \32700 , \32701 , \32702 , \32703 , \32704 ,
         \32705 , \32706 , \32707 , \32708 , \32709 , \32710 , \32711 , \32712 , \32713 , \32714 ,
         \32715 , \32716 , \32717 , \32718 , \32719 , \32720 , \32721 , \32722 , \32723 , \32724 ,
         \32725 , \32726 , \32727 , \32728 , \32729 , \32730 , \32731 , \32732 , \32733 , \32734 ,
         \32735 , \32736 , \32737 , \32738 , \32739 , \32740 , \32741 , \32742 , \32743 , \32744 ,
         \32745 , \32746 , \32747 , \32748 , \32749 , \32750 , \32751 , \32752 , \32753 , \32754 ,
         \32755 , \32756 , \32757 , \32758 , \32759 , \32760 , \32761 , \32762 , \32763 , \32764 ,
         \32765 , \32766 , \32767 , \32768 , \32769 , \32770 , \32771 , \32772 , \32773 , \32774 ,
         \32775 , \32776 , \32777 , \32778 , \32779 , \32780 , \32781 , \32782 , \32783 , \32784 ,
         \32785 , \32786 , \32787 , \32788 , \32789 , \32790 , \32791 , \32792 , \32793 , \32794 ,
         \32795 , \32796 , \32797 , \32798 , \32799 , \32800 , \32801 , \32802 , \32803 , \32804 ,
         \32805 , \32806 , \32807 , \32808 , \32809 , \32810 , \32811 , \32812 , \32813 , \32814 ,
         \32815 , \32816 , \32817 , \32818 , \32819 , \32820 , \32821 , \32822 , \32823 , \32824 ,
         \32825 , \32826 , \32827 , \32828 , \32829 , \32830 , \32831 , \32832 , \32833 , \32834 ,
         \32835 , \32836 , \32837 , \32838 , \32839 , \32840 , \32841 , \32842 , \32843 , \32844 ,
         \32845 , \32846 , \32847 , \32848 , \32849 , \32850 , \32851 , \32852 , \32853 , \32854 ,
         \32855 , \32856 , \32857 , \32858 , \32859 , \32860 , \32861 , \32862 , \32863 , \32864 ,
         \32865 , \32866 , \32867 , \32868 , \32869 , \32870 , \32871 , \32872 , \32873 , \32874 ,
         \32875 , \32876 , \32877 , \32878 , \32879 , \32880 , \32881 , \32882 , \32883 , \32884 ,
         \32885 , \32886 , \32887 , \32888 , \32889 , \32890 , \32891 , \32892 , \32893 , \32894 ,
         \32895 , \32896 , \32897 , \32898 , \32899 , \32900 , \32901 , \32902 , \32903 , \32904 ,
         \32905 , \32906 , \32907 , \32908 , \32909 , \32910 , \32911 , \32912 , \32913 , \32914 ,
         \32915 , \32916 , \32917 , \32918 , \32919 , \32920 , \32921 , \32922 , \32923 , \32924 ,
         \32925 , \32926 , \32927 , \32928 , \32929 , \32930 , \32931 , \32932 , \32933 , \32934 ,
         \32935 , \32936 , \32937 , \32938 , \32939 , \32940 , \32941 , \32942 , \32943 , \32944 ,
         \32945 , \32946 , \32947 , \32948 , \32949 , \32950 , \32951 , \32952 , \32953 , \32954 ,
         \32955 , \32956 , \32957 , \32958 , \32959 , \32960 , \32961 , \32962 , \32963 , \32964 ,
         \32965 , \32966 , \32967 , \32968 , \32969 , \32970 , \32971 , \32972 , \32973 , \32974 ,
         \32975 , \32976 , \32977 , \32978 , \32979 , \32980 , \32981 , \32982 , \32983 , \32984 ,
         \32985 , \32986 , \32987 , \32988 , \32989 , \32990 , \32991 , \32992 , \32993 , \32994 ,
         \32995 , \32996 , \32997 , \32998 , \32999 , \33000 , \33001 , \33002 , \33003 , \33004 ,
         \33005 , \33006 , \33007 , \33008 , \33009 , \33010 , \33011 , \33012 , \33013 , \33014 ,
         \33015 , \33016 , \33017 , \33018 , \33019 , \33020 , \33021 , \33022 , \33023 , \33024 ,
         \33025 , \33026 , \33027 , \33028 , \33029 , \33030 , \33031 , \33032 , \33033 , \33034 ,
         \33035 , \33036 , \33037 , \33038 , \33039 , \33040 , \33041 , \33042 , \33043 , \33044 ,
         \33045 , \33046 , \33047 , \33048 , \33049 , \33050 , \33051 , \33052 , \33053 , \33054 ,
         \33055 , \33056 , \33057 , \33058 , \33059 , \33060 , \33061 , \33062 , \33063 , \33064 ,
         \33065 , \33066 , \33067 , \33068 , \33069 , \33070 , \33071 , \33072 , \33073 , \33074 ,
         \33075 , \33076 , \33077 , \33078 , \33079 , \33080 , \33081 , \33082 , \33083 , \33084 ,
         \33085 , \33086 , \33087 , \33088 , \33089 , \33090 , \33091 , \33092 , \33093 , \33094 ,
         \33095 , \33096 , \33097 , \33098 , \33099 , \33100 , \33101 , \33102 , \33103 , \33104 ,
         \33105 , \33106 , \33107 , \33108 , \33109 , \33110 , \33111 , \33112 , \33113 , \33114 ,
         \33115 , \33116 , \33117 , \33118 , \33119 , \33120 , \33121 , \33122 , \33123 , \33124 ,
         \33125 , \33126 , \33127 , \33128 , \33129 , \33130 , \33131 , \33132 , \33133 , \33134 ,
         \33135 , \33136 , \33137 , \33138 , \33139 , \33140 , \33141 , \33142 , \33143 , \33144 ,
         \33145 , \33146 , \33147 , \33148 , \33149 , \33150 , \33151 , \33152 , \33153 , \33154 ,
         \33155 , \33156 , \33157 , \33158 , \33159 , \33160 , \33161 , \33162 , \33163 , \33164 ,
         \33165 , \33166 , \33167 , \33168 , \33169 , \33170 , \33171 , \33172 , \33173 , \33174 ,
         \33175 , \33176 , \33177 , \33178 , \33179 , \33180 , \33181 , \33182 , \33183 , \33184 ,
         \33185 , \33186 , \33187 , \33188 , \33189 , \33190 , \33191 , \33192 , \33193 , \33194 ,
         \33195 , \33196 , \33197 , \33198 , \33199 , \33200 , \33201 , \33202 , \33203 , \33204 ,
         \33205 , \33206 , \33207 , \33208 , \33209 , \33210 , \33211 , \33212 , \33213 , \33214 ,
         \33215 , \33216 , \33217 , \33218 , \33219 , \33220 , \33221 , \33222 , \33223 , \33224 ,
         \33225 , \33226 , \33227 , \33228 , \33229 , \33230 , \33231 , \33232 , \33233 , \33234 ,
         \33235 , \33236 , \33237 , \33238 , \33239 , \33240 , \33241 , \33242 , \33243 , \33244 ,
         \33245 , \33246 , \33247 , \33248 , \33249 , \33250 , \33251 , \33252 , \33253 , \33254 ,
         \33255 , \33256 , \33257 , \33258 , \33259 , \33260 , \33261 , \33262 , \33263 , \33264 ,
         \33265 , \33266 , \33267 , \33268 , \33269 , \33270 , \33271 , \33272 , \33273 , \33274 ,
         \33275 , \33276 , \33277 , \33278 , \33279 , \33280 , \33281 , \33282 , \33283 , \33284 ,
         \33285 , \33286 , \33287 , \33288 , \33289 , \33290 , \33291 , \33292 , \33293 , \33294 ,
         \33295 , \33296 , \33297 , \33298 , \33299 , \33300 , \33301 , \33302 , \33303 , \33304 ,
         \33305 , \33306 , \33307 , \33308 , \33309 , \33310 , \33311 , \33312 , \33313 , \33314 ,
         \33315 , \33316 , \33317 , \33318 , \33319 , \33320 , \33321 , \33322 , \33323 , \33324 ,
         \33325 , \33326 , \33327 , \33328 , \33329 , \33330 , \33331 , \33332 , \33333 , \33334 ,
         \33335 , \33336 , \33337 , \33338 , \33339 , \33340 , \33341 , \33342 , \33343 , \33344 ,
         \33345 , \33346 , \33347 , \33348 , \33349 , \33350 , \33351 , \33352 , \33353 , \33354 ,
         \33355 , \33356 , \33357 , \33358 , \33359 , \33360 , \33361 , \33362 , \33363 , \33364 ,
         \33365 , \33366 , \33367 , \33368 , \33369 , \33370 , \33371 , \33372 , \33373 , \33374 ,
         \33375 , \33376 , \33377 , \33378 , \33379 , \33380 , \33381 , \33382 , \33383 , \33384 ,
         \33385 , \33386 , \33387 , \33388 , \33389 , \33390 , \33391 , \33392 , \33393 , \33394 ,
         \33395 , \33396 , \33397 , \33398 , \33399 , \33400 , \33401 , \33402 , \33403 , \33404 ,
         \33405 , \33406 , \33407 , \33408 , \33409 , \33410 , \33411 , \33412 , \33413 , \33414 ,
         \33415 , \33416 , \33417 , \33418 , \33419 , \33420 , \33421 , \33422 , \33423 , \33424 ,
         \33425 , \33426 , \33427 , \33428 , \33429 , \33430 , \33431 , \33432 , \33433 , \33434 ,
         \33435 , \33436 , \33437 , \33438 , \33439 , \33440 , \33441 , \33442 , \33443 , \33444 ,
         \33445 , \33446 , \33447 , \33448 , \33449 , \33450 , \33451 , \33452 , \33453 , \33454 ,
         \33455 , \33456 , \33457 , \33458 , \33459 , \33460 , \33461 , \33462 , \33463 , \33464 ,
         \33465 , \33466 , \33467 , \33468 , \33469 , \33470 , \33471 , \33472 , \33473 , \33474 ,
         \33475 , \33476 , \33477 , \33478 , \33479 , \33480 , \33481 , \33482 , \33483 , \33484 ,
         \33485 , \33486 , \33487 , \33488 , \33489 , \33490 , \33491 , \33492 , \33493 , \33494 ,
         \33495 , \33496 , \33497 , \33498 , \33499 , \33500 , \33501 , \33502 , \33503 , \33504 ,
         \33505 , \33506 , \33507 , \33508 , \33509 , \33510 , \33511 , \33512 , \33513 , \33514 ,
         \33515 , \33516 , \33517 , \33518 , \33519 , \33520 , \33521 , \33522 , \33523 , \33524 ,
         \33525 , \33526 , \33527 , \33528 , \33529 , \33530 , \33531 , \33532 , \33533 , \33534 ,
         \33535 , \33536 , \33537 , \33538 , \33539 , \33540 , \33541 , \33542 , \33543 , \33544 ,
         \33545 , \33546 , \33547 , \33548 , \33549 , \33550 , \33551 , \33552 , \33553 , \33554 ,
         \33555 , \33556 , \33557 , \33558 , \33559 , \33560 , \33561 , \33562 , \33563 , \33564 ,
         \33565 , \33566 , \33567 , \33568 , \33569 , \33570 , \33571 , \33572 , \33573 , \33574 ,
         \33575 , \33576 , \33577 , \33578 , \33579 , \33580 , \33581 , \33582 , \33583 , \33584 ,
         \33585 , \33586 , \33587 , \33588 , \33589 , \33590 , \33591 , \33592 , \33593 , \33594 ,
         \33595 , \33596 , \33597 , \33598 , \33599 , \33600 , \33601 , \33602 , \33603 , \33604 ,
         \33605 , \33606 , \33607 , \33608 , \33609 , \33610 , \33611 , \33612 , \33613 , \33614 ,
         \33615 , \33616 , \33617 , \33618 , \33619 , \33620 , \33621 , \33622 , \33623 , \33624 ,
         \33625 , \33626 , \33627 , \33628 , \33629 , \33630 , \33631 , \33632 , \33633 , \33634 ,
         \33635 , \33636 , \33637 , \33638 , \33639 , \33640 , \33641 , \33642 , \33643 , \33644 ,
         \33645 , \33646 , \33647 , \33648 , \33649 , \33650 , \33651 , \33652 , \33653 , \33654 ,
         \33655 , \33656 , \33657 , \33658 , \33659 , \33660 , \33661 , \33662 , \33663 , \33664 ,
         \33665 , \33666 , \33667 , \33668 , \33669 , \33670 , \33671 , \33672 , \33673 , \33674 ,
         \33675 , \33676 , \33677 , \33678 , \33679 , \33680 , \33681 , \33682 , \33683 , \33684 ,
         \33685 , \33686 , \33687 , \33688 , \33689 , \33690 , \33691 , \33692 , \33693 , \33694 ,
         \33695 , \33696 , \33697 , \33698 , \33699 , \33700 , \33701 , \33702 , \33703 , \33704 ,
         \33705 , \33706 , \33707 , \33708 , \33709 , \33710 , \33711 , \33712 , \33713 , \33714 ,
         \33715 , \33716 , \33717 , \33718 , \33719 , \33720 , \33721 , \33722 , \33723 , \33724 ,
         \33725 , \33726 , \33727 , \33728 , \33729 , \33730 , \33731 , \33732 , \33733 , \33734 ,
         \33735 , \33736 , \33737 , \33738 , \33739 , \33740 , \33741 , \33742 , \33743 , \33744 ,
         \33745 , \33746 , \33747 , \33748 , \33749 , \33750 , \33751 , \33752 , \33753 , \33754 ,
         \33755 , \33756 , \33757 , \33758 , \33759 , \33760 , \33761 , \33762 , \33763 , \33764 ,
         \33765 , \33766 , \33767 , \33768 , \33769 , \33770 , \33771 , \33772 , \33773 , \33774 ,
         \33775 , \33776 , \33777 , \33778 , \33779 , \33780 , \33781 , \33782 , \33783 , \33784 ,
         \33785 , \33786 , \33787 , \33788 , \33789 , \33790 , \33791 , \33792 , \33793 , \33794 ,
         \33795 , \33796 , \33797 , \33798 , \33799 , \33800 , \33801 , \33802 , \33803 , \33804 ,
         \33805 , \33806 , \33807 , \33808 , \33809 , \33810 , \33811 , \33812 , \33813 , \33814 ,
         \33815 , \33816 , \33817 , \33818 , \33819 , \33820 , \33821 , \33822 , \33823 , \33824 ,
         \33825 , \33826 , \33827 , \33828 , \33829 , \33830 , \33831 , \33832 , \33833 , \33834 ,
         \33835 , \33836 , \33837 , \33838 , \33839 , \33840 , \33841 , \33842 , \33843 , \33844 ,
         \33845 , \33846 , \33847 , \33848 , \33849 , \33850 , \33851 , \33852 , \33853 , \33854 ,
         \33855 , \33856 , \33857 , \33858 , \33859 , \33860 , \33861 , \33862 , \33863 , \33864 ,
         \33865 , \33866 , \33867 , \33868 , \33869 , \33870 , \33871 , \33872 , \33873 , \33874 ,
         \33875 , \33876 , \33877 , \33878 , \33879 , \33880 , \33881 , \33882 , \33883 , \33884 ,
         \33885 , \33886 , \33887 , \33888 , \33889 , \33890 , \33891 , \33892 , \33893 , \33894 ,
         \33895 , \33896 , \33897 , \33898 , \33899 , \33900 , \33901 , \33902 , \33903 , \33904 ,
         \33905 , \33906 , \33907 , \33908 , \33909 , \33910 , \33911 , \33912 , \33913 , \33914 ,
         \33915 , \33916 , \33917 , \33918 , \33919 , \33920 , \33921 , \33922 , \33923 , \33924 ,
         \33925 , \33926 , \33927 , \33928 , \33929 , \33930 , \33931 , \33932 , \33933 , \33934 ,
         \33935 , \33936 , \33937 , \33938 , \33939 , \33940 , \33941 , \33942 , \33943 , \33944 ,
         \33945 , \33946 , \33947 , \33948 , \33949 , \33950 , \33951 , \33952 , \33953 , \33954 ,
         \33955 , \33956 , \33957 , \33958 , \33959 , \33960 , \33961 , \33962 , \33963 , \33964 ,
         \33965 , \33966 , \33967 , \33968 , \33969 , \33970 , \33971 , \33972 , \33973 , \33974 ,
         \33975 , \33976 , \33977 , \33978 , \33979 , \33980 , \33981 , \33982 , \33983 , \33984 ,
         \33985 , \33986 , \33987 , \33988 , \33989 , \33990 , \33991 , \33992 , \33993 , \33994 ,
         \33995 , \33996 , \33997 , \33998 , \33999 , \34000 , \34001 , \34002 , \34003 , \34004 ,
         \34005 , \34006 , \34007 , \34008 , \34009 , \34010 , \34011 , \34012 , \34013 , \34014 ,
         \34015 , \34016 , \34017 , \34018 , \34019 , \34020 , \34021 , \34022 , \34023 , \34024 ,
         \34025 , \34026 , \34027 , \34028 , \34029 , \34030 , \34031 , \34032 , \34033 , \34034 ,
         \34035 , \34036 , \34037 , \34038 , \34039 , \34040 , \34041 , \34042 , \34043 , \34044 ,
         \34045 , \34046 , \34047 , \34048 , \34049 , \34050 , \34051 , \34052 , \34053 , \34054 ,
         \34055 , \34056 , \34057 , \34058 , \34059 , \34060 , \34061 , \34062 , \34063 , \34064 ,
         \34065 , \34066 , \34067 , \34068 , \34069 , \34070 , \34071 , \34072 , \34073 , \34074 ,
         \34075 , \34076 , \34077 , \34078 , \34079 , \34080 , \34081 , \34082 , \34083 , \34084 ,
         \34085 , \34086 , \34087 , \34088 , \34089 , \34090 , \34091 , \34092 , \34093 , \34094 ,
         \34095 , \34096 , \34097 , \34098 , \34099 , \34100 , \34101 , \34102 , \34103 , \34104 ,
         \34105 , \34106 , \34107 , \34108 , \34109 , \34110 , \34111 , \34112 , \34113 , \34114 ,
         \34115 , \34116 , \34117 , \34118 , \34119 , \34120 , \34121 , \34122 , \34123 , \34124 ,
         \34125 , \34126 , \34127 , \34128 , \34129 , \34130 , \34131 , \34132 , \34133 , \34134 ,
         \34135 , \34136 , \34137 , \34138 , \34139 , \34140 , \34141 , \34142 , \34143 , \34144 ,
         \34145 , \34146 , \34147 , \34148 , \34149 , \34150 , \34151 , \34152 , \34153 , \34154 ,
         \34155 , \34156 , \34157 , \34158 , \34159 , \34160 , \34161 , \34162 , \34163 , \34164 ,
         \34165 , \34166 , \34167 , \34168 , \34169 , \34170 , \34171 , \34172 , \34173 , \34174 ,
         \34175 , \34176 , \34177 , \34178 , \34179 , \34180 , \34181 , \34182 , \34183 , \34184 ,
         \34185 , \34186 , \34187 , \34188 , \34189 , \34190 , \34191 , \34192 , \34193 , \34194 ,
         \34195 , \34196 , \34197 , \34198 , \34199 , \34200 , \34201 , \34202 , \34203 , \34204 ,
         \34205 , \34206 , \34207 , \34208 , \34209 , \34210 , \34211 , \34212 , \34213 , \34214 ,
         \34215 , \34216 , \34217 , \34218 , \34219 , \34220 , \34221 , \34222 , \34223 , \34224 ,
         \34225 , \34226 , \34227 , \34228 , \34229 , \34230 , \34231 , \34232 , \34233 , \34234 ,
         \34235 , \34236 , \34237 , \34238 , \34239 , \34240 , \34241 , \34242 , \34243 , \34244 ,
         \34245 , \34246 , \34247 , \34248 , \34249 , \34250 , \34251 , \34252 , \34253 , \34254 ,
         \34255 , \34256 , \34257 , \34258 , \34259 , \34260 , \34261 , \34262 , \34263 , \34264 ,
         \34265 , \34266 , \34267 , \34268 , \34269 , \34270 , \34271 , \34272 , \34273 , \34274 ,
         \34275 , \34276 , \34277 , \34278 , \34279 , \34280 , \34281 , \34282 , \34283 , \34284 ,
         \34285 , \34286 , \34287 , \34288 , \34289 , \34290 , \34291 , \34292 , \34293 , \34294 ,
         \34295 , \34296 , \34297 , \34298 , \34299 , \34300 , \34301 , \34302 , \34303 , \34304 ,
         \34305 , \34306 , \34307 , \34308 , \34309 , \34310 , \34311 , \34312 , \34313 , \34314 ,
         \34315 , \34316 , \34317 , \34318 , \34319 , \34320 , \34321 , \34322 , \34323 , \34324 ,
         \34325 , \34326 , \34327 , \34328 , \34329 , \34330 , \34331 , \34332 , \34333 , \34334 ,
         \34335 , \34336 , \34337 , \34338 , \34339 , \34340 , \34341 , \34342 , \34343 , \34344 ,
         \34345 , \34346 , \34347 , \34348 , \34349 , \34350 , \34351 , \34352 , \34353 , \34354 ,
         \34355 , \34356 , \34357 , \34358 , \34359 , \34360 , \34361 , \34362 , \34363 , \34364 ,
         \34365 , \34366 , \34367 , \34368 , \34369 , \34370 , \34371 , \34372 , \34373 , \34374 ,
         \34375 , \34376 , \34377 , \34378 , \34379 , \34380 , \34381 , \34382 , \34383 , \34384 ,
         \34385 , \34386 , \34387 , \34388 , \34389 , \34390 , \34391 , \34392 , \34393 , \34394 ,
         \34395 , \34396 , \34397 , \34398 , \34399 , \34400 , \34401 , \34402 , \34403 , \34404 ,
         \34405 , \34406 , \34407 , \34408 , \34409 , \34410 , \34411 , \34412 , \34413 , \34414 ,
         \34415 , \34416 , \34417 , \34418 , \34419 , \34420 , \34421 , \34422 , \34423 , \34424 ,
         \34425 , \34426 , \34427 , \34428 , \34429 , \34430 , \34431 , \34432 , \34433 , \34434 ,
         \34435 , \34436 , \34437 , \34438 , \34439 , \34440 , \34441 , \34442 , \34443 , \34444 ,
         \34445 , \34446 , \34447 , \34448 , \34449 , \34450 , \34451 , \34452 , \34453 , \34454 ,
         \34455 , \34456 , \34457 , \34458 , \34459 , \34460 , \34461 , \34462 , \34463 , \34464 ,
         \34465 , \34466 , \34467 , \34468 , \34469 , \34470 , \34471 , \34472 , \34473 , \34474 ,
         \34475 , \34476 , \34477 , \34478 , \34479 , \34480 , \34481 , \34482 , \34483 , \34484 ,
         \34485 , \34486 , \34487 , \34488 , \34489 , \34490 , \34491 , \34492 , \34493 , \34494 ,
         \34495 , \34496 , \34497 , \34498 , \34499 , \34500 , \34501 , \34502 , \34503 , \34504 ,
         \34505 , \34506 , \34507 , \34508 , \34509 , \34510 , \34511 , \34512 , \34513 , \34514 ,
         \34515 , \34516 , \34517 , \34518 , \34519 , \34520 , \34521 , \34522 , \34523 , \34524 ,
         \34525 , \34526 , \34527 , \34528 , \34529 , \34530 , \34531 , \34532 , \34533 , \34534 ,
         \34535 , \34536 , \34537 , \34538 , \34539 , \34540 , \34541 , \34542 , \34543 , \34544 ,
         \34545 , \34546 , \34547 , \34548 , \34549 , \34550 , \34551 , \34552 , \34553 , \34554 ,
         \34555 , \34556 , \34557 , \34558 , \34559 , \34560 , \34561 , \34562 , \34563 , \34564 ,
         \34565 , \34566 , \34567 , \34568 , \34569 , \34570 , \34571 , \34572 , \34573 , \34574 ,
         \34575 , \34576 , \34577 , \34578 , \34579 , \34580 , \34581 , \34582 , \34583 , \34584 ,
         \34585 , \34586 , \34587 , \34588 , \34589 , \34590 , \34591 , \34592 , \34593 , \34594 ,
         \34595 , \34596 , \34597 , \34598 , \34599 , \34600 , \34601 , \34602 , \34603 , \34604 ,
         \34605 , \34606 , \34607 , \34608 , \34609 , \34610 , \34611 , \34612 , \34613 , \34614 ,
         \34615 , \34616 , \34617 , \34618 , \34619 , \34620 , \34621 , \34622 , \34623 , \34624 ,
         \34625 , \34626 , \34627 , \34628 , \34629 , \34630 , \34631 , \34632 , \34633 , \34634 ,
         \34635 , \34636 , \34637 , \34638 , \34639 , \34640 , \34641 , \34642 , \34643 , \34644 ,
         \34645 , \34646 , \34647 , \34648 , \34649 , \34650 , \34651 , \34652 , \34653 , \34654 ,
         \34655 , \34656 , \34657 , \34658 , \34659 , \34660 , \34661 , \34662 , \34663 , \34664 ,
         \34665 , \34666 , \34667 , \34668 , \34669 , \34670 , \34671 , \34672 , \34673 , \34674 ,
         \34675 , \34676 , \34677 , \34678 , \34679 , \34680 , \34681 , \34682 , \34683 , \34684 ,
         \34685 , \34686 , \34687 , \34688 , \34689 , \34690 , \34691 , \34692 , \34693 , \34694 ,
         \34695 , \34696 , \34697 , \34698 , \34699 , \34700 , \34701 , \34702 , \34703 , \34704 ,
         \34705 , \34706 , \34707 , \34708 , \34709 , \34710 , \34711 , \34712 , \34713 , \34714 ,
         \34715 , \34716 , \34717 , \34718 , \34719 , \34720 , \34721 , \34722 , \34723 , \34724 ,
         \34725 , \34726 , \34727 , \34728 , \34729 , \34730 , \34731 , \34732 , \34733 , \34734 ,
         \34735 , \34736 , \34737 , \34738 , \34739 , \34740 , \34741 , \34742 , \34743 , \34744 ,
         \34745 , \34746 , \34747 , \34748 , \34749 , \34750 , \34751 , \34752 , \34753 , \34754 ,
         \34755 , \34756 , \34757 , \34758 , \34759 , \34760 , \34761 , \34762 , \34763 , \34764 ,
         \34765 , \34766 , \34767 , \34768 , \34769 , \34770 , \34771 , \34772 , \34773 , \34774 ,
         \34775 , \34776 , \34777 , \34778 , \34779 , \34780 , \34781 , \34782 , \34783 , \34784 ,
         \34785 , \34786 , \34787 , \34788 , \34789 , \34790 , \34791 , \34792 , \34793 , \34794 ,
         \34795 , \34796 , \34797 , \34798 , \34799 , \34800 , \34801 , \34802 , \34803 , \34804 ,
         \34805 , \34806 , \34807 , \34808 , \34809 , \34810 , \34811 , \34812 , \34813 , \34814 ,
         \34815 , \34816 , \34817 , \34818 , \34819 , \34820 , \34821 , \34822 , \34823 , \34824 ,
         \34825 , \34826 , \34827 , \34828 , \34829 , \34830 , \34831 , \34832 , \34833 , \34834 ,
         \34835 , \34836 , \34837 , \34838 , \34839 , \34840 , \34841 , \34842 , \34843 , \34844 ,
         \34845 , \34846 , \34847 , \34848 , \34849 , \34850 , \34851 , \34852 , \34853 , \34854 ,
         \34855 , \34856 , \34857 , \34858 , \34859 , \34860 , \34861 , \34862 , \34863 , \34864 ,
         \34865 , \34866 , \34867 , \34868 , \34869 , \34870 , \34871 , \34872 , \34873 , \34874 ,
         \34875 , \34876 , \34877 , \34878 , \34879 , \34880 , \34881 , \34882 , \34883 , \34884 ,
         \34885 , \34886 , \34887 , \34888 , \34889 , \34890 , \34891 , \34892 , \34893 , \34894 ,
         \34895 , \34896 , \34897 , \34898 , \34899 , \34900 , \34901 , \34902 , \34903 , \34904 ,
         \34905 , \34906 , \34907 , \34908 , \34909 , \34910 , \34911 , \34912 , \34913 , \34914 ,
         \34915 , \34916 , \34917 , \34918 , \34919 , \34920 , \34921 , \34922 , \34923 , \34924 ,
         \34925 , \34926 , \34927 , \34928 , \34929 , \34930 , \34931 , \34932 , \34933 , \34934 ,
         \34935 , \34936 , \34937 , \34938 , \34939 , \34940 , \34941 , \34942 , \34943 , \34944 ,
         \34945 , \34946 , \34947 , \34948 , \34949 , \34950 , \34951 , \34952 , \34953 , \34954 ,
         \34955 , \34956 , \34957 , \34958 , \34959 , \34960 , \34961 , \34962 , \34963 , \34964 ,
         \34965 , \34966 , \34967 , \34968 , \34969 , \34970 , \34971 , \34972 , \34973 , \34974 ,
         \34975 , \34976 , \34977 , \34978 , \34979 , \34980 , \34981 , \34982 , \34983 , \34984 ,
         \34985 , \34986 , \34987 , \34988 , \34989 , \34990 , \34991 , \34992 , \34993 , \34994 ,
         \34995 , \34996 , \34997 , \34998 , \34999 , \35000 , \35001 , \35002 , \35003 , \35004 ,
         \35005 , \35006 , \35007 , \35008 , \35009 , \35010 , \35011 , \35012 , \35013 , \35014 ,
         \35015 , \35016 , \35017 , \35018 , \35019 , \35020 , \35021 , \35022 , \35023 , \35024 ,
         \35025 , \35026 , \35027 , \35028 , \35029 , \35030 , \35031 , \35032 , \35033 , \35034 ,
         \35035 , \35036 , \35037 , \35038 , \35039 , \35040 , \35041 , \35042 , \35043 , \35044 ,
         \35045 , \35046 , \35047 , \35048 , \35049 , \35050 , \35051 , \35052 , \35053 , \35054 ,
         \35055 , \35056 , \35057 , \35058 , \35059 , \35060 , \35061 , \35062 , \35063 , \35064 ,
         \35065 , \35066 , \35067 , \35068 , \35069 , \35070 , \35071 , \35072 , \35073 , \35074 ,
         \35075 , \35076 , \35077 , \35078 , \35079 , \35080 , \35081 , \35082 , \35083 , \35084 ,
         \35085 , \35086 , \35087 , \35088 , \35089 , \35090 , \35091 , \35092 , \35093 , \35094 ,
         \35095 , \35096 , \35097 , \35098 , \35099 , \35100 , \35101 , \35102 , \35103 , \35104 ,
         \35105 , \35106 , \35107 , \35108 , \35109 , \35110 , \35111 , \35112 , \35113 , \35114 ,
         \35115 , \35116 , \35117 , \35118 , \35119 , \35120 , \35121 , \35122 , \35123 , \35124 ,
         \35125 , \35126 , \35127 , \35128 , \35129 , \35130 , \35131 , \35132 , \35133 , \35134 ,
         \35135 , \35136 , \35137 , \35138 , \35139 , \35140 , \35141 , \35142 , \35143 , \35144 ,
         \35145 , \35146 , \35147 , \35148 , \35149 , \35150 , \35151 , \35152 , \35153 , \35154 ,
         \35155 , \35156 , \35157 , \35158 , \35159 , \35160 , \35161 , \35162 , \35163 , \35164 ,
         \35165 , \35166 , \35167 , \35168 , \35169 , \35170 , \35171 , \35172 , \35173 , \35174 ,
         \35175 , \35176 , \35177 , \35178 , \35179 , \35180 , \35181 , \35182 , \35183 , \35184 ,
         \35185 , \35186 , \35187 , \35188 , \35189 , \35190 , \35191 , \35192 , \35193 , \35194 ,
         \35195 , \35196 , \35197 , \35198 , \35199 , \35200 , \35201 , \35202 , \35203 , \35204 ,
         \35205 , \35206 , \35207 , \35208 , \35209 , \35210 , \35211 , \35212 , \35213 , \35214 ,
         \35215 , \35216 , \35217 , \35218 , \35219 , \35220 , \35221 , \35222 , \35223 , \35224 ,
         \35225 , \35226 , \35227 , \35228 , \35229 , \35230 , \35231 , \35232 , \35233 , \35234 ,
         \35235 , \35236 , \35237 , \35238 , \35239 , \35240 , \35241 , \35242 , \35243 , \35244 ,
         \35245 , \35246 , \35247 , \35248 , \35249 , \35250 , \35251 , \35252 , \35253 , \35254 ,
         \35255 , \35256 , \35257 , \35258 , \35259 , \35260 , \35261 , \35262 , \35263 , \35264 ,
         \35265 , \35266 , \35267 , \35268 , \35269 , \35270 , \35271 , \35272 , \35273 , \35274 ,
         \35275 , \35276 , \35277 , \35278 , \35279 , \35280 , \35281 , \35282 , \35283 , \35284 ,
         \35285 , \35286 , \35287 , \35288 , \35289 , \35290 , \35291 , \35292 , \35293 , \35294 ,
         \35295 , \35296 , \35297 , \35298 , \35299 , \35300 , \35301 , \35302 , \35303 , \35304 ,
         \35305 , \35306 , \35307 , \35308 , \35309 , \35310 , \35311 , \35312 , \35313 , \35314 ,
         \35315 , \35316 , \35317 , \35318 , \35319 , \35320 , \35321 , \35322 , \35323 , \35324 ,
         \35325 , \35326 , \35327 , \35328 , \35329 , \35330 , \35331 , \35332 , \35333 , \35334 ,
         \35335 , \35336 , \35337 , \35338 , \35339 , \35340 , \35341 , \35342 , \35343 , \35344 ,
         \35345 , \35346 , \35347 , \35348 , \35349 , \35350 , \35351 , \35352 , \35353 , \35354 ,
         \35355 , \35356 , \35357 , \35358 , \35359 , \35360 , \35361 , \35362 , \35363 , \35364 ,
         \35365 , \35366 , \35367 , \35368 , \35369 , \35370 , \35371 , \35372 , \35373 , \35374 ,
         \35375 , \35376 , \35377 , \35378 , \35379 , \35380 , \35381 , \35382 , \35383 , \35384 ,
         \35385 , \35386 , \35387 , \35388 , \35389 , \35390 , \35391 , \35392 , \35393 , \35394 ,
         \35395 , \35396 , \35397 , \35398 , \35399 , \35400 , \35401 , \35402 , \35403 , \35404 ,
         \35405 , \35406 , \35407 , \35408 , \35409 , \35410 , \35411 , \35412 , \35413 , \35414 ,
         \35415 , \35416 , \35417 , \35418 , \35419 , \35420 , \35421 , \35422 , \35423 , \35424 ,
         \35425 , \35426 , \35427 , \35428 , \35429 , \35430 , \35431 , \35432 , \35433 , \35434 ,
         \35435 , \35436 , \35437 , \35438 , \35439 , \35440 , \35441 , \35442 , \35443 , \35444 ,
         \35445 , \35446 , \35447 , \35448 , \35449 , \35450 , \35451 , \35452 , \35453 , \35454 ,
         \35455 , \35456 , \35457 , \35458 , \35459 , \35460 , \35461 , \35462 , \35463 , \35464 ,
         \35465 , \35466 , \35467 , \35468 , \35469 , \35470 , \35471 , \35472 , \35473 , \35474 ,
         \35475 , \35476 , \35477 , \35478 , \35479 , \35480 , \35481 , \35482 , \35483 , \35484 ,
         \35485 , \35486 , \35487 , \35488 , \35489 , \35490 , \35491 , \35492 , \35493 , \35494 ,
         \35495 , \35496 , \35497 , \35498 , \35499 , \35500 , \35501 , \35502 , \35503 , \35504 ,
         \35505 , \35506 , \35507 , \35508 , \35509 , \35510 , \35511 , \35512 , \35513 , \35514 ,
         \35515 , \35516 , \35517 , \35518 , \35519 , \35520 , \35521 , \35522 , \35523 , \35524 ,
         \35525 , \35526 , \35527 , \35528 , \35529 , \35530 , \35531 , \35532 , \35533 , \35534 ,
         \35535 , \35536 , \35537 , \35538 , \35539 , \35540 , \35541 , \35542 , \35543 , \35544 ,
         \35545 , \35546 , \35547 , \35548 , \35549 , \35550 , \35551 , \35552 , \35553 , \35554 ,
         \35555 , \35556 , \35557 , \35558 , \35559 , \35560 , \35561 , \35562 , \35563 , \35564 ,
         \35565 , \35566 , \35567 , \35568 , \35569 , \35570 , \35571 , \35572 , \35573 , \35574 ,
         \35575 , \35576 , \35577 , \35578 , \35579 , \35580 , \35581 , \35582 , \35583 , \35584 ,
         \35585 , \35586 , \35587 , \35588 , \35589 , \35590 , \35591 , \35592 , \35593 , \35594 ,
         \35595 , \35596 , \35597 , \35598 , \35599 , \35600 , \35601 , \35602 , \35603 , \35604 ,
         \35605 , \35606 , \35607 , \35608 , \35609 , \35610 , \35611 , \35612 , \35613 , \35614 ,
         \35615 , \35616 , \35617 , \35618 , \35619 , \35620 , \35621 , \35622 , \35623 , \35624 ,
         \35625 , \35626 , \35627 , \35628 , \35629 , \35630 , \35631 , \35632 , \35633 , \35634 ,
         \35635 , \35636 , \35637 , \35638 , \35639 , \35640 , \35641 , \35642 , \35643 , \35644 ,
         \35645 , \35646 , \35647 , \35648 , \35649 , \35650 , \35651 , \35652 , \35653 , \35654 ,
         \35655 , \35656 , \35657 , \35658 , \35659 , \35660 , \35661 , \35662 , \35663 , \35664 ,
         \35665 , \35666 , \35667 , \35668 , \35669 , \35670 , \35671 , \35672 , \35673 , \35674 ,
         \35675 , \35676 , \35677 , \35678 , \35679 , \35680 , \35681 , \35682 , \35683 , \35684 ,
         \35685 , \35686 , \35687 , \35688 , \35689 , \35690 , \35691 , \35692 , \35693 , \35694 ,
         \35695 , \35696 , \35697 , \35698 , \35699 , \35700 , \35701 , \35702 , \35703 , \35704 ,
         \35705 , \35706 , \35707 , \35708 , \35709 , \35710 , \35711 , \35712 , \35713 , \35714 ,
         \35715 , \35716 , \35717 , \35718 , \35719 , \35720 , \35721 , \35722 , \35723 , \35724 ,
         \35725 , \35726 , \35727 , \35728 , \35729 , \35730 , \35731 , \35732 , \35733 , \35734 ,
         \35735 , \35736 , \35737 , \35738 , \35739 , \35740 , \35741 , \35742 , \35743 , \35744 ,
         \35745 , \35746 , \35747 , \35748 , \35749 , \35750 , \35751 , \35752 , \35753 , \35754 ,
         \35755 , \35756 , \35757 , \35758 , \35759 , \35760 , \35761 , \35762 , \35763 , \35764 ,
         \35765 , \35766 , \35767 , \35768 , \35769 , \35770 , \35771 , \35772 , \35773 , \35774 ,
         \35775 , \35776 , \35777 , \35778 , \35779 , \35780 , \35781 , \35782 , \35783 , \35784 ,
         \35785 , \35786 , \35787 , \35788 , \35789 , \35790 , \35791 , \35792 , \35793 , \35794 ,
         \35795 , \35796 , \35797 , \35798 , \35799 , \35800 , \35801 , \35802 , \35803 , \35804 ,
         \35805 , \35806 , \35807 , \35808 , \35809 , \35810 , \35811 , \35812 , \35813 , \35814 ,
         \35815 , \35816 , \35817 , \35818 , \35819 , \35820 , \35821 , \35822 , \35823 , \35824 ,
         \35825 , \35826 , \35827 , \35828 , \35829 , \35830 , \35831 , \35832 , \35833 , \35834 ,
         \35835 , \35836 , \35837 , \35838 , \35839 , \35840 , \35841 , \35842 , \35843 , \35844 ,
         \35845 , \35846 , \35847 , \35848 , \35849 , \35850 , \35851 , \35852 , \35853 , \35854 ,
         \35855 , \35856 , \35857 , \35858 , \35859 , \35860 , \35861 , \35862 , \35863 , \35864 ,
         \35865 , \35866 , \35867 , \35868 , \35869 , \35870 , \35871 , \35872 , \35873 , \35874 ,
         \35875 , \35876 , \35877 , \35878 , \35879 , \35880 , \35881 , \35882 , \35883 , \35884 ,
         \35885 , \35886 , \35887 , \35888 , \35889 , \35890 , \35891 , \35892 , \35893 , \35894 ,
         \35895 , \35896 , \35897 , \35898 , \35899 , \35900 , \35901 , \35902 , \35903 , \35904 ,
         \35905 , \35906 , \35907 , \35908 , \35909 , \35910 , \35911 , \35912 , \35913 , \35914 ,
         \35915 , \35916 , \35917 , \35918 , \35919 , \35920 , \35921 , \35922 , \35923 , \35924 ,
         \35925 , \35926 , \35927 , \35928 , \35929 , \35930 , \35931 , \35932 , \35933 , \35934 ,
         \35935 , \35936 , \35937 , \35938 , \35939 , \35940 , \35941 , \35942 , \35943 , \35944 ,
         \35945 , \35946 , \35947 , \35948 , \35949 , \35950 , \35951 , \35952 , \35953 , \35954 ,
         \35955 , \35956 , \35957 , \35958 , \35959 , \35960 , \35961 , \35962 , \35963 , \35964 ,
         \35965 , \35966 , \35967 , \35968 , \35969 , \35970 , \35971 , \35972 , \35973 , \35974 ,
         \35975 , \35976 , \35977 , \35978 , \35979 , \35980 , \35981 , \35982 , \35983 , \35984 ,
         \35985 , \35986 , \35987 , \35988 , \35989 , \35990 , \35991 , \35992 , \35993 , \35994 ,
         \35995 , \35996 , \35997 , \35998 , \35999 , \36000 , \36001 , \36002 , \36003 , \36004 ,
         \36005 , \36006 , \36007 , \36008 , \36009 , \36010 , \36011 , \36012 , \36013 , \36014 ,
         \36015 , \36016 , \36017 , \36018 , \36019 , \36020 , \36021 , \36022 , \36023 , \36024 ,
         \36025 , \36026 , \36027 , \36028 , \36029 , \36030 , \36031 , \36032 , \36033 , \36034 ,
         \36035 , \36036 , \36037 , \36038 , \36039 , \36040 , \36041 , \36042 , \36043 , \36044 ,
         \36045 , \36046 , \36047 , \36048 , \36049 , \36050 , \36051 , \36052 , \36053 , \36054 ,
         \36055 , \36056 , \36057 , \36058 , \36059 , \36060 , \36061 , \36062 , \36063 , \36064 ,
         \36065 , \36066 , \36067 , \36068 , \36069 , \36070 , \36071 , \36072 , \36073 , \36074 ,
         \36075 , \36076 , \36077 , \36078 , \36079 , \36080 , \36081 , \36082 , \36083 , \36084 ,
         \36085 , \36086 , \36087 , \36088 , \36089 , \36090 , \36091 , \36092 , \36093 , \36094 ,
         \36095 , \36096 , \36097 , \36098 , \36099 , \36100 , \36101 , \36102 , \36103 , \36104 ,
         \36105 , \36106 , \36107 , \36108 , \36109 , \36110 , \36111 , \36112 , \36113 , \36114 ,
         \36115 , \36116 , \36117 , \36118 , \36119 , \36120 , \36121 , \36122 , \36123 , \36124 ,
         \36125 , \36126 , \36127 , \36128 , \36129 , \36130 , \36131 , \36132 , \36133 , \36134 ,
         \36135 , \36136 , \36137 , \36138 , \36139 , \36140 , \36141 , \36142 , \36143 , \36144 ,
         \36145 , \36146 , \36147 , \36148 , \36149 , \36150 , \36151 , \36152 , \36153 , \36154 ,
         \36155 , \36156 , \36157 , \36158 , \36159 , \36160 , \36161 , \36162 , \36163 , \36164 ,
         \36165 , \36166 , \36167 , \36168 , \36169 , \36170 , \36171 , \36172 , \36173 , \36174 ,
         \36175 , \36176 , \36177 , \36178 , \36179 , \36180 , \36181 , \36182 , \36183 , \36184 ,
         \36185 , \36186 , \36187 , \36188 , \36189 , \36190 , \36191 , \36192 , \36193 , \36194 ,
         \36195 , \36196 , \36197 , \36198 , \36199 , \36200 , \36201 , \36202 , \36203 , \36204 ,
         \36205 , \36206 , \36207 , \36208 , \36209 , \36210 , \36211 , \36212 , \36213 , \36214 ,
         \36215 , \36216 , \36217 , \36218 , \36219 , \36220 , \36221 , \36222 , \36223 , \36224 ,
         \36225 , \36226 , \36227 , \36228 , \36229 , \36230 , \36231 , \36232 , \36233 , \36234 ,
         \36235 , \36236 , \36237 , \36238 , \36239 , \36240 , \36241 , \36242 , \36243 , \36244 ,
         \36245 , \36246 , \36247 , \36248 , \36249 , \36250 , \36251 , \36252 , \36253 , \36254 ,
         \36255 , \36256 , \36257 , \36258 , \36259 , \36260 , \36261 , \36262 , \36263 , \36264 ,
         \36265 , \36266 , \36267 , \36268 , \36269 , \36270 , \36271 , \36272 , \36273 , \36274 ,
         \36275 , \36276 , \36277 , \36278 , \36279 , \36280 , \36281 , \36282 , \36283 , \36284 ,
         \36285 , \36286 , \36287 , \36288 , \36289 , \36290 , \36291 , \36292 , \36293 , \36294 ,
         \36295 , \36296 , \36297 , \36298 , \36299 , \36300 , \36301 , \36302 , \36303 , \36304 ,
         \36305 , \36306 , \36307 , \36308 , \36309 , \36310 , \36311 , \36312 , \36313 , \36314 ,
         \36315 , \36316 , \36317 , \36318 , \36319 , \36320 , \36321 , \36322 , \36323 , \36324 ,
         \36325 , \36326 , \36327 , \36328 , \36329 , \36330 , \36331 , \36332 , \36333 , \36334 ,
         \36335 , \36336 , \36337 , \36338 , \36339 , \36340 , \36341 , \36342 , \36343 , \36344 ,
         \36345 , \36346 , \36347 , \36348 , \36349 , \36350 , \36351 , \36352 , \36353 , \36354 ,
         \36355 , \36356 , \36357 , \36358 , \36359 , \36360 , \36361 , \36362 , \36363 , \36364 ,
         \36365 , \36366 , \36367 , \36368 , \36369 , \36370 , \36371 , \36372 , \36373 , \36374 ,
         \36375 , \36376 , \36377 , \36378 , \36379 , \36380 , \36381 , \36382 , \36383 , \36384 ,
         \36385 , \36386 , \36387 , \36388 , \36389 , \36390 , \36391 , \36392 , \36393 , \36394 ,
         \36395 , \36396 , \36397 , \36398 , \36399 , \36400 , \36401 , \36402 , \36403 , \36404 ,
         \36405 , \36406 , \36407 , \36408 , \36409 , \36410 , \36411 , \36412 , \36413 , \36414 ,
         \36415 , \36416 , \36417 , \36418 , \36419 , \36420 , \36421 , \36422 , \36423 , \36424 ,
         \36425 , \36426 , \36427 , \36428 , \36429 , \36430 , \36431 , \36432 , \36433 , \36434 ,
         \36435 , \36436 , \36437 , \36438 , \36439 , \36440 , \36441 , \36442 , \36443 , \36444 ,
         \36445 , \36446 , \36447 , \36448 , \36449 , \36450 , \36451 , \36452 , \36453 , \36454 ,
         \36455 , \36456 , \36457 , \36458 , \36459 , \36460 , \36461 , \36462 , \36463 , \36464 ,
         \36465 , \36466 , \36467 , \36468 , \36469 , \36470 , \36471 , \36472 , \36473 , \36474 ,
         \36475 , \36476 , \36477 , \36478 , \36479 , \36480 , \36481 , \36482 , \36483 , \36484 ,
         \36485 , \36486 , \36487 , \36488 , \36489 , \36490 , \36491 , \36492 , \36493 , \36494 ,
         \36495 , \36496 , \36497 , \36498 , \36499 , \36500 , \36501 , \36502 , \36503 , \36504 ,
         \36505 , \36506 , \36507 , \36508 , \36509 , \36510 , \36511 , \36512 , \36513 , \36514 ,
         \36515 , \36516 , \36517 , \36518 , \36519 , \36520 , \36521 , \36522 , \36523 , \36524 ,
         \36525 , \36526 , \36527 , \36528 , \36529 , \36530 , \36531 , \36532 , \36533 , \36534 ,
         \36535 , \36536 , \36537 , \36538 , \36539 , \36540 , \36541 , \36542 , \36543 , \36544 ,
         \36545 , \36546 , \36547 , \36548 , \36549 , \36550 , \36551 , \36552 , \36553 , \36554 ,
         \36555 , \36556 , \36557 , \36558 , \36559 , \36560 , \36561 , \36562 , \36563 , \36564 ,
         \36565 , \36566 , \36567 , \36568 , \36569 , \36570 , \36571 , \36572 , \36573 , \36574 ,
         \36575 , \36576 , \36577 , \36578 , \36579 , \36580 , \36581 , \36582 , \36583 , \36584 ,
         \36585 , \36586 , \36587 , \36588 , \36589 , \36590 , \36591 , \36592 , \36593 , \36594 ,
         \36595 , \36596 , \36597 , \36598 , \36599 , \36600 , \36601 , \36602 , \36603 , \36604 ,
         \36605 , \36606 , \36607 , \36608 , \36609 , \36610 , \36611 , \36612 , \36613 , \36614 ,
         \36615 , \36616 , \36617 , \36618 , \36619 , \36620 , \36621 , \36622 , \36623 , \36624 ,
         \36625 , \36626 , \36627 , \36628 , \36629 , \36630 , \36631 , \36632 , \36633 , \36634 ,
         \36635 , \36636 , \36637 , \36638 , \36639 , \36640 , \36641 , \36642 , \36643 , \36644 ,
         \36645 , \36646 , \36647 , \36648 , \36649 , \36650 , \36651 , \36652 , \36653 , \36654 ,
         \36655 , \36656 , \36657 , \36658 , \36659 , \36660 , \36661 , \36662 , \36663 , \36664 ,
         \36665 , \36666 , \36667 , \36668 , \36669 , \36670 , \36671 , \36672 , \36673 , \36674 ,
         \36675 , \36676 , \36677 , \36678 , \36679 , \36680 , \36681 , \36682 , \36683 , \36684 ,
         \36685 , \36686 , \36687 , \36688 , \36689 , \36690 , \36691 , \36692 , \36693 , \36694 ,
         \36695 , \36696 , \36697 , \36698 , \36699 , \36700 , \36701 , \36702 , \36703 , \36704 ,
         \36705 , \36706 , \36707 , \36708 , \36709 , \36710 , \36711 , \36712 , \36713 , \36714 ,
         \36715 , \36716 , \36717 , \36718 , \36719 , \36720 , \36721 , \36722 , \36723 , \36724 ,
         \36725 , \36726 , \36727 , \36728 , \36729 , \36730 , \36731 , \36732 , \36733 , \36734 ,
         \36735 , \36736 , \36737 , \36738 , \36739 , \36740 , \36741 , \36742 , \36743 , \36744 ,
         \36745 , \36746 , \36747 , \36748 , \36749 , \36750 , \36751 , \36752 , \36753 , \36754 ,
         \36755 , \36756 , \36757 , \36758 , \36759 , \36760 , \36761 , \36762 , \36763 , \36764 ,
         \36765 , \36766 , \36767 , \36768 , \36769 , \36770 , \36771 , \36772 , \36773 , \36774 ,
         \36775 , \36776 , \36777 , \36778 , \36779 , \36780 , \36781 , \36782 , \36783 , \36784 ,
         \36785 , \36786 , \36787 , \36788 , \36789 , \36790 , \36791 , \36792 , \36793 , \36794 ,
         \36795 , \36796 , \36797 , \36798 , \36799 , \36800 , \36801 , \36802 , \36803 , \36804 ,
         \36805 , \36806 , \36807 , \36808 , \36809 , \36810 , \36811 , \36812 , \36813 , \36814 ,
         \36815 , \36816 , \36817 , \36818 , \36819 , \36820 , \36821 , \36822 , \36823 , \36824 ,
         \36825 , \36826 , \36827 , \36828 , \36829 , \36830 , \36831 , \36832 , \36833 , \36834 ,
         \36835 , \36836 , \36837 , \36838 , \36839 , \36840 , \36841 , \36842 , \36843 , \36844 ,
         \36845 , \36846 , \36847 , \36848 , \36849 , \36850 , \36851 , \36852 , \36853 , \36854 ,
         \36855 , \36856 , \36857 , \36858 , \36859 , \36860 , \36861 , \36862 , \36863 , \36864 ,
         \36865 , \36866 , \36867 , \36868 , \36869 , \36870 , \36871 , \36872 , \36873 , \36874 ,
         \36875 , \36876 , \36877 , \36878 , \36879 , \36880 , \36881 , \36882 , \36883 , \36884 ,
         \36885 , \36886 , \36887 , \36888 , \36889 , \36890 , \36891 , \36892 , \36893 , \36894 ,
         \36895 , \36896 , \36897 , \36898 , \36899 , \36900 , \36901 , \36902 , \36903 , \36904 ,
         \36905 , \36906 , \36907 , \36908 , \36909 , \36910 , \36911 , \36912 , \36913 , \36914 ,
         \36915 , \36916 , \36917 , \36918 , \36919 , \36920 , \36921 , \36922 , \36923 , \36924 ,
         \36925 , \36926 , \36927 , \36928 , \36929 , \36930 , \36931 , \36932 , \36933 , \36934 ,
         \36935 , \36936 , \36937 , \36938 , \36939 , \36940 , \36941 , \36942 , \36943 , \36944 ,
         \36945 , \36946 , \36947 , \36948 , \36949 , \36950 , \36951 , \36952 , \36953 , \36954 ,
         \36955 , \36956 , \36957 , \36958 , \36959 , \36960 , \36961 , \36962 , \36963 , \36964 ,
         \36965 , \36966 , \36967 , \36968 , \36969 , \36970 , \36971 , \36972 , \36973 , \36974 ,
         \36975 , \36976 , \36977 , \36978 , \36979 , \36980 , \36981 , \36982 , \36983 , \36984 ,
         \36985 , \36986 , \36987 , \36988 , \36989 , \36990 , \36991 , \36992 , \36993 , \36994 ,
         \36995 , \36996 , \36997 , \36998 , \36999 , \37000 , \37001 , \37002 , \37003 , \37004 ,
         \37005 , \37006 , \37007 , \37008 , \37009 , \37010 , \37011 , \37012 , \37013 , \37014 ,
         \37015 , \37016 , \37017 , \37018 , \37019 , \37020 , \37021 , \37022 , \37023 , \37024 ,
         \37025 , \37026 , \37027 , \37028 , \37029 , \37030 , \37031 , \37032 , \37033 , \37034 ,
         \37035 , \37036 , \37037 , \37038 , \37039 , \37040 , \37041 , \37042 , \37043 , \37044 ,
         \37045 , \37046 , \37047 , \37048 , \37049 , \37050 , \37051 , \37052 , \37053 , \37054 ,
         \37055 , \37056 , \37057 , \37058 , \37059 , \37060 , \37061 , \37062 , \37063 , \37064 ,
         \37065 , \37066 , \37067 , \37068 , \37069 , \37070 , \37071 , \37072 , \37073 , \37074 ,
         \37075 , \37076 , \37077 , \37078 , \37079 , \37080 , \37081 , \37082 , \37083 , \37084 ,
         \37085 , \37086 , \37087 , \37088 , \37089 , \37090 , \37091 , \37092 , \37093 , \37094 ,
         \37095 , \37096 , \37097 , \37098 , \37099 , \37100 , \37101 , \37102 , \37103 , \37104 ,
         \37105 , \37106 , \37107 , \37108 , \37109 , \37110 , \37111 , \37112 , \37113 , \37114 ,
         \37115 , \37116 , \37117 , \37118 , \37119 , \37120 , \37121 , \37122 , \37123 , \37124 ,
         \37125 , \37126 , \37127 , \37128 , \37129 , \37130 , \37131 , \37132 , \37133 , \37134 ,
         \37135 , \37136 , \37137 , \37138 , \37139 , \37140 , \37141 , \37142 , \37143 , \37144 ,
         \37145 , \37146 , \37147 , \37148 , \37149 , \37150 , \37151 , \37152 , \37153 , \37154 ,
         \37155 , \37156 , \37157 , \37158 , \37159 , \37160 , \37161 , \37162 , \37163 , \37164 ,
         \37165 , \37166 , \37167 , \37168 , \37169 , \37170 , \37171 , \37172 , \37173 , \37174 ,
         \37175 , \37176 , \37177 , \37178 , \37179 , \37180 , \37181 , \37182 , \37183 , \37184 ,
         \37185 , \37186 , \37187 , \37188 , \37189 , \37190 , \37191 , \37192 , \37193 , \37194 ,
         \37195 , \37196 , \37197 , \37198 , \37199 , \37200 , \37201 , \37202 , \37203 , \37204 ,
         \37205 , \37206 , \37207 , \37208 , \37209 , \37210 , \37211 , \37212 , \37213 , \37214 ,
         \37215 , \37216 , \37217 , \37218 , \37219 , \37220 , \37221 , \37222 , \37223 , \37224 ,
         \37225 , \37226 , \37227 , \37228 , \37229 , \37230 , \37231 , \37232 , \37233 , \37234 ,
         \37235 , \37236 , \37237 , \37238 , \37239 , \37240 , \37241 , \37242 , \37243 , \37244 ,
         \37245 , \37246 , \37247 , \37248 , \37249 , \37250 , \37251 , \37252 , \37253 , \37254 ,
         \37255 , \37256 , \37257 , \37258 , \37259 , \37260 , \37261 , \37262 , \37263 , \37264 ,
         \37265 , \37266 , \37267 , \37268 , \37269 , \37270 , \37271 , \37272 , \37273 , \37274 ,
         \37275 , \37276 , \37277 , \37278 , \37279 , \37280 , \37281 , \37282 , \37283 , \37284 ,
         \37285 , \37286 , \37287 , \37288 , \37289 , \37290 , \37291 , \37292 , \37293 , \37294 ,
         \37295 , \37296 , \37297 , \37298 , \37299 , \37300 , \37301 , \37302 , \37303 , \37304 ,
         \37305 , \37306 , \37307 , \37308 , \37309 , \37310 , \37311 , \37312 , \37313 , \37314 ,
         \37315 , \37316 , \37317 , \37318 , \37319 , \37320 , \37321 , \37322 , \37323 , \37324 ,
         \37325 , \37326 , \37327 , \37328 , \37329 , \37330 , \37331 , \37332 , \37333 , \37334 ,
         \37335 , \37336 , \37337 , \37338 , \37339 , \37340 , \37341 , \37342 , \37343 , \37344 ,
         \37345 , \37346 , \37347 , \37348 , \37349 , \37350 , \37351 , \37352 , \37353 , \37354 ,
         \37355 , \37356 , \37357 , \37358 , \37359 , \37360 , \37361 , \37362 , \37363 , \37364 ,
         \37365 , \37366 , \37367 , \37368 , \37369 , \37370 , \37371 , \37372 , \37373 , \37374 ,
         \37375 , \37376 , \37377 , \37378 , \37379 , \37380 , \37381 , \37382 , \37383 , \37384 ,
         \37385 , \37386 , \37387 , \37388 , \37389 , \37390 , \37391 , \37392 , \37393 , \37394 ,
         \37395 , \37396 , \37397 , \37398 , \37399 , \37400 , \37401 , \37402 , \37403 , \37404 ,
         \37405 , \37406 , \37407 , \37408 , \37409 , \37410 , \37411 , \37412 , \37413 , \37414 ,
         \37415 , \37416 , \37417 , \37418 , \37419 , \37420 , \37421 , \37422 , \37423 , \37424 ,
         \37425 , \37426 , \37427 , \37428 , \37429 , \37430 , \37431 , \37432 , \37433 , \37434 ,
         \37435 , \37436 , \37437 , \37438 , \37439 , \37440 , \37441 , \37442 , \37443 , \37444 ,
         \37445 , \37446 , \37447 , \37448 , \37449 , \37450 , \37451 , \37452 , \37453 , \37454 ,
         \37455 , \37456 , \37457 , \37458 , \37459 , \37460 , \37461 , \37462 , \37463 , \37464 ,
         \37465 , \37466 , \37467 , \37468 , \37469 , \37470 , \37471 , \37472 , \37473 , \37474 ,
         \37475 , \37476 , \37477 , \37478 , \37479 , \37480 , \37481 , \37482 , \37483 , \37484 ,
         \37485 , \37486 , \37487 , \37488 , \37489 , \37490 , \37491 , \37492 , \37493 , \37494 ,
         \37495 , \37496 , \37497 , \37498 , \37499 , \37500 , \37501 , \37502 , \37503 , \37504 ,
         \37505 , \37506 , \37507 , \37508 , \37509 , \37510 , \37511 , \37512 , \37513 , \37514 ,
         \37515 , \37516 , \37517 , \37518 , \37519 , \37520 , \37521 , \37522 , \37523 , \37524 ,
         \37525 , \37526 , \37527 , \37528 , \37529 , \37530 , \37531 , \37532 , \37533 , \37534 ,
         \37535 , \37536 , \37537 , \37538 , \37539 , \37540 , \37541 , \37542 , \37543 , \37544 ,
         \37545 , \37546 , \37547 , \37548 , \37549 , \37550 , \37551 , \37552 , \37553 , \37554 ,
         \37555 , \37556 , \37557 , \37558 , \37559 , \37560 , \37561 , \37562 , \37563 , \37564 ,
         \37565 , \37566 , \37567 , \37568 , \37569 , \37570 , \37571 , \37572 , \37573 , \37574 ,
         \37575 , \37576 , \37577 , \37578 , \37579 , \37580 , \37581 , \37582 , \37583 , \37584 ,
         \37585 , \37586 , \37587 , \37588 , \37589 , \37590 , \37591 , \37592 , \37593 , \37594 ,
         \37595 , \37596 , \37597 , \37598 , \37599 , \37600 , \37601 , \37602 , \37603 , \37604 ,
         \37605 , \37606 , \37607 , \37608 , \37609 , \37610 , \37611 , \37612 , \37613 , \37614 ,
         \37615 , \37616 , \37617 , \37618 , \37619 , \37620 , \37621 , \37622 , \37623 , \37624 ,
         \37625 , \37626 , \37627 , \37628 , \37629 , \37630 , \37631 , \37632 , \37633 , \37634 ,
         \37635 , \37636 , \37637 , \37638 , \37639 , \37640 , \37641 , \37642 , \37643 , \37644 ,
         \37645 , \37646 , \37647 , \37648 , \37649 , \37650 , \37651 , \37652 , \37653 , \37654 ,
         \37655 , \37656 , \37657 , \37658 , \37659 , \37660 , \37661 , \37662 , \37663 , \37664 ,
         \37665 , \37666 , \37667 , \37668 , \37669 , \37670 , \37671 , \37672 , \37673 , \37674 ,
         \37675 , \37676 , \37677 , \37678 , \37679 , \37680 , \37681 , \37682 , \37683 , \37684 ,
         \37685 , \37686 , \37687 , \37688 , \37689 , \37690 , \37691 , \37692 , \37693 , \37694 ,
         \37695 , \37696 , \37697 , \37698 , \37699 , \37700 , \37701 , \37702 , \37703 , \37704 ,
         \37705 , \37706 , \37707 , \37708 , \37709 , \37710 , \37711 , \37712 , \37713 , \37714 ,
         \37715 , \37716 , \37717 , \37718 , \37719 , \37720 , \37721 , \37722 , \37723 , \37724 ,
         \37725 , \37726 , \37727 , \37728 , \37729 , \37730 , \37731 , \37732 , \37733 , \37734 ,
         \37735 , \37736 , \37737 , \37738 , \37739 , \37740 , \37741 , \37742 , \37743 , \37744 ,
         \37745 , \37746 , \37747 , \37748 , \37749 , \37750 , \37751 , \37752 , \37753 , \37754 ,
         \37755 , \37756 , \37757 , \37758 , \37759 , \37760 , \37761 , \37762 , \37763 , \37764 ,
         \37765 , \37766 , \37767 , \37768 , \37769 , \37770 , \37771 , \37772 , \37773 , \37774 ,
         \37775 , \37776 , \37777 , \37778 , \37779 , \37780 , \37781 , \37782 , \37783 , \37784 ,
         \37785 , \37786 , \37787 , \37788 , \37789 , \37790 , \37791 , \37792 , \37793 , \37794 ,
         \37795 , \37796 , \37797 , \37798 , \37799 , \37800 , \37801 , \37802 , \37803 , \37804 ,
         \37805 , \37806 , \37807 , \37808 , \37809 , \37810 , \37811 , \37812 , \37813 , \37814 ,
         \37815 , \37816 , \37817 , \37818 , \37819 , \37820 , \37821 , \37822 , \37823 , \37824 ,
         \37825 , \37826 , \37827 , \37828 , \37829 , \37830 , \37831 , \37832 , \37833 , \37834 ,
         \37835 , \37836 , \37837 , \37838 , \37839 , \37840 , \37841 , \37842 , \37843 , \37844 ,
         \37845 , \37846 , \37847 , \37848 , \37849 , \37850 , \37851 , \37852 , \37853 , \37854 ,
         \37855 , \37856 , \37857 , \37858 , \37859 , \37860 , \37861 , \37862 , \37863 , \37864 ,
         \37865 , \37866 , \37867 , \37868 , \37869 , \37870 , \37871 , \37872 , \37873 , \37874 ,
         \37875 , \37876 , \37877 , \37878 , \37879 , \37880 , \37881 , \37882 , \37883 , \37884 ,
         \37885 , \37886 , \37887 , \37888 , \37889 , \37890 , \37891 , \37892 , \37893 , \37894 ,
         \37895 , \37896 , \37897 , \37898 , \37899 , \37900 , \37901 , \37902 , \37903 , \37904 ,
         \37905 , \37906 , \37907 , \37908 , \37909 , \37910 , \37911 , \37912 , \37913 , \37914 ,
         \37915 , \37916 , \37917 , \37918 , \37919 , \37920 , \37921 , \37922 , \37923 , \37924 ,
         \37925 , \37926 , \37927 , \37928 , \37929 , \37930 , \37931 , \37932 , \37933 , \37934 ,
         \37935 , \37936 , \37937 , \37938 , \37939 , \37940 , \37941 , \37942 , \37943 , \37944 ,
         \37945 , \37946 , \37947 , \37948 , \37949 , \37950 , \37951 , \37952 , \37953 , \37954 ,
         \37955 , \37956 , \37957 , \37958 , \37959 , \37960 , \37961 , \37962 , \37963 , \37964 ,
         \37965 , \37966 , \37967 , \37968 , \37969 , \37970 , \37971 , \37972 , \37973 , \37974 ,
         \37975 , \37976 , \37977 , \37978 , \37979 , \37980 , \37981 , \37982 , \37983 , \37984 ,
         \37985 , \37986 , \37987 , \37988 , \37989 , \37990 , \37991 , \37992 , \37993 , \37994 ,
         \37995 , \37996 , \37997 , \37998 , \37999 , \38000 , \38001 , \38002 , \38003 , \38004 ,
         \38005 , \38006 , \38007 , \38008 , \38009 , \38010 , \38011 , \38012 , \38013 , \38014 ,
         \38015 , \38016 , \38017 , \38018 , \38019 , \38020 , \38021 , \38022 , \38023 , \38024 ,
         \38025 , \38026 , \38027 , \38028 , \38029 , \38030 , \38031 , \38032 , \38033 , \38034 ,
         \38035 , \38036 , \38037 , \38038 , \38039 , \38040 , \38041 , \38042 , \38043 , \38044 ,
         \38045 , \38046 , \38047 , \38048 , \38049 , \38050 , \38051 , \38052 , \38053 , \38054 ,
         \38055 , \38056 , \38057 , \38058 , \38059 , \38060 , \38061 , \38062 , \38063 , \38064 ,
         \38065 , \38066 , \38067 , \38068 , \38069 , \38070 , \38071 , \38072 , \38073 , \38074 ,
         \38075 , \38076 , \38077 , \38078 , \38079 , \38080 , \38081 , \38082 , \38083 , \38084 ,
         \38085 , \38086 , \38087 , \38088 , \38089 , \38090 , \38091 , \38092 , \38093 , \38094 ,
         \38095 , \38096 , \38097 , \38098 , \38099 , \38100 , \38101 , \38102 , \38103 , \38104 ,
         \38105 , \38106 , \38107 , \38108 , \38109 , \38110 , \38111 , \38112 , \38113 , \38114 ,
         \38115 , \38116 , \38117 , \38118 , \38119 , \38120 , \38121 , \38122 , \38123 , \38124 ,
         \38125 , \38126 , \38127 , \38128 , \38129 , \38130 , \38131 , \38132 , \38133 , \38134 ,
         \38135 , \38136 , \38137 , \38138 , \38139 , \38140 , \38141 , \38142 , \38143 , \38144 ,
         \38145 , \38146 , \38147 , \38148 , \38149 , \38150 , \38151 , \38152 , \38153 , \38154 ,
         \38155 , \38156 , \38157 , \38158 , \38159 , \38160 , \38161 , \38162 , \38163 , \38164 ,
         \38165 , \38166 , \38167 , \38168 , \38169 , \38170 , \38171 , \38172 , \38173 , \38174 ,
         \38175 , \38176 , \38177 , \38178 , \38179 , \38180 , \38181 , \38182 , \38183 , \38184 ,
         \38185 , \38186 , \38187 , \38188 , \38189 , \38190 , \38191 , \38192 , \38193 , \38194 ,
         \38195 , \38196 , \38197 , \38198 , \38199 , \38200 , \38201 , \38202 , \38203 , \38204 ,
         \38205 , \38206 , \38207 , \38208 , \38209 , \38210 , \38211 , \38212 , \38213 , \38214 ,
         \38215 , \38216 , \38217 , \38218 , \38219 , \38220 , \38221 , \38222 , \38223 , \38224 ,
         \38225 , \38226 , \38227 , \38228 , \38229 , \38230 , \38231 , \38232 , \38233 , \38234 ,
         \38235 , \38236 , \38237 , \38238 , \38239 , \38240 , \38241 , \38242 , \38243 , \38244 ,
         \38245 , \38246 , \38247 , \38248 , \38249 , \38250 , \38251 , \38252 , \38253 , \38254 ,
         \38255 , \38256 , \38257 , \38258 , \38259 , \38260 , \38261 , \38262 , \38263 , \38264 ,
         \38265 , \38266 , \38267 , \38268 , \38269 , \38270 , \38271 , \38272 , \38273 , \38274 ,
         \38275 , \38276 , \38277 , \38278 , \38279 , \38280 , \38281 , \38282 , \38283 , \38284 ,
         \38285 , \38286 , \38287 , \38288 , \38289 , \38290 , \38291 , \38292 , \38293 , \38294 ,
         \38295 , \38296 , \38297 , \38298 , \38299 , \38300 , \38301 , \38302 , \38303 , \38304 ,
         \38305 , \38306 , \38307 , \38308 , \38309 , \38310 , \38311 , \38312 , \38313 , \38314 ,
         \38315 , \38316 , \38317 , \38318 , \38319 , \38320 , \38321 , \38322 , \38323 , \38324 ,
         \38325 , \38326 , \38327 , \38328 , \38329 , \38330 , \38331 , \38332 , \38333 , \38334 ,
         \38335 , \38336 , \38337 , \38338 , \38339 , \38340 , \38341 , \38342 , \38343 , \38344 ,
         \38345 , \38346 , \38347 , \38348 , \38349 , \38350 , \38351 , \38352 , \38353 , \38354 ,
         \38355 , \38356 , \38357 , \38358 , \38359 , \38360 , \38361 , \38362 , \38363 , \38364 ,
         \38365 , \38366 , \38367 , \38368 , \38369 , \38370 , \38371 , \38372 , \38373 , \38374 ,
         \38375 , \38376 , \38377 , \38378 , \38379 , \38380 , \38381 , \38382 , \38383 , \38384 ,
         \38385 , \38386 , \38387 , \38388 , \38389 , \38390 , \38391 , \38392 , \38393 , \38394 ,
         \38395 , \38396 , \38397 , \38398 , \38399 , \38400 , \38401 , \38402 , \38403 , \38404 ,
         \38405 , \38406 , \38407 , \38408 , \38409 , \38410 , \38411 , \38412 , \38413 , \38414 ,
         \38415 , \38416 , \38417 , \38418 , \38419 , \38420 , \38421 , \38422 , \38423 , \38424 ,
         \38425 , \38426 , \38427 , \38428 , \38429 , \38430 , \38431 , \38432 , \38433 , \38434 ,
         \38435 , \38436 , \38437 , \38438 , \38439 , \38440 , \38441 , \38442 , \38443 , \38444 ,
         \38445 , \38446 , \38447 , \38448 , \38449 , \38450 , \38451 , \38452 , \38453 , \38454 ,
         \38455 , \38456 , \38457 , \38458 , \38459 , \38460 , \38461 , \38462 , \38463 , \38464 ,
         \38465 , \38466 , \38467 , \38468 , \38469 , \38470 , \38471 , \38472 , \38473 , \38474 ,
         \38475 , \38476 , \38477 , \38478 , \38479 , \38480 , \38481 , \38482 , \38483 , \38484 ,
         \38485 , \38486 , \38487 , \38488 , \38489 , \38490 , \38491 , \38492 , \38493 , \38494 ,
         \38495 , \38496 , \38497 , \38498 , \38499 , \38500 , \38501 , \38502 , \38503 , \38504 ,
         \38505 , \38506 , \38507 , \38508 , \38509 , \38510 , \38511 , \38512 , \38513 , \38514 ,
         \38515 , \38516 , \38517 , \38518 , \38519 , \38520 , \38521 , \38522 , \38523 , \38524 ,
         \38525 , \38526 , \38527 , \38528 , \38529 , \38530 , \38531 , \38532 , \38533 , \38534 ,
         \38535 , \38536 , \38537 , \38538 , \38539 , \38540 , \38541 , \38542 , \38543 , \38544 ,
         \38545 , \38546 , \38547 , \38548 , \38549 , \38550 , \38551 , \38552 , \38553 , \38554 ,
         \38555 , \38556 , \38557 , \38558 , \38559 , \38560 , \38561 , \38562 , \38563 , \38564 ,
         \38565 , \38566 , \38567 , \38568 , \38569 , \38570 , \38571 , \38572 , \38573 , \38574 ,
         \38575 , \38576 , \38577 , \38578 , \38579 , \38580 , \38581 , \38582 , \38583 , \38584 ,
         \38585 , \38586 , \38587 , \38588 , \38589 , \38590 , \38591 , \38592 , \38593 , \38594 ,
         \38595 , \38596 , \38597 , \38598 , \38599 , \38600 , \38601 , \38602 , \38603 , \38604 ,
         \38605 , \38606 , \38607 , \38608 , \38609 , \38610 , \38611 , \38612 , \38613 , \38614 ,
         \38615 , \38616 , \38617 , \38618 , \38619 , \38620 , \38621 , \38622 , \38623 , \38624 ,
         \38625 , \38626 , \38627 , \38628 , \38629 , \38630 , \38631 , \38632 , \38633 , \38634 ,
         \38635 , \38636 , \38637 , \38638 , \38639 , \38640 , \38641 , \38642 , \38643 , \38644 ,
         \38645 , \38646 , \38647 , \38648 , \38649 , \38650 , \38651 , \38652 , \38653 , \38654 ,
         \38655 , \38656 , \38657 , \38658 , \38659 , \38660 , \38661 , \38662 , \38663 , \38664 ,
         \38665 , \38666 , \38667 , \38668 , \38669 , \38670 , \38671 , \38672 , \38673 , \38674 ,
         \38675 , \38676 , \38677 , \38678 , \38679 , \38680 , \38681 , \38682 , \38683 , \38684 ,
         \38685 , \38686 , \38687 , \38688 , \38689 , \38690 , \38691 , \38692 , \38693 , \38694 ,
         \38695 , \38696 , \38697 , \38698 , \38699 , \38700 , \38701 , \38702 , \38703 , \38704 ,
         \38705 , \38706 , \38707 , \38708 , \38709 , \38710 , \38711 , \38712 , \38713 , \38714 ,
         \38715 , \38716 , \38717 , \38718 , \38719 , \38720 , \38721 , \38722 , \38723 , \38724 ,
         \38725 , \38726 , \38727 , \38728 , \38729 , \38730 , \38731 , \38732 , \38733 , \38734 ,
         \38735 , \38736 , \38737 , \38738 , \38739 , \38740 , \38741 , \38742 , \38743 , \38744 ,
         \38745 , \38746 , \38747 , \38748 , \38749 , \38750 , \38751 , \38752 , \38753 , \38754 ,
         \38755 , \38756 , \38757 , \38758 , \38759 , \38760 , \38761 , \38762 , \38763 , \38764 ,
         \38765 , \38766 , \38767 , \38768 , \38769 , \38770 , \38771 , \38772 , \38773 , \38774 ,
         \38775 , \38776 , \38777 , \38778 , \38779 , \38780 , \38781 , \38782 , \38783 , \38784 ,
         \38785 , \38786 , \38787 , \38788 , \38789 , \38790 , \38791 , \38792 , \38793 , \38794 ,
         \38795 , \38796 , \38797 , \38798 , \38799 , \38800 , \38801 , \38802 , \38803 , \38804 ,
         \38805 , \38806 , \38807 , \38808 , \38809 , \38810 , \38811 , \38812 , \38813 , \38814 ,
         \38815 , \38816 , \38817 , \38818 , \38819 , \38820 , \38821 , \38822 , \38823 , \38824 ,
         \38825 , \38826 , \38827 , \38828 , \38829 , \38830 , \38831 , \38832 , \38833 , \38834 ,
         \38835 , \38836 , \38837 , \38838 , \38839 , \38840 , \38841 , \38842 , \38843 , \38844 ,
         \38845 , \38846 , \38847 , \38848 , \38849 , \38850 , \38851 , \38852 , \38853 , \38854 ,
         \38855 , \38856 , \38857 , \38858 , \38859 , \38860 , \38861 , \38862 , \38863 , \38864 ,
         \38865 , \38866 , \38867 , \38868 , \38869 , \38870 , \38871 , \38872 , \38873 , \38874 ,
         \38875 , \38876 , \38877 , \38878 , \38879 , \38880 , \38881 , \38882 , \38883 , \38884 ,
         \38885 , \38886 , \38887 , \38888 , \38889 , \38890 , \38891 , \38892 , \38893 , \38894 ,
         \38895 , \38896 , \38897 , \38898 , \38899 , \38900 , \38901 , \38902 , \38903 , \38904 ,
         \38905 , \38906 , \38907 , \38908 , \38909 , \38910 , \38911 , \38912 , \38913 , \38914 ,
         \38915 , \38916 , \38917 , \38918 , \38919 , \38920 , \38921 , \38922 , \38923 , \38924 ,
         \38925 , \38926 , \38927 , \38928 , \38929 , \38930 , \38931 , \38932 , \38933 , \38934 ,
         \38935 , \38936 , \38937 , \38938 , \38939 , \38940 , \38941 , \38942 , \38943 , \38944 ,
         \38945 , \38946 , \38947 , \38948 , \38949 , \38950 , \38951 , \38952 , \38953 , \38954 ,
         \38955 , \38956 , \38957 , \38958 , \38959 , \38960 , \38961 , \38962 , \38963 , \38964 ,
         \38965 , \38966 , \38967 , \38968 , \38969 , \38970 , \38971 , \38972 , \38973 , \38974 ,
         \38975 , \38976 , \38977 , \38978 , \38979 , \38980 , \38981 , \38982 , \38983 , \38984 ,
         \38985 , \38986 , \38987 , \38988 , \38989 , \38990 , \38991 , \38992 , \38993 , \38994 ,
         \38995 , \38996 , \38997 , \38998 , \38999 , \39000 , \39001 , \39002 , \39003 , \39004 ,
         \39005 , \39006 , \39007 , \39008 , \39009 , \39010 , \39011 , \39012 , \39013 , \39014 ,
         \39015 , \39016 , \39017 , \39018 , \39019 , \39020 , \39021 , \39022 , \39023 , \39024 ,
         \39025 , \39026 , \39027 , \39028 , \39029 , \39030 , \39031 , \39032 , \39033 , \39034 ,
         \39035 , \39036 , \39037 , \39038 , \39039 , \39040 , \39041 , \39042 , \39043 , \39044 ,
         \39045 , \39046 , \39047 , \39048 , \39049 , \39050 , \39051 , \39052 , \39053 , \39054 ,
         \39055 , \39056 , \39057 , \39058 , \39059 , \39060 , \39061 , \39062 , \39063 , \39064 ,
         \39065 , \39066 , \39067 , \39068 , \39069 , \39070 , \39071 , \39072 , \39073 , \39074 ,
         \39075 , \39076 , \39077 , \39078 , \39079 , \39080 , \39081 , \39082 , \39083 , \39084 ,
         \39085 , \39086 , \39087 , \39088 , \39089 , \39090 , \39091 , \39092 , \39093 , \39094 ,
         \39095 , \39096 , \39097 , \39098 , \39099 , \39100 , \39101 , \39102 , \39103 , \39104 ,
         \39105 , \39106 , \39107 , \39108 , \39109 , \39110 , \39111 , \39112 , \39113 , \39114 ,
         \39115 , \39116 , \39117 , \39118 , \39119 , \39120 , \39121 , \39122 , \39123 , \39124 ,
         \39125 , \39126 , \39127 , \39128 , \39129 , \39130 , \39131 , \39132 , \39133 , \39134 ,
         \39135 , \39136 , \39137 , \39138 , \39139 , \39140 , \39141 , \39142 , \39143 , \39144 ,
         \39145 , \39146 , \39147 , \39148 , \39149 , \39150 , \39151 , \39152 , \39153 , \39154 ,
         \39155 , \39156 , \39157 , \39158 , \39159 , \39160 , \39161 , \39162 , \39163 , \39164 ,
         \39165 , \39166 , \39167 , \39168 , \39169 , \39170 , \39171 , \39172 , \39173 , \39174 ,
         \39175 , \39176 , \39177 , \39178 , \39179 , \39180 , \39181 , \39182 , \39183 , \39184 ,
         \39185 , \39186 , \39187 , \39188 , \39189 , \39190 , \39191 , \39192 , \39193 , \39194 ,
         \39195 , \39196 , \39197 , \39198 , \39199 , \39200 , \39201 , \39202 , \39203 , \39204 ,
         \39205 , \39206 , \39207 , \39208 , \39209 , \39210 , \39211 , \39212 , \39213 , \39214 ,
         \39215 , \39216 , \39217 , \39218 , \39219 , \39220 , \39221 , \39222 , \39223 , \39224 ,
         \39225 , \39226 , \39227 , \39228 , \39229 , \39230 , \39231 , \39232 , \39233 , \39234 ,
         \39235 , \39236 , \39237 , \39238 , \39239 , \39240 , \39241 , \39242 , \39243 , \39244 ,
         \39245 , \39246 , \39247 , \39248 , \39249 , \39250 , \39251 , \39252 , \39253 , \39254 ,
         \39255 , \39256 , \39257 , \39258 , \39259 , \39260 , \39261 , \39262 , \39263 , \39264 ,
         \39265 , \39266 , \39267 , \39268 , \39269 , \39270 , \39271 , \39272 , \39273 , \39274 ,
         \39275 , \39276 , \39277 , \39278 , \39279 , \39280 , \39281 , \39282 , \39283 , \39284 ,
         \39285 , \39286 , \39287 , \39288 , \39289 , \39290 , \39291 , \39292 , \39293 , \39294 ,
         \39295 , \39296 , \39297 , \39298 , \39299 , \39300 , \39301 , \39302 , \39303 , \39304 ,
         \39305 , \39306 , \39307 , \39308 , \39309 , \39310 , \39311 , \39312 , \39313 , \39314 ,
         \39315 , \39316 , \39317 , \39318 , \39319 , \39320 , \39321 , \39322 , \39323 , \39324 ,
         \39325 , \39326 , \39327 , \39328 , \39329 , \39330 , \39331 , \39332 , \39333 , \39334 ,
         \39335 , \39336 , \39337 , \39338 , \39339 , \39340 , \39341 , \39342 , \39343 , \39344 ,
         \39345 , \39346 , \39347 , \39348 , \39349 , \39350 , \39351 , \39352 , \39353 , \39354 ,
         \39355 , \39356 , \39357 , \39358 , \39359 , \39360 , \39361 , \39362 , \39363 , \39364 ,
         \39365 , \39366 , \39367 , \39368 , \39369 , \39370 , \39371 , \39372 , \39373 , \39374 ,
         \39375 , \39376 , \39377 , \39378 , \39379 , \39380 , \39381 , \39382 , \39383 , \39384 ,
         \39385 , \39386 , \39387 , \39388 , \39389 , \39390 , \39391 , \39392 , \39393 , \39394 ,
         \39395 , \39396 , \39397 , \39398 , \39399 , \39400 , \39401 , \39402 , \39403 , \39404 ,
         \39405 , \39406 , \39407 , \39408 , \39409 , \39410 , \39411 , \39412 , \39413 , \39414 ,
         \39415 , \39416 , \39417 , \39418 , \39419 , \39420 , \39421 , \39422 , \39423 , \39424 ,
         \39425 , \39426 , \39427 , \39428 , \39429 , \39430 , \39431 , \39432 , \39433 , \39434 ,
         \39435 , \39436 , \39437 , \39438 , \39439 , \39440 , \39441 , \39442 , \39443 , \39444 ,
         \39445 , \39446 , \39447 , \39448 , \39449 , \39450 , \39451 , \39452 , \39453 , \39454 ,
         \39455 , \39456 , \39457 , \39458 , \39459 , \39460 , \39461 , \39462 , \39463 , \39464 ,
         \39465 , \39466 , \39467 , \39468 , \39469 , \39470 , \39471 , \39472 , \39473 , \39474 ,
         \39475 , \39476 , \39477 , \39478 , \39479 , \39480 , \39481 , \39482 , \39483 , \39484 ,
         \39485 , \39486 , \39487 , \39488 , \39489 , \39490 , \39491 , \39492 , \39493 , \39494 ,
         \39495 , \39496 , \39497 , \39498 , \39499 , \39500 , \39501 , \39502 , \39503 , \39504 ,
         \39505 , \39506 , \39507 , \39508 , \39509 , \39510 , \39511 , \39512 , \39513 , \39514 ,
         \39515 , \39516 , \39517 , \39518 , \39519 , \39520 , \39521 , \39522 , \39523 , \39524 ,
         \39525 , \39526 , \39527 , \39528 , \39529 , \39530 , \39531 , \39532 , \39533 , \39534 ,
         \39535 , \39536 , \39537 , \39538 , \39539 , \39540 , \39541 , \39542 , \39543 , \39544 ,
         \39545 , \39546 , \39547 , \39548 , \39549 , \39550 , \39551 , \39552 , \39553 , \39554 ,
         \39555 , \39556 , \39557 , \39558 , \39559 , \39560 , \39561 , \39562 , \39563 , \39564 ,
         \39565 , \39566 , \39567 , \39568 , \39569 , \39570 , \39571 , \39572 , \39573 , \39574 ,
         \39575 , \39576 , \39577 , \39578 , \39579 , \39580 , \39581 , \39582 , \39583 , \39584 ,
         \39585 , \39586 , \39587 , \39588 , \39589 , \39590 , \39591 , \39592 , \39593 , \39594 ,
         \39595 , \39596 , \39597 , \39598 , \39599 , \39600 , \39601 , \39602 , \39603 , \39604 ,
         \39605 , \39606 , \39607 , \39608 , \39609 , \39610 , \39611 , \39612 , \39613 , \39614 ,
         \39615 , \39616 , \39617 , \39618 , \39619 , \39620 , \39621 , \39622 , \39623 , \39624 ,
         \39625 , \39626 , \39627 , \39628 , \39629 , \39630 , \39631 , \39632 , \39633 , \39634 ,
         \39635 , \39636 , \39637 , \39638 , \39639 , \39640 , \39641 , \39642 , \39643 , \39644 ,
         \39645 , \39646 , \39647 , \39648 , \39649 , \39650 , \39651 , \39652 , \39653 , \39654 ,
         \39655 , \39656 , \39657 , \39658 , \39659 , \39660 , \39661 , \39662 , \39663 , \39664 ,
         \39665 , \39666 , \39667 , \39668 , \39669 , \39670 , \39671 , \39672 , \39673 , \39674 ,
         \39675 , \39676 , \39677 , \39678 , \39679 , \39680 , \39681 , \39682 , \39683 , \39684 ,
         \39685 , \39686 , \39687 , \39688 , \39689 , \39690 , \39691 , \39692 , \39693 , \39694 ,
         \39695 , \39696 , \39697 , \39698 , \39699 , \39700 , \39701 , \39702 , \39703 , \39704 ,
         \39705 , \39706 , \39707 , \39708 , \39709 , \39710 , \39711 , \39712 , \39713 , \39714 ,
         \39715 , \39716 , \39717 , \39718 , \39719 , \39720 , \39721 , \39722 , \39723 , \39724 ,
         \39725 , \39726 , \39727 , \39728 , \39729 , \39730 , \39731 , \39732 , \39733 , \39734 ,
         \39735 , \39736 , \39737 , \39738 , \39739 , \39740 , \39741 , \39742 , \39743 , \39744 ,
         \39745 , \39746 , \39747 , \39748 , \39749 , \39750 , \39751 , \39752 , \39753 , \39754 ,
         \39755 , \39756 , \39757 , \39758 , \39759 , \39760 , \39761 , \39762 , \39763 , \39764 ,
         \39765 , \39766 , \39767 , \39768 , \39769 , \39770 , \39771 , \39772 , \39773 , \39774 ,
         \39775 , \39776 , \39777 , \39778 , \39779 , \39780 , \39781 , \39782 , \39783 , \39784 ,
         \39785 , \39786 , \39787 , \39788 , \39789 , \39790 , \39791 , \39792 , \39793 , \39794 ,
         \39795 , \39796 , \39797 , \39798 , \39799 , \39800 , \39801 , \39802 , \39803 , \39804 ,
         \39805 , \39806 , \39807 , \39808 , \39809 , \39810 , \39811 , \39812 , \39813 , \39814 ,
         \39815 , \39816 , \39817 , \39818 , \39819 , \39820 , \39821 , \39822 , \39823 , \39824 ,
         \39825 , \39826 , \39827 , \39828 , \39829 , \39830 , \39831 , \39832 , \39833 , \39834 ,
         \39835 , \39836 , \39837 , \39838 , \39839 , \39840 , \39841 , \39842 , \39843 , \39844 ,
         \39845 , \39846 , \39847 , \39848 , \39849 , \39850 , \39851 , \39852 , \39853 , \39854 ,
         \39855 , \39856 , \39857 , \39858 , \39859 , \39860 , \39861 , \39862 , \39863 , \39864 ,
         \39865 , \39866 , \39867 , \39868 , \39869 , \39870 , \39871 , \39872 , \39873 , \39874 ,
         \39875 , \39876 , \39877 , \39878 , \39879 , \39880 , \39881 , \39882 , \39883 , \39884 ,
         \39885 , \39886 , \39887 , \39888 , \39889 , \39890 , \39891 , \39892 , \39893 , \39894 ,
         \39895 , \39896 , \39897 , \39898 , \39899 , \39900 , \39901 , \39902 , \39903 , \39904 ,
         \39905 , \39906 , \39907 , \39908 , \39909 , \39910 , \39911 , \39912 , \39913 , \39914 ,
         \39915 , \39916 , \39917 , \39918 , \39919 , \39920 , \39921 , \39922 , \39923 , \39924 ,
         \39925 , \39926 , \39927 , \39928 , \39929 , \39930 , \39931 , \39932 , \39933 , \39934 ,
         \39935 , \39936 , \39937 , \39938 , \39939 , \39940 , \39941 , \39942 , \39943 , \39944 ,
         \39945 , \39946 , \39947 , \39948 , \39949 , \39950 , \39951 , \39952 , \39953 , \39954 ,
         \39955 , \39956 , \39957 , \39958 , \39959 , \39960 , \39961 , \39962 , \39963 , \39964 ,
         \39965 , \39966 , \39967 , \39968 , \39969 , \39970 , \39971 , \39972 , \39973 , \39974 ,
         \39975 , \39976 , \39977 , \39978 , \39979 , \39980 , \39981 , \39982 , \39983 , \39984 ,
         \39985 , \39986 , \39987 , \39988 , \39989 , \39990 , \39991 , \39992 , \39993 , \39994 ,
         \39995 , \39996 , \39997 , \39998 , \39999 , \40000 , \40001 , \40002 , \40003 , \40004 ,
         \40005 , \40006 , \40007 , \40008 , \40009 , \40010 , \40011 , \40012 , \40013 , \40014 ,
         \40015 , \40016 , \40017 , \40018 , \40019 , \40020 , \40021 , \40022 , \40023 , \40024 ,
         \40025 , \40026 , \40027 , \40028 , \40029 , \40030 , \40031 , \40032 , \40033 , \40034 ,
         \40035 , \40036 , \40037 , \40038 , \40039 , \40040 , \40041 , \40042 , \40043 , \40044 ,
         \40045 , \40046 , \40047 , \40048 , \40049 , \40050 , \40051 , \40052 , \40053 , \40054 ,
         \40055 , \40056 , \40057 , \40058 , \40059 , \40060 , \40061 , \40062 , \40063 , \40064 ,
         \40065 , \40066 , \40067 , \40068 , \40069 , \40070 , \40071 , \40072 , \40073 , \40074 ,
         \40075 , \40076 , \40077 , \40078 , \40079 , \40080 , \40081 , \40082 , \40083 , \40084 ,
         \40085 , \40086 , \40087 , \40088 , \40089 , \40090 , \40091 , \40092 , \40093 , \40094 ,
         \40095 , \40096 , \40097 , \40098 , \40099 , \40100 , \40101 , \40102 , \40103 , \40104 ,
         \40105 , \40106 , \40107 , \40108 , \40109 , \40110 , \40111 , \40112 , \40113 , \40114 ,
         \40115 , \40116 , \40117 , \40118 , \40119 , \40120 , \40121 , \40122 , \40123 , \40124 ,
         \40125 , \40126 , \40127 , \40128 , \40129 , \40130 , \40131 , \40132 , \40133 , \40134 ,
         \40135 , \40136 , \40137 , \40138 , \40139 , \40140 , \40141 , \40142 , \40143 , \40144 ,
         \40145 , \40146 , \40147 , \40148 , \40149 , \40150 , \40151 , \40152 , \40153 , \40154 ,
         \40155 , \40156 , \40157 , \40158 , \40159 , \40160 , \40161 , \40162 , \40163 , \40164 ,
         \40165 , \40166 , \40167 , \40168 , \40169 , \40170 , \40171 , \40172 , \40173 , \40174 ,
         \40175 , \40176 , \40177 , \40178 , \40179 , \40180 , \40181 , \40182 , \40183 , \40184 ,
         \40185 , \40186 , \40187 , \40188 , \40189 , \40190 , \40191 , \40192 , \40193 , \40194 ,
         \40195 , \40196 , \40197 , \40198 , \40199 , \40200 , \40201 , \40202 , \40203 , \40204 ,
         \40205 , \40206 , \40207 , \40208 , \40209 , \40210 , \40211 , \40212 , \40213 , \40214 ,
         \40215 , \40216 , \40217 , \40218 , \40219 , \40220 , \40221 , \40222 , \40223 , \40224 ,
         \40225 , \40226 , \40227 , \40228 , \40229 , \40230 , \40231 , \40232 , \40233 , \40234 ,
         \40235 , \40236 , \40237 , \40238 , \40239 , \40240 , \40241 , \40242 , \40243 , \40244 ,
         \40245 , \40246 , \40247 , \40248 , \40249 , \40250 , \40251 , \40252 , \40253 , \40254 ,
         \40255 , \40256 , \40257 , \40258 , \40259 , \40260 , \40261 , \40262 , \40263 , \40264 ,
         \40265 , \40266 , \40267 , \40268 , \40269 , \40270 , \40271 , \40272 , \40273 , \40274 ,
         \40275 , \40276 , \40277 , \40278 , \40279 , \40280 , \40281 , \40282 , \40283 , \40284 ,
         \40285 , \40286 , \40287 , \40288 , \40289 , \40290 , \40291 , \40292 , \40293 , \40294 ,
         \40295 , \40296 , \40297 , \40298 , \40299 , \40300 , \40301 , \40302 , \40303 , \40304 ,
         \40305 , \40306 , \40307 , \40308 , \40309 , \40310 , \40311 , \40312 , \40313 , \40314 ,
         \40315 , \40316 , \40317 , \40318 , \40319 , \40320 , \40321 , \40322 , \40323 , \40324 ,
         \40325 , \40326 , \40327 , \40328 , \40329 , \40330 , \40331 , \40332 , \40333 , \40334 ,
         \40335 , \40336 , \40337 , \40338 , \40339 , \40340 , \40341 , \40342 , \40343 , \40344 ,
         \40345 , \40346 , \40347 , \40348 , \40349 , \40350 , \40351 , \40352 , \40353 , \40354 ,
         \40355 , \40356 , \40357 , \40358 , \40359 , \40360 , \40361 , \40362 , \40363 , \40364 ,
         \40365 , \40366 , \40367 , \40368 , \40369 , \40370 , \40371 , \40372 , \40373 , \40374 ,
         \40375 , \40376 , \40377 , \40378 , \40379 , \40380 , \40381 , \40382 , \40383 , \40384 ,
         \40385 , \40386 , \40387 , \40388 , \40389 , \40390 , \40391 , \40392 , \40393 , \40394 ,
         \40395 , \40396 , \40397 , \40398 , \40399 , \40400 , \40401 , \40402 , \40403 , \40404 ,
         \40405 , \40406 , \40407 , \40408 , \40409 , \40410 , \40411 , \40412 , \40413 , \40414 ,
         \40415 , \40416 , \40417 , \40418 , \40419 , \40420 , \40421 , \40422 , \40423 , \40424 ,
         \40425 , \40426 , \40427 , \40428 , \40429 , \40430 , \40431 , \40432 , \40433 , \40434 ,
         \40435 , \40436 , \40437 , \40438 , \40439 , \40440 , \40441 , \40442 , \40443 , \40444 ,
         \40445 , \40446 , \40447 , \40448 , \40449 , \40450 , \40451 , \40452 , \40453 , \40454 ,
         \40455 , \40456 , \40457 , \40458 , \40459 , \40460 , \40461 , \40462 , \40463 , \40464 ,
         \40465 , \40466 , \40467 , \40468 , \40469 , \40470 , \40471 , \40472 , \40473 , \40474 ,
         \40475 , \40476 , \40477 , \40478 , \40479 , \40480 , \40481 , \40482 , \40483 , \40484 ,
         \40485 , \40486 , \40487 , \40488 , \40489 , \40490 , \40491 , \40492 , \40493 , \40494 ,
         \40495 , \40496 , \40497 , \40498 , \40499 , \40500 , \40501 , \40502 , \40503 , \40504 ,
         \40505 , \40506 , \40507 , \40508 , \40509 , \40510 , \40511 , \40512 , \40513 , \40514 ,
         \40515 , \40516 , \40517 , \40518 , \40519 , \40520 , \40521 , \40522 , \40523 , \40524 ,
         \40525 , \40526 , \40527 , \40528 , \40529 , \40530 , \40531 , \40532 , \40533 , \40534 ,
         \40535 , \40536 , \40537 , \40538 , \40539 , \40540 , \40541 , \40542 , \40543 , \40544 ,
         \40545 , \40546 , \40547 , \40548 , \40549 , \40550 , \40551 , \40552 , \40553 , \40554 ,
         \40555 , \40556 , \40557 , \40558 , \40559 , \40560 , \40561 , \40562 , \40563 , \40564 ,
         \40565 , \40566 , \40567 , \40568 , \40569 , \40570 , \40571 , \40572 , \40573 , \40574 ,
         \40575 , \40576 , \40577 , \40578 , \40579 , \40580 , \40581 , \40582 , \40583 , \40584 ,
         \40585 , \40586 , \40587 , \40588 , \40589 , \40590 , \40591 , \40592 , \40593 , \40594 ,
         \40595 , \40596 , \40597 , \40598 , \40599 , \40600 , \40601 , \40602 , \40603 , \40604 ,
         \40605 , \40606 , \40607 , \40608 , \40609 , \40610 , \40611 , \40612 , \40613 , \40614 ,
         \40615 , \40616 , \40617 , \40618 , \40619 , \40620 , \40621 , \40622 , \40623 , \40624 ,
         \40625 , \40626 , \40627 , \40628 , \40629 , \40630 , \40631 , \40632 , \40633 , \40634 ,
         \40635 , \40636 , \40637 , \40638 , \40639 , \40640 , \40641 , \40642 , \40643 , \40644 ,
         \40645 , \40646 , \40647 , \40648 , \40649 , \40650 , \40651 , \40652 , \40653 , \40654 ,
         \40655 , \40656 , \40657 , \40658 , \40659 , \40660 , \40661 , \40662 , \40663 , \40664 ,
         \40665 , \40666 , \40667 , \40668 , \40669 , \40670 , \40671 , \40672 , \40673 , \40674 ,
         \40675 , \40676 , \40677 , \40678 , \40679 , \40680 , \40681 , \40682 , \40683 , \40684 ,
         \40685 , \40686 , \40687 , \40688 , \40689 , \40690 , \40691 , \40692 , \40693 , \40694 ,
         \40695 , \40696 , \40697 , \40698 , \40699 , \40700 , \40701 , \40702 , \40703 , \40704 ,
         \40705 , \40706 , \40707 , \40708 , \40709 , \40710 , \40711 , \40712 , \40713 , \40714 ,
         \40715 , \40716 , \40717 , \40718 , \40719 , \40720 , \40721 , \40722 , \40723 , \40724 ,
         \40725 , \40726 , \40727 , \40728 , \40729 , \40730 , \40731 , \40732 , \40733 , \40734 ,
         \40735 , \40736 , \40737 , \40738 , \40739 , \40740 , \40741 , \40742 , \40743 , \40744 ,
         \40745 , \40746 , \40747 , \40748 , \40749 , \40750 , \40751 , \40752 , \40753 , \40754 ,
         \40755 , \40756 , \40757 , \40758 , \40759 , \40760 , \40761 , \40762 , \40763 , \40764 ,
         \40765 , \40766 , \40767 , \40768 , \40769 , \40770 , \40771 , \40772 , \40773 , \40774 ,
         \40775 , \40776 , \40777 , \40778 , \40779 , \40780 , \40781 , \40782 , \40783 , \40784 ,
         \40785 , \40786 , \40787 , \40788 , \40789 , \40790 , \40791 , \40792 , \40793 , \40794 ,
         \40795 , \40796 , \40797 , \40798 , \40799 , \40800 , \40801 , \40802 , \40803 , \40804 ,
         \40805 , \40806 , \40807 , \40808 , \40809 , \40810 , \40811 , \40812 , \40813 , \40814 ,
         \40815 , \40816 , \40817 , \40818 , \40819 , \40820 , \40821 , \40822 , \40823 , \40824 ,
         \40825 , \40826 , \40827 , \40828 , \40829 , \40830 , \40831 , \40832 , \40833 , \40834 ,
         \40835 , \40836 , \40837 , \40838 , \40839 , \40840 , \40841 , \40842 , \40843 , \40844 ,
         \40845 , \40846 , \40847 , \40848 , \40849 , \40850 , \40851 , \40852 , \40853 , \40854 ,
         \40855 , \40856 , \40857 , \40858 , \40859 , \40860 , \40861 , \40862 , \40863 , \40864 ,
         \40865 , \40866 , \40867 , \40868 , \40869 , \40870 , \40871 , \40872 , \40873 , \40874 ,
         \40875 , \40876 , \40877 , \40878 , \40879 , \40880 , \40881 , \40882 , \40883 , \40884 ,
         \40885 , \40886 , \40887 , \40888 , \40889 , \40890 , \40891 , \40892 , \40893 , \40894 ,
         \40895 , \40896 , \40897 , \40898 , \40899 , \40900 , \40901 , \40902 , \40903 , \40904 ,
         \40905 , \40906 , \40907 , \40908 , \40909 , \40910 , \40911 , \40912 , \40913 , \40914 ,
         \40915 , \40916 , \40917 , \40918 , \40919 , \40920 , \40921 , \40922 , \40923 , \40924 ,
         \40925 , \40926 , \40927 , \40928 , \40929 , \40930 , \40931 , \40932 , \40933 , \40934 ,
         \40935 , \40936 , \40937 , \40938 , \40939 , \40940 , \40941 , \40942 , \40943 , \40944 ,
         \40945 , \40946 , \40947 , \40948 , \40949 , \40950 , \40951 , \40952 , \40953 , \40954 ,
         \40955 , \40956 , \40957 , \40958 , \40959 , \40960 , \40961 , \40962 , \40963 , \40964 ,
         \40965 , \40966 , \40967 , \40968 , \40969 , \40970 , \40971 , \40972 , \40973 , \40974 ,
         \40975 , \40976 , \40977 , \40978 , \40979 , \40980 , \40981 , \40982 , \40983 , \40984 ,
         \40985 , \40986 , \40987 , \40988 , \40989 , \40990 , \40991 , \40992 , \40993 , \40994 ,
         \40995 , \40996 , \40997 , \40998 , \40999 , \41000 , \41001 , \41002 , \41003 , \41004 ,
         \41005 , \41006 , \41007 , \41008 , \41009 , \41010 , \41011 , \41012 , \41013 , \41014 ,
         \41015 , \41016 , \41017 , \41018 , \41019 , \41020 , \41021 , \41022 , \41023 , \41024 ,
         \41025 , \41026 , \41027 , \41028 , \41029 , \41030 , \41031 , \41032 , \41033 , \41034 ,
         \41035 , \41036 , \41037 , \41038 , \41039 , \41040 , \41041 , \41042 , \41043 , \41044 ,
         \41045 , \41046 , \41047 , \41048 , \41049 , \41050 , \41051 , \41052 , \41053 , \41054 ,
         \41055 , \41056 , \41057 , \41058 , \41059 , \41060 , \41061 , \41062 , \41063 , \41064 ,
         \41065 , \41066 , \41067 , \41068 , \41069 , \41070 , \41071 , \41072 , \41073 , \41074 ,
         \41075 , \41076 , \41077 , \41078 , \41079 , \41080 , \41081 , \41082 , \41083 , \41084 ,
         \41085 , \41086 , \41087 , \41088 , \41089 , \41090 , \41091 , \41092 , \41093 , \41094 ,
         \41095 , \41096 , \41097 , \41098 , \41099 , \41100 , \41101 , \41102 , \41103 , \41104 ,
         \41105 , \41106 , \41107 , \41108 , \41109 , \41110 , \41111 , \41112 , \41113 , \41114 ,
         \41115 , \41116 , \41117 , \41118 , \41119 , \41120 , \41121 , \41122 , \41123 , \41124 ,
         \41125 , \41126 , \41127 , \41128 , \41129 , \41130 , \41131 , \41132 , \41133 , \41134 ,
         \41135 , \41136 , \41137 , \41138 , \41139 , \41140 , \41141 , \41142 , \41143 , \41144 ,
         \41145 , \41146 , \41147 , \41148 , \41149 , \41150 , \41151 , \41152 , \41153 , \41154 ,
         \41155 , \41156 , \41157 , \41158 , \41159 , \41160 , \41161 , \41162 , \41163 , \41164 ,
         \41165 , \41166 , \41167 , \41168 , \41169 , \41170 , \41171 , \41172 , \41173 , \41174 ,
         \41175 , \41176 , \41177 , \41178 , \41179 , \41180 , \41181 , \41182 , \41183 , \41184 ,
         \41185 , \41186 , \41187 , \41188 , \41189 , \41190 , \41191 , \41192 , \41193 , \41194 ,
         \41195 , \41196 , \41197 , \41198 , \41199 , \41200 , \41201 , \41202 , \41203 , \41204 ,
         \41205 , \41206 , \41207 , \41208 , \41209 , \41210 , \41211 , \41212 , \41213 , \41214 ,
         \41215 , \41216 , \41217 , \41218 , \41219 , \41220 , \41221 , \41222 , \41223 , \41224 ,
         \41225 , \41226 , \41227 , \41228 , \41229 , \41230 , \41231 , \41232 , \41233 , \41234 ,
         \41235 , \41236 , \41237 , \41238 , \41239 , \41240 , \41241 , \41242 , \41243 , \41244 ,
         \41245 , \41246 , \41247 , \41248 , \41249 , \41250 , \41251 , \41252 , \41253 , \41254 ,
         \41255 , \41256 , \41257 , \41258 , \41259 , \41260 , \41261 , \41262 , \41263 , \41264 ,
         \41265 , \41266 , \41267 , \41268 , \41269 , \41270 , \41271 , \41272 , \41273 , \41274 ,
         \41275 , \41276 , \41277 , \41278 , \41279 , \41280 , \41281 , \41282 , \41283 , \41284 ,
         \41285 , \41286 , \41287 , \41288 , \41289 , \41290 , \41291 , \41292 , \41293 , \41294 ,
         \41295 , \41296 , \41297 , \41298 , \41299 , \41300 , \41301 , \41302 , \41303 , \41304 ,
         \41305 , \41306 , \41307 , \41308 , \41309 , \41310 , \41311 , \41312 , \41313 , \41314 ,
         \41315 , \41316 , \41317 , \41318 , \41319 , \41320 , \41321 , \41322 , \41323 , \41324 ,
         \41325 , \41326 , \41327 , \41328 , \41329 , \41330 , \41331 , \41332 , \41333 , \41334 ,
         \41335 , \41336 , \41337 , \41338 , \41339 , \41340 , \41341 , \41342 , \41343 , \41344 ,
         \41345 , \41346 , \41347 , \41348 , \41349 , \41350 , \41351 , \41352 , \41353 , \41354 ,
         \41355 , \41356 , \41357 , \41358 , \41359 , \41360 , \41361 , \41362 , \41363 , \41364 ,
         \41365 , \41366 , \41367 , \41368 , \41369 , \41370 , \41371 , \41372 , \41373 , \41374 ,
         \41375 , \41376 , \41377 , \41378 , \41379 , \41380 , \41381 , \41382 , \41383 , \41384 ,
         \41385 , \41386 , \41387 , \41388 , \41389 , \41390 , \41391 , \41392 , \41393 , \41394 ,
         \41395 , \41396 , \41397 , \41398 , \41399 , \41400 , \41401 , \41402 , \41403 , \41404 ,
         \41405 , \41406 , \41407 , \41408 , \41409 , \41410 , \41411 , \41412 , \41413 , \41414 ,
         \41415 , \41416 , \41417 , \41418 , \41419 , \41420 , \41421 , \41422 , \41423 , \41424 ,
         \41425 , \41426 , \41427 , \41428 , \41429 , \41430 , \41431 , \41432 , \41433 , \41434 ,
         \41435 , \41436 , \41437 , \41438 , \41439 , \41440 , \41441 , \41442 , \41443 , \41444 ,
         \41445 , \41446 , \41447 , \41448 , \41449 , \41450 , \41451 , \41452 , \41453 , \41454 ,
         \41455 , \41456 , \41457 , \41458 , \41459 , \41460 , \41461 , \41462 , \41463 , \41464 ,
         \41465 , \41466 , \41467 , \41468 , \41469 , \41470 , \41471 , \41472 , \41473 , \41474 ,
         \41475 , \41476 , \41477 , \41478 , \41479 , \41480 , \41481 , \41482 , \41483 , \41484 ,
         \41485 , \41486 , \41487 , \41488 , \41489 , \41490 , \41491 , \41492 , \41493 , \41494 ,
         \41495 , \41496 , \41497 , \41498 , \41499 , \41500 , \41501 , \41502 , \41503 , \41504 ,
         \41505 , \41506 , \41507 , \41508 , \41509 , \41510 , \41511 , \41512 , \41513 , \41514 ,
         \41515 , \41516 , \41517 , \41518 , \41519 , \41520 , \41521 , \41522 , \41523 , \41524 ,
         \41525 , \41526 , \41527 , \41528 , \41529 , \41530 , \41531 , \41532 , \41533 , \41534 ,
         \41535 , \41536 , \41537 , \41538 , \41539 , \41540 , \41541 , \41542 , \41543 , \41544 ,
         \41545 , \41546 , \41547 , \41548 , \41549 , \41550 , \41551 , \41552 , \41553 , \41554 ,
         \41555 , \41556 , \41557 , \41558 , \41559 , \41560 , \41561 , \41562 , \41563 , \41564 ,
         \41565 , \41566 , \41567 , \41568 , \41569 , \41570 , \41571 , \41572 , \41573 , \41574 ,
         \41575 , \41576 , \41577 , \41578 , \41579 , \41580 , \41581 , \41582 , \41583 , \41584 ,
         \41585 , \41586 , \41587 , \41588 , \41589 , \41590 , \41591 , \41592 , \41593 , \41594 ,
         \41595 , \41596 , \41597 , \41598 , \41599 , \41600 , \41601 , \41602 , \41603 , \41604 ,
         \41605 , \41606 , \41607 , \41608 , \41609 , \41610 , \41611 , \41612 , \41613 , \41614 ,
         \41615 , \41616 , \41617 , \41618 , \41619 , \41620 , \41621 , \41622 , \41623 , \41624 ,
         \41625 , \41626 , \41627 , \41628 , \41629 , \41630 , \41631 , \41632 , \41633 , \41634 ,
         \41635 , \41636 , \41637 , \41638 , \41639 , \41640 , \41641 , \41642 , \41643 , \41644 ,
         \41645 , \41646 , \41647 , \41648 , \41649 , \41650 , \41651 , \41652 , \41653 , \41654 ,
         \41655 , \41656 , \41657 , \41658 , \41659 , \41660 , \41661 , \41662 , \41663 , \41664 ,
         \41665 , \41666 , \41667 , \41668 , \41669 , \41670 , \41671 , \41672 , \41673 , \41674 ,
         \41675 , \41676 , \41677 , \41678 , \41679 , \41680 , \41681 , \41682 , \41683 , \41684 ,
         \41685 , \41686 , \41687 , \41688 , \41689 , \41690 , \41691 , \41692 , \41693 , \41694 ,
         \41695 , \41696 , \41697 , \41698 , \41699 , \41700 , \41701 , \41702 , \41703 , \41704 ,
         \41705 , \41706 , \41707 , \41708 , \41709 , \41710 , \41711 , \41712 , \41713 , \41714 ,
         \41715 , \41716 , \41717 , \41718 , \41719 , \41720 , \41721 , \41722 , \41723 , \41724 ,
         \41725 , \41726 , \41727 , \41728 , \41729 , \41730 , \41731 , \41732 , \41733 , \41734 ,
         \41735 , \41736 , \41737 , \41738 , \41739 , \41740 , \41741 , \41742 , \41743 , \41744 ,
         \41745 , \41746 , \41747 , \41748 , \41749 , \41750 , \41751 , \41752 , \41753 , \41754 ,
         \41755 , \41756 , \41757 , \41758 , \41759 , \41760 , \41761 , \41762 , \41763 , \41764 ,
         \41765 , \41766 , \41767 , \41768 , \41769 , \41770 , \41771 , \41772 , \41773 , \41774 ,
         \41775 , \41776 , \41777 , \41778 , \41779 , \41780 , \41781 , \41782 , \41783 , \41784 ,
         \41785 , \41786 , \41787 , \41788 , \41789 , \41790 , \41791 , \41792 , \41793 , \41794 ,
         \41795 , \41796 , \41797 , \41798 , \41799 , \41800 , \41801 , \41802 , \41803 , \41804 ,
         \41805 , \41806 , \41807 , \41808 , \41809 , \41810 , \41811 , \41812 , \41813 , \41814 ,
         \41815 , \41816 , \41817 , \41818 , \41819 , \41820 , \41821 , \41822 , \41823 , \41824 ,
         \41825 , \41826 , \41827 , \41828 , \41829 , \41830 , \41831 , \41832 , \41833 , \41834 ,
         \41835 , \41836 , \41837 , \41838 , \41839 , \41840 , \41841 , \41842 , \41843 , \41844 ,
         \41845 , \41846 , \41847 , \41848 , \41849 , \41850 , \41851 , \41852 , \41853 , \41854 ,
         \41855 , \41856 , \41857 , \41858 , \41859 , \41860 , \41861 , \41862 , \41863 , \41864 ,
         \41865 , \41866 , \41867 , \41868 , \41869 , \41870 , \41871 , \41872 , \41873 , \41874 ,
         \41875 , \41876 , \41877 , \41878 , \41879 , \41880 , \41881 , \41882 , \41883 , \41884 ,
         \41885 , \41886 , \41887 , \41888 , \41889 , \41890 , \41891 , \41892 , \41893 , \41894 ,
         \41895 , \41896 , \41897 , \41898 , \41899 , \41900 , \41901 , \41902 , \41903 , \41904 ,
         \41905 , \41906 , \41907 , \41908 , \41909 , \41910 , \41911 , \41912 , \41913 , \41914 ,
         \41915 , \41916 , \41917 , \41918 , \41919 , \41920 , \41921 , \41922 , \41923 , \41924 ,
         \41925 , \41926 , \41927 , \41928 , \41929 , \41930 , \41931 , \41932 , \41933 , \41934 ,
         \41935 , \41936 , \41937 , \41938 , \41939 , \41940 , \41941 , \41942 , \41943 , \41944 ,
         \41945 , \41946 , \41947 , \41948 , \41949 , \41950 , \41951 , \41952 , \41953 , \41954 ,
         \41955 , \41956 , \41957 , \41958 , \41959 , \41960 , \41961 , \41962 , \41963 , \41964 ,
         \41965 , \41966 , \41967 , \41968 , \41969 , \41970 , \41971 , \41972 , \41973 , \41974 ,
         \41975 , \41976 , \41977 , \41978 , \41979 , \41980 , \41981 , \41982 , \41983 , \41984 ,
         \41985 , \41986 , \41987 , \41988 , \41989 , \41990 , \41991 , \41992 , \41993 , \41994 ,
         \41995 , \41996 , \41997 , \41998 , \41999 , \42000 , \42001 , \42002 , \42003 , \42004 ,
         \42005 , \42006 , \42007 , \42008 , \42009 , \42010 , \42011 , \42012 , \42013 , \42014 ,
         \42015 , \42016 , \42017 , \42018 , \42019 , \42020 , \42021 , \42022 , \42023 , \42024 ,
         \42025 , \42026 , \42027 , \42028 , \42029 , \42030 , \42031 , \42032 , \42033 , \42034 ,
         \42035 , \42036 , \42037 , \42038 , \42039 , \42040 , \42041 , \42042 , \42043 , \42044 ,
         \42045 , \42046 , \42047 , \42048 , \42049 , \42050 , \42051 , \42052 , \42053 , \42054 ,
         \42055 , \42056 , \42057 , \42058 , \42059 , \42060 , \42061 , \42062 , \42063 , \42064 ,
         \42065 , \42066 , \42067 , \42068 , \42069 , \42070 , \42071 , \42072 , \42073 , \42074 ,
         \42075 , \42076 , \42077 , \42078 , \42079 , \42080 , \42081 , \42082 , \42083 , \42084 ,
         \42085 , \42086 , \42087 , \42088 , \42089 , \42090 , \42091 , \42092 , \42093 , \42094 ,
         \42095 , \42096 , \42097 , \42098 , \42099 , \42100 , \42101 , \42102 , \42103 , \42104 ,
         \42105 , \42106 , \42107 , \42108 , \42109 , \42110 , \42111 , \42112 , \42113 , \42114 ,
         \42115 , \42116 , \42117 , \42118 , \42119 , \42120 , \42121 , \42122 , \42123 , \42124 ,
         \42125 , \42126 , \42127 , \42128 , \42129 , \42130 , \42131 , \42132 , \42133 , \42134 ,
         \42135 , \42136 , \42137 , \42138 , \42139 , \42140 , \42141 , \42142 , \42143 , \42144 ,
         \42145 , \42146 , \42147 , \42148 , \42149 , \42150 , \42151 , \42152 , \42153 , \42154 ,
         \42155 , \42156 , \42157 , \42158 , \42159 , \42160 , \42161 , \42162 , \42163 , \42164 ,
         \42165 , \42166 , \42167 , \42168 , \42169 , \42170 , \42171 , \42172 , \42173 , \42174 ,
         \42175 , \42176 , \42177 , \42178 , \42179 , \42180 , \42181 , \42182 , \42183 , \42184 ,
         \42185 , \42186 , \42187 , \42188 , \42189 , \42190 , \42191 , \42192 , \42193 , \42194 ,
         \42195 , \42196 , \42197 , \42198 , \42199 , \42200 , \42201 , \42202 , \42203 , \42204 ,
         \42205 , \42206 , \42207 , \42208 , \42209 , \42210 , \42211 , \42212 , \42213 , \42214 ,
         \42215 , \42216 , \42217 , \42218 , \42219 , \42220 , \42221 , \42222 , \42223 , \42224 ,
         \42225 , \42226 , \42227 , \42228 , \42229 , \42230 , \42231 , \42232 , \42233 , \42234 ,
         \42235 , \42236 , \42237 , \42238 , \42239 , \42240 , \42241 , \42242 , \42243 , \42244 ,
         \42245 , \42246 , \42247 , \42248 , \42249 , \42250 , \42251 , \42252 , \42253 , \42254 ,
         \42255 , \42256 , \42257 , \42258 , \42259 , \42260 , \42261 , \42262 , \42263 , \42264 ,
         \42265 , \42266 , \42267 , \42268 , \42269 , \42270 , \42271 , \42272 , \42273 , \42274 ,
         \42275 , \42276 , \42277 , \42278 , \42279 , \42280 , \42281 , \42282 , \42283 , \42284 ,
         \42285 , \42286 , \42287 , \42288 , \42289 , \42290 , \42291 , \42292 , \42293 , \42294 ,
         \42295 , \42296 , \42297 , \42298 , \42299 , \42300 , \42301 , \42302 , \42303 , \42304 ,
         \42305 , \42306 , \42307 , \42308 , \42309 , \42310 , \42311 , \42312 , \42313 , \42314 ,
         \42315 , \42316 , \42317 , \42318 , \42319 , \42320 , \42321 , \42322 , \42323 , \42324 ,
         \42325 , \42326 , \42327 , \42328 , \42329 , \42330 , \42331 , \42332 , \42333 , \42334 ,
         \42335 , \42336 , \42337 , \42338 , \42339 , \42340 , \42341 , \42342 , \42343 , \42344 ,
         \42345 , \42346 , \42347 , \42348 , \42349 , \42350 , \42351 , \42352 , \42353 , \42354 ,
         \42355 , \42356 , \42357 , \42358 , \42359 , \42360 , \42361 , \42362 , \42363 , \42364 ,
         \42365 , \42366 , \42367 , \42368 , \42369 , \42370 , \42371 , \42372 , \42373 , \42374 ,
         \42375 , \42376 , \42377 , \42378 , \42379 , \42380 , \42381 , \42382 , \42383 , \42384 ,
         \42385 , \42386 , \42387 , \42388 , \42389 , \42390 , \42391 , \42392 , \42393 , \42394 ,
         \42395 , \42396 , \42397 , \42398 , \42399 , \42400 , \42401 , \42402 , \42403 , \42404 ,
         \42405 , \42406 , \42407 , \42408 , \42409 , \42410 , \42411 , \42412 , \42413 , \42414 ,
         \42415 , \42416 , \42417 , \42418 , \42419 , \42420 , \42421 , \42422 , \42423 , \42424 ,
         \42425 , \42426 , \42427 , \42428 , \42429 , \42430 , \42431 , \42432 , \42433 , \42434 ,
         \42435 , \42436 , \42437 , \42438 , \42439 , \42440 , \42441 , \42442 , \42443 , \42444 ,
         \42445 , \42446 , \42447 , \42448 , \42449 , \42450 , \42451 , \42452 , \42453 , \42454 ,
         \42455 , \42456 , \42457 , \42458 , \42459 , \42460 , \42461 , \42462 , \42463 , \42464 ,
         \42465 , \42466 , \42467 , \42468 , \42469 , \42470 , \42471 , \42472 , \42473 , \42474 ,
         \42475 , \42476 , \42477 , \42478 , \42479 , \42480 , \42481 , \42482 , \42483 , \42484 ,
         \42485 , \42486 , \42487 , \42488 , \42489 , \42490 , \42491 , \42492 , \42493 , \42494 ,
         \42495 , \42496 , \42497 , \42498 , \42499 , \42500 , \42501 , \42502 , \42503 , \42504 ,
         \42505 , \42506 , \42507 , \42508 , \42509 , \42510 , \42511 , \42512 , \42513 , \42514 ,
         \42515 , \42516 , \42517 , \42518 , \42519 , \42520 , \42521 , \42522 , \42523 , \42524 ,
         \42525 , \42526 , \42527 , \42528 , \42529 , \42530 , \42531 , \42532 , \42533 , \42534 ,
         \42535 , \42536 , \42537 , \42538 , \42539 , \42540 , \42541 , \42542 , \42543 , \42544 ,
         \42545 , \42546 , \42547 , \42548 , \42549 , \42550 , \42551 , \42552 , \42553 , \42554 ,
         \42555 , \42556 , \42557 , \42558 , \42559 , \42560 , \42561 , \42562 , \42563 , \42564 ,
         \42565 , \42566 , \42567 , \42568 , \42569 , \42570 , \42571 , \42572 , \42573 , \42574 ,
         \42575 , \42576 , \42577 , \42578 , \42579 , \42580 , \42581 , \42582 , \42583 , \42584 ,
         \42585 , \42586 , \42587 , \42588 , \42589 , \42590 , \42591 , \42592 , \42593 , \42594 ,
         \42595 , \42596 , \42597 , \42598 , \42599 , \42600 , \42601 , \42602 , \42603 , \42604 ,
         \42605 , \42606 , \42607 , \42608 , \42609 , \42610 , \42611 , \42612 , \42613 , \42614 ,
         \42615 , \42616 , \42617 , \42618 , \42619 , \42620 , \42621 , \42622 , \42623 , \42624 ,
         \42625 , \42626 , \42627 , \42628 , \42629 , \42630 , \42631 , \42632 , \42633 , \42634 ,
         \42635 , \42636 , \42637 , \42638 , \42639 , \42640 , \42641 , \42642 , \42643 , \42644 ,
         \42645 , \42646 , \42647 , \42648 , \42649 , \42650 , \42651 , \42652 , \42653 , \42654 ,
         \42655 , \42656 , \42657 , \42658 , \42659 , \42660 , \42661 , \42662 , \42663 , \42664 ,
         \42665 , \42666 , \42667 , \42668 , \42669 , \42670 , \42671 , \42672 , \42673 , \42674 ,
         \42675 , \42676 , \42677 , \42678 , \42679 , \42680 , \42681 , \42682 , \42683 , \42684 ,
         \42685 , \42686 , \42687 , \42688 , \42689 , \42690 , \42691 , \42692 , \42693 , \42694 ,
         \42695 , \42696 , \42697 , \42698 , \42699 , \42700 , \42701 , \42702 , \42703 , \42704 ,
         \42705 , \42706 , \42707 , \42708 , \42709 , \42710 , \42711 , \42712 , \42713 , \42714 ,
         \42715 , \42716 , \42717 , \42718 , \42719 , \42720 , \42721 , \42722 , \42723 , \42724 ,
         \42725 , \42726 , \42727 , \42728 , \42729 , \42730 , \42731 , \42732 , \42733 , \42734 ,
         \42735 , \42736 , \42737 , \42738 , \42739 , \42740 , \42741 , \42742 , \42743 , \42744 ,
         \42745 , \42746 , \42747 , \42748 , \42749 , \42750 , \42751 , \42752 , \42753 , \42754 ,
         \42755 , \42756 , \42757 , \42758 , \42759 , \42760 , \42761 , \42762 , \42763 , \42764 ,
         \42765 , \42766 , \42767 , \42768 , \42769 , \42770 , \42771 , \42772 , \42773 , \42774 ,
         \42775 , \42776 , \42777 , \42778 , \42779 , \42780 , \42781 , \42782 , \42783 , \42784 ,
         \42785 , \42786 , \42787 , \42788 , \42789 , \42790 , \42791 , \42792 , \42793 , \42794 ,
         \42795 , \42796 , \42797 , \42798 , \42799 , \42800 , \42801 , \42802 , \42803 , \42804 ,
         \42805 , \42806 , \42807 , \42808 , \42809 , \42810 , \42811 , \42812 , \42813 , \42814 ,
         \42815 , \42816 , \42817 , \42818 , \42819 , \42820 , \42821 , \42822 , \42823 , \42824 ,
         \42825 , \42826 , \42827 , \42828 , \42829 , \42830 , \42831 , \42832 , \42833 , \42834 ,
         \42835 , \42836 , \42837 , \42838 , \42839 , \42840 , \42841 , \42842 , \42843 , \42844 ,
         \42845 , \42846 , \42847 , \42848 , \42849 , \42850 , \42851 , \42852 , \42853 , \42854 ,
         \42855 , \42856 , \42857 , \42858 , \42859 , \42860 , \42861 , \42862 , \42863 , \42864 ,
         \42865 , \42866 , \42867 , \42868 , \42869 , \42870 , \42871 , \42872 , \42873 , \42874 ,
         \42875 , \42876 , \42877 , \42878 , \42879 , \42880 , \42881 , \42882 , \42883 , \42884 ,
         \42885 , \42886 , \42887 , \42888 , \42889 , \42890 , \42891 , \42892 , \42893 , \42894 ,
         \42895 , \42896 , \42897 , \42898 , \42899 , \42900 , \42901 , \42902 , \42903 , \42904 ,
         \42905 , \42906 , \42907 , \42908 , \42909 , \42910 , \42911 , \42912 , \42913 , \42914 ,
         \42915 , \42916 , \42917 , \42918 , \42919 , \42920 , \42921 , \42922 , \42923 , \42924 ,
         \42925 , \42926 , \42927 , \42928 , \42929 , \42930 , \42931 , \42932 , \42933 , \42934 ,
         \42935 , \42936 , \42937 , \42938 , \42939 , \42940 , \42941 , \42942 , \42943 , \42944 ,
         \42945 , \42946 , \42947 , \42948 , \42949 , \42950 , \42951 , \42952 , \42953 , \42954 ,
         \42955 , \42956 , \42957 , \42958 , \42959 , \42960 , \42961 , \42962 , \42963 , \42964 ,
         \42965 , \42966 , \42967 , \42968 , \42969 , \42970 , \42971 , \42972 , \42973 , \42974 ,
         \42975 , \42976 , \42977 , \42978 , \42979 , \42980 , \42981 , \42982 , \42983 , \42984 ,
         \42985 , \42986 , \42987 , \42988 , \42989 , \42990 , \42991 , \42992 , \42993 , \42994 ,
         \42995 , \42996 , \42997 , \42998 , \42999 , \43000 , \43001 , \43002 , \43003 , \43004 ,
         \43005 , \43006 , \43007 , \43008 , \43009 , \43010 , \43011 , \43012 , \43013 , \43014 ,
         \43015 , \43016 , \43017 , \43018 , \43019 , \43020 , \43021 , \43022 , \43023 , \43024 ,
         \43025 , \43026 , \43027 , \43028 , \43029 , \43030 , \43031 , \43032 , \43033 , \43034 ,
         \43035 , \43036 , \43037 , \43038 , \43039 , \43040 , \43041 , \43042 , \43043 , \43044 ,
         \43045 , \43046 , \43047 , \43048 , \43049 , \43050 , \43051 , \43052 , \43053 , \43054 ,
         \43055 , \43056 , \43057 , \43058 , \43059 , \43060 , \43061 , \43062 , \43063 , \43064 ,
         \43065 , \43066 , \43067 , \43068 , \43069 , \43070 , \43071 , \43072 , \43073 , \43074 ,
         \43075 , \43076 , \43077 , \43078 , \43079 , \43080 , \43081 , \43082 , \43083 , \43084 ,
         \43085 , \43086 , \43087 , \43088 , \43089 , \43090 , \43091 , \43092 , \43093 , \43094 ,
         \43095 , \43096 , \43097 , \43098 , \43099 , \43100 , \43101 , \43102 , \43103 , \43104 ,
         \43105 , \43106 , \43107 , \43108 , \43109 , \43110 , \43111 , \43112 , \43113 , \43114 ,
         \43115 , \43116 , \43117 , \43118 , \43119 , \43120 , \43121 , \43122 , \43123 , \43124 ,
         \43125 , \43126 , \43127 , \43128 , \43129 , \43130 , \43131 , \43132 , \43133 , \43134 ,
         \43135 , \43136 , \43137 , \43138 , \43139 , \43140 , \43141 , \43142 , \43143 , \43144 ,
         \43145 , \43146 , \43147 , \43148 , \43149 , \43150 , \43151 , \43152 , \43153 , \43154 ,
         \43155 , \43156 , \43157 , \43158 , \43159 , \43160 , \43161 , \43162 , \43163 , \43164 ,
         \43165 , \43166 , \43167 , \43168 , \43169 , \43170 , \43171 , \43172 , \43173 , \43174 ,
         \43175 , \43176 , \43177 , \43178 , \43179 , \43180 , \43181 , \43182 , \43183 , \43184 ,
         \43185 , \43186 , \43187 , \43188 , \43189 , \43190 , \43191 , \43192 , \43193 , \43194 ,
         \43195 , \43196 , \43197 , \43198 , \43199 , \43200 , \43201 , \43202 , \43203 , \43204 ,
         \43205 , \43206 , \43207 , \43208 , \43209 , \43210 , \43211 , \43212 , \43213 , \43214 ,
         \43215 , \43216 , \43217 , \43218 , \43219 , \43220 , \43221 , \43222 , \43223 , \43224 ,
         \43225 , \43226 , \43227 , \43228 , \43229 , \43230 , \43231 , \43232 , \43233 , \43234 ,
         \43235 , \43236 , \43237 , \43238 , \43239 , \43240 , \43241 , \43242 , \43243 , \43244 ,
         \43245 , \43246 , \43247 , \43248 , \43249 , \43250 , \43251 , \43252 , \43253 , \43254 ,
         \43255 , \43256 , \43257 , \43258 , \43259 , \43260 , \43261 , \43262 , \43263 , \43264 ,
         \43265 , \43266 , \43267 , \43268 , \43269 , \43270 , \43271 , \43272 , \43273 , \43274 ,
         \43275 , \43276 , \43277 , \43278 , \43279 , \43280 , \43281 , \43282 , \43283 , \43284 ,
         \43285 , \43286 , \43287 , \43288 , \43289 , \43290 , \43291 , \43292 , \43293 , \43294 ,
         \43295 , \43296 , \43297 , \43298 , \43299 , \43300 , \43301 , \43302 , \43303 , \43304 ,
         \43305 , \43306 , \43307 , \43308 , \43309 , \43310 , \43311 , \43312 , \43313 , \43314 ,
         \43315 , \43316 , \43317 , \43318 , \43319 , \43320 , \43321 , \43322 , \43323 , \43324 ,
         \43325 , \43326 , \43327 , \43328 , \43329 , \43330 , \43331 , \43332 , \43333 , \43334 ,
         \43335 , \43336 , \43337 , \43338 , \43339 , \43340 , \43341 , \43342 , \43343 , \43344 ,
         \43345 , \43346 , \43347 , \43348 , \43349 , \43350 , \43351 , \43352 , \43353 , \43354 ,
         \43355 , \43356 , \43357 , \43358 , \43359 , \43360 , \43361 , \43362 , \43363 , \43364 ,
         \43365 , \43366 , \43367 , \43368 , \43369 , \43370 , \43371 , \43372 , \43373 , \43374 ,
         \43375 , \43376 , \43377 , \43378 , \43379 , \43380 , \43381 , \43382 , \43383 , \43384 ,
         \43385 , \43386 , \43387 , \43388 , \43389 , \43390 , \43391 , \43392 , \43393 , \43394 ,
         \43395 , \43396 , \43397 , \43398 , \43399 , \43400 , \43401 , \43402 , \43403 , \43404 ,
         \43405 , \43406 , \43407 , \43408 , \43409 , \43410 , \43411 , \43412 , \43413 , \43414 ,
         \43415 , \43416 , \43417 , \43418 , \43419 , \43420 , \43421 , \43422 , \43423 , \43424 ,
         \43425 , \43426 , \43427 , \43428 , \43429 , \43430 , \43431 , \43432 , \43433 , \43434 ,
         \43435 , \43436 , \43437 , \43438 , \43439 , \43440 , \43441 , \43442 , \43443 , \43444 ,
         \43445 , \43446 , \43447 , \43448 , \43449 , \43450 , \43451 , \43452 , \43453 , \43454 ,
         \43455 , \43456 , \43457 , \43458 , \43459 , \43460 , \43461 , \43462 , \43463 , \43464 ,
         \43465 , \43466 , \43467 , \43468 , \43469 , \43470 , \43471 , \43472 , \43473 , \43474 ,
         \43475 , \43476 , \43477 , \43478 , \43479 , \43480 , \43481 , \43482 , \43483 , \43484 ,
         \43485 , \43486 , \43487 , \43488 , \43489 , \43490 , \43491 , \43492 , \43493 , \43494 ,
         \43495 , \43496 , \43497 , \43498 , \43499 , \43500 , \43501 , \43502 , \43503 , \43504 ,
         \43505 , \43506 , \43507 , \43508 , \43509 , \43510 , \43511 , \43512 , \43513 , \43514 ,
         \43515 , \43516 , \43517 , \43518 , \43519 , \43520 , \43521 , \43522 , \43523 , \43524 ,
         \43525 , \43526 , \43527 , \43528 , \43529 , \43530 , \43531 , \43532 , \43533 , \43534 ,
         \43535 , \43536 , \43537 , \43538 , \43539 , \43540 , \43541 , \43542 , \43543 , \43544 ,
         \43545 , \43546 , \43547 , \43548 , \43549 , \43550 , \43551 , \43552 , \43553 , \43554 ,
         \43555 , \43556 , \43557 , \43558 , \43559 , \43560 , \43561 , \43562 , \43563 , \43564 ,
         \43565 , \43566 , \43567 , \43568 , \43569 , \43570 , \43571 , \43572 , \43573 , \43574 ,
         \43575 , \43576 , \43577 , \43578 , \43579 , \43580 , \43581 , \43582 , \43583 , \43584 ,
         \43585 , \43586 , \43587 , \43588 , \43589 , \43590 , \43591 , \43592 , \43593 , \43594 ,
         \43595 , \43596 , \43597 , \43598 , \43599 , \43600 , \43601 , \43602 , \43603 , \43604 ,
         \43605 , \43606 , \43607 , \43608 , \43609 , \43610 , \43611 , \43612 , \43613 , \43614 ,
         \43615 , \43616 , \43617 , \43618 , \43619 , \43620 , \43621 , \43622 , \43623 , \43624 ,
         \43625 , \43626 , \43627 , \43628 , \43629 , \43630 , \43631 , \43632 , \43633 , \43634 ,
         \43635 , \43636 , \43637 , \43638 , \43639 , \43640 , \43641 , \43642 , \43643 , \43644 ,
         \43645 , \43646 , \43647 , \43648 , \43649 , \43650 , \43651 , \43652 , \43653 , \43654 ,
         \43655 , \43656 , \43657 , \43658 , \43659 , \43660 , \43661 , \43662 , \43663 , \43664 ,
         \43665 , \43666 , \43667 , \43668 , \43669 , \43670 , \43671 , \43672 , \43673 , \43674 ,
         \43675 , \43676 , \43677 , \43678 , \43679 , \43680 , \43681 , \43682 , \43683 , \43684 ,
         \43685 , \43686 , \43687 , \43688 , \43689 , \43690 , \43691 , \43692 , \43693 , \43694 ,
         \43695 , \43696 , \43697 , \43698 , \43699 , \43700 , \43701 , \43702 , \43703 , \43704 ,
         \43705 , \43706 , \43707 , \43708 , \43709 , \43710 , \43711 , \43712 , \43713 , \43714 ,
         \43715 , \43716 , \43717 , \43718 , \43719 , \43720 , \43721 , \43722 , \43723 , \43724 ,
         \43725 , \43726 , \43727 , \43728 , \43729 , \43730 , \43731 , \43732 , \43733 , \43734 ,
         \43735 , \43736 , \43737 , \43738 , \43739 , \43740 , \43741 , \43742 , \43743 , \43744 ,
         \43745 , \43746 , \43747 , \43748 , \43749 , \43750 , \43751 , \43752 , \43753 , \43754 ,
         \43755 , \43756 , \43757 , \43758 , \43759 , \43760 , \43761 , \43762 , \43763 , \43764 ,
         \43765 , \43766 , \43767 , \43768 , \43769 , \43770 , \43771 , \43772 , \43773 , \43774 ,
         \43775 , \43776 , \43777 , \43778 , \43779 , \43780 , \43781 , \43782 , \43783 , \43784 ,
         \43785 , \43786 , \43787 , \43788 , \43789 , \43790 , \43791 , \43792 , \43793 , \43794 ,
         \43795 , \43796 , \43797 , \43798 , \43799 , \43800 , \43801 , \43802 , \43803 , \43804 ,
         \43805 , \43806 , \43807 , \43808 , \43809 , \43810 , \43811 , \43812 , \43813 , \43814 ,
         \43815 , \43816 , \43817 , \43818 , \43819 , \43820 , \43821 , \43822 , \43823 , \43824 ,
         \43825 , \43826 , \43827 , \43828 , \43829 , \43830 , \43831 , \43832 , \43833 , \43834 ,
         \43835 , \43836 , \43837 , \43838 , \43839 , \43840 , \43841 , \43842 , \43843 , \43844 ,
         \43845 , \43846 , \43847 , \43848 , \43849 , \43850 , \43851 , \43852 , \43853 , \43854 ,
         \43855 , \43856 , \43857 , \43858 , \43859 , \43860 , \43861 , \43862 , \43863 , \43864 ,
         \43865 , \43866 , \43867 , \43868 , \43869 , \43870 , \43871 , \43872 , \43873 , \43874 ,
         \43875 , \43876 , \43877 , \43878 , \43879 , \43880 , \43881 , \43882 , \43883 , \43884 ,
         \43885 , \43886 , \43887 , \43888 , \43889 , \43890 , \43891 , \43892 , \43893 , \43894 ,
         \43895 , \43896 , \43897 , \43898 , \43899 , \43900 , \43901 , \43902 , \43903 , \43904 ,
         \43905 , \43906 , \43907 , \43908 , \43909 , \43910 , \43911 , \43912 , \43913 , \43914 ,
         \43915 , \43916 , \43917 , \43918 , \43919 , \43920 , \43921 , \43922 , \43923 , \43924 ,
         \43925 , \43926 , \43927 , \43928 , \43929 , \43930 , \43931 , \43932 , \43933 , \43934 ,
         \43935 , \43936 , \43937 , \43938 , \43939 , \43940 , \43941 , \43942 , \43943 , \43944 ,
         \43945 , \43946 , \43947 , \43948 , \43949 , \43950 , \43951 , \43952 , \43953 , \43954 ,
         \43955 , \43956 , \43957 , \43958 , \43959 , \43960 , \43961 , \43962 , \43963 , \43964 ,
         \43965 , \43966 , \43967 , \43968 , \43969 , \43970 , \43971 , \43972 , \43973 , \43974 ,
         \43975 , \43976 , \43977 , \43978 , \43979 , \43980 , \43981 , \43982 , \43983 , \43984 ,
         \43985 , \43986 , \43987 , \43988 , \43989 , \43990 , \43991 , \43992 , \43993 , \43994 ,
         \43995 , \43996 , \43997 , \43998 , \43999 , \44000 , \44001 , \44002 , \44003 , \44004 ,
         \44005 , \44006 , \44007 , \44008 , \44009 , \44010 , \44011 , \44012 , \44013 , \44014 ,
         \44015 , \44016 , \44017 , \44018 , \44019 , \44020 , \44021 , \44022 , \44023 , \44024 ,
         \44025 , \44026 , \44027 , \44028 , \44029 , \44030 , \44031 , \44032 , \44033 , \44034 ,
         \44035 , \44036 , \44037 , \44038 , \44039 , \44040 , \44041 , \44042 , \44043 , \44044 ,
         \44045 , \44046 , \44047 , \44048 , \44049 , \44050 , \44051 , \44052 , \44053 , \44054 ,
         \44055 , \44056 , \44057 , \44058 , \44059 , \44060 , \44061 , \44062 , \44063 , \44064 ,
         \44065 , \44066 , \44067 , \44068 , \44069 , \44070 , \44071 , \44072 , \44073 , \44074 ,
         \44075 , \44076 , \44077 , \44078 , \44079 , \44080 , \44081 , \44082 , \44083 , \44084 ,
         \44085 , \44086 , \44087 , \44088 , \44089 , \44090 , \44091 , \44092 , \44093 , \44094 ,
         \44095 , \44096 , \44097 , \44098 , \44099 , \44100 , \44101 , \44102 , \44103 , \44104 ,
         \44105 , \44106 , \44107 , \44108 , \44109 , \44110 , \44111 , \44112 , \44113 , \44114 ,
         \44115 , \44116 , \44117 , \44118 , \44119 , \44120 , \44121 , \44122 , \44123 , \44124 ,
         \44125 , \44126 , \44127 , \44128 , \44129 , \44130 , \44131 , \44132 , \44133 , \44134 ,
         \44135 , \44136 , \44137 , \44138 , \44139 , \44140 , \44141 , \44142 , \44143 , \44144 ,
         \44145 , \44146 , \44147 , \44148 , \44149 , \44150 , \44151 , \44152 , \44153 , \44154 ,
         \44155 , \44156 , \44157 , \44158 , \44159 , \44160 , \44161 , \44162 , \44163 , \44164 ,
         \44165 , \44166 , \44167 , \44168 , \44169 , \44170 , \44171 , \44172 , \44173 , \44174 ,
         \44175 , \44176 , \44177 , \44178 , \44179 , \44180 , \44181 , \44182 , \44183 , \44184 ,
         \44185 , \44186 , \44187 , \44188 , \44189 , \44190 , \44191 , \44192 , \44193 , \44194 ,
         \44195 , \44196 , \44197 , \44198 , \44199 , \44200 , \44201 , \44202 , \44203 , \44204 ,
         \44205 , \44206 , \44207 , \44208 , \44209 , \44210 , \44211 , \44212 , \44213 , \44214 ,
         \44215 , \44216 , \44217 , \44218 , \44219 , \44220 , \44221 , \44222 , \44223 , \44224 ,
         \44225 , \44226 , \44227 , \44228 , \44229 , \44230 , \44231 , \44232 , \44233 , \44234 ,
         \44235 , \44236 , \44237 , \44238 , \44239 , \44240 , \44241 , \44242 , \44243 , \44244 ,
         \44245 , \44246 , \44247 , \44248 , \44249 , \44250 , \44251 , \44252 , \44253 , \44254 ,
         \44255 , \44256 , \44257 , \44258 , \44259 , \44260 , \44261 , \44262 , \44263 , \44264 ,
         \44265 , \44266 , \44267 , \44268 , \44269 , \44270 , \44271 , \44272 , \44273 , \44274 ,
         \44275 , \44276 , \44277 , \44278 , \44279 , \44280 , \44281 , \44282 , \44283 , \44284 ,
         \44285 , \44286 , \44287 , \44288 , \44289 , \44290 , \44291 , \44292 , \44293 , \44294 ,
         \44295 , \44296 , \44297 , \44298 , \44299 , \44300 , \44301 , \44302 , \44303 , \44304 ,
         \44305 , \44306 , \44307 , \44308 , \44309 , \44310 , \44311 , \44312 , \44313 , \44314 ,
         \44315 , \44316 , \44317 , \44318 , \44319 , \44320 , \44321 , \44322 , \44323 , \44324 ,
         \44325 , \44326 , \44327 , \44328 , \44329 , \44330 , \44331 , \44332 , \44333 , \44334 ,
         \44335 , \44336 , \44337 , \44338 , \44339 , \44340 , \44341 , \44342 , \44343 , \44344 ,
         \44345 , \44346 , \44347 , \44348 , \44349 , \44350 , \44351 , \44352 , \44353 , \44354 ,
         \44355 , \44356 , \44357 , \44358 , \44359 , \44360 , \44361 , \44362 , \44363 , \44364 ,
         \44365 , \44366 , \44367 , \44368 , \44369 , \44370 , \44371 , \44372 , \44373 , \44374 ,
         \44375 , \44376 , \44377 , \44378 , \44379 , \44380 , \44381 , \44382 , \44383 , \44384 ,
         \44385 , \44386 , \44387 , \44388 , \44389 , \44390 , \44391 , \44392 , \44393 , \44394 ,
         \44395 , \44396 , \44397 , \44398 , \44399 , \44400 , \44401 , \44402 , \44403 , \44404 ,
         \44405 , \44406 , \44407 , \44408 , \44409 , \44410 , \44411 , \44412 , \44413 , \44414 ,
         \44415 , \44416 , \44417 , \44418 , \44419 , \44420 , \44421 , \44422 , \44423 , \44424 ,
         \44425 , \44426 , \44427 , \44428 , \44429 , \44430 , \44431 , \44432 , \44433 , \44434 ,
         \44435 , \44436 , \44437 , \44438 , \44439 , \44440 , \44441 , \44442 , \44443 , \44444 ,
         \44445 , \44446 , \44447 , \44448 , \44449 , \44450 , \44451 , \44452 , \44453 , \44454 ,
         \44455 , \44456 , \44457 , \44458 , \44459 , \44460 , \44461 , \44462 , \44463 , \44464 ,
         \44465 , \44466 , \44467 , \44468 , \44469 , \44470 , \44471 , \44472 , \44473 , \44474 ,
         \44475 , \44476 , \44477 , \44478 , \44479 , \44480 , \44481 , \44482 , \44483 , \44484 ,
         \44485 , \44486 , \44487 , \44488 , \44489 , \44490 , \44491 , \44492 , \44493 , \44494 ,
         \44495 , \44496 , \44497 , \44498 , \44499 , \44500 , \44501 , \44502 , \44503 , \44504 ,
         \44505 , \44506 , \44507 , \44508 , \44509 , \44510 , \44511 , \44512 , \44513 , \44514 ,
         \44515 , \44516 , \44517 , \44518 , \44519 , \44520 , \44521 , \44522 , \44523 , \44524 ,
         \44525 , \44526 , \44527 , \44528 , \44529 , \44530 , \44531 , \44532 , \44533 , \44534 ,
         \44535 , \44536 , \44537 , \44538 , \44539 , \44540 , \44541 , \44542 , \44543 , \44544 ,
         \44545 , \44546 , \44547 , \44548 , \44549 , \44550 , \44551 , \44552 , \44553 , \44554 ,
         \44555 , \44556 , \44557 , \44558 , \44559 , \44560 , \44561 , \44562 , \44563 , \44564 ,
         \44565 , \44566 , \44567 , \44568 , \44569 , \44570 , \44571 , \44572 , \44573 , \44574 ,
         \44575 , \44576 , \44577 , \44578 , \44579 , \44580 , \44581 , \44582 , \44583 , \44584 ,
         \44585 , \44586 , \44587 , \44588 , \44589 , \44590 , \44591 , \44592 , \44593 , \44594 ,
         \44595 , \44596 , \44597 , \44598 , \44599 , \44600 , \44601 , \44602 , \44603 , \44604 ,
         \44605 , \44606 , \44607 , \44608 , \44609 , \44610 , \44611 , \44612 , \44613 , \44614 ,
         \44615 , \44616 , \44617 , \44618 , \44619 , \44620 , \44621 , \44622 , \44623 , \44624 ,
         \44625 , \44626 , \44627 , \44628 , \44629 , \44630 , \44631 , \44632 , \44633 , \44634 ,
         \44635 , \44636 , \44637 , \44638 , \44639 , \44640 , \44641 , \44642 , \44643 , \44644 ,
         \44645 , \44646 , \44647 , \44648 , \44649 , \44650 , \44651 , \44652 , \44653 , \44654 ,
         \44655 , \44656 , \44657 , \44658 , \44659 , \44660 , \44661 , \44662 , \44663 , \44664 ,
         \44665 , \44666 , \44667 , \44668 , \44669 , \44670 , \44671 , \44672 , \44673 , \44674 ,
         \44675 , \44676 , \44677 , \44678 , \44679 , \44680 , \44681 , \44682 , \44683 , \44684 ,
         \44685 , \44686 , \44687 , \44688 , \44689 , \44690 , \44691 , \44692 , \44693 , \44694 ,
         \44695 , \44696 , \44697 , \44698 , \44699 , \44700 , \44701 , \44702 , \44703 , \44704 ,
         \44705 , \44706 , \44707 , \44708 , \44709 , \44710 , \44711 , \44712 , \44713 , \44714 ,
         \44715 , \44716 , \44717 , \44718 , \44719 , \44720 , \44721 , \44722 , \44723 , \44724 ,
         \44725 , \44726 , \44727 , \44728 , \44729 , \44730 , \44731 , \44732 , \44733 , \44734 ,
         \44735 , \44736 , \44737 , \44738 , \44739 , \44740 , \44741 , \44742 , \44743 , \44744 ,
         \44745 , \44746 , \44747 , \44748 , \44749 , \44750 , \44751 , \44752 , \44753 , \44754 ,
         \44755 , \44756 , \44757 , \44758 , \44759 , \44760 , \44761 , \44762 , \44763 , \44764 ,
         \44765 , \44766 , \44767 , \44768 , \44769 , \44770 , \44771 , \44772 , \44773 , \44774 ,
         \44775 , \44776 , \44777 , \44778 , \44779 , \44780 , \44781 , \44782 , \44783 , \44784 ,
         \44785 , \44786 , \44787 , \44788 , \44789 , \44790 , \44791 , \44792 , \44793 , \44794 ,
         \44795 , \44796 , \44797 , \44798 , \44799 , \44800 , \44801 , \44802 , \44803 , \44804 ,
         \44805 , \44806 , \44807 , \44808 , \44809 , \44810 , \44811 , \44812 , \44813 , \44814 ,
         \44815 , \44816 , \44817 , \44818 , \44819 , \44820 , \44821 , \44822 , \44823 , \44824 ,
         \44825 , \44826 , \44827 , \44828 , \44829 , \44830 , \44831 , \44832 , \44833 , \44834 ,
         \44835 , \44836 , \44837 , \44838 , \44839 , \44840 , \44841 , \44842 , \44843 , \44844 ,
         \44845 , \44846 , \44847 , \44848 , \44849 , \44850 , \44851 , \44852 , \44853 , \44854 ,
         \44855 , \44856 , \44857 , \44858 , \44859 , \44860 , \44861 , \44862 , \44863 , \44864 ,
         \44865 , \44866 , \44867 , \44868 , \44869 , \44870 , \44871 , \44872 , \44873 , \44874 ,
         \44875 , \44876 , \44877 , \44878 , \44879 , \44880 , \44881 , \44882 , \44883 , \44884 ,
         \44885 , \44886 , \44887 , \44888 , \44889 , \44890 , \44891 , \44892 , \44893 , \44894 ,
         \44895 , \44896 , \44897 , \44898 , \44899 , \44900 , \44901 , \44902 , \44903 , \44904 ,
         \44905 , \44906 , \44907 , \44908 , \44909 , \44910 , \44911 , \44912 , \44913 , \44914 ,
         \44915 , \44916 , \44917 , \44918 , \44919 , \44920 , \44921 , \44922 , \44923 , \44924 ,
         \44925 , \44926 , \44927 , \44928 , \44929 , \44930 , \44931 , \44932 , \44933 , \44934 ,
         \44935 , \44936 , \44937 , \44938 , \44939 , \44940 , \44941 , \44942 , \44943 , \44944 ,
         \44945 , \44946 , \44947 , \44948 , \44949 , \44950 , \44951 , \44952 , \44953 , \44954 ,
         \44955 , \44956 , \44957 , \44958 , \44959 , \44960 , \44961 , \44962 , \44963 , \44964 ,
         \44965 , \44966 , \44967 , \44968 , \44969 , \44970 , \44971 , \44972 , \44973 , \44974 ,
         \44975 , \44976 , \44977 , \44978 , \44979 , \44980 , \44981 , \44982 , \44983 , \44984 ,
         \44985 , \44986 , \44987 , \44988 , \44989 , \44990 , \44991 , \44992 , \44993 , \44994 ,
         \44995 , \44996 , \44997 , \44998 , \44999 , \45000 , \45001 , \45002 , \45003 , \45004 ,
         \45005 , \45006 , \45007 , \45008 , \45009 , \45010 , \45011 , \45012 , \45013 , \45014 ,
         \45015 , \45016 , \45017 , \45018 , \45019 , \45020 , \45021 , \45022 , \45023 , \45024 ,
         \45025 , \45026 , \45027 , \45028 , \45029 , \45030 , \45031 , \45032 , \45033 , \45034 ,
         \45035 , \45036 , \45037 , \45038 , \45039 , \45040 , \45041 , \45042 , \45043 , \45044 ,
         \45045 , \45046 , \45047 , \45048 , \45049 , \45050 , \45051 , \45052 , \45053 , \45054 ,
         \45055 , \45056 , \45057 , \45058 , \45059 , \45060 , \45061 , \45062 , \45063 , \45064 ,
         \45065 , \45066 , \45067 , \45068 , \45069 , \45070 , \45071 , \45072 , \45073 , \45074 ,
         \45075 , \45076 , \45077 , \45078 , \45079 , \45080 , \45081 , \45082 , \45083 , \45084 ,
         \45085 , \45086 , \45087 , \45088 , \45089 , \45090 , \45091 , \45092 , \45093 , \45094 ,
         \45095 , \45096 , \45097 , \45098 , \45099 , \45100 , \45101 , \45102 , \45103 , \45104 ,
         \45105 , \45106 , \45107 , \45108 , \45109 , \45110 , \45111 , \45112 , \45113 , \45114 ,
         \45115 , \45116 , \45117 , \45118 , \45119 , \45120 , \45121 , \45122 , \45123 , \45124 ,
         \45125 , \45126 , \45127 , \45128 , \45129 , \45130 , \45131 , \45132 , \45133 , \45134 ,
         \45135 , \45136 , \45137 , \45138 , \45139 , \45140 , \45141 , \45142 , \45143 , \45144 ,
         \45145 , \45146 , \45147 , \45148 , \45149 , \45150 , \45151 , \45152 , \45153 , \45154 ,
         \45155 , \45156 , \45157 , \45158 , \45159 , \45160 , \45161 , \45162 , \45163 , \45164 ,
         \45165 , \45166 , \45167 , \45168 , \45169 , \45170 , \45171 , \45172 , \45173 , \45174 ,
         \45175 , \45176 , \45177 , \45178 , \45179 , \45180 , \45181 , \45182 , \45183 , \45184 ,
         \45185 , \45186 , \45187 , \45188 , \45189 , \45190 , \45191 , \45192 , \45193 , \45194 ,
         \45195 , \45196 , \45197 , \45198 , \45199 , \45200 , \45201 , \45202 , \45203 , \45204 ,
         \45205 , \45206 , \45207 , \45208 , \45209 , \45210 , \45211 , \45212 , \45213 , \45214 ,
         \45215 , \45216 , \45217 , \45218 , \45219 , \45220 , \45221 , \45222 , \45223 , \45224 ,
         \45225 , \45226 , \45227 , \45228 , \45229 , \45230 , \45231 , \45232 , \45233 , \45234 ,
         \45235 , \45236 , \45237 , \45238 , \45239 , \45240 , \45241 , \45242 , \45243 , \45244 ,
         \45245 , \45246 , \45247 , \45248 , \45249 , \45250 , \45251 , \45252 , \45253 , \45254 ,
         \45255 , \45256 , \45257 , \45258 , \45259 , \45260 , \45261 , \45262 , \45263 , \45264 ,
         \45265 , \45266 , \45267 , \45268 , \45269 , \45270 , \45271 , \45272 , \45273 , \45274 ,
         \45275 , \45276 , \45277 , \45278 , \45279 , \45280 , \45281 , \45282 , \45283 , \45284 ,
         \45285 , \45286 , \45287 , \45288 , \45289 , \45290 , \45291 , \45292 , \45293 , \45294 ,
         \45295 , \45296 , \45297 , \45298 , \45299 , \45300 , \45301 , \45302 , \45303 , \45304 ,
         \45305 , \45306 , \45307 , \45308 , \45309 , \45310 , \45311 , \45312 , \45313 , \45314 ,
         \45315 , \45316 , \45317 , \45318 , \45319 , \45320 , \45321 , \45322 , \45323 , \45324 ,
         \45325 , \45326 , \45327 , \45328 , \45329 , \45330 , \45331 , \45332 , \45333 , \45334 ,
         \45335 , \45336 , \45337 , \45338 , \45339 , \45340 , \45341 , \45342 , \45343 , \45344 ,
         \45345 , \45346 , \45347 , \45348 , \45349 , \45350 , \45351 , \45352 , \45353 , \45354 ,
         \45355 , \45356 , \45357 , \45358 , \45359 , \45360 , \45361 , \45362 , \45363 , \45364 ,
         \45365 , \45366 , \45367 , \45368 , \45369 , \45370 , \45371 , \45372 , \45373 , \45374 ,
         \45375 , \45376 , \45377 , \45378 , \45379 , \45380 , \45381 , \45382 , \45383 , \45384 ,
         \45385 , \45386 , \45387 , \45388 , \45389 , \45390 , \45391 , \45392 , \45393 , \45394 ,
         \45395 , \45396 , \45397 , \45398 , \45399 , \45400 , \45401 , \45402 , \45403 , \45404 ,
         \45405 , \45406 , \45407 , \45408 , \45409 , \45410 , \45411 , \45412 , \45413 , \45414 ,
         \45415 , \45416 , \45417 , \45418 , \45419 , \45420 , \45421 , \45422 , \45423 , \45424 ,
         \45425 , \45426 , \45427 , \45428 , \45429 , \45430 , \45431 , \45432 , \45433 , \45434 ,
         \45435 , \45436 , \45437 , \45438 , \45439 , \45440 , \45441 , \45442 , \45443 , \45444 ,
         \45445 , \45446 , \45447 , \45448 , \45449 , \45450 , \45451 , \45452 , \45453 , \45454 ,
         \45455 , \45456 , \45457 , \45458 , \45459 , \45460 , \45461 , \45462 , \45463 , \45464 ,
         \45465 , \45466 , \45467 , \45468 , \45469 , \45470 , \45471 , \45472 , \45473 , \45474 ,
         \45475 , \45476 , \45477 , \45478 , \45479 , \45480 , \45481 , \45482 , \45483 , \45484 ,
         \45485 , \45486 , \45487 , \45488 , \45489 , \45490 , \45491 , \45492 , \45493 , \45494 ,
         \45495 , \45496 , \45497 , \45498 , \45499 , \45500 , \45501 , \45502 , \45503 , \45504 ,
         \45505 , \45506 , \45507 , \45508 , \45509 , \45510 , \45511 , \45512 , \45513 , \45514 ,
         \45515 , \45516 , \45517 , \45518 , \45519 , \45520 , \45521 , \45522 , \45523 , \45524 ,
         \45525 , \45526 , \45527 , \45528 , \45529 , \45530 , \45531 , \45532 , \45533 , \45534 ,
         \45535 , \45536 , \45537 , \45538 , \45539 , \45540 , \45541 , \45542 , \45543 , \45544 ,
         \45545 , \45546 , \45547 , \45548 , \45549 , \45550 , \45551 , \45552 , \45553 , \45554 ,
         \45555 , \45556 , \45557 , \45558 , \45559 , \45560 , \45561 , \45562 , \45563 , \45564 ,
         \45565 , \45566 , \45567 , \45568 , \45569 , \45570 , \45571 , \45572 , \45573 , \45574 ,
         \45575 , \45576 , \45577 , \45578 , \45579 , \45580 , \45581 , \45582 , \45583 , \45584 ,
         \45585 , \45586 , \45587 , \45588 , \45589 , \45590 , \45591 , \45592 , \45593 , \45594 ,
         \45595 , \45596 , \45597 , \45598 , \45599 , \45600 , \45601 , \45602 , \45603 , \45604 ,
         \45605 , \45606 , \45607 , \45608 , \45609 , \45610 , \45611 , \45612 , \45613 , \45614 ,
         \45615 , \45616 , \45617 , \45618 , \45619 , \45620 , \45621 , \45622 , \45623 , \45624 ,
         \45625 , \45626 , \45627 , \45628 , \45629 , \45630 , \45631 , \45632 , \45633 , \45634 ,
         \45635 , \45636 , \45637 , \45638 , \45639 , \45640 , \45641 , \45642 , \45643 , \45644 ,
         \45645 , \45646 , \45647 , \45648 , \45649 , \45650 , \45651 , \45652 , \45653 , \45654 ,
         \45655 , \45656 , \45657 , \45658 , \45659 , \45660 , \45661 , \45662 , \45663 , \45664 ,
         \45665 , \45666 , \45667 , \45668 , \45669 , \45670 , \45671 , \45672 , \45673 , \45674 ,
         \45675 , \45676 , \45677 , \45678 , \45679 , \45680 , \45681 , \45682 , \45683 , \45684 ,
         \45685 , \45686 , \45687 , \45688 , \45689 , \45690 , \45691 , \45692 , \45693 , \45694 ,
         \45695 , \45696 , \45697 , \45698 , \45699 , \45700 , \45701 , \45702 , \45703 , \45704 ,
         \45705 , \45706 , \45707 , \45708 , \45709 , \45710 , \45711 , \45712 , \45713 , \45714 ,
         \45715 , \45716 , \45717 , \45718 , \45719 , \45720 , \45721 , \45722 , \45723 , \45724 ,
         \45725 , \45726 , \45727 , \45728 , \45729 , \45730 , \45731 , \45732 , \45733 , \45734 ,
         \45735 , \45736 , \45737 , \45738 , \45739 , \45740 , \45741 , \45742 , \45743 , \45744 ,
         \45745 , \45746 , \45747 , \45748 , \45749 , \45750 , \45751 , \45752 , \45753 , \45754 ,
         \45755 , \45756 , \45757 , \45758 , \45759 , \45760 , \45761 , \45762 , \45763 , \45764 ,
         \45765 , \45766 , \45767 , \45768 , \45769 , \45770 , \45771 , \45772 , \45773 , \45774 ,
         \45775 , \45776 , \45777 , \45778 , \45779 , \45780 , \45781 , \45782 , \45783 , \45784 ,
         \45785 , \45786 , \45787 , \45788 , \45789 , \45790 , \45791 , \45792 , \45793 , \45794 ,
         \45795 , \45796 , \45797 , \45798 , \45799 , \45800 , \45801 , \45802 , \45803 , \45804 ,
         \45805 , \45806 , \45807 , \45808 , \45809 , \45810 , \45811 , \45812 , \45813 , \45814 ,
         \45815 , \45816 , \45817 , \45818 , \45819 , \45820 , \45821 , \45822 , \45823 , \45824 ,
         \45825 , \45826 , \45827 , \45828 , \45829 , \45830 , \45831 , \45832 , \45833 , \45834 ,
         \45835 , \45836 , \45837 , \45838 , \45839 , \45840 , \45841 , \45842 , \45843 , \45844 ,
         \45845 , \45846 , \45847 , \45848 , \45849 , \45850 , \45851 , \45852 , \45853 , \45854 ,
         \45855 , \45856 , \45857 , \45858 , \45859 , \45860 , \45861 , \45862 , \45863 , \45864 ,
         \45865 , \45866 , \45867 , \45868 , \45869 , \45870 , \45871 , \45872 , \45873 , \45874 ,
         \45875 , \45876 , \45877 , \45878 , \45879 , \45880 , \45881 , \45882 , \45883 , \45884 ,
         \45885 , \45886 , \45887 , \45888 , \45889 , \45890 , \45891 , \45892 , \45893 , \45894 ,
         \45895 , \45896 , \45897 , \45898 , \45899 , \45900 , \45901 , \45902 , \45903 , \45904 ,
         \45905 , \45906 , \45907 , \45908 , \45909 , \45910 , \45911 , \45912 , \45913 , \45914 ,
         \45915 , \45916 , \45917 , \45918 , \45919 , \45920 , \45921 , \45922 , \45923 , \45924 ,
         \45925 , \45926 , \45927 , \45928 , \45929 , \45930 , \45931 , \45932 , \45933 , \45934 ,
         \45935 , \45936 , \45937 , \45938 , \45939 , \45940 , \45941 , \45942 , \45943 , \45944 ,
         \45945 , \45946 , \45947 , \45948 , \45949 , \45950 , \45951 , \45952 , \45953 , \45954 ,
         \45955 , \45956 , \45957 , \45958 , \45959 , \45960 , \45961 , \45962 , \45963 , \45964 ,
         \45965 , \45966 , \45967 , \45968 , \45969 , \45970 , \45971 , \45972 , \45973 , \45974 ,
         \45975 , \45976 , \45977 , \45978 , \45979 , \45980 , \45981 , \45982 , \45983 , \45984 ,
         \45985 , \45986 , \45987 , \45988 , \45989 , \45990 , \45991 , \45992 , \45993 , \45994 ,
         \45995 , \45996 , \45997 , \45998 , \45999 , \46000 , \46001 , \46002 , \46003 , \46004 ,
         \46005 , \46006 , \46007 , \46008 , \46009 , \46010 , \46011 , \46012 , \46013 , \46014 ,
         \46015 , \46016 , \46017 , \46018 , \46019 , \46020 , \46021 , \46022 , \46023 , \46024 ,
         \46025 , \46026 , \46027 , \46028 , \46029 , \46030 , \46031 , \46032 , \46033 , \46034 ,
         \46035 , \46036 , \46037 , \46038 , \46039 , \46040 , \46041 , \46042 , \46043 , \46044 ,
         \46045 , \46046 , \46047 , \46048 , \46049 , \46050 , \46051 , \46052 , \46053 , \46054 ,
         \46055 , \46056 , \46057 , \46058 , \46059 , \46060 , \46061 , \46062 , \46063 , \46064 ,
         \46065 , \46066 , \46067 , \46068 , \46069 , \46070 , \46071 , \46072 , \46073 , \46074 ,
         \46075 , \46076 , \46077 , \46078 , \46079 , \46080 , \46081 , \46082 , \46083 , \46084 ,
         \46085 , \46086 , \46087 , \46088 , \46089 , \46090 , \46091 , \46092 , \46093 , \46094 ,
         \46095 , \46096 , \46097 , \46098 , \46099 , \46100 , \46101 , \46102 , \46103 , \46104 ,
         \46105 , \46106 , \46107 , \46108 , \46109 , \46110 , \46111 , \46112 , \46113 , \46114 ,
         \46115 , \46116 , \46117 , \46118 , \46119 , \46120 , \46121 , \46122 , \46123 , \46124 ,
         \46125 , \46126 , \46127 , \46128 , \46129 , \46130 , \46131 , \46132 , \46133 , \46134 ,
         \46135 , \46136 , \46137 , \46138 , \46139 , \46140 , \46141 , \46142 , \46143 , \46144 ,
         \46145 , \46146 , \46147 , \46148 , \46149 , \46150 , \46151 , \46152 , \46153 , \46154 ,
         \46155 , \46156 , \46157 , \46158 , \46159 , \46160 , \46161 , \46162 , \46163 , \46164 ,
         \46165 , \46166 , \46167 , \46168 , \46169 , \46170 , \46171 , \46172 , \46173 , \46174 ,
         \46175 , \46176 , \46177 , \46178 , \46179 , \46180 , \46181 , \46182 , \46183 , \46184 ,
         \46185 , \46186 , \46187 , \46188 , \46189 , \46190 , \46191 , \46192 , \46193 , \46194 ,
         \46195 , \46196 , \46197 , \46198 , \46199 , \46200 , \46201 , \46202 , \46203 , \46204 ,
         \46205 , \46206 , \46207 , \46208 , \46209 , \46210 , \46211 , \46212 , \46213 , \46214 ,
         \46215 , \46216 , \46217 , \46218 , \46219 , \46220 , \46221 , \46222 , \46223 , \46224 ,
         \46225 , \46226 , \46227 , \46228 , \46229 , \46230 , \46231 , \46232 , \46233 , \46234 ,
         \46235 , \46236 , \46237 , \46238 , \46239 , \46240 , \46241 , \46242 , \46243 , \46244 ,
         \46245 , \46246 , \46247 , \46248 , \46249 , \46250 , \46251 , \46252 , \46253 , \46254 ,
         \46255 , \46256 , \46257 , \46258 , \46259 , \46260 , \46261 , \46262 , \46263 , \46264 ,
         \46265 , \46266 , \46267 , \46268 , \46269 , \46270 , \46271 , \46272 , \46273 , \46274 ,
         \46275 , \46276 , \46277 , \46278 , \46279 , \46280 , \46281 , \46282 , \46283 , \46284 ,
         \46285 , \46286 , \46287 , \46288 , \46289 , \46290 , \46291 , \46292 , \46293 , \46294 ,
         \46295 , \46296 , \46297 , \46298 , \46299 , \46300 , \46301 , \46302 , \46303 , \46304 ,
         \46305 , \46306 , \46307 , \46308 , \46309 , \46310 , \46311 , \46312 , \46313 , \46314 ,
         \46315 , \46316 , \46317 , \46318 , \46319 , \46320 , \46321 , \46322 , \46323 , \46324 ,
         \46325 , \46326 , \46327 , \46328 , \46329 , \46330 , \46331 , \46332 , \46333 , \46334 ,
         \46335 , \46336 , \46337 , \46338 , \46339 , \46340 , \46341 , \46342 , \46343 , \46344 ,
         \46345 , \46346 , \46347 , \46348 , \46349 , \46350 , \46351 , \46352 , \46353 , \46354 ,
         \46355 , \46356 , \46357 , \46358 , \46359 , \46360 , \46361 , \46362 , \46363 , \46364 ,
         \46365 , \46366 , \46367 , \46368 , \46369 , \46370 , \46371 , \46372 , \46373 , \46374 ,
         \46375 , \46376 , \46377 , \46378 , \46379 , \46380 , \46381 , \46382 , \46383 , \46384 ,
         \46385 , \46386 , \46387 , \46388 , \46389 , \46390 , \46391 , \46392 , \46393 , \46394 ,
         \46395 , \46396 , \46397 , \46398 , \46399 , \46400 , \46401 , \46402 , \46403 , \46404 ,
         \46405 , \46406 , \46407 , \46408 , \46409 , \46410 , \46411 , \46412 , \46413 , \46414 ,
         \46415 , \46416 , \46417 , \46418 , \46419 , \46420 , \46421 , \46422 , \46423 , \46424 ,
         \46425 , \46426 , \46427 , \46428 , \46429 , \46430 , \46431 , \46432 , \46433 , \46434 ,
         \46435 , \46436 , \46437 , \46438 , \46439 , \46440 , \46441 , \46442 , \46443 , \46444 ,
         \46445 , \46446 , \46447 , \46448 , \46449 , \46450 , \46451 , \46452 , \46453 , \46454 ,
         \46455 , \46456 , \46457 , \46458 , \46459 , \46460 , \46461 , \46462 , \46463 , \46464 ,
         \46465 , \46466 , \46467 , \46468 , \46469 , \46470 , \46471 , \46472 , \46473 , \46474 ,
         \46475 , \46476 , \46477 , \46478 , \46479 , \46480 , \46481 , \46482 , \46483 , \46484 ,
         \46485 , \46486 , \46487 , \46488 , \46489 , \46490 , \46491 , \46492 , \46493 , \46494 ,
         \46495 , \46496 , \46497 , \46498 , \46499 , \46500 , \46501 , \46502 , \46503 , \46504 ,
         \46505 , \46506 , \46507 , \46508 , \46509 , \46510 , \46511 , \46512 , \46513 , \46514 ,
         \46515 , \46516 , \46517 , \46518 , \46519 , \46520 , \46521 , \46522 , \46523 , \46524 ,
         \46525 , \46526 , \46527 , \46528 , \46529 , \46530 , \46531 , \46532 , \46533 , \46534 ,
         \46535 , \46536 , \46537 , \46538 , \46539 , \46540 , \46541 , \46542 , \46543 , \46544 ,
         \46545 , \46546 , \46547 , \46548 , \46549 , \46550 , \46551 , \46552 , \46553 , \46554 ,
         \46555 , \46556 , \46557 , \46558 , \46559 , \46560 , \46561 , \46562 , \46563 , \46564 ,
         \46565 , \46566 , \46567 , \46568 , \46569 , \46570 , \46571 , \46572 , \46573 , \46574 ,
         \46575 , \46576 , \46577 , \46578 , \46579 , \46580 , \46581 , \46582 , \46583 , \46584 ,
         \46585 , \46586 , \46587 , \46588 , \46589 , \46590 , \46591 , \46592 , \46593 , \46594 ,
         \46595 , \46596 , \46597 , \46598 , \46599 , \46600 , \46601 , \46602 , \46603 , \46604 ,
         \46605 , \46606 , \46607 , \46608 , \46609 , \46610 , \46611 , \46612 , \46613 , \46614 ,
         \46615 , \46616 , \46617 , \46618 , \46619 , \46620 , \46621 , \46622 , \46623 , \46624 ,
         \46625 , \46626 , \46627 , \46628 , \46629 , \46630 , \46631 , \46632 , \46633 , \46634 ,
         \46635 , \46636 , \46637 , \46638 , \46639 , \46640 , \46641 , \46642 , \46643 , \46644 ,
         \46645 , \46646 , \46647 , \46648 , \46649 , \46650 , \46651 , \46652 , \46653 , \46654 ,
         \46655 , \46656 , \46657 , \46658 , \46659 , \46660 , \46661 , \46662 , \46663 , \46664 ,
         \46665 , \46666 , \46667 , \46668 , \46669 , \46670 , \46671 , \46672 , \46673 , \46674 ,
         \46675 , \46676 , \46677 , \46678 , \46679 , \46680 , \46681 , \46682 , \46683 , \46684 ,
         \46685 , \46686 , \46687 , \46688 , \46689 , \46690 , \46691 , \46692 , \46693 , \46694 ,
         \46695 , \46696 , \46697 , \46698 , \46699 , \46700 , \46701 , \46702 , \46703 , \46704 ,
         \46705 , \46706 , \46707 , \46708 , \46709 , \46710 , \46711 , \46712 , \46713 , \46714 ,
         \46715 , \46716 , \46717 , \46718 , \46719 , \46720 , \46721 , \46722 , \46723 , \46724 ,
         \46725 , \46726 , \46727 , \46728 , \46729 , \46730 , \46731 , \46732 , \46733 , \46734 ,
         \46735 , \46736 , \46737 , \46738 , \46739 , \46740 , \46741 , \46742 , \46743 , \46744 ,
         \46745 , \46746 , \46747 , \46748 , \46749 , \46750 , \46751 , \46752 , \46753 , \46754 ,
         \46755 , \46756 , \46757 , \46758 , \46759 , \46760 , \46761 , \46762 , \46763 , \46764 ,
         \46765 , \46766 , \46767 , \46768 , \46769 , \46770 , \46771 , \46772 , \46773 , \46774 ,
         \46775 , \46776 , \46777 , \46778 , \46779 , \46780 , \46781 , \46782 , \46783 , \46784 ,
         \46785 , \46786 ;
buf \U$labajz4723 ( R_101_77c8620, \45206 );
buf \U$labajz4724 ( R_102_af8fd30, \45240 );
buf \U$labajz4725 ( R_103_af901c8, \45255 );
buf \U$labajz4726 ( R_104_af9a140, \45267 );
buf \U$labajz4727 ( R_105_af99768, \45284 );
buf \U$labajz4728 ( R_106_af8be30, \45296 );
buf \U$labajz4729 ( R_107_77c1150, \45310 );
buf \U$labajz4730 ( R_108_af8ddb0, \45314 );
buf \U$labajz4731 ( R_109_af8f010, \45325 );
buf \U$labajz4732 ( R_10a_af996c0, \45353 );
buf \U$labajz4733 ( R_10b_77c34c0, \45367 );
buf \U$labajz4734 ( R_10c_77c28f0, \45376 );
buf \U$labajz4735 ( R_10d_af8d090, \45402 );
buf \U$labajz4736 ( R_10e_77ca5a0, \45406 );
buf \U$labajz4737 ( R_10f_77ce4a0, \45414 );
buf \U$labajz4738 ( R_110_77cd780, \45419 );
buf \U$labajz4739 ( R_111_af8f2b0, \45446 );
buf \U$labajz4740 ( R_112_77c6550, \45466 );
buf \U$labajz4741 ( R_113_af98ee0, \45474 );
buf \U$labajz4742 ( R_114_77c2068, \45482 );
buf \U$labajz4743 ( R_115_af99ea0, \45506 );
buf \U$labajz4744 ( R_116_77c0eb0, \45510 );
buf \U$labajz4745 ( R_117_77cc280, \45519 );
buf \U$labajz4746 ( R_118_77bf860, \45523 );
buf \U$labajz4747 ( R_119_77c9f10, \45537 );
buf \U$labajz4748 ( R_11a_af8bf80, \45548 );
buf \U$labajz4749 ( R_11b_77bf320, \45556 );
buf \U$labajz4750 ( R_11c_77c4fa8, \45560 );
buf \U$labajz4751 ( R_11d_af99ab0, \45574 );
buf \U$labajz4752 ( R_11e_77ca258, \45583 );
buf \U$labajz4753 ( R_11f_af92880, \45592 );
buf \U$labajz4754 ( R_120_af91c08, \45596 );
buf \U$labajz4755 ( R_121_af92298, \45628 );
buf \U$labajz4756 ( R_122_af99ca8, \45641 );
buf \U$labajz4757 ( R_123_af990d8, \45655 );
buf \U$labajz4758 ( R_124_77c5638, \45659 );
buf \U$labajz4759 ( R_125_af8e6e0, \45683 );
buf \U$labajz4760 ( R_126_77c3aa8, \45691 );
buf \U$labajz4761 ( R_127_77c8d58, \45705 );
buf \U$labajz4762 ( R_128_77c1fc0, \45710 );
buf \U$labajz4763 ( R_129_77c6748, \45740 );
buf \U$labajz4764 ( R_12a_77c3370, \45748 );
buf \U$labajz4765 ( R_12b_af99d50, \45764 );
buf \U$labajz4766 ( R_12c_77c5248, \45768 );
buf \U$labajz4767 ( R_12d_77ca840, \45789 );
buf \U$labajz4768 ( R_12e_af8eec0, \45803 );
buf \U$labajz4769 ( R_12f_77c1498, \45815 );
buf \U$labajz4770 ( R_130_77c5398, \45823 );
buf \U$labajz4771 ( R_131_77c0820, \45871 );
buf \U$labajz4772 ( R_132_af8d480, \45876 );
buf \U$labajz4773 ( R_133_77ce890, \45888 );
buf \U$labajz4774 ( R_134_af97c80, \45897 );
buf \U$labajz4775 ( R_135_77c65f8, \45914 );
buf \U$labajz4776 ( R_136_af8d678, \45927 );
buf \U$labajz4777 ( R_137_77c3e98, \45942 );
buf \U$labajz4778 ( R_138_af8e0f8, \45946 );
buf \U$labajz4779 ( R_139_af99378, \45972 );
buf \U$labajz4780 ( R_13a_77c7078, \45980 );
buf \U$labajz4781 ( R_13b_77ce740, \45994 );
buf \U$labajz4782 ( R_13c_af97fc8, \46002 );
buf \U$labajz4783 ( R_13d_77c62b0, \46021 );
buf \U$labajz4784 ( R_13e_77c27a0, \46025 );
buf \U$labajz4785 ( R_13f_af979e0, \46034 );
buf \U$labajz4786 ( R_140_77c25a8, \46042 );
buf \U$labajz4787 ( R_141_af921f0, \46076 );
buf \U$labajz4788 ( R_142_af8b7a0, \46082 );
buf \U$labajz4789 ( R_143_77bfcf8, \46097 );
buf \U$labajz4790 ( R_144_af92148, \46104 );
buf \U$labajz4791 ( R_145_77c1c78, \46124 );
buf \U$labajz4792 ( R_146_77cb560, \46135 );
buf \U$labajz4793 ( R_147_af99960, \46149 );
buf \U$labajz4794 ( R_148_af92490, \46159 );
buf \U$labajz4795 ( R_149_77c9298, \46189 );
buf \U$labajz4796 ( R_14a_77cb170, \46200 );
buf \U$labajz4797 ( R_14b_af98268, \46216 );
buf \U$labajz4798 ( R_14c_77bf9b0, \46226 );
buf \U$labajz4799 ( R_14d_af91b60, \46248 );
buf \U$labajz4800 ( R_14e_af8f208, \46259 );
buf \U$labajz4801 ( R_14f_77c7a50, \46271 );
buf \U$labajz4802 ( R_150_af99030, \46277 );
buf \U$labajz4803 ( R_151_77c67f0, \46306 );
buf \U$labajz4804 ( R_152_af8c370, \46312 );
buf \U$labajz4805 ( R_153_77c8818, \46319 );
buf \U$labajz4806 ( R_154_77c6d30, \46326 );
buf \U$labajz4807 ( R_155_af98c40, \46352 );
buf \U$labajz4808 ( R_156_77c9538, \46363 );
buf \U$labajz4809 ( R_157_af96f60, \46379 );
buf \U$labajz4810 ( R_158_af96d68, \46386 );
buf \U$labajz4811 ( R_159_af8d870, \46412 );
buf \U$labajz4812 ( R_15a_af8e830, \46422 );
buf \U$labajz4813 ( R_15b_77ccbb0, \46437 );
buf \U$labajz4814 ( R_15c_af8c610, \46447 );
buf \U$labajz4815 ( R_15d_77c6898, \46467 );
buf \U$labajz4816 ( R_15e_af8cb50, \46477 );
buf \U$labajz4817 ( R_15f_af92538, \46488 );
buf \U$labajz4818 ( R_160_af975f0, \46494 );
buf \U$labajz4819 ( R_161_77c71c8, \46518 );
buf \U$labajz4820 ( R_162_af8d720, \46528 );
buf \U$labajz4821 ( R_163_77cb608, \46542 );
buf \U$labajz4822 ( R_164_af8b650, \46552 );
buf \U$labajz4823 ( R_165_af988f8, \46575 );
buf \U$labajz4824 ( R_166_77c41e0, \46585 );
buf \U$labajz4825 ( R_167_af8e398, \46600 );
buf \U$labajz4826 ( R_168_af974a0, \46610 );
buf \U$labajz4827 ( R_169_af8d330, \46628 );
buf \U$labajz4828 ( R_16a_af8c0d0, \46639 );
buf \U$labajz4829 ( R_16b_77cc520, \46655 );
buf \U$labajz4830 ( R_16c_77cb8a8, \46665 );
buf \U$labajz4831 ( R_16d_77ccda8, \46681 );
buf \U$labajz4832 ( R_16e_af973f8, \46691 );
buf \U$labajz4833 ( R_16f_77cd6d8, \46703 );
buf \U$labajz4834 ( R_170_af99ff0, \46710 );
buf \U$labajz4835 ( R_171_77c54e8, \46732 );
buf \U$labajz4836 ( R_172_77c3808, \46742 );
buf \U$labajz4837 ( R_173_77c0580, \46758 );
buf \U$labajz4838 ( R_174_af99618, \46764 );
buf \U$labajz4839 ( R_175_77cd198, \46773 );
buf \U$labajz4840 ( R_176_77c0628, \46780 );
buf \U$labajz4841 ( R_177_af97698, \46786 );
nor \U$1 ( \378 , RIae76b68_57, RIae76be0_58);
nor \U$2 ( \379 , RIae78a58_123, RIae78ad0_124);
nor \U$3 ( \380 , \378 , \379 );
not \U$4 ( \381 , \380 );
nor \U$5 ( \382 , RIae76028_33, RIae760a0_34);
nor \U$6 ( \383 , RIae76118_35, RIae76190_36);
nor \U$7 ( \384 , \382 , \383 );
or \U$8 ( \385 , RIae762f8_39, RIae76370_40);
or \U$9 ( \386 , RIae76208_37, RIae76280_38);
and \U$10 ( \387 , \384 , \385 , \386 );
nor \U$11 ( \388 , RIae763e8_41, RIae76460_42);
nor \U$12 ( \389 , RIae764d8_43, RIae76550_44);
nor \U$13 ( \390 , \388 , \389 );
or \U$14 ( \391 , RIae76730_48, RIae766b8_47);
or \U$15 ( \392 , RIae76640_46, RIae765c8_45);
and \U$16 ( \393 , \390 , \391 , \392 );
nor \U$17 ( \394 , RIae76988_53, RIae76a00_54);
nor \U$18 ( \395 , RIae76a78_55, RIae76af0_56);
nor \U$19 ( \396 , \394 , \395 );
or \U$20 ( \397 , RIae767a8_49, RIae76820_50);
or \U$21 ( \398 , RIae76898_51, RIae76910_52);
and \U$22 ( \399 , \396 , \397 , \398 );
and \U$23 ( \400 , \387 , \393 , \399 );
not \U$24 ( \401 , \400 );
nor \U$25 ( \402 , RIae77798_83, RIae77810_84);
nor \U$26 ( \403 , RIae77888_85, RIae77900_86);
nor \U$27 ( \404 , \402 , \403 );
not \U$28 ( \405 , \404 );
nand \U$29 ( \406 , RIae77a68_89, RIae77ae0_90);
nor \U$30 ( \407 , RIae77978_87, RIae779f0_88);
or \U$31 ( \408 , \406 , \407 );
nand \U$32 ( \409 , RIae77978_87, RIae779f0_88);
nand \U$33 ( \410 , \408 , \409 );
not \U$34 ( \411 , \410 );
or \U$35 ( \412 , \405 , \411 );
nor \U$36 ( \413 , RIae77888_85, RIae77900_86);
nand \U$37 ( \414 , RIae77798_83, RIae77810_84);
or \U$38 ( \415 , \413 , \414 );
nand \U$39 ( \416 , RIae77888_85, RIae77900_86);
nand \U$40 ( \417 , \415 , \416 );
not \U$41 ( \418 , \417 );
nand \U$42 ( \419 , \412 , \418 );
nor \U$43 ( \420 , RIae77108_69, RIae77180_70);
nor \U$44 ( \421 , RIae77018_67, RIae77090_68);
nor \U$45 ( \422 , \420 , \421 );
nor \U$46 ( \423 , RIae772e8_73, RIae77360_74);
nor \U$47 ( \424 , RIae771f8_71, RIae77270_72);
nor \U$48 ( \425 , \423 , \424 );
nand \U$49 ( \426 , \422 , \425 );
not \U$50 ( \427 , \426 );
nor \U$51 ( \428 , RIae76c58_59, RIae76cd0_60);
nor \U$52 ( \429 , RIae76d48_61, RIae76dc0_62);
nor \U$53 ( \430 , \428 , \429 );
nor \U$54 ( \431 , RIae76f28_65, RIae76fa0_66);
nor \U$55 ( \432 , RIae76e38_63, RIae76eb0_64);
nor \U$56 ( \433 , \431 , \432 );
nand \U$57 ( \434 , \430 , \433 );
not \U$58 ( \435 , \434 );
nand \U$59 ( \436 , \419 , \427 , \435 );
nor \U$60 ( \437 , RIae77018_67, RIae77090_68);
nand \U$61 ( \438 , RIae77108_69, RIae77180_70);
or \U$62 ( \439 , \437 , \438 );
nand \U$63 ( \440 , RIae77018_67, RIae77090_68);
nand \U$64 ( \441 , \439 , \440 );
not \U$65 ( \442 , \441 );
not \U$66 ( \443 , \425 );
or \U$67 ( \444 , \442 , \443 );
nor \U$68 ( \445 , RIae772e8_73, RIae77360_74);
not \U$69 ( \446 , \445 );
nand \U$70 ( \447 , RIae771f8_71, RIae77270_72);
not \U$71 ( \448 , \447 );
and \U$72 ( \449 , \446 , \448 );
and \U$73 ( \450 , RIae772e8_73, RIae77360_74);
nor \U$74 ( \451 , \449 , \450 );
nand \U$75 ( \452 , \444 , \451 );
not \U$76 ( \453 , \452 );
nor \U$77 ( \454 , RIae780f8_103, RIae78170_104);
nand \U$78 ( \455 , RIae782d8_107, RIae78350_108);
or \U$79 ( \456 , \454 , \455 );
nand \U$80 ( \457 , RIae780f8_103, RIae78170_104);
nand \U$81 ( \458 , \456 , \457 );
nand \U$82 ( \459 , RIae77f18_99, RIae77f90_100);
nand \U$83 ( \460 , RIae78008_101, RIae78080_102);
nand \U$84 ( \461 , \459 , \460 );
nor \U$85 ( \462 , \458 , \461 );
nand \U$86 ( \463 , \436 , \453 , \462 );
nor \U$87 ( \464 , RIae77e28_97, RIae77ea0_98);
nor \U$88 ( \465 , RIae78698_115, RIae78710_116);
nor \U$89 ( \466 , \464 , \465 );
not \U$90 ( \467 , \466 );
not \U$91 ( \468 , RIae78968_121);
not \U$92 ( \469 , RIae789e0_122);
nand \U$93 ( \470 , \468 , \469 );
nor \U$94 ( \471 , RIae78878_119, RIae788f0_120);
not \U$95 ( \472 , \471 );
not \U$96 ( \473 , RIae78788_117);
not \U$97 ( \474 , RIae78800_118);
nand \U$98 ( \475 , \473 , \474 );
nand \U$99 ( \476 , \470 , \472 , \475 );
nor \U$100 ( \477 , \467 , \476 );
nor \U$101 ( \478 , RIae77b58_91, RIae77bd0_92);
not \U$102 ( \479 , \478 );
not \U$103 ( \480 , RIae77c48_93);
not \U$104 ( \481 , RIae77cc0_94);
nand \U$105 ( \482 , \480 , \481 );
not \U$106 ( \483 , RIae77d38_95);
not \U$107 ( \484 , RIae77db0_96);
nand \U$108 ( \485 , \483 , \484 );
and \U$109 ( \486 , \479 , \482 , \485 );
nand \U$110 ( \487 , \477 , \486 );
not \U$111 ( \488 , \487 );
nor \U$112 ( \489 , RIae77f18_99, RIae77f90_100);
nor \U$113 ( \490 , RIae78008_101, RIae78080_102);
nor \U$114 ( \491 , \489 , \490 );
not \U$115 ( \492 , RIae780f8_103);
not \U$116 ( \493 , RIae78170_104);
and \U$117 ( \494 , \492 , \493 );
nor \U$118 ( \495 , RIae782d8_107, RIae78350_108);
nor \U$119 ( \496 , \494 , \495 );
nand \U$120 ( \497 , \491 , \496 );
and \U$121 ( \498 , RIae780f8_103, RIae78170_104);
and \U$122 ( \499 , RIae77f18_99, RIae77f90_100);
nor \U$123 ( \500 , \498 , \499 );
nand \U$124 ( \501 , \497 , \500 );
not \U$125 ( \502 , \501 );
not \U$126 ( \503 , \491 );
or \U$127 ( \504 , \502 , \503 );
nand \U$128 ( \505 , \504 , \460 );
not \U$129 ( \506 , RIae785a8_113);
not \U$130 ( \507 , RIae78620_114);
and \U$131 ( \508 , \506 , \507 );
nor \U$132 ( \509 , RIae781e8_105, RIae78260_106);
nor \U$133 ( \510 , \508 , \509 );
nor \U$134 ( \511 , RIae784b8_111, RIae78530_112);
nor \U$135 ( \512 , RIae783c8_109, RIae78440_110);
nor \U$136 ( \513 , \511 , \512 );
nand \U$137 ( \514 , \510 , \513 );
not \U$138 ( \515 , \514 );
nand \U$139 ( \516 , \463 , \488 , \505 , \515 );
not \U$140 ( \517 , \516 );
nor \U$141 ( \518 , RIae774c8_77, RIae77540_78);
nor \U$142 ( \519 , RIae776a8_81, RIae77720_82);
nor \U$143 ( \520 , \518 , \519 );
not \U$144 ( \521 , RIae77450_76);
not \U$145 ( \522 , RIae773d8_75);
nand \U$146 ( \523 , \521 , \522 );
not \U$147 ( \524 , RIae774c8_77);
not \U$148 ( \525 , RIae77540_78);
or \U$149 ( \526 , \524 , \525 );
nand \U$150 ( \527 , RIae775b8_79, RIae77630_80);
nand \U$151 ( \528 , \526 , \527 );
nand \U$152 ( \529 , \520 , \523 , \528 );
nand \U$153 ( \530 , RIae776a8_81, RIae77720_82);
not \U$154 ( \531 , \530 );
nand \U$155 ( \532 , \531 , \523 );
nand \U$156 ( \533 , RIae773d8_75, RIae77450_76);
nand \U$157 ( \534 , \529 , \532 , \533 );
not \U$158 ( \535 , \534 );
nor \U$159 ( \536 , RIae77a68_89, RIae77ae0_90);
nor \U$160 ( \537 , RIae77978_87, RIae779f0_88);
nor \U$161 ( \538 , \536 , \537 );
nand \U$162 ( \539 , \404 , \538 );
nor \U$163 ( \540 , \434 , \539 , \426 );
not \U$164 ( \541 , \540 );
or \U$165 ( \542 , \535 , \541 );
nand \U$166 ( \543 , RIae76c58_59, RIae76cd0_60);
nand \U$167 ( \544 , RIae76d48_61, RIae76dc0_62);
nand \U$168 ( \545 , \543 , \544 );
or \U$169 ( \546 , RIae76c58_59, RIae76cd0_60);
nand \U$170 ( \547 , \545 , \546 );
not \U$171 ( \548 , \547 );
nor \U$172 ( \549 , RIae76e38_63, RIae76eb0_64);
nand \U$173 ( \550 , RIae76f28_65, RIae76fa0_66);
or \U$174 ( \551 , \549 , \550 );
nand \U$175 ( \552 , RIae76e38_63, RIae76eb0_64);
nand \U$176 ( \553 , \551 , \552 );
nand \U$177 ( \554 , \553 , \430 );
not \U$178 ( \555 , \554 );
or \U$179 ( \556 , \548 , \555 );
nand \U$180 ( \557 , \556 , \427 );
nand \U$181 ( \558 , \542 , \557 );
not \U$182 ( \559 , \558 );
not \U$183 ( \560 , \477 );
not \U$184 ( \561 , \514 );
not \U$185 ( \562 , \497 );
nand \U$186 ( \563 , \561 , \486 , \562 );
nor \U$187 ( \564 , \560 , \563 );
not \U$188 ( \565 , \564 );
or \U$189 ( \566 , \559 , \565 );
not \U$190 ( \567 , \513 );
nand \U$191 ( \568 , RIae781e8_105, RIae78260_106);
not \U$192 ( \569 , \568 );
not \U$193 ( \570 , \569 );
nand \U$194 ( \571 , \506 , \507 );
not \U$195 ( \572 , \571 );
or \U$196 ( \573 , \570 , \572 );
nand \U$197 ( \574 , RIae785a8_113, RIae78620_114);
nand \U$198 ( \575 , \573 , \574 );
not \U$199 ( \576 , \575 );
or \U$200 ( \577 , \567 , \576 );
nand \U$201 ( \578 , RIae783c8_109, RIae78440_110);
or \U$202 ( \579 , \511 , \578 );
nand \U$203 ( \580 , RIae784b8_111, RIae78530_112);
nand \U$204 ( \581 , \579 , \580 );
not \U$205 ( \582 , \581 );
nand \U$206 ( \583 , \577 , \582 );
and \U$207 ( \584 , \488 , \583 );
nand \U$208 ( \585 , RIae77d38_95, RIae77db0_96);
nand \U$209 ( \586 , RIae77e28_97, RIae77ea0_98);
and \U$210 ( \587 , \585 , \586 );
not \U$211 ( \588 , \587 );
nand \U$212 ( \589 , RIae77c48_93, RIae77cc0_94);
or \U$213 ( \590 , \478 , \589 );
nand \U$214 ( \591 , RIae77b58_91, RIae77bd0_92);
nand \U$215 ( \592 , \590 , \591 );
nand \U$216 ( \593 , \592 , \485 );
not \U$217 ( \594 , \593 );
or \U$218 ( \595 , \588 , \594 );
nand \U$219 ( \596 , \595 , \477 );
not \U$220 ( \597 , \475 );
nand \U$221 ( \598 , RIae78968_121, RIae789e0_122);
nor \U$222 ( \599 , RIae78878_119, RIae788f0_120);
or \U$223 ( \600 , \598 , \599 );
nand \U$224 ( \601 , RIae78878_119, RIae788f0_120);
nand \U$225 ( \602 , \600 , \601 );
not \U$226 ( \603 , \602 );
or \U$227 ( \604 , \597 , \603 );
nand \U$228 ( \605 , RIae78788_117, RIae78800_118);
nand \U$229 ( \606 , \604 , \605 );
not \U$230 ( \607 , \465 );
nand \U$231 ( \608 , \606 , \607 );
nand \U$232 ( \609 , RIae78698_115, RIae78710_116);
nand \U$233 ( \610 , \596 , \608 , \609 );
nor \U$234 ( \611 , \584 , \610 );
nand \U$235 ( \612 , \566 , \611 );
or \U$236 ( \613 , \517 , \612 );
or \U$237 ( \614 , RIae755d8_11, RIae75650_12);
nor \U$238 ( \615 , RIae754e8_9, RIae75560_10);
not \U$239 ( \616 , \615 );
or \U$240 ( \617 , RIae75830_16, RIae757b8_15);
or \U$241 ( \618 , RIae756c8_13, RIae75740_14);
and \U$242 ( \619 , \614 , \616 , \617 , \618 );
or \U$243 ( \620 , RIae75380_6, RIae75308_5);
or \U$244 ( \621 , RIae75218_3, RIae75290_4);
nor \U$245 ( \622 , RIae75128_1, RIae751a0_2);
not \U$246 ( \623 , \622 );
or \U$247 ( \624 , RIae753f8_7, RIae75470_8);
and \U$248 ( \625 , \620 , \621 , \623 , \624 );
nand \U$249 ( \626 , \619 , \625 );
or \U$250 ( \627 , RIae75998_19, RIae75a10_20);
or \U$251 ( \628 , RIae758a8_17, RIae75920_18);
nand \U$252 ( \629 , \627 , \628 );
or \U$253 ( \630 , RIae75b78_23, RIae75bf0_24);
or \U$254 ( \631 , RIae75a88_21, RIae75b00_22);
nand \U$255 ( \632 , \630 , \631 );
nor \U$256 ( \633 , \629 , \632 );
nor \U$257 ( \634 , RIae75e48_29, RIae75ec0_30);
nor \U$258 ( \635 , RIae75f38_31, RIae75fb0_32);
nor \U$259 ( \636 , \634 , \635 );
or \U$260 ( \637 , RIae75c68_25, RIae75ce0_26);
and \U$261 ( \638 , \636 , \637 );
nor \U$262 ( \639 , RIae75d58_27, RIae75dd0_28);
not \U$263 ( \640 , \639 );
nand \U$264 ( \641 , \633 , \638 , \640 );
nor \U$265 ( \642 , \626 , \641 );
nand \U$266 ( \643 , \613 , \642 );
nor \U$267 ( \644 , RIae75a88_21, RIae75b00_22);
nand \U$268 ( \645 , RIae75b78_23, RIae75bf0_24);
or \U$269 ( \646 , \644 , \645 );
nand \U$270 ( \647 , RIae75a88_21, RIae75b00_22);
nand \U$271 ( \648 , \646 , \647 );
and \U$272 ( \649 , RIae75998_19, RIae75a10_20);
or \U$273 ( \650 , \648 , \649 );
or \U$274 ( \651 , RIae75a10_20, RIae75998_19);
nand \U$275 ( \652 , \650 , \651 );
not \U$276 ( \653 , \652 );
nand \U$277 ( \654 , RIae758a8_17, RIae75920_18);
not \U$278 ( \655 , \654 );
or \U$279 ( \656 , \653 , \655 );
nor \U$280 ( \657 , RIae758a8_17, RIae75920_18);
nor \U$281 ( \658 , \657 , \639 );
and \U$282 ( \659 , \636 , \658 , \637 );
nand \U$283 ( \660 , \656 , \659 );
not \U$284 ( \661 , \637 );
nand \U$285 ( \662 , RIae75f38_31, RIae75fb0_32);
or \U$286 ( \663 , \634 , \662 );
nand \U$287 ( \664 , RIae75e48_29, RIae75ec0_30);
nand \U$288 ( \665 , \663 , \664 );
not \U$289 ( \666 , \665 );
or \U$290 ( \667 , \661 , \666 );
nand \U$291 ( \668 , RIae75c68_25, RIae75ce0_26);
nand \U$292 ( \669 , \667 , \668 );
nand \U$293 ( \670 , \669 , \640 );
nand \U$294 ( \671 , RIae75d58_27, RIae75dd0_28);
nand \U$295 ( \672 , \660 , \670 , \671 );
and \U$296 ( \673 , \619 , \625 );
nand \U$297 ( \674 , \672 , \673 );
not \U$298 ( \675 , \625 );
not \U$299 ( \676 , \618 );
not \U$300 ( \677 , \617 );
nand \U$301 ( \678 , RIae755d8_11, RIae75650_12);
or \U$302 ( \679 , \678 , \615 );
nand \U$303 ( \680 , RIae754e8_9, RIae75560_10);
nand \U$304 ( \681 , \679 , \680 );
not \U$305 ( \682 , \681 );
or \U$306 ( \683 , \677 , \682 );
nand \U$307 ( \684 , RIae757b8_15, RIae75830_16);
nand \U$308 ( \685 , \683 , \684 );
not \U$309 ( \686 , \685 );
or \U$310 ( \687 , \676 , \686 );
nand \U$311 ( \688 , RIae756c8_13, RIae75740_14);
nand \U$312 ( \689 , \687 , \688 );
not \U$313 ( \690 , \689 );
or \U$314 ( \691 , \675 , \690 );
not \U$315 ( \692 , \624 );
not \U$316 ( \693 , \620 );
nand \U$317 ( \694 , RIae75218_3, RIae75290_4);
or \U$318 ( \695 , \622 , \694 );
nand \U$319 ( \696 , RIae75128_1, RIae751a0_2);
nand \U$320 ( \697 , \695 , \696 );
not \U$321 ( \698 , \697 );
or \U$322 ( \699 , \693 , \698 );
nand \U$323 ( \700 , RIae75308_5, RIae75380_6);
nand \U$324 ( \701 , \699 , \700 );
not \U$325 ( \702 , \701 );
or \U$326 ( \703 , \692 , \702 );
nand \U$327 ( \704 , RIae753f8_7, RIae75470_8);
nand \U$328 ( \705 , \703 , \704 );
not \U$329 ( \706 , \705 );
nand \U$330 ( \707 , \691 , \706 );
not \U$331 ( \708 , \707 );
and \U$332 ( \709 , \674 , \708 );
nand \U$333 ( \710 , \643 , \709 );
not \U$334 ( \711 , \710 );
or \U$335 ( \712 , \401 , \711 );
not \U$336 ( \713 , \399 );
not \U$337 ( \714 , \387 );
not \U$338 ( \715 , \392 );
not \U$339 ( \716 , \391 );
nand \U$340 ( \717 , RIae763e8_41, RIae76460_42);
or \U$341 ( \718 , \389 , \717 );
nand \U$342 ( \719 , RIae764d8_43, RIae76550_44);
nand \U$343 ( \720 , \718 , \719 );
not \U$344 ( \721 , \720 );
or \U$345 ( \722 , \716 , \721 );
nand \U$346 ( \723 , RIae766b8_47, RIae76730_48);
nand \U$347 ( \724 , \722 , \723 );
not \U$348 ( \725 , \724 );
or \U$349 ( \726 , \715 , \725 );
nand \U$350 ( \727 , RIae765c8_45, RIae76640_46);
nand \U$351 ( \728 , \726 , \727 );
not \U$352 ( \729 , \728 );
or \U$353 ( \730 , \714 , \729 );
not \U$354 ( \731 , \385 );
nand \U$355 ( \732 , RIae76118_35, RIae76190_36);
or \U$356 ( \733 , \382 , \732 );
nand \U$357 ( \734 , RIae76028_33, RIae760a0_34);
nand \U$358 ( \735 , \733 , \734 );
not \U$359 ( \736 , \735 );
or \U$360 ( \737 , \731 , \736 );
nand \U$361 ( \738 , RIae762f8_39, RIae76370_40);
nand \U$362 ( \739 , \737 , \738 );
and \U$363 ( \740 , \739 , \386 );
and \U$364 ( \741 , RIae76208_37, RIae76280_38);
nor \U$365 ( \742 , \740 , \741 );
nand \U$366 ( \743 , \730 , \742 );
not \U$367 ( \744 , \743 );
or \U$368 ( \745 , \713 , \744 );
not \U$369 ( \746 , \398 );
not \U$370 ( \747 , \397 );
nand \U$371 ( \748 , RIae76a78_55, RIae76af0_56);
or \U$372 ( \749 , \394 , \748 );
nand \U$373 ( \750 , RIae76988_53, RIae76a00_54);
nand \U$374 ( \751 , \749 , \750 );
not \U$375 ( \752 , \751 );
or \U$376 ( \753 , \747 , \752 );
nand \U$377 ( \754 , RIae767a8_49, RIae76820_50);
nand \U$378 ( \755 , \753 , \754 );
not \U$379 ( \756 , \755 );
or \U$380 ( \757 , \746 , \756 );
nand \U$381 ( \758 , RIae76898_51, RIae76910_52);
nand \U$382 ( \759 , \757 , \758 );
not \U$383 ( \760 , \759 );
nand \U$384 ( \761 , \745 , \760 );
not \U$385 ( \762 , \761 );
nand \U$386 ( \763 , \712 , \762 );
not \U$387 ( \764 , \763 );
or \U$388 ( \765 , \381 , \764 );
nand \U$389 ( \766 , RIae76b68_57, RIae76be0_58);
or \U$390 ( \767 , \379 , \766 );
nand \U$391 ( \768 , RIae78a58_123, RIae78ad0_124);
nand \U$392 ( \769 , \767 , \768 );
not \U$393 ( \770 , \769 );
nand \U$394 ( \771 , \765 , \770 );
or \U$395 ( \772 , RIae78cb0_128, RIae78d28_129);
nand \U$396 ( \773 , RIae78cb0_128, RIae78d28_129);
and \U$397 ( \774 , \772 , \773 );
not \U$398 ( \775 , \774 );
and \U$399 ( \776 , \771 , \775 );
not \U$400 ( \777 , \771 );
and \U$401 ( \778 , \777 , \774 );
nor \U$402 ( \779 , \776 , \778 );
buf \U$403 ( \780 , \779 );
not \U$404 ( \781 , \780 );
buf \U$405 ( \782 , \781 );
not \U$406 ( \783 , \782 );
xor \U$407 ( \784 , \783 , RIae78f80_134);
not \U$408 ( \785 , \784 );
nand \U$409 ( \786 , RIae79070_136, RIae790e8_137);
not \U$410 ( \787 , \786 );
nor \U$411 ( \788 , RIae79070_136, RIae790e8_137);
nor \U$412 ( \789 , \787 , \788 );
not \U$413 ( \790 , \789 );
and \U$414 ( \791 , RIae78f80_134, RIae790e8_137);
not \U$415 ( \792 , RIae78f80_134);
not \U$416 ( \793 , RIae790e8_137);
and \U$417 ( \794 , \792 , \793 );
nor \U$418 ( \795 , \791 , \794 );
and \U$419 ( \796 , \790 , \795 );
buf \U$420 ( \797 , \796 );
not \U$421 ( \798 , \797 );
not \U$422 ( \799 , \798 );
and \U$423 ( \800 , \785 , \799 );
and \U$424 ( \801 , \380 , \772 );
and \U$425 ( \802 , \801 , \399 );
not \U$426 ( \803 , \802 );
and \U$427 ( \804 , \387 , \393 );
not \U$428 ( \805 , \804 );
not \U$429 ( \806 , \710 );
or \U$430 ( \807 , \805 , \806 );
not \U$431 ( \808 , \743 );
nand \U$432 ( \809 , \807 , \808 );
not \U$433 ( \810 , \809 );
or \U$434 ( \811 , \803 , \810 );
nand \U$435 ( \812 , \759 , \801 );
and \U$436 ( \813 , \769 , \772 );
not \U$437 ( \814 , \773 );
nor \U$438 ( \815 , \813 , \814 );
and \U$439 ( \816 , \812 , \815 );
nand \U$440 ( \817 , \811 , \816 );
or \U$441 ( \818 , RIae78da0_130, RIae78e18_131);
nand \U$442 ( \819 , RIae78da0_130, RIae78e18_131);
nand \U$443 ( \820 , \818 , \819 );
and \U$444 ( \821 , \817 , \820 );
not \U$445 ( \822 , \817 );
not \U$446 ( \823 , \820 );
and \U$447 ( \824 , \822 , \823 );
nor \U$448 ( \825 , \821 , \824 );
not \U$449 ( \826 , \825 );
not \U$450 ( \827 , \826 );
buf \U$451 ( \828 , \827 );
buf \U$452 ( \829 , \828 );
not \U$453 ( \830 , \829 );
and \U$454 ( \831 , RIae78f80_134, \830 );
not \U$455 ( \832 , RIae78f80_134);
not \U$456 ( \833 , \825 );
not \U$457 ( \834 , \833 );
buf \U$458 ( \835 , \834 );
and \U$459 ( \836 , \832 , \835 );
nor \U$460 ( \837 , \831 , \836 );
buf \U$461 ( \838 , \789 );
buf \U$462 ( \839 , \838 );
buf \U$463 ( \840 , \839 );
and \U$464 ( \841 , \837 , \840 );
nor \U$465 ( \842 , \800 , \841 );
not \U$466 ( \843 , \395 );
not \U$467 ( \844 , \843 );
not \U$468 ( \845 , \809 );
or \U$469 ( \846 , \844 , \845 );
nand \U$470 ( \847 , \846 , \748 );
xor \U$471 ( \848 , RIae76988_53, RIae76a00_54);
and \U$472 ( \849 , \847 , \848 );
not \U$473 ( \850 , \847 );
not \U$474 ( \851 , \848 );
and \U$475 ( \852 , \850 , \851 );
nor \U$476 ( \853 , \849 , \852 );
buf \U$477 ( \854 , \853 );
not \U$478 ( \855 , \854 );
not \U$479 ( \856 , \855 );
not \U$480 ( \857 , \856 );
not \U$481 ( \858 , \857 );
nand \U$482 ( \859 , \858 , RIae78b48_125);
not \U$483 ( \860 , RIae78b48_125);
nand \U$484 ( \861 , \857 , \860 );
and \U$485 ( \862 , \859 , \861 );
nand \U$486 ( \863 , RIae78bc0_126, RIae78c38_127);
not \U$487 ( \864 , \863 );
nor \U$488 ( \865 , RIae78bc0_126, RIae78c38_127);
nor \U$489 ( \866 , \864 , \865 );
buf \U$490 ( \867 , \866 );
buf \U$491 ( \868 , \867 );
and \U$492 ( \869 , \862 , \868 );
buf \U$493 ( \870 , \809 );
not \U$494 ( \871 , \870 );
nand \U$495 ( \872 , \843 , \748 );
not \U$496 ( \873 , \872 );
and \U$497 ( \874 , \871 , \873 );
and \U$498 ( \875 , \870 , \872 );
nor \U$499 ( \876 , \874 , \875 );
buf \U$500 ( \877 , \876 );
buf \U$501 ( \878 , \877 );
buf \U$502 ( \879 , \878 );
not \U$503 ( \880 , \879 );
and \U$504 ( \881 , RIae78b48_125, \880 );
not \U$505 ( \882 , RIae78b48_125);
not \U$506 ( \883 , \877 );
not \U$507 ( \884 , \883 );
and \U$508 ( \885 , \882 , \884 );
nor \U$509 ( \886 , \881 , \885 );
or \U$510 ( \887 , RIae78b48_125, RIae78c38_127);
not \U$511 ( \888 , RIae78c38_127);
or \U$512 ( \889 , \888 , \860 );
not \U$513 ( \890 , \866 );
nand \U$514 ( \891 , \887 , \889 , \890 );
not \U$515 ( \892 , \891 );
buf \U$516 ( \893 , \892 );
and \U$517 ( \894 , \886 , \893 );
nor \U$518 ( \895 , \869 , \894 );
xnor \U$519 ( \896 , \842 , \895 );
not \U$520 ( \897 , \397 );
and \U$521 ( \898 , \387 , \393 , \396 );
not \U$522 ( \899 , \898 );
not \U$523 ( \900 , \710 );
or \U$524 ( \901 , \899 , \900 );
not \U$525 ( \902 , \396 );
not \U$526 ( \903 , \743 );
or \U$527 ( \904 , \902 , \903 );
not \U$528 ( \905 , \751 );
nand \U$529 ( \906 , \904 , \905 );
not \U$530 ( \907 , \906 );
nand \U$531 ( \908 , \901 , \907 );
not \U$532 ( \909 , \908 );
or \U$533 ( \910 , \897 , \909 );
nand \U$534 ( \911 , \910 , \754 );
nand \U$535 ( \912 , \398 , \758 );
not \U$536 ( \913 , \912 );
and \U$537 ( \914 , \911 , \913 );
not \U$538 ( \915 , \911 );
and \U$539 ( \916 , \915 , \912 );
nor \U$540 ( \917 , \914 , \916 );
buf \U$541 ( \918 , \917 );
not \U$542 ( \919 , \918 );
xnor \U$543 ( \920 , \919 , RIae78bc0_126);
not \U$544 ( \921 , RIae78e90_132);
not \U$545 ( \922 , RIae78ff8_135);
and \U$546 ( \923 , \921 , \922 );
and \U$547 ( \924 , RIae78e90_132, RIae78ff8_135);
nor \U$548 ( \925 , \923 , \924 );
buf \U$549 ( \926 , \925 );
buf \U$550 ( \927 , \926 );
not \U$551 ( \928 , \927 );
not \U$552 ( \929 , \928 );
and \U$553 ( \930 , \920 , \929 );
nand \U$554 ( \931 , \397 , \754 );
and \U$555 ( \932 , \908 , \931 );
not \U$556 ( \933 , \908 );
not \U$557 ( \934 , \931 );
and \U$558 ( \935 , \933 , \934 );
nor \U$559 ( \936 , \932 , \935 );
not \U$560 ( \937 , \936 );
not \U$561 ( \938 , \937 );
not \U$562 ( \939 , \938 );
not \U$563 ( \940 , \939 );
not \U$564 ( \941 , \940 );
and \U$565 ( \942 , RIae78bc0_126, \941 );
not \U$566 ( \943 , RIae78bc0_126);
buf \U$567 ( \944 , \940 );
and \U$568 ( \945 , \943 , \944 );
nor \U$569 ( \946 , \942 , \945 );
and \U$570 ( \947 , RIae78bc0_126, RIae78ff8_135);
nor \U$571 ( \948 , RIae78bc0_126, RIae78ff8_135);
nor \U$572 ( \949 , \947 , \925 , \948 );
not \U$573 ( \950 , \949 );
not \U$574 ( \951 , \950 );
buf \U$575 ( \952 , \951 );
buf \U$576 ( \953 , \952 );
and \U$577 ( \954 , \946 , \953 );
nor \U$578 ( \955 , \930 , \954 );
xor \U$579 ( \956 , \896 , \955 );
not \U$580 ( \957 , \956 );
not \U$581 ( \958 , \384 );
and \U$582 ( \959 , \710 , \393 );
not \U$583 ( \960 , \959 );
or \U$584 ( \961 , \958 , \960 );
not \U$585 ( \962 , \384 );
not \U$586 ( \963 , \728 );
or \U$587 ( \964 , \962 , \963 );
not \U$588 ( \965 , \735 );
nand \U$589 ( \966 , \964 , \965 );
not \U$590 ( \967 , \966 );
nand \U$591 ( \968 , \961 , \967 );
not \U$592 ( \969 , \968 );
nand \U$593 ( \970 , \385 , \738 );
not \U$594 ( \971 , \970 );
and \U$595 ( \972 , \969 , \971 );
and \U$596 ( \973 , \968 , \970 );
nor \U$597 ( \974 , \972 , \973 );
buf \U$598 ( \975 , \974 );
not \U$599 ( \976 , \975 );
not \U$600 ( \977 , \976 );
buf \U$601 ( \978 , \977 );
not \U$602 ( \979 , \978 );
nand \U$603 ( \980 , \979 , RIae78b48_125);
not \U$604 ( \981 , \980 );
not \U$605 ( \982 , \818 );
not \U$606 ( \983 , \801 );
buf \U$607 ( \984 , \763 );
not \U$608 ( \985 , \984 );
or \U$609 ( \986 , \983 , \985 );
nand \U$610 ( \987 , \986 , \815 );
not \U$611 ( \988 , \987 );
or \U$612 ( \989 , \982 , \988 );
nand \U$613 ( \990 , \989 , \819 );
buf \U$614 ( \991 , \990 );
buf \U$615 ( \992 , \991 );
not \U$616 ( \993 , \992 );
not \U$617 ( \994 , \993 );
and \U$618 ( \995 , \994 , RIae79160_138);
not \U$619 ( \996 , \994 );
not \U$620 ( \997 , RIae79160_138);
and \U$621 ( \998 , \996 , \997 );
nor \U$622 ( \999 , \995 , \998 );
xor \U$623 ( \1000 , RIae791d8_139, RIae79250_140);
not \U$624 ( \1001 , \1000 );
and \U$625 ( \1002 , RIae79160_138, RIae791d8_139);
not \U$626 ( \1003 , RIae79160_138);
not \U$627 ( \1004 , RIae791d8_139);
and \U$628 ( \1005 , \1003 , \1004 );
nor \U$629 ( \1006 , \1002 , \1005 );
and \U$630 ( \1007 , \1001 , \1006 );
buf \U$631 ( \1008 , \1007 );
buf \U$632 ( \1009 , \1008 );
buf \U$633 ( \1010 , \1009 );
nand \U$634 ( \1011 , \999 , \1010 );
buf \U$635 ( \1012 , \1000 );
buf \U$636 ( \1013 , \1012 );
nand \U$637 ( \1014 , \1013 , RIae79160_138);
and \U$638 ( \1015 , \1011 , \1014 );
not \U$639 ( \1016 , \1015 );
not \U$640 ( \1017 , \1016 );
or \U$641 ( \1018 , \981 , \1017 );
or \U$642 ( \1019 , \1016 , \980 );
nand \U$643 ( \1020 , \1018 , \1019 );
not \U$644 ( \1021 , \1020 );
not \U$645 ( \1022 , \854 );
not \U$646 ( \1023 , \1022 );
not \U$647 ( \1024 , \1023 );
xor \U$648 ( \1025 , \1024 , RIae78bc0_126);
not \U$649 ( \1026 , \1025 );
buf \U$650 ( \1027 , \926 );
buf \U$651 ( \1028 , \1027 );
not \U$652 ( \1029 , \1028 );
not \U$653 ( \1030 , \1029 );
and \U$654 ( \1031 , \1026 , \1030 );
and \U$655 ( \1032 , RIae78bc0_126, \880 );
not \U$656 ( \1033 , RIae78bc0_126);
and \U$657 ( \1034 , \1033 , \879 );
nor \U$658 ( \1035 , \1032 , \1034 );
buf \U$659 ( \1036 , \951 );
and \U$660 ( \1037 , \1035 , \1036 );
nor \U$661 ( \1038 , \1031 , \1037 );
not \U$662 ( \1039 , RIae79070_136);
and \U$663 ( \1040 , \1039 , \835 );
not \U$664 ( \1041 , \1039 );
and \U$665 ( \1042 , \1041 , \830 );
nor \U$666 ( \1043 , \1040 , \1042 );
and \U$667 ( \1044 , RIae79160_138, RIae792c8_141);
not \U$668 ( \1045 , RIae79160_138);
not \U$669 ( \1046 , RIae792c8_141);
and \U$670 ( \1047 , \1045 , \1046 );
nor \U$671 ( \1048 , \1044 , \1047 );
buf \U$672 ( \1049 , \1048 );
and \U$673 ( \1050 , \1043 , \1049 );
not \U$674 ( \1051 , \782 );
not \U$675 ( \1052 , RIae79070_136);
and \U$676 ( \1053 , \1051 , \1052 );
and \U$677 ( \1054 , \782 , RIae79070_136);
nor \U$678 ( \1055 , \1053 , \1054 );
nand \U$679 ( \1056 , RIae79160_138, RIae792c8_141);
and \U$680 ( \1057 , \1039 , \1056 );
not \U$681 ( \1058 , \1039 );
nand \U$682 ( \1059 , \997 , \1046 );
and \U$683 ( \1060 , \1058 , \1059 );
nor \U$684 ( \1061 , \1057 , \1060 );
buf \U$685 ( \1062 , \1061 );
and \U$686 ( \1063 , \1055 , \1062 );
nor \U$687 ( \1064 , \1050 , \1063 );
xor \U$688 ( \1065 , \1038 , \1064 );
not \U$689 ( \1066 , RIae78e90_132);
and \U$690 ( \1067 , \919 , \1066 );
not \U$691 ( \1068 , \919 );
and \U$692 ( \1069 , \1068 , RIae78e90_132);
nor \U$693 ( \1070 , \1067 , \1069 );
xor \U$694 ( \1071 , RIae78f08_133, RIae78f80_134);
buf \U$695 ( \1072 , \1071 );
not \U$696 ( \1073 , \1072 );
not \U$697 ( \1074 , \1073 );
and \U$698 ( \1075 , \1070 , \1074 );
and \U$699 ( \1076 , \944 , \921 );
not \U$700 ( \1077 , \944 );
and \U$701 ( \1078 , \1077 , RIae78e90_132);
nor \U$702 ( \1079 , \1076 , \1078 );
not \U$703 ( \1080 , \1071 );
and \U$704 ( \1081 , RIae78e90_132, RIae78f08_133);
not \U$705 ( \1082 , RIae78e90_132);
not \U$706 ( \1083 , RIae78f08_133);
and \U$707 ( \1084 , \1082 , \1083 );
nor \U$708 ( \1085 , \1081 , \1084 );
and \U$709 ( \1086 , \1080 , \1085 );
buf \U$710 ( \1087 , \1086 );
and \U$711 ( \1088 , \1079 , \1087 );
nor \U$712 ( \1089 , \1075 , \1088 );
and \U$713 ( \1090 , \1065 , \1089 );
and \U$714 ( \1091 , \1038 , \1064 );
nor \U$715 ( \1092 , \1090 , \1091 );
not \U$716 ( \1093 , \1092 );
or \U$717 ( \1094 , \1021 , \1093 );
or \U$718 ( \1095 , \1015 , \980 );
nand \U$719 ( \1096 , \1094 , \1095 );
not \U$720 ( \1097 , \1096 );
or \U$721 ( \1098 , \957 , \1097 );
not \U$722 ( \1099 , \741 );
nand \U$723 ( \1100 , \1099 , \386 );
not \U$724 ( \1101 , \1100 );
not \U$725 ( \1102 , \1101 );
and \U$726 ( \1103 , \384 , \385 );
not \U$727 ( \1104 , \1103 );
not \U$728 ( \1105 , \959 );
or \U$729 ( \1106 , \1104 , \1105 );
not \U$730 ( \1107 , \385 );
not \U$731 ( \1108 , \966 );
or \U$732 ( \1109 , \1107 , \1108 );
nand \U$733 ( \1110 , \1109 , \738 );
not \U$734 ( \1111 , \1110 );
nand \U$735 ( \1112 , \1106 , \1111 );
not \U$736 ( \1113 , \1112 );
not \U$737 ( \1114 , \1113 );
or \U$738 ( \1115 , \1102 , \1114 );
nand \U$739 ( \1116 , \1112 , \1100 );
nand \U$740 ( \1117 , \1115 , \1116 );
buf \U$741 ( \1118 , \1117 );
not \U$742 ( \1119 , \1118 );
not \U$743 ( \1120 , \1119 );
xor \U$744 ( \1121 , RIae78b48_125, \1120 );
buf \U$745 ( \1122 , \868 );
and \U$746 ( \1123 , \1121 , \1122 );
not \U$747 ( \1124 , \974 );
not \U$748 ( \1125 , \1124 );
nand \U$749 ( \1126 , \1125 , \860 );
and \U$750 ( \1127 , \980 , \1126 );
not \U$751 ( \1128 , \892 );
not \U$752 ( \1129 , \1128 );
and \U$753 ( \1130 , \1127 , \1129 );
nor \U$754 ( \1131 , \1123 , \1130 );
not \U$755 ( \1132 , RIae78f80_134);
not \U$756 ( \1133 , \378 );
not \U$757 ( \1134 , \1133 );
not \U$758 ( \1135 , \763 );
or \U$759 ( \1136 , \1134 , \1135 );
nand \U$760 ( \1137 , \1136 , \766 );
not \U$761 ( \1138 , \379 );
nand \U$762 ( \1139 , \1138 , \768 );
xnor \U$763 ( \1140 , \1137 , \1139 );
buf \U$764 ( \1141 , \1140 );
not \U$765 ( \1142 , \1141 );
buf \U$766 ( \1143 , \1142 );
and \U$767 ( \1144 , \1132 , \1143 );
not \U$768 ( \1145 , \1132 );
not \U$769 ( \1146 , \1141 );
not \U$770 ( \1147 , \1146 );
and \U$771 ( \1148 , \1145 , \1147 );
nor \U$772 ( \1149 , \1144 , \1148 );
and \U$773 ( \1150 , \1149 , \840 );
not \U$774 ( \1151 , \763 );
nand \U$775 ( \1152 , \1133 , \766 );
not \U$776 ( \1153 , \1152 );
and \U$777 ( \1154 , \1151 , \1153 );
and \U$778 ( \1155 , \984 , \1152 );
nor \U$779 ( \1156 , \1154 , \1155 );
not \U$780 ( \1157 , \1156 );
not \U$781 ( \1158 , \1157 );
not \U$782 ( \1159 , \1158 );
and \U$783 ( \1160 , RIae78f80_134, \1159 );
not \U$784 ( \1161 , RIae78f80_134);
not \U$785 ( \1162 , \1159 );
and \U$786 ( \1163 , \1161 , \1162 );
nor \U$787 ( \1164 , \1160 , \1163 );
and \U$788 ( \1165 , \1164 , \797 );
nor \U$789 ( \1166 , \1150 , \1165 );
not \U$790 ( \1167 , \383 );
not \U$791 ( \1168 , \1167 );
not \U$792 ( \1169 , \393 );
and \U$793 ( \1170 , \674 , \708 );
nand \U$794 ( \1171 , \643 , \1170 );
not \U$795 ( \1172 , \1171 );
or \U$796 ( \1173 , \1169 , \1172 );
not \U$797 ( \1174 , \728 );
nand \U$798 ( \1175 , \1173 , \1174 );
not \U$799 ( \1176 , \1175 );
or \U$800 ( \1177 , \1168 , \1176 );
nand \U$801 ( \1178 , \1177 , \732 );
not \U$802 ( \1179 , \382 );
nand \U$803 ( \1180 , \1179 , \734 );
and \U$804 ( \1181 , \1178 , \1180 );
not \U$805 ( \1182 , \1178 );
not \U$806 ( \1183 , \1180 );
and \U$807 ( \1184 , \1182 , \1183 );
nor \U$808 ( \1185 , \1181 , \1184 );
buf \U$809 ( \1186 , \1185 );
buf \U$810 ( \1187 , \1186 );
not \U$811 ( \1188 , \1187 );
nand \U$812 ( \1189 , \1188 , RIae78b48_125);
xnor \U$813 ( \1190 , \1166 , \1189 );
or \U$814 ( \1191 , \1131 , \1190 );
or \U$815 ( \1192 , \1166 , \1189 );
nand \U$816 ( \1193 , \1191 , \1192 );
not \U$817 ( \1194 , \991 );
buf \U$818 ( \1195 , \1194 );
not \U$819 ( \1196 , \1195 );
buf \U$820 ( \1197 , \1196 );
and \U$821 ( \1198 , \1197 , \1039 );
not \U$822 ( \1199 , \1197 );
and \U$823 ( \1200 , \1199 , RIae79070_136);
nor \U$824 ( \1201 , \1198 , \1200 );
not \U$825 ( \1202 , \1201 );
not \U$826 ( \1203 , \1049 );
not \U$827 ( \1204 , \1203 );
and \U$828 ( \1205 , \1202 , \1204 );
and \U$829 ( \1206 , \1043 , \1062 );
nor \U$830 ( \1207 , \1205 , \1206 );
not \U$831 ( \1208 , \1009 );
buf \U$832 ( \1209 , \1012 );
not \U$833 ( \1210 , \1209 );
and \U$834 ( \1211 , \1208 , \1210 );
nor \U$835 ( \1212 , \1211 , \997 );
xnor \U$836 ( \1213 , \1207 , \1212 );
and \U$837 ( \1214 , RIae78e90_132, \1159 );
not \U$838 ( \1215 , RIae78e90_132);
and \U$839 ( \1216 , \1215 , \1162 );
nor \U$840 ( \1217 , \1214 , \1216 );
and \U$841 ( \1218 , \1217 , \1074 );
and \U$842 ( \1219 , \1070 , \1087 );
nor \U$843 ( \1220 , \1218 , \1219 );
xor \U$844 ( \1221 , \1213 , \1220 );
xor \U$845 ( \1222 , \1193 , \1221 );
and \U$846 ( \1223 , \886 , \1122 );
and \U$847 ( \1224 , \1121 , \1129 );
nor \U$848 ( \1225 , \1223 , \1224 );
not \U$849 ( \1226 , \784 );
not \U$850 ( \1227 , \840 );
not \U$851 ( \1228 , \1227 );
and \U$852 ( \1229 , \1226 , \1228 );
and \U$853 ( \1230 , \1149 , \797 );
nor \U$854 ( \1231 , \1229 , \1230 );
not \U$855 ( \1232 , \1025 );
not \U$856 ( \1233 , \953 );
not \U$857 ( \1234 , \1233 );
and \U$858 ( \1235 , \1232 , \1234 );
and \U$859 ( \1236 , \946 , \929 );
nor \U$860 ( \1237 , \1235 , \1236 );
xnor \U$861 ( \1238 , \1231 , \1237 );
xor \U$862 ( \1239 , \1225 , \1238 );
and \U$863 ( \1240 , \1222 , \1239 );
and \U$864 ( \1241 , \1193 , \1221 );
nor \U$865 ( \1242 , \1240 , \1241 );
not \U$866 ( \1243 , \1242 );
xor \U$867 ( \1244 , \956 , \1096 );
nand \U$868 ( \1245 , \1243 , \1244 );
nand \U$869 ( \1246 , \1098 , \1245 );
and \U$870 ( \1247 , RIae78b48_125, \1120 );
not \U$871 ( \1248 , \1201 );
not \U$872 ( \1249 , \1062 );
not \U$873 ( \1250 , \1249 );
and \U$874 ( \1251 , \1248 , \1250 );
and \U$875 ( \1252 , \1049 , RIae79070_136);
nor \U$876 ( \1253 , \1251 , \1252 );
and \U$877 ( \1254 , \1247 , \1253 );
not \U$878 ( \1255 , \1247 );
not \U$879 ( \1256 , \1253 );
and \U$880 ( \1257 , \1255 , \1256 );
nor \U$881 ( \1258 , \1254 , \1257 );
buf \U$882 ( \1259 , \1086 );
not \U$883 ( \1260 , \1259 );
not \U$884 ( \1261 , \1217 );
or \U$885 ( \1262 , \1260 , \1261 );
xnor \U$886 ( \1263 , \1147 , RIae78e90_132);
or \U$887 ( \1264 , \1263 , \1073 );
nand \U$888 ( \1265 , \1262 , \1264 );
xor \U$889 ( \1266 , \1258 , \1265 );
or \U$890 ( \1267 , \1213 , \1220 );
or \U$891 ( \1268 , \1207 , \1212 );
nand \U$892 ( \1269 , \1267 , \1268 );
and \U$893 ( \1270 , \1266 , \1269 );
xor \U$894 ( \1271 , \1266 , \1269 );
or \U$895 ( \1272 , \1238 , \1225 );
or \U$896 ( \1273 , \1231 , \1237 );
nand \U$897 ( \1274 , \1272 , \1273 );
and \U$898 ( \1275 , \1271 , \1274 );
nor \U$899 ( \1276 , \1270 , \1275 );
and \U$900 ( \1277 , \1246 , \1276 );
not \U$901 ( \1278 , \1246 );
not \U$902 ( \1279 , \1276 );
and \U$903 ( \1280 , \1278 , \1279 );
nor \U$904 ( \1281 , \1277 , \1280 );
not \U$905 ( \1282 , \1281 );
and \U$906 ( \1283 , \1258 , \1265 );
and \U$907 ( \1284 , \1253 , \1247 );
nor \U$908 ( \1285 , \1283 , \1284 );
not \U$909 ( \1286 , RIae78bc0_126);
and \U$910 ( \1287 , \1162 , \1286 );
buf \U$911 ( \1288 , \1156 );
not \U$912 ( \1289 , \1288 );
not \U$913 ( \1290 , \1289 );
not \U$914 ( \1291 , \1290 );
and \U$915 ( \1292 , \1291 , RIae78bc0_126);
nor \U$916 ( \1293 , \1287 , \1292 );
and \U$917 ( \1294 , \1293 , \1027 );
and \U$918 ( \1295 , \920 , \953 );
nor \U$919 ( \1296 , \1294 , \1295 );
and \U$920 ( \1297 , \1056 , RIae79070_136);
xor \U$921 ( \1298 , \1296 , \1297 );
and \U$922 ( \1299 , \837 , \797 );
xor \U$923 ( \1300 , \994 , RIae78f80_134);
and \U$924 ( \1301 , \1300 , \840 );
nor \U$925 ( \1302 , \1299 , \1301 );
xor \U$926 ( \1303 , \1298 , \1302 );
xor \U$927 ( \1304 , \1285 , \1303 );
or \U$928 ( \1305 , \896 , \955 );
or \U$929 ( \1306 , \895 , \842 );
nand \U$930 ( \1307 , \1305 , \1306 );
and \U$931 ( \1308 , \1307 , \1256 );
not \U$932 ( \1309 , \1307 );
and \U$933 ( \1310 , \1309 , \1253 );
nor \U$934 ( \1311 , \1308 , \1310 );
not \U$935 ( \1312 , \1263 );
not \U$936 ( \1313 , \1087 );
not \U$937 ( \1314 , \1313 );
and \U$938 ( \1315 , \1312 , \1314 );
and \U$939 ( \1316 , \1066 , \783 );
not \U$940 ( \1317 , \1066 );
and \U$941 ( \1318 , \1317 , \782 );
nor \U$942 ( \1319 , \1316 , \1318 );
buf \U$943 ( \1320 , \1072 );
buf \U$944 ( \1321 , \1320 );
buf \U$945 ( \1322 , \1321 );
and \U$946 ( \1323 , \1319 , \1322 );
nor \U$947 ( \1324 , \1315 , \1323 );
nand \U$948 ( \1325 , \880 , RIae78b48_125);
xnor \U$949 ( \1326 , \1324 , \1325 );
and \U$950 ( \1327 , \944 , \860 );
and \U$951 ( \1328 , \941 , RIae78b48_125);
nor \U$952 ( \1329 , \1327 , \1328 );
and \U$953 ( \1330 , \1329 , \1122 );
and \U$954 ( \1331 , \862 , \1129 );
nor \U$955 ( \1332 , \1330 , \1331 );
xor \U$956 ( \1333 , \1326 , \1332 );
xnor \U$957 ( \1334 , \1311 , \1333 );
xor \U$958 ( \1335 , \1304 , \1334 );
not \U$959 ( \1336 , \1335 );
and \U$960 ( \1337 , \1282 , \1336 );
and \U$961 ( \1338 , \1246 , \1279 );
nor \U$962 ( \1339 , \1337 , \1338 );
and \U$963 ( \1340 , RIae78e90_132, \830 );
not \U$964 ( \1341 , RIae78e90_132);
and \U$965 ( \1342 , \1341 , \829 );
nor \U$966 ( \1343 , \1340 , \1342 );
and \U$967 ( \1344 , \1343 , \1322 );
and \U$968 ( \1345 , \1319 , \1087 );
nor \U$969 ( \1346 , \1344 , \1345 );
xnor \U$970 ( \1347 , \1346 , \859 );
and \U$971 ( \1348 , \919 , \860 );
and \U$972 ( \1349 , \1068 , RIae78b48_125);
nor \U$973 ( \1350 , \1348 , \1349 );
and \U$974 ( \1351 , \1350 , \1122 );
and \U$975 ( \1352 , \1329 , \1129 );
nor \U$976 ( \1353 , \1351 , \1352 );
xor \U$977 ( \1354 , \1347 , \1353 );
xor \U$978 ( \1355 , \1296 , \1297 );
and \U$979 ( \1356 , \1355 , \1302 );
and \U$980 ( \1357 , \1296 , \1297 );
nor \U$981 ( \1358 , \1356 , \1357 );
xor \U$982 ( \1359 , \1354 , \1358 );
or \U$983 ( \1360 , \1326 , \1332 );
or \U$984 ( \1361 , \1324 , \1325 );
nand \U$985 ( \1362 , \1360 , \1361 );
nand \U$986 ( \1363 , \1300 , \797 );
nand \U$987 ( \1364 , \840 , RIae78f80_134);
and \U$988 ( \1365 , \1363 , \1364 );
not \U$989 ( \1366 , \1143 );
and \U$990 ( \1367 , RIae78bc0_126, \1366 );
not \U$991 ( \1368 , RIae78bc0_126);
and \U$992 ( \1369 , \1368 , \1143 );
nor \U$993 ( \1370 , \1367 , \1369 );
and \U$994 ( \1371 , \1370 , \929 );
and \U$995 ( \1372 , \1293 , \953 );
nor \U$996 ( \1373 , \1371 , \1372 );
not \U$997 ( \1374 , \1373 );
and \U$998 ( \1375 , \1365 , \1374 );
not \U$999 ( \1376 , \1365 );
and \U$1000 ( \1377 , \1376 , \1373 );
nor \U$1001 ( \1378 , \1375 , \1377 );
xor \U$1002 ( \1379 , \1362 , \1378 );
xnor \U$1003 ( \1380 , \1359 , \1379 );
and \U$1004 ( \1381 , \1307 , \1256 );
and \U$1005 ( \1382 , \1311 , \1333 );
nor \U$1006 ( \1383 , \1381 , \1382 );
xor \U$1007 ( \1384 , \1380 , \1383 );
xor \U$1008 ( \1385 , \1285 , \1303 );
and \U$1009 ( \1386 , \1385 , \1334 );
and \U$1010 ( \1387 , \1285 , \1303 );
or \U$1011 ( \1388 , \1386 , \1387 );
xor \U$1012 ( \1389 , \1384 , \1388 );
nand \U$1013 ( \1390 , \1339 , \1389 );
not \U$1014 ( \1391 , \1049 );
not \U$1015 ( \1392 , \1055 );
or \U$1016 ( \1393 , \1391 , \1392 );
xnor \U$1017 ( \1394 , \1143 , RIae79070_136);
nand \U$1018 ( \1395 , \1394 , \1062 );
nand \U$1019 ( \1396 , \1393 , \1395 );
buf \U$1020 ( \1397 , \1175 );
nand \U$1021 ( \1398 , \1167 , \732 );
not \U$1022 ( \1399 , \1398 );
and \U$1023 ( \1400 , \1397 , \1399 );
not \U$1024 ( \1401 , \1397 );
and \U$1025 ( \1402 , \1401 , \1398 );
nor \U$1026 ( \1403 , \1400 , \1402 );
buf \U$1027 ( \1404 , \1403 );
not \U$1028 ( \1405 , \1404 );
not \U$1029 ( \1406 , \1405 );
and \U$1030 ( \1407 , RIae78b48_125, \1406 );
xor \U$1031 ( \1408 , \1396 , \1407 );
not \U$1032 ( \1409 , \1322 );
not \U$1033 ( \1410 , \1079 );
or \U$1034 ( \1411 , \1409 , \1410 );
xor \U$1035 ( \1412 , RIae78e90_132, \857 );
not \U$1036 ( \1413 , \1259 );
or \U$1037 ( \1414 , \1412 , \1413 );
nand \U$1038 ( \1415 , \1411 , \1414 );
and \U$1039 ( \1416 , \1408 , \1415 );
and \U$1040 ( \1417 , \1396 , \1407 );
nor \U$1041 ( \1418 , \1416 , \1417 );
not \U$1042 ( \1419 , \1418 );
not \U$1043 ( \1420 , \1419 );
not \U$1044 ( \1421 , \1013 );
not \U$1045 ( \1422 , \999 );
or \U$1046 ( \1423 , \1421 , \1422 );
not \U$1047 ( \1424 , \835 );
not \U$1048 ( \1425 , \1424 );
not \U$1049 ( \1426 , RIae79160_138);
and \U$1050 ( \1427 , \1425 , \1426 );
and \U$1051 ( \1428 , \830 , RIae79160_138);
nor \U$1052 ( \1429 , \1427 , \1428 );
buf \U$1053 ( \1430 , \1009 );
nand \U$1054 ( \1431 , \1429 , \1430 );
nand \U$1055 ( \1432 , \1423 , \1431 );
not \U$1056 ( \1433 , \1432 );
nand \U$1057 ( \1434 , RIae79340_142, RIae793b8_143);
and \U$1058 ( \1435 , \1434 , RIae79250_140);
or \U$1059 ( \1436 , \1433 , \1435 );
and \U$1060 ( \1437 , \1164 , \840 );
not \U$1061 ( \1438 , \917 );
buf \U$1062 ( \1439 , \1438 );
buf \U$1063 ( \1440 , \1439 );
not \U$1064 ( \1441 , \1440 );
and \U$1065 ( \1442 , RIae78f80_134, \1441 );
not \U$1066 ( \1443 , RIae78f80_134);
and \U$1067 ( \1444 , \1443 , \919 );
nor \U$1068 ( \1445 , \1442 , \1444 );
and \U$1069 ( \1446 , \1445 , \797 );
nor \U$1070 ( \1447 , \1437 , \1446 );
not \U$1071 ( \1448 , \1447 );
not \U$1072 ( \1449 , \1435 );
not \U$1073 ( \1450 , \1432 );
or \U$1074 ( \1451 , \1449 , \1450 );
or \U$1075 ( \1452 , \1432 , \1435 );
nand \U$1076 ( \1453 , \1451 , \1452 );
nand \U$1077 ( \1454 , \1448 , \1453 );
nand \U$1078 ( \1455 , \1436 , \1454 );
and \U$1079 ( \1456 , \1455 , \1015 );
not \U$1080 ( \1457 , \1455 );
and \U$1081 ( \1458 , \1457 , \1016 );
nor \U$1082 ( \1459 , \1456 , \1458 );
not \U$1083 ( \1460 , \1459 );
or \U$1084 ( \1461 , \1420 , \1460 );
nand \U$1085 ( \1462 , \1455 , \1015 );
nand \U$1086 ( \1463 , \1461 , \1462 );
not \U$1087 ( \1464 , \1463 );
xnor \U$1088 ( \1465 , \1092 , \1020 );
or \U$1089 ( \1466 , \1464 , \1465 );
not \U$1090 ( \1467 , \1463 );
not \U$1091 ( \1468 , \1465 );
and \U$1092 ( \1469 , \1467 , \1468 );
and \U$1093 ( \1470 , \1463 , \1465 );
nor \U$1094 ( \1471 , \1469 , \1470 );
not \U$1095 ( \1472 , \1118 );
not \U$1096 ( \1473 , \1472 );
and \U$1097 ( \1474 , RIae78bc0_126, \1473 );
not \U$1098 ( \1475 , RIae78bc0_126);
and \U$1099 ( \1476 , \1475 , \1119 );
nor \U$1100 ( \1477 , \1474 , \1476 );
not \U$1101 ( \1478 , \1477 );
not \U$1102 ( \1479 , \1478 );
not \U$1103 ( \1480 , \1233 );
and \U$1104 ( \1481 , \1479 , \1480 );
and \U$1105 ( \1482 , \1035 , \1027 );
nor \U$1106 ( \1483 , \1481 , \1482 );
not \U$1107 ( \1484 , \1197 );
not \U$1108 ( \1485 , RIae79250_140);
and \U$1109 ( \1486 , \1484 , \1485 );
and \U$1110 ( \1487 , \994 , RIae79250_140);
nor \U$1111 ( \1488 , \1486 , \1487 );
xor \U$1112 ( \1489 , RIae79340_142, RIae793b8_143);
not \U$1113 ( \1490 , \1489 );
and \U$1114 ( \1491 , RIae79250_140, RIae79340_142);
not \U$1115 ( \1492 , RIae79250_140);
not \U$1116 ( \1493 , RIae79340_142);
and \U$1117 ( \1494 , \1492 , \1493 );
nor \U$1118 ( \1495 , \1491 , \1494 );
nand \U$1119 ( \1496 , \1490 , \1495 );
not \U$1120 ( \1497 , \1496 );
not \U$1121 ( \1498 , \1497 );
not \U$1122 ( \1499 , \1498 );
and \U$1123 ( \1500 , \1488 , \1499 );
buf \U$1124 ( \1501 , \1489 );
not \U$1125 ( \1502 , \1501 );
not \U$1126 ( \1503 , RIae79250_140);
nor \U$1127 ( \1504 , \1502 , \1503 );
nor \U$1128 ( \1505 , \1500 , \1504 );
not \U$1129 ( \1506 , \1505 );
and \U$1130 ( \1507 , \1483 , \1506 );
not \U$1131 ( \1508 , \1483 );
and \U$1132 ( \1509 , \1508 , \1505 );
nor \U$1133 ( \1510 , \1507 , \1509 );
and \U$1134 ( \1511 , \1127 , \1122 );
xor \U$1135 ( \1512 , \1188 , RIae78b48_125);
and \U$1136 ( \1513 , \1512 , \1129 );
nor \U$1137 ( \1514 , \1511 , \1513 );
or \U$1138 ( \1515 , \1510 , \1514 );
or \U$1139 ( \1516 , \1483 , \1505 );
nand \U$1140 ( \1517 , \1515 , \1516 );
xor \U$1141 ( \1518 , \1190 , \1131 );
xor \U$1142 ( \1519 , \1517 , \1518 );
xor \U$1143 ( \1520 , \1038 , \1064 );
xor \U$1144 ( \1521 , \1520 , \1089 );
not \U$1145 ( \1522 , \1521 );
and \U$1146 ( \1523 , \1519 , \1522 );
and \U$1147 ( \1524 , \1517 , \1518 );
nor \U$1148 ( \1525 , \1523 , \1524 );
or \U$1149 ( \1526 , \1471 , \1525 );
nand \U$1150 ( \1527 , \1466 , \1526 );
xor \U$1151 ( \1528 , \1271 , \1274 );
not \U$1152 ( \1529 , \1528 );
not \U$1153 ( \1530 , \1242 );
not \U$1154 ( \1531 , \1244 );
and \U$1155 ( \1532 , \1530 , \1531 );
and \U$1156 ( \1533 , \1242 , \1244 );
nor \U$1157 ( \1534 , \1532 , \1533 );
nand \U$1158 ( \1535 , \1529 , \1534 );
and \U$1159 ( \1536 , \1527 , \1535 );
not \U$1160 ( \1537 , \1534 );
and \U$1161 ( \1538 , \1537 , \1528 );
nor \U$1162 ( \1539 , \1536 , \1538 );
xnor \U$1163 ( \1540 , \1281 , \1335 );
nand \U$1164 ( \1541 , \1539 , \1540 );
and \U$1165 ( \1542 , \1390 , \1541 );
xor \U$1166 ( \1543 , \1380 , \1383 );
and \U$1167 ( \1544 , \1543 , \1388 );
and \U$1168 ( \1545 , \1380 , \1383 );
or \U$1169 ( \1546 , \1544 , \1545 );
not \U$1170 ( \1547 , \1328 );
xnor \U$1171 ( \1548 , \1365 , \1547 );
xnor \U$1172 ( \1549 , \783 , RIae78bc0_126);
and \U$1173 ( \1550 , \1549 , \929 );
and \U$1174 ( \1551 , \1370 , \953 );
nor \U$1175 ( \1552 , \1550 , \1551 );
xor \U$1176 ( \1553 , \1548 , \1552 );
or \U$1177 ( \1554 , \1347 , \1353 );
or \U$1178 ( \1555 , \1346 , \859 );
nand \U$1179 ( \1556 , \1554 , \1555 );
xor \U$1180 ( \1557 , \1553 , \1556 );
and \U$1181 ( \1558 , \1343 , \1259 );
xor \U$1182 ( \1559 , \1197 , RIae78e90_132);
and \U$1183 ( \1560 , \1559 , \1074 );
nor \U$1184 ( \1561 , \1558 , \1560 );
and \U$1185 ( \1562 , \798 , \1227 );
nor \U$1186 ( \1563 , \1562 , \1132 );
xnor \U$1187 ( \1564 , \1561 , \1563 );
and \U$1188 ( \1565 , \1290 , \860 );
nor \U$1189 ( \1566 , \1290 , \860 );
nor \U$1190 ( \1567 , \1565 , \1566 );
and \U$1191 ( \1568 , \1567 , \1122 );
and \U$1192 ( \1569 , \1350 , \1129 );
nor \U$1193 ( \1570 , \1568 , \1569 );
xor \U$1194 ( \1571 , \1564 , \1570 );
xnor \U$1195 ( \1572 , \1557 , \1571 );
and \U$1196 ( \1573 , \1362 , \1378 );
and \U$1197 ( \1574 , \1365 , \1374 );
nor \U$1198 ( \1575 , \1573 , \1574 );
xor \U$1199 ( \1576 , \1572 , \1575 );
and \U$1200 ( \1577 , \1354 , \1358 );
and \U$1201 ( \1578 , \1359 , \1379 );
nor \U$1202 ( \1579 , \1577 , \1578 );
xor \U$1203 ( \1580 , \1576 , \1579 );
nand \U$1204 ( \1581 , \1546 , \1580 );
and \U$1205 ( \1582 , \1542 , \1581 );
or \U$1206 ( \1583 , \1564 , \1570 );
or \U$1207 ( \1584 , \1561 , \1563 );
nand \U$1208 ( \1585 , \1583 , \1584 );
and \U$1209 ( \1586 , \1559 , \1259 );
and \U$1210 ( \1587 , \1322 , RIae78e90_132);
nor \U$1211 ( \1588 , \1586 , \1587 );
and \U$1212 ( \1589 , \1585 , \1588 );
not \U$1213 ( \1590 , \1585 );
not \U$1214 ( \1591 , \1588 );
and \U$1215 ( \1592 , \1590 , \1591 );
nor \U$1216 ( \1593 , \1589 , \1592 );
or \U$1217 ( \1594 , \1548 , \1552 );
or \U$1218 ( \1595 , \1365 , \1547 );
nand \U$1219 ( \1596 , \1594 , \1595 );
xnor \U$1220 ( \1597 , \1593 , \1596 );
or \U$1221 ( \1598 , \1366 , RIae78b48_125);
and \U$1222 ( \1599 , \1366 , RIae78b48_125);
not \U$1223 ( \1600 , \1599 );
nand \U$1224 ( \1601 , \1598 , \1600 );
not \U$1225 ( \1602 , \1601 );
not \U$1226 ( \1603 , \1122 );
not \U$1227 ( \1604 , \1603 );
and \U$1228 ( \1605 , \1602 , \1604 );
and \U$1229 ( \1606 , \1567 , \1129 );
nor \U$1230 ( \1607 , \1605 , \1606 );
not \U$1231 ( \1608 , \1349 );
xor \U$1232 ( \1609 , \1607 , \1608 );
xnor \U$1233 ( \1610 , \829 , RIae78bc0_126);
and \U$1234 ( \1611 , \1610 , \929 );
and \U$1235 ( \1612 , \1549 , \953 );
nor \U$1236 ( \1613 , \1611 , \1612 );
xor \U$1237 ( \1614 , \1609 , \1613 );
xor \U$1238 ( \1615 , \1597 , \1614 );
and \U$1239 ( \1616 , \1553 , \1556 );
and \U$1240 ( \1617 , \1557 , \1571 );
nor \U$1241 ( \1618 , \1616 , \1617 );
xor \U$1242 ( \1619 , \1615 , \1618 );
xor \U$1243 ( \1620 , \1572 , \1575 );
and \U$1244 ( \1621 , \1620 , \1579 );
and \U$1245 ( \1622 , \1572 , \1575 );
or \U$1246 ( \1623 , \1621 , \1622 );
nand \U$1247 ( \1624 , \1619 , \1623 );
and \U$1248 ( \1625 , \1582 , \1624 );
xor \U$1249 ( \1626 , \1607 , \1608 );
and \U$1250 ( \1627 , \1626 , \1613 );
and \U$1251 ( \1628 , \1607 , \1608 );
nor \U$1252 ( \1629 , \1627 , \1628 );
or \U$1253 ( \1630 , \782 , RIae78b48_125);
nand \U$1254 ( \1631 , \782 , RIae78b48_125);
nand \U$1255 ( \1632 , \1630 , \1631 );
or \U$1256 ( \1633 , \1632 , \1603 );
or \U$1257 ( \1634 , \1601 , \1128 );
nand \U$1258 ( \1635 , \1633 , \1634 );
and \U$1259 ( \1636 , \1635 , \1591 );
not \U$1260 ( \1637 , \1635 );
and \U$1261 ( \1638 , \1637 , \1588 );
nor \U$1262 ( \1639 , \1636 , \1638 );
xnor \U$1263 ( \1640 , \1629 , \1639 );
and \U$1264 ( \1641 , \1610 , \953 );
xor \U$1265 ( \1642 , \1197 , RIae78bc0_126);
and \U$1266 ( \1643 , \1642 , \929 );
nor \U$1267 ( \1644 , \1641 , \1643 );
not \U$1268 ( \1645 , \1566 );
not \U$1269 ( \1646 , \1322 );
and \U$1270 ( \1647 , \1413 , \1646 );
nor \U$1271 ( \1648 , \1647 , \1066 );
xnor \U$1272 ( \1649 , \1645 , \1648 );
xnor \U$1273 ( \1650 , \1644 , \1649 );
xor \U$1274 ( \1651 , \1640 , \1650 );
and \U$1275 ( \1652 , \1593 , \1596 );
and \U$1276 ( \1653 , \1585 , \1588 );
nor \U$1277 ( \1654 , \1652 , \1653 );
xor \U$1278 ( \1655 , \1651 , \1654 );
xor \U$1279 ( \1656 , \1597 , \1614 );
and \U$1280 ( \1657 , \1656 , \1618 );
and \U$1281 ( \1658 , \1597 , \1614 );
or \U$1282 ( \1659 , \1657 , \1658 );
nand \U$1283 ( \1660 , \1655 , \1659 );
not \U$1284 ( \1661 , \1660 );
xor \U$1285 ( \1662 , \1640 , \1650 );
and \U$1286 ( \1663 , \1662 , \1654 );
and \U$1287 ( \1664 , \1640 , \1650 );
or \U$1288 ( \1665 , \1663 , \1664 );
not \U$1289 ( \1666 , \1665 );
and \U$1290 ( \1667 , \1642 , \953 );
and \U$1291 ( \1668 , \929 , RIae78bc0_126);
nor \U$1292 ( \1669 , \1667 , \1668 );
xor \U$1293 ( \1670 , \1669 , \1599 );
not \U$1294 ( \1671 , \1122 );
and \U$1295 ( \1672 , \829 , \860 );
nand \U$1296 ( \1673 , \830 , RIae78b48_125);
not \U$1297 ( \1674 , \1673 );
nor \U$1298 ( \1675 , \1672 , \1674 );
not \U$1299 ( \1676 , \1675 );
or \U$1300 ( \1677 , \1671 , \1676 );
or \U$1301 ( \1678 , \1632 , \1128 );
nand \U$1302 ( \1679 , \1677 , \1678 );
xor \U$1303 ( \1680 , \1670 , \1679 );
not \U$1304 ( \1681 , \1680 );
and \U$1305 ( \1682 , \1629 , \1639 );
and \U$1306 ( \1683 , \1635 , \1591 );
nor \U$1307 ( \1684 , \1682 , \1683 );
not \U$1308 ( \1685 , \1684 );
or \U$1309 ( \1686 , \1644 , \1649 );
or \U$1310 ( \1687 , \1645 , \1648 );
nand \U$1311 ( \1688 , \1686 , \1687 );
not \U$1312 ( \1689 , \1688 );
and \U$1313 ( \1690 , \1685 , \1689 );
and \U$1314 ( \1691 , \1684 , \1688 );
nor \U$1315 ( \1692 , \1690 , \1691 );
not \U$1316 ( \1693 , \1692 );
or \U$1317 ( \1694 , \1681 , \1693 );
or \U$1318 ( \1695 , \1692 , \1680 );
nand \U$1319 ( \1696 , \1694 , \1695 );
nor \U$1320 ( \1697 , \1666 , \1696 );
nor \U$1321 ( \1698 , \1661 , \1697 );
and \U$1322 ( \1699 , \1680 , \1688 );
not \U$1323 ( \1700 , \1680 );
not \U$1324 ( \1701 , \1688 );
and \U$1325 ( \1702 , \1700 , \1701 );
nor \U$1326 ( \1703 , \1702 , \1684 );
nor \U$1327 ( \1704 , \1699 , \1703 );
nand \U$1328 ( \1705 , RIae78e90_132, RIae78ff8_135);
and \U$1329 ( \1706 , \1705 , RIae78bc0_126);
xor \U$1330 ( \1707 , \1631 , \1706 );
and \U$1331 ( \1708 , \1675 , \1129 );
xor \U$1332 ( \1709 , \1197 , RIae78b48_125);
and \U$1333 ( \1710 , \1709 , \1122 );
nor \U$1334 ( \1711 , \1708 , \1710 );
xor \U$1335 ( \1712 , \1707 , \1711 );
and \U$1336 ( \1713 , \1670 , \1679 );
and \U$1337 ( \1714 , \1669 , \1599 );
nor \U$1338 ( \1715 , \1713 , \1714 );
xor \U$1339 ( \1716 , \1669 , \1715 );
xor \U$1340 ( \1717 , \1712 , \1716 );
nand \U$1341 ( \1718 , \1704 , \1717 );
and \U$1342 ( \1719 , \1625 , \1698 , \1718 );
not \U$1343 ( \1720 , \1719 );
not \U$1344 ( \1721 , \839 );
not \U$1345 ( \1722 , \614 );
nor \U$1346 ( \1723 , \517 , \612 );
buf \U$1347 ( \1724 , \641 );
or \U$1348 ( \1725 , \1723 , \1724 );
buf \U$1349 ( \1726 , \672 );
not \U$1350 ( \1727 , \1726 );
nand \U$1351 ( \1728 , \1725 , \1727 );
not \U$1352 ( \1729 , \1728 );
or \U$1353 ( \1730 , \1722 , \1729 );
buf \U$1354 ( \1731 , \678 );
nand \U$1355 ( \1732 , \1730 , \1731 );
not \U$1356 ( \1733 , \1732 );
nand \U$1357 ( \1734 , \616 , \680 );
not \U$1358 ( \1735 , \1734 );
and \U$1359 ( \1736 , \1733 , \1735 );
and \U$1360 ( \1737 , \1732 , \1734 );
nor \U$1361 ( \1738 , \1736 , \1737 );
buf \U$1362 ( \1739 , \1738 );
not \U$1363 ( \1740 , \1739 );
not \U$1364 ( \1741 , \1740 );
not \U$1365 ( \1742 , RIae78f80_134);
xor \U$1366 ( \1743 , \1741 , \1742 );
not \U$1367 ( \1744 , \1743 );
or \U$1368 ( \1745 , \1721 , \1744 );
buf \U$1369 ( \1746 , \1728 );
not \U$1370 ( \1747 , \1746 );
nand \U$1371 ( \1748 , \614 , \1731 );
not \U$1372 ( \1749 , \1748 );
and \U$1373 ( \1750 , \1747 , \1749 );
and \U$1374 ( \1751 , \1746 , \1748 );
nor \U$1375 ( \1752 , \1750 , \1751 );
not \U$1376 ( \1753 , \1752 );
not \U$1377 ( \1754 , \1753 );
not \U$1378 ( \1755 , \1754 );
and \U$1379 ( \1756 , RIae78f80_134, \1755 );
not \U$1380 ( \1757 , RIae78f80_134);
xor \U$1381 ( \1758 , \1746 , \1748 );
not \U$1382 ( \1759 , \1758 );
not \U$1383 ( \1760 , \1759 );
and \U$1384 ( \1761 , \1757 , \1760 );
nor \U$1385 ( \1762 , \1756 , \1761 );
nand \U$1386 ( \1763 , \1762 , \797 );
nand \U$1387 ( \1764 , \1745 , \1763 );
not \U$1388 ( \1765 , \1259 );
not \U$1389 ( \1766 , \636 );
not \U$1390 ( \1767 , \633 );
not \U$1391 ( \1768 , \516 );
or \U$1392 ( \1769 , \612 , \1768 );
not \U$1393 ( \1770 , \1769 );
or \U$1394 ( \1771 , \1767 , \1770 );
not \U$1395 ( \1772 , \652 );
not \U$1396 ( \1773 , \654 );
or \U$1397 ( \1774 , \1772 , \1773 );
not \U$1398 ( \1775 , \657 );
nand \U$1399 ( \1776 , \1774 , \1775 );
nand \U$1400 ( \1777 , \1771 , \1776 );
not \U$1401 ( \1778 , \1777 );
or \U$1402 ( \1779 , \1766 , \1778 );
not \U$1403 ( \1780 , \665 );
nand \U$1404 ( \1781 , \1779 , \1780 );
not \U$1405 ( \1782 , \1781 );
nand \U$1406 ( \1783 , \637 , \668 );
not \U$1407 ( \1784 , \1783 );
and \U$1408 ( \1785 , \1782 , \1784 );
and \U$1409 ( \1786 , \1781 , \1783 );
nor \U$1410 ( \1787 , \1785 , \1786 );
buf \U$1411 ( \1788 , \1787 );
buf \U$1412 ( \1789 , \1788 );
buf \U$1413 ( \1790 , \1789 );
and \U$1414 ( \1791 , \1790 , \921 );
not \U$1415 ( \1792 , \1790 );
and \U$1416 ( \1793 , \1792 , RIae78e90_132);
nor \U$1417 ( \1794 , \1791 , \1793 );
not \U$1418 ( \1795 , \1794 );
or \U$1419 ( \1796 , \1765 , \1795 );
not \U$1420 ( \1797 , \638 );
not \U$1421 ( \1798 , \1777 );
or \U$1422 ( \1799 , \1797 , \1798 );
not \U$1423 ( \1800 , \669 );
nand \U$1424 ( \1801 , \1799 , \1800 );
nand \U$1425 ( \1802 , \640 , \671 );
not \U$1426 ( \1803 , \1802 );
and \U$1427 ( \1804 , \1801 , \1803 );
not \U$1428 ( \1805 , \1801 );
and \U$1429 ( \1806 , \1805 , \1802 );
nor \U$1430 ( \1807 , \1804 , \1806 );
buf \U$1431 ( \1808 , \1807 );
not \U$1432 ( \1809 , \1808 );
xnor \U$1433 ( \1810 , \1809 , RIae78e90_132);
nand \U$1434 ( \1811 , \1810 , \1321 );
nand \U$1435 ( \1812 , \1796 , \1811 );
xor \U$1436 ( \1813 , \1764 , \1812 );
and \U$1437 ( \1814 , RIae79ac0_158, RIae79b38_159);
not \U$1438 ( \1815 , RIae79ac0_158);
not \U$1439 ( \1816 , RIae79b38_159);
and \U$1440 ( \1817 , \1815 , \1816 );
nor \U$1441 ( \1818 , \1814 , \1817 );
not \U$1442 ( \1819 , \1818 );
not \U$1443 ( \1820 , \1819 );
buf \U$1444 ( \1821 , \1820 );
buf \U$1445 ( \1822 , \1821 );
not \U$1446 ( \1823 , \1822 );
and \U$1447 ( \1824 , RIae79688_149, \1186 );
not \U$1448 ( \1825 , RIae79688_149);
not \U$1449 ( \1826 , \1186 );
and \U$1450 ( \1827 , \1825 , \1826 );
or \U$1451 ( \1828 , \1824 , \1827 );
not \U$1452 ( \1829 , \1828 );
or \U$1453 ( \1830 , \1823 , \1829 );
and \U$1454 ( \1831 , RIae79688_149, \1405 );
not \U$1455 ( \1832 , RIae79688_149);
not \U$1456 ( \1833 , \1404 );
buf \U$1457 ( \1834 , \1833 );
not \U$1458 ( \1835 , \1834 );
and \U$1459 ( \1836 , \1832 , \1835 );
or \U$1460 ( \1837 , \1831 , \1836 );
and \U$1461 ( \1838 , RIae79688_149, RIae79b38_159);
not \U$1462 ( \1839 , RIae79688_149);
and \U$1463 ( \1840 , \1839 , \1816 );
nor \U$1464 ( \1841 , \1838 , \1840 );
and \U$1465 ( \1842 , \1819 , \1841 );
buf \U$1466 ( \1843 , \1842 );
buf \U$1467 ( \1844 , \1843 );
nand \U$1468 ( \1845 , \1837 , \1844 );
nand \U$1469 ( \1846 , \1830 , \1845 );
and \U$1470 ( \1847 , \1813 , \1846 );
and \U$1471 ( \1848 , \1764 , \1812 );
or \U$1472 ( \1849 , \1847 , \1848 );
not \U$1473 ( \1850 , RIae78b48_125);
not \U$1474 ( \1851 , \1723 );
not \U$1475 ( \1852 , \1851 );
nor \U$1476 ( \1853 , RIae75b78_23, RIae75bf0_24);
or \U$1477 ( \1854 , \1852 , \1853 );
nand \U$1478 ( \1855 , \1854 , \645 );
not \U$1479 ( \1856 , \644 );
nand \U$1480 ( \1857 , \1856 , \647 );
xor \U$1481 ( \1858 , \1855 , \1857 );
buf \U$1482 ( \1859 , \1858 );
buf \U$1483 ( \1860 , \1859 );
nor \U$1484 ( \1861 , \1850 , \1860 );
xnor \U$1485 ( \1862 , RIae799d0_156, RIae79610_148);
not \U$1486 ( \1863 , \1862 );
buf \U$1487 ( \1864 , \1863 );
not \U$1488 ( \1865 , \1864 );
not \U$1489 ( \1866 , \388 );
not \U$1490 ( \1867 , \1866 );
not \U$1491 ( \1868 , \1171 );
or \U$1492 ( \1869 , \1867 , \1868 );
nand \U$1493 ( \1870 , \1869 , \717 );
not \U$1494 ( \1871 , \389 );
nand \U$1495 ( \1872 , \1871 , \719 );
and \U$1496 ( \1873 , \1870 , \1872 );
not \U$1497 ( \1874 , \1870 );
not \U$1498 ( \1875 , \1872 );
and \U$1499 ( \1876 , \1874 , \1875 );
nor \U$1500 ( \1877 , \1873 , \1876 );
buf \U$1501 ( \1878 , \1877 );
not \U$1502 ( \1879 , \1878 );
not \U$1503 ( \1880 , \1879 );
xnor \U$1504 ( \1881 , \1880 , RIae793b8_143);
not \U$1505 ( \1882 , \1881 );
or \U$1506 ( \1883 , \1865 , \1882 );
not \U$1507 ( \1884 , RIae793b8_143);
not \U$1508 ( \1885 , \1884 );
and \U$1509 ( \1886 , \1866 , \717 );
not \U$1510 ( \1887 , \1886 );
not \U$1511 ( \1888 , \1171 );
not \U$1512 ( \1889 , \1888 );
or \U$1513 ( \1890 , \1887 , \1889 );
not \U$1514 ( \1891 , \1866 );
not \U$1515 ( \1892 , \717 );
or \U$1516 ( \1893 , \1891 , \1892 );
not \U$1517 ( \1894 , \1888 );
nand \U$1518 ( \1895 , \1893 , \1894 );
nand \U$1519 ( \1896 , \1890 , \1895 );
buf \U$1520 ( \1897 , \1896 );
buf \U$1521 ( \1898 , \1897 );
buf \U$1522 ( \1899 , \1898 );
not \U$1523 ( \1900 , \1899 );
or \U$1524 ( \1901 , \1885 , \1900 );
not \U$1525 ( \1902 , RIae793b8_143);
or \U$1526 ( \1903 , \1899 , \1902 );
nand \U$1527 ( \1904 , \1901 , \1903 );
not \U$1528 ( \1905 , RIae799d0_156);
and \U$1529 ( \1906 , \1902 , \1905 );
and \U$1530 ( \1907 , RIae793b8_143, RIae799d0_156);
nor \U$1531 ( \1908 , \1906 , \1907 );
and \U$1532 ( \1909 , \1862 , \1908 );
buf \U$1533 ( \1910 , \1909 );
nand \U$1534 ( \1911 , \1904 , \1910 );
nand \U$1535 ( \1912 , \1883 , \1911 );
xor \U$1536 ( \1913 , \1861 , \1912 );
nand \U$1537 ( \1914 , RIae798e0_154, RIae79958_155);
not \U$1538 ( \1915 , \1914 );
nor \U$1539 ( \1916 , RIae798e0_154, RIae79958_155);
nor \U$1540 ( \1917 , \1915 , \1916 );
buf \U$1541 ( \1918 , \1917 );
buf \U$1542 ( \1919 , \1918 );
not \U$1543 ( \1920 , \1919 );
not \U$1544 ( \1921 , \919 );
xor \U$1545 ( \1922 , RIae794a8_145, \1921 );
not \U$1546 ( \1923 , \1922 );
or \U$1547 ( \1924 , \1920 , \1923 );
xnor \U$1548 ( \1925 , \938 , RIae794a8_145);
not \U$1549 ( \1926 , RIae79958_155);
and \U$1550 ( \1927 , RIae794a8_145, \1926 );
not \U$1551 ( \1928 , RIae794a8_145);
and \U$1552 ( \1929 , \1928 , RIae79958_155);
nor \U$1553 ( \1930 , \1927 , \1929 );
nor \U$1554 ( \1931 , \1917 , \1930 );
buf \U$1555 ( \1932 , \1931 );
buf \U$1556 ( \1933 , \1932 );
nand \U$1557 ( \1934 , \1925 , \1933 );
nand \U$1558 ( \1935 , \1924 , \1934 );
and \U$1559 ( \1936 , \1913 , \1935 );
and \U$1560 ( \1937 , \1861 , \1912 );
or \U$1561 ( \1938 , \1936 , \1937 );
xor \U$1562 ( \1939 , \1849 , \1938 );
not \U$1563 ( \1940 , \651 );
or \U$1564 ( \1941 , \1723 , \632 );
not \U$1565 ( \1942 , \648 );
nand \U$1566 ( \1943 , \1941 , \1942 );
not \U$1567 ( \1944 , \1943 );
or \U$1568 ( \1945 , \1940 , \1944 );
not \U$1569 ( \1946 , \649 );
nand \U$1570 ( \1947 , \1945 , \1946 );
nand \U$1571 ( \1948 , \1775 , \654 );
not \U$1572 ( \1949 , \1948 );
and \U$1573 ( \1950 , \1947 , \1949 );
not \U$1574 ( \1951 , \1947 );
and \U$1575 ( \1952 , \1951 , \1948 );
nor \U$1576 ( \1953 , \1950 , \1952 );
not \U$1577 ( \1954 , \1953 );
buf \U$1578 ( \1955 , \1954 );
not \U$1579 ( \1956 , \1955 );
xor \U$1580 ( \1957 , RIae78b48_125, \1956 );
not \U$1581 ( \1958 , \1957 );
not \U$1582 ( \1959 , \868 );
or \U$1583 ( \1960 , \1958 , \1959 );
buf \U$1584 ( \1961 , \1943 );
not \U$1585 ( \1962 , \1961 );
not \U$1586 ( \1963 , \649 );
nand \U$1587 ( \1964 , \1963 , \651 );
not \U$1588 ( \1965 , \1964 );
and \U$1589 ( \1966 , \1962 , \1965 );
and \U$1590 ( \1967 , \1961 , \1964 );
nor \U$1591 ( \1968 , \1966 , \1967 );
buf \U$1592 ( \1969 , \1968 );
buf \U$1593 ( \1970 , \1969 );
and \U$1594 ( \1971 , RIae78b48_125, \1970 );
not \U$1595 ( \1972 , RIae78b48_125);
not \U$1596 ( \1973 , \1970 );
and \U$1597 ( \1974 , \1972 , \1973 );
nor \U$1598 ( \1975 , \1971 , \1974 );
not \U$1599 ( \1976 , \893 );
or \U$1600 ( \1977 , \1975 , \1976 );
nand \U$1601 ( \1978 , \1960 , \1977 );
not \U$1602 ( \1979 , \1978 );
or \U$1603 ( \1980 , RIae79700_150, RIae797f0_152);
not \U$1604 ( \1981 , RIae79700_150);
not \U$1605 ( \1982 , RIae797f0_152);
or \U$1606 ( \1983 , \1981 , \1982 );
xor \U$1607 ( \1984 , RIae79700_150, RIae79778_151);
not \U$1608 ( \1985 , \1984 );
nand \U$1609 ( \1986 , \1980 , \1983 , \1985 );
not \U$1610 ( \1987 , \1986 );
buf \U$1611 ( \1988 , \1987 );
buf \U$1612 ( \1989 , \1988 );
not \U$1613 ( \1990 , \1989 );
not \U$1614 ( \1991 , RIae797f0_152);
not \U$1615 ( \1992 , \1991 );
buf \U$1616 ( \1993 , \779 );
not \U$1617 ( \1994 , \1993 );
not \U$1618 ( \1995 , \1994 );
or \U$1619 ( \1996 , \1992 , \1995 );
not \U$1620 ( \1997 , RIae797f0_152);
or \U$1621 ( \1998 , \1994 , \1997 );
nand \U$1622 ( \1999 , \1996 , \1998 );
not \U$1623 ( \2000 , \1999 );
or \U$1624 ( \2001 , \1990 , \2000 );
and \U$1625 ( \2002 , RIae797f0_152, \835 );
not \U$1626 ( \2003 , RIae797f0_152);
not \U$1627 ( \2004 , \827 );
and \U$1628 ( \2005 , \2003 , \2004 );
or \U$1629 ( \2006 , \2002 , \2005 );
buf \U$1630 ( \2007 , \1984 );
nand \U$1631 ( \2008 , \2006 , \2007 );
nand \U$1632 ( \2009 , \2001 , \2008 );
xor \U$1633 ( \2010 , RIae79598_147, RIae79688_149);
buf \U$1634 ( \2011 , \2010 );
not \U$1635 ( \2012 , \2011 );
and \U$1636 ( \2013 , \390 , \391 );
not \U$1637 ( \2014 , \2013 );
not \U$1638 ( \2015 , \1171 );
or \U$1639 ( \2016 , \2014 , \2015 );
not \U$1640 ( \2017 , \724 );
nand \U$1641 ( \2018 , \2016 , \2017 );
nand \U$1642 ( \2019 , \392 , \727 );
not \U$1643 ( \2020 , \2019 );
and \U$1644 ( \2021 , \2018 , \2020 );
not \U$1645 ( \2022 , \2018 );
and \U$1646 ( \2023 , \2022 , \2019 );
nor \U$1647 ( \2024 , \2021 , \2023 );
buf \U$1648 ( \2025 , \2024 );
not \U$1649 ( \2026 , \2025 );
buf \U$1650 ( \2027 , \2026 );
and \U$1651 ( \2028 , RIae79610_148, \2027 );
not \U$1652 ( \2029 , RIae79610_148);
not \U$1653 ( \2030 , \2025 );
not \U$1654 ( \2031 , \2030 );
and \U$1655 ( \2032 , \2029 , \2031 );
or \U$1656 ( \2033 , \2028 , \2032 );
not \U$1657 ( \2034 , \2033 );
or \U$1658 ( \2035 , \2012 , \2034 );
not \U$1659 ( \2036 , \390 );
not \U$1660 ( \2037 , \1171 );
or \U$1661 ( \2038 , \2036 , \2037 );
not \U$1662 ( \2039 , \720 );
nand \U$1663 ( \2040 , \2038 , \2039 );
nand \U$1664 ( \2041 , \391 , \723 );
and \U$1665 ( \2042 , \2040 , \2041 );
not \U$1666 ( \2043 , \2040 );
not \U$1667 ( \2044 , \2041 );
and \U$1668 ( \2045 , \2043 , \2044 );
nor \U$1669 ( \2046 , \2042 , \2045 );
buf \U$1670 ( \2047 , \2046 );
not \U$1671 ( \2048 , \2047 );
not \U$1672 ( \2049 , \2048 );
not \U$1673 ( \2050 , \2049 );
and \U$1674 ( \2051 , \2050 , RIae79610_148);
not \U$1675 ( \2052 , \2050 );
not \U$1676 ( \2053 , RIae79610_148);
and \U$1677 ( \2054 , \2052 , \2053 );
nor \U$1678 ( \2055 , \2051 , \2054 );
not \U$1679 ( \2056 , RIae79610_148);
not \U$1680 ( \2057 , RIae79598_147);
and \U$1681 ( \2058 , \2056 , \2057 );
and \U$1682 ( \2059 , RIae79598_147, RIae79610_148);
nor \U$1683 ( \2060 , \2058 , \2059 );
not \U$1684 ( \2061 , \2060 );
nor \U$1685 ( \2062 , \2061 , \2010 );
buf \U$1686 ( \2063 , \2062 );
nand \U$1687 ( \2064 , \2055 , \2063 );
nand \U$1688 ( \2065 , \2035 , \2064 );
xor \U$1689 ( \2066 , \2009 , \2065 );
not \U$1690 ( \2067 , \2066 );
or \U$1691 ( \2068 , \1979 , \2067 );
buf \U$1692 ( \2069 , \2009 );
nand \U$1693 ( \2070 , \2069 , \2065 );
nand \U$1694 ( \2071 , \2068 , \2070 );
xor \U$1695 ( \2072 , \1939 , \2071 );
nor \U$1696 ( \2073 , \1970 , \860 );
not \U$1697 ( \2074 , \893 );
not \U$1698 ( \2075 , \1957 );
or \U$1699 ( \2076 , \2074 , \2075 );
or \U$1700 ( \2077 , RIae75f38_31, RIae75fb0_32);
buf \U$1701 ( \2078 , \662 );
nand \U$1702 ( \2079 , \2077 , \2078 );
not \U$1703 ( \2080 , \2079 );
not \U$1704 ( \2081 , \1777 );
or \U$1705 ( \2082 , \2080 , \2081 );
not \U$1706 ( \2083 , \1777 );
not \U$1707 ( \2084 , \635 );
and \U$1708 ( \2085 , \2084 , \2078 );
nand \U$1709 ( \2086 , \2083 , \2085 );
nand \U$1710 ( \2087 , \2082 , \2086 );
buf \U$1711 ( \2088 , \2087 );
buf \U$1712 ( \2089 , \2088 );
not \U$1713 ( \2090 , \2089 );
and \U$1714 ( \2091 , RIae78b48_125, \2090 );
not \U$1715 ( \2092 , RIae78b48_125);
buf \U$1716 ( \2093 , \2087 );
and \U$1717 ( \2094 , \2092 , \2093 );
or \U$1718 ( \2095 , \2091 , \2094 );
buf \U$1719 ( \2096 , \867 );
nand \U$1720 ( \2097 , \2095 , \2096 );
nand \U$1721 ( \2098 , \2076 , \2097 );
xor \U$1722 ( \2099 , \2073 , \2098 );
not \U$1723 ( \2100 , \2011 );
not \U$1724 ( \2101 , \1404 );
not \U$1725 ( \2102 , \2101 );
and \U$1726 ( \2103 , RIae79610_148, \2102 );
not \U$1727 ( \2104 , RIae79610_148);
and \U$1728 ( \2105 , \2104 , \1834 );
nor \U$1729 ( \2106 , \2103 , \2105 );
not \U$1730 ( \2107 , \2106 );
or \U$1731 ( \2108 , \2100 , \2107 );
nand \U$1732 ( \2109 , \2033 , \2063 );
nand \U$1733 ( \2110 , \2108 , \2109 );
xor \U$1734 ( \2111 , \2099 , \2110 );
not \U$1735 ( \2112 , \1013 );
buf \U$1736 ( \2113 , \621 );
not \U$1737 ( \2114 , \2113 );
not \U$1738 ( \2115 , \619 );
not \U$1739 ( \2116 , \1724 );
not \U$1740 ( \2117 , \2116 );
not \U$1741 ( \2118 , \1769 );
or \U$1742 ( \2119 , \2117 , \2118 );
nand \U$1743 ( \2120 , \2119 , \1727 );
not \U$1744 ( \2121 , \2120 );
or \U$1745 ( \2122 , \2115 , \2121 );
not \U$1746 ( \2123 , \689 );
nand \U$1747 ( \2124 , \2122 , \2123 );
not \U$1748 ( \2125 , \2124 );
or \U$1749 ( \2126 , \2114 , \2125 );
buf \U$1750 ( \2127 , \694 );
nand \U$1751 ( \2128 , \2126 , \2127 );
not \U$1752 ( \2129 , \2128 );
nand \U$1753 ( \2130 , \623 , \696 );
not \U$1754 ( \2131 , \2130 );
and \U$1755 ( \2132 , \2129 , \2131 );
and \U$1756 ( \2133 , \2128 , \2130 );
nor \U$1757 ( \2134 , \2132 , \2133 );
not \U$1758 ( \2135 , \2134 );
not \U$1759 ( \2136 , \2135 );
buf \U$1760 ( \2137 , \2136 );
and \U$1761 ( \2138 , RIae79160_138, \2137 );
not \U$1762 ( \2139 , RIae79160_138);
not \U$1763 ( \2140 , \2135 );
buf \U$1764 ( \2141 , \2140 );
not \U$1765 ( \2142 , \2141 );
and \U$1766 ( \2143 , \2139 , \2142 );
or \U$1767 ( \2144 , \2138 , \2143 );
not \U$1768 ( \2145 , \2144 );
or \U$1769 ( \2146 , \2112 , \2145 );
not \U$1770 ( \2147 , \2124 );
nand \U$1771 ( \2148 , \621 , \2127 );
not \U$1772 ( \2149 , \2148 );
and \U$1773 ( \2150 , \2147 , \2149 );
and \U$1774 ( \2151 , \2124 , \2148 );
nor \U$1775 ( \2152 , \2150 , \2151 );
buf \U$1776 ( \2153 , \2152 );
not \U$1777 ( \2154 , \2153 );
not \U$1778 ( \2155 , \2154 );
xnor \U$1779 ( \2156 , RIae79160_138, \2155 );
buf \U$1780 ( \2157 , \1008 );
nand \U$1781 ( \2158 , \2156 , \2157 );
nand \U$1782 ( \2159 , \2146 , \2158 );
not \U$1783 ( \2160 , \2159 );
xor \U$1784 ( \2161 , RIae79430_144, RIae794a8_145);
buf \U$1785 ( \2162 , \2161 );
buf \U$1786 ( \2163 , \2162 );
not \U$1787 ( \2164 , \2163 );
not \U$1788 ( \2165 , RIae79520_146);
not \U$1789 ( \2166 , \854 );
not \U$1790 ( \2167 , \2166 );
or \U$1791 ( \2168 , \2165 , \2167 );
not \U$1792 ( \2169 , \854 );
or \U$1793 ( \2170 , \2169 , RIae79520_146);
nand \U$1794 ( \2171 , \2168 , \2170 );
not \U$1795 ( \2172 , \2171 );
or \U$1796 ( \2173 , \2164 , \2172 );
not \U$1797 ( \2174 , RIae79520_146);
buf \U$1798 ( \2175 , \877 );
not \U$1799 ( \2176 , \2175 );
or \U$1800 ( \2177 , \2174 , \2176 );
not \U$1801 ( \2178 , \877 );
not \U$1802 ( \2179 , \2178 );
or \U$1803 ( \2180 , \2179 , RIae79520_146);
nand \U$1804 ( \2181 , \2177 , \2180 );
not \U$1805 ( \2182 , \2161 );
not \U$1806 ( \2183 , RIae79520_146);
not \U$1807 ( \2184 , RIae79430_144);
and \U$1808 ( \2185 , \2183 , \2184 );
and \U$1809 ( \2186 , RIae79430_144, RIae79520_146);
nor \U$1810 ( \2187 , \2185 , \2186 );
and \U$1811 ( \2188 , \2182 , \2187 );
buf \U$1812 ( \2189 , \2188 );
nand \U$1813 ( \2190 , \2181 , \2189 );
nand \U$1814 ( \2191 , \2173 , \2190 );
not \U$1815 ( \2192 , \1501 );
not \U$1816 ( \2193 , RIae79250_140);
and \U$1817 ( \2194 , \623 , \621 );
and \U$1818 ( \2195 , \2194 , \620 );
not \U$1819 ( \2196 , \2195 );
not \U$1820 ( \2197 , \2124 );
or \U$1821 ( \2198 , \2196 , \2197 );
not \U$1822 ( \2199 , \701 );
nand \U$1823 ( \2200 , \2198 , \2199 );
nand \U$1824 ( \2201 , \624 , \704 );
not \U$1825 ( \2202 , \2201 );
and \U$1826 ( \2203 , \2200 , \2202 );
not \U$1827 ( \2204 , \2200 );
and \U$1828 ( \2205 , \2204 , \2201 );
nor \U$1829 ( \2206 , \2203 , \2205 );
buf \U$1830 ( \2207 , \2206 );
not \U$1831 ( \2208 , \2207 );
not \U$1832 ( \2209 , \2208 );
or \U$1833 ( \2210 , \2193 , \2209 );
buf \U$1834 ( \2211 , \2207 );
not \U$1835 ( \2212 , \2211 );
or \U$1836 ( \2213 , \2212 , RIae79250_140);
nand \U$1837 ( \2214 , \2210 , \2213 );
not \U$1838 ( \2215 , \2214 );
or \U$1839 ( \2216 , \2192 , \2215 );
not \U$1840 ( \2217 , RIae79250_140);
not \U$1841 ( \2218 , \2217 );
not \U$1842 ( \2219 , \2194 );
not \U$1843 ( \2220 , \2124 );
or \U$1844 ( \2221 , \2219 , \2220 );
not \U$1845 ( \2222 , \697 );
nand \U$1846 ( \2223 , \2221 , \2222 );
not \U$1847 ( \2224 , \2223 );
nand \U$1848 ( \2225 , \620 , \700 );
not \U$1849 ( \2226 , \2225 );
and \U$1850 ( \2227 , \2224 , \2226 );
and \U$1851 ( \2228 , \2223 , \2225 );
nor \U$1852 ( \2229 , \2227 , \2228 );
buf \U$1853 ( \2230 , \2229 );
not \U$1854 ( \2231 , \2230 );
not \U$1855 ( \2232 , \2231 );
or \U$1856 ( \2233 , \2218 , \2232 );
nand \U$1857 ( \2234 , \2230 , RIae79250_140);
nand \U$1858 ( \2235 , \2233 , \2234 );
nand \U$1859 ( \2236 , \2235 , \1499 );
nand \U$1860 ( \2237 , \2216 , \2236 );
xor \U$1861 ( \2238 , \2191 , \2237 );
not \U$1862 ( \2239 , \2238 );
or \U$1863 ( \2240 , \2160 , \2239 );
nand \U$1864 ( \2241 , \2237 , \2191 );
nand \U$1865 ( \2242 , \2240 , \2241 );
xor \U$1866 ( \2243 , \2111 , \2242 );
and \U$1867 ( \2244 , RIae79520_146, RIae79a48_157);
not \U$1868 ( \2245 , RIae79520_146);
not \U$1869 ( \2246 , RIae79a48_157);
and \U$1870 ( \2247 , \2245 , \2246 );
nor \U$1871 ( \2248 , \2244 , \2247 );
buf \U$1872 ( \2249 , \2248 );
not \U$1873 ( \2250 , \2249 );
not \U$1874 ( \2251 , \2250 );
buf \U$1875 ( \2252 , \2251 );
not \U$1876 ( \2253 , \2252 );
not \U$1877 ( \2254 , RIae79ac0_158);
not \U$1878 ( \2255 , \1119 );
or \U$1879 ( \2256 , \2254 , \2255 );
or \U$1880 ( \2257 , \1119 , RIae79ac0_158);
nand \U$1881 ( \2258 , \2256 , \2257 );
not \U$1882 ( \2259 , \2258 );
or \U$1883 ( \2260 , \2253 , \2259 );
not \U$1884 ( \2261 , RIae79ac0_158);
not \U$1885 ( \2262 , \975 );
not \U$1886 ( \2263 , \2262 );
not \U$1887 ( \2264 , \2263 );
or \U$1888 ( \2265 , \2261 , \2264 );
or \U$1889 ( \2266 , \2263 , RIae79ac0_158);
nand \U$1890 ( \2267 , \2265 , \2266 );
not \U$1891 ( \2268 , RIae79ac0_158);
and \U$1892 ( \2269 , \2268 , \2246 );
and \U$1893 ( \2270 , RIae79a48_157, RIae79ac0_158);
nor \U$1894 ( \2271 , \2269 , \2270 , \2248 );
buf \U$1895 ( \2272 , \2271 );
nand \U$1896 ( \2273 , \2267 , \2272 );
nand \U$1897 ( \2274 , \2260 , \2273 );
not \U$1898 ( \2275 , \2274 );
buf \U$1899 ( \2276 , \1062 );
not \U$1900 ( \2277 , \614 );
nor \U$1901 ( \2278 , \2277 , \615 );
not \U$1902 ( \2279 , \2278 );
not \U$1903 ( \2280 , \2120 );
or \U$1904 ( \2281 , \2279 , \2280 );
not \U$1905 ( \2282 , \681 );
nand \U$1906 ( \2283 , \2281 , \2282 );
nand \U$1907 ( \2284 , \617 , \684 );
xor \U$1908 ( \2285 , \2283 , \2284 );
buf \U$1909 ( \2286 , \2285 );
buf \U$1910 ( \2287 , \2286 );
and \U$1911 ( \2288 , \2287 , \1039 );
not \U$1912 ( \2289 , \2287 );
and \U$1913 ( \2290 , \2289 , RIae79070_136);
nor \U$1914 ( \2291 , \2288 , \2290 );
and \U$1915 ( \2292 , \2276 , \2291 );
and \U$1916 ( \2293 , \2278 , \617 );
not \U$1917 ( \2294 , \2293 );
not \U$1918 ( \2295 , \1728 );
or \U$1919 ( \2296 , \2294 , \2295 );
not \U$1920 ( \2297 , \685 );
nand \U$1921 ( \2298 , \2296 , \2297 );
not \U$1922 ( \2299 , \2298 );
nand \U$1923 ( \2300 , \618 , \688 );
not \U$1924 ( \2301 , \2300 );
and \U$1925 ( \2302 , \2299 , \2301 );
and \U$1926 ( \2303 , \2298 , \2300 );
nor \U$1927 ( \2304 , \2302 , \2303 );
buf \U$1928 ( \2305 , \2304 );
and \U$1929 ( \2306 , RIae79070_136, \2305 );
not \U$1930 ( \2307 , RIae79070_136);
xnor \U$1931 ( \2308 , \2298 , \2300 );
buf \U$1932 ( \2309 , \2308 );
buf \U$1933 ( \2310 , \2309 );
and \U$1934 ( \2311 , \2307 , \2310 );
or \U$1935 ( \2312 , \2306 , \2311 );
and \U$1936 ( \2313 , \2312 , \1049 );
nor \U$1937 ( \2314 , \2292 , \2313 );
not \U$1938 ( \2315 , \2314 );
and \U$1939 ( \2316 , \2275 , \2315 );
and \U$1940 ( \2317 , \2274 , \2314 );
nor \U$1941 ( \2318 , \2316 , \2317 );
and \U$1942 ( \2319 , RIae797f0_152, RIae79868_153);
nor \U$1943 ( \2320 , RIae797f0_152, RIae79868_153);
nor \U$1944 ( \2321 , \2319 , \2320 );
buf \U$1945 ( \2322 , \2321 );
buf \U$1946 ( \2323 , \1140 );
not \U$1947 ( \2324 , \2323 );
xnor \U$1948 ( \2325 , RIae798e0_154, \2324 );
and \U$1949 ( \2326 , \2322 , \2325 );
not \U$1950 ( \2327 , RIae798e0_154);
not \U$1951 ( \2328 , \1158 );
or \U$1952 ( \2329 , \2327 , \2328 );
buf \U$1953 ( \2330 , \1157 );
not \U$1954 ( \2331 , \2330 );
or \U$1955 ( \2332 , \2331 , RIae798e0_154);
nand \U$1956 ( \2333 , \2329 , \2332 );
not \U$1957 ( \2334 , RIae798e0_154);
not \U$1958 ( \2335 , RIae79868_153);
and \U$1959 ( \2336 , \2334 , \2335 );
and \U$1960 ( \2337 , RIae79868_153, RIae798e0_154);
nor \U$1961 ( \2338 , \2336 , \2337 , \2321 );
buf \U$1962 ( \2339 , \2338 );
buf \U$1963 ( \2340 , \2339 );
buf \U$1964 ( \2341 , \2340 );
and \U$1965 ( \2342 , \2333 , \2341 );
nor \U$1966 ( \2343 , \2326 , \2342 );
or \U$1967 ( \2344 , \2318 , \2343 );
not \U$1968 ( \2345 , \2314 );
nand \U$1969 ( \2346 , \2345 , \2274 );
nand \U$1970 ( \2347 , \2344 , \2346 );
xor \U$1971 ( \2348 , \2243 , \2347 );
xor \U$1972 ( \2349 , \2072 , \2348 );
not \U$1973 ( \2350 , \952 );
not \U$1974 ( \2351 , \1947 );
not \U$1975 ( \2352 , \1948 );
and \U$1976 ( \2353 , \2351 , \2352 );
and \U$1977 ( \2354 , \1947 , \1948 );
nor \U$1978 ( \2355 , \2353 , \2354 );
not \U$1979 ( \2356 , \2355 );
not \U$1980 ( \2357 , \2356 );
buf \U$1981 ( \2358 , \2357 );
and \U$1982 ( \2359 , \2358 , \1286 );
not \U$1983 ( \2360 , \2358 );
and \U$1984 ( \2361 , \2360 , RIae78bc0_126);
nor \U$1985 ( \2362 , \2359 , \2361 );
not \U$1986 ( \2363 , \2362 );
or \U$1987 ( \2364 , \2350 , \2363 );
and \U$1988 ( \2365 , RIae78bc0_126, \2093 );
not \U$1989 ( \2366 , RIae78bc0_126);
and \U$1990 ( \2367 , \2366 , \2090 );
nor \U$1991 ( \2368 , \2365 , \2367 );
nand \U$1992 ( \2369 , \1027 , \2368 );
nand \U$1993 ( \2370 , \2364 , \2369 );
not \U$1994 ( \2371 , \1822 );
not \U$1995 ( \2372 , \1837 );
or \U$1996 ( \2373 , \2371 , \2372 );
not \U$1997 ( \2374 , \2031 );
and \U$1998 ( \2375 , RIae79688_149, \2374 );
not \U$1999 ( \2376 , RIae79688_149);
and \U$2000 ( \2377 , \2376 , \2031 );
or \U$2001 ( \2378 , \2375 , \2377 );
nand \U$2002 ( \2379 , \2378 , \1844 );
nand \U$2003 ( \2380 , \2373 , \2379 );
xor \U$2004 ( \2381 , \2370 , \2380 );
or \U$2005 ( \2382 , \1975 , \1959 );
and \U$2006 ( \2383 , RIae78b48_125, \1860 );
not \U$2007 ( \2384 , RIae78b48_125);
not \U$2008 ( \2385 , \1859 );
and \U$2009 ( \2386 , \2384 , \2385 );
nor \U$2010 ( \2387 , \2383 , \2386 );
or \U$2011 ( \2388 , \2387 , \1128 );
nand \U$2012 ( \2389 , \2382 , \2388 );
and \U$2013 ( \2390 , \2381 , \2389 );
and \U$2014 ( \2391 , \2370 , \2380 );
nor \U$2015 ( \2392 , \2390 , \2391 );
not \U$2016 ( \2393 , \2392 );
not \U$2017 ( \2394 , \2393 );
not \U$2018 ( \2395 , \1852 );
not \U$2019 ( \2396 , \645 );
nor \U$2020 ( \2397 , \2396 , \1853 );
not \U$2021 ( \2398 , \2397 );
and \U$2022 ( \2399 , \2395 , \2398 );
and \U$2023 ( \2400 , \1852 , \2397 );
nor \U$2024 ( \2401 , \2399 , \2400 );
buf \U$2025 ( \2402 , \2401 );
buf \U$2026 ( \2403 , \2402 );
not \U$2027 ( \2404 , \2403 );
and \U$2028 ( \2405 , \2404 , RIae78b48_125);
not \U$2029 ( \2406 , RIae79ca0_162);
not \U$2030 ( \2407 , RIae79d18_163);
nand \U$2031 ( \2408 , \2406 , \2407 );
nand \U$2032 ( \2409 , RIae79ca0_162, RIae79d18_163);
nand \U$2033 ( \2410 , \2408 , \2409 );
not \U$2034 ( \2411 , \2410 );
and \U$2035 ( \2412 , RIae79c28_161, \2407 );
not \U$2036 ( \2413 , RIae79c28_161);
and \U$2037 ( \2414 , \2413 , RIae79d18_163);
nor \U$2038 ( \2415 , \2412 , \2414 );
nor \U$2039 ( \2416 , \2411 , \2415 );
buf \U$2040 ( \2417 , \2416 );
not \U$2041 ( \2418 , \2410 );
or \U$2042 ( \2419 , \2417 , \2418 );
nand \U$2043 ( \2420 , \2419 , RIae79c28_161);
xnor \U$2044 ( \2421 , \2405 , \2420 );
not \U$2045 ( \2422 , \2421 );
xor \U$2046 ( \2423 , RIae79bb0_160, RIae79c28_161);
not \U$2047 ( \2424 , \2423 );
and \U$2048 ( \2425 , RIae79778_151, RIae79bb0_160);
not \U$2049 ( \2426 , RIae79778_151);
not \U$2050 ( \2427 , RIae79bb0_160);
and \U$2051 ( \2428 , \2426 , \2427 );
nor \U$2052 ( \2429 , \2425 , \2428 );
nand \U$2053 ( \2430 , \2424 , \2429 );
not \U$2054 ( \2431 , \2430 );
buf \U$2055 ( \2432 , \2431 );
buf \U$2056 ( \2433 , \2432 );
not \U$2057 ( \2434 , \2433 );
not \U$2058 ( \2435 , RIae79778_151);
not \U$2059 ( \2436 , \828 );
or \U$2060 ( \2437 , \2435 , \2436 );
or \U$2061 ( \2438 , \835 , RIae79778_151);
nand \U$2062 ( \2439 , \2437 , \2438 );
not \U$2063 ( \2440 , \2439 );
or \U$2064 ( \2441 , \2434 , \2440 );
not \U$2065 ( \2442 , RIae79778_151);
not \U$2066 ( \2443 , \2442 );
not \U$2067 ( \2444 , \1194 );
not \U$2068 ( \2445 , \2444 );
or \U$2069 ( \2446 , \2443 , \2445 );
not \U$2070 ( \2447 , RIae79778_151);
or \U$2071 ( \2448 , \2444 , \2447 );
nand \U$2072 ( \2449 , \2446 , \2448 );
buf \U$2073 ( \2450 , \2423 );
nand \U$2074 ( \2451 , \2449 , \2450 );
nand \U$2075 ( \2452 , \2441 , \2451 );
and \U$2076 ( \2453 , \2422 , \2452 );
and \U$2077 ( \2454 , \2405 , \2420 );
nor \U$2078 ( \2455 , \2453 , \2454 );
not \U$2079 ( \2456 , \2455 );
buf \U$2080 ( \2457 , \1932 );
buf \U$2081 ( \2458 , \2457 );
not \U$2082 ( \2459 , \2458 );
not \U$2083 ( \2460 , RIae794a8_145);
not \U$2084 ( \2461 , \2169 );
or \U$2085 ( \2462 , \2460 , \2461 );
or \U$2086 ( \2463 , \855 , RIae794a8_145);
nand \U$2087 ( \2464 , \2462 , \2463 );
not \U$2088 ( \2465 , \2464 );
or \U$2089 ( \2466 , \2459 , \2465 );
buf \U$2090 ( \2467 , \1919 );
nand \U$2091 ( \2468 , \1925 , \2467 );
nand \U$2092 ( \2469 , \2466 , \2468 );
not \U$2093 ( \2470 , \2341 );
not \U$2094 ( \2471 , \1439 );
and \U$2095 ( \2472 , \2471 , RIae798e0_154);
not \U$2096 ( \2473 , \2471 );
and \U$2097 ( \2474 , \2473 , \2334 );
nor \U$2098 ( \2475 , \2472 , \2474 );
not \U$2099 ( \2476 , \2475 );
or \U$2100 ( \2477 , \2470 , \2476 );
nand \U$2101 ( \2478 , \2333 , \2322 );
nand \U$2102 ( \2479 , \2477 , \2478 );
xor \U$2103 ( \2480 , \2469 , \2479 );
and \U$2104 ( \2481 , \2011 , \2055 );
and \U$2105 ( \2482 , \1880 , \2056 );
not \U$2106 ( \2483 , \1880 );
and \U$2107 ( \2484 , \2483 , RIae79610_148);
nor \U$2108 ( \2485 , \2482 , \2484 );
and \U$2109 ( \2486 , \2485 , \2063 );
nor \U$2110 ( \2487 , \2481 , \2486 );
not \U$2111 ( \2488 , \2487 );
and \U$2112 ( \2489 , \2480 , \2488 );
and \U$2113 ( \2490 , \2469 , \2479 );
nor \U$2114 ( \2491 , \2489 , \2490 );
not \U$2115 ( \2492 , \2491 );
not \U$2116 ( \2493 , \2492 );
or \U$2117 ( \2494 , \2456 , \2493 );
or \U$2118 ( \2495 , \2492 , \2455 );
nand \U$2119 ( \2496 , \2494 , \2495 );
not \U$2120 ( \2497 , \2496 );
or \U$2121 ( \2498 , \2394 , \2497 );
not \U$2122 ( \2499 , \2455 );
nand \U$2123 ( \2500 , \2499 , \2492 );
nand \U$2124 ( \2501 , \2498 , \2500 );
xor \U$2125 ( \2502 , \2349 , \2501 );
and \U$2126 ( \2503 , RIae79bb0_160, RIae79c28_161);
not \U$2127 ( \2504 , RIae79778_151);
nor \U$2128 ( \2505 , \2503 , \2504 );
not \U$2129 ( \2506 , \2505 );
not \U$2130 ( \2507 , \1933 );
not \U$2131 ( \2508 , \1922 );
or \U$2132 ( \2509 , \2507 , \2508 );
not \U$2133 ( \2510 , \1289 );
and \U$2134 ( \2511 , RIae794a8_145, \2510 );
not \U$2135 ( \2512 , RIae794a8_145);
and \U$2136 ( \2513 , \2512 , \1159 );
or \U$2137 ( \2514 , \2511 , \2513 );
nand \U$2138 ( \2515 , \2514 , \1919 );
nand \U$2139 ( \2516 , \2509 , \2515 );
xor \U$2140 ( \2517 , \2506 , \2516 );
not \U$2141 ( \2518 , \2007 );
not \U$2142 ( \2519 , \2518 );
not \U$2143 ( \2520 , \2519 );
not \U$2144 ( \2521 , RIae797f0_152);
not \U$2145 ( \2522 , \2521 );
not \U$2146 ( \2523 , \992 );
or \U$2147 ( \2524 , \2522 , \2523 );
or \U$2148 ( \2525 , \992 , \2521 );
nand \U$2149 ( \2526 , \2524 , \2525 );
not \U$2150 ( \2527 , \2526 );
or \U$2151 ( \2528 , \2520 , \2527 );
buf \U$2152 ( \2529 , \1989 );
nand \U$2153 ( \2530 , \2006 , \2529 );
nand \U$2154 ( \2531 , \2528 , \2530 );
xnor \U$2155 ( \2532 , \2517 , \2531 );
not \U$2156 ( \2533 , \2532 );
not \U$2157 ( \2534 , \1259 );
not \U$2158 ( \2535 , \1810 );
or \U$2159 ( \2536 , \2534 , \2535 );
not \U$2160 ( \2537 , \1759 );
not \U$2161 ( \2538 , \1066 );
and \U$2162 ( \2539 , \2537 , \2538 );
and \U$2163 ( \2540 , \1755 , \921 );
nor \U$2164 ( \2541 , \2539 , \2540 );
not \U$2165 ( \2542 , \2541 );
nand \U$2166 ( \2543 , \2542 , \1074 );
nand \U$2167 ( \2544 , \2536 , \2543 );
buf \U$2168 ( \2545 , \2431 );
not \U$2169 ( \2546 , \2545 );
not \U$2170 ( \2547 , \2449 );
or \U$2171 ( \2548 , \2546 , \2547 );
nand \U$2172 ( \2549 , \2450 , RIae79778_151);
nand \U$2173 ( \2550 , \2548 , \2549 );
xor \U$2174 ( \2551 , \2544 , \2550 );
not \U$2175 ( \2552 , \2084 );
not \U$2176 ( \2553 , \1777 );
or \U$2177 ( \2554 , \2552 , \2553 );
nand \U$2178 ( \2555 , \2554 , \2078 );
not \U$2179 ( \2556 , \664 );
nor \U$2180 ( \2557 , \2556 , \634 );
and \U$2181 ( \2558 , \2555 , \2557 );
not \U$2182 ( \2559 , \2555 );
not \U$2183 ( \2560 , \2557 );
and \U$2184 ( \2561 , \2559 , \2560 );
nor \U$2185 ( \2562 , \2558 , \2561 );
not \U$2186 ( \2563 , \2562 );
buf \U$2187 ( \2564 , \2563 );
not \U$2188 ( \2565 , \2564 );
and \U$2189 ( \2566 , RIae78bc0_126, \2565 );
not \U$2190 ( \2567 , RIae78bc0_126);
and \U$2191 ( \2568 , \2567 , \2564 );
nor \U$2192 ( \2569 , \2566 , \2568 );
not \U$2193 ( \2570 , \2569 );
not \U$2194 ( \2571 , \1036 );
or \U$2195 ( \2572 , \2570 , \2571 );
not \U$2196 ( \2573 , \1789 );
and \U$2197 ( \2574 , \1286 , \2573 );
not \U$2198 ( \2575 , \1286 );
not \U$2199 ( \2576 , \1788 );
not \U$2200 ( \2577 , \2576 );
and \U$2201 ( \2578 , \2575 , \2577 );
nor \U$2202 ( \2579 , \2574 , \2578 );
not \U$2203 ( \2580 , \2579 );
nand \U$2204 ( \2581 , \2580 , \1028 );
nand \U$2205 ( \2582 , \2572 , \2581 );
xnor \U$2206 ( \2583 , \2551 , \2582 );
and \U$2207 ( \2584 , \2533 , \2583 );
not \U$2208 ( \2585 , \2533 );
not \U$2209 ( \2586 , \2583 );
and \U$2210 ( \2587 , \2585 , \2586 );
or \U$2211 ( \2588 , \2584 , \2587 );
not \U$2212 ( \2589 , \1910 );
not \U$2213 ( \2590 , \1881 );
or \U$2214 ( \2591 , \2589 , \2590 );
not \U$2215 ( \2592 , \2047 );
not \U$2216 ( \2593 , \2592 );
buf \U$2217 ( \2594 , \2593 );
not \U$2218 ( \2595 , \2594 );
and \U$2219 ( \2596 , RIae793b8_143, \2595 );
not \U$2220 ( \2597 , RIae793b8_143);
and \U$2221 ( \2598 , \2597 , \2594 );
nor \U$2222 ( \2599 , \2596 , \2598 );
nand \U$2223 ( \2600 , \2599 , \1864 );
nand \U$2224 ( \2601 , \2591 , \2600 );
buf \U$2225 ( \2602 , \2188 );
not \U$2226 ( \2603 , \2602 );
not \U$2227 ( \2604 , \2171 );
or \U$2228 ( \2605 , \2603 , \2604 );
and \U$2229 ( \2606 , \938 , \2183 );
not \U$2230 ( \2607 , \938 );
and \U$2231 ( \2608 , \2607 , RIae79520_146);
nor \U$2232 ( \2609 , \2606 , \2608 );
buf \U$2233 ( \2610 , \2163 );
nand \U$2234 ( \2611 , \2609 , \2610 );
nand \U$2235 ( \2612 , \2605 , \2611 );
xor \U$2236 ( \2613 , \2601 , \2612 );
not \U$2237 ( \2614 , \1499 );
not \U$2238 ( \2615 , \2214 );
or \U$2239 ( \2616 , \2614 , \2615 );
xnor \U$2240 ( \2617 , RIae79250_140, \1899 );
not \U$2241 ( \2618 , \2617 );
nand \U$2242 ( \2619 , \2618 , \1501 );
nand \U$2243 ( \2620 , \2616 , \2619 );
xor \U$2244 ( \2621 , \2613 , \2620 );
xor \U$2245 ( \2622 , \2588 , \2621 );
not \U$2246 ( \2623 , \2622 );
xor \U$2247 ( \2624 , \1978 , \2065 );
xor \U$2248 ( \2625 , \2624 , \2069 );
not \U$2249 ( \2626 , \2625 );
not \U$2250 ( \2627 , \1910 );
buf \U$2251 ( \2628 , \2206 );
not \U$2252 ( \2629 , \2628 );
and \U$2253 ( \2630 , \2629 , \1902 );
not \U$2254 ( \2631 , \2629 );
and \U$2255 ( \2632 , \2631 , RIae793b8_143);
nor \U$2256 ( \2633 , \2630 , \2632 );
not \U$2257 ( \2634 , \2633 );
or \U$2258 ( \2635 , \2627 , \2634 );
nand \U$2259 ( \2636 , \1904 , \1864 );
nand \U$2260 ( \2637 , \2635 , \2636 );
not \U$2261 ( \2638 , \2637 );
not \U$2262 ( \2639 , \2529 );
buf \U$2263 ( \2640 , \1141 );
and \U$2264 ( \2641 , \2640 , RIae797f0_152);
not \U$2265 ( \2642 , \2640 );
and \U$2266 ( \2643 , \2642 , \2521 );
nor \U$2267 ( \2644 , \2641 , \2643 );
not \U$2268 ( \2645 , \2644 );
or \U$2269 ( \2646 , \2639 , \2645 );
nand \U$2270 ( \2647 , \1999 , \2007 );
nand \U$2271 ( \2648 , \2646 , \2647 );
not \U$2272 ( \2649 , \2648 );
buf \U$2273 ( \2650 , \1499 );
not \U$2274 ( \2651 , \2650 );
not \U$2275 ( \2652 , RIae79250_140);
and \U$2276 ( \2653 , \2141 , \2652 );
not \U$2277 ( \2654 , \2141 );
and \U$2278 ( \2655 , \2654 , RIae79250_140);
nor \U$2279 ( \2656 , \2653 , \2655 );
not \U$2280 ( \2657 , \2656 );
or \U$2281 ( \2658 , \2651 , \2657 );
nand \U$2282 ( \2659 , \2235 , \1501 );
nand \U$2283 ( \2660 , \2658 , \2659 );
not \U$2284 ( \2661 , \2660 );
not \U$2285 ( \2662 , \2661 );
or \U$2286 ( \2663 , \2649 , \2662 );
or \U$2287 ( \2664 , \2661 , \2648 );
nand \U$2288 ( \2665 , \2663 , \2664 );
not \U$2289 ( \2666 , \2665 );
or \U$2290 ( \2667 , \2638 , \2666 );
nand \U$2291 ( \2668 , \2660 , \2648 );
nand \U$2292 ( \2669 , \2667 , \2668 );
not \U$2293 ( \2670 , \2669 );
not \U$2294 ( \2671 , \1321 );
not \U$2295 ( \2672 , \1794 );
or \U$2296 ( \2673 , \2671 , \2672 );
not \U$2297 ( \2674 , RIae78e90_132);
buf \U$2298 ( \2675 , \2562 );
not \U$2299 ( \2676 , \2675 );
not \U$2300 ( \2677 , \2676 );
or \U$2301 ( \2678 , \2674 , \2677 );
or \U$2302 ( \2679 , \2676 , RIae78e90_132);
nand \U$2303 ( \2680 , \2678 , \2679 );
nand \U$2304 ( \2681 , \2680 , \1259 );
nand \U$2305 ( \2682 , \2673 , \2681 );
not \U$2306 ( \2683 , \2272 );
not \U$2307 ( \2684 , RIae79ac0_158);
not \U$2308 ( \2685 , \1186 );
or \U$2309 ( \2686 , \2684 , \2685 );
or \U$2310 ( \2687 , \1186 , RIae79ac0_158);
nand \U$2311 ( \2688 , \2686 , \2687 );
not \U$2312 ( \2689 , \2688 );
or \U$2313 ( \2690 , \2683 , \2689 );
nand \U$2314 ( \2691 , \2267 , \2252 );
nand \U$2315 ( \2692 , \2690 , \2691 );
xor \U$2316 ( \2693 , \2682 , \2692 );
not \U$2317 ( \2694 , \797 );
not \U$2318 ( \2695 , RIae78f80_134);
not \U$2319 ( \2696 , \1808 );
buf \U$2320 ( \2697 , \2696 );
not \U$2321 ( \2698 , \2697 );
or \U$2322 ( \2699 , \2695 , \2698 );
or \U$2323 ( \2700 , \2697 , RIae78f80_134);
nand \U$2324 ( \2701 , \2699 , \2700 );
not \U$2325 ( \2702 , \2701 );
or \U$2326 ( \2703 , \2694 , \2702 );
nand \U$2327 ( \2704 , \1762 , \839 );
nand \U$2328 ( \2705 , \2703 , \2704 );
and \U$2329 ( \2706 , \2693 , \2705 );
and \U$2330 ( \2707 , \2682 , \2692 );
nor \U$2331 ( \2708 , \2706 , \2707 );
not \U$2332 ( \2709 , \2708 );
or \U$2333 ( \2710 , \2670 , \2709 );
or \U$2334 ( \2711 , \2669 , \2708 );
nand \U$2335 ( \2712 , \2710 , \2711 );
not \U$2336 ( \2713 , \2712 );
or \U$2337 ( \2714 , \2626 , \2713 );
not \U$2338 ( \2715 , \2708 );
nand \U$2339 ( \2716 , \2715 , \2669 );
nand \U$2340 ( \2717 , \2714 , \2716 );
not \U$2341 ( \2718 , \2717 );
xor \U$2342 ( \2719 , \1764 , \1812 );
xor \U$2343 ( \2720 , \2719 , \1846 );
not \U$2344 ( \2721 , \2720 );
xor \U$2345 ( \2722 , \1861 , \1912 );
xor \U$2346 ( \2723 , \2722 , \1935 );
not \U$2347 ( \2724 , \2723 );
not \U$2348 ( \2725 , \2724 );
not \U$2349 ( \2726 , \2159 );
and \U$2350 ( \2727 , \2238 , \2726 );
not \U$2351 ( \2728 , \2238 );
and \U$2352 ( \2729 , \2728 , \2159 );
nor \U$2353 ( \2730 , \2727 , \2729 );
not \U$2354 ( \2731 , \2730 );
not \U$2355 ( \2732 , \2731 );
or \U$2356 ( \2733 , \2725 , \2732 );
nand \U$2357 ( \2734 , \2730 , \2723 );
nand \U$2358 ( \2735 , \2733 , \2734 );
not \U$2359 ( \2736 , \2735 );
or \U$2360 ( \2737 , \2721 , \2736 );
nand \U$2361 ( \2738 , \2731 , \2723 );
nand \U$2362 ( \2739 , \2737 , \2738 );
not \U$2363 ( \2740 , \2739 );
not \U$2364 ( \2741 , \2740 );
and \U$2365 ( \2742 , \2718 , \2741 );
and \U$2366 ( \2743 , \2717 , \2740 );
nor \U$2367 ( \2744 , \2742 , \2743 );
not \U$2368 ( \2745 , \2744 );
or \U$2369 ( \2746 , \2623 , \2745 );
or \U$2370 ( \2747 , \2744 , \2622 );
nand \U$2371 ( \2748 , \2746 , \2747 );
xor \U$2372 ( \2749 , \2502 , \2748 );
xor \U$2373 ( \2750 , \2682 , \2705 );
xor \U$2374 ( \2751 , \2750 , \2692 );
not \U$2375 ( \2752 , \2751 );
not \U$2376 ( \2753 , \797 );
not \U$2377 ( \2754 , RIae78f80_134);
not \U$2378 ( \2755 , \2577 );
or \U$2379 ( \2756 , \2754 , \2755 );
not \U$2380 ( \2757 , \1789 );
not \U$2381 ( \2758 , \2757 );
not \U$2382 ( \2759 , \2758 );
nand \U$2383 ( \2760 , \2759 , \1132 );
nand \U$2384 ( \2761 , \2756 , \2760 );
not \U$2385 ( \2762 , \2761 );
or \U$2386 ( \2763 , \2753 , \2762 );
nand \U$2387 ( \2764 , \2701 , \839 );
nand \U$2388 ( \2765 , \2763 , \2764 );
not \U$2389 ( \2766 , \2765 );
buf \U$2390 ( \2767 , \2417 );
not \U$2391 ( \2768 , \2767 );
not \U$2392 ( \2769 , \991 );
not \U$2393 ( \2770 , RIae79c28_161);
and \U$2394 ( \2771 , \2769 , \2770 );
and \U$2395 ( \2772 , \991 , RIae79c28_161);
nor \U$2396 ( \2773 , \2771 , \2772 );
not \U$2397 ( \2774 , \2773 );
or \U$2398 ( \2775 , \2768 , \2774 );
buf \U$2399 ( \2776 , \2418 );
nand \U$2400 ( \2777 , \2776 , RIae79c28_161);
nand \U$2401 ( \2778 , \2775 , \2777 );
not \U$2402 ( \2779 , \2778 );
not \U$2403 ( \2780 , \1072 );
not \U$2404 ( \2781 , \2680 );
or \U$2405 ( \2782 , \2780 , \2781 );
and \U$2406 ( \2783 , RIae78e90_132, \2093 );
not \U$2407 ( \2784 , RIae78e90_132);
not \U$2408 ( \2785 , \2088 );
buf \U$2409 ( \2786 , \2785 );
and \U$2410 ( \2787 , \2784 , \2786 );
nor \U$2411 ( \2788 , \2783 , \2787 );
nand \U$2412 ( \2789 , \2788 , \1086 );
nand \U$2413 ( \2790 , \2782 , \2789 );
not \U$2414 ( \2791 , \2790 );
and \U$2415 ( \2792 , \2779 , \2791 );
and \U$2416 ( \2793 , \2778 , \2790 );
nor \U$2417 ( \2794 , \2792 , \2793 );
not \U$2418 ( \2795 , \2794 );
not \U$2419 ( \2796 , \2795 );
or \U$2420 ( \2797 , \2766 , \2796 );
not \U$2421 ( \2798 , \2778 );
nand \U$2422 ( \2799 , \2798 , \2790 );
nand \U$2423 ( \2800 , \2797 , \2799 );
not \U$2424 ( \2801 , \2800 );
not \U$2425 ( \2802 , \2801 );
not \U$2426 ( \2803 , \2637 );
not \U$2427 ( \2804 , \2803 );
not \U$2428 ( \2805 , \2665 );
or \U$2429 ( \2806 , \2804 , \2805 );
not \U$2430 ( \2807 , \2665 );
nand \U$2431 ( \2808 , \2807 , \2637 );
nand \U$2432 ( \2809 , \2806 , \2808 );
not \U$2433 ( \2810 , \2809 );
or \U$2434 ( \2811 , \2802 , \2810 );
or \U$2435 ( \2812 , \2809 , \2801 );
nand \U$2436 ( \2813 , \2811 , \2812 );
not \U$2437 ( \2814 , \2813 );
or \U$2438 ( \2815 , \2752 , \2814 );
nand \U$2439 ( \2816 , \2809 , \2800 );
nand \U$2440 ( \2817 , \2815 , \2816 );
not \U$2441 ( \2818 , \2817 );
not \U$2442 ( \2819 , \2818 );
not \U$2443 ( \2820 , \2480 );
not \U$2444 ( \2821 , \2487 );
and \U$2445 ( \2822 , \2820 , \2821 );
and \U$2446 ( \2823 , \2480 , \2487 );
nor \U$2447 ( \2824 , \2822 , \2823 );
not \U$2448 ( \2825 , \1013 );
and \U$2449 ( \2826 , RIae79160_138, \2305 );
not \U$2450 ( \2827 , RIae79160_138);
and \U$2451 ( \2828 , \2827 , \2310 );
or \U$2452 ( \2829 , \2826 , \2828 );
not \U$2453 ( \2830 , \2829 );
or \U$2454 ( \2831 , \2825 , \2830 );
not \U$2455 ( \2832 , RIae79160_138);
not \U$2456 ( \2833 , \2287 );
or \U$2457 ( \2834 , \2832 , \2833 );
buf \U$2458 ( \2835 , \2285 );
buf \U$2459 ( \2836 , \2835 );
or \U$2460 ( \2837 , \2836 , RIae79160_138);
nand \U$2461 ( \2838 , \2834 , \2837 );
nand \U$2462 ( \2839 , \2838 , \1009 );
nand \U$2463 ( \2840 , \2831 , \2839 );
not \U$2464 ( \2841 , \2840 );
not \U$2465 ( \2842 , \2252 );
not \U$2466 ( \2843 , \2688 );
or \U$2467 ( \2844 , \2842 , \2843 );
and \U$2468 ( \2845 , RIae79ac0_158, \1405 );
not \U$2469 ( \2846 , RIae79ac0_158);
not \U$2470 ( \2847 , \1403 );
not \U$2471 ( \2848 , \2847 );
not \U$2472 ( \2849 , \2848 );
not \U$2473 ( \2850 , \2849 );
and \U$2474 ( \2851 , \2846 , \2850 );
or \U$2475 ( \2852 , \2845 , \2851 );
nand \U$2476 ( \2853 , \2852 , \2272 );
nand \U$2477 ( \2854 , \2844 , \2853 );
not \U$2478 ( \2855 , \2854 );
or \U$2479 ( \2856 , \2841 , \2855 );
buf \U$2480 ( \2857 , \1739 );
not \U$2481 ( \2858 , \2857 );
and \U$2482 ( \2859 , \2858 , RIae79070_136);
not \U$2483 ( \2860 , \2858 );
and \U$2484 ( \2861 , \2860 , \1039 );
nor \U$2485 ( \2862 , \2859 , \2861 );
and \U$2486 ( \2863 , \2862 , \1049 );
xnor \U$2487 ( \2864 , \1760 , RIae79070_136);
and \U$2488 ( \2865 , \2864 , \1062 );
nor \U$2489 ( \2866 , \2863 , \2865 );
nand \U$2490 ( \2867 , \2856 , \2866 );
or \U$2491 ( \2868 , \2854 , \2840 );
nand \U$2492 ( \2869 , \2867 , \2868 );
nand \U$2493 ( \2870 , \2824 , \2869 );
not \U$2494 ( \2871 , \2870 );
xor \U$2495 ( \2872 , \2370 , \2380 );
xor \U$2496 ( \2873 , \2872 , \2389 );
not \U$2497 ( \2874 , \2873 );
or \U$2498 ( \2875 , \2871 , \2874 );
not \U$2499 ( \2876 , \2824 );
not \U$2500 ( \2877 , \2869 );
nand \U$2501 ( \2878 , \2876 , \2877 );
nand \U$2502 ( \2879 , \2875 , \2878 );
nor \U$2503 ( \2880 , \2819 , \2879 );
not \U$2504 ( \2881 , \2720 );
and \U$2505 ( \2882 , \2735 , \2881 );
not \U$2506 ( \2883 , \2735 );
and \U$2507 ( \2884 , \2883 , \2720 );
nor \U$2508 ( \2885 , \2882 , \2884 );
or \U$2509 ( \2886 , \2880 , \2885 );
not \U$2510 ( \2887 , \2879 );
or \U$2511 ( \2888 , \2818 , \2887 );
nand \U$2512 ( \2889 , \2886 , \2888 );
and \U$2513 ( \2890 , \2749 , \2889 );
and \U$2514 ( \2891 , \2502 , \2748 );
or \U$2515 ( \2892 , \2890 , \2891 );
not \U$2516 ( \2893 , \2892 );
xor \U$2517 ( \2894 , \2072 , \2348 );
and \U$2518 ( \2895 , \2894 , \2501 );
and \U$2519 ( \2896 , \2072 , \2348 );
or \U$2520 ( \2897 , \2895 , \2896 );
not \U$2521 ( \2898 , \1027 );
not \U$2522 ( \2899 , \2569 );
or \U$2523 ( \2900 , \2898 , \2899 );
nand \U$2524 ( \2901 , \1036 , \2368 );
nand \U$2525 ( \2902 , \2900 , \2901 );
buf \U$2526 ( \2903 , \2550 );
not \U$2527 ( \2904 , \2903 );
xor \U$2528 ( \2905 , \2902 , \2904 );
not \U$2529 ( \2906 , \2905 );
not \U$2530 ( \2907 , \1209 );
not \U$2531 ( \2908 , \2156 );
or \U$2532 ( \2909 , \2907 , \2908 );
nand \U$2533 ( \2910 , \2829 , \1009 );
nand \U$2534 ( \2911 , \2909 , \2910 );
not \U$2535 ( \2912 , \2911 );
not \U$2536 ( \2913 , \2602 );
not \U$2537 ( \2914 , RIae79520_146);
not \U$2538 ( \2915 , \1472 );
or \U$2539 ( \2916 , \2914 , \2915 );
buf \U$2540 ( \2917 , \1117 );
not \U$2541 ( \2918 , \2917 );
or \U$2542 ( \2919 , \2918 , RIae79520_146);
nand \U$2543 ( \2920 , \2916 , \2919 );
not \U$2544 ( \2921 , \2920 );
or \U$2545 ( \2922 , \2913 , \2921 );
not \U$2546 ( \2923 , \2163 );
not \U$2547 ( \2924 , \2923 );
nand \U$2548 ( \2925 , \2181 , \2924 );
nand \U$2549 ( \2926 , \2922 , \2925 );
not \U$2550 ( \2927 , \1049 );
not \U$2551 ( \2928 , \2291 );
or \U$2552 ( \2929 , \2927 , \2928 );
nand \U$2553 ( \2930 , \2862 , \2276 );
nand \U$2554 ( \2931 , \2929 , \2930 );
xor \U$2555 ( \2932 , \2926 , \2931 );
not \U$2556 ( \2933 , \2932 );
or \U$2557 ( \2934 , \2912 , \2933 );
buf \U$2558 ( \2935 , \2926 );
nand \U$2559 ( \2936 , \2935 , \2931 );
nand \U$2560 ( \2937 , \2934 , \2936 );
not \U$2561 ( \2938 , \2937 );
or \U$2562 ( \2939 , \2906 , \2938 );
not \U$2563 ( \2940 , \2903 );
nand \U$2564 ( \2941 , \2940 , \2902 );
nand \U$2565 ( \2942 , \2939 , \2941 );
not \U$2566 ( \2943 , \2942 );
not \U$2567 ( \2944 , \797 );
not \U$2568 ( \2945 , \1743 );
or \U$2569 ( \2946 , \2944 , \2945 );
and \U$2570 ( \2947 , \2287 , \1132 );
not \U$2571 ( \2948 , \2287 );
and \U$2572 ( \2949 , \2948 , RIae78f80_134);
nor \U$2573 ( \2950 , \2947 , \2949 );
nand \U$2574 ( \2951 , \2950 , \839 );
nand \U$2575 ( \2952 , \2946 , \2951 );
not \U$2576 ( \2953 , \1049 );
buf \U$2577 ( \2954 , \2152 );
not \U$2578 ( \2955 , \2954 );
not \U$2579 ( \2956 , \2955 );
and \U$2580 ( \2957 , \2956 , \1039 );
not \U$2581 ( \2958 , \2956 );
and \U$2582 ( \2959 , \2958 , RIae79070_136);
nor \U$2583 ( \2960 , \2957 , \2959 );
not \U$2584 ( \2961 , \2960 );
or \U$2585 ( \2962 , \2953 , \2961 );
nand \U$2586 ( \2963 , \2312 , \1062 );
nand \U$2587 ( \2964 , \2962 , \2963 );
xor \U$2588 ( \2965 , \2952 , \2964 );
buf \U$2589 ( \2966 , \1843 );
not \U$2590 ( \2967 , \2966 );
not \U$2591 ( \2968 , \1828 );
or \U$2592 ( \2969 , \2967 , \2968 );
not \U$2593 ( \2970 , RIae79688_149);
and \U$2594 ( \2971 , \978 , \2970 );
not \U$2595 ( \2972 , \978 );
and \U$2596 ( \2973 , \2972 , RIae79688_149);
nor \U$2597 ( \2974 , \2971 , \2973 );
nand \U$2598 ( \2975 , \2974 , \1822 );
nand \U$2599 ( \2976 , \2969 , \2975 );
xor \U$2600 ( \2977 , \2965 , \2976 );
not \U$2601 ( \2978 , \2341 );
not \U$2602 ( \2979 , \2325 );
or \U$2603 ( \2980 , \2978 , \2979 );
not \U$2604 ( \2981 , RIae798e0_154);
not \U$2605 ( \2982 , \2981 );
not \U$2606 ( \2983 , \781 );
or \U$2607 ( \2984 , \2982 , \2983 );
nand \U$2608 ( \2985 , \1993 , RIae798e0_154);
nand \U$2609 ( \2986 , \2984 , \2985 );
nand \U$2610 ( \2987 , \2986 , \2322 );
nand \U$2611 ( \2988 , \2980 , \2987 );
not \U$2612 ( \2989 , \1430 );
not \U$2613 ( \2990 , \2144 );
or \U$2614 ( \2991 , \2989 , \2990 );
not \U$2615 ( \2992 , \997 );
buf \U$2616 ( \2993 , \2229 );
not \U$2617 ( \2994 , \2993 );
buf \U$2618 ( \2995 , \2994 );
not \U$2619 ( \2996 , \2995 );
or \U$2620 ( \2997 , \2992 , \2996 );
nand \U$2621 ( \2998 , \2993 , RIae79160_138);
nand \U$2622 ( \2999 , \2997 , \2998 );
nand \U$2623 ( \3000 , \2999 , \1209 );
nand \U$2624 ( \3001 , \2991 , \3000 );
and \U$2625 ( \3002 , \2988 , \3001 );
not \U$2626 ( \3003 , \2988 );
not \U$2627 ( \3004 , \3001 );
and \U$2628 ( \3005 , \3003 , \3004 );
nor \U$2629 ( \3006 , \3002 , \3005 );
not \U$2630 ( \3007 , \2272 );
not \U$2631 ( \3008 , \2258 );
or \U$2632 ( \3009 , \3007 , \3008 );
and \U$2633 ( \3010 , \2268 , \883 );
not \U$2634 ( \3011 , \2268 );
and \U$2635 ( \3012 , \3011 , \879 );
nor \U$2636 ( \3013 , \3010 , \3012 );
buf \U$2637 ( \3014 , \2249 );
buf \U$2638 ( \3015 , \3014 );
not \U$2639 ( \3016 , \3015 );
or \U$2640 ( \3017 , \3013 , \3016 );
nand \U$2641 ( \3018 , \3009 , \3017 );
not \U$2642 ( \3019 , \3018 );
and \U$2643 ( \3020 , \3006 , \3019 );
not \U$2644 ( \3021 , \3006 );
and \U$2645 ( \3022 , \3021 , \3018 );
nor \U$2646 ( \3023 , \3020 , \3022 );
or \U$2647 ( \3024 , \2977 , \3023 );
nand \U$2648 ( \3025 , \3023 , \2977 );
nand \U$2649 ( \3026 , \3024 , \3025 );
not \U$2650 ( \3027 , \3026 );
or \U$2651 ( \3028 , \2943 , \3027 );
not \U$2652 ( \3029 , \3023 );
nand \U$2653 ( \3030 , \3029 , \2977 );
nand \U$2654 ( \3031 , \3028 , \3030 );
not \U$2655 ( \3032 , \3031 );
not \U$2656 ( \3033 , \3032 );
and \U$2657 ( \3034 , \2551 , \2582 );
and \U$2658 ( \3035 , \2544 , \2550 );
nor \U$2659 ( \3036 , \3034 , \3035 );
not \U$2660 ( \3037 , \3036 );
not \U$2661 ( \3038 , \1919 );
not \U$2662 ( \3039 , RIae794a8_145);
and \U$2663 ( \3040 , \2324 , \3039 );
not \U$2664 ( \3041 , \2324 );
and \U$2665 ( \3042 , \3041 , RIae794a8_145);
nor \U$2666 ( \3043 , \3040 , \3042 );
not \U$2667 ( \3044 , \3043 );
or \U$2668 ( \3045 , \3038 , \3044 );
nand \U$2669 ( \3046 , \2514 , \1933 );
nand \U$2670 ( \3047 , \3045 , \3046 );
not \U$2671 ( \3048 , \3047 );
not \U$2672 ( \3049 , \3048 );
not \U$2673 ( \3050 , \1209 );
not \U$2674 ( \3051 , \2207 );
buf \U$2675 ( \3052 , \3051 );
and \U$2676 ( \3053 , RIae79160_138, \3052 );
not \U$2677 ( \3054 , RIae79160_138);
not \U$2678 ( \3055 , \2212 );
and \U$2679 ( \3056 , \3054 , \3055 );
or \U$2680 ( \3057 , \3053 , \3056 );
not \U$2681 ( \3058 , \3057 );
or \U$2682 ( \3059 , \3050 , \3058 );
nand \U$2683 ( \3060 , \2999 , \1010 );
nand \U$2684 ( \3061 , \3059 , \3060 );
not \U$2685 ( \3062 , \3061 );
or \U$2686 ( \3063 , \3049 , \3062 );
or \U$2687 ( \3064 , \3061 , \3048 );
nand \U$2688 ( \3065 , \3063 , \3064 );
not \U$2689 ( \3066 , \3065 );
not \U$2690 ( \3067 , \1049 );
not \U$2691 ( \3068 , RIae79070_136);
buf \U$2692 ( \3069 , \2134 );
not \U$2693 ( \3070 , \3069 );
not \U$2694 ( \3071 , \3070 );
buf \U$2695 ( \3072 , \3071 );
not \U$2696 ( \3073 , \3072 );
or \U$2697 ( \3074 , \3068 , \3073 );
nand \U$2698 ( \3075 , \2142 , \1039 );
nand \U$2699 ( \3076 , \3074 , \3075 );
not \U$2700 ( \3077 , \3076 );
or \U$2701 ( \3078 , \3067 , \3077 );
nand \U$2702 ( \3079 , \2960 , \1062 );
nand \U$2703 ( \3080 , \3078 , \3079 );
not \U$2704 ( \3081 , \3080 );
not \U$2705 ( \3082 , \3081 );
and \U$2706 ( \3083 , \3066 , \3082 );
and \U$2707 ( \3084 , \3065 , \3081 );
nor \U$2708 ( \3085 , \3083 , \3084 );
not \U$2709 ( \3086 , \3085 );
not \U$2710 ( \3087 , \3086 );
or \U$2711 ( \3088 , \3037 , \3087 );
not \U$2712 ( \3089 , \3036 );
nand \U$2713 ( \3090 , \3089 , \3085 );
nand \U$2714 ( \3091 , \3088 , \3090 );
buf \U$2715 ( \3092 , \1738 );
not \U$2716 ( \3093 , \3092 );
buf \U$2717 ( \3094 , \3093 );
not \U$2718 ( \3095 , \3094 );
and \U$2719 ( \3096 , RIae78e90_132, \3095 );
not \U$2720 ( \3097 , RIae78e90_132);
buf \U$2721 ( \3098 , \3092 );
not \U$2722 ( \3099 , \3098 );
and \U$2723 ( \3100 , \3097 , \3099 );
nor \U$2724 ( \3101 , \3096 , \3100 );
or \U$2725 ( \3102 , \3101 , \1073 );
or \U$2726 ( \3103 , \2541 , \1313 );
nand \U$2727 ( \3104 , \3102 , \3103 );
not \U$2728 ( \3105 , RIae78f80_134);
not \U$2729 ( \3106 , \3105 );
not \U$2730 ( \3107 , \2309 );
or \U$2731 ( \3108 , \3106 , \3107 );
nand \U$2732 ( \3109 , \2305 , RIae78f80_134);
nand \U$2733 ( \3110 , \3108 , \3109 );
not \U$2734 ( \3111 , \3110 );
not \U$2735 ( \3112 , \839 );
or \U$2736 ( \3113 , \3111 , \3112 );
not \U$2737 ( \3114 , \2950 );
or \U$2738 ( \3115 , \3114 , \798 );
nand \U$2739 ( \3116 , \3113 , \3115 );
xor \U$2740 ( \3117 , \3104 , \3116 );
not \U$2741 ( \3118 , \1822 );
xor \U$2742 ( \3119 , \1473 , RIae79688_149);
not \U$2743 ( \3120 , \3119 );
or \U$2744 ( \3121 , \3118 , \3120 );
nand \U$2745 ( \3122 , \2974 , \2966 );
nand \U$2746 ( \3123 , \3121 , \3122 );
xor \U$2747 ( \3124 , \3117 , \3123 );
not \U$2748 ( \3125 , \3124 );
and \U$2749 ( \3126 , \3091 , \3125 );
not \U$2750 ( \3127 , \3091 );
and \U$2751 ( \3128 , \3127 , \3124 );
nor \U$2752 ( \3129 , \3126 , \3128 );
not \U$2753 ( \3130 , \3129 );
not \U$2754 ( \3131 , \3130 );
or \U$2755 ( \3132 , \3033 , \3131 );
nand \U$2756 ( \3133 , \3129 , \3031 );
nand \U$2757 ( \3134 , \3132 , \3133 );
xnor \U$2758 ( \3135 , \2897 , \3134 );
not \U$2759 ( \3136 , \3135 );
not \U$2760 ( \3137 , \1822 );
not \U$2761 ( \3138 , \2378 );
or \U$2762 ( \3139 , \3137 , \3138 );
not \U$2763 ( \3140 , RIae79688_149);
not \U$2764 ( \3141 , \2592 );
not \U$2765 ( \3142 , \3141 );
or \U$2766 ( \3143 , \3140 , \3142 );
not \U$2767 ( \3144 , \2046 );
not \U$2768 ( \3145 , \3144 );
not \U$2769 ( \3146 , \3145 );
not \U$2770 ( \3147 , RIae79688_149);
nand \U$2771 ( \3148 , \3146 , \3147 );
nand \U$2772 ( \3149 , \3143 , \3148 );
nand \U$2773 ( \3150 , \3149 , \2966 );
nand \U$2774 ( \3151 , \3139 , \3150 );
not \U$2775 ( \3152 , \3151 );
nand \U$2776 ( \3153 , \607 , \609 );
not \U$2777 ( \3154 , \3153 );
buf \U$2778 ( \3155 , \470 );
and \U$2779 ( \3156 , \472 , \3155 );
buf \U$2780 ( \3157 , \475 );
and \U$2781 ( \3158 , \3156 , \3157 );
not \U$2782 ( \3159 , \3158 );
not \U$2783 ( \3160 , \486 );
nor \U$2784 ( \3161 , \3160 , \464 );
not \U$2785 ( \3162 , \3161 );
not \U$2786 ( \3163 , \562 );
not \U$2787 ( \3164 , \515 );
nor \U$2788 ( \3165 , \3163 , \3164 );
not \U$2789 ( \3166 , \3165 );
not \U$2790 ( \3167 , \558 );
and \U$2791 ( \3168 , \427 , \435 , \419 );
nor \U$2792 ( \3169 , \3168 , \452 );
nand \U$2793 ( \3170 , \3167 , \3169 );
not \U$2794 ( \3171 , \3170 );
or \U$2795 ( \3172 , \3166 , \3171 );
not \U$2796 ( \3173 , \491 );
not \U$2797 ( \3174 , \460 );
not \U$2798 ( \3175 , \3174 );
and \U$2799 ( \3176 , \3173 , \3175 );
nor \U$2800 ( \3177 , \3176 , \462 );
not \U$2801 ( \3178 , \3177 );
or \U$2802 ( \3179 , \3178 , \3164 );
not \U$2803 ( \3180 , \583 );
nand \U$2804 ( \3181 , \3179 , \3180 );
not \U$2805 ( \3182 , \3181 );
nand \U$2806 ( \3183 , \3172 , \3182 );
not \U$2807 ( \3184 , \3183 );
or \U$2808 ( \3185 , \3162 , \3184 );
not \U$2809 ( \3186 , \464 );
not \U$2810 ( \3187 , \3186 );
buf \U$2811 ( \3188 , \485 );
not \U$2812 ( \3189 , \3188 );
buf \U$2813 ( \3190 , \592 );
not \U$2814 ( \3191 , \3190 );
or \U$2815 ( \3192 , \3189 , \3191 );
nand \U$2816 ( \3193 , \3192 , \585 );
not \U$2817 ( \3194 , \3193 );
or \U$2818 ( \3195 , \3187 , \3194 );
nand \U$2819 ( \3196 , \3195 , \586 );
not \U$2820 ( \3197 , \3196 );
nand \U$2821 ( \3198 , \3185 , \3197 );
not \U$2822 ( \3199 , \3198 );
or \U$2823 ( \3200 , \3159 , \3199 );
not \U$2824 ( \3201 , \606 );
nand \U$2825 ( \3202 , \3200 , \3201 );
not \U$2826 ( \3203 , \3202 );
or \U$2827 ( \3204 , \3154 , \3203 );
or \U$2828 ( \3205 , \3153 , \3202 );
nand \U$2829 ( \3206 , \3204 , \3205 );
buf \U$2830 ( \3207 , \3206 );
buf \U$2831 ( \3208 , \3207 );
and \U$2832 ( \3209 , RIae78b48_125, \3208 );
not \U$2833 ( \3210 , \3209 );
not \U$2834 ( \3211 , \1027 );
not \U$2835 ( \3212 , \2362 );
or \U$2836 ( \3213 , \3211 , \3212 );
and \U$2837 ( \3214 , RIae78bc0_126, \1970 );
not \U$2838 ( \3215 , RIae78bc0_126);
buf \U$2839 ( \3216 , \1968 );
not \U$2840 ( \3217 , \3216 );
and \U$2841 ( \3218 , \3215 , \3217 );
or \U$2842 ( \3219 , \3214 , \3218 );
nand \U$2843 ( \3220 , \3219 , \951 );
nand \U$2844 ( \3221 , \3213 , \3220 );
not \U$2845 ( \3222 , \3221 );
not \U$2846 ( \3223 , \3222 );
or \U$2847 ( \3224 , \3210 , \3223 );
or \U$2848 ( \3225 , \3222 , \3209 );
nand \U$2849 ( \3226 , \3224 , \3225 );
not \U$2850 ( \3227 , \3226 );
or \U$2851 ( \3228 , \3152 , \3227 );
not \U$2852 ( \3229 , \3222 );
nand \U$2853 ( \3230 , \3229 , \3209 );
nand \U$2854 ( \3231 , \3228 , \3230 );
not \U$2855 ( \3232 , \2322 );
not \U$2856 ( \3233 , \2475 );
or \U$2857 ( \3234 , \3232 , \3233 );
buf \U$2858 ( \3235 , \936 );
not \U$2859 ( \3236 , \3235 );
xor \U$2860 ( \3237 , RIae798e0_154, \3236 );
nand \U$2861 ( \3238 , \3237 , \2341 );
nand \U$2862 ( \3239 , \3234 , \3238 );
not \U$2863 ( \3240 , \1864 );
not \U$2864 ( \3241 , \2633 );
or \U$2865 ( \3242 , \3240 , \3241 );
not \U$2866 ( \3243 , \1902 );
buf \U$2867 ( \3244 , \2230 );
not \U$2868 ( \3245 , \3244 );
not \U$2869 ( \3246 , \3245 );
or \U$2870 ( \3247 , \3243 , \3246 );
nand \U$2871 ( \3248 , \3244 , RIae793b8_143);
nand \U$2872 ( \3249 , \3247 , \3248 );
nand \U$2873 ( \3250 , \3249 , \1910 );
nand \U$2874 ( \3251 , \3242 , \3250 );
xor \U$2875 ( \3252 , \3239 , \3251 );
not \U$2876 ( \3253 , \1919 );
not \U$2877 ( \3254 , \2464 );
or \U$2878 ( \3255 , \3253 , \3254 );
not \U$2879 ( \3256 , \2179 );
and \U$2880 ( \3257 , RIae794a8_145, \3256 );
not \U$2881 ( \3258 , RIae794a8_145);
and \U$2882 ( \3259 , \3258 , \884 );
nor \U$2883 ( \3260 , \3257 , \3259 );
nand \U$2884 ( \3261 , \3260 , \2458 );
nand \U$2885 ( \3262 , \3255 , \3261 );
and \U$2886 ( \3263 , \3252 , \3262 );
and \U$2887 ( \3264 , \3239 , \3251 );
or \U$2888 ( \3265 , \3263 , \3264 );
xor \U$2889 ( \3266 , \3231 , \3265 );
not \U$2890 ( \3267 , \2096 );
or \U$2891 ( \3268 , \2387 , \3267 );
not \U$2892 ( \3269 , \2401 );
not \U$2893 ( \3270 , \3269 );
and \U$2894 ( \3271 , RIae78b48_125, \3270 );
not \U$2895 ( \3272 , RIae78b48_125);
not \U$2896 ( \3273 , \2402 );
and \U$2897 ( \3274 , \3272 , \3273 );
nor \U$2898 ( \3275 , \3271 , \3274 );
or \U$2899 ( \3276 , \3275 , \1976 );
nand \U$2900 ( \3277 , \3268 , \3276 );
not \U$2901 ( \3278 , \3277 );
not \U$2902 ( \3279 , \2450 );
not \U$2903 ( \3280 , \2439 );
or \U$2904 ( \3281 , \3279 , \3280 );
not \U$2905 ( \3282 , \2442 );
not \U$2906 ( \3283 , \1993 );
not \U$2907 ( \3284 , \3283 );
or \U$2908 ( \3285 , \3282 , \3284 );
not \U$2909 ( \3286 , \3283 );
nand \U$2910 ( \3287 , \3286 , RIae79778_151);
nand \U$2911 ( \3288 , \3285 , \3287 );
nand \U$2912 ( \3289 , \3288 , \2545 );
nand \U$2913 ( \3290 , \3281 , \3289 );
not \U$2914 ( \3291 , \2011 );
not \U$2915 ( \3292 , \2485 );
or \U$2916 ( \3293 , \3291 , \3292 );
buf \U$2917 ( \3294 , \1897 );
xor \U$2918 ( \3295 , RIae79610_148, \3294 );
nand \U$2919 ( \3296 , \3295 , \2063 );
nand \U$2920 ( \3297 , \3293 , \3296 );
or \U$2921 ( \3298 , \3290 , \3297 );
not \U$2922 ( \3299 , \3298 );
or \U$2923 ( \3300 , \3278 , \3299 );
nand \U$2924 ( \3301 , \3290 , \3297 );
nand \U$2925 ( \3302 , \3300 , \3301 );
and \U$2926 ( \3303 , \3266 , \3302 );
and \U$2927 ( \3304 , \3231 , \3265 );
or \U$2928 ( \3305 , \3303 , \3304 );
xor \U$2929 ( \3306 , \2455 , \2392 );
xnor \U$2930 ( \3307 , \3306 , \2491 );
xor \U$2931 ( \3308 , \3305 , \3307 );
xor \U$2932 ( \3309 , \2625 , \2712 );
and \U$2933 ( \3310 , \3308 , \3309 );
and \U$2934 ( \3311 , \3305 , \3307 );
nor \U$2935 ( \3312 , \3310 , \3311 );
not \U$2936 ( \3313 , \3312 );
not \U$2937 ( \3314 , \3313 );
not \U$2938 ( \3315 , \2452 );
not \U$2939 ( \3316 , \2421 );
and \U$2940 ( \3317 , \3315 , \3316 );
and \U$2941 ( \3318 , \2452 , \2421 );
nor \U$2942 ( \3319 , \3317 , \3318 );
nor \U$2943 ( \3320 , \3319 , \2798 );
not \U$2944 ( \3321 , \2007 );
not \U$2945 ( \3322 , \2644 );
or \U$2946 ( \3323 , \3321 , \3322 );
and \U$2947 ( \3324 , RIae797f0_152, \2330 );
not \U$2948 ( \3325 , RIae797f0_152);
buf \U$2949 ( \3326 , \1288 );
and \U$2950 ( \3327 , \3325 , \3326 );
nor \U$2951 ( \3328 , \3324 , \3327 );
nand \U$2952 ( \3329 , \3328 , \1989 );
nand \U$2953 ( \3330 , \3323 , \3329 );
not \U$2954 ( \3331 , \3330 );
not \U$2955 ( \3332 , \3331 );
not \U$2956 ( \3333 , \1501 );
not \U$2957 ( \3334 , \2656 );
or \U$2958 ( \3335 , \3333 , \3334 );
not \U$2959 ( \3336 , \1503 );
not \U$2960 ( \3337 , \2955 );
or \U$2961 ( \3338 , \3336 , \3337 );
nand \U$2962 ( \3339 , \2155 , RIae79250_140);
nand \U$2963 ( \3340 , \3338 , \3339 );
nand \U$2964 ( \3341 , \3340 , \1499 );
nand \U$2965 ( \3342 , \3335 , \3341 );
not \U$2966 ( \3343 , \3342 );
not \U$2967 ( \3344 , \3343 );
or \U$2968 ( \3345 , \3332 , \3344 );
not \U$2969 ( \3346 , \2163 );
not \U$2970 ( \3347 , \2920 );
or \U$2971 ( \3348 , \3346 , \3347 );
not \U$2972 ( \3349 , \2183 );
not \U$2973 ( \3350 , \2262 );
or \U$2974 ( \3351 , \3349 , \3350 );
nand \U$2975 ( \3352 , \2263 , RIae79520_146);
nand \U$2976 ( \3353 , \3351 , \3352 );
nand \U$2977 ( \3354 , \3353 , \2189 );
nand \U$2978 ( \3355 , \3348 , \3354 );
nand \U$2979 ( \3356 , \3345 , \3355 );
nand \U$2980 ( \3357 , \3342 , \3330 );
nand \U$2981 ( \3358 , \3356 , \3357 );
or \U$2982 ( \3359 , \3320 , \3358 );
nand \U$2983 ( \3360 , \3319 , \2798 );
nand \U$2984 ( \3361 , \3359 , \3360 );
xnor \U$2985 ( \3362 , \2343 , \2318 );
and \U$2986 ( \3363 , \3361 , \3362 );
xnor \U$2987 ( \3364 , \2937 , \2905 );
or \U$2988 ( \3365 , \3363 , \3364 );
or \U$2989 ( \3366 , \3361 , \3362 );
nand \U$2990 ( \3367 , \3365 , \3366 );
not \U$2991 ( \3368 , \2942 );
and \U$2992 ( \3369 , \3026 , \3368 );
not \U$2993 ( \3370 , \3026 );
and \U$2994 ( \3371 , \3370 , \2942 );
nor \U$2995 ( \3372 , \3369 , \3371 );
xnor \U$2996 ( \3373 , \3367 , \3372 );
not \U$2997 ( \3374 , \3373 );
or \U$2998 ( \3375 , \3314 , \3374 );
not \U$2999 ( \3376 , \3372 );
nand \U$3000 ( \3377 , \3376 , \3367 );
nand \U$3001 ( \3378 , \3375 , \3377 );
not \U$3002 ( \3379 , \3378 );
or \U$3003 ( \3380 , \3136 , \3379 );
or \U$3004 ( \3381 , \3378 , \3135 );
nand \U$3005 ( \3382 , \3380 , \3381 );
not \U$3006 ( \3383 , \3382 );
or \U$3007 ( \3384 , \2893 , \3383 );
not \U$3008 ( \3385 , \3135 );
nand \U$3009 ( \3386 , \3385 , \3378 );
nand \U$3010 ( \3387 , \3384 , \3386 );
not \U$3011 ( \3388 , \3387 );
not \U$3012 ( \3389 , \3388 );
xor \U$3013 ( \3390 , \2952 , \2964 );
and \U$3014 ( \3391 , \3390 , \2976 );
and \U$3015 ( \3392 , \2952 , \2964 );
or \U$3016 ( \3393 , \3391 , \3392 );
xor \U$3017 ( \3394 , \2601 , \2612 );
and \U$3018 ( \3395 , \3394 , \2620 );
and \U$3019 ( \3396 , \2601 , \2612 );
or \U$3020 ( \3397 , \3395 , \3396 );
xor \U$3021 ( \3398 , \3393 , \3397 );
not \U$3022 ( \3399 , \2988 );
not \U$3023 ( \3400 , \3001 );
or \U$3024 ( \3401 , \3399 , \3400 );
or \U$3025 ( \3402 , \3001 , \2988 );
nand \U$3026 ( \3403 , \3402 , \3018 );
nand \U$3027 ( \3404 , \3401 , \3403 );
and \U$3028 ( \3405 , \3398 , \3404 );
and \U$3029 ( \3406 , \3393 , \3397 );
or \U$3030 ( \3407 , \3405 , \3406 );
not \U$3031 ( \3408 , \3407 );
not \U$3032 ( \3409 , \868 );
xor \U$3033 ( \3410 , RIae78b48_125, \2573 );
not \U$3034 ( \3411 , \3410 );
or \U$3035 ( \3412 , \3409 , \3411 );
and \U$3036 ( \3413 , \2555 , \2557 );
not \U$3037 ( \3414 , \2555 );
and \U$3038 ( \3415 , \3414 , \2560 );
or \U$3039 ( \3416 , \3413 , \3415 );
buf \U$3040 ( \3417 , \3416 );
xnor \U$3041 ( \3418 , \3417 , RIae78b48_125);
not \U$3042 ( \3419 , \3418 );
or \U$3043 ( \3420 , \3419 , \1128 );
nand \U$3044 ( \3421 , \3412 , \3420 );
not \U$3045 ( \3422 , \1989 );
not \U$3046 ( \3423 , \2526 );
or \U$3047 ( \3424 , \3422 , \3423 );
nand \U$3048 ( \3425 , \2007 , RIae797f0_152);
nand \U$3049 ( \3426 , \3424 , \3425 );
xor \U$3050 ( \3427 , \3421 , \3426 );
not \U$3051 ( \3428 , \2322 );
and \U$3052 ( \3429 , RIae798e0_154, \1424 );
not \U$3053 ( \3430 , RIae798e0_154);
not \U$3054 ( \3431 , \2004 );
and \U$3055 ( \3432 , \3430 , \3431 );
nor \U$3056 ( \3433 , \3429 , \3432 );
not \U$3057 ( \3434 , \3433 );
or \U$3058 ( \3435 , \3428 , \3434 );
nand \U$3059 ( \3436 , \2986 , \2341 );
nand \U$3060 ( \3437 , \3435 , \3436 );
not \U$3061 ( \3438 , \3437 );
and \U$3062 ( \3439 , RIae78b48_125, \1956 );
buf \U$3063 ( \3440 , \2163 );
not \U$3064 ( \3441 , \3440 );
not \U$3065 ( \3442 , RIae79520_146);
not \U$3066 ( \3443 , \918 );
not \U$3067 ( \3444 , \3443 );
or \U$3068 ( \3445 , \3442 , \3444 );
or \U$3069 ( \3446 , \3443 , RIae79520_146);
nand \U$3070 ( \3447 , \3445 , \3446 );
not \U$3071 ( \3448 , \3447 );
or \U$3072 ( \3449 , \3441 , \3448 );
nand \U$3073 ( \3450 , \2609 , \2189 );
nand \U$3074 ( \3451 , \3449 , \3450 );
xor \U$3075 ( \3452 , \3439 , \3451 );
not \U$3076 ( \3453 , \3452 );
or \U$3077 ( \3454 , \3438 , \3453 );
nand \U$3078 ( \3455 , \3451 , \3439 );
nand \U$3079 ( \3456 , \3454 , \3455 );
xor \U$3080 ( \3457 , \3427 , \3456 );
not \U$3081 ( \3458 , \3457 );
not \U$3082 ( \3459 , \2516 );
not \U$3083 ( \3460 , \2531 );
nand \U$3084 ( \3461 , \3460 , \2505 );
not \U$3085 ( \3462 , \3461 );
or \U$3086 ( \3463 , \3459 , \3462 );
nand \U$3087 ( \3464 , \2531 , \2506 );
nand \U$3088 ( \3465 , \3463 , \3464 );
not \U$3089 ( \3466 , \3426 );
or \U$3090 ( \3467 , \3465 , \3466 );
not \U$3091 ( \3468 , \3465 );
not \U$3092 ( \3469 , \3466 );
or \U$3093 ( \3470 , \3468 , \3469 );
xor \U$3094 ( \3471 , \2073 , \2098 );
and \U$3095 ( \3472 , \3471 , \2110 );
and \U$3096 ( \3473 , \2073 , \2098 );
or \U$3097 ( \3474 , \3472 , \3473 );
not \U$3098 ( \3475 , \3474 );
nand \U$3099 ( \3476 , \3470 , \3475 );
nand \U$3100 ( \3477 , \3467 , \3476 );
not \U$3101 ( \3478 , \3477 );
or \U$3102 ( \3479 , \3458 , \3478 );
or \U$3103 ( \3480 , \3477 , \3457 );
nand \U$3104 ( \3481 , \3479 , \3480 );
not \U$3105 ( \3482 , \3481 );
or \U$3106 ( \3483 , \3408 , \3482 );
or \U$3107 ( \3484 , \3481 , \3407 );
nand \U$3108 ( \3485 , \3483 , \3484 );
xor \U$3109 ( \3486 , \3437 , \3452 );
not \U$3110 ( \3487 , \1910 );
not \U$3111 ( \3488 , \2599 );
or \U$3112 ( \3489 , \3487 , \3488 );
and \U$3113 ( \3490 , RIae793b8_143, \2031 );
not \U$3114 ( \3491 , RIae793b8_143);
and \U$3115 ( \3492 , \3491 , \2027 );
or \U$3116 ( \3493 , \3490 , \3492 );
not \U$3117 ( \3494 , \1864 );
or \U$3118 ( \3495 , \3493 , \3494 );
nand \U$3119 ( \3496 , \3489 , \3495 );
xor \U$3120 ( \3497 , RIae79250_140, \1880 );
or \U$3121 ( \3498 , \3497 , \1502 );
not \U$3122 ( \3499 , \2650 );
or \U$3123 ( \3500 , \2617 , \3499 );
nand \U$3124 ( \3501 , \3498 , \3500 );
xor \U$3125 ( \3502 , \3496 , \3501 );
not \U$3126 ( \3503 , RIae79ac0_158);
not \U$3127 ( \3504 , \1024 );
or \U$3128 ( \3505 , \3503 , \3504 );
or \U$3129 ( \3506 , \857 , RIae79ac0_158);
nand \U$3130 ( \3507 , \3505 , \3506 );
not \U$3131 ( \3508 , \3507 );
or \U$3132 ( \3509 , \3508 , \3016 );
not \U$3133 ( \3510 , \2272 );
or \U$3134 ( \3511 , \3013 , \3510 );
nand \U$3135 ( \3512 , \3509 , \3511 );
xor \U$3136 ( \3513 , \3502 , \3512 );
xor \U$3137 ( \3514 , \3486 , \3513 );
not \U$3138 ( \3515 , \2096 );
not \U$3139 ( \3516 , \3418 );
or \U$3140 ( \3517 , \3515 , \3516 );
nand \U$3141 ( \3518 , \2095 , \893 );
nand \U$3142 ( \3519 , \3517 , \3518 );
not \U$3143 ( \3520 , \1036 );
not \U$3144 ( \3521 , \3520 );
not \U$3145 ( \3522 , \2579 );
and \U$3146 ( \3523 , \3521 , \3522 );
not \U$3147 ( \3524 , \1808 );
buf \U$3148 ( \3525 , \3524 );
and \U$3149 ( \3526 , RIae78bc0_126, \3525 );
not \U$3150 ( \3527 , RIae78bc0_126);
not \U$3151 ( \3528 , \1808 );
not \U$3152 ( \3529 , \3528 );
buf \U$3153 ( \3530 , \3529 );
and \U$3154 ( \3531 , \3527 , \3530 );
or \U$3155 ( \3532 , \3526 , \3531 );
and \U$3156 ( \3533 , \3532 , \929 );
nor \U$3157 ( \3534 , \3523 , \3533 );
xor \U$3158 ( \3535 , \3519 , \3534 );
not \U$3159 ( \3536 , \2011 );
not \U$3160 ( \3537 , RIae79610_148);
not \U$3161 ( \3538 , \1185 );
not \U$3162 ( \3539 , \3538 );
not \U$3163 ( \3540 , \3539 );
or \U$3164 ( \3541 , \3537 , \3540 );
or \U$3165 ( \3542 , \1186 , RIae79610_148);
nand \U$3166 ( \3543 , \3541 , \3542 );
not \U$3167 ( \3544 , \3543 );
or \U$3168 ( \3545 , \3536 , \3544 );
nand \U$3169 ( \3546 , \2106 , \2063 );
nand \U$3170 ( \3547 , \3545 , \3546 );
xnor \U$3171 ( \3548 , \3535 , \3547 );
xor \U$3172 ( \3549 , \3514 , \3548 );
not \U$3173 ( \3550 , \3549 );
not \U$3174 ( \3551 , \2533 );
not \U$3175 ( \3552 , \2586 );
or \U$3176 ( \3553 , \3551 , \3552 );
not \U$3177 ( \3554 , \2583 );
not \U$3178 ( \3555 , \2532 );
or \U$3179 ( \3556 , \3554 , \3555 );
nand \U$3180 ( \3557 , \3556 , \2621 );
nand \U$3181 ( \3558 , \3553 , \3557 );
xor \U$3182 ( \3559 , \2111 , \2242 );
and \U$3183 ( \3560 , \3559 , \2347 );
and \U$3184 ( \3561 , \2111 , \2242 );
or \U$3185 ( \3562 , \3560 , \3561 );
xor \U$3186 ( \3563 , \3558 , \3562 );
not \U$3187 ( \3564 , \3563 );
or \U$3188 ( \3565 , \3550 , \3564 );
nand \U$3189 ( \3566 , \3562 , \3558 );
nand \U$3190 ( \3567 , \3565 , \3566 );
not \U$3191 ( \3568 , \3567 );
xor \U$3192 ( \3569 , \3485 , \3568 );
xor \U$3193 ( \3570 , \3486 , \3513 );
and \U$3194 ( \3571 , \3570 , \3548 );
and \U$3195 ( \3572 , \3486 , \3513 );
or \U$3196 ( \3573 , \3571 , \3572 );
not \U$3197 ( \3574 , \3124 );
not \U$3198 ( \3575 , \3091 );
or \U$3199 ( \3576 , \3574 , \3575 );
not \U$3200 ( \3577 , \3036 );
nand \U$3201 ( \3578 , \3577 , \3086 );
nand \U$3202 ( \3579 , \3576 , \3578 );
xor \U$3203 ( \3580 , \3573 , \3579 );
not \U$3204 ( \3581 , \3080 );
not \U$3205 ( \3582 , \3065 );
or \U$3206 ( \3583 , \3581 , \3582 );
nand \U$3207 ( \3584 , \3061 , \3047 );
nand \U$3208 ( \3585 , \3583 , \3584 );
xor \U$3209 ( \3586 , \3496 , \3501 );
and \U$3210 ( \3587 , \3586 , \3512 );
and \U$3211 ( \3588 , \3496 , \3501 );
or \U$3212 ( \3589 , \3587 , \3588 );
xor \U$3213 ( \3590 , \3585 , \3589 );
not \U$3214 ( \3591 , \3116 );
xor \U$3215 ( \3592 , \3123 , \3104 );
not \U$3216 ( \3593 , \3592 );
or \U$3217 ( \3594 , \3591 , \3593 );
nand \U$3218 ( \3595 , \3123 , \3104 );
nand \U$3219 ( \3596 , \3594 , \3595 );
xnor \U$3220 ( \3597 , \3590 , \3596 );
and \U$3221 ( \3598 , \3580 , \3597 );
not \U$3222 ( \3599 , \3580 );
xor \U$3223 ( \3600 , \3590 , \3596 );
and \U$3224 ( \3601 , \3599 , \3600 );
nor \U$3225 ( \3602 , \3598 , \3601 );
xor \U$3226 ( \3603 , \3569 , \3602 );
not \U$3227 ( \3604 , \3603 );
not \U$3228 ( \3605 , \3604 );
xor \U$3229 ( \3606 , \1849 , \1938 );
and \U$3230 ( \3607 , \3606 , \2071 );
and \U$3231 ( \3608 , \1849 , \1938 );
or \U$3232 ( \3609 , \3607 , \3608 );
xor \U$3233 ( \3610 , \3393 , \3397 );
xor \U$3234 ( \3611 , \3610 , \3404 );
xor \U$3235 ( \3612 , \3609 , \3611 );
xor \U$3236 ( \3613 , \3426 , \3475 );
xor \U$3237 ( \3614 , \3613 , \3465 );
xnor \U$3238 ( \3615 , \3612 , \3614 );
not \U$3239 ( \3616 , \3615 );
xnor \U$3240 ( \3617 , \3563 , \3549 );
not \U$3241 ( \3618 , \3617 );
or \U$3242 ( \3619 , \3616 , \3618 );
not \U$3243 ( \3620 , \2717 );
not \U$3244 ( \3621 , \2739 );
or \U$3245 ( \3622 , \3620 , \3621 );
not \U$3246 ( \3623 , \2744 );
nand \U$3247 ( \3624 , \3623 , \2622 );
nand \U$3248 ( \3625 , \3622 , \3624 );
nand \U$3249 ( \3626 , \3619 , \3625 );
or \U$3250 ( \3627 , \3617 , \3615 );
nand \U$3251 ( \3628 , \3626 , \3627 );
not \U$3252 ( \3629 , \3628 );
not \U$3253 ( \3630 , \3134 );
not \U$3254 ( \3631 , \2897 );
or \U$3255 ( \3632 , \3630 , \3631 );
nand \U$3256 ( \3633 , \3130 , \3031 );
nand \U$3257 ( \3634 , \3632 , \3633 );
not \U$3258 ( \3635 , \3634 );
not \U$3259 ( \3636 , \3611 );
and \U$3260 ( \3637 , \3614 , \3609 );
not \U$3261 ( \3638 , \3614 );
not \U$3262 ( \3639 , \3609 );
and \U$3263 ( \3640 , \3638 , \3639 );
nor \U$3264 ( \3641 , \3637 , \3640 );
not \U$3265 ( \3642 , \3641 );
or \U$3266 ( \3643 , \3636 , \3642 );
nand \U$3267 ( \3644 , \3614 , \3609 );
nand \U$3268 ( \3645 , \3643 , \3644 );
not \U$3269 ( \3646 , \3645 );
xor \U$3270 ( \3647 , \3547 , \3519 );
not \U$3271 ( \3648 , \3534 );
and \U$3272 ( \3649 , \3647 , \3648 );
and \U$3273 ( \3650 , \3547 , \3519 );
or \U$3274 ( \3651 , \3649 , \3650 );
not \U$3275 ( \3652 , \3651 );
not \U$3276 ( \3653 , RIae79700_150);
not \U$3277 ( \3654 , RIae79778_151);
or \U$3278 ( \3655 , \3653 , \3654 );
nand \U$3279 ( \3656 , \3655 , RIae797f0_152);
not \U$3280 ( \3657 , \2189 );
not \U$3281 ( \3658 , \3447 );
or \U$3282 ( \3659 , \3657 , \3658 );
not \U$3283 ( \3660 , \2923 );
not \U$3284 ( \3661 , \2183 );
not \U$3285 ( \3662 , \1289 );
or \U$3286 ( \3663 , \3661 , \3662 );
or \U$3287 ( \3664 , \1291 , \2183 );
nand \U$3288 ( \3665 , \3663 , \3664 );
nand \U$3289 ( \3666 , \3660 , \3665 );
nand \U$3290 ( \3667 , \3659 , \3666 );
xor \U$3291 ( \3668 , \3656 , \3667 );
not \U$3292 ( \3669 , \2322 );
not \U$3293 ( \3670 , \2334 );
not \U$3294 ( \3671 , \1196 );
or \U$3295 ( \3672 , \3670 , \3671 );
or \U$3296 ( \3673 , \1196 , \2334 );
nand \U$3297 ( \3674 , \3672 , \3673 );
not \U$3298 ( \3675 , \3674 );
or \U$3299 ( \3676 , \3669 , \3675 );
nand \U$3300 ( \3677 , \3433 , \2341 );
nand \U$3301 ( \3678 , \3676 , \3677 );
xnor \U$3302 ( \3679 , \3668 , \3678 );
not \U$3303 ( \3680 , \3679 );
or \U$3304 ( \3681 , \3652 , \3680 );
or \U$3305 ( \3682 , \3651 , \3679 );
nand \U$3306 ( \3683 , \3681 , \3682 );
not \U$3307 ( \3684 , \3683 );
nand \U$3308 ( \3685 , \2093 , RIae78b48_125);
not \U$3309 ( \3686 , \3685 );
not \U$3310 ( \3687 , \1864 );
not \U$3311 ( \3688 , \2848 );
not \U$3312 ( \3689 , \3688 );
and \U$3313 ( \3690 , RIae793b8_143, \3689 );
not \U$3314 ( \3691 , RIae793b8_143);
and \U$3315 ( \3692 , \3691 , \2849 );
nor \U$3316 ( \3693 , \3690 , \3692 );
not \U$3317 ( \3694 , \3693 );
or \U$3318 ( \3695 , \3687 , \3694 );
not \U$3319 ( \3696 , \3493 );
nand \U$3320 ( \3697 , \3696 , \1910 );
nand \U$3321 ( \3698 , \3695 , \3697 );
xor \U$3322 ( \3699 , \3686 , \3698 );
and \U$3323 ( \3700 , \3141 , \1503 );
not \U$3324 ( \3701 , \3141 );
and \U$3325 ( \3702 , \3701 , RIae79250_140);
nor \U$3326 ( \3703 , \3700 , \3702 );
not \U$3327 ( \3704 , \3703 );
nor \U$3328 ( \3705 , \3704 , \1502 );
nor \U$3329 ( \3706 , \3497 , \1498 );
or \U$3330 ( \3707 , \3705 , \3706 );
xnor \U$3331 ( \3708 , \3699 , \3707 );
not \U$3332 ( \3709 , \3708 );
and \U$3333 ( \3710 , \3684 , \3709 );
and \U$3334 ( \3711 , \3683 , \3708 );
nor \U$3335 ( \3712 , \3710 , \3711 );
not \U$3336 ( \3713 , \3712 );
not \U$3337 ( \3714 , \2063 );
not \U$3338 ( \3715 , \3543 );
or \U$3339 ( \3716 , \3714 , \3715 );
not \U$3340 ( \3717 , \2056 );
not \U$3341 ( \3718 , \1125 );
not \U$3342 ( \3719 , \3718 );
or \U$3343 ( \3720 , \3717 , \3719 );
not \U$3344 ( \3721 , \976 );
buf \U$3345 ( \3722 , \3721 );
nand \U$3346 ( \3723 , \3722 , RIae79610_148);
nand \U$3347 ( \3724 , \3720 , \3723 );
nand \U$3348 ( \3725 , \3724 , \2011 );
nand \U$3349 ( \3726 , \3716 , \3725 );
not \U$3350 ( \3727 , \3726 );
not \U$3351 ( \3728 , \953 );
not \U$3352 ( \3729 , \3532 );
or \U$3353 ( \3730 , \3728 , \3729 );
and \U$3354 ( \3731 , \1755 , RIae78bc0_126);
not \U$3355 ( \3732 , \1755 );
and \U$3356 ( \3733 , \3732 , \1286 );
nor \U$3357 ( \3734 , \3731 , \3733 );
nand \U$3358 ( \3735 , \3734 , \1027 );
nand \U$3359 ( \3736 , \3730 , \3735 );
not \U$3360 ( \3737 , \3736 );
not \U$3361 ( \3738 , \3101 );
not \U$3362 ( \3739 , \1413 );
and \U$3363 ( \3740 , \3738 , \3739 );
and \U$3364 ( \3741 , RIae78e90_132, \2287 );
not \U$3365 ( \3742 , RIae78e90_132);
not \U$3366 ( \3743 , \2284 );
and \U$3367 ( \3744 , \2283 , \3743 );
not \U$3368 ( \3745 , \2283 );
and \U$3369 ( \3746 , \3745 , \2284 );
nor \U$3370 ( \3747 , \3744 , \3746 );
buf \U$3371 ( \3748 , \3747 );
and \U$3372 ( \3749 , \3742 , \3748 );
or \U$3373 ( \3750 , \3741 , \3749 );
and \U$3374 ( \3751 , \3750 , \1321 );
nor \U$3375 ( \3752 , \3740 , \3751 );
not \U$3376 ( \3753 , \3752 );
and \U$3377 ( \3754 , \3737 , \3753 );
and \U$3378 ( \3755 , \3736 , \3752 );
nor \U$3379 ( \3756 , \3754 , \3755 );
not \U$3380 ( \3757 , \3756 );
or \U$3381 ( \3758 , \3727 , \3757 );
or \U$3382 ( \3759 , \3756 , \3726 );
nand \U$3383 ( \3760 , \3758 , \3759 );
not \U$3384 ( \3761 , \3760 );
not \U$3385 ( \3762 , \1062 );
not \U$3386 ( \3763 , \3076 );
or \U$3387 ( \3764 , \3762 , \3763 );
not \U$3388 ( \3765 , \2993 );
xor \U$3389 ( \3766 , RIae79070_136, \3765 );
nand \U$3390 ( \3767 , \3766 , \1049 );
nand \U$3391 ( \3768 , \3764 , \3767 );
not \U$3392 ( \3769 , \2272 );
not \U$3393 ( \3770 , \3507 );
or \U$3394 ( \3771 , \3769 , \3770 );
not \U$3395 ( \3772 , RIae79ac0_158);
not \U$3396 ( \3773 , \940 );
or \U$3397 ( \3774 , \3772 , \3773 );
not \U$3398 ( \3775 , \3236 );
or \U$3399 ( \3776 , \3775 , RIae79ac0_158);
nand \U$3400 ( \3777 , \3774 , \3776 );
nand \U$3401 ( \3778 , \3777 , \2252 );
nand \U$3402 ( \3779 , \3771 , \3778 );
xor \U$3403 ( \3780 , \3768 , \3779 );
not \U$3404 ( \3781 , \3780 );
not \U$3405 ( \3782 , \1430 );
not \U$3406 ( \3783 , \3057 );
or \U$3407 ( \3784 , \3782 , \3783 );
not \U$3408 ( \3785 , \3294 );
and \U$3409 ( \3786 , RIae79160_138, \3785 );
not \U$3410 ( \3787 , RIae79160_138);
and \U$3411 ( \3788 , \3787 , \1899 );
nor \U$3412 ( \3789 , \3786 , \3788 );
not \U$3413 ( \3790 , \3789 );
nand \U$3414 ( \3791 , \3790 , \1013 );
nand \U$3415 ( \3792 , \3784 , \3791 );
not \U$3416 ( \3793 , \3792 );
not \U$3417 ( \3794 , \3793 );
and \U$3418 ( \3795 , \3781 , \3794 );
and \U$3419 ( \3796 , \3780 , \3793 );
nor \U$3420 ( \3797 , \3795 , \3796 );
not \U$3421 ( \3798 , \839 );
and \U$3422 ( \3799 , \2956 , \1132 );
not \U$3423 ( \3800 , \2956 );
and \U$3424 ( \3801 , \3800 , RIae78f80_134);
nor \U$3425 ( \3802 , \3799 , \3801 );
not \U$3426 ( \3803 , \3802 );
or \U$3427 ( \3804 , \3798 , \3803 );
nand \U$3428 ( \3805 , \3110 , \797 );
nand \U$3429 ( \3806 , \3804 , \3805 );
not \U$3430 ( \3807 , \1933 );
not \U$3431 ( \3808 , \3043 );
or \U$3432 ( \3809 , \3807 , \3808 );
not \U$3433 ( \3810 , RIae794a8_145);
not \U$3434 ( \3811 , \3810 );
not \U$3435 ( \3812 , \3283 );
or \U$3436 ( \3813 , \3811 , \3812 );
not \U$3437 ( \3814 , \781 );
nand \U$3438 ( \3815 , \3814 , RIae794a8_145);
nand \U$3439 ( \3816 , \3813 , \3815 );
nand \U$3440 ( \3817 , \3816 , \1919 );
nand \U$3441 ( \3818 , \3809 , \3817 );
xor \U$3442 ( \3819 , \3806 , \3818 );
not \U$3443 ( \3820 , \2966 );
not \U$3444 ( \3821 , \3119 );
or \U$3445 ( \3822 , \3820 , \3821 );
and \U$3446 ( \3823 , \2179 , \3147 );
not \U$3447 ( \3824 , \2179 );
and \U$3448 ( \3825 , \3824 , RIae79688_149);
nor \U$3449 ( \3826 , \3823 , \3825 );
buf \U$3450 ( \3827 , \1821 );
nand \U$3451 ( \3828 , \3826 , \3827 );
nand \U$3452 ( \3829 , \3822 , \3828 );
xor \U$3453 ( \3830 , \3819 , \3829 );
not \U$3454 ( \3831 , \3830 );
and \U$3455 ( \3832 , \3797 , \3831 );
not \U$3456 ( \3833 , \3797 );
and \U$3457 ( \3834 , \3833 , \3830 );
nor \U$3458 ( \3835 , \3832 , \3834 );
not \U$3459 ( \3836 , \3835 );
not \U$3460 ( \3837 , \3836 );
or \U$3461 ( \3838 , \3761 , \3837 );
not \U$3462 ( \3839 , \3760 );
nand \U$3463 ( \3840 , \3839 , \3835 );
nand \U$3464 ( \3841 , \3838 , \3840 );
not \U$3465 ( \3842 , \3841 );
or \U$3466 ( \3843 , \3713 , \3842 );
or \U$3467 ( \3844 , \3841 , \3712 );
nand \U$3468 ( \3845 , \3843 , \3844 );
not \U$3469 ( \3846 , \3845 );
not \U$3470 ( \3847 , \3846 );
or \U$3471 ( \3848 , \3646 , \3847 );
not \U$3472 ( \3849 , \3645 );
nand \U$3473 ( \3850 , \3845 , \3849 );
nand \U$3474 ( \3851 , \3848 , \3850 );
not \U$3475 ( \3852 , \3851 );
not \U$3476 ( \3853 , \3852 );
or \U$3477 ( \3854 , \3635 , \3853 );
not \U$3478 ( \3855 , \3634 );
nand \U$3479 ( \3856 , \3855 , \3851 );
nand \U$3480 ( \3857 , \3854 , \3856 );
not \U$3481 ( \3858 , \3857 );
not \U$3482 ( \3859 , \3858 );
or \U$3483 ( \3860 , \3629 , \3859 );
not \U$3484 ( \3861 , \3628 );
nand \U$3485 ( \3862 , \3861 , \3857 );
nand \U$3486 ( \3863 , \3860 , \3862 );
not \U$3487 ( \3864 , \3863 );
not \U$3488 ( \3865 , \3864 );
or \U$3489 ( \3866 , \3605 , \3865 );
nand \U$3490 ( \3867 , \3863 , \3603 );
nand \U$3491 ( \3868 , \3866 , \3867 );
not \U$3492 ( \3869 , \3868 );
or \U$3493 ( \3870 , \3389 , \3869 );
or \U$3494 ( \3871 , \3388 , \3868 );
nand \U$3495 ( \3872 , \3870 , \3871 );
xor \U$3496 ( \3873 , \2892 , \3382 );
xor \U$3497 ( \3874 , \3615 , \3617 );
xor \U$3498 ( \3875 , \3874 , \3625 );
or \U$3499 ( \3876 , \3873 , \3875 );
xor \U$3500 ( \3877 , \2887 , \2885 );
xnor \U$3501 ( \3878 , \3877 , \2818 );
not \U$3502 ( \3879 , \3878 );
xor \U$3503 ( \3880 , \3297 , \3277 );
xnor \U$3504 ( \3881 , \3880 , \3290 );
not \U$3505 ( \3882 , \3881 );
not \U$3506 ( \3883 , \3882 );
not \U$3507 ( \3884 , \2765 );
not \U$3508 ( \3885 , \2794 );
or \U$3509 ( \3886 , \3884 , \3885 );
or \U$3510 ( \3887 , \2794 , \2765 );
nand \U$3511 ( \3888 , \3886 , \3887 );
not \U$3512 ( \3889 , \3226 );
not \U$3513 ( \3890 , \3151 );
not \U$3514 ( \3891 , \3890 );
and \U$3515 ( \3892 , \3889 , \3891 );
and \U$3516 ( \3893 , \3226 , \3890 );
nor \U$3517 ( \3894 , \3892 , \3893 );
and \U$3518 ( \3895 , \3888 , \3894 );
not \U$3519 ( \3896 , \3888 );
not \U$3520 ( \3897 , \3894 );
and \U$3521 ( \3898 , \3896 , \3897 );
or \U$3522 ( \3899 , \3895 , \3898 );
not \U$3523 ( \3900 , \3899 );
or \U$3524 ( \3901 , \3883 , \3900 );
nand \U$3525 ( \3902 , \3888 , \3897 );
nand \U$3526 ( \3903 , \3901 , \3902 );
nand \U$3527 ( \3904 , \2878 , \2870 );
not \U$3528 ( \3905 , \2873 );
and \U$3529 ( \3906 , \3904 , \3905 );
not \U$3530 ( \3907 , \3904 );
and \U$3531 ( \3908 , \3907 , \2873 );
nor \U$3532 ( \3909 , \3906 , \3908 );
nor \U$3533 ( \3910 , \3903 , \3909 );
not \U$3534 ( \3911 , \3910 );
nand \U$3535 ( \3912 , \3903 , \3909 );
xnor \U$3536 ( \3913 , \2813 , \2751 );
nand \U$3537 ( \3914 , \3912 , \3913 );
nand \U$3538 ( \3915 , \3911 , \3914 );
not \U$3539 ( \3916 , \3915 );
not \U$3540 ( \3917 , \3916 );
or \U$3541 ( \3918 , \3879 , \3917 );
not \U$3542 ( \3919 , \3915 );
not \U$3543 ( \3920 , \3878 );
not \U$3544 ( \3921 , \3920 );
or \U$3545 ( \3922 , \3919 , \3921 );
xor \U$3546 ( \3923 , \3308 , \3309 );
nand \U$3547 ( \3924 , \3922 , \3923 );
nand \U$3548 ( \3925 , \3918 , \3924 );
not \U$3549 ( \3926 , \3925 );
not \U$3550 ( \3927 , \3373 );
not \U$3551 ( \3928 , \3312 );
or \U$3552 ( \3929 , \3927 , \3928 );
or \U$3553 ( \3930 , \3373 , \3312 );
nand \U$3554 ( \3931 , \3929 , \3930 );
not \U$3555 ( \3932 , \3364 );
not \U$3556 ( \3933 , \3362 );
not \U$3557 ( \3934 , \3361 );
or \U$3558 ( \3935 , \3933 , \3934 );
or \U$3559 ( \3936 , \3362 , \3361 );
nand \U$3560 ( \3937 , \3935 , \3936 );
not \U$3561 ( \3938 , \3937 );
or \U$3562 ( \3939 , \3932 , \3938 );
or \U$3563 ( \3940 , \3937 , \3364 );
nand \U$3564 ( \3941 , \3939 , \3940 );
not \U$3565 ( \3942 , \3941 );
not \U$3566 ( \3943 , \3942 );
xor \U$3567 ( \3944 , \2421 , \2798 );
xnor \U$3568 ( \3945 , \3944 , \2452 );
and \U$3569 ( \3946 , \3945 , \3358 );
not \U$3570 ( \3947 , \3945 );
not \U$3571 ( \3948 , \3358 );
and \U$3572 ( \3949 , \3947 , \3948 );
nor \U$3573 ( \3950 , \3946 , \3949 );
not \U$3574 ( \3951 , \3950 );
xor \U$3575 ( \3952 , \3239 , \3251 );
xor \U$3576 ( \3953 , \3952 , \3262 );
not \U$3577 ( \3954 , \3355 );
not \U$3578 ( \3955 , \3343 );
or \U$3579 ( \3956 , \3954 , \3955 );
not \U$3580 ( \3957 , \3342 );
or \U$3581 ( \3958 , \3355 , \3957 );
nand \U$3582 ( \3959 , \3956 , \3958 );
and \U$3583 ( \3960 , \3959 , \3330 );
not \U$3584 ( \3961 , \3959 );
and \U$3585 ( \3962 , \3961 , \3331 );
nor \U$3586 ( \3963 , \3960 , \3962 );
nand \U$3587 ( \3964 , \3953 , \3963 );
or \U$3588 ( \3965 , \3963 , \3953 );
xor \U$3589 ( \3966 , \2866 , \2840 );
xnor \U$3590 ( \3967 , \3966 , \2854 );
nand \U$3591 ( \3968 , \3965 , \3967 );
nand \U$3592 ( \3969 , \3964 , \3968 );
not \U$3593 ( \3970 , \3969 );
or \U$3594 ( \3971 , \3951 , \3970 );
or \U$3595 ( \3972 , \3969 , \3950 );
nand \U$3596 ( \3973 , \3971 , \3972 );
not \U$3597 ( \3974 , \3973 );
xor \U$3598 ( \3975 , \3231 , \3265 );
xor \U$3599 ( \3976 , \3975 , \3302 );
not \U$3600 ( \3977 , \3976 );
or \U$3601 ( \3978 , \3974 , \3977 );
not \U$3602 ( \3979 , \3950 );
nand \U$3603 ( \3980 , \3979 , \3969 );
nand \U$3604 ( \3981 , \3978 , \3980 );
not \U$3605 ( \3982 , \3981 );
or \U$3606 ( \3983 , \3943 , \3982 );
not \U$3607 ( \3984 , \3941 );
not \U$3608 ( \3985 , \3981 );
not \U$3609 ( \3986 , \3985 );
or \U$3610 ( \3987 , \3984 , \3986 );
not \U$3611 ( \3988 , \1501 );
not \U$3612 ( \3989 , \3340 );
or \U$3613 ( \3990 , \3988 , \3989 );
not \U$3614 ( \3991 , \2652 );
not \U$3615 ( \3992 , \2310 );
or \U$3616 ( \3993 , \3991 , \3992 );
nand \U$3617 ( \3994 , \2305 , RIae79250_140);
nand \U$3618 ( \3995 , \3993 , \3994 );
nand \U$3619 ( \3996 , \3995 , \2650 );
nand \U$3620 ( \3997 , \3990 , \3996 );
not \U$3621 ( \3998 , \2433 );
not \U$3622 ( \3999 , \1141 );
and \U$3623 ( \4000 , RIae79778_151, \3999 );
not \U$3624 ( \4001 , RIae79778_151);
and \U$3625 ( \4002 , \4001 , \2640 );
or \U$3626 ( \4003 , \4000 , \4002 );
not \U$3627 ( \4004 , \4003 );
or \U$3628 ( \4005 , \3998 , \4004 );
nand \U$3629 ( \4006 , \3288 , \2450 );
nand \U$3630 ( \4007 , \4005 , \4006 );
xor \U$3631 ( \4008 , \3997 , \4007 );
not \U$3632 ( \4009 , \1933 );
and \U$3633 ( \4010 , \3039 , \1119 );
not \U$3634 ( \4011 , \3039 );
and \U$3635 ( \4012 , \4011 , \1120 );
nor \U$3636 ( \4013 , \4010 , \4012 );
not \U$3637 ( \4014 , \4013 );
or \U$3638 ( \4015 , \4009 , \4014 );
nand \U$3639 ( \4016 , \3260 , \2467 );
nand \U$3640 ( \4017 , \4015 , \4016 );
and \U$3641 ( \4018 , \4008 , \4017 );
and \U$3642 ( \4019 , \3997 , \4007 );
or \U$3643 ( \4020 , \4018 , \4019 );
and \U$3644 ( \4021 , RIae79160_138, \3099 );
not \U$3645 ( \4022 , RIae79160_138);
not \U$3646 ( \4023 , \3092 );
not \U$3647 ( \4024 , \4023 );
and \U$3648 ( \4025 , \4022 , \4024 );
nor \U$3649 ( \4026 , \4021 , \4025 );
not \U$3650 ( \4027 , \4026 );
not \U$3651 ( \4028 , \2157 );
or \U$3652 ( \4029 , \4027 , \4028 );
nand \U$3653 ( \4030 , \2838 , \1013 );
nand \U$3654 ( \4031 , \4029 , \4030 );
not \U$3655 ( \4032 , \4031 );
not \U$3656 ( \4033 , \2276 );
and \U$3657 ( \4034 , RIae79070_136, \1809 );
not \U$3658 ( \4035 , RIae79070_136);
not \U$3659 ( \4036 , \2696 );
and \U$3660 ( \4037 , \4035 , \4036 );
or \U$3661 ( \4038 , \4034 , \4037 );
not \U$3662 ( \4039 , \4038 );
or \U$3663 ( \4040 , \4033 , \4039 );
nand \U$3664 ( \4041 , \2864 , \1049 );
nand \U$3665 ( \4042 , \4040 , \4041 );
not \U$3666 ( \4043 , \4042 );
nand \U$3667 ( \4044 , \4032 , \4043 );
not \U$3668 ( \4045 , \4044 );
not \U$3669 ( \4046 , \2189 );
and \U$3670 ( \4047 , \1826 , RIae79520_146);
not \U$3671 ( \4048 , \1826 );
and \U$3672 ( \4049 , \4048 , \2183 );
nor \U$3673 ( \4050 , \4047 , \4049 );
not \U$3674 ( \4051 , \4050 );
or \U$3675 ( \4052 , \4046 , \4051 );
nand \U$3676 ( \4053 , \3353 , \2163 );
nand \U$3677 ( \4054 , \4052 , \4053 );
not \U$3678 ( \4055 , \4054 );
or \U$3679 ( \4056 , \4045 , \4055 );
nand \U$3680 ( \4057 , \4042 , \4031 );
nand \U$3681 ( \4058 , \4056 , \4057 );
xor \U$3682 ( \4059 , \4020 , \4058 );
not \U$3683 ( \4060 , \2063 );
not \U$3684 ( \4061 , RIae79610_148);
not \U$3685 ( \4062 , \2212 );
or \U$3686 ( \4063 , \4061 , \4062 );
not \U$3687 ( \4064 , \2207 );
not \U$3688 ( \4065 , \4064 );
nand \U$3689 ( \4066 , \4065 , \2056 );
nand \U$3690 ( \4067 , \4063 , \4066 );
not \U$3691 ( \4068 , \4067 );
or \U$3692 ( \4069 , \4060 , \4068 );
nand \U$3693 ( \4070 , \3295 , \2011 );
nand \U$3694 ( \4071 , \4069 , \4070 );
not \U$3695 ( \4072 , \2341 );
xor \U$3696 ( \4073 , \1023 , RIae798e0_154);
not \U$3697 ( \4074 , \4073 );
or \U$3698 ( \4075 , \4072 , \4074 );
nand \U$3699 ( \4076 , \3237 , \2322 );
nand \U$3700 ( \4077 , \4075 , \4076 );
xor \U$3701 ( \4078 , \4071 , \4077 );
not \U$3702 ( \4079 , \1910 );
not \U$3703 ( \4080 , \2140 );
buf \U$3704 ( \4081 , \4080 );
and \U$3705 ( \4082 , RIae793b8_143, \4081 );
not \U$3706 ( \4083 , RIae793b8_143);
and \U$3707 ( \4084 , \4083 , \2137 );
nor \U$3708 ( \4085 , \4082 , \4084 );
not \U$3709 ( \4086 , \4085 );
or \U$3710 ( \4087 , \4079 , \4086 );
nand \U$3711 ( \4088 , \3249 , \1864 );
nand \U$3712 ( \4089 , \4087 , \4088 );
and \U$3713 ( \4090 , \4078 , \4089 );
and \U$3714 ( \4091 , \4071 , \4077 );
or \U$3715 ( \4092 , \4090 , \4091 );
and \U$3716 ( \4093 , \4059 , \4092 );
and \U$3717 ( \4094 , \4020 , \4058 );
or \U$3718 ( \4095 , \4093 , \4094 );
not \U$3719 ( \4096 , \4095 );
xor \U$3720 ( \4097 , \2931 , \2911 );
xor \U$3721 ( \4098 , \4097 , \2935 );
not \U$3722 ( \4099 , \952 );
not \U$3723 ( \4100 , \2385 );
and \U$3724 ( \4101 , RIae78bc0_126, \4100 );
not \U$3725 ( \4102 , RIae78bc0_126);
not \U$3726 ( \4103 , \1860 );
and \U$3727 ( \4104 , \4102 , \4103 );
or \U$3728 ( \4105 , \4101 , \4104 );
not \U$3729 ( \4106 , \4105 );
or \U$3730 ( \4107 , \4099 , \4106 );
nand \U$3731 ( \4108 , \3219 , \1027 );
nand \U$3732 ( \4109 , \4107 , \4108 );
not \U$3733 ( \4110 , \4109 );
not \U$3734 ( \4111 , \1087 );
buf \U$3735 ( \4112 , \2355 );
buf \U$3736 ( \4113 , \4112 );
and \U$3737 ( \4114 , \4113 , \1066 );
not \U$3738 ( \4115 , \4113 );
and \U$3739 ( \4116 , \4115 , RIae78e90_132);
nor \U$3740 ( \4117 , \4114 , \4116 );
not \U$3741 ( \4118 , \4117 );
or \U$3742 ( \4119 , \4111 , \4118 );
nand \U$3743 ( \4120 , \2788 , \1320 );
nand \U$3744 ( \4121 , \4119 , \4120 );
not \U$3745 ( \4122 , \4121 );
or \U$3746 ( \4123 , \4110 , \4122 );
or \U$3747 ( \4124 , \4121 , \4109 );
not \U$3748 ( \4125 , \3015 );
not \U$3749 ( \4126 , \2852 );
or \U$3750 ( \4127 , \4125 , \4126 );
and \U$3751 ( \4128 , \2031 , RIae79ac0_158);
not \U$3752 ( \4129 , \2031 );
and \U$3753 ( \4130 , \4129 , \2268 );
nor \U$3754 ( \4131 , \4128 , \4130 );
nand \U$3755 ( \4132 , \4131 , \2272 );
nand \U$3756 ( \4133 , \4127 , \4132 );
nand \U$3757 ( \4134 , \4124 , \4133 );
nand \U$3758 ( \4135 , \4123 , \4134 );
not \U$3759 ( \4136 , \4135 );
not \U$3760 ( \4137 , \1129 );
xor \U$3761 ( \4138 , RIae78b48_125, \3208 );
not \U$3762 ( \4139 , \4138 );
or \U$3763 ( \4140 , \4137 , \4139 );
or \U$3764 ( \4141 , \3275 , \1959 );
nand \U$3765 ( \4142 , \4140 , \4141 );
not \U$3766 ( \4143 , \4142 );
nand \U$3767 ( \4144 , RIae79d90_164, RIae79e08_165);
not \U$3768 ( \4145 , \4144 );
nor \U$3769 ( \4146 , RIae79d90_164, RIae79e08_165);
nor \U$3770 ( \4147 , \4145 , \4146 );
not \U$3771 ( \4148 , \4147 );
and \U$3772 ( \4149 , RIae79ca0_162, RIae79e08_165);
not \U$3773 ( \4150 , RIae79ca0_162);
not \U$3774 ( \4151 , RIae79e08_165);
and \U$3775 ( \4152 , \4150 , \4151 );
nor \U$3776 ( \4153 , \4149 , \4152 );
and \U$3777 ( \4154 , \4148 , \4153 );
buf \U$3778 ( \4155 , \4147 );
or \U$3779 ( \4156 , \4154 , \4155 );
nand \U$3780 ( \4157 , \4156 , RIae79ca0_162);
not \U$3781 ( \4158 , \4157 );
not \U$3782 ( \4159 , \3156 );
not \U$3783 ( \4160 , \3198 );
or \U$3784 ( \4161 , \4159 , \4160 );
not \U$3785 ( \4162 , \602 );
nand \U$3786 ( \4163 , \4161 , \4162 );
nand \U$3787 ( \4164 , \3157 , \605 );
nor \U$3788 ( \4165 , \4163 , \4164 );
not \U$3789 ( \4166 , \4165 );
nand \U$3790 ( \4167 , \4163 , \4164 );
nand \U$3791 ( \4168 , \4166 , \4167 );
buf \U$3792 ( \4169 , \4168 );
buf \U$3793 ( \4170 , \4169 );
nand \U$3794 ( \4171 , \4170 , RIae78b48_125);
not \U$3795 ( \4172 , \4171 );
or \U$3796 ( \4173 , \4158 , \4172 );
not \U$3797 ( \4174 , \4157 );
nand \U$3798 ( \4175 , \4174 , \4170 , RIae78b48_125);
nand \U$3799 ( \4176 , \4173 , \4175 );
not \U$3800 ( \4177 , \4176 );
or \U$3801 ( \4178 , \4143 , \4177 );
nand \U$3802 ( \4179 , \4170 , \4157 , RIae78b48_125);
nand \U$3803 ( \4180 , \4178 , \4179 );
not \U$3804 ( \4181 , \2776 );
not \U$3805 ( \4182 , \2773 );
or \U$3806 ( \4183 , \4181 , \4182 );
and \U$3807 ( \4184 , RIae79c28_161, \834 );
not \U$3808 ( \4185 , RIae79c28_161);
and \U$3809 ( \4186 , \4185 , \2004 );
or \U$3810 ( \4187 , \4184 , \4186 );
nand \U$3811 ( \4188 , \4187 , \2767 );
nand \U$3812 ( \4189 , \4183 , \4188 );
not \U$3813 ( \4190 , \4189 );
not \U$3814 ( \4191 , \1821 );
not \U$3815 ( \4192 , \3149 );
or \U$3816 ( \4193 , \4191 , \4192 );
not \U$3817 ( \4194 , \1878 );
and \U$3818 ( \4195 , RIae79688_149, \4194 );
not \U$3819 ( \4196 , RIae79688_149);
buf \U$3820 ( \4197 , \1877 );
not \U$3821 ( \4198 , \4197 );
not \U$3822 ( \4199 , \4198 );
and \U$3823 ( \4200 , \4196 , \4199 );
nor \U$3824 ( \4201 , \4195 , \4200 );
nand \U$3825 ( \4202 , \4201 , \1844 );
nand \U$3826 ( \4203 , \4193 , \4202 );
not \U$3827 ( \4204 , \4203 );
or \U$3828 ( \4205 , \4190 , \4204 );
or \U$3829 ( \4206 , \4189 , \4203 );
not \U$3830 ( \4207 , \1989 );
not \U$3831 ( \4208 , RIae797f0_152);
not \U$3832 ( \4209 , \1439 );
or \U$3833 ( \4210 , \4208 , \4209 );
or \U$3834 ( \4211 , \1439 , RIae797f0_152);
nand \U$3835 ( \4212 , \4210 , \4211 );
not \U$3836 ( \4213 , \4212 );
or \U$3837 ( \4214 , \4207 , \4213 );
nand \U$3838 ( \4215 , \3328 , \2007 );
nand \U$3839 ( \4216 , \4214 , \4215 );
nand \U$3840 ( \4217 , \4206 , \4216 );
nand \U$3841 ( \4218 , \4205 , \4217 );
and \U$3842 ( \4219 , \4180 , \4218 );
not \U$3843 ( \4220 , \4180 );
not \U$3844 ( \4221 , \4218 );
and \U$3845 ( \4222 , \4220 , \4221 );
nor \U$3846 ( \4223 , \4219 , \4222 );
not \U$3847 ( \4224 , \4223 );
or \U$3848 ( \4225 , \4136 , \4224 );
not \U$3849 ( \4226 , \4221 );
nand \U$3850 ( \4227 , \4226 , \4180 );
nand \U$3851 ( \4228 , \4225 , \4227 );
and \U$3852 ( \4229 , \4098 , \4228 );
not \U$3853 ( \4230 , \4098 );
not \U$3854 ( \4231 , \4228 );
and \U$3855 ( \4232 , \4230 , \4231 );
nor \U$3856 ( \4233 , \4229 , \4232 );
not \U$3857 ( \4234 , \4233 );
or \U$3858 ( \4235 , \4096 , \4234 );
not \U$3859 ( \4236 , \4231 );
nand \U$3860 ( \4237 , \4236 , \4098 );
nand \U$3861 ( \4238 , \4235 , \4237 );
nand \U$3862 ( \4239 , \3987 , \4238 );
nand \U$3863 ( \4240 , \3983 , \4239 );
or \U$3864 ( \4241 , \3931 , \4240 );
not \U$3865 ( \4242 , \4241 );
or \U$3866 ( \4243 , \3926 , \4242 );
nand \U$3867 ( \4244 , \3931 , \4240 );
nand \U$3868 ( \4245 , \4243 , \4244 );
nand \U$3869 ( \4246 , \3876 , \4245 );
nand \U$3870 ( \4247 , \3873 , \3875 );
nand \U$3871 ( \4248 , \4246 , \4247 );
or \U$3872 ( \4249 , \3872 , \4248 );
buf \U$3873 ( \4250 , \4249 );
not \U$3874 ( \4251 , \3387 );
not \U$3875 ( \4252 , \3868 );
or \U$3876 ( \4253 , \4251 , \4252 );
nand \U$3877 ( \4254 , \3604 , \3863 );
nand \U$3878 ( \4255 , \4253 , \4254 );
not \U$3879 ( \4256 , \3857 );
not \U$3880 ( \4257 , \3628 );
or \U$3881 ( \4258 , \4256 , \4257 );
nand \U$3882 ( \4259 , \3851 , \3634 );
nand \U$3883 ( \4260 , \4258 , \4259 );
not \U$3884 ( \4261 , \4260 );
not \U$3885 ( \4262 , \4261 );
not \U$3886 ( \4263 , \3678 );
not \U$3887 ( \4264 , \3668 );
or \U$3888 ( \4265 , \4263 , \4264 );
nand \U$3889 ( \4266 , RIae79700_150, RIae79778_151);
and \U$3890 ( \4267 , \4266 , RIae797f0_152);
not \U$3891 ( \4268 , \4267 );
nand \U$3892 ( \4269 , \4268 , \3667 );
nand \U$3893 ( \4270 , \4265 , \4269 );
not \U$3894 ( \4271 , \3707 );
not \U$3895 ( \4272 , \3685 );
not \U$3896 ( \4273 , \3698 );
or \U$3897 ( \4274 , \4272 , \4273 );
or \U$3898 ( \4275 , \3698 , \3685 );
nand \U$3899 ( \4276 , \4274 , \4275 );
not \U$3900 ( \4277 , \4276 );
or \U$3901 ( \4278 , \4271 , \4277 );
nand \U$3902 ( \4279 , \3698 , \3686 );
nand \U$3903 ( \4280 , \4278 , \4279 );
xor \U$3904 ( \4281 , \4270 , \4280 );
not \U$3905 ( \4282 , \4281 );
not \U$3906 ( \4283 , \3792 );
not \U$3907 ( \4284 , \3780 );
or \U$3908 ( \4285 , \4283 , \4284 );
nand \U$3909 ( \4286 , \3779 , \3768 );
nand \U$3910 ( \4287 , \4285 , \4286 );
not \U$3911 ( \4288 , \4287 );
not \U$3912 ( \4289 , \4288 );
and \U$3913 ( \4290 , \4282 , \4289 );
and \U$3914 ( \4291 , \4281 , \4288 );
nor \U$3915 ( \4292 , \4290 , \4291 );
not \U$3916 ( \4293 , \3806 );
or \U$3917 ( \4294 , \3829 , \3818 );
not \U$3918 ( \4295 , \4294 );
or \U$3919 ( \4296 , \4293 , \4295 );
nand \U$3920 ( \4297 , \3829 , \3818 );
nand \U$3921 ( \4298 , \4296 , \4297 );
nand \U$3922 ( \4299 , \2565 , RIae78b48_125);
not \U$3923 ( \4300 , \893 );
not \U$3924 ( \4301 , \3410 );
or \U$3925 ( \4302 , \4300 , \4301 );
and \U$3926 ( \4303 , RIae78b48_125, \3525 );
not \U$3927 ( \4304 , RIae78b48_125);
not \U$3928 ( \4305 , \3525 );
and \U$3929 ( \4306 , \4304 , \4305 );
or \U$3930 ( \4307 , \4303 , \4306 );
nand \U$3931 ( \4308 , \4307 , \868 );
nand \U$3932 ( \4309 , \4302 , \4308 );
xor \U$3933 ( \4310 , \4299 , \4309 );
not \U$3934 ( \4311 , \2341 );
not \U$3935 ( \4312 , \3674 );
or \U$3936 ( \4313 , \4311 , \4312 );
nand \U$3937 ( \4314 , \2322 , RIae798e0_154);
nand \U$3938 ( \4315 , \4313 , \4314 );
not \U$3939 ( \4316 , \4315 );
xnor \U$3940 ( \4317 , \4310 , \4316 );
xor \U$3941 ( \4318 , \4298 , \4317 );
not \U$3942 ( \4319 , \4318 );
not \U$3943 ( \4320 , \3756 );
nand \U$3944 ( \4321 , \4320 , \3726 );
not \U$3945 ( \4322 , \3752 );
nand \U$3946 ( \4323 , \4322 , \3736 );
and \U$3947 ( \4324 , \4321 , \4323 );
not \U$3948 ( \4325 , \4324 );
and \U$3949 ( \4326 , \4319 , \4325 );
and \U$3950 ( \4327 , \4318 , \4324 );
nor \U$3951 ( \4328 , \4326 , \4327 );
xor \U$3952 ( \4329 , \4292 , \4328 );
not \U$3953 ( \4330 , \3797 );
not \U$3954 ( \4331 , \3831 );
and \U$3955 ( \4332 , \4330 , \4331 );
and \U$3956 ( \4333 , \3835 , \3760 );
nor \U$3957 ( \4334 , \4332 , \4333 );
xor \U$3958 ( \4335 , \4329 , \4334 );
not \U$3959 ( \4336 , \4335 );
not \U$3960 ( \4337 , \2011 );
and \U$3961 ( \4338 , RIae79610_148, \1473 );
not \U$3962 ( \4339 , RIae79610_148);
and \U$3963 ( \4340 , \4339 , \1472 );
nor \U$3964 ( \4341 , \4338 , \4340 );
not \U$3965 ( \4342 , \4341 );
or \U$3966 ( \4343 , \4337 , \4342 );
buf \U$3967 ( \4344 , \2063 );
nand \U$3968 ( \4345 , \3724 , \4344 );
nand \U$3969 ( \4346 , \4343 , \4345 );
not \U$3970 ( \4347 , \2924 );
and \U$3971 ( \4348 , \1146 , \2183 );
not \U$3972 ( \4349 , \1146 );
and \U$3973 ( \4350 , \4349 , RIae79520_146);
nor \U$3974 ( \4351 , \4348 , \4350 );
not \U$3975 ( \4352 , \4351 );
or \U$3976 ( \4353 , \4347 , \4352 );
nand \U$3977 ( \4354 , \2602 , \3665 );
nand \U$3978 ( \4355 , \4353 , \4354 );
xor \U$3979 ( \4356 , \4346 , \4355 );
not \U$3980 ( \4357 , \840 );
not \U$3981 ( \4358 , \4081 );
xnor \U$3982 ( \4359 , \4358 , RIae78f80_134);
not \U$3983 ( \4360 , \4359 );
or \U$3984 ( \4361 , \4357 , \4360 );
not \U$3985 ( \4362 , \3802 );
or \U$3986 ( \4363 , \4362 , \798 );
nand \U$3987 ( \4364 , \4361 , \4363 );
xor \U$3988 ( \4365 , \4356 , \4364 );
xor \U$3989 ( \4366 , \3421 , \3426 );
and \U$3990 ( \4367 , \4366 , \3456 );
and \U$3991 ( \4368 , \3421 , \3426 );
or \U$3992 ( \4369 , \4367 , \4368 );
xor \U$3993 ( \4370 , \4365 , \4369 );
not \U$3994 ( \4371 , \3596 );
not \U$3995 ( \4372 , \3590 );
or \U$3996 ( \4373 , \4371 , \4372 );
nand \U$3997 ( \4374 , \3585 , \3589 );
nand \U$3998 ( \4375 , \4373 , \4374 );
xor \U$3999 ( \4376 , \4370 , \4375 );
and \U$4000 ( \4377 , \3580 , \3600 );
and \U$4001 ( \4378 , \3573 , \3579 );
nor \U$4002 ( \4379 , \4377 , \4378 );
xnor \U$4003 ( \4380 , \4376 , \4379 );
not \U$4004 ( \4381 , \4380 );
or \U$4005 ( \4382 , \4336 , \4381 );
or \U$4006 ( \4383 , \4380 , \4335 );
nand \U$4007 ( \4384 , \4382 , \4383 );
not \U$4008 ( \4385 , \4384 );
not \U$4009 ( \4386 , \3845 );
not \U$4010 ( \4387 , \3645 );
or \U$4011 ( \4388 , \4386 , \4387 );
not \U$4012 ( \4389 , \3712 );
nand \U$4013 ( \4390 , \4389 , \3841 );
nand \U$4014 ( \4391 , \4388 , \4390 );
not \U$4015 ( \4392 , \4391 );
not \U$4016 ( \4393 , \3708 );
not \U$4017 ( \4394 , \4393 );
not \U$4018 ( \4395 , \3683 );
or \U$4019 ( \4396 , \4394 , \4395 );
not \U$4020 ( \4397 , \3679 );
nand \U$4021 ( \4398 , \4397 , \3651 );
nand \U$4022 ( \4399 , \4396 , \4398 );
not \U$4023 ( \4400 , \4399 );
not \U$4024 ( \4401 , \1501 );
xnor \U$4025 ( \4402 , \2027 , RIae79250_140);
not \U$4026 ( \4403 , \4402 );
or \U$4027 ( \4404 , \4401 , \4403 );
nand \U$4028 ( \4405 , \3703 , \1499 );
nand \U$4029 ( \4406 , \4404 , \4405 );
not \U$4030 ( \4407 , \1933 );
not \U$4031 ( \4408 , \3816 );
or \U$4032 ( \4409 , \4407 , \4408 );
not \U$4033 ( \4410 , \3039 );
not \U$4034 ( \4411 , \2004 );
or \U$4035 ( \4412 , \4410 , \4411 );
not \U$4036 ( \4413 , \833 );
nand \U$4037 ( \4414 , \4413 , RIae794a8_145);
nand \U$4038 ( \4415 , \4412 , \4414 );
nand \U$4039 ( \4416 , \4415 , \1919 );
nand \U$4040 ( \4417 , \4409 , \4416 );
xor \U$4041 ( \4418 , \4406 , \4417 );
not \U$4042 ( \4419 , \3015 );
not \U$4043 ( \4420 , RIae79ac0_158);
not \U$4044 ( \4421 , \919 );
or \U$4045 ( \4422 , \4420 , \4421 );
nand \U$4046 ( \4423 , \918 , \2268 );
nand \U$4047 ( \4424 , \4422 , \4423 );
not \U$4048 ( \4425 , \4424 );
or \U$4049 ( \4426 , \4419 , \4425 );
nand \U$4050 ( \4427 , \3777 , \2272 );
nand \U$4051 ( \4428 , \4426 , \4427 );
xnor \U$4052 ( \4429 , \4418 , \4428 );
not \U$4053 ( \4430 , \929 );
not \U$4054 ( \4431 , \1739 );
xor \U$4055 ( \4432 , RIae78bc0_126, \4431 );
not \U$4056 ( \4433 , \4432 );
or \U$4057 ( \4434 , \4430 , \4433 );
nand \U$4058 ( \4435 , \3734 , \952 );
nand \U$4059 ( \4436 , \4434 , \4435 );
not \U$4060 ( \4437 , \1259 );
not \U$4061 ( \4438 , \3750 );
or \U$4062 ( \4439 , \4437 , \4438 );
and \U$4063 ( \4440 , \2309 , RIae78e90_132);
not \U$4064 ( \4441 , \2309 );
and \U$4065 ( \4442 , \4441 , \1066 );
nor \U$4066 ( \4443 , \4440 , \4442 );
nand \U$4067 ( \4444 , \4443 , \1321 );
nand \U$4068 ( \4445 , \4439 , \4444 );
xor \U$4069 ( \4446 , \4436 , \4445 );
and \U$4070 ( \4447 , RIae793b8_143, \1188 );
not \U$4071 ( \4448 , RIae793b8_143);
and \U$4072 ( \4449 , \4448 , \1187 );
or \U$4073 ( \4450 , \4447 , \4449 );
not \U$4074 ( \4451 , \4450 );
not \U$4075 ( \4452 , \3494 );
and \U$4076 ( \4453 , \4451 , \4452 );
and \U$4077 ( \4454 , \3693 , \1910 );
nor \U$4078 ( \4455 , \4453 , \4454 );
xor \U$4079 ( \4456 , \4446 , \4455 );
xor \U$4080 ( \4457 , \4429 , \4456 );
not \U$4081 ( \4458 , \1879 );
and \U$4082 ( \4459 , \4458 , \997 );
not \U$4083 ( \4460 , \4458 );
and \U$4084 ( \4461 , \4460 , RIae79160_138);
nor \U$4085 ( \4462 , \4459 , \4461 );
not \U$4086 ( \4463 , \4462 );
or \U$4087 ( \4464 , \4463 , \1210 );
not \U$4088 ( \4465 , \2157 );
or \U$4089 ( \4466 , \3789 , \4465 );
nand \U$4090 ( \4467 , \4464 , \4466 );
not \U$4091 ( \4468 , \3827 );
and \U$4092 ( \4469 , RIae79688_149, \856 );
not \U$4093 ( \4470 , RIae79688_149);
and \U$4094 ( \4471 , \4470 , \857 );
nor \U$4095 ( \4472 , \4469 , \4471 );
not \U$4096 ( \4473 , \4472 );
or \U$4097 ( \4474 , \4468 , \4473 );
nand \U$4098 ( \4475 , \3826 , \1844 );
nand \U$4099 ( \4476 , \4474 , \4475 );
xor \U$4100 ( \4477 , \4467 , \4476 );
not \U$4101 ( \4478 , \1049 );
not \U$4102 ( \4479 , \3052 );
not \U$4103 ( \4480 , \4479 );
and \U$4104 ( \4481 , \4480 , \1039 );
not \U$4105 ( \4482 , \4480 );
and \U$4106 ( \4483 , \4482 , RIae79070_136);
nor \U$4107 ( \4484 , \4481 , \4483 );
not \U$4108 ( \4485 , \4484 );
or \U$4109 ( \4486 , \4478 , \4485 );
nand \U$4110 ( \4487 , \3766 , \1062 );
nand \U$4111 ( \4488 , \4486 , \4487 );
buf \U$4112 ( \4489 , \4488 );
xnor \U$4113 ( \4490 , \4477 , \4489 );
xor \U$4114 ( \4491 , \4457 , \4490 );
not \U$4115 ( \4492 , \4491 );
or \U$4116 ( \4493 , \4400 , \4492 );
or \U$4117 ( \4494 , \4399 , \4491 );
nand \U$4118 ( \4495 , \4493 , \4494 );
not \U$4119 ( \4496 , \3477 );
nand \U$4120 ( \4497 , \4496 , \3407 );
not \U$4121 ( \4498 , \3407 );
not \U$4122 ( \4499 , \4498 );
not \U$4123 ( \4500 , \3477 );
or \U$4124 ( \4501 , \4499 , \4500 );
nand \U$4125 ( \4502 , \4501 , \3457 );
nand \U$4126 ( \4503 , \4497 , \4502 );
xnor \U$4127 ( \4504 , \4495 , \4503 );
not \U$4128 ( \4505 , \4504 );
or \U$4129 ( \4506 , \4392 , \4505 );
or \U$4130 ( \4507 , \4391 , \4504 );
nand \U$4131 ( \4508 , \4506 , \4507 );
not \U$4132 ( \4509 , \4508 );
xor \U$4133 ( \4510 , \3485 , \3568 );
and \U$4134 ( \4511 , \4510 , \3602 );
and \U$4135 ( \4512 , \3485 , \3568 );
or \U$4136 ( \4513 , \4511 , \4512 );
not \U$4137 ( \4514 , \4513 );
and \U$4138 ( \4515 , \4509 , \4514 );
and \U$4139 ( \4516 , \4508 , \4513 );
nor \U$4140 ( \4517 , \4515 , \4516 );
not \U$4141 ( \4518 , \4517 );
or \U$4142 ( \4519 , \4385 , \4518 );
buf \U$4143 ( \4520 , \4384 );
or \U$4144 ( \4521 , \4520 , \4517 );
nand \U$4145 ( \4522 , \4519 , \4521 );
not \U$4146 ( \4523 , \4522 );
or \U$4147 ( \4524 , \4262 , \4523 );
or \U$4148 ( \4525 , \4522 , \4261 );
nand \U$4149 ( \4526 , \4524 , \4525 );
nor \U$4150 ( \4527 , \4255 , \4526 );
not \U$4151 ( \4528 , \4527 );
not \U$4152 ( \4529 , \4335 );
not \U$4153 ( \4530 , \4529 );
not \U$4154 ( \4531 , \4380 );
or \U$4155 ( \4532 , \4530 , \4531 );
not \U$4156 ( \4533 , \4379 );
nand \U$4157 ( \4534 , \4533 , \4376 );
nand \U$4158 ( \4535 , \4532 , \4534 );
not \U$4159 ( \4536 , \4503 );
not \U$4160 ( \4537 , \4495 );
or \U$4161 ( \4538 , \4536 , \4537 );
not \U$4162 ( \4539 , \4491 );
nand \U$4163 ( \4540 , \4539 , \4399 );
nand \U$4164 ( \4541 , \4538 , \4540 );
and \U$4165 ( \4542 , RIae78bc0_126, \2287 );
not \U$4166 ( \4543 , RIae78bc0_126);
and \U$4167 ( \4544 , \4543 , \3748 );
nor \U$4168 ( \4545 , \4542 , \4544 );
not \U$4169 ( \4546 , \4545 );
not \U$4170 ( \4547 , \928 );
and \U$4171 ( \4548 , \4546 , \4547 );
and \U$4172 ( \4549 , \4432 , \953 );
nor \U$4173 ( \4550 , \4548 , \4549 );
not \U$4174 ( \4551 , \4550 );
not \U$4175 ( \4552 , \1087 );
not \U$4176 ( \4553 , \4443 );
or \U$4177 ( \4554 , \4552 , \4553 );
buf \U$4178 ( \4555 , \2155 );
and \U$4179 ( \4556 , \4555 , \921 );
not \U$4180 ( \4557 , \4555 );
and \U$4181 ( \4558 , \4557 , RIae78e90_132);
nor \U$4182 ( \4559 , \4556 , \4558 );
nand \U$4183 ( \4560 , \4559 , \1321 );
nand \U$4184 ( \4561 , \4554 , \4560 );
not \U$4185 ( \4562 , \4561 );
or \U$4186 ( \4563 , \4551 , \4562 );
or \U$4187 ( \4564 , \4561 , \4550 );
nand \U$4188 ( \4565 , \4563 , \4564 );
not \U$4189 ( \4566 , \2063 );
not \U$4190 ( \4567 , \4341 );
or \U$4191 ( \4568 , \4566 , \4567 );
and \U$4192 ( \4569 , RIae79610_148, \880 );
not \U$4193 ( \4570 , RIae79610_148);
and \U$4194 ( \4571 , \4570 , \879 );
nor \U$4195 ( \4572 , \4569 , \4571 );
nand \U$4196 ( \4573 , \4572 , \2011 );
nand \U$4197 ( \4574 , \4568 , \4573 );
xor \U$4198 ( \4575 , \4565 , \4574 );
not \U$4199 ( \4576 , \4575 );
not \U$4200 ( \4577 , \4576 );
and \U$4201 ( \4578 , RIae78b48_125, \2573 );
not \U$4202 ( \4579 , \893 );
not \U$4203 ( \4580 , \4307 );
or \U$4204 ( \4581 , \4579 , \4580 );
not \U$4205 ( \4582 , \1752 );
not \U$4206 ( \4583 , \4582 );
not \U$4207 ( \4584 , \4583 );
not \U$4208 ( \4585 , \4584 );
and \U$4209 ( \4586 , RIae78b48_125, \4585 );
not \U$4210 ( \4587 , RIae78b48_125);
and \U$4211 ( \4588 , \4587 , \4584 );
nor \U$4212 ( \4589 , \4586 , \4588 );
or \U$4213 ( \4590 , \4589 , \1959 );
nand \U$4214 ( \4591 , \4581 , \4590 );
xor \U$4215 ( \4592 , \4578 , \4591 );
not \U$4216 ( \4593 , RIae793b8_143);
not \U$4217 ( \4594 , \3722 );
or \U$4218 ( \4595 , \4593 , \4594 );
not \U$4219 ( \4596 , \978 );
nand \U$4220 ( \4597 , \4596 , \1884 );
nand \U$4221 ( \4598 , \4595 , \4597 );
not \U$4222 ( \4599 , \4598 );
not \U$4223 ( \4600 , \1864 );
or \U$4224 ( \4601 , \4599 , \4600 );
not \U$4225 ( \4602 , \4450 );
nand \U$4226 ( \4603 , \4602 , \1910 );
nand \U$4227 ( \4604 , \4601 , \4603 );
xnor \U$4228 ( \4605 , \4592 , \4604 );
nor \U$4229 ( \4606 , \2341 , \2322 );
nor \U$4230 ( \4607 , \4606 , \2334 );
not \U$4231 ( \4608 , \2272 );
not \U$4232 ( \4609 , \4424 );
or \U$4233 ( \4610 , \4608 , \4609 );
and \U$4234 ( \4611 , RIae79ac0_158, \1162 );
not \U$4235 ( \4612 , RIae79ac0_158);
and \U$4236 ( \4613 , \4612 , \1291 );
nor \U$4237 ( \4614 , \4611 , \4613 );
or \U$4238 ( \4615 , \4614 , \3016 );
nand \U$4239 ( \4616 , \4610 , \4615 );
xor \U$4240 ( \4617 , \4607 , \4616 );
not \U$4241 ( \4618 , \1919 );
not \U$4242 ( \4619 , \992 );
not \U$4243 ( \4620 , RIae794a8_145);
and \U$4244 ( \4621 , \4619 , \4620 );
and \U$4245 ( \4622 , \1196 , RIae794a8_145);
nor \U$4246 ( \4623 , \4621 , \4622 );
not \U$4247 ( \4624 , \4623 );
or \U$4248 ( \4625 , \4618 , \4624 );
nand \U$4249 ( \4626 , \4415 , \2458 );
nand \U$4250 ( \4627 , \4625 , \4626 );
xor \U$4251 ( \4628 , \4617 , \4627 );
not \U$4252 ( \4629 , \4628 );
and \U$4253 ( \4630 , \4605 , \4629 );
not \U$4254 ( \4631 , \4605 );
and \U$4255 ( \4632 , \4631 , \4628 );
or \U$4256 ( \4633 , \4630 , \4632 );
not \U$4257 ( \4634 , \4633 );
or \U$4258 ( \4635 , \4577 , \4634 );
or \U$4259 ( \4636 , \4633 , \4576 );
nand \U$4260 ( \4637 , \4635 , \4636 );
xor \U$4261 ( \4638 , \4429 , \4456 );
and \U$4262 ( \4639 , \4638 , \4490 );
and \U$4263 ( \4640 , \4429 , \4456 );
or \U$4264 ( \4641 , \4639 , \4640 );
not \U$4265 ( \4642 , \4641 );
xor \U$4266 ( \4643 , \4637 , \4642 );
not \U$4267 ( \4644 , \4299 );
xor \U$4268 ( \4645 , \4644 , \4316 );
and \U$4269 ( \4646 , \4645 , \4309 );
and \U$4270 ( \4647 , \4644 , \4316 );
nor \U$4271 ( \4648 , \4646 , \4647 );
not \U$4272 ( \4649 , \4648 );
not \U$4273 ( \4650 , \2189 );
not \U$4274 ( \4651 , \4351 );
or \U$4275 ( \4652 , \4650 , \4651 );
not \U$4276 ( \4653 , RIae79520_146);
not \U$4277 ( \4654 , \4653 );
not \U$4278 ( \4655 , \781 );
or \U$4279 ( \4656 , \4654 , \4655 );
nand \U$4280 ( \4657 , \3814 , RIae79520_146);
nand \U$4281 ( \4658 , \4656 , \4657 );
nand \U$4282 ( \4659 , \4658 , \2924 );
nand \U$4283 ( \4660 , \4652 , \4659 );
not \U$4284 ( \4661 , \1062 );
not \U$4285 ( \4662 , \4484 );
or \U$4286 ( \4663 , \4661 , \4662 );
and \U$4287 ( \4664 , RIae79070_136, \1899 );
not \U$4288 ( \4665 , RIae79070_136);
and \U$4289 ( \4666 , \4665 , \3785 );
nor \U$4290 ( \4667 , \4664 , \4666 );
nand \U$4291 ( \4668 , \4667 , \1049 );
nand \U$4292 ( \4669 , \4663 , \4668 );
xor \U$4293 ( \4670 , \4660 , \4669 );
not \U$4294 ( \4671 , \4670 );
not \U$4295 ( \4672 , \797 );
not \U$4296 ( \4673 , \4359 );
or \U$4297 ( \4674 , \4672 , \4673 );
not \U$4298 ( \4675 , \2231 );
and \U$4299 ( \4676 , \4675 , \1132 );
not \U$4300 ( \4677 , \4675 );
and \U$4301 ( \4678 , \4677 , RIae78f80_134);
nor \U$4302 ( \4679 , \4676 , \4678 );
nand \U$4303 ( \4680 , \4679 , \840 );
nand \U$4304 ( \4681 , \4674 , \4680 );
not \U$4305 ( \4682 , \4681 );
not \U$4306 ( \4683 , \4682 );
or \U$4307 ( \4684 , \4671 , \4683 );
or \U$4308 ( \4685 , \4682 , \4670 );
nand \U$4309 ( \4686 , \4684 , \4685 );
not \U$4310 ( \4687 , \4686 );
or \U$4311 ( \4688 , \4649 , \4687 );
or \U$4312 ( \4689 , \4648 , \4686 );
nand \U$4313 ( \4690 , \4688 , \4689 );
not \U$4314 ( \4691 , \4287 );
not \U$4315 ( \4692 , \4281 );
or \U$4316 ( \4693 , \4691 , \4692 );
nand \U$4317 ( \4694 , \4270 , \4280 );
nand \U$4318 ( \4695 , \4693 , \4694 );
xor \U$4319 ( \4696 , \4690 , \4695 );
xor \U$4320 ( \4697 , \4643 , \4696 );
nor \U$4321 ( \4698 , \4541 , \4697 );
not \U$4322 ( \4699 , \4698 );
nand \U$4323 ( \4700 , \4541 , \4697 );
nand \U$4324 ( \4701 , \4699 , \4700 );
xor \U$4325 ( \4702 , \4535 , \4701 );
not \U$4326 ( \4703 , \4702 );
not \U$4327 ( \4704 , \4703 );
xor \U$4328 ( \4705 , \4365 , \4369 );
and \U$4329 ( \4706 , \4705 , \4375 );
and \U$4330 ( \4707 , \4365 , \4369 );
or \U$4331 ( \4708 , \4706 , \4707 );
xor \U$4332 ( \4709 , \4292 , \4328 );
and \U$4333 ( \4710 , \4709 , \4334 );
and \U$4334 ( \4711 , \4292 , \4328 );
or \U$4335 ( \4712 , \4710 , \4711 );
xnor \U$4336 ( \4713 , \4708 , \4712 );
not \U$4337 ( \4714 , \4324 );
not \U$4338 ( \4715 , \4714 );
not \U$4339 ( \4716 , \4318 );
or \U$4340 ( \4717 , \4715 , \4716 );
nand \U$4341 ( \4718 , \4298 , \4317 );
nand \U$4342 ( \4719 , \4717 , \4718 );
not \U$4343 ( \4720 , \4406 );
not \U$4344 ( \4721 , \4417 );
or \U$4345 ( \4722 , \4720 , \4721 );
or \U$4346 ( \4723 , \4417 , \4406 );
nand \U$4347 ( \4724 , \4723 , \4428 );
nand \U$4348 ( \4725 , \4722 , \4724 );
xor \U$4349 ( \4726 , \4315 , \4725 );
not \U$4350 ( \4727 , \4467 );
xor \U$4351 ( \4728 , \4476 , \4488 );
not \U$4352 ( \4729 , \4728 );
or \U$4353 ( \4730 , \4727 , \4729 );
nand \U$4354 ( \4731 , \4489 , \4476 );
nand \U$4355 ( \4732 , \4730 , \4731 );
xnor \U$4356 ( \4733 , \4726 , \4732 );
xor \U$4357 ( \4734 , \4719 , \4733 );
not \U$4358 ( \4735 , \1209 );
and \U$4359 ( \4736 , \2594 , \997 );
not \U$4360 ( \4737 , \2594 );
and \U$4361 ( \4738 , \4737 , RIae79160_138);
nor \U$4362 ( \4739 , \4736 , \4738 );
not \U$4363 ( \4740 , \4739 );
or \U$4364 ( \4741 , \4735 , \4740 );
nand \U$4365 ( \4742 , \4462 , \1009 );
nand \U$4366 ( \4743 , \4741 , \4742 );
not \U$4367 ( \4744 , \1501 );
and \U$4368 ( \4745 , RIae79250_140, \1835 );
not \U$4369 ( \4746 , RIae79250_140);
and \U$4370 ( \4747 , \4746 , \2101 );
nor \U$4371 ( \4748 , \4745 , \4747 );
not \U$4372 ( \4749 , \4748 );
or \U$4373 ( \4750 , \4744 , \4749 );
nand \U$4374 ( \4751 , \4402 , \2650 );
nand \U$4375 ( \4752 , \4750 , \4751 );
xor \U$4376 ( \4753 , \4743 , \4752 );
not \U$4377 ( \4754 , \1844 );
not \U$4378 ( \4755 , \4472 );
or \U$4379 ( \4756 , \4754 , \4755 );
and \U$4380 ( \4757 , RIae79688_149, \940 );
not \U$4381 ( \4758 , RIae79688_149);
and \U$4382 ( \4759 , \4758 , \3236 );
or \U$4383 ( \4760 , \4757 , \4759 );
nand \U$4384 ( \4761 , \4760 , \1822 );
nand \U$4385 ( \4762 , \4756 , \4761 );
xor \U$4386 ( \4763 , \4753 , \4762 );
not \U$4387 ( \4764 , \4455 );
or \U$4388 ( \4765 , \4764 , \4445 );
nand \U$4389 ( \4766 , \4765 , \4436 );
nand \U$4390 ( \4767 , \4764 , \4445 );
nand \U$4391 ( \4768 , \4766 , \4767 );
xor \U$4392 ( \4769 , \4763 , \4768 );
not \U$4393 ( \4770 , \4364 );
not \U$4394 ( \4771 , \4356 );
or \U$4395 ( \4772 , \4770 , \4771 );
nand \U$4396 ( \4773 , \4346 , \4355 );
nand \U$4397 ( \4774 , \4772 , \4773 );
xnor \U$4398 ( \4775 , \4769 , \4774 );
not \U$4399 ( \4776 , \4775 );
xor \U$4400 ( \4777 , \4734 , \4776 );
and \U$4401 ( \4778 , \4713 , \4777 );
not \U$4402 ( \4779 , \4713 );
not \U$4403 ( \4780 , \4777 );
and \U$4404 ( \4781 , \4779 , \4780 );
or \U$4405 ( \4782 , \4778 , \4781 );
not \U$4406 ( \4783 , \4782 );
not \U$4407 ( \4784 , \4513 );
not \U$4408 ( \4785 , \4784 );
not \U$4409 ( \4786 , \4508 );
or \U$4410 ( \4787 , \4785 , \4786 );
not \U$4411 ( \4788 , \4504 );
nand \U$4412 ( \4789 , \4788 , \4391 );
nand \U$4413 ( \4790 , \4787 , \4789 );
not \U$4414 ( \4791 , \4790 );
not \U$4415 ( \4792 , \4791 );
or \U$4416 ( \4793 , \4783 , \4792 );
not \U$4417 ( \4794 , \4782 );
nand \U$4418 ( \4795 , \4794 , \4790 );
nand \U$4419 ( \4796 , \4793 , \4795 );
not \U$4420 ( \4797 , \4796 );
or \U$4421 ( \4798 , \4704 , \4797 );
or \U$4422 ( \4799 , \4796 , \4703 );
nand \U$4423 ( \4800 , \4798 , \4799 );
not \U$4424 ( \4801 , \4261 );
not \U$4425 ( \4802 , \4520 );
not \U$4426 ( \4803 , \4802 );
or \U$4427 ( \4804 , \4801 , \4803 );
not \U$4428 ( \4805 , \4260 );
not \U$4429 ( \4806 , \4520 );
or \U$4430 ( \4807 , \4805 , \4806 );
nand \U$4431 ( \4808 , \4807 , \4517 );
nand \U$4432 ( \4809 , \4804 , \4808 );
nand \U$4433 ( \4810 , \4800 , \4809 );
and \U$4434 ( \4811 , \4250 , \4528 , \4810 );
xnor \U$4435 ( \4812 , \3973 , \3976 );
not \U$4436 ( \4813 , \3910 );
nand \U$4437 ( \4814 , \4813 , \3912 );
not \U$4438 ( \4815 , \3913 );
and \U$4439 ( \4816 , \4814 , \4815 );
not \U$4440 ( \4817 , \4814 );
and \U$4441 ( \4818 , \4817 , \3913 );
nor \U$4442 ( \4819 , \4816 , \4818 );
xor \U$4443 ( \4820 , \4812 , \4819 );
not \U$4444 ( \4821 , \3899 );
not \U$4445 ( \4822 , \3881 );
and \U$4446 ( \4823 , \4821 , \4822 );
and \U$4447 ( \4824 , \3899 , \3881 );
nor \U$4448 ( \4825 , \4823 , \4824 );
not \U$4449 ( \4826 , \4825 );
xor \U$4450 ( \4827 , \3997 , \4007 );
xor \U$4451 ( \4828 , \4827 , \4017 );
xor \U$4452 ( \4829 , \4071 , \4077 );
xor \U$4453 ( \4830 , \4829 , \4089 );
xor \U$4454 ( \4831 , \4828 , \4830 );
not \U$4455 ( \4832 , \839 );
not \U$4456 ( \4833 , \2761 );
or \U$4457 ( \4834 , \4832 , \4833 );
and \U$4458 ( \4835 , RIae78f80_134, \2564 );
not \U$4459 ( \4836 , RIae78f80_134);
not \U$4460 ( \4837 , \3417 );
and \U$4461 ( \4838 , \4836 , \4837 );
or \U$4462 ( \4839 , \4835 , \4838 );
nand \U$4463 ( \4840 , \4839 , \797 );
nand \U$4464 ( \4841 , \4834 , \4840 );
buf \U$4465 ( \4842 , \4154 );
not \U$4466 ( \4843 , \4842 );
not \U$4467 ( \4844 , RIae79ca0_162);
not \U$4468 ( \4845 , \4844 );
not \U$4469 ( \4846 , \992 );
or \U$4470 ( \4847 , \4845 , \4846 );
or \U$4471 ( \4848 , \2444 , \4844 );
nand \U$4472 ( \4849 , \4847 , \4848 );
not \U$4473 ( \4850 , \4849 );
or \U$4474 ( \4851 , \4843 , \4850 );
not \U$4475 ( \4852 , \4155 );
not \U$4476 ( \4853 , \4852 );
nand \U$4477 ( \4854 , \4853 , RIae79ca0_162);
nand \U$4478 ( \4855 , \4851 , \4854 );
xor \U$4479 ( \4856 , \4841 , \4855 );
xor \U$4480 ( \4857 , \4176 , \4142 );
xor \U$4481 ( \4858 , \4856 , \4857 );
and \U$4482 ( \4859 , \4831 , \4858 );
and \U$4483 ( \4860 , \4828 , \4830 );
or \U$4484 ( \4861 , \4859 , \4860 );
not \U$4485 ( \4862 , \4861 );
not \U$4486 ( \4863 , \4862 );
and \U$4487 ( \4864 , \4826 , \4863 );
not \U$4488 ( \4865 , \4861 );
not \U$4489 ( \4866 , \4825 );
or \U$4490 ( \4867 , \4865 , \4866 );
or \U$4491 ( \4868 , \4825 , \4861 );
nand \U$4492 ( \4869 , \4867 , \4868 );
or \U$4493 ( \4870 , \3963 , \3953 );
nand \U$4494 ( \4871 , \4870 , \3964 );
not \U$4495 ( \4872 , \3967 );
and \U$4496 ( \4873 , \4871 , \4872 );
not \U$4497 ( \4874 , \4871 );
and \U$4498 ( \4875 , \4874 , \3967 );
nor \U$4499 ( \4876 , \4873 , \4875 );
and \U$4500 ( \4877 , \4869 , \4876 );
nor \U$4501 ( \4878 , \4864 , \4877 );
xor \U$4502 ( \4879 , \4820 , \4878 );
and \U$4503 ( \4880 , \4223 , \4135 );
not \U$4504 ( \4881 , \4223 );
not \U$4505 ( \4882 , \4135 );
and \U$4506 ( \4883 , \4881 , \4882 );
nor \U$4507 ( \4884 , \4880 , \4883 );
xor \U$4508 ( \4885 , \4109 , \4121 );
xnor \U$4509 ( \4886 , \4885 , \4133 );
not \U$4510 ( \4887 , \4886 );
not \U$4511 ( \4888 , \4887 );
xor \U$4512 ( \4889 , \4031 , \4043 );
xor \U$4513 ( \4890 , \4889 , \4054 );
not \U$4514 ( \4891 , \4890 );
not \U$4515 ( \4892 , \4891 );
or \U$4516 ( \4893 , \4888 , \4892 );
not \U$4517 ( \4894 , \4886 );
not \U$4518 ( \4895 , \4890 );
or \U$4519 ( \4896 , \4894 , \4895 );
not \U$4520 ( \4897 , \4203 );
xor \U$4521 ( \4898 , \4216 , \4897 );
not \U$4522 ( \4899 , \4189 );
xnor \U$4523 ( \4900 , \4898 , \4899 );
not \U$4524 ( \4901 , \4900 );
nand \U$4525 ( \4902 , \4896 , \4901 );
nand \U$4526 ( \4903 , \4893 , \4902 );
xor \U$4527 ( \4904 , \4884 , \4903 );
xor \U$4528 ( \4905 , \4020 , \4058 );
xor \U$4529 ( \4906 , \4905 , \4092 );
xor \U$4530 ( \4907 , \4904 , \4906 );
xor \U$4531 ( \4908 , \4828 , \4830 );
xor \U$4532 ( \4909 , \4908 , \4858 );
not \U$4533 ( \4910 , \4909 );
and \U$4534 ( \4911 , \4900 , \4891 );
not \U$4535 ( \4912 , \4900 );
and \U$4536 ( \4913 , \4912 , \4890 );
or \U$4537 ( \4914 , \4911 , \4913 );
and \U$4538 ( \4915 , \4914 , \4887 );
not \U$4539 ( \4916 , \4914 );
and \U$4540 ( \4917 , \4916 , \4886 );
nor \U$4541 ( \4918 , \4915 , \4917 );
not \U$4542 ( \4919 , \4918 );
or \U$4543 ( \4920 , \4910 , \4919 );
not \U$4544 ( \4921 , \1129 );
not \U$4545 ( \4922 , \4163 );
not \U$4546 ( \4923 , \4164 );
and \U$4547 ( \4924 , \4922 , \4923 );
and \U$4548 ( \4925 , \4163 , \4164 );
nor \U$4549 ( \4926 , \4924 , \4925 );
not \U$4550 ( \4927 , \4926 );
not \U$4551 ( \4928 , \4927 );
buf \U$4552 ( \4929 , \4928 );
and \U$4553 ( \4930 , RIae78b48_125, \4929 );
not \U$4554 ( \4931 , RIae78b48_125);
and \U$4555 ( \4932 , \4931 , \4169 );
or \U$4556 ( \4933 , \4930 , \4932 );
not \U$4557 ( \4934 , \4933 );
or \U$4558 ( \4935 , \4921 , \4934 );
nand \U$4559 ( \4936 , \4138 , \868 );
nand \U$4560 ( \4937 , \4935 , \4936 );
not \U$4561 ( \4938 , \2252 );
not \U$4562 ( \4939 , \4131 );
or \U$4563 ( \4940 , \4938 , \4939 );
not \U$4564 ( \4941 , RIae79ac0_158);
not \U$4565 ( \4942 , \3141 );
or \U$4566 ( \4943 , \4941 , \4942 );
or \U$4567 ( \4944 , \2594 , RIae79ac0_158);
nand \U$4568 ( \4945 , \4943 , \4944 );
nand \U$4569 ( \4946 , \4945 , \2272 );
nand \U$4570 ( \4947 , \4940 , \4946 );
xor \U$4571 ( \4948 , \4937 , \4947 );
not \U$4572 ( \4949 , \3155 );
not \U$4573 ( \4950 , \3198 );
or \U$4574 ( \4951 , \4949 , \4950 );
buf \U$4575 ( \4952 , \598 );
nand \U$4576 ( \4953 , \4951 , \4952 );
not \U$4577 ( \4954 , \4953 );
xnor \U$4578 ( \4955 , RIae788f0_120, RIae78878_119);
not \U$4579 ( \4956 , \4955 );
and \U$4580 ( \4957 , \4954 , \4956 );
and \U$4581 ( \4958 , \4953 , \4955 );
nor \U$4582 ( \4959 , \4957 , \4958 );
buf \U$4583 ( \4960 , \4959 );
not \U$4584 ( \4961 , \4960 );
nand \U$4585 ( \4962 , \4961 , RIae78b48_125);
not \U$4586 ( \4963 , \4962 );
xor \U$4587 ( \4964 , \4948 , \4963 );
not \U$4588 ( \4965 , \4855 );
not \U$4589 ( \4966 , \4965 );
and \U$4590 ( \4967 , RIae79e80_166, RIae79ef8_167);
not \U$4591 ( \4968 , RIae79d90_164);
nor \U$4592 ( \4969 , \4967 , \4968 );
not \U$4593 ( \4970 , \4969 );
not \U$4594 ( \4971 , \893 );
not \U$4595 ( \4972 , \4960 );
xor \U$4596 ( \4973 , \4972 , RIae78b48_125);
not \U$4597 ( \4974 , \4973 );
or \U$4598 ( \4975 , \4971 , \4974 );
nand \U$4599 ( \4976 , \4933 , \2096 );
nand \U$4600 ( \4977 , \4975 , \4976 );
not \U$4601 ( \4978 , \4977 );
not \U$4602 ( \4979 , \4978 );
or \U$4603 ( \4980 , \4970 , \4979 );
not \U$4604 ( \4981 , \952 );
buf \U$4605 ( \4982 , \3206 );
xor \U$4606 ( \4983 , \4982 , RIae78bc0_126);
not \U$4607 ( \4984 , \4983 );
or \U$4608 ( \4985 , \4981 , \4984 );
and \U$4609 ( \4986 , \1286 , \2403 );
not \U$4610 ( \4987 , \1286 );
and \U$4611 ( \4988 , \4987 , \3269 );
nor \U$4612 ( \4989 , \4986 , \4988 );
nand \U$4613 ( \4990 , \4989 , \1027 );
nand \U$4614 ( \4991 , \4985 , \4990 );
nand \U$4615 ( \4992 , \4980 , \4991 );
not \U$4616 ( \4993 , \4969 );
nand \U$4617 ( \4994 , \4977 , \4993 );
nand \U$4618 ( \4995 , \4992 , \4994 );
not \U$4619 ( \4996 , \4995 );
not \U$4620 ( \4997 , \4996 );
or \U$4621 ( \4998 , \4966 , \4997 );
not \U$4622 ( \4999 , \4994 );
not \U$4623 ( \5000 , \4992 );
or \U$4624 ( \5001 , \4999 , \5000 );
nand \U$4625 ( \5002 , \5001 , \4855 );
nand \U$4626 ( \5003 , \4998 , \5002 );
xor \U$4627 ( \5004 , \4964 , \5003 );
not \U$4628 ( \5005 , \2157 );
and \U$4629 ( \5006 , \3525 , \997 );
not \U$4630 ( \5007 , \3525 );
and \U$4631 ( \5008 , \5007 , RIae79160_138);
nor \U$4632 ( \5009 , \5006 , \5008 );
not \U$4633 ( \5010 , \5009 );
or \U$4634 ( \5011 , \5005 , \5010 );
and \U$4635 ( \5012 , RIae79160_138, \4584 );
not \U$4636 ( \5013 , RIae79160_138);
and \U$4637 ( \5014 , \5013 , \4585 );
nor \U$4638 ( \5015 , \5012 , \5014 );
nand \U$4639 ( \5016 , \5015 , \1209 );
nand \U$4640 ( \5017 , \5011 , \5016 );
not \U$4641 ( \5018 , \5017 );
not \U$4642 ( \5019 , \1049 );
buf \U$4643 ( \5020 , \1789 );
and \U$4644 ( \5021 , \5020 , \1039 );
not \U$4645 ( \5022 , \5020 );
and \U$4646 ( \5023 , \5022 , RIae79070_136);
nor \U$4647 ( \5024 , \5021 , \5023 );
not \U$4648 ( \5025 , \5024 );
or \U$4649 ( \5026 , \5019 , \5025 );
xnor \U$4650 ( \5027 , RIae79070_136, \3417 );
nand \U$4651 ( \5028 , \5027 , \2276 );
nand \U$4652 ( \5029 , \5026 , \5028 );
not \U$4653 ( \5030 , RIae79e80_166);
and \U$4654 ( \5031 , RIae79ef8_167, \5030 );
not \U$4655 ( \5032 , RIae79ef8_167);
and \U$4656 ( \5033 , \5032 , RIae79e80_166);
nor \U$4657 ( \5034 , \5031 , \5033 );
and \U$4658 ( \5035 , RIae79d90_164, RIae79e80_166);
not \U$4659 ( \5036 , RIae79d90_164);
and \U$4660 ( \5037 , \5036 , \5030 );
nor \U$4661 ( \5038 , \5035 , \5037 );
and \U$4662 ( \5039 , \5034 , \5038 );
buf \U$4663 ( \5040 , \5039 );
not \U$4664 ( \5041 , \5040 );
and \U$4665 ( \5042 , RIae79d90_164, \1194 );
not \U$4666 ( \5043 , RIae79d90_164);
and \U$4667 ( \5044 , \5043 , \991 );
or \U$4668 ( \5045 , \5042 , \5044 );
not \U$4669 ( \5046 , \5045 );
or \U$4670 ( \5047 , \5041 , \5046 );
not \U$4671 ( \5048 , \5034 );
buf \U$4672 ( \5049 , \5048 );
nand \U$4673 ( \5050 , \5049 , RIae79d90_164);
nand \U$4674 ( \5051 , \5047 , \5050 );
buf \U$4675 ( \5052 , \5051 );
xor \U$4676 ( \5053 , \5029 , \5052 );
not \U$4677 ( \5054 , \5053 );
or \U$4678 ( \5055 , \5018 , \5054 );
nand \U$4679 ( \5056 , \5052 , \5029 );
nand \U$4680 ( \5057 , \5055 , \5056 );
not \U$4681 ( \5058 , \5057 );
not \U$4682 ( \5059 , \2650 );
not \U$4683 ( \5060 , RIae79250_140);
not \U$4684 ( \5061 , \2287 );
or \U$4685 ( \5062 , \5060 , \5061 );
nand \U$4686 ( \5063 , \3748 , \1503 );
nand \U$4687 ( \5064 , \5062 , \5063 );
not \U$4688 ( \5065 , \5064 );
or \U$4689 ( \5066 , \5059 , \5065 );
nand \U$4690 ( \5067 , \3995 , \1501 );
nand \U$4691 ( \5068 , \5066 , \5067 );
not \U$4692 ( \5069 , \1013 );
not \U$4693 ( \5070 , \4026 );
or \U$4694 ( \5071 , \5069 , \5070 );
nand \U$4695 ( \5072 , \5015 , \1009 );
nand \U$4696 ( \5073 , \5071 , \5072 );
xor \U$4697 ( \5074 , \5068 , \5073 );
not \U$4698 ( \5075 , \1919 );
not \U$4699 ( \5076 , \4013 );
or \U$4700 ( \5077 , \5075 , \5076 );
not \U$4701 ( \5078 , RIae794a8_145);
not \U$4702 ( \5079 , \1125 );
or \U$4703 ( \5080 , \5078 , \5079 );
buf \U$4704 ( \5081 , \974 );
not \U$4705 ( \5082 , \5081 );
nand \U$4706 ( \5083 , \5082 , \3810 );
nand \U$4707 ( \5084 , \5080 , \5083 );
nand \U$4708 ( \5085 , \5084 , \1933 );
nand \U$4709 ( \5086 , \5077 , \5085 );
not \U$4710 ( \5087 , \5086 );
xor \U$4711 ( \5088 , \5074 , \5087 );
nand \U$4712 ( \5089 , \5058 , \5088 );
and \U$4713 ( \5090 , \5004 , \5089 );
nor \U$4714 ( \5091 , \5058 , \5088 );
nor \U$4715 ( \5092 , \5090 , \5091 );
nand \U$4716 ( \5093 , \4920 , \5092 );
not \U$4717 ( \5094 , \4909 );
not \U$4718 ( \5095 , \4918 );
nand \U$4719 ( \5096 , \5094 , \5095 );
nand \U$4720 ( \5097 , \5093 , \5096 );
xor \U$4721 ( \5098 , \4907 , \5097 );
xor \U$4722 ( \5099 , \4869 , \4876 );
xor \U$4723 ( \5100 , \5098 , \5099 );
nand \U$4724 ( \5101 , \3155 , \4952 );
buf \U$4725 ( \5102 , \3198 );
or \U$4726 ( \5103 , \5101 , \5102 );
nand \U$4727 ( \5104 , \3155 , \4952 );
nand \U$4728 ( \5105 , \5102 , \5104 );
nand \U$4729 ( \5106 , \5103 , \5105 );
buf \U$4730 ( \5107 , \5106 );
not \U$4731 ( \5108 , \5107 );
not \U$4732 ( \5109 , \5108 );
and \U$4733 ( \5110 , RIae78b48_125, \5109 );
not \U$4734 ( \5111 , \797 );
not \U$4735 ( \5112 , RIae78f80_134);
not \U$4736 ( \5113 , \2358 );
or \U$4737 ( \5114 , \5112 , \5113 );
not \U$4738 ( \5115 , \1955 );
nand \U$4739 ( \5116 , \5115 , \3105 );
nand \U$4740 ( \5117 , \5114 , \5116 );
not \U$4741 ( \5118 , \5117 );
or \U$4742 ( \5119 , \5111 , \5118 );
and \U$4743 ( \5120 , RIae78f80_134, \2093 );
not \U$4744 ( \5121 , RIae78f80_134);
and \U$4745 ( \5122 , \5121 , \2786 );
nor \U$4746 ( \5123 , \5120 , \5122 );
buf \U$4747 ( \5124 , \839 );
nand \U$4748 ( \5125 , \5123 , \5124 );
nand \U$4749 ( \5126 , \5119 , \5125 );
xor \U$4750 ( \5127 , \5110 , \5126 );
and \U$4751 ( \5128 , RIae79520_146, \1405 );
not \U$4752 ( \5129 , RIae79520_146);
and \U$4753 ( \5130 , \5129 , \2102 );
nor \U$4754 ( \5131 , \5128 , \5130 );
not \U$4755 ( \5132 , \3440 );
or \U$4756 ( \5133 , \5131 , \5132 );
not \U$4757 ( \5134 , \2025 );
and \U$4758 ( \5135 , RIae79520_146, \5134 );
not \U$4759 ( \5136 , RIae79520_146);
not \U$4760 ( \5137 , \2027 );
and \U$4761 ( \5138 , \5136 , \5137 );
nor \U$4762 ( \5139 , \5135 , \5138 );
not \U$4763 ( \5140 , \2602 );
or \U$4764 ( \5141 , \5139 , \5140 );
nand \U$4765 ( \5142 , \5133 , \5141 );
and \U$4766 ( \5143 , \5127 , \5142 );
and \U$4767 ( \5144 , \5110 , \5126 );
or \U$4768 ( \5145 , \5143 , \5144 );
not \U$4769 ( \5146 , \5145 );
not \U$4770 ( \5147 , \5146 );
not \U$4771 ( \5148 , \1259 );
and \U$4772 ( \5149 , RIae78e90_132, \1860 );
not \U$4773 ( \5150 , RIae78e90_132);
and \U$4774 ( \5151 , \5150 , \2385 );
or \U$4775 ( \5152 , \5149 , \5151 );
not \U$4776 ( \5153 , \5152 );
or \U$4777 ( \5154 , \5148 , \5153 );
and \U$4778 ( \5155 , RIae78e90_132, \3216 );
not \U$4779 ( \5156 , RIae78e90_132);
and \U$4780 ( \5157 , \5156 , \1973 );
or \U$4781 ( \5158 , \5155 , \5157 );
nand \U$4782 ( \5159 , \5158 , \1074 );
nand \U$4783 ( \5160 , \5154 , \5159 );
not \U$4784 ( \5161 , \2272 );
not \U$4785 ( \5162 , \1878 );
xor \U$4786 ( \5163 , \5162 , RIae79ac0_158);
not \U$4787 ( \5164 , \5163 );
or \U$4788 ( \5165 , \5161 , \5164 );
nand \U$4789 ( \5166 , \4945 , \3014 );
nand \U$4790 ( \5167 , \5165 , \5166 );
xor \U$4791 ( \5168 , \5160 , \5167 );
not \U$4792 ( \5169 , \4842 );
not \U$4793 ( \5170 , RIae79ca0_162);
not \U$4794 ( \5171 , \4413 );
or \U$4795 ( \5172 , \5170 , \5171 );
or \U$4796 ( \5173 , \3431 , RIae79ca0_162);
nand \U$4797 ( \5174 , \5172 , \5173 );
not \U$4798 ( \5175 , \5174 );
or \U$4799 ( \5176 , \5169 , \5175 );
nand \U$4800 ( \5177 , \4849 , \4853 );
nand \U$4801 ( \5178 , \5176 , \5177 );
and \U$4802 ( \5179 , \5168 , \5178 );
and \U$4803 ( \5180 , \5160 , \5167 );
or \U$4804 ( \5181 , \5179 , \5180 );
not \U$4805 ( \5182 , \5181 );
not \U$4806 ( \5183 , \5182 );
or \U$4807 ( \5184 , \5147 , \5183 );
not \U$4808 ( \5185 , \5145 );
not \U$4809 ( \5186 , \5181 );
or \U$4810 ( \5187 , \5185 , \5186 );
not \U$4811 ( \5188 , \2529 );
and \U$4812 ( \5189 , RIae797f0_152, \1024 );
not \U$4813 ( \5190 , RIae797f0_152);
not \U$4814 ( \5191 , \2169 );
and \U$4815 ( \5192 , \5190 , \5191 );
or \U$4816 ( \5193 , \5189 , \5192 );
not \U$4817 ( \5194 , \5193 );
or \U$4818 ( \5195 , \5188 , \5194 );
not \U$4819 ( \5196 , \1991 );
not \U$4820 ( \5197 , \3236 );
or \U$4821 ( \5198 , \5196 , \5197 );
nand \U$4822 ( \5199 , \940 , RIae797f0_152);
nand \U$4823 ( \5200 , \5198 , \5199 );
nand \U$4824 ( \5201 , \5200 , \2519 );
nand \U$4825 ( \5202 , \5195 , \5201 );
not \U$4826 ( \5203 , \2433 );
not \U$4827 ( \5204 , RIae79778_151);
not \U$4828 ( \5205 , \1439 );
or \U$4829 ( \5206 , \5204 , \5205 );
or \U$4830 ( \5207 , \919 , RIae79778_151);
nand \U$4831 ( \5208 , \5206 , \5207 );
not \U$4832 ( \5209 , \5208 );
or \U$4833 ( \5210 , \5203 , \5209 );
not \U$4834 ( \5211 , \2447 );
not \U$4835 ( \5212 , \1291 );
or \U$4836 ( \5213 , \5211 , \5212 );
nand \U$4837 ( \5214 , \1158 , RIae79778_151);
nand \U$4838 ( \5215 , \5213 , \5214 );
nand \U$4839 ( \5216 , \5215 , \2450 );
nand \U$4840 ( \5217 , \5210 , \5216 );
nand \U$4841 ( \5218 , \5202 , \5217 );
not \U$4842 ( \5219 , \5218 );
and \U$4843 ( \5220 , RIae79688_149, \4479 );
not \U$4844 ( \5221 , RIae79688_149);
not \U$4845 ( \5222 , \3055 );
and \U$4846 ( \5223 , \5221 , \5222 );
nor \U$4847 ( \5224 , \5220 , \5223 );
and \U$4848 ( \5225 , \5224 , \2966 );
not \U$4849 ( \5226 , \3147 );
not \U$4850 ( \5227 , \3294 );
or \U$4851 ( \5228 , \5226 , \5227 );
not \U$4852 ( \5229 , RIae79688_149);
or \U$4853 ( \5230 , \1899 , \5229 );
nand \U$4854 ( \5231 , \5228 , \5230 );
and \U$4855 ( \5232 , \5231 , \3827 );
nor \U$4856 ( \5233 , \5225 , \5232 );
not \U$4857 ( \5234 , \5233 );
or \U$4858 ( \5235 , \5219 , \5234 );
or \U$4859 ( \5236 , \5202 , \5217 );
nand \U$4860 ( \5237 , \5235 , \5236 );
nand \U$4861 ( \5238 , \5187 , \5237 );
nand \U$4862 ( \5239 , \5184 , \5238 );
not \U$4863 ( \5240 , \5239 );
not \U$4864 ( \5241 , \4964 );
not \U$4865 ( \5242 , \5003 );
or \U$4866 ( \5243 , \5241 , \5242 );
nand \U$4867 ( \5244 , \4995 , \4965 );
nand \U$4868 ( \5245 , \5243 , \5244 );
not \U$4869 ( \5246 , \5245 );
not \U$4870 ( \5247 , \5246 );
or \U$4871 ( \5248 , \5240 , \5247 );
not \U$4872 ( \5249 , \5239 );
not \U$4873 ( \5250 , \5249 );
not \U$4874 ( \5251 , \5245 );
or \U$4875 ( \5252 , \5250 , \5251 );
not \U$4876 ( \5253 , \2650 );
not \U$4877 ( \5254 , RIae79250_140);
not \U$4878 ( \5255 , \4024 );
or \U$4879 ( \5256 , \5254 , \5255 );
nand \U$4880 ( \5257 , \3099 , \1503 );
nand \U$4881 ( \5258 , \5256 , \5257 );
not \U$4882 ( \5259 , \5258 );
or \U$4883 ( \5260 , \5253 , \5259 );
nand \U$4884 ( \5261 , \5064 , \1501 );
nand \U$4885 ( \5262 , \5260 , \5261 );
not \U$4886 ( \5263 , \1864 );
and \U$4887 ( \5264 , \2154 , RIae793b8_143);
not \U$4888 ( \5265 , \2154 );
and \U$4889 ( \5266 , \5265 , \1902 );
nor \U$4890 ( \5267 , \5264 , \5266 );
not \U$4891 ( \5268 , \5267 );
or \U$4892 ( \5269 , \5263 , \5268 );
and \U$4893 ( \5270 , \2310 , RIae793b8_143);
not \U$4894 ( \5271 , \2310 );
and \U$4895 ( \5272 , \5271 , \1884 );
nor \U$4896 ( \5273 , \5270 , \5272 );
nand \U$4897 ( \5274 , \5273 , \1910 );
nand \U$4898 ( \5275 , \5269 , \5274 );
xor \U$4899 ( \5276 , \5262 , \5275 );
not \U$4900 ( \5277 , \1933 );
not \U$4901 ( \5278 , RIae794a8_145);
not \U$4902 ( \5279 , \1186 );
or \U$4903 ( \5280 , \5278 , \5279 );
nand \U$4904 ( \5281 , \1826 , \3039 );
nand \U$4905 ( \5282 , \5280 , \5281 );
not \U$4906 ( \5283 , \5282 );
or \U$4907 ( \5284 , \5277 , \5283 );
buf \U$4908 ( \5285 , \2467 );
nand \U$4909 ( \5286 , \5084 , \5285 );
nand \U$4910 ( \5287 , \5284 , \5286 );
and \U$4911 ( \5288 , \5276 , \5287 );
and \U$4912 ( \5289 , \5262 , \5275 );
or \U$4913 ( \5290 , \5288 , \5289 );
not \U$4914 ( \5291 , \5290 );
not \U$4915 ( \5292 , \839 );
not \U$4916 ( \5293 , \4839 );
or \U$4917 ( \5294 , \5292 , \5293 );
nand \U$4918 ( \5295 , \5123 , \797 );
nand \U$4919 ( \5296 , \5294 , \5295 );
not \U$4920 ( \5297 , \1062 );
not \U$4921 ( \5298 , \5024 );
or \U$4922 ( \5299 , \5297 , \5298 );
nand \U$4923 ( \5300 , \4038 , \1049 );
nand \U$4924 ( \5301 , \5299 , \5300 );
xor \U$4925 ( \5302 , \5296 , \5301 );
not \U$4926 ( \5303 , \2610 );
not \U$4927 ( \5304 , \4050 );
or \U$4928 ( \5305 , \5303 , \5304 );
not \U$4929 ( \5306 , \5131 );
nand \U$4930 ( \5307 , \5306 , \2602 );
nand \U$4931 ( \5308 , \5305 , \5307 );
xor \U$4932 ( \5309 , \5302 , \5308 );
not \U$4933 ( \5310 , \5309 );
or \U$4934 ( \5311 , \5291 , \5310 );
not \U$4935 ( \5312 , \2767 );
and \U$4936 ( \5313 , RIae79c28_161, \1147 );
not \U$4937 ( \5314 , RIae79c28_161);
and \U$4938 ( \5315 , \5314 , \1146 );
nor \U$4939 ( \5316 , \5313 , \5315 );
not \U$4940 ( \5317 , \5316 );
or \U$4941 ( \5318 , \5312 , \5317 );
and \U$4942 ( \5319 , RIae79c28_161, \780 );
not \U$4943 ( \5320 , RIae79c28_161);
and \U$4944 ( \5321 , \5320 , \3283 );
or \U$4945 ( \5322 , \5319 , \5321 );
not \U$4946 ( \5323 , \2776 );
not \U$4947 ( \5324 , \5323 );
nand \U$4948 ( \5325 , \5322 , \5324 );
nand \U$4949 ( \5326 , \5318 , \5325 );
not \U$4950 ( \5327 , \2011 );
and \U$4951 ( \5328 , RIae79610_148, \2995 );
not \U$4952 ( \5329 , RIae79610_148);
not \U$4953 ( \5330 , \3245 );
and \U$4954 ( \5331 , \5329 , \5330 );
nor \U$4955 ( \5332 , \5328 , \5331 );
not \U$4956 ( \5333 , \5332 );
or \U$4957 ( \5334 , \5327 , \5333 );
not \U$4958 ( \5335 , \2137 );
and \U$4959 ( \5336 , RIae79610_148, \5335 );
not \U$4960 ( \5337 , RIae79610_148);
and \U$4961 ( \5338 , \5337 , \2137 );
nor \U$4962 ( \5339 , \5336 , \5338 );
nand \U$4963 ( \5340 , \5339 , \4344 );
nand \U$4964 ( \5341 , \5334 , \5340 );
xor \U$4965 ( \5342 , \5326 , \5341 );
not \U$4966 ( \5343 , \2341 );
not \U$4967 ( \5344 , RIae798e0_154);
and \U$4968 ( \5345 , \5344 , \1472 );
not \U$4969 ( \5346 , \5344 );
and \U$4970 ( \5347 , \5346 , \1120 );
nor \U$4971 ( \5348 , \5345 , \5347 );
not \U$4972 ( \5349 , \5348 );
or \U$4973 ( \5350 , \5343 , \5349 );
not \U$4974 ( \5351 , \2175 );
xor \U$4975 ( \5352 , \5351 , RIae798e0_154);
nand \U$4976 ( \5353 , \5352 , \2322 );
nand \U$4977 ( \5354 , \5350 , \5353 );
and \U$4978 ( \5355 , \5342 , \5354 );
and \U$4979 ( \5356 , \5326 , \5341 );
or \U$4980 ( \5357 , \5355 , \5356 );
not \U$4981 ( \5358 , \5357 );
nand \U$4982 ( \5359 , \5311 , \5358 );
not \U$4983 ( \5360 , \5290 );
not \U$4984 ( \5361 , \5309 );
nand \U$4985 ( \5362 , \5360 , \5361 );
nand \U$4986 ( \5363 , \5359 , \5362 );
nand \U$4987 ( \5364 , \5252 , \5363 );
nand \U$4988 ( \5365 , \5248 , \5364 );
not \U$4989 ( \5366 , \5365 );
not \U$4990 ( \5367 , \4841 );
not \U$4991 ( \5368 , \4857 );
nand \U$4992 ( \5369 , \5368 , \4965 );
not \U$4993 ( \5370 , \5369 );
or \U$4994 ( \5371 , \5367 , \5370 );
nand \U$4995 ( \5372 , \4857 , \4855 );
nand \U$4996 ( \5373 , \5371 , \5372 );
not \U$4997 ( \5374 , \1321 );
not \U$4998 ( \5375 , \4117 );
or \U$4999 ( \5376 , \5374 , \5375 );
nand \U$5000 ( \5377 , \5158 , \1259 );
nand \U$5001 ( \5378 , \5376 , \5377 );
not \U$5002 ( \5379 , \5378 );
and \U$5003 ( \5380 , \4105 , \929 );
and \U$5004 ( \5381 , \4989 , \952 );
nor \U$5005 ( \5382 , \5380 , \5381 );
nand \U$5006 ( \5383 , \5379 , \5382 );
not \U$5007 ( \5384 , \5383 );
not \U$5008 ( \5385 , \2767 );
not \U$5009 ( \5386 , \5322 );
or \U$5010 ( \5387 , \5385 , \5386 );
nand \U$5011 ( \5388 , \4187 , \5324 );
nand \U$5012 ( \5389 , \5387 , \5388 );
not \U$5013 ( \5390 , \5389 );
or \U$5014 ( \5391 , \5384 , \5390 );
not \U$5015 ( \5392 , \5382 );
nand \U$5016 ( \5393 , \5378 , \5392 );
nand \U$5017 ( \5394 , \5391 , \5393 );
not \U$5018 ( \5395 , \3827 );
not \U$5019 ( \5396 , \4201 );
or \U$5020 ( \5397 , \5395 , \5396 );
nand \U$5021 ( \5398 , \5231 , \2966 );
nand \U$5022 ( \5399 , \5397 , \5398 );
not \U$5023 ( \5400 , \5399 );
not \U$5024 ( \5401 , \2322 );
not \U$5025 ( \5402 , \4073 );
or \U$5026 ( \5403 , \5401 , \5402 );
nand \U$5027 ( \5404 , \5352 , \2341 );
nand \U$5028 ( \5405 , \5403 , \5404 );
not \U$5029 ( \5406 , \5405 );
or \U$5030 ( \5407 , \5400 , \5406 );
or \U$5031 ( \5408 , \5405 , \5399 );
not \U$5032 ( \5409 , \2007 );
not \U$5033 ( \5410 , \4212 );
or \U$5034 ( \5411 , \5409 , \5410 );
nand \U$5035 ( \5412 , \5200 , \2529 );
nand \U$5036 ( \5413 , \5411 , \5412 );
nand \U$5037 ( \5414 , \5408 , \5413 );
nand \U$5038 ( \5415 , \5407 , \5414 );
xor \U$5039 ( \5416 , \5394 , \5415 );
xor \U$5040 ( \5417 , \4937 , \4947 );
not \U$5041 ( \5418 , \4962 );
and \U$5042 ( \5419 , \5417 , \5418 );
and \U$5043 ( \5420 , \4937 , \4947 );
or \U$5044 ( \5421 , \5419 , \5420 );
and \U$5045 ( \5422 , \5416 , \5421 );
and \U$5046 ( \5423 , \5394 , \5415 );
or \U$5047 ( \5424 , \5422 , \5423 );
xor \U$5048 ( \5425 , \5373 , \5424 );
not \U$5049 ( \5426 , \5425 );
xor \U$5050 ( \5427 , \5296 , \5301 );
and \U$5051 ( \5428 , \5427 , \5308 );
and \U$5052 ( \5429 , \5296 , \5301 );
or \U$5053 ( \5430 , \5428 , \5429 );
not \U$5054 ( \5431 , \5430 );
or \U$5055 ( \5432 , \5073 , \5068 );
not \U$5056 ( \5433 , \5432 );
not \U$5057 ( \5434 , \5086 );
or \U$5058 ( \5435 , \5433 , \5434 );
nand \U$5059 ( \5436 , \5073 , \5068 );
nand \U$5060 ( \5437 , \5435 , \5436 );
not \U$5061 ( \5438 , \5437 );
or \U$5062 ( \5439 , \5431 , \5438 );
or \U$5063 ( \5440 , \5437 , \5430 );
not \U$5064 ( \5441 , \2450 );
not \U$5065 ( \5442 , \4003 );
or \U$5066 ( \5443 , \5441 , \5442 );
nand \U$5067 ( \5444 , \5215 , \2545 );
nand \U$5068 ( \5445 , \5443 , \5444 );
not \U$5069 ( \5446 , \1864 );
not \U$5070 ( \5447 , \4085 );
or \U$5071 ( \5448 , \5446 , \5447 );
nand \U$5072 ( \5449 , \5267 , \1910 );
nand \U$5073 ( \5450 , \5448 , \5449 );
xor \U$5074 ( \5451 , \5445 , \5450 );
not \U$5075 ( \5452 , \4344 );
not \U$5076 ( \5453 , \5332 );
or \U$5077 ( \5454 , \5452 , \5453 );
nand \U$5078 ( \5455 , \4067 , \2011 );
nand \U$5079 ( \5456 , \5454 , \5455 );
and \U$5080 ( \5457 , \5451 , \5456 );
and \U$5081 ( \5458 , \5445 , \5450 );
or \U$5082 ( \5459 , \5457 , \5458 );
nand \U$5083 ( \5460 , \5440 , \5459 );
nand \U$5084 ( \5461 , \5439 , \5460 );
not \U$5085 ( \5462 , \5461 );
not \U$5086 ( \5463 , \5462 );
or \U$5087 ( \5464 , \5426 , \5463 );
or \U$5088 ( \5465 , \5425 , \5462 );
nand \U$5089 ( \5466 , \5464 , \5465 );
xor \U$5090 ( \5467 , \5366 , \5466 );
xor \U$5091 ( \5468 , \5394 , \5415 );
xor \U$5092 ( \5469 , \5468 , \5421 );
xor \U$5093 ( \5470 , \5445 , \5450 );
xor \U$5094 ( \5471 , \5470 , \5456 );
not \U$5095 ( \5472 , \5471 );
buf \U$5096 ( \5473 , \5378 );
xor \U$5097 ( \5474 , \5392 , \5473 );
xnor \U$5098 ( \5475 , \5474 , \5389 );
and \U$5099 ( \5476 , \5405 , \5399 );
not \U$5100 ( \5477 , \5405 );
not \U$5101 ( \5478 , \5399 );
and \U$5102 ( \5479 , \5477 , \5478 );
nor \U$5103 ( \5480 , \5476 , \5479 );
not \U$5104 ( \5481 , \5413 );
and \U$5105 ( \5482 , \5480 , \5481 );
not \U$5106 ( \5483 , \5480 );
and \U$5107 ( \5484 , \5483 , \5413 );
nor \U$5108 ( \5485 , \5482 , \5484 );
nand \U$5109 ( \5486 , \5475 , \5485 );
not \U$5110 ( \5487 , \5486 );
or \U$5111 ( \5488 , \5472 , \5487 );
not \U$5112 ( \5489 , \5485 );
not \U$5113 ( \5490 , \5475 );
nand \U$5114 ( \5491 , \5489 , \5490 );
nand \U$5115 ( \5492 , \5488 , \5491 );
nand \U$5116 ( \5493 , \5469 , \5492 );
not \U$5117 ( \5494 , \5493 );
buf \U$5118 ( \5495 , \5459 );
not \U$5119 ( \5496 , \5495 );
not \U$5120 ( \5497 , \5430 );
not \U$5121 ( \5498 , \5497 );
not \U$5122 ( \5499 , \5437 );
or \U$5123 ( \5500 , \5498 , \5499 );
or \U$5124 ( \5501 , \5437 , \5497 );
nand \U$5125 ( \5502 , \5500 , \5501 );
not \U$5126 ( \5503 , \5502 );
or \U$5127 ( \5504 , \5496 , \5503 );
or \U$5128 ( \5505 , \5502 , \5495 );
nand \U$5129 ( \5506 , \5504 , \5505 );
not \U$5130 ( \5507 , \5506 );
or \U$5131 ( \5508 , \5494 , \5507 );
not \U$5132 ( \5509 , \5469 );
not \U$5133 ( \5510 , \5492 );
nand \U$5134 ( \5511 , \5509 , \5510 );
nand \U$5135 ( \5512 , \5508 , \5511 );
not \U$5136 ( \5513 , \5512 );
xor \U$5137 ( \5514 , \5467 , \5513 );
not \U$5138 ( \5515 , \5514 );
nand \U$5139 ( \5516 , \5100 , \5515 );
not \U$5140 ( \5517 , \5145 );
not \U$5141 ( \5518 , \5237 );
or \U$5142 ( \5519 , \5517 , \5518 );
or \U$5143 ( \5520 , \5237 , \5145 );
nand \U$5144 ( \5521 , \5519 , \5520 );
xnor \U$5145 ( \5522 , \5182 , \5521 );
not \U$5146 ( \5523 , \1864 );
not \U$5147 ( \5524 , \5273 );
or \U$5148 ( \5525 , \5523 , \5524 );
and \U$5149 ( \5526 , \3748 , RIae793b8_143);
not \U$5150 ( \5527 , \3748 );
and \U$5151 ( \5528 , \5527 , \1902 );
nor \U$5152 ( \5529 , \5526 , \5528 );
nand \U$5153 ( \5530 , \5529 , \1910 );
nand \U$5154 ( \5531 , \5525 , \5530 );
not \U$5155 ( \5532 , \5531 );
not \U$5156 ( \5533 , \5324 );
not \U$5157 ( \5534 , \5316 );
or \U$5158 ( \5535 , \5533 , \5534 );
not \U$5159 ( \5536 , RIae79c28_161);
not \U$5160 ( \5537 , \2510 );
or \U$5161 ( \5538 , \5536 , \5537 );
or \U$5162 ( \5539 , \2331 , RIae79c28_161);
nand \U$5163 ( \5540 , \5538 , \5539 );
nand \U$5164 ( \5541 , \5540 , \2767 );
nand \U$5165 ( \5542 , \5535 , \5541 );
not \U$5166 ( \5543 , \5542 );
or \U$5167 ( \5544 , \5532 , \5543 );
not \U$5168 ( \5545 , \2322 );
not \U$5169 ( \5546 , \5348 );
or \U$5170 ( \5547 , \5545 , \5546 );
not \U$5171 ( \5548 , \3721 );
and \U$5172 ( \5549 , RIae798e0_154, \5548 );
not \U$5173 ( \5550 , RIae798e0_154);
and \U$5174 ( \5551 , \5550 , \2263 );
nor \U$5175 ( \5552 , \5549 , \5551 );
nand \U$5176 ( \5553 , \5552 , \2341 );
nand \U$5177 ( \5554 , \5547 , \5553 );
not \U$5178 ( \5555 , \5554 );
nand \U$5179 ( \5556 , \5544 , \5555 );
not \U$5180 ( \5557 , \5531 );
not \U$5181 ( \5558 , \5542 );
nand \U$5182 ( \5559 , \5557 , \5558 );
and \U$5183 ( \5560 , \5556 , \5559 );
xor \U$5184 ( \5561 , \5160 , \5167 );
xor \U$5185 ( \5562 , \5561 , \5178 );
xor \U$5186 ( \5563 , \5560 , \5562 );
xor \U$5187 ( \5564 , \5217 , \5202 );
xnor \U$5188 ( \5565 , \5564 , \5233 );
and \U$5189 ( \5566 , \5563 , \5565 );
and \U$5190 ( \5567 , \5560 , \5562 );
or \U$5191 ( \5568 , \5566 , \5567 );
xor \U$5192 ( \5569 , \5522 , \5568 );
xor \U$5193 ( \5570 , \5110 , \5126 );
xor \U$5194 ( \5571 , \5570 , \5142 );
xor \U$5195 ( \5572 , \5326 , \5341 );
xor \U$5196 ( \5573 , \5572 , \5354 );
xor \U$5197 ( \5574 , \5571 , \5573 );
xor \U$5198 ( \5575 , \5017 , \5029 );
xor \U$5199 ( \5576 , \5575 , \5052 );
and \U$5200 ( \5577 , \5574 , \5576 );
and \U$5201 ( \5578 , \5571 , \5573 );
or \U$5202 ( \5579 , \5577 , \5578 );
and \U$5203 ( \5580 , \5569 , \5579 );
and \U$5204 ( \5581 , \5522 , \5568 );
or \U$5205 ( \5582 , \5580 , \5581 );
not \U$5206 ( \5583 , \5582 );
not \U$5207 ( \5584 , \3014 );
not \U$5208 ( \5585 , \5163 );
or \U$5209 ( \5586 , \5584 , \5585 );
not \U$5210 ( \5587 , \2268 );
not \U$5211 ( \5588 , \1899 );
or \U$5212 ( \5589 , \5587 , \5588 );
or \U$5213 ( \5590 , \3294 , \2268 );
nand \U$5214 ( \5591 , \5589 , \5590 );
nand \U$5215 ( \5592 , \5591 , \2272 );
nand \U$5216 ( \5593 , \5586 , \5592 );
not \U$5217 ( \5594 , \2450 );
not \U$5218 ( \5595 , \5208 );
or \U$5219 ( \5596 , \5594 , \5595 );
and \U$5220 ( \5597 , RIae79778_151, \3775 );
not \U$5221 ( \5598 , RIae79778_151);
and \U$5222 ( \5599 , \5598 , \3236 );
or \U$5223 ( \5600 , \5597 , \5599 );
nand \U$5224 ( \5601 , \5600 , \2433 );
nand \U$5225 ( \5602 , \5596 , \5601 );
xor \U$5226 ( \5603 , \5593 , \5602 );
not \U$5227 ( \5604 , \4853 );
not \U$5228 ( \5605 , \5174 );
or \U$5229 ( \5606 , \5604 , \5605 );
and \U$5230 ( \5607 , RIae79ca0_162, \781 );
not \U$5231 ( \5608 , RIae79ca0_162);
and \U$5232 ( \5609 , \5608 , \780 );
nor \U$5233 ( \5610 , \5607 , \5609 );
nand \U$5234 ( \5611 , \5610 , \4842 );
nand \U$5235 ( \5612 , \5606 , \5611 );
and \U$5236 ( \5613 , \5603 , \5612 );
and \U$5237 ( \5614 , \5593 , \5602 );
or \U$5238 ( \5615 , \5613 , \5614 );
not \U$5239 ( \5616 , \5615 );
not \U$5240 ( \5617 , \2007 );
not \U$5241 ( \5618 , \5193 );
or \U$5242 ( \5619 , \5617 , \5618 );
and \U$5243 ( \5620 , \2179 , \1997 );
not \U$5244 ( \5621 , \2179 );
and \U$5245 ( \5622 , \5621 , RIae797f0_152);
nor \U$5246 ( \5623 , \5620 , \5622 );
nand \U$5247 ( \5624 , \5623 , \1989 );
nand \U$5248 ( \5625 , \5619 , \5624 );
not \U$5249 ( \5626 , \2011 );
not \U$5250 ( \5627 , \5339 );
or \U$5251 ( \5628 , \5626 , \5627 );
and \U$5252 ( \5629 , RIae79610_148, \2155 );
not \U$5253 ( \5630 , RIae79610_148);
not \U$5254 ( \5631 , \2153 );
and \U$5255 ( \5632 , \5630 , \5631 );
or \U$5256 ( \5633 , \5629 , \5632 );
nand \U$5257 ( \5634 , \5633 , \4344 );
nand \U$5258 ( \5635 , \5628 , \5634 );
xor \U$5259 ( \5636 , \5625 , \5635 );
not \U$5260 ( \5637 , \3827 );
not \U$5261 ( \5638 , \5224 );
or \U$5262 ( \5639 , \5637 , \5638 );
not \U$5263 ( \5640 , \3244 );
xor \U$5264 ( \5641 , RIae79688_149, \5640 );
nand \U$5265 ( \5642 , \5641 , \2966 );
nand \U$5266 ( \5643 , \5639 , \5642 );
and \U$5267 ( \5644 , \5636 , \5643 );
and \U$5268 ( \5645 , \5625 , \5635 );
or \U$5269 ( \5646 , \5644 , \5645 );
not \U$5270 ( \5647 , \5646 );
or \U$5271 ( \5648 , \5616 , \5647 );
not \U$5272 ( \5649 , \2602 );
not \U$5273 ( \5650 , RIae79520_146);
not \U$5274 ( \5651 , \2047 );
or \U$5275 ( \5652 , \5650 , \5651 );
or \U$5276 ( \5653 , \3141 , RIae79520_146);
nand \U$5277 ( \5654 , \5652 , \5653 );
not \U$5278 ( \5655 , \5654 );
or \U$5279 ( \5656 , \5649 , \5655 );
not \U$5280 ( \5657 , \5139 );
nand \U$5281 ( \5658 , \5657 , \2924 );
nand \U$5282 ( \5659 , \5656 , \5658 );
not \U$5283 ( \5660 , \5659 );
not \U$5284 ( \5661 , \5124 );
not \U$5285 ( \5662 , \5117 );
or \U$5286 ( \5663 , \5661 , \5662 );
and \U$5287 ( \5664 , RIae78f80_134, \1970 );
not \U$5288 ( \5665 , RIae78f80_134);
and \U$5289 ( \5666 , \5665 , \3217 );
or \U$5290 ( \5667 , \5664 , \5666 );
nand \U$5291 ( \5668 , \5667 , \797 );
nand \U$5292 ( \5669 , \5663 , \5668 );
not \U$5293 ( \5670 , \1321 );
not \U$5294 ( \5671 , \5152 );
or \U$5295 ( \5672 , \5670 , \5671 );
not \U$5296 ( \5673 , \2402 );
not \U$5297 ( \5674 , \5673 );
and \U$5298 ( \5675 , \5674 , \1066 );
not \U$5299 ( \5676 , \5674 );
and \U$5300 ( \5677 , \5676 , RIae78e90_132);
nor \U$5301 ( \5678 , \5675 , \5677 );
nand \U$5302 ( \5679 , \5678 , \1086 );
nand \U$5303 ( \5680 , \5672 , \5679 );
xor \U$5304 ( \5681 , \5669 , \5680 );
not \U$5305 ( \5682 , \5681 );
or \U$5306 ( \5683 , \5660 , \5682 );
nand \U$5307 ( \5684 , \5669 , \5680 );
nand \U$5308 ( \5685 , \5683 , \5684 );
not \U$5309 ( \5686 , \5685 );
nand \U$5310 ( \5687 , \5648 , \5686 );
or \U$5311 ( \5688 , \5646 , \5615 );
nand \U$5312 ( \5689 , \5687 , \5688 );
not \U$5313 ( \5690 , \5689 );
not \U$5314 ( \5691 , \5690 );
not \U$5315 ( \5692 , \5290 );
not \U$5316 ( \5693 , \5358 );
or \U$5317 ( \5694 , \5692 , \5693 );
not \U$5318 ( \5695 , \5290 );
nand \U$5319 ( \5696 , \5695 , \5357 );
nand \U$5320 ( \5697 , \5694 , \5696 );
and \U$5321 ( \5698 , \5697 , \5361 );
not \U$5322 ( \5699 , \5697 );
and \U$5323 ( \5700 , \5699 , \5309 );
nor \U$5324 ( \5701 , \5698 , \5700 );
not \U$5325 ( \5702 , \5701 );
not \U$5326 ( \5703 , \5702 );
or \U$5327 ( \5704 , \5691 , \5703 );
not \U$5328 ( \5705 , \5689 );
not \U$5329 ( \5706 , \5701 );
or \U$5330 ( \5707 , \5705 , \5706 );
xor \U$5331 ( \5708 , \4993 , \4991 );
xnor \U$5332 ( \5709 , \5708 , \4977 );
not \U$5333 ( \5710 , \3160 );
not \U$5334 ( \5711 , \5710 );
not \U$5335 ( \5712 , \3183 );
or \U$5336 ( \5713 , \5711 , \5712 );
not \U$5337 ( \5714 , \3193 );
nand \U$5338 ( \5715 , \5713 , \5714 );
nand \U$5339 ( \5716 , \3186 , \586 );
not \U$5340 ( \5717 , \5716 );
and \U$5341 ( \5718 , \5715 , \5717 );
not \U$5342 ( \5719 , \5715 );
and \U$5343 ( \5720 , \5719 , \5716 );
nor \U$5344 ( \5721 , \5718 , \5720 );
buf \U$5345 ( \5722 , \5721 );
and \U$5346 ( \5723 , RIae78b48_125, \5722 );
not \U$5347 ( \5724 , \868 );
not \U$5348 ( \5725 , \4973 );
or \U$5349 ( \5726 , \5724 , \5725 );
xor \U$5350 ( \5727 , RIae78b48_125, \5109 );
nand \U$5351 ( \5728 , \5727 , \893 );
nand \U$5352 ( \5729 , \5726 , \5728 );
or \U$5353 ( \5730 , \5723 , \5729 );
not \U$5354 ( \5731 , \929 );
not \U$5355 ( \5732 , \4983 );
or \U$5356 ( \5733 , \5731 , \5732 );
not \U$5357 ( \5734 , RIae78bc0_126);
not \U$5358 ( \5735 , \4929 );
or \U$5359 ( \5736 , \5734 , \5735 );
nand \U$5360 ( \5737 , \4169 , \1286 );
nand \U$5361 ( \5738 , \5736 , \5737 );
nand \U$5362 ( \5739 , \5738 , \1036 );
nand \U$5363 ( \5740 , \5733 , \5739 );
nand \U$5364 ( \5741 , \5730 , \5740 );
nand \U$5365 ( \5742 , \5729 , \5723 );
nand \U$5366 ( \5743 , \5741 , \5742 );
and \U$5367 ( \5744 , \5709 , \5743 );
not \U$5368 ( \5745 , \5709 );
not \U$5369 ( \5746 , \5743 );
and \U$5370 ( \5747 , \5745 , \5746 );
or \U$5371 ( \5748 , \5744 , \5747 );
not \U$5372 ( \5749 , \5748 );
not \U$5373 ( \5750 , \5749 );
not \U$5374 ( \5751 , \1501 );
not \U$5375 ( \5752 , \5258 );
or \U$5376 ( \5753 , \5751 , \5752 );
and \U$5377 ( \5754 , RIae79250_140, \1755 );
not \U$5378 ( \5755 , RIae79250_140);
and \U$5379 ( \5756 , \5755 , \1760 );
nor \U$5380 ( \5757 , \5754 , \5756 );
nand \U$5381 ( \5758 , \5757 , \2650 );
nand \U$5382 ( \5759 , \5753 , \5758 );
not \U$5383 ( \5760 , \1010 );
not \U$5384 ( \5761 , RIae79160_138);
not \U$5385 ( \5762 , \2577 );
or \U$5386 ( \5763 , \5761 , \5762 );
or \U$5387 ( \5764 , \5020 , RIae79160_138);
nand \U$5388 ( \5765 , \5763 , \5764 );
not \U$5389 ( \5766 , \5765 );
or \U$5390 ( \5767 , \5760 , \5766 );
nand \U$5391 ( \5768 , \5009 , \1013 );
nand \U$5392 ( \5769 , \5767 , \5768 );
xor \U$5393 ( \5770 , \5759 , \5769 );
not \U$5394 ( \5771 , \1919 );
not \U$5395 ( \5772 , \5282 );
or \U$5396 ( \5773 , \5771 , \5772 );
and \U$5397 ( \5774 , RIae794a8_145, \3689 );
not \U$5398 ( \5775 , RIae794a8_145);
and \U$5399 ( \5776 , \5775 , \1405 );
nor \U$5400 ( \5777 , \5774 , \5776 );
nand \U$5401 ( \5778 , \5777 , \1933 );
nand \U$5402 ( \5779 , \5773 , \5778 );
and \U$5403 ( \5780 , \5770 , \5779 );
and \U$5404 ( \5781 , \5759 , \5769 );
or \U$5405 ( \5782 , \5780 , \5781 );
not \U$5406 ( \5783 , \5782 );
not \U$5407 ( \5784 , \5783 );
and \U$5408 ( \5785 , \5750 , \5784 );
not \U$5409 ( \5786 , \5709 );
and \U$5410 ( \5787 , \5786 , \5743 );
nor \U$5411 ( \5788 , \5785 , \5787 );
not \U$5412 ( \5789 , \5788 );
nand \U$5413 ( \5790 , \5707 , \5789 );
nand \U$5414 ( \5791 , \5704 , \5790 );
not \U$5415 ( \5792 , \5791 );
or \U$5416 ( \5793 , \5583 , \5792 );
or \U$5417 ( \5794 , \5791 , \5582 );
xor \U$5418 ( \5795 , \5239 , \5363 );
xnor \U$5419 ( \5796 , \5795 , \5246 );
nand \U$5420 ( \5797 , \5794 , \5796 );
nand \U$5421 ( \5798 , \5793 , \5797 );
and \U$5422 ( \5799 , \5516 , \5798 );
nor \U$5423 ( \5800 , \5100 , \5515 );
nor \U$5424 ( \5801 , \5799 , \5800 );
xor \U$5425 ( \5802 , \4879 , \5801 );
xor \U$5426 ( \5803 , \5366 , \5466 );
and \U$5427 ( \5804 , \5803 , \5513 );
and \U$5428 ( \5805 , \5366 , \5466 );
or \U$5429 ( \5806 , \5804 , \5805 );
xor \U$5430 ( \5807 , \4884 , \4903 );
and \U$5431 ( \5808 , \5807 , \4906 );
and \U$5432 ( \5809 , \4884 , \4903 );
or \U$5433 ( \5810 , \5808 , \5809 );
not \U$5434 ( \5811 , \5810 );
and \U$5435 ( \5812 , \5425 , \5461 );
and \U$5436 ( \5813 , \5373 , \5424 );
nor \U$5437 ( \5814 , \5812 , \5813 );
not \U$5438 ( \5815 , \5814 );
not \U$5439 ( \5816 , \4095 );
not \U$5440 ( \5817 , \5816 );
not \U$5441 ( \5818 , \4233 );
or \U$5442 ( \5819 , \5817 , \5818 );
not \U$5443 ( \5820 , \4233 );
nand \U$5444 ( \5821 , \5820 , \4095 );
nand \U$5445 ( \5822 , \5819 , \5821 );
not \U$5446 ( \5823 , \5822 );
or \U$5447 ( \5824 , \5815 , \5823 );
or \U$5448 ( \5825 , \5822 , \5814 );
nand \U$5449 ( \5826 , \5824 , \5825 );
not \U$5450 ( \5827 , \5826 );
not \U$5451 ( \5828 , \5827 );
or \U$5452 ( \5829 , \5811 , \5828 );
not \U$5453 ( \5830 , \5810 );
nand \U$5454 ( \5831 , \5830 , \5826 );
nand \U$5455 ( \5832 , \5829 , \5831 );
xor \U$5456 ( \5833 , \5806 , \5832 );
not \U$5457 ( \5834 , \4907 );
nand \U$5458 ( \5835 , \5834 , \5097 );
not \U$5459 ( \5836 , \5835 );
not \U$5460 ( \5837 , \5099 );
or \U$5461 ( \5838 , \5836 , \5837 );
not \U$5462 ( \5839 , \5097 );
nand \U$5463 ( \5840 , \5839 , \4907 );
nand \U$5464 ( \5841 , \5838 , \5840 );
xnor \U$5465 ( \5842 , \5833 , \5841 );
xor \U$5466 ( \5843 , \5802 , \5842 );
and \U$5467 ( \5844 , \5092 , \4918 );
not \U$5468 ( \5845 , \5092 );
and \U$5469 ( \5846 , \5845 , \5095 );
nor \U$5470 ( \5847 , \5844 , \5846 );
xnor \U$5471 ( \5848 , \4909 , \5847 );
not \U$5472 ( \5849 , \5848 );
nand \U$5473 ( \5850 , \5491 , \5486 );
not \U$5474 ( \5851 , \5471 );
and \U$5475 ( \5852 , \5850 , \5851 );
not \U$5476 ( \5853 , \5850 );
and \U$5477 ( \5854 , \5853 , \5471 );
nor \U$5478 ( \5855 , \5852 , \5854 );
xor \U$5479 ( \5856 , \5262 , \5275 );
xor \U$5480 ( \5857 , \5856 , \5287 );
buf \U$5481 ( \5858 , \1086 );
not \U$5482 ( \5859 , \5858 );
not \U$5483 ( \5860 , \3207 );
not \U$5484 ( \5861 , \5860 );
xor \U$5485 ( \5862 , RIae78e90_132, \5861 );
not \U$5486 ( \5863 , \5862 );
or \U$5487 ( \5864 , \5859 , \5863 );
nand \U$5488 ( \5865 , \5678 , \1321 );
nand \U$5489 ( \5866 , \5864 , \5865 );
not \U$5490 ( \5867 , RIae79fe8_169);
not \U$5491 ( \5868 , RIae79f70_168);
or \U$5492 ( \5869 , \5867 , \5868 );
nand \U$5493 ( \5870 , \5869 , RIae79ef8_167);
or \U$5494 ( \5871 , \5866 , \5870 );
not \U$5495 ( \5872 , \952 );
and \U$5496 ( \5873 , \4960 , \1286 );
not \U$5497 ( \5874 , \4960 );
and \U$5498 ( \5875 , \5874 , RIae78bc0_126);
nor \U$5499 ( \5876 , \5873 , \5875 );
not \U$5500 ( \5877 , \5876 );
or \U$5501 ( \5878 , \5872 , \5877 );
nand \U$5502 ( \5879 , \5738 , \927 );
nand \U$5503 ( \5880 , \5878 , \5879 );
nand \U$5504 ( \5881 , \5871 , \5880 );
nand \U$5505 ( \5882 , \5866 , \5870 );
nand \U$5506 ( \5883 , \5881 , \5882 );
not \U$5507 ( \5884 , \5883 );
not \U$5508 ( \5885 , \1049 );
not \U$5509 ( \5886 , \5027 );
or \U$5510 ( \5887 , \5885 , \5886 );
and \U$5511 ( \5888 , RIae79070_136, \2090 );
not \U$5512 ( \5889 , RIae79070_136);
not \U$5513 ( \5890 , \2088 );
not \U$5514 ( \5891 , \5890 );
and \U$5515 ( \5892 , \5889 , \5891 );
or \U$5516 ( \5893 , \5888 , \5892 );
nand \U$5517 ( \5894 , \5893 , \1062 );
nand \U$5518 ( \5895 , \5887 , \5894 );
not \U$5519 ( \5896 , \5895 );
not \U$5520 ( \5897 , \5051 );
or \U$5521 ( \5898 , \5896 , \5897 );
or \U$5522 ( \5899 , \5051 , \5895 );
nand \U$5523 ( \5900 , \5898 , \5899 );
not \U$5524 ( \5901 , \5900 );
or \U$5525 ( \5902 , \5884 , \5901 );
not \U$5526 ( \5903 , \5052 );
nand \U$5527 ( \5904 , \5903 , \5895 );
nand \U$5528 ( \5905 , \5902 , \5904 );
xor \U$5529 ( \5906 , \5857 , \5905 );
not \U$5530 ( \5907 , \5906 );
not \U$5531 ( \5908 , \1062 );
and \U$5532 ( \5909 , RIae79070_136, \4113 );
not \U$5533 ( \5910 , RIae79070_136);
buf \U$5534 ( \5911 , \1953 );
buf \U$5535 ( \5912 , \5911 );
and \U$5536 ( \5913 , \5910 , \5912 );
or \U$5537 ( \5914 , \5909 , \5913 );
not \U$5538 ( \5915 , \5914 );
or \U$5539 ( \5916 , \5908 , \5915 );
nand \U$5540 ( \5917 , \5893 , \1049 );
nand \U$5541 ( \5918 , \5916 , \5917 );
not \U$5542 ( \5919 , \839 );
not \U$5543 ( \5920 , \5667 );
or \U$5544 ( \5921 , \5919 , \5920 );
and \U$5545 ( \5922 , RIae78f80_134, \2385 );
not \U$5546 ( \5923 , RIae78f80_134);
and \U$5547 ( \5924 , \5923 , \1859 );
nor \U$5548 ( \5925 , \5922 , \5924 );
nand \U$5549 ( \5926 , \5925 , \797 );
nand \U$5550 ( \5927 , \5921 , \5926 );
or \U$5551 ( \5928 , \5918 , \5927 );
not \U$5552 ( \5929 , \5928 );
not \U$5553 ( \5930 , \5040 );
xor \U$5554 ( \5931 , RIae79d90_164, \2004 );
not \U$5555 ( \5932 , \5931 );
or \U$5556 ( \5933 , \5930 , \5932 );
nand \U$5557 ( \5934 , \5045 , \5049 );
nand \U$5558 ( \5935 , \5933 , \5934 );
not \U$5559 ( \5936 , \5935 );
or \U$5560 ( \5937 , \5929 , \5936 );
nand \U$5561 ( \5938 , \5918 , \5927 );
nand \U$5562 ( \5939 , \5937 , \5938 );
not \U$5563 ( \5940 , \3440 );
not \U$5564 ( \5941 , \5654 );
or \U$5565 ( \5942 , \5940 , \5941 );
not \U$5566 ( \5943 , RIae79520_146);
not \U$5567 ( \5944 , \4197 );
not \U$5568 ( \5945 , \5944 );
not \U$5569 ( \5946 , \5945 );
or \U$5570 ( \5947 , \5943 , \5946 );
or \U$5571 ( \5948 , \4199 , RIae79520_146);
nand \U$5572 ( \5949 , \5947 , \5948 );
buf \U$5573 ( \5950 , \2602 );
nand \U$5574 ( \5951 , \5949 , \5950 );
nand \U$5575 ( \5952 , \5942 , \5951 );
not \U$5576 ( \5953 , \2767 );
not \U$5577 ( \5954 , RIae79c28_161);
not \U$5578 ( \5955 , \1439 );
or \U$5579 ( \5956 , \5954 , \5955 );
not \U$5580 ( \5957 , \1438 );
not \U$5581 ( \5958 , \5957 );
or \U$5582 ( \5959 , \5958 , RIae79c28_161);
nand \U$5583 ( \5960 , \5956 , \5959 );
not \U$5584 ( \5961 , \5960 );
or \U$5585 ( \5962 , \5953 , \5961 );
nand \U$5586 ( \5963 , \5540 , \2776 );
nand \U$5587 ( \5964 , \5962 , \5963 );
xor \U$5588 ( \5965 , \5952 , \5964 );
not \U$5589 ( \5966 , \2252 );
not \U$5590 ( \5967 , \5591 );
or \U$5591 ( \5968 , \5966 , \5967 );
and \U$5592 ( \5969 , RIae79ac0_158, \2208 );
not \U$5593 ( \5970 , RIae79ac0_158);
not \U$5594 ( \5971 , \2629 );
and \U$5595 ( \5972 , \5970 , \5971 );
or \U$5596 ( \5973 , \5969 , \5972 );
not \U$5597 ( \5974 , \5973 );
or \U$5598 ( \5975 , \5974 , \3510 );
nand \U$5599 ( \5976 , \5968 , \5975 );
and \U$5600 ( \5977 , \5965 , \5976 );
and \U$5601 ( \5978 , \5952 , \5964 );
or \U$5602 ( \5979 , \5977 , \5978 );
xor \U$5603 ( \5980 , \5939 , \5979 );
not \U$5604 ( \5981 , \3827 );
not \U$5605 ( \5982 , \5641 );
or \U$5606 ( \5983 , \5981 , \5982 );
not \U$5607 ( \5984 , \2970 );
not \U$5608 ( \5985 , \2141 );
not \U$5609 ( \5986 , \5985 );
or \U$5610 ( \5987 , \5984 , \5986 );
nand \U$5611 ( \5988 , \3071 , RIae79688_149);
nand \U$5612 ( \5989 , \5987 , \5988 );
nand \U$5613 ( \5990 , \5989 , \2966 );
nand \U$5614 ( \5991 , \5983 , \5990 );
not \U$5615 ( \5992 , \4842 );
and \U$5616 ( \5993 , RIae79ca0_162, \2640 );
not \U$5617 ( \5994 , RIae79ca0_162);
and \U$5618 ( \5995 , \5994 , \3999 );
nor \U$5619 ( \5996 , \5993 , \5995 );
not \U$5620 ( \5997 , \5996 );
or \U$5621 ( \5998 , \5992 , \5997 );
nand \U$5622 ( \5999 , \5610 , \4853 );
nand \U$5623 ( \6000 , \5998 , \5999 );
nor \U$5624 ( \6001 , \5991 , \6000 );
not \U$5625 ( \6002 , \2442 );
not \U$5626 ( \6003 , \5191 );
or \U$5627 ( \6004 , \6002 , \6003 );
nand \U$5628 ( \6005 , \2169 , RIae79778_151);
nand \U$5629 ( \6006 , \6004 , \6005 );
and \U$5630 ( \6007 , \2545 , \6006 );
and \U$5631 ( \6008 , \5600 , \2450 );
nor \U$5632 ( \6009 , \6007 , \6008 );
or \U$5633 ( \6010 , \6001 , \6009 );
nand \U$5634 ( \6011 , \5991 , \6000 );
nand \U$5635 ( \6012 , \6010 , \6011 );
and \U$5636 ( \6013 , \5980 , \6012 );
and \U$5637 ( \6014 , \5939 , \5979 );
or \U$5638 ( \6015 , \6013 , \6014 );
not \U$5639 ( \6016 , \6015 );
or \U$5640 ( \6017 , \5907 , \6016 );
nand \U$5641 ( \6018 , \5905 , \5857 );
nand \U$5642 ( \6019 , \6017 , \6018 );
xor \U$5643 ( \6020 , \5855 , \6019 );
xor \U$5644 ( \6021 , \5057 , \5088 );
xnor \U$5645 ( \6022 , \6021 , \5004 );
and \U$5646 ( \6023 , \6020 , \6022 );
and \U$5647 ( \6024 , \5855 , \6019 );
or \U$5648 ( \6025 , \6023 , \6024 );
not \U$5649 ( \6026 , \6025 );
or \U$5650 ( \6027 , \5849 , \6026 );
or \U$5651 ( \6028 , \6025 , \5848 );
nand \U$5652 ( \6029 , \5493 , \5511 );
not \U$5653 ( \6030 , \5506 );
and \U$5654 ( \6031 , \6029 , \6030 );
not \U$5655 ( \6032 , \6029 );
and \U$5656 ( \6033 , \6032 , \5506 );
nor \U$5657 ( \6034 , \6031 , \6033 );
not \U$5658 ( \6035 , \6034 );
nand \U$5659 ( \6036 , \6028 , \6035 );
nand \U$5660 ( \6037 , \6027 , \6036 );
not \U$5661 ( \6038 , \6037 );
not \U$5662 ( \6039 , \5798 );
not \U$5663 ( \6040 , \5515 );
or \U$5664 ( \6041 , \6039 , \6040 );
not \U$5665 ( \6042 , \5798 );
nand \U$5666 ( \6043 , \5514 , \6042 );
nand \U$5667 ( \6044 , \6041 , \6043 );
buf \U$5668 ( \6045 , \5100 );
not \U$5669 ( \6046 , \6045 );
and \U$5670 ( \6047 , \6044 , \6046 );
not \U$5671 ( \6048 , \6044 );
and \U$5672 ( \6049 , \6048 , \6045 );
nor \U$5673 ( \6050 , \6047 , \6049 );
not \U$5674 ( \6051 , \6050 );
or \U$5675 ( \6052 , \6038 , \6051 );
or \U$5676 ( \6053 , \6050 , \6037 );
xor \U$5677 ( \6054 , \5522 , \5568 );
xor \U$5678 ( \6055 , \6054 , \5579 );
xor \U$5679 ( \6056 , \5906 , \6015 );
xor \U$5680 ( \6057 , \5571 , \5573 );
xor \U$5681 ( \6058 , \6057 , \5576 );
xor \U$5682 ( \6059 , \6056 , \6058 );
buf \U$5683 ( \6060 , \5900 );
xor \U$5684 ( \6061 , \5883 , \6060 );
not \U$5685 ( \6062 , \6061 );
not \U$5686 ( \6063 , \839 );
not \U$5687 ( \6064 , \5925 );
or \U$5688 ( \6065 , \6063 , \6064 );
xnor \U$5689 ( \6066 , \3270 , RIae78f80_134);
nand \U$5690 ( \6067 , \797 , \6066 );
nand \U$5691 ( \6068 , \6065 , \6067 );
not \U$5692 ( \6069 , \2610 );
not \U$5693 ( \6070 , \5949 );
or \U$5694 ( \6071 , \6069 , \6070 );
not \U$5695 ( \6072 , \4653 );
not \U$5696 ( \6073 , \1899 );
or \U$5697 ( \6074 , \6072 , \6073 );
or \U$5698 ( \6075 , \3294 , \4653 );
nand \U$5699 ( \6076 , \6074 , \6075 );
nand \U$5700 ( \6077 , \6076 , \2602 );
nand \U$5701 ( \6078 , \6071 , \6077 );
xor \U$5702 ( \6079 , \6068 , \6078 );
buf \U$5703 ( \6080 , \5048 );
not \U$5704 ( \6081 , \6080 );
not \U$5705 ( \6082 , \5931 );
or \U$5706 ( \6083 , \6081 , \6082 );
not \U$5707 ( \6084 , RIae79d90_164);
not \U$5708 ( \6085 , \6084 );
not \U$5709 ( \6086 , \780 );
not \U$5710 ( \6087 , \6086 );
or \U$5711 ( \6088 , \6085 , \6087 );
or \U$5712 ( \6089 , \1994 , \4968 );
nand \U$5713 ( \6090 , \6088 , \6089 );
buf \U$5714 ( \6091 , \5039 );
nand \U$5715 ( \6092 , \6090 , \6091 );
nand \U$5716 ( \6093 , \6083 , \6092 );
and \U$5717 ( \6094 , \6079 , \6093 );
and \U$5718 ( \6095 , \6068 , \6078 );
or \U$5719 ( \6096 , \6094 , \6095 );
not \U$5720 ( \6097 , \6096 );
not \U$5721 ( \6098 , \2450 );
not \U$5722 ( \6099 , \6006 );
or \U$5723 ( \6100 , \6098 , \6099 );
not \U$5724 ( \6101 , \5351 );
not \U$5725 ( \6102 , \2447 );
and \U$5726 ( \6103 , \6101 , \6102 );
not \U$5727 ( \6104 , \878 );
and \U$5728 ( \6105 , \6104 , \2447 );
nor \U$5729 ( \6106 , \6103 , \6105 );
not \U$5730 ( \6107 , \6106 );
nand \U$5731 ( \6108 , \6107 , \2545 );
nand \U$5732 ( \6109 , \6100 , \6108 );
not \U$5733 ( \6110 , \6109 );
not \U$5734 ( \6111 , \5324 );
not \U$5735 ( \6112 , \5960 );
or \U$5736 ( \6113 , \6111 , \6112 );
xor \U$5737 ( \6114 , \3236 , RIae79c28_161);
nand \U$5738 ( \6115 , \6114 , \2767 );
nand \U$5739 ( \6116 , \6113 , \6115 );
not \U$5740 ( \6117 , \6116 );
not \U$5741 ( \6118 , \6117 );
not \U$5742 ( \6119 , \2272 );
and \U$5743 ( \6120 , RIae79ac0_158, \3244 );
not \U$5744 ( \6121 , RIae79ac0_158);
and \U$5745 ( \6122 , \6121 , \2231 );
or \U$5746 ( \6123 , \6120 , \6122 );
not \U$5747 ( \6124 , \6123 );
or \U$5748 ( \6125 , \6119 , \6124 );
nand \U$5749 ( \6126 , \5973 , \3014 );
nand \U$5750 ( \6127 , \6125 , \6126 );
not \U$5751 ( \6128 , \6127 );
or \U$5752 ( \6129 , \6118 , \6128 );
or \U$5753 ( \6130 , \6127 , \6117 );
nand \U$5754 ( \6131 , \6129 , \6130 );
not \U$5755 ( \6132 , \6131 );
or \U$5756 ( \6133 , \6110 , \6132 );
nand \U$5757 ( \6134 , \6127 , \6116 );
nand \U$5758 ( \6135 , \6133 , \6134 );
not \U$5759 ( \6136 , \6135 );
or \U$5760 ( \6137 , \6097 , \6136 );
or \U$5761 ( \6138 , \6135 , \6096 );
not \U$5762 ( \6139 , \2322 );
not \U$5763 ( \6140 , RIae798e0_154);
not \U$5764 ( \6141 , \1186 );
or \U$5765 ( \6142 , \6140 , \6141 );
or \U$5766 ( \6143 , \1187 , RIae798e0_154);
nand \U$5767 ( \6144 , \6142 , \6143 );
not \U$5768 ( \6145 , \6144 );
or \U$5769 ( \6146 , \6139 , \6145 );
buf \U$5770 ( \6147 , \2847 );
not \U$5771 ( \6148 , \6147 );
and \U$5772 ( \6149 , RIae798e0_154, \6148 );
not \U$5773 ( \6150 , RIae798e0_154);
and \U$5774 ( \6151 , \6150 , \1405 );
nor \U$5775 ( \6152 , \6149 , \6151 );
nand \U$5776 ( \6153 , \6152 , \2341 );
nand \U$5777 ( \6154 , \6146 , \6153 );
not \U$5778 ( \6155 , \2063 );
and \U$5779 ( \6156 , RIae79610_148, \2287 );
not \U$5780 ( \6157 , RIae79610_148);
and \U$5781 ( \6158 , \6157 , \3748 );
or \U$5782 ( \6159 , \6156 , \6158 );
not \U$5783 ( \6160 , \6159 );
or \U$5784 ( \6161 , \6155 , \6160 );
and \U$5785 ( \6162 , \2309 , RIae79610_148);
not \U$5786 ( \6163 , \2309 );
and \U$5787 ( \6164 , \6163 , \2053 );
nor \U$5788 ( \6165 , \6162 , \6164 );
nand \U$5789 ( \6166 , \6165 , \2011 );
nand \U$5790 ( \6167 , \6161 , \6166 );
nor \U$5791 ( \6168 , \6154 , \6167 );
and \U$5792 ( \6169 , RIae793b8_143, \1741 );
not \U$5793 ( \6170 , RIae793b8_143);
not \U$5794 ( \6171 , \1739 );
and \U$5795 ( \6172 , \6170 , \6171 );
or \U$5796 ( \6173 , \6169 , \6172 );
and \U$5797 ( \6174 , \1864 , \6173 );
and \U$5798 ( \6175 , RIae793b8_143, \1759 );
not \U$5799 ( \6176 , RIae793b8_143);
and \U$5800 ( \6177 , \6176 , \1760 );
nor \U$5801 ( \6178 , \6175 , \6177 );
and \U$5802 ( \6179 , \6178 , \1910 );
nor \U$5803 ( \6180 , \6174 , \6179 );
or \U$5804 ( \6181 , \6168 , \6180 );
nand \U$5805 ( \6182 , \6154 , \6167 );
nand \U$5806 ( \6183 , \6181 , \6182 );
nand \U$5807 ( \6184 , \6138 , \6183 );
nand \U$5808 ( \6185 , \6137 , \6184 );
not \U$5809 ( \6186 , \6185 );
or \U$5810 ( \6187 , \6062 , \6186 );
or \U$5811 ( \6188 , \6185 , \6061 );
not \U$5812 ( \6189 , RIae79f70_168);
and \U$5813 ( \6190 , RIae79fe8_169, \6189 );
not \U$5814 ( \6191 , RIae79fe8_169);
and \U$5815 ( \6192 , \6191 , RIae79f70_168);
nor \U$5816 ( \6193 , \6190 , \6192 );
and \U$5817 ( \6194 , RIae79ef8_167, RIae79f70_168);
not \U$5818 ( \6195 , RIae79ef8_167);
and \U$5819 ( \6196 , \6195 , \6189 );
nor \U$5820 ( \6197 , \6194 , \6196 );
nand \U$5821 ( \6198 , \6193 , \6197 );
not \U$5822 ( \6199 , \6198 );
buf \U$5823 ( \6200 , \6199 );
buf \U$5824 ( \6201 , \6200 );
not \U$5825 ( \6202 , \6201 );
not \U$5826 ( \6203 , RIae79ef8_167);
not \U$5827 ( \6204 , \6203 );
not \U$5828 ( \6205 , \992 );
or \U$5829 ( \6206 , \6204 , \6205 );
not \U$5830 ( \6207 , RIae79ef8_167);
or \U$5831 ( \6208 , \992 , \6207 );
nand \U$5832 ( \6209 , \6206 , \6208 );
not \U$5833 ( \6210 , \6209 );
or \U$5834 ( \6211 , \6202 , \6210 );
not \U$5835 ( \6212 , \6193 );
not \U$5836 ( \6213 , \6212 );
not \U$5837 ( \6214 , \6213 );
nand \U$5838 ( \6215 , \6214 , RIae79ef8_167);
nand \U$5839 ( \6216 , \6211 , \6215 );
buf \U$5840 ( \6217 , \482 );
not \U$5841 ( \6218 , \6217 );
not \U$5842 ( \6219 , \3183 );
or \U$5843 ( \6220 , \6218 , \6219 );
nand \U$5844 ( \6221 , \6220 , \589 );
not \U$5845 ( \6222 , \6221 );
buf \U$5846 ( \6223 , \479 );
nand \U$5847 ( \6224 , \6223 , \591 );
not \U$5848 ( \6225 , \6224 );
and \U$5849 ( \6226 , \6222 , \6225 );
and \U$5850 ( \6227 , \6221 , \6224 );
nor \U$5851 ( \6228 , \6226 , \6227 );
not \U$5852 ( \6229 , \6228 );
buf \U$5853 ( \6230 , \6229 );
not \U$5854 ( \6231 , \6230 );
not \U$5855 ( \6232 , \6231 );
and \U$5856 ( \6233 , RIae78b48_125, \6232 );
not \U$5857 ( \6234 , \6233 );
not \U$5858 ( \6235 , \1074 );
not \U$5859 ( \6236 , \5862 );
or \U$5860 ( \6237 , \6235 , \6236 );
buf \U$5861 ( \6238 , \4926 );
not \U$5862 ( \6239 , \6238 );
not \U$5863 ( \6240 , RIae78e90_132);
and \U$5864 ( \6241 , \6239 , \6240 );
buf \U$5865 ( \6242 , \4926 );
not \U$5866 ( \6243 , \6242 );
not \U$5867 ( \6244 , \6243 );
and \U$5868 ( \6245 , \6244 , RIae78e90_132);
nor \U$5869 ( \6246 , \6241 , \6245 );
not \U$5870 ( \6247 , \6246 );
nand \U$5871 ( \6248 , \6247 , \5858 );
nand \U$5872 ( \6249 , \6237 , \6248 );
not \U$5873 ( \6250 , \6249 );
or \U$5874 ( \6251 , \6234 , \6250 );
or \U$5875 ( \6252 , \6249 , \6233 );
not \U$5876 ( \6253 , \1027 );
not \U$5877 ( \6254 , \5876 );
or \U$5878 ( \6255 , \6253 , \6254 );
buf \U$5879 ( \6256 , \5106 );
not \U$5880 ( \6257 , \6256 );
and \U$5881 ( \6258 , RIae78bc0_126, \6257 );
not \U$5882 ( \6259 , RIae78bc0_126);
and \U$5883 ( \6260 , \6259 , \6256 );
or \U$5884 ( \6261 , \6258 , \6260 );
nand \U$5885 ( \6262 , \6261 , \1036 );
nand \U$5886 ( \6263 , \6255 , \6262 );
nand \U$5887 ( \6264 , \6252 , \6263 );
nand \U$5888 ( \6265 , \6251 , \6264 );
xor \U$5889 ( \6266 , \6216 , \6265 );
not \U$5890 ( \6267 , \4853 );
not \U$5891 ( \6268 , \5996 );
or \U$5892 ( \6269 , \6267 , \6268 );
not \U$5893 ( \6270 , RIae79ca0_162);
not \U$5894 ( \6271 , \6270 );
not \U$5895 ( \6272 , \1289 );
or \U$5896 ( \6273 , \6271 , \6272 );
nand \U$5897 ( \6274 , \3326 , RIae79ca0_162);
nand \U$5898 ( \6275 , \6273 , \6274 );
buf \U$5899 ( \6276 , \4154 );
nand \U$5900 ( \6277 , \6275 , \6276 );
nand \U$5901 ( \6278 , \6269 , \6277 );
not \U$5902 ( \6279 , \3827 );
not \U$5903 ( \6280 , \5989 );
or \U$5904 ( \6281 , \6279 , \6280 );
and \U$5905 ( \6282 , RIae79688_149, \5631 );
not \U$5906 ( \6283 , RIae79688_149);
and \U$5907 ( \6284 , \6283 , \2155 );
nor \U$5908 ( \6285 , \6282 , \6284 );
nand \U$5909 ( \6286 , \6285 , \1844 );
nand \U$5910 ( \6287 , \6281 , \6286 );
xor \U$5911 ( \6288 , \6278 , \6287 );
not \U$5912 ( \6289 , \2007 );
not \U$5913 ( \6290 , RIae797f0_152);
not \U$5914 ( \6291 , \1472 );
or \U$5915 ( \6292 , \6290 , \6291 );
or \U$5916 ( \6293 , \2918 , RIae797f0_152);
nand \U$5917 ( \6294 , \6292 , \6293 );
not \U$5918 ( \6295 , \6294 );
or \U$5919 ( \6296 , \6289 , \6295 );
not \U$5920 ( \6297 , RIae797f0_152);
not \U$5921 ( \6298 , \2263 );
or \U$5922 ( \6299 , \6297 , \6298 );
or \U$5923 ( \6300 , \3721 , RIae797f0_152);
nand \U$5924 ( \6301 , \6299 , \6300 );
nand \U$5925 ( \6302 , \6301 , \1989 );
nand \U$5926 ( \6303 , \6296 , \6302 );
and \U$5927 ( \6304 , \6288 , \6303 );
and \U$5928 ( \6305 , \6278 , \6287 );
or \U$5929 ( \6306 , \6304 , \6305 );
and \U$5930 ( \6307 , \6266 , \6306 );
and \U$5931 ( \6308 , \6216 , \6265 );
or \U$5932 ( \6309 , \6307 , \6308 );
nand \U$5933 ( \6310 , \6188 , \6309 );
nand \U$5934 ( \6311 , \6187 , \6310 );
and \U$5935 ( \6312 , \6059 , \6311 );
and \U$5936 ( \6313 , \6056 , \6058 );
or \U$5937 ( \6314 , \6312 , \6313 );
xor \U$5938 ( \6315 , \6055 , \6314 );
xor \U$5939 ( \6316 , \5855 , \6019 );
xor \U$5940 ( \6317 , \6316 , \6022 );
and \U$5941 ( \6318 , \6315 , \6317 );
and \U$5942 ( \6319 , \6055 , \6314 );
or \U$5943 ( \6320 , \6318 , \6319 );
xor \U$5944 ( \6321 , \5560 , \5562 );
xor \U$5945 ( \6322 , \6321 , \5565 );
and \U$5946 ( \6323 , \5748 , \5782 );
not \U$5947 ( \6324 , \5748 );
and \U$5948 ( \6325 , \6324 , \5783 );
nor \U$5949 ( \6326 , \6323 , \6325 );
or \U$5950 ( \6327 , \6322 , \6326 );
xor \U$5951 ( \6328 , \5685 , \5615 );
xor \U$5952 ( \6329 , \6328 , \5646 );
nand \U$5953 ( \6330 , \6327 , \6329 );
nand \U$5954 ( \6331 , \6322 , \6326 );
nand \U$5955 ( \6332 , \6330 , \6331 );
and \U$5956 ( \6333 , \6217 , \6223 );
not \U$5957 ( \6334 , \6333 );
not \U$5958 ( \6335 , \3183 );
or \U$5959 ( \6336 , \6334 , \6335 );
not \U$5960 ( \6337 , \3190 );
nand \U$5961 ( \6338 , \6336 , \6337 );
nand \U$5962 ( \6339 , \3188 , \585 );
not \U$5963 ( \6340 , \6339 );
and \U$5964 ( \6341 , \6338 , \6340 );
not \U$5965 ( \6342 , \6338 );
and \U$5966 ( \6343 , \6342 , \6339 );
nor \U$5967 ( \6344 , \6341 , \6343 );
buf \U$5968 ( \6345 , \6344 );
not \U$5969 ( \6346 , \6345 );
not \U$5970 ( \6347 , \6346 );
nand \U$5971 ( \6348 , \6347 , RIae78b48_125);
and \U$5972 ( \6349 , \868 , \5727 );
xor \U$5973 ( \6350 , RIae78b48_125, \5722 );
and \U$5974 ( \6351 , \6350 , \893 );
nor \U$5975 ( \6352 , \6349 , \6351 );
xor \U$5976 ( \6353 , \6348 , \6352 );
not \U$5977 ( \6354 , \5285 );
not \U$5978 ( \6355 , \5777 );
or \U$5979 ( \6356 , \6354 , \6355 );
and \U$5980 ( \6357 , RIae794a8_145, \2026 );
not \U$5981 ( \6358 , RIae794a8_145);
not \U$5982 ( \6359 , \5134 );
and \U$5983 ( \6360 , \6358 , \6359 );
or \U$5984 ( \6361 , \6357 , \6360 );
nand \U$5985 ( \6362 , \6361 , \1933 );
nand \U$5986 ( \6363 , \6356 , \6362 );
not \U$5987 ( \6364 , \6363 );
and \U$5988 ( \6365 , \6353 , \6364 );
and \U$5989 ( \6366 , \6348 , \6352 );
nor \U$5990 ( \6367 , \6365 , \6366 );
not \U$5991 ( \6368 , \6367 );
not \U$5992 ( \6369 , \1910 );
not \U$5993 ( \6370 , \6173 );
or \U$5994 ( \6371 , \6369 , \6370 );
nand \U$5995 ( \6372 , \5529 , \1864 );
nand \U$5996 ( \6373 , \6371 , \6372 );
not \U$5997 ( \6374 , \2011 );
not \U$5998 ( \6375 , \5633 );
or \U$5999 ( \6376 , \6374 , \6375 );
nand \U$6000 ( \6377 , \6165 , \2063 );
nand \U$6001 ( \6378 , \6376 , \6377 );
xor \U$6002 ( \6379 , \6373 , \6378 );
not \U$6003 ( \6380 , \2529 );
not \U$6004 ( \6381 , \6294 );
or \U$6005 ( \6382 , \6380 , \6381 );
nand \U$6006 ( \6383 , \5623 , \2007 );
nand \U$6007 ( \6384 , \6382 , \6383 );
and \U$6008 ( \6385 , \6379 , \6384 );
and \U$6009 ( \6386 , \6373 , \6378 );
or \U$6010 ( \6387 , \6385 , \6386 );
not \U$6011 ( \6388 , \6387 );
or \U$6012 ( \6389 , \6368 , \6388 );
xor \U$6013 ( \6390 , \5723 , \5729 );
xnor \U$6014 ( \6391 , \6390 , \5740 );
nand \U$6015 ( \6392 , \6389 , \6391 );
not \U$6016 ( \6393 , \6387 );
not \U$6017 ( \6394 , \6367 );
nand \U$6018 ( \6395 , \6393 , \6394 );
and \U$6019 ( \6396 , \6392 , \6395 );
not \U$6020 ( \6397 , \1499 );
not \U$6021 ( \6398 , \2697 );
and \U$6022 ( \6399 , RIae79250_140, \6398 );
not \U$6023 ( \6400 , RIae79250_140);
and \U$6024 ( \6401 , \6400 , \3525 );
nor \U$6025 ( \6402 , \6399 , \6401 );
not \U$6026 ( \6403 , \6402 );
or \U$6027 ( \6404 , \6397 , \6403 );
nand \U$6028 ( \6405 , \5757 , \1501 );
nand \U$6029 ( \6406 , \6404 , \6405 );
not \U$6030 ( \6407 , \1209 );
not \U$6031 ( \6408 , \5765 );
or \U$6032 ( \6409 , \6407 , \6408 );
not \U$6033 ( \6410 , RIae79160_138);
not \U$6034 ( \6411 , \2564 );
or \U$6035 ( \6412 , \6410 , \6411 );
not \U$6036 ( \6413 , \2563 );
not \U$6037 ( \6414 , RIae79160_138);
nand \U$6038 ( \6415 , \6413 , \6414 );
nand \U$6039 ( \6416 , \6412 , \6415 );
nand \U$6040 ( \6417 , \6416 , \1009 );
nand \U$6041 ( \6418 , \6409 , \6417 );
xor \U$6042 ( \6419 , \6406 , \6418 );
not \U$6043 ( \6420 , \2341 );
not \U$6044 ( \6421 , \6144 );
or \U$6045 ( \6422 , \6420 , \6421 );
nand \U$6046 ( \6423 , \5552 , \2322 );
nand \U$6047 ( \6424 , \6422 , \6423 );
and \U$6048 ( \6425 , \6419 , \6424 );
and \U$6049 ( \6426 , \6406 , \6418 );
or \U$6050 ( \6427 , \6425 , \6426 );
xor \U$6051 ( \6428 , \5593 , \5602 );
xor \U$6052 ( \6429 , \6428 , \5612 );
xor \U$6053 ( \6430 , \6427 , \6429 );
xor \U$6054 ( \6431 , \5625 , \5635 );
xor \U$6055 ( \6432 , \6431 , \5643 );
and \U$6056 ( \6433 , \6430 , \6432 );
and \U$6057 ( \6434 , \6427 , \6429 );
or \U$6058 ( \6435 , \6433 , \6434 );
xor \U$6059 ( \6436 , \6396 , \6435 );
xor \U$6060 ( \6437 , \5681 , \5659 );
xor \U$6061 ( \6438 , \5759 , \5769 );
xor \U$6062 ( \6439 , \6438 , \5779 );
xor \U$6063 ( \6440 , \6437 , \6439 );
xor \U$6064 ( \6441 , \5531 , \5554 );
not \U$6065 ( \6442 , \5558 );
xor \U$6066 ( \6443 , \6441 , \6442 );
and \U$6067 ( \6444 , \6440 , \6443 );
and \U$6068 ( \6445 , \6437 , \6439 );
or \U$6069 ( \6446 , \6444 , \6445 );
and \U$6070 ( \6447 , \6436 , \6446 );
and \U$6071 ( \6448 , \6396 , \6435 );
or \U$6072 ( \6449 , \6447 , \6448 );
xor \U$6073 ( \6450 , \6332 , \6449 );
xnor \U$6074 ( \6451 , \5690 , \5788 );
and \U$6075 ( \6452 , \6451 , \5702 );
not \U$6076 ( \6453 , \6451 );
and \U$6077 ( \6454 , \6453 , \5701 );
nor \U$6078 ( \6455 , \6452 , \6454 );
and \U$6079 ( \6456 , \6450 , \6455 );
and \U$6080 ( \6457 , \6332 , \6449 );
or \U$6081 ( \6458 , \6456 , \6457 );
and \U$6082 ( \6459 , \6320 , \6458 );
xor \U$6083 ( \6460 , \5796 , \5791 );
xor \U$6084 ( \6461 , \6460 , \5582 );
nor \U$6085 ( \6462 , \6459 , \6461 );
nor \U$6086 ( \6463 , \6320 , \6458 );
nor \U$6087 ( \6464 , \6462 , \6463 );
nand \U$6088 ( \6465 , \6053 , \6464 );
nand \U$6089 ( \6466 , \6052 , \6465 );
not \U$6090 ( \6467 , \6466 );
nand \U$6091 ( \6468 , \5843 , \6467 );
not \U$6092 ( \6469 , \3981 );
not \U$6093 ( \6470 , \4238 );
not \U$6094 ( \6471 , \3941 );
or \U$6095 ( \6472 , \6470 , \6471 );
or \U$6096 ( \6473 , \4238 , \3941 );
nand \U$6097 ( \6474 , \6472 , \6473 );
not \U$6098 ( \6475 , \6474 );
or \U$6099 ( \6476 , \6469 , \6475 );
or \U$6100 ( \6477 , \6474 , \3981 );
nand \U$6101 ( \6478 , \6476 , \6477 );
not \U$6102 ( \6479 , \6478 );
not \U$6103 ( \6480 , \5810 );
not \U$6104 ( \6481 , \5826 );
or \U$6105 ( \6482 , \6480 , \6481 );
not \U$6106 ( \6483 , \5814 );
nand \U$6107 ( \6484 , \6483 , \5822 );
nand \U$6108 ( \6485 , \6482 , \6484 );
not \U$6109 ( \6486 , \6485 );
and \U$6110 ( \6487 , \6479 , \6486 );
and \U$6111 ( \6488 , \6485 , \6478 );
nor \U$6112 ( \6489 , \6487 , \6488 );
not \U$6113 ( \6490 , \6489 );
not \U$6114 ( \6491 , \3916 );
not \U$6115 ( \6492 , \3878 );
or \U$6116 ( \6493 , \6491 , \6492 );
or \U$6117 ( \6494 , \3878 , \3916 );
nand \U$6118 ( \6495 , \6493 , \6494 );
xor \U$6119 ( \6496 , \6495 , \3923 );
not \U$6120 ( \6497 , \6496 );
or \U$6121 ( \6498 , \6490 , \6497 );
or \U$6122 ( \6499 , \6496 , \6489 );
nand \U$6123 ( \6500 , \6498 , \6499 );
not \U$6124 ( \6501 , \6500 );
not \U$6125 ( \6502 , \5841 );
not \U$6126 ( \6503 , \5832 );
or \U$6127 ( \6504 , \6502 , \6503 );
not \U$6128 ( \6505 , \5806 );
nand \U$6129 ( \6506 , \6504 , \6505 );
not \U$6130 ( \6507 , \5841 );
not \U$6131 ( \6508 , \5832 );
nand \U$6132 ( \6509 , \6507 , \6508 );
nand \U$6133 ( \6510 , \6506 , \6509 );
not \U$6134 ( \6511 , \6510 );
xor \U$6135 ( \6512 , \4812 , \4819 );
and \U$6136 ( \6513 , \6512 , \4878 );
and \U$6137 ( \6514 , \4812 , \4819 );
or \U$6138 ( \6515 , \6513 , \6514 );
not \U$6139 ( \6516 , \6515 );
not \U$6140 ( \6517 , \6516 );
and \U$6141 ( \6518 , \6511 , \6517 );
and \U$6142 ( \6519 , \6510 , \6516 );
nor \U$6143 ( \6520 , \6518 , \6519 );
not \U$6144 ( \6521 , \6520 );
or \U$6145 ( \6522 , \6501 , \6521 );
or \U$6146 ( \6523 , \6520 , \6500 );
nand \U$6147 ( \6524 , \6522 , \6523 );
xor \U$6148 ( \6525 , \4879 , \5801 );
and \U$6149 ( \6526 , \6525 , \5842 );
and \U$6150 ( \6527 , \4879 , \5801 );
or \U$6151 ( \6528 , \6526 , \6527 );
nand \U$6152 ( \6529 , \6524 , \6528 );
and \U$6153 ( \6530 , \6468 , \6529 );
not \U$6154 ( \6531 , \6489 );
not \U$6155 ( \6532 , \6531 );
not \U$6156 ( \6533 , \6496 );
or \U$6157 ( \6534 , \6532 , \6533 );
not \U$6158 ( \6535 , \6485 );
nand \U$6159 ( \6536 , \6535 , \6478 );
nand \U$6160 ( \6537 , \6534 , \6536 );
not \U$6161 ( \6538 , \6537 );
xor \U$6162 ( \6539 , \2502 , \2748 );
xor \U$6163 ( \6540 , \6539 , \2889 );
not \U$6164 ( \6541 , \6540 );
xor \U$6165 ( \6542 , \3931 , \4240 );
not \U$6166 ( \6543 , \3925 );
and \U$6167 ( \6544 , \6542 , \6543 );
not \U$6168 ( \6545 , \6542 );
and \U$6169 ( \6546 , \6545 , \3925 );
nor \U$6170 ( \6547 , \6544 , \6546 );
not \U$6171 ( \6548 , \6547 );
or \U$6172 ( \6549 , \6541 , \6548 );
or \U$6173 ( \6550 , \6540 , \6547 );
nand \U$6174 ( \6551 , \6549 , \6550 );
not \U$6175 ( \6552 , \6551 );
not \U$6176 ( \6553 , \6552 );
or \U$6177 ( \6554 , \6538 , \6553 );
not \U$6178 ( \6555 , \6537 );
nand \U$6179 ( \6556 , \6555 , \6551 );
nand \U$6180 ( \6557 , \6554 , \6556 );
not \U$6181 ( \6558 , \6500 );
not \U$6182 ( \6559 , \6520 );
not \U$6183 ( \6560 , \6559 );
or \U$6184 ( \6561 , \6558 , \6560 );
not \U$6185 ( \6562 , \6516 );
nand \U$6186 ( \6563 , \6562 , \6510 );
nand \U$6187 ( \6564 , \6561 , \6563 );
nand \U$6188 ( \6565 , \6557 , \6564 );
not \U$6189 ( \6566 , \6540 );
nand \U$6190 ( \6567 , \6566 , \6547 );
not \U$6191 ( \6568 , \6567 );
nand \U$6192 ( \6569 , \6551 , \6537 );
not \U$6193 ( \6570 , \6569 );
or \U$6194 ( \6571 , \6568 , \6570 );
xor \U$6195 ( \6572 , \4245 , \3875 );
xnor \U$6196 ( \6573 , \6572 , \3873 );
nand \U$6197 ( \6574 , \6571 , \6573 );
and \U$6198 ( \6575 , \6530 , \6565 , \6574 );
not \U$6199 ( \6576 , \4782 );
nand \U$6200 ( \6577 , \6576 , \4791 );
not \U$6201 ( \6578 , \6577 );
nand \U$6202 ( \6579 , \4796 , \4702 );
not \U$6203 ( \6580 , \6579 );
or \U$6204 ( \6581 , \6578 , \6580 );
not \U$6205 ( \6582 , \4777 );
not \U$6206 ( \6583 , \4713 );
or \U$6207 ( \6584 , \6582 , \6583 );
not \U$6208 ( \6585 , \4708 );
nand \U$6209 ( \6586 , \6585 , \4712 );
nand \U$6210 ( \6587 , \6584 , \6586 );
not \U$6211 ( \6588 , \4698 );
not \U$6212 ( \6589 , \6588 );
not \U$6213 ( \6590 , \4535 );
or \U$6214 ( \6591 , \6589 , \6590 );
nand \U$6215 ( \6592 , \6591 , \4700 );
xor \U$6216 ( \6593 , \6587 , \6592 );
not \U$6217 ( \6594 , \4763 );
or \U$6218 ( \6595 , \4774 , \4768 );
not \U$6219 ( \6596 , \6595 );
or \U$6220 ( \6597 , \6594 , \6596 );
nand \U$6221 ( \6598 , \4774 , \4768 );
nand \U$6222 ( \6599 , \6597 , \6598 );
not \U$6223 ( \6600 , \4604 );
not \U$6224 ( \6601 , \4592 );
or \U$6225 ( \6602 , \6600 , \6601 );
nand \U$6226 ( \6603 , \4591 , \4578 );
nand \U$6227 ( \6604 , \6602 , \6603 );
and \U$6228 ( \6605 , RIae79160_138, \2027 );
not \U$6229 ( \6606 , RIae79160_138);
and \U$6230 ( \6607 , \6606 , \2031 );
nor \U$6231 ( \6608 , \6605 , \6607 );
or \U$6232 ( \6609 , \1210 , \6608 );
not \U$6233 ( \6610 , \4739 );
not \U$6234 ( \6611 , \1010 );
or \U$6235 ( \6612 , \6610 , \6611 );
nand \U$6236 ( \6613 , \6609 , \6612 );
not \U$6237 ( \6614 , \4760 );
not \U$6238 ( \6615 , \2966 );
or \U$6239 ( \6616 , \6614 , \6615 );
and \U$6240 ( \6617 , RIae79688_149, \1068 );
not \U$6241 ( \6618 , RIae79688_149);
and \U$6242 ( \6619 , \6618 , \3443 );
nor \U$6243 ( \6620 , \6617 , \6619 );
not \U$6244 ( \6621 , \6620 );
not \U$6245 ( \6622 , \1822 );
or \U$6246 ( \6623 , \6621 , \6622 );
nand \U$6247 ( \6624 , \6616 , \6623 );
xor \U$6248 ( \6625 , \6613 , \6624 );
not \U$6249 ( \6626 , RIae79520_146);
not \U$6250 ( \6627 , \835 );
or \U$6251 ( \6628 , \6626 , \6627 );
or \U$6252 ( \6629 , \829 , RIae79520_146);
nand \U$6253 ( \6630 , \6628 , \6629 );
not \U$6254 ( \6631 , \6630 );
not \U$6255 ( \6632 , \2610 );
or \U$6256 ( \6633 , \6631 , \6632 );
not \U$6257 ( \6634 , \4658 );
not \U$6258 ( \6635 , \2189 );
or \U$6259 ( \6636 , \6634 , \6635 );
nand \U$6260 ( \6637 , \6633 , \6636 );
xor \U$6261 ( \6638 , \6625 , \6637 );
xor \U$6262 ( \6639 , \6604 , \6638 );
nand \U$6263 ( \6640 , \4305 , RIae78b48_125);
not \U$6264 ( \6641 , \868 );
not \U$6265 ( \6642 , \3095 );
xor \U$6266 ( \6643 , RIae78b48_125, \6642 );
not \U$6267 ( \6644 , \6643 );
or \U$6268 ( \6645 , \6641 , \6644 );
or \U$6269 ( \6646 , \4589 , \1976 );
nand \U$6270 ( \6647 , \6645 , \6646 );
xor \U$6271 ( \6648 , \6640 , \6647 );
not \U$6272 ( \6649 , \3015 );
not \U$6273 ( \6650 , RIae79ac0_158);
not \U$6274 ( \6651 , \1146 );
or \U$6275 ( \6652 , \6650 , \6651 );
or \U$6276 ( \6653 , \1143 , RIae79ac0_158);
nand \U$6277 ( \6654 , \6652 , \6653 );
not \U$6278 ( \6655 , \6654 );
or \U$6279 ( \6656 , \6649 , \6655 );
or \U$6280 ( \6657 , \4614 , \3510 );
nand \U$6281 ( \6658 , \6656 , \6657 );
xnor \U$6282 ( \6659 , \6648 , \6658 );
xor \U$6283 ( \6660 , \6639 , \6659 );
xor \U$6284 ( \6661 , \6599 , \6660 );
not \U$6285 ( \6662 , \797 );
not \U$6286 ( \6663 , \4679 );
or \U$6287 ( \6664 , \6662 , \6663 );
not \U$6288 ( \6665 , \4480 );
and \U$6289 ( \6666 , RIae78f80_134, \6665 );
not \U$6290 ( \6667 , RIae78f80_134);
buf \U$6291 ( \6668 , \3052 );
and \U$6292 ( \6669 , \6667 , \6668 );
nor \U$6293 ( \6670 , \6666 , \6669 );
nand \U$6294 ( \6671 , \840 , \6670 );
nand \U$6295 ( \6672 , \6664 , \6671 );
not \U$6296 ( \6673 , \2011 );
not \U$6297 ( \6674 , RIae79610_148);
not \U$6298 ( \6675 , \6674 );
not \U$6299 ( \6676 , \856 );
or \U$6300 ( \6677 , \6675 , \6676 );
nand \U$6301 ( \6678 , \857 , RIae79610_148);
nand \U$6302 ( \6679 , \6677 , \6678 );
not \U$6303 ( \6680 , \6679 );
or \U$6304 ( \6681 , \6673 , \6680 );
nand \U$6305 ( \6682 , \4572 , \2063 );
nand \U$6306 ( \6683 , \6681 , \6682 );
not \U$6307 ( \6684 , \1049 );
and \U$6308 ( \6685 , RIae79070_136, \1879 );
not \U$6309 ( \6686 , RIae79070_136);
and \U$6310 ( \6687 , \6686 , \1880 );
nor \U$6311 ( \6688 , \6685 , \6687 );
not \U$6312 ( \6689 , \6688 );
or \U$6313 ( \6690 , \6684 , \6689 );
nand \U$6314 ( \6691 , \4667 , \1062 );
nand \U$6315 ( \6692 , \6690 , \6691 );
xor \U$6316 ( \6693 , \6683 , \6692 );
xor \U$6317 ( \6694 , \6672 , \6693 );
not \U$6318 ( \6695 , \6694 );
not \U$6319 ( \6696 , \4545 );
not \U$6320 ( \6697 , \3520 );
and \U$6321 ( \6698 , \6696 , \6697 );
xor \U$6322 ( \6699 , \2310 , RIae78bc0_126);
and \U$6323 ( \6700 , \6699 , \1028 );
nor \U$6324 ( \6701 , \6698 , \6700 );
not \U$6325 ( \6702 , \6701 );
not \U$6326 ( \6703 , \1864 );
not \U$6327 ( \6704 , RIae793b8_143);
not \U$6328 ( \6705 , \1119 );
or \U$6329 ( \6706 , \6704 , \6705 );
or \U$6330 ( \6707 , \1472 , RIae793b8_143);
nand \U$6331 ( \6708 , \6706 , \6707 );
not \U$6332 ( \6709 , \6708 );
or \U$6333 ( \6710 , \6703 , \6709 );
nand \U$6334 ( \6711 , \4598 , \1910 );
nand \U$6335 ( \6712 , \6710 , \6711 );
not \U$6336 ( \6713 , \6712 );
or \U$6337 ( \6714 , \6702 , \6713 );
or \U$6338 ( \6715 , \6701 , \6712 );
nand \U$6339 ( \6716 , \6714 , \6715 );
not \U$6340 ( \6717 , \6716 );
not \U$6341 ( \6718 , \921 );
not \U$6342 ( \6719 , \3072 );
not \U$6343 ( \6720 , \6719 );
or \U$6344 ( \6721 , \6718 , \6720 );
nand \U$6345 ( \6722 , \4358 , RIae78e90_132);
nand \U$6346 ( \6723 , \6721 , \6722 );
and \U$6347 ( \6724 , \6723 , \1322 );
and \U$6348 ( \6725 , \4559 , \1259 );
nor \U$6349 ( \6726 , \6724 , \6725 );
not \U$6350 ( \6727 , \6726 );
and \U$6351 ( \6728 , \6717 , \6727 );
and \U$6352 ( \6729 , \6716 , \6726 );
nor \U$6353 ( \6730 , \6728 , \6729 );
not \U$6354 ( \6731 , \6730 );
or \U$6355 ( \6732 , \6695 , \6731 );
or \U$6356 ( \6733 , \6730 , \6694 );
nand \U$6357 ( \6734 , \6732 , \6733 );
not \U$6358 ( \6735 , \4725 );
not \U$6359 ( \6736 , \4732 );
not \U$6360 ( \6737 , \4316 );
or \U$6361 ( \6738 , \6736 , \6737 );
or \U$6362 ( \6739 , \4732 , \4316 );
nand \U$6363 ( \6740 , \6738 , \6739 );
not \U$6364 ( \6741 , \6740 );
or \U$6365 ( \6742 , \6735 , \6741 );
nand \U$6366 ( \6743 , \4732 , \4315 );
nand \U$6367 ( \6744 , \6742 , \6743 );
xor \U$6368 ( \6745 , \6734 , \6744 );
xor \U$6369 ( \6746 , \6661 , \6745 );
xor \U$6370 ( \6747 , \4637 , \4642 );
and \U$6371 ( \6748 , \6747 , \4696 );
and \U$6372 ( \6749 , \4637 , \4642 );
or \U$6373 ( \6750 , \6748 , \6749 );
xor \U$6374 ( \6751 , \6746 , \6750 );
not \U$6375 ( \6752 , \4690 );
not \U$6376 ( \6753 , \4695 );
or \U$6377 ( \6754 , \6752 , \6753 );
not \U$6378 ( \6755 , \4648 );
nand \U$6379 ( \6756 , \6755 , \4686 );
nand \U$6380 ( \6757 , \6754 , \6756 );
not \U$6381 ( \6758 , \6757 );
not \U$6382 ( \6759 , \4776 );
not \U$6383 ( \6760 , \4733 );
not \U$6384 ( \6761 , \6760 );
or \U$6385 ( \6762 , \6759 , \6761 );
not \U$6386 ( \6763 , \4775 );
not \U$6387 ( \6764 , \4733 );
or \U$6388 ( \6765 , \6763 , \6764 );
nand \U$6389 ( \6766 , \6765 , \4719 );
nand \U$6390 ( \6767 , \6762 , \6766 );
xor \U$6391 ( \6768 , \6758 , \6767 );
not \U$6392 ( \6769 , \1933 );
not \U$6393 ( \6770 , \4623 );
or \U$6394 ( \6771 , \6769 , \6770 );
nand \U$6395 ( \6772 , \1919 , RIae794a8_145);
nand \U$6396 ( \6773 , \6771 , \6772 );
not \U$6397 ( \6774 , \6773 );
not \U$6398 ( \6775 , \1501 );
xnor \U$6399 ( \6776 , \1187 , RIae79250_140);
not \U$6400 ( \6777 , \6776 );
or \U$6401 ( \6778 , \6775 , \6777 );
nand \U$6402 ( \6779 , \4748 , \1499 );
nand \U$6403 ( \6780 , \6778 , \6779 );
xor \U$6404 ( \6781 , \6774 , \6780 );
not \U$6405 ( \6782 , \4574 );
not \U$6406 ( \6783 , \4565 );
or \U$6407 ( \6784 , \6782 , \6783 );
not \U$6408 ( \6785 , \4550 );
nand \U$6409 ( \6786 , \6785 , \4561 );
nand \U$6410 ( \6787 , \6784 , \6786 );
xor \U$6411 ( \6788 , \6781 , \6787 );
xor \U$6412 ( \6789 , \4743 , \4752 );
and \U$6413 ( \6790 , \6789 , \4762 );
and \U$6414 ( \6791 , \4743 , \4752 );
or \U$6415 ( \6792 , \6790 , \6791 );
not \U$6416 ( \6793 , \4616 );
not \U$6417 ( \6794 , \4607 );
not \U$6418 ( \6795 , \4627 );
or \U$6419 ( \6796 , \6794 , \6795 );
or \U$6420 ( \6797 , \4627 , \4607 );
nand \U$6421 ( \6798 , \6796 , \6797 );
not \U$6422 ( \6799 , \6798 );
or \U$6423 ( \6800 , \6793 , \6799 );
not \U$6424 ( \6801 , \4607 );
nand \U$6425 ( \6802 , \6801 , \4627 );
nand \U$6426 ( \6803 , \6800 , \6802 );
xor \U$6427 ( \6804 , \6792 , \6803 );
not \U$6428 ( \6805 , \4681 );
not \U$6429 ( \6806 , \4670 );
or \U$6430 ( \6807 , \6805 , \6806 );
nand \U$6431 ( \6808 , \4669 , \4660 );
nand \U$6432 ( \6809 , \6807 , \6808 );
xor \U$6433 ( \6810 , \6804 , \6809 );
xor \U$6434 ( \6811 , \6788 , \6810 );
not \U$6435 ( \6812 , \4575 );
not \U$6436 ( \6813 , \4633 );
or \U$6437 ( \6814 , \6812 , \6813 );
not \U$6438 ( \6815 , \4605 );
nand \U$6439 ( \6816 , \6815 , \4629 );
nand \U$6440 ( \6817 , \6814 , \6816 );
not \U$6441 ( \6818 , \6817 );
xor \U$6442 ( \6819 , \6811 , \6818 );
xor \U$6443 ( \6820 , \6768 , \6819 );
xor \U$6444 ( \6821 , \6751 , \6820 );
xor \U$6445 ( \6822 , \6593 , \6821 );
nand \U$6446 ( \6823 , \6581 , \6822 );
buf \U$6447 ( \6824 , \6823 );
and \U$6448 ( \6825 , \4811 , \6575 , \6824 );
not \U$6449 ( \6826 , \1322 );
and \U$6450 ( \6827 , \6668 , \1066 );
not \U$6451 ( \6828 , \6668 );
and \U$6452 ( \6829 , \6828 , RIae78e90_132);
nor \U$6453 ( \6830 , \6827 , \6829 );
not \U$6454 ( \6831 , \6830 );
or \U$6455 ( \6832 , \6826 , \6831 );
xor \U$6456 ( \6833 , RIae78e90_132, \2231 );
not \U$6457 ( \6834 , \6833 );
or \U$6458 ( \6835 , \6834 , \1413 );
nand \U$6459 ( \6836 , \6832 , \6835 );
and \U$6460 ( \6837 , RIae793b8_143, \1024 );
not \U$6461 ( \6838 , RIae793b8_143);
and \U$6462 ( \6839 , \6838 , \858 );
nor \U$6463 ( \6840 , \6837 , \6839 );
or \U$6464 ( \6841 , \6840 , \3494 );
and \U$6465 ( \6842 , RIae793b8_143, \879 );
not \U$6466 ( \6843 , RIae793b8_143);
and \U$6467 ( \6844 , \6843 , \883 );
nor \U$6468 ( \6845 , \6842 , \6844 );
not \U$6469 ( \6846 , \1910 );
or \U$6470 ( \6847 , \6845 , \6846 );
nand \U$6471 ( \6848 , \6841 , \6847 );
and \U$6472 ( \6849 , \6836 , \6848 );
not \U$6473 ( \6850 , \6836 );
not \U$6474 ( \6851 , \6848 );
and \U$6475 ( \6852 , \6850 , \6851 );
nor \U$6476 ( \6853 , \6849 , \6852 );
not \U$6477 ( \6854 , \840 );
not \U$6478 ( \6855 , \1880 );
xor \U$6479 ( \6856 , \6855 , RIae78f80_134);
not \U$6480 ( \6857 , \6856 );
or \U$6481 ( \6858 , \6854 , \6857 );
and \U$6482 ( \6859 , \3785 , RIae78f80_134);
and \U$6483 ( \6860 , \3294 , \1132 );
nor \U$6484 ( \6861 , \6859 , \6860 );
or \U$6485 ( \6862 , \6861 , \798 );
nand \U$6486 ( \6863 , \6858 , \6862 );
xor \U$6487 ( \6864 , \6853 , \6863 );
not \U$6488 ( \6865 , \6864 );
not \U$6489 ( \6866 , \1501 );
and \U$6490 ( \6867 , RIae79250_140, \1120 );
not \U$6491 ( \6868 , RIae79250_140);
and \U$6492 ( \6869 , \6868 , \1472 );
nor \U$6493 ( \6870 , \6867 , \6869 );
not \U$6494 ( \6871 , \6870 );
or \U$6495 ( \6872 , \6866 , \6871 );
and \U$6496 ( \6873 , RIae79250_140, \3718 );
not \U$6497 ( \6874 , RIae79250_140);
and \U$6498 ( \6875 , \6874 , \3722 );
nor \U$6499 ( \6876 , \6873 , \6875 );
nand \U$6500 ( \6877 , \6876 , \2650 );
nand \U$6501 ( \6878 , \6872 , \6877 );
not \U$6502 ( \6879 , \6878 );
xor \U$6503 ( \6880 , RIae78b48_125, \2309 );
nand \U$6504 ( \6881 , \6880 , \868 );
and \U$6505 ( \6882 , RIae78b48_125, \2287 );
not \U$6506 ( \6883 , RIae78b48_125);
and \U$6507 ( \6884 , \6883 , \3748 );
nor \U$6508 ( \6885 , \6882 , \6884 );
not \U$6509 ( \6886 , \6885 );
nand \U$6510 ( \6887 , \6886 , \1129 );
and \U$6511 ( \6888 , \6881 , \6887 );
not \U$6512 ( \6889 , \6888 );
and \U$6513 ( \6890 , \6879 , \6889 );
and \U$6514 ( \6891 , \6878 , \6888 );
nor \U$6515 ( \6892 , \6890 , \6891 );
and \U$6516 ( \6893 , RIae78bc0_126, \4358 );
not \U$6517 ( \6894 , RIae78bc0_126);
and \U$6518 ( \6895 , \6894 , \6719 );
nor \U$6519 ( \6896 , \6893 , \6895 );
not \U$6520 ( \6897 , \6896 );
not \U$6521 ( \6898 , \1029 );
and \U$6522 ( \6899 , \6897 , \6898 );
and \U$6523 ( \6900 , \1286 , \4555 );
not \U$6524 ( \6901 , \1286 );
not \U$6525 ( \6902 , \4555 );
and \U$6526 ( \6903 , \6901 , \6902 );
nor \U$6527 ( \6904 , \6900 , \6903 );
and \U$6528 ( \6905 , \6904 , \1036 );
nor \U$6529 ( \6906 , \6899 , \6905 );
not \U$6530 ( \6907 , \6906 );
and \U$6531 ( \6908 , \6892 , \6907 );
not \U$6532 ( \6909 , \6892 );
and \U$6533 ( \6910 , \6909 , \6906 );
nor \U$6534 ( \6911 , \6908 , \6910 );
not \U$6535 ( \6912 , \6911 );
not \U$6536 ( \6913 , \3443 );
and \U$6537 ( \6914 , RIae79610_148, \6913 );
not \U$6538 ( \6915 , RIae79610_148);
and \U$6539 ( \6916 , \6915 , \1440 );
nor \U$6540 ( \6917 , \6914 , \6916 );
and \U$6541 ( \6918 , \6917 , \2011 );
xnor \U$6542 ( \6919 , \3775 , RIae79610_148);
and \U$6543 ( \6920 , \6919 , \4344 );
nor \U$6544 ( \6921 , \6918 , \6920 );
not \U$6545 ( \6922 , \6921 );
not \U$6546 ( \6923 , \3015 );
and \U$6547 ( \6924 , \835 , \2268 );
not \U$6548 ( \6925 , \835 );
and \U$6549 ( \6926 , \6925 , RIae79ac0_158);
nor \U$6550 ( \6927 , \6924 , \6926 );
not \U$6551 ( \6928 , \6927 );
or \U$6552 ( \6929 , \6923 , \6928 );
not \U$6553 ( \6930 , RIae79ac0_158);
not \U$6554 ( \6931 , \1993 );
or \U$6555 ( \6932 , \6930 , \6931 );
or \U$6556 ( \6933 , \3286 , RIae79ac0_158);
nand \U$6557 ( \6934 , \6932 , \6933 );
nand \U$6558 ( \6935 , \6934 , \2272 );
nand \U$6559 ( \6936 , \6929 , \6935 );
not \U$6560 ( \6937 , \6936 );
or \U$6561 ( \6938 , \6922 , \6937 );
or \U$6562 ( \6939 , \6936 , \6921 );
nand \U$6563 ( \6940 , \6938 , \6939 );
not \U$6564 ( \6941 , \1062 );
and \U$6565 ( \6942 , RIae79070_136, \2050 );
not \U$6566 ( \6943 , RIae79070_136);
and \U$6567 ( \6944 , \6943 , \2049 );
nor \U$6568 ( \6945 , \6942 , \6944 );
not \U$6569 ( \6946 , \6945 );
or \U$6570 ( \6947 , \6941 , \6946 );
and \U$6571 ( \6948 , RIae79070_136, \2027 );
not \U$6572 ( \6949 , RIae79070_136);
and \U$6573 ( \6950 , \6949 , \5137 );
nor \U$6574 ( \6951 , \6948 , \6950 );
or \U$6575 ( \6952 , \6951 , \1203 );
nand \U$6576 ( \6953 , \6947 , \6952 );
xor \U$6577 ( \6954 , \6940 , \6953 );
not \U$6578 ( \6955 , \6954 );
or \U$6579 ( \6956 , \6912 , \6955 );
or \U$6580 ( \6957 , \6954 , \6911 );
nand \U$6581 ( \6958 , \6956 , \6957 );
not \U$6582 ( \6959 , \6958 );
or \U$6583 ( \6960 , \6865 , \6959 );
not \U$6584 ( \6961 , \6911 );
nand \U$6585 ( \6962 , \6961 , \6954 );
nand \U$6586 ( \6963 , \6960 , \6962 );
not \U$6587 ( \6964 , \6963 );
and \U$6588 ( \6965 , \6904 , \1028 );
and \U$6589 ( \6966 , \6699 , \953 );
nor \U$6590 ( \6967 , \6965 , \6966 );
not \U$6591 ( \6968 , \6967 );
not \U$6592 ( \6969 , \6968 );
not \U$6593 ( \6970 , \893 );
not \U$6594 ( \6971 , \6643 );
or \U$6595 ( \6972 , \6970 , \6971 );
or \U$6596 ( \6973 , \6885 , \1959 );
nand \U$6597 ( \6974 , \6972 , \6973 );
not \U$6598 ( \6975 , \1910 );
not \U$6599 ( \6976 , \6708 );
or \U$6600 ( \6977 , \6975 , \6976 );
not \U$6601 ( \6978 , \6845 );
nand \U$6602 ( \6979 , \6978 , \1864 );
nand \U$6603 ( \6980 , \6977 , \6979 );
xor \U$6604 ( \6981 , \6974 , \6980 );
not \U$6605 ( \6982 , \6981 );
or \U$6606 ( \6983 , \6969 , \6982 );
nand \U$6607 ( \6984 , \6980 , \6974 );
nand \U$6608 ( \6985 , \6983 , \6984 );
not \U$6609 ( \6986 , \6985 );
not \U$6610 ( \6987 , \3827 );
and \U$6611 ( \6988 , RIae79688_149, \1159 );
not \U$6612 ( \6989 , RIae79688_149);
and \U$6613 ( \6990 , \6989 , \1162 );
nor \U$6614 ( \6991 , \6988 , \6990 );
not \U$6615 ( \6992 , \6991 );
or \U$6616 ( \6993 , \6987 , \6992 );
nand \U$6617 ( \6994 , \6620 , \2966 );
nand \U$6618 ( \6995 , \6993 , \6994 );
not \U$6619 ( \6996 , \6995 );
and \U$6620 ( \6997 , \1914 , RIae794a8_145);
not \U$6621 ( \6998 , \6997 );
not \U$6622 ( \6999 , RIae79520_146);
not \U$6623 ( \7000 , \1196 );
or \U$6624 ( \7001 , \6999 , \7000 );
or \U$6625 ( \7002 , \992 , RIae79520_146);
nand \U$6626 ( \7003 , \7001 , \7002 );
or \U$6627 ( \7004 , \7003 , \6632 );
nand \U$6628 ( \7005 , \6630 , \2189 );
nand \U$6629 ( \7006 , \7004 , \7005 );
not \U$6630 ( \7007 , \7006 );
or \U$6631 ( \7008 , \6998 , \7007 );
or \U$6632 ( \7009 , \7006 , \6997 );
nand \U$6633 ( \7010 , \7008 , \7009 );
not \U$6634 ( \7011 , \7010 );
or \U$6635 ( \7012 , \6996 , \7011 );
not \U$6636 ( \7013 , \6997 );
nand \U$6637 ( \7014 , \7013 , \7006 );
nand \U$6638 ( \7015 , \7012 , \7014 );
and \U$6639 ( \7016 , RIae78b48_125, \6642 );
not \U$6640 ( \7017 , \3827 );
and \U$6641 ( \7018 , RIae79688_149, \1146 );
not \U$6642 ( \7019 , RIae79688_149);
and \U$6643 ( \7020 , \7019 , \1147 );
or \U$6644 ( \7021 , \7018 , \7020 );
not \U$6645 ( \7022 , \7021 );
or \U$6646 ( \7023 , \7017 , \7022 );
nand \U$6647 ( \7024 , \6991 , \1844 );
nand \U$6648 ( \7025 , \7023 , \7024 );
xor \U$6649 ( \7026 , \7016 , \7025 );
not \U$6650 ( \7027 , \7026 );
not \U$6651 ( \7028 , \1013 );
and \U$6652 ( \7029 , \1187 , \997 );
not \U$6653 ( \7030 , \1187 );
and \U$6654 ( \7031 , \7030 , RIae79160_138);
nor \U$6655 ( \7032 , \7029 , \7031 );
not \U$6656 ( \7033 , \7032 );
or \U$6657 ( \7034 , \7028 , \7033 );
and \U$6658 ( \7035 , RIae79160_138, \1835 );
not \U$6659 ( \7036 , RIae79160_138);
and \U$6660 ( \7037 , \7036 , \6147 );
nor \U$6661 ( \7038 , \7035 , \7037 );
nand \U$6662 ( \7039 , \1430 , \7038 );
nand \U$6663 ( \7040 , \7034 , \7039 );
not \U$6664 ( \7041 , \7040 );
not \U$6665 ( \7042 , \7041 );
and \U$6666 ( \7043 , \7027 , \7042 );
and \U$6667 ( \7044 , \7026 , \7041 );
nor \U$6668 ( \7045 , \7043 , \7044 );
and \U$6669 ( \7046 , \7015 , \7045 );
not \U$6670 ( \7047 , \7015 );
not \U$6671 ( \7048 , \7045 );
and \U$6672 ( \7049 , \7047 , \7048 );
or \U$6673 ( \7050 , \7046 , \7049 );
not \U$6674 ( \7051 , \7050 );
or \U$6675 ( \7052 , \6986 , \7051 );
nand \U$6676 ( \7053 , \7015 , \7048 );
nand \U$6677 ( \7054 , \7052 , \7053 );
not \U$6678 ( \7055 , \7054 );
or \U$6679 ( \7056 , \6892 , \6906 );
not \U$6680 ( \7057 , \6888 );
nand \U$6681 ( \7058 , \7057 , \6878 );
nand \U$6682 ( \7059 , \7056 , \7058 );
not \U$6683 ( \7060 , \7059 );
and \U$6684 ( \7061 , \7026 , \7040 );
and \U$6685 ( \7062 , \7016 , \7025 );
nor \U$6686 ( \7063 , \7061 , \7062 );
not \U$6687 ( \7064 , \7063 );
and \U$6688 ( \7065 , \7060 , \7064 );
and \U$6689 ( \7066 , \7059 , \7063 );
nor \U$6690 ( \7067 , \7065 , \7066 );
not \U$6691 ( \7068 , \7067 );
not \U$6692 ( \7069 , \6953 );
not \U$6693 ( \7070 , \6940 );
or \U$6694 ( \7071 , \7069 , \7070 );
not \U$6695 ( \7072 , \6921 );
nand \U$6696 ( \7073 , \7072 , \6936 );
nand \U$6697 ( \7074 , \7071 , \7073 );
not \U$6698 ( \7075 , \7074 );
and \U$6699 ( \7076 , \7068 , \7075 );
and \U$6700 ( \7077 , \7067 , \7074 );
nor \U$6701 ( \7078 , \7076 , \7077 );
not \U$6702 ( \7079 , \7078 );
or \U$6703 ( \7080 , \7055 , \7079 );
or \U$6704 ( \7081 , \7054 , \7078 );
nand \U$6705 ( \7082 , \7080 , \7081 );
not \U$6706 ( \7083 , \7082 );
or \U$6707 ( \7084 , \6964 , \7083 );
not \U$6708 ( \7085 , \7078 );
nand \U$6709 ( \7086 , \7085 , \7054 );
nand \U$6710 ( \7087 , \7084 , \7086 );
not \U$6711 ( \7088 , \7074 );
not \U$6712 ( \7089 , \7067 );
not \U$6713 ( \7090 , \7089 );
or \U$6714 ( \7091 , \7088 , \7090 );
not \U$6715 ( \7092 , \7063 );
nand \U$6716 ( \7093 , \7092 , \7059 );
nand \U$6717 ( \7094 , \7091 , \7093 );
not \U$6718 ( \7095 , \7094 );
not \U$6719 ( \7096 , \1910 );
not \U$6720 ( \7097 , \6840 );
not \U$6721 ( \7098 , \7097 );
or \U$6722 ( \7099 , \7096 , \7098 );
and \U$6723 ( \7100 , RIae793b8_143, \940 );
not \U$6724 ( \7101 , RIae793b8_143);
and \U$6725 ( \7102 , \7101 , \941 );
nor \U$6726 ( \7103 , \7100 , \7102 );
not \U$6727 ( \7104 , \7103 );
nand \U$6728 ( \7105 , \7104 , \1864 );
nand \U$6729 ( \7106 , \7099 , \7105 );
and \U$6730 ( \7107 , \1039 , \1406 );
not \U$6731 ( \7108 , \1039 );
and \U$6732 ( \7109 , \7108 , \1834 );
nor \U$6733 ( \7110 , \7107 , \7109 );
or \U$6734 ( \7111 , \7110 , \1203 );
or \U$6735 ( \7112 , \6951 , \1249 );
nand \U$6736 ( \7113 , \7111 , \7112 );
xor \U$6737 ( \7114 , \7106 , \7113 );
and \U$6738 ( \7115 , \2594 , \1132 );
and \U$6739 ( \7116 , \2595 , RIae78f80_134);
nor \U$6740 ( \7117 , \7115 , \7116 );
and \U$6741 ( \7118 , \7117 , \840 );
and \U$6742 ( \7119 , \6856 , \797 );
nor \U$6743 ( \7120 , \7118 , \7119 );
not \U$6744 ( \7121 , \7120 );
and \U$6745 ( \7122 , \7114 , \7121 );
not \U$6746 ( \7123 , \7114 );
and \U$6747 ( \7124 , \7123 , \7120 );
nor \U$6748 ( \7125 , \7122 , \7124 );
not \U$6749 ( \7126 , \7125 );
not \U$6750 ( \7127 , \2272 );
not \U$6751 ( \7128 , \6927 );
or \U$6752 ( \7129 , \7127 , \7128 );
and \U$6753 ( \7130 , \992 , RIae79ac0_158);
not \U$6754 ( \7131 , \992 );
and \U$6755 ( \7132 , \7131 , \2268 );
nor \U$6756 ( \7133 , \7130 , \7132 );
nand \U$6757 ( \7134 , \7133 , \3015 );
nand \U$6758 ( \7135 , \7129 , \7134 );
or \U$6759 ( \7136 , \2602 , \3440 );
nand \U$6760 ( \7137 , \7136 , RIae79520_146);
xor \U$6761 ( \7138 , \7135 , \7137 );
and \U$6762 ( \7139 , \1162 , \2056 );
and \U$6763 ( \7140 , \1159 , RIae79610_148);
nor \U$6764 ( \7141 , \7139 , \7140 );
and \U$6765 ( \7142 , \7141 , \2011 );
and \U$6766 ( \7143 , \6917 , \2063 );
nor \U$6767 ( \7144 , \7142 , \7143 );
not \U$6768 ( \7145 , \7144 );
xor \U$6769 ( \7146 , \7138 , \7145 );
not \U$6770 ( \7147 , \7146 );
not \U$6771 ( \7148 , \7147 );
not \U$6772 ( \7149 , \929 );
xor \U$6773 ( \7150 , \2995 , RIae78bc0_126);
not \U$6774 ( \7151 , \7150 );
or \U$6775 ( \7152 , \7149 , \7151 );
not \U$6776 ( \7153 , \6896 );
nand \U$6777 ( \7154 , \7153 , \1036 );
nand \U$6778 ( \7155 , \7152 , \7154 );
not \U$6779 ( \7156 , \2966 );
not \U$6780 ( \7157 , \7021 );
or \U$6781 ( \7158 , \7156 , \7157 );
and \U$6782 ( \7159 , RIae79688_149, \3814 );
not \U$6783 ( \7160 , RIae79688_149);
and \U$6784 ( \7161 , \7160 , \782 );
nor \U$6785 ( \7162 , \7159 , \7161 );
not \U$6786 ( \7163 , \3827 );
or \U$6787 ( \7164 , \7162 , \7163 );
nand \U$6788 ( \7165 , \7158 , \7164 );
xor \U$6789 ( \7166 , \7155 , \7165 );
xor \U$6790 ( \7167 , \1899 , RIae78e90_132);
and \U$6791 ( \7168 , \7167 , \1322 );
and \U$6792 ( \7169 , \6830 , \1259 );
nor \U$6793 ( \7170 , \7168 , \7169 );
not \U$6794 ( \7171 , \7170 );
xor \U$6795 ( \7172 , \7166 , \7171 );
not \U$6796 ( \7173 , \7172 );
or \U$6797 ( \7174 , \7148 , \7173 );
or \U$6798 ( \7175 , \7172 , \7147 );
nand \U$6799 ( \7176 , \7174 , \7175 );
not \U$6800 ( \7177 , \7176 );
or \U$6801 ( \7178 , \7126 , \7177 );
not \U$6802 ( \7179 , \7147 );
nand \U$6803 ( \7180 , \7179 , \7172 );
nand \U$6804 ( \7181 , \7178 , \7180 );
not \U$6805 ( \7182 , \7181 );
not \U$6806 ( \7183 , \7182 );
or \U$6807 ( \7184 , \7095 , \7183 );
not \U$6808 ( \7185 , \7094 );
nand \U$6809 ( \7186 , \7185 , \7181 );
nand \U$6810 ( \7187 , \7184 , \7186 );
xor \U$6811 ( \7188 , \7135 , \7137 );
not \U$6812 ( \7189 , \7144 );
and \U$6813 ( \7190 , \7188 , \7189 );
and \U$6814 ( \7191 , \7135 , \7137 );
or \U$6815 ( \7192 , \7190 , \7191 );
not \U$6816 ( \7193 , \7192 );
not \U$6817 ( \7194 , \7193 );
and \U$6818 ( \7195 , RIae78b48_125, \4555 );
not \U$6819 ( \7196 , RIae78b48_125);
and \U$6820 ( \7197 , \7196 , \6902 );
nor \U$6821 ( \7198 , \7195 , \7197 );
or \U$6822 ( \7199 , \7198 , \1603 );
not \U$6823 ( \7200 , \6880 );
or \U$6824 ( \7201 , \7200 , \1128 );
nand \U$6825 ( \7202 , \7199 , \7201 );
not \U$6826 ( \7203 , \7202 );
nand \U$6827 ( \7204 , \3748 , RIae78b48_125);
not \U$6828 ( \7205 , \6870 );
not \U$6829 ( \7206 , \7205 );
not \U$6830 ( \7207 , \1498 );
and \U$6831 ( \7208 , \7206 , \7207 );
and \U$6832 ( \7209 , RIae79250_140, \3256 );
not \U$6833 ( \7210 , RIae79250_140);
and \U$6834 ( \7211 , \7210 , \884 );
nor \U$6835 ( \7212 , \7209 , \7211 );
and \U$6836 ( \7213 , \7212 , \1501 );
nor \U$6837 ( \7214 , \7208 , \7213 );
xor \U$6838 ( \7215 , \7204 , \7214 );
not \U$6839 ( \7216 , \7215 );
or \U$6840 ( \7217 , \7203 , \7216 );
or \U$6841 ( \7218 , \7214 , \7204 );
nand \U$6842 ( \7219 , \7217 , \7218 );
not \U$6843 ( \7220 , \7219 );
and \U$6844 ( \7221 , \7194 , \7220 );
and \U$6845 ( \7222 , \7219 , \7193 );
nor \U$6846 ( \7223 , \7221 , \7222 );
not \U$6847 ( \7224 , \7223 );
xor \U$6848 ( \7225 , \7155 , \7165 );
not \U$6849 ( \7226 , \7170 );
and \U$6850 ( \7227 , \7225 , \7226 );
and \U$6851 ( \7228 , \7155 , \7165 );
or \U$6852 ( \7229 , \7227 , \7228 );
not \U$6853 ( \7230 , \7229 );
and \U$6854 ( \7231 , \7224 , \7230 );
and \U$6855 ( \7232 , \7223 , \7229 );
nor \U$6856 ( \7233 , \7231 , \7232 );
not \U$6857 ( \7234 , \7233 );
and \U$6858 ( \7235 , \7187 , \7234 );
not \U$6859 ( \7236 , \7187 );
and \U$6860 ( \7237 , \7236 , \7233 );
nor \U$6861 ( \7238 , \7235 , \7237 );
nor \U$6862 ( \7239 , \7087 , \7238 );
not \U$6863 ( \7240 , \7239 );
not \U$6864 ( \7241 , \7240 );
and \U$6865 ( \7242 , \6945 , \1049 );
and \U$6866 ( \7243 , \6688 , \1062 );
nor \U$6867 ( \7244 , \7242 , \7243 );
not \U$6868 ( \7245 , \7244 );
not \U$6869 ( \7246 , \1013 );
not \U$6870 ( \7247 , \7038 );
or \U$6871 ( \7248 , \7246 , \7247 );
not \U$6872 ( \7249 , \6608 );
nand \U$6873 ( \7250 , \7249 , \1430 );
nand \U$6874 ( \7251 , \7248 , \7250 );
not \U$6875 ( \7252 , \7251 );
or \U$6876 ( \7253 , \7245 , \7252 );
or \U$6877 ( \7254 , \7251 , \7244 );
nand \U$6878 ( \7255 , \7253 , \7254 );
and \U$6879 ( \7256 , \6919 , \2011 );
and \U$6880 ( \7257 , \6679 , \2063 );
nor \U$6881 ( \7258 , \7256 , \7257 );
not \U$6882 ( \7259 , \7258 );
and \U$6883 ( \7260 , \7255 , \7259 );
not \U$6884 ( \7261 , \7255 );
and \U$6885 ( \7262 , \7261 , \7258 );
nor \U$6886 ( \7263 , \7260 , \7262 );
not \U$6887 ( \7264 , \7263 );
not \U$6888 ( \7265 , \6640 );
xor \U$6889 ( \7266 , \7265 , \6658 );
and \U$6890 ( \7267 , \7266 , \6647 );
and \U$6891 ( \7268 , \7265 , \6658 );
nor \U$6892 ( \7269 , \7267 , \7268 );
not \U$6893 ( \7270 , \7269 );
not \U$6894 ( \7271 , \1499 );
not \U$6895 ( \7272 , \6776 );
or \U$6896 ( \7273 , \7271 , \7272 );
not \U$6897 ( \7274 , \6876 );
or \U$6898 ( \7275 , \7274 , \1502 );
nand \U$6899 ( \7276 , \7273 , \7275 );
nand \U$6900 ( \7277 , \4584 , RIae78b48_125);
not \U$6901 ( \7278 , \7277 );
not \U$6902 ( \7279 , \6773 );
or \U$6903 ( \7280 , \7278 , \7279 );
or \U$6904 ( \7281 , \6773 , \7277 );
nand \U$6905 ( \7282 , \7280 , \7281 );
xor \U$6906 ( \7283 , \7276 , \7282 );
not \U$6907 ( \7284 , \7283 );
or \U$6908 ( \7285 , \7270 , \7284 );
or \U$6909 ( \7286 , \7283 , \7269 );
nand \U$6910 ( \7287 , \7285 , \7286 );
not \U$6911 ( \7288 , \7287 );
or \U$6912 ( \7289 , \7264 , \7288 );
not \U$6913 ( \7290 , \7269 );
nand \U$6914 ( \7291 , \7290 , \7283 );
nand \U$6915 ( \7292 , \7289 , \7291 );
not \U$6916 ( \7293 , \7292 );
not \U$6917 ( \7294 , \6985 );
not \U$6918 ( \7295 , \7294 );
not \U$6919 ( \7296 , \7050 );
or \U$6920 ( \7297 , \7295 , \7296 );
or \U$6921 ( \7298 , \7050 , \7294 );
nand \U$6922 ( \7299 , \7297 , \7298 );
not \U$6923 ( \7300 , \6967 );
not \U$6924 ( \7301 , \6981 );
or \U$6925 ( \7302 , \7300 , \7301 );
or \U$6926 ( \7303 , \6981 , \6967 );
nand \U$6927 ( \7304 , \7302 , \7303 );
not \U$6928 ( \7305 , \7304 );
xnor \U$6929 ( \7306 , \7010 , \6995 );
not \U$6930 ( \7307 , \7306 );
not \U$6931 ( \7308 , \797 );
not \U$6932 ( \7309 , \6670 );
or \U$6933 ( \7310 , \7308 , \7309 );
or \U$6934 ( \7311 , \6861 , \1227 );
nand \U$6935 ( \7312 , \7310 , \7311 );
not \U$6936 ( \7313 , \7312 );
not \U$6937 ( \7314 , \7313 );
not \U$6938 ( \7315 , \2272 );
not \U$6939 ( \7316 , \6654 );
or \U$6940 ( \7317 , \7315 , \7316 );
nand \U$6941 ( \7318 , \6934 , \3015 );
nand \U$6942 ( \7319 , \7317 , \7318 );
not \U$6943 ( \7320 , \1074 );
not \U$6944 ( \7321 , \6833 );
or \U$6945 ( \7322 , \7320 , \7321 );
nand \U$6946 ( \7323 , \6723 , \1087 );
nand \U$6947 ( \7324 , \7322 , \7323 );
xor \U$6948 ( \7325 , \7319 , \7324 );
not \U$6949 ( \7326 , \7325 );
or \U$6950 ( \7327 , \7314 , \7326 );
not \U$6951 ( \7328 , \7325 );
nand \U$6952 ( \7329 , \7328 , \7312 );
nand \U$6953 ( \7330 , \7327 , \7329 );
not \U$6954 ( \7331 , \7330 );
or \U$6955 ( \7332 , \7307 , \7331 );
or \U$6956 ( \7333 , \7306 , \7330 );
nand \U$6957 ( \7334 , \7332 , \7333 );
not \U$6958 ( \7335 , \7334 );
or \U$6959 ( \7336 , \7305 , \7335 );
not \U$6960 ( \7337 , \7306 );
nand \U$6961 ( \7338 , \7337 , \7330 );
nand \U$6962 ( \7339 , \7336 , \7338 );
xor \U$6963 ( \7340 , \7299 , \7339 );
not \U$6964 ( \7341 , \7340 );
or \U$6965 ( \7342 , \7293 , \7341 );
nand \U$6966 ( \7343 , \7299 , \7339 );
nand \U$6967 ( \7344 , \7342 , \7343 );
not \U$6968 ( \7345 , \7344 );
xor \U$6969 ( \7346 , \7176 , \7125 );
nand \U$6970 ( \7347 , \7325 , \7312 );
nand \U$6971 ( \7348 , \7324 , \7319 );
and \U$6972 ( \7349 , \7347 , \7348 );
not \U$6973 ( \7350 , \7244 );
not \U$6974 ( \7351 , \7350 );
not \U$6975 ( \7352 , \7251 );
or \U$6976 ( \7353 , \7351 , \7352 );
nand \U$6977 ( \7354 , \7255 , \7259 );
nand \U$6978 ( \7355 , \7353 , \7354 );
not \U$6979 ( \7356 , \7003 );
not \U$6980 ( \7357 , \6635 );
and \U$6981 ( \7358 , \7356 , \7357 );
and \U$6982 ( \7359 , \2610 , RIae79520_146);
nor \U$6983 ( \7360 , \7358 , \7359 );
not \U$6984 ( \7361 , \7360 );
and \U$6985 ( \7362 , \7355 , \7361 );
not \U$6986 ( \7363 , \7355 );
and \U$6987 ( \7364 , \7363 , \7360 );
or \U$6988 ( \7365 , \7362 , \7364 );
xnor \U$6989 ( \7366 , \7349 , \7365 );
not \U$6990 ( \7367 , \7366 );
not \U$6991 ( \7368 , \6774 );
not \U$6992 ( \7369 , \7277 );
and \U$6993 ( \7370 , \7368 , \7369 );
and \U$6994 ( \7371 , \7282 , \7276 );
nor \U$6995 ( \7372 , \7370 , \7371 );
not \U$6996 ( \7373 , \7372 );
not \U$6997 ( \7374 , \7373 );
xor \U$6998 ( \7375 , \6613 , \6624 );
and \U$6999 ( \7376 , \7375 , \6637 );
and \U$7000 ( \7377 , \6613 , \6624 );
or \U$7001 ( \7378 , \7376 , \7377 );
not \U$7002 ( \7379 , \6672 );
not \U$7003 ( \7380 , \6693 );
or \U$7004 ( \7381 , \7379 , \7380 );
nand \U$7005 ( \7382 , \6683 , \6692 );
nand \U$7006 ( \7383 , \7381 , \7382 );
xor \U$7007 ( \7384 , \7378 , \7383 );
not \U$7008 ( \7385 , \7384 );
not \U$7009 ( \7386 , \6723 );
or \U$7010 ( \7387 , \7386 , \1646 );
not \U$7011 ( \7388 , \4559 );
or \U$7012 ( \7389 , \7388 , \1413 );
nand \U$7013 ( \7390 , \7387 , \7389 );
not \U$7014 ( \7391 , \7390 );
not \U$7015 ( \7392 , \6716 );
or \U$7016 ( \7393 , \7391 , \7392 );
not \U$7017 ( \7394 , \6701 );
nand \U$7018 ( \7395 , \7394 , \6712 );
nand \U$7019 ( \7396 , \7393 , \7395 );
not \U$7020 ( \7397 , \7396 );
or \U$7021 ( \7398 , \7385 , \7397 );
nand \U$7022 ( \7399 , \7383 , \7378 );
nand \U$7023 ( \7400 , \7398 , \7399 );
not \U$7024 ( \7401 , \7400 );
not \U$7025 ( \7402 , \7401 );
or \U$7026 ( \7403 , \7374 , \7402 );
nand \U$7027 ( \7404 , \7400 , \7372 );
nand \U$7028 ( \7405 , \7403 , \7404 );
not \U$7029 ( \7406 , \7405 );
or \U$7030 ( \7407 , \7367 , \7406 );
nand \U$7031 ( \7408 , \7400 , \7373 );
nand \U$7032 ( \7409 , \7407 , \7408 );
xor \U$7033 ( \7410 , \7346 , \7409 );
not \U$7034 ( \7411 , \7410 );
or \U$7035 ( \7412 , \7345 , \7411 );
nand \U$7036 ( \7413 , \7409 , \7346 );
nand \U$7037 ( \7414 , \7412 , \7413 );
not \U$7038 ( \7415 , \7414 );
or \U$7039 ( \7416 , \7241 , \7415 );
nand \U$7040 ( \7417 , \7087 , \7238 );
nand \U$7041 ( \7418 , \7416 , \7417 );
not \U$7042 ( \7419 , \7418 );
not \U$7043 ( \7420 , \7360 );
not \U$7044 ( \7421 , \7355 );
or \U$7045 ( \7422 , \7420 , \7421 );
not \U$7046 ( \7423 , \7349 );
nand \U$7047 ( \7424 , \7423 , \7365 );
nand \U$7048 ( \7425 , \7422 , \7424 );
not \U$7049 ( \7426 , \7425 );
not \U$7050 ( \7427 , \7032 );
not \U$7051 ( \7428 , \7427 );
not \U$7052 ( \7429 , \1430 );
not \U$7053 ( \7430 , \7429 );
and \U$7054 ( \7431 , \7428 , \7430 );
and \U$7055 ( \7432 , RIae79160_138, \3718 );
not \U$7056 ( \7433 , RIae79160_138);
and \U$7057 ( \7434 , \7433 , \1125 );
nor \U$7058 ( \7435 , \7432 , \7434 );
and \U$7059 ( \7436 , \7435 , \1013 );
nor \U$7060 ( \7437 , \7431 , \7436 );
and \U$7061 ( \7438 , \7437 , \7361 );
not \U$7062 ( \7439 , \7437 );
and \U$7063 ( \7440 , \7439 , \7360 );
nor \U$7064 ( \7441 , \7438 , \7440 );
not \U$7065 ( \7442 , \7441 );
not \U$7066 ( \7443 , \6863 );
not \U$7067 ( \7444 , \6853 );
or \U$7068 ( \7445 , \7443 , \7444 );
nand \U$7069 ( \7446 , \6836 , \6848 );
nand \U$7070 ( \7447 , \7445 , \7446 );
not \U$7071 ( \7448 , \7447 );
or \U$7072 ( \7449 , \7442 , \7448 );
or \U$7073 ( \7450 , \7447 , \7441 );
nand \U$7074 ( \7451 , \7449 , \7450 );
xnor \U$7075 ( \7452 , \7215 , \7202 );
xor \U$7076 ( \7453 , \7451 , \7452 );
not \U$7077 ( \7454 , \7453 );
not \U$7078 ( \7455 , \7454 );
or \U$7079 ( \7456 , \7426 , \7455 );
not \U$7080 ( \7457 , \7452 );
nand \U$7081 ( \7458 , \7457 , \7451 );
nand \U$7082 ( \7459 , \7456 , \7458 );
not \U$7083 ( \7460 , \7459 );
and \U$7084 ( \7461 , \2053 , \1143 );
not \U$7085 ( \7462 , \2053 );
and \U$7086 ( \7463 , \7462 , \1366 );
nor \U$7087 ( \7464 , \7461 , \7463 );
and \U$7088 ( \7465 , \7464 , \2011 );
and \U$7089 ( \7466 , \7141 , \2063 );
nor \U$7090 ( \7467 , \7465 , \7466 );
not \U$7091 ( \7468 , \7467 );
and \U$7092 ( \7469 , RIae78b48_125, \2309 );
not \U$7093 ( \7470 , \868 );
xor \U$7094 ( \7471 , RIae78b48_125, \4081 );
not \U$7095 ( \7472 , \7471 );
or \U$7096 ( \7473 , \7470 , \7472 );
not \U$7097 ( \7474 , \7198 );
nand \U$7098 ( \7475 , \7474 , \893 );
nand \U$7099 ( \7476 , \7473 , \7475 );
xor \U$7100 ( \7477 , \7469 , \7476 );
not \U$7101 ( \7478 , \7477 );
or \U$7102 ( \7479 , \7468 , \7478 );
or \U$7103 ( \7480 , \7477 , \7467 );
nand \U$7104 ( \7481 , \7479 , \7480 );
not \U$7105 ( \7482 , \7481 );
and \U$7106 ( \7483 , \7114 , \7121 );
and \U$7107 ( \7484 , \7106 , \7113 );
nor \U$7108 ( \7485 , \7483 , \7484 );
not \U$7109 ( \7486 , \7485 );
or \U$7110 ( \7487 , \7482 , \7486 );
or \U$7111 ( \7488 , \7481 , \7485 );
nand \U$7112 ( \7489 , \7487 , \7488 );
xnor \U$7113 ( \7490 , \1119 , RIae79160_138);
and \U$7114 ( \7491 , \7490 , \1209 );
and \U$7115 ( \7492 , \7435 , \1430 );
nor \U$7116 ( \7493 , \7491 , \7492 );
not \U$7117 ( \7494 , \1049 );
xor \U$7118 ( \7495 , \1188 , RIae79070_136);
not \U$7119 ( \7496 , \7495 );
or \U$7120 ( \7497 , \7494 , \7496 );
not \U$7121 ( \7498 , \7110 );
nand \U$7122 ( \7499 , \7498 , \1062 );
nand \U$7123 ( \7500 , \7497 , \7499 );
not \U$7124 ( \7501 , \2272 );
not \U$7125 ( \7502 , \7133 );
or \U$7126 ( \7503 , \7501 , \7502 );
nand \U$7127 ( \7504 , \3015 , RIae79ac0_158);
nand \U$7128 ( \7505 , \7503 , \7504 );
and \U$7129 ( \7506 , \7500 , \7505 );
not \U$7130 ( \7507 , \7500 );
not \U$7131 ( \7508 , \7505 );
and \U$7132 ( \7509 , \7507 , \7508 );
nor \U$7133 ( \7510 , \7506 , \7509 );
xor \U$7134 ( \7511 , \7493 , \7510 );
xor \U$7135 ( \7512 , \7489 , \7511 );
not \U$7136 ( \7513 , \7447 );
or \U$7137 ( \7514 , \7513 , \7441 );
or \U$7138 ( \7515 , \7437 , \7360 );
nand \U$7139 ( \7516 , \7514 , \7515 );
xor \U$7140 ( \7517 , RIae79250_140, \858 );
and \U$7141 ( \7518 , \7517 , \1501 );
and \U$7142 ( \7519 , \7212 , \1499 );
nor \U$7143 ( \7520 , \7518 , \7519 );
not \U$7144 ( \7521 , \7520 );
and \U$7145 ( \7522 , RIae78e90_132, \4458 );
not \U$7146 ( \7523 , RIae78e90_132);
and \U$7147 ( \7524 , \7523 , \6855 );
nor \U$7148 ( \7525 , \7522 , \7524 );
not \U$7149 ( \7526 , \7525 );
not \U$7150 ( \7527 , \1646 );
and \U$7151 ( \7528 , \7526 , \7527 );
and \U$7152 ( \7529 , \7167 , \1087 );
nor \U$7153 ( \7530 , \7528 , \7529 );
not \U$7154 ( \7531 , \1036 );
not \U$7155 ( \7532 , \7150 );
or \U$7156 ( \7533 , \7531 , \7532 );
and \U$7157 ( \7534 , RIae78bc0_126, \6665 );
not \U$7158 ( \7535 , RIae78bc0_126);
and \U$7159 ( \7536 , \7535 , \6668 );
nor \U$7160 ( \7537 , \7534 , \7536 );
nand \U$7161 ( \7538 , \7537 , \1028 );
nand \U$7162 ( \7539 , \7533 , \7538 );
not \U$7163 ( \7540 , \7539 );
and \U$7164 ( \7541 , \7530 , \7540 );
not \U$7165 ( \7542 , \7530 );
and \U$7166 ( \7543 , \7542 , \7539 );
nor \U$7167 ( \7544 , \7541 , \7543 );
not \U$7168 ( \7545 , \7544 );
or \U$7169 ( \7546 , \7521 , \7545 );
or \U$7170 ( \7547 , \7520 , \7544 );
nand \U$7171 ( \7548 , \7546 , \7547 );
and \U$7172 ( \7549 , RIae78f80_134, \5137 );
not \U$7173 ( \7550 , RIae78f80_134);
and \U$7174 ( \7551 , \7550 , \2374 );
nor \U$7175 ( \7552 , \7549 , \7551 );
and \U$7176 ( \7553 , \7552 , \839 );
and \U$7177 ( \7554 , \7117 , \797 );
nor \U$7178 ( \7555 , \7553 , \7554 );
and \U$7179 ( \7556 , \1884 , \1441 );
not \U$7180 ( \7557 , \1884 );
not \U$7181 ( \7558 , \1068 );
and \U$7182 ( \7559 , \7557 , \7558 );
nor \U$7183 ( \7560 , \7556 , \7559 );
or \U$7184 ( \7561 , \7560 , \3494 );
or \U$7185 ( \7562 , \7103 , \6846 );
nand \U$7186 ( \7563 , \7561 , \7562 );
and \U$7187 ( \7564 , \7555 , \7563 );
not \U$7188 ( \7565 , \7555 );
not \U$7189 ( \7566 , \7563 );
and \U$7190 ( \7567 , \7565 , \7566 );
or \U$7191 ( \7568 , \7564 , \7567 );
and \U$7192 ( \7569 , \835 , \3147 );
not \U$7193 ( \7570 , \835 );
and \U$7194 ( \7571 , \7570 , RIae79688_149);
nor \U$7195 ( \7572 , \7569 , \7571 );
not \U$7196 ( \7573 , \7572 );
or \U$7197 ( \7574 , \7573 , \6622 );
not \U$7198 ( \7575 , \2966 );
or \U$7199 ( \7576 , \7162 , \7575 );
nand \U$7200 ( \7577 , \7574 , \7576 );
not \U$7201 ( \7578 , \7577 );
and \U$7202 ( \7579 , \7568 , \7578 );
not \U$7203 ( \7580 , \7568 );
and \U$7204 ( \7581 , \7580 , \7577 );
nor \U$7205 ( \7582 , \7579 , \7581 );
xor \U$7206 ( \7583 , \7548 , \7582 );
xnor \U$7207 ( \7584 , \7516 , \7583 );
xor \U$7208 ( \7585 , \7512 , \7584 );
not \U$7209 ( \7586 , \7585 );
or \U$7210 ( \7587 , \7460 , \7586 );
nand \U$7211 ( \7588 , \7584 , \7512 );
nand \U$7212 ( \7589 , \7587 , \7588 );
and \U$7213 ( \7590 , RIae79250_140, \939 );
not \U$7214 ( \7591 , RIae79250_140);
and \U$7215 ( \7592 , \7591 , \944 );
nor \U$7216 ( \7593 , \7590 , \7592 );
and \U$7217 ( \7594 , \7593 , \1501 );
and \U$7218 ( \7595 , \7517 , \1499 );
nor \U$7219 ( \7596 , \7594 , \7595 );
not \U$7220 ( \7597 , \7596 );
not \U$7221 ( \7598 , \7525 );
not \U$7222 ( \7599 , \1413 );
and \U$7223 ( \7600 , \7598 , \7599 );
xnor \U$7224 ( \7601 , \2049 , RIae78e90_132);
and \U$7225 ( \7602 , \7601 , \1074 );
nor \U$7226 ( \7603 , \7600 , \7602 );
and \U$7227 ( \7604 , RIae78f80_134, \1834 );
not \U$7228 ( \7605 , RIae78f80_134);
and \U$7229 ( \7606 , \7605 , \6148 );
nor \U$7230 ( \7607 , \7604 , \7606 );
not \U$7231 ( \7608 , \7607 );
not \U$7232 ( \7609 , \3112 );
and \U$7233 ( \7610 , \7608 , \7609 );
and \U$7234 ( \7611 , \7552 , \797 );
nor \U$7235 ( \7612 , \7610 , \7611 );
xor \U$7236 ( \7613 , \7603 , \7612 );
not \U$7237 ( \7614 , \7613 );
or \U$7238 ( \7615 , \7597 , \7614 );
or \U$7239 ( \7616 , \7613 , \7596 );
nand \U$7240 ( \7617 , \7615 , \7616 );
and \U$7241 ( \7618 , \1162 , RIae793b8_143);
and \U$7242 ( \7619 , \1291 , \1902 );
nor \U$7243 ( \7620 , \7618 , \7619 );
or \U$7244 ( \7621 , \7620 , \3494 );
or \U$7245 ( \7622 , \7560 , \6846 );
nand \U$7246 ( \7623 , \7621 , \7622 );
nand \U$7247 ( \7624 , RIae79520_146, RIae79a48_157);
and \U$7248 ( \7625 , \7624 , RIae79ac0_158);
not \U$7249 ( \7626 , \1822 );
not \U$7250 ( \7627 , \992 );
not \U$7251 ( \7628 , RIae79688_149);
and \U$7252 ( \7629 , \7627 , \7628 );
and \U$7253 ( \7630 , \994 , RIae79688_149);
nor \U$7254 ( \7631 , \7629 , \7630 );
not \U$7255 ( \7632 , \7631 );
or \U$7256 ( \7633 , \7626 , \7632 );
nand \U$7257 ( \7634 , \7572 , \2966 );
nand \U$7258 ( \7635 , \7633 , \7634 );
and \U$7259 ( \7636 , \7625 , \7635 );
not \U$7260 ( \7637 , \7625 );
not \U$7261 ( \7638 , \7635 );
and \U$7262 ( \7639 , \7637 , \7638 );
or \U$7263 ( \7640 , \7636 , \7639 );
xor \U$7264 ( \7641 , \7623 , \7640 );
xor \U$7265 ( \7642 , \7617 , \7641 );
not \U$7266 ( \7643 , \1129 );
not \U$7267 ( \7644 , \7471 );
or \U$7268 ( \7645 , \7643 , \7644 );
and \U$7269 ( \7646 , RIae78b48_125, \4675 );
not \U$7270 ( \7647 , RIae78b48_125);
and \U$7271 ( \7648 , \7647 , \2231 );
nor \U$7272 ( \7649 , \7646 , \7648 );
not \U$7273 ( \7650 , \7649 );
nand \U$7274 ( \7651 , \7650 , \868 );
nand \U$7275 ( \7652 , \7645 , \7651 );
not \U$7276 ( \7653 , \1036 );
not \U$7277 ( \7654 , \7537 );
or \U$7278 ( \7655 , \7653 , \7654 );
and \U$7279 ( \7656 , RIae78bc0_126, \3785 );
not \U$7280 ( \7657 , RIae78bc0_126);
and \U$7281 ( \7658 , \7657 , \1899 );
nor \U$7282 ( \7659 , \7656 , \7658 );
or \U$7283 ( \7660 , \7659 , \928 );
nand \U$7284 ( \7661 , \7655 , \7660 );
xor \U$7285 ( \7662 , \7652 , \7661 );
xnor \U$7286 ( \7663 , \1993 , RIae79610_148);
and \U$7287 ( \7664 , \7663 , \2011 );
and \U$7288 ( \7665 , \7464 , \2063 );
nor \U$7289 ( \7666 , \7664 , \7665 );
not \U$7290 ( \7667 , \7666 );
and \U$7291 ( \7668 , \7662 , \7667 );
not \U$7292 ( \7669 , \7662 );
and \U$7293 ( \7670 , \7669 , \7666 );
nor \U$7294 ( \7671 , \7668 , \7670 );
and \U$7295 ( \7672 , \7642 , \7671 );
not \U$7296 ( \7673 , \7642 );
not \U$7297 ( \7674 , \7671 );
and \U$7298 ( \7675 , \7673 , \7674 );
nor \U$7299 ( \7676 , \7672 , \7675 );
not \U$7300 ( \7677 , \7583 );
nand \U$7301 ( \7678 , \7677 , \7516 );
not \U$7302 ( \7679 , \7582 );
nand \U$7303 ( \7680 , \7679 , \7548 );
and \U$7304 ( \7681 , \7678 , \7680 );
xor \U$7305 ( \7682 , \7676 , \7681 );
not \U$7306 ( \7683 , \7544 );
or \U$7307 ( \7684 , \7683 , \7520 );
or \U$7308 ( \7685 , \7540 , \7530 );
nand \U$7309 ( \7686 , \7684 , \7685 );
not \U$7310 ( \7687 , \7686 );
not \U$7311 ( \7688 , \7510 );
not \U$7312 ( \7689 , \7493 );
and \U$7313 ( \7690 , \7688 , \7689 );
and \U$7314 ( \7691 , \7500 , \7508 );
nor \U$7315 ( \7692 , \7690 , \7691 );
not \U$7316 ( \7693 , \7692 );
or \U$7317 ( \7694 , \7687 , \7693 );
or \U$7318 ( \7695 , \7692 , \7686 );
nand \U$7319 ( \7696 , \7694 , \7695 );
not \U$7320 ( \7697 , \1062 );
not \U$7321 ( \7698 , \7495 );
or \U$7322 ( \7699 , \7697 , \7698 );
and \U$7323 ( \7700 , RIae79070_136, \3722 );
not \U$7324 ( \7701 , RIae79070_136);
not \U$7325 ( \7702 , \3722 );
and \U$7326 ( \7703 , \7701 , \7702 );
nor \U$7327 ( \7704 , \7700 , \7703 );
not \U$7328 ( \7705 , \7704 );
nand \U$7329 ( \7706 , \7705 , \1049 );
nand \U$7330 ( \7707 , \7699 , \7706 );
and \U$7331 ( \7708 , \6902 , RIae78b48_125);
and \U$7332 ( \7709 , \7707 , \7708 );
not \U$7333 ( \7710 , \7707 );
not \U$7334 ( \7711 , \7708 );
and \U$7335 ( \7712 , \7710 , \7711 );
nor \U$7336 ( \7713 , \7709 , \7712 );
not \U$7337 ( \7714 , \1010 );
not \U$7338 ( \7715 , \7490 );
or \U$7339 ( \7716 , \7714 , \7715 );
and \U$7340 ( \7717 , RIae79160_138, \879 );
not \U$7341 ( \7718 , RIae79160_138);
and \U$7342 ( \7719 , \7718 , \3256 );
nor \U$7343 ( \7720 , \7717 , \7719 );
or \U$7344 ( \7721 , \7720 , \1210 );
nand \U$7345 ( \7722 , \7716 , \7721 );
xor \U$7346 ( \7723 , \7713 , \7722 );
and \U$7347 ( \7724 , \7696 , \7723 );
not \U$7348 ( \7725 , \7696 );
not \U$7349 ( \7726 , \7723 );
and \U$7350 ( \7727 , \7725 , \7726 );
nor \U$7351 ( \7728 , \7724 , \7727 );
xnor \U$7352 ( \7729 , \7682 , \7728 );
xor \U$7353 ( \7730 , \7589 , \7729 );
nand \U$7354 ( \7731 , \7182 , \7233 );
and \U$7355 ( \7732 , \7731 , \7094 );
nor \U$7356 ( \7733 , \7233 , \7182 );
nor \U$7357 ( \7734 , \7732 , \7733 );
not \U$7358 ( \7735 , \7734 );
not \U$7359 ( \7736 , \7193 );
not \U$7360 ( \7737 , \7736 );
not \U$7361 ( \7738 , \7219 );
or \U$7362 ( \7739 , \7737 , \7738 );
not \U$7363 ( \7740 , \7229 );
or \U$7364 ( \7741 , \7223 , \7740 );
nand \U$7365 ( \7742 , \7739 , \7741 );
not \U$7366 ( \7743 , \7742 );
not \U$7367 ( \7744 , \7566 );
not \U$7368 ( \7745 , \7555 );
and \U$7369 ( \7746 , \7744 , \7745 );
and \U$7370 ( \7747 , \7568 , \7577 );
nor \U$7371 ( \7748 , \7746 , \7747 );
not \U$7372 ( \7749 , \7748 );
not \U$7373 ( \7750 , \7467 );
not \U$7374 ( \7751 , \7750 );
not \U$7375 ( \7752 , \7477 );
or \U$7376 ( \7753 , \7751 , \7752 );
nand \U$7377 ( \7754 , \7476 , \7469 );
nand \U$7378 ( \7755 , \7753 , \7754 );
and \U$7379 ( \7756 , \7755 , \7505 );
not \U$7380 ( \7757 , \7755 );
and \U$7381 ( \7758 , \7757 , \7508 );
nor \U$7382 ( \7759 , \7756 , \7758 );
not \U$7383 ( \7760 , \7759 );
or \U$7384 ( \7761 , \7749 , \7760 );
or \U$7385 ( \7762 , \7759 , \7748 );
nand \U$7386 ( \7763 , \7761 , \7762 );
not \U$7387 ( \7764 , \7511 );
not \U$7388 ( \7765 , \7489 );
or \U$7389 ( \7766 , \7764 , \7765 );
not \U$7390 ( \7767 , \7485 );
nand \U$7391 ( \7768 , \7767 , \7481 );
nand \U$7392 ( \7769 , \7766 , \7768 );
xor \U$7393 ( \7770 , \7763 , \7769 );
not \U$7394 ( \7771 , \7770 );
not \U$7395 ( \7772 , \7771 );
or \U$7396 ( \7773 , \7743 , \7772 );
not \U$7397 ( \7774 , \7742 );
nand \U$7398 ( \7775 , \7774 , \7770 );
nand \U$7399 ( \7776 , \7773 , \7775 );
not \U$7400 ( \7777 , \7776 );
or \U$7401 ( \7778 , \7735 , \7777 );
or \U$7402 ( \7779 , \7776 , \7734 );
nand \U$7403 ( \7780 , \7778 , \7779 );
buf \U$7404 ( \7781 , \7780 );
xor \U$7405 ( \7782 , \7730 , \7781 );
not \U$7406 ( \7783 , \7782 );
or \U$7407 ( \7784 , \7419 , \7783 );
xor \U$7408 ( \7785 , \7781 , \7729 );
nand \U$7409 ( \7786 , \7785 , \7589 );
nand \U$7410 ( \7787 , \7784 , \7786 );
not \U$7411 ( \7788 , \7667 );
not \U$7412 ( \7789 , \7662 );
or \U$7413 ( \7790 , \7788 , \7789 );
nand \U$7414 ( \7791 , \7652 , \7661 );
nand \U$7415 ( \7792 , \7790 , \7791 );
xor \U$7416 ( \7793 , \1188 , RIae78f80_134);
and \U$7417 ( \7794 , \7793 , \840 );
not \U$7418 ( \7795 , \7607 );
and \U$7419 ( \7796 , \7795 , \797 );
nor \U$7420 ( \7797 , \7794 , \7796 );
not \U$7421 ( \7798 , \7163 );
not \U$7422 ( \7799 , \3147 );
and \U$7423 ( \7800 , \7798 , \7799 );
and \U$7424 ( \7801 , \7631 , \2966 );
nor \U$7425 ( \7802 , \7800 , \7801 );
not \U$7426 ( \7803 , \7802 );
and \U$7427 ( \7804 , \7797 , \7803 );
not \U$7428 ( \7805 , \7797 );
and \U$7429 ( \7806 , \7805 , \7802 );
nor \U$7430 ( \7807 , \7804 , \7806 );
not \U$7431 ( \7808 , \7807 );
and \U$7432 ( \7809 , \7792 , \7808 );
not \U$7433 ( \7810 , \7792 );
and \U$7434 ( \7811 , \7810 , \7807 );
nor \U$7435 ( \7812 , \7809 , \7811 );
not \U$7436 ( \7813 , \7671 );
not \U$7437 ( \7814 , \7642 );
or \U$7438 ( \7815 , \7813 , \7814 );
nand \U$7439 ( \7816 , \7641 , \7617 );
nand \U$7440 ( \7817 , \7815 , \7816 );
xor \U$7441 ( \7818 , \7812 , \7817 );
not \U$7442 ( \7819 , \7748 );
not \U$7443 ( \7820 , \7819 );
not \U$7444 ( \7821 , \7759 );
or \U$7445 ( \7822 , \7820 , \7821 );
nand \U$7446 ( \7823 , \7755 , \7505 );
nand \U$7447 ( \7824 , \7822 , \7823 );
xnor \U$7448 ( \7825 , \7818 , \7824 );
not \U$7449 ( \7826 , \7742 );
not \U$7450 ( \7827 , \7770 );
or \U$7451 ( \7828 , \7826 , \7827 );
nand \U$7452 ( \7829 , \7763 , \7769 );
nand \U$7453 ( \7830 , \7828 , \7829 );
xor \U$7454 ( \7831 , \7825 , \7830 );
and \U$7455 ( \7832 , \1286 , \1879 );
not \U$7456 ( \7833 , \1286 );
and \U$7457 ( \7834 , \7833 , \4458 );
nor \U$7458 ( \7835 , \7832 , \7834 );
or \U$7459 ( \7836 , \7835 , \1029 );
or \U$7460 ( \7837 , \7659 , \3520 );
nand \U$7461 ( \7838 , \7836 , \7837 );
and \U$7462 ( \7839 , \997 , \858 );
not \U$7463 ( \7840 , \997 );
and \U$7464 ( \7841 , \7840 , \857 );
nor \U$7465 ( \7842 , \7839 , \7841 );
or \U$7466 ( \7843 , \7842 , \1210 );
or \U$7467 ( \7844 , \7720 , \6611 );
nand \U$7468 ( \7845 , \7843 , \7844 );
xor \U$7469 ( \7846 , \7838 , \7845 );
and \U$7470 ( \7847 , RIae78b48_125, \6668 );
not \U$7471 ( \7848 , RIae78b48_125);
and \U$7472 ( \7849 , \7848 , \6665 );
nor \U$7473 ( \7850 , \7847 , \7849 );
or \U$7474 ( \7851 , \7850 , \1959 );
or \U$7475 ( \7852 , \7649 , \1976 );
nand \U$7476 ( \7853 , \7851 , \7852 );
xnor \U$7477 ( \7854 , \7846 , \7853 );
not \U$7478 ( \7855 , \7854 );
and \U$7479 ( \7856 , \1143 , RIae793b8_143);
and \U$7480 ( \7857 , \1147 , \1902 );
nor \U$7481 ( \7858 , \7856 , \7857 );
or \U$7482 ( \7859 , \7858 , \3494 );
or \U$7483 ( \7860 , \7620 , \6846 );
nand \U$7484 ( \7861 , \7859 , \7860 );
and \U$7485 ( \7862 , RIae78b48_125, \4081 );
not \U$7486 ( \7863 , \1473 );
xor \U$7487 ( \7864 , RIae79070_136, \7863 );
or \U$7488 ( \7865 , \7864 , \1203 );
or \U$7489 ( \7866 , \1249 , \7704 );
nand \U$7490 ( \7867 , \7865 , \7866 );
xor \U$7491 ( \7868 , \7862 , \7867 );
xor \U$7492 ( \7869 , \7861 , \7868 );
not \U$7493 ( \7870 , \7869 );
or \U$7494 ( \7871 , \7855 , \7870 );
or \U$7495 ( \7872 , \7869 , \7854 );
nand \U$7496 ( \7873 , \7871 , \7872 );
and \U$7497 ( \7874 , \7558 , \1503 );
and \U$7498 ( \7875 , \6913 , RIae79250_140);
nor \U$7499 ( \7876 , \7874 , \7875 );
and \U$7500 ( \7877 , \7876 , \1501 );
and \U$7501 ( \7878 , \7593 , \2650 );
nor \U$7502 ( \7879 , \7877 , \7878 );
not \U$7503 ( \7880 , \4344 );
not \U$7504 ( \7881 , \7663 );
or \U$7505 ( \7882 , \7880 , \7881 );
and \U$7506 ( \7883 , RIae79610_148, \3431 );
not \U$7507 ( \7884 , RIae79610_148);
and \U$7508 ( \7885 , \7884 , \830 );
nor \U$7509 ( \7886 , \7883 , \7885 );
not \U$7510 ( \7887 , \2011 );
or \U$7511 ( \7888 , \7886 , \7887 );
nand \U$7512 ( \7889 , \7882 , \7888 );
and \U$7513 ( \7890 , \7879 , \7889 );
not \U$7514 ( \7891 , \7879 );
not \U$7515 ( \7892 , \7889 );
and \U$7516 ( \7893 , \7891 , \7892 );
nor \U$7517 ( \7894 , \7890 , \7893 );
and \U$7518 ( \7895 , \2027 , RIae78e90_132);
and \U$7519 ( \7896 , \5137 , \1066 );
nor \U$7520 ( \7897 , \7895 , \7896 );
not \U$7521 ( \7898 , \7897 );
and \U$7522 ( \7899 , \7898 , \1322 );
and \U$7523 ( \7900 , \7601 , \1087 );
nor \U$7524 ( \7901 , \7899 , \7900 );
xor \U$7525 ( \7902 , \7894 , \7901 );
xnor \U$7526 ( \7903 , \7873 , \7902 );
nand \U$7527 ( \7904 , \7696 , \7723 );
not \U$7528 ( \7905 , \7692 );
nand \U$7529 ( \7906 , \7905 , \7686 );
and \U$7530 ( \7907 , \7904 , \7906 );
not \U$7531 ( \7908 , \7722 );
not \U$7532 ( \7909 , \7713 );
or \U$7533 ( \7910 , \7908 , \7909 );
nand \U$7534 ( \7911 , \7707 , \7708 );
nand \U$7535 ( \7912 , \7910 , \7911 );
not \U$7536 ( \7913 , \7623 );
not \U$7537 ( \7914 , \7640 );
or \U$7538 ( \7915 , \7913 , \7914 );
or \U$7539 ( \7916 , \7638 , \7625 );
nand \U$7540 ( \7917 , \7915 , \7916 );
and \U$7541 ( \7918 , \7912 , \7917 );
not \U$7542 ( \7919 , \7912 );
not \U$7543 ( \7920 , \7917 );
and \U$7544 ( \7921 , \7919 , \7920 );
nor \U$7545 ( \7922 , \7918 , \7921 );
not \U$7546 ( \7923 , \7613 );
or \U$7547 ( \7924 , \7923 , \7596 );
or \U$7548 ( \7925 , \7612 , \7603 );
nand \U$7549 ( \7926 , \7924 , \7925 );
and \U$7550 ( \7927 , \7922 , \7926 );
not \U$7551 ( \7928 , \7922 );
not \U$7552 ( \7929 , \7926 );
and \U$7553 ( \7930 , \7928 , \7929 );
nor \U$7554 ( \7931 , \7927 , \7930 );
not \U$7555 ( \7932 , \7931 );
and \U$7556 ( \7933 , \7907 , \7932 );
not \U$7557 ( \7934 , \7907 );
and \U$7558 ( \7935 , \7934 , \7931 );
nor \U$7559 ( \7936 , \7933 , \7935 );
not \U$7560 ( \7937 , \7936 );
xor \U$7561 ( \7938 , \7903 , \7937 );
xnor \U$7562 ( \7939 , \7831 , \7938 );
not \U$7563 ( \7940 , \7939 );
not \U$7564 ( \7941 , \7676 );
not \U$7565 ( \7942 , \7681 );
not \U$7566 ( \7943 , \7728 );
or \U$7567 ( \7944 , \7942 , \7943 );
or \U$7568 ( \7945 , \7728 , \7681 );
nand \U$7569 ( \7946 , \7944 , \7945 );
not \U$7570 ( \7947 , \7946 );
or \U$7571 ( \7948 , \7941 , \7947 );
not \U$7572 ( \7949 , \7681 );
nand \U$7573 ( \7950 , \7949 , \7728 );
nand \U$7574 ( \7951 , \7948 , \7950 );
not \U$7575 ( \7952 , \7951 );
not \U$7576 ( \7953 , \7952 );
not \U$7577 ( \7954 , \7729 );
not \U$7578 ( \7955 , \7780 );
or \U$7579 ( \7956 , \7954 , \7955 );
not \U$7580 ( \7957 , \7734 );
nand \U$7581 ( \7958 , \7957 , \7776 );
nand \U$7582 ( \7959 , \7956 , \7958 );
not \U$7583 ( \7960 , \7959 );
or \U$7584 ( \7961 , \7953 , \7960 );
or \U$7585 ( \7962 , \7959 , \7952 );
nand \U$7586 ( \7963 , \7961 , \7962 );
not \U$7587 ( \7964 , \7963 );
or \U$7588 ( \7965 , \7940 , \7964 );
or \U$7589 ( \7966 , \7939 , \7963 );
nand \U$7590 ( \7967 , \7965 , \7966 );
nor \U$7591 ( \7968 , \7787 , \7967 );
not \U$7592 ( \7969 , \7968 );
xor \U$7593 ( \7970 , \7418 , \7782 );
and \U$7594 ( \7971 , \7585 , \7459 );
not \U$7595 ( \7972 , \7585 );
not \U$7596 ( \7973 , \7459 );
and \U$7597 ( \7974 , \7972 , \7973 );
nor \U$7598 ( \7975 , \7971 , \7974 );
not \U$7599 ( \7976 , \7975 );
not \U$7600 ( \7977 , \7239 );
nand \U$7601 ( \7978 , \7977 , \7417 );
xor \U$7602 ( \7979 , \7978 , \7414 );
xor \U$7603 ( \7980 , \7976 , \7979 );
not \U$7604 ( \7981 , \7453 );
not \U$7605 ( \7982 , \7425 );
and \U$7606 ( \7983 , \7981 , \7982 );
and \U$7607 ( \7984 , \7453 , \7425 );
nor \U$7608 ( \7985 , \7983 , \7984 );
not \U$7609 ( \7986 , \7985 );
xor \U$7610 ( \7987 , \6963 , \7082 );
not \U$7611 ( \7988 , \7987 );
not \U$7612 ( \7989 , \7988 );
or \U$7613 ( \7990 , \7986 , \7989 );
not \U$7614 ( \7991 , \7349 );
not \U$7615 ( \7992 , \7365 );
or \U$7616 ( \7993 , \7991 , \7992 );
or \U$7617 ( \7994 , \7365 , \7349 );
nand \U$7618 ( \7995 , \7993 , \7994 );
and \U$7619 ( \7996 , \7405 , \7995 );
not \U$7620 ( \7997 , \7405 );
not \U$7621 ( \7998 , \7995 );
and \U$7622 ( \7999 , \7997 , \7998 );
nor \U$7623 ( \8000 , \7996 , \7999 );
not \U$7624 ( \8001 , \8000 );
xnor \U$7625 ( \8002 , \6958 , \6864 );
nand \U$7626 ( \8003 , \8001 , \8002 );
not \U$7627 ( \8004 , \8003 );
xor \U$7628 ( \8005 , \7396 , \7384 );
not \U$7629 ( \8006 , \8005 );
xor \U$7630 ( \8007 , \6774 , \6780 );
and \U$7631 ( \8008 , \8007 , \6787 );
and \U$7632 ( \8009 , \6774 , \6780 );
nor \U$7633 ( \8010 , \8008 , \8009 );
not \U$7634 ( \8011 , \8010 );
xor \U$7635 ( \8012 , \6792 , \6803 );
and \U$7636 ( \8013 , \8012 , \6809 );
and \U$7637 ( \8014 , \6792 , \6803 );
nor \U$7638 ( \8015 , \8013 , \8014 );
not \U$7639 ( \8016 , \8015 );
not \U$7640 ( \8017 , \8016 );
or \U$7641 ( \8018 , \8011 , \8017 );
or \U$7642 ( \8019 , \8016 , \8010 );
nand \U$7643 ( \8020 , \8018 , \8019 );
not \U$7644 ( \8021 , \8020 );
or \U$7645 ( \8022 , \8006 , \8021 );
not \U$7646 ( \8023 , \8010 );
nand \U$7647 ( \8024 , \8023 , \8016 );
nand \U$7648 ( \8025 , \8022 , \8024 );
not \U$7649 ( \8026 , \8025 );
or \U$7650 ( \8027 , \8004 , \8026 );
not \U$7651 ( \8028 , \8002 );
nand \U$7652 ( \8029 , \8028 , \8000 );
nand \U$7653 ( \8030 , \8027 , \8029 );
nand \U$7654 ( \8031 , \7990 , \8030 );
not \U$7655 ( \8032 , \7985 );
nand \U$7656 ( \8033 , \7987 , \8032 );
and \U$7657 ( \8034 , \8031 , \8033 );
and \U$7658 ( \8035 , \7980 , \8034 );
and \U$7659 ( \8036 , \7976 , \7979 );
nor \U$7660 ( \8037 , \8035 , \8036 );
or \U$7661 ( \8038 , \7970 , \8037 );
not \U$7662 ( \8039 , \7938 );
not \U$7663 ( \8040 , \7831 );
or \U$7664 ( \8041 , \8039 , \8040 );
nand \U$7665 ( \8042 , \7830 , \7825 );
nand \U$7666 ( \8043 , \8041 , \8042 );
not \U$7667 ( \8044 , \8043 );
and \U$7668 ( \8045 , RIae78f80_134, \7702 );
not \U$7669 ( \8046 , RIae78f80_134);
not \U$7670 ( \8047 , \979 );
and \U$7671 ( \8048 , \8046 , \8047 );
nor \U$7672 ( \8049 , \8045 , \8048 );
and \U$7673 ( \8050 , \8049 , \840 );
and \U$7674 ( \8051 , \7793 , \797 );
nor \U$7675 ( \8052 , \8050 , \8051 );
not \U$7676 ( \8053 , \8052 );
not \U$7677 ( \8054 , \7864 );
nand \U$7678 ( \8055 , \8054 , \1062 );
and \U$7679 ( \8056 , \1039 , \883 );
not \U$7680 ( \8057 , \1039 );
and \U$7681 ( \8058 , \8057 , \879 );
nor \U$7682 ( \8059 , \8056 , \8058 );
not \U$7683 ( \8060 , \8059 );
nand \U$7684 ( \8061 , \8060 , \1049 );
nand \U$7685 ( \8062 , \8055 , \8061 );
xnor \U$7686 ( \8063 , \8062 , \7802 );
not \U$7687 ( \8064 , \8063 );
and \U$7688 ( \8065 , \8053 , \8064 );
and \U$7689 ( \8066 , \8052 , \8063 );
nor \U$7690 ( \8067 , \8065 , \8066 );
not \U$7691 ( \8068 , \8067 );
not \U$7692 ( \8069 , \7807 );
not \U$7693 ( \8070 , \7792 );
or \U$7694 ( \8071 , \8069 , \8070 );
not \U$7695 ( \8072 , \7797 );
nand \U$7696 ( \8073 , \8072 , \7802 );
nand \U$7697 ( \8074 , \8071 , \8073 );
not \U$7698 ( \8075 , \8074 );
or \U$7699 ( \8076 , \8068 , \8075 );
or \U$7700 ( \8077 , \8067 , \8074 );
nand \U$7701 ( \8078 , \8076 , \8077 );
not \U$7702 ( \8079 , \7926 );
not \U$7703 ( \8080 , \7922 );
or \U$7704 ( \8081 , \8079 , \8080 );
nand \U$7705 ( \8082 , \7912 , \7917 );
nand \U$7706 ( \8083 , \8081 , \8082 );
xor \U$7707 ( \8084 , \8078 , \8083 );
not \U$7708 ( \8085 , \7817 );
not \U$7709 ( \8086 , \7812 );
not \U$7710 ( \8087 , \7824 );
or \U$7711 ( \8088 , \8086 , \8087 );
or \U$7712 ( \8089 , \7824 , \7812 );
nand \U$7713 ( \8090 , \8088 , \8089 );
not \U$7714 ( \8091 , \8090 );
or \U$7715 ( \8092 , \8085 , \8091 );
not \U$7716 ( \8093 , \7812 );
nand \U$7717 ( \8094 , \8093 , \7824 );
nand \U$7718 ( \8095 , \8092 , \8094 );
xor \U$7719 ( \8096 , \8084 , \8095 );
or \U$7720 ( \8097 , \7894 , \7901 );
or \U$7721 ( \8098 , \7892 , \7879 );
nand \U$7722 ( \8099 , \8097 , \8098 );
not \U$7723 ( \8100 , \8099 );
not \U$7724 ( \8101 , \8100 );
and \U$7725 ( \8102 , \7846 , \7853 );
and \U$7726 ( \8103 , \7838 , \7845 );
nor \U$7727 ( \8104 , \8102 , \8103 );
not \U$7728 ( \8105 , \8104 );
not \U$7729 ( \8106 , \7861 );
not \U$7730 ( \8107 , \7868 );
or \U$7731 ( \8108 , \8106 , \8107 );
nand \U$7732 ( \8109 , \7862 , \7867 );
nand \U$7733 ( \8110 , \8108 , \8109 );
not \U$7734 ( \8111 , \8110 );
or \U$7735 ( \8112 , \8105 , \8111 );
or \U$7736 ( \8113 , \8110 , \8104 );
nand \U$7737 ( \8114 , \8112 , \8113 );
not \U$7738 ( \8115 , \8114 );
or \U$7739 ( \8116 , \8101 , \8115 );
or \U$7740 ( \8117 , \8114 , \8100 );
nand \U$7741 ( \8118 , \8116 , \8117 );
not \U$7742 ( \8119 , \8118 );
not \U$7743 ( \8120 , \7902 );
not \U$7744 ( \8121 , \7873 );
or \U$7745 ( \8122 , \8120 , \8121 );
not \U$7746 ( \8123 , \7854 );
nand \U$7747 ( \8124 , \8123 , \7869 );
nand \U$7748 ( \8125 , \8122 , \8124 );
not \U$7749 ( \8126 , \8125 );
not \U$7750 ( \8127 , \8126 );
or \U$7751 ( \8128 , \8119 , \8127 );
or \U$7752 ( \8129 , \8118 , \8126 );
nand \U$7753 ( \8130 , \8128 , \8129 );
not \U$7754 ( \8131 , \1074 );
and \U$7755 ( \8132 , RIae78e90_132, \1406 );
not \U$7756 ( \8133 , RIae78e90_132);
and \U$7757 ( \8134 , \8133 , \3688 );
nor \U$7758 ( \8135 , \8132 , \8134 );
not \U$7759 ( \8136 , \8135 );
or \U$7760 ( \8137 , \8131 , \8136 );
or \U$7761 ( \8138 , \7897 , \1413 );
nand \U$7762 ( \8139 , \8137 , \8138 );
and \U$7763 ( \8140 , \1286 , \2050 );
not \U$7764 ( \8141 , \1286 );
and \U$7765 ( \8142 , \8141 , \2049 );
nor \U$7766 ( \8143 , \8140 , \8142 );
not \U$7767 ( \8144 , \1027 );
or \U$7768 ( \8145 , \8143 , \8144 );
not \U$7769 ( \8146 , \952 );
or \U$7770 ( \8147 , \7835 , \8146 );
nand \U$7771 ( \8148 , \8145 , \8147 );
xor \U$7772 ( \8149 , \8139 , \8148 );
not \U$7773 ( \8150 , \7842 );
not \U$7774 ( \8151 , \7429 );
and \U$7775 ( \8152 , \8150 , \8151 );
and \U$7776 ( \8153 , RIae79160_138, \941 );
not \U$7777 ( \8154 , RIae79160_138);
and \U$7778 ( \8155 , \8154 , \940 );
nor \U$7779 ( \8156 , \8153 , \8155 );
and \U$7780 ( \8157 , \8156 , \1013 );
nor \U$7781 ( \8158 , \8152 , \8157 );
not \U$7782 ( \8159 , \8158 );
xor \U$7783 ( \8160 , \8149 , \8159 );
and \U$7784 ( \8161 , \7575 , \7163 );
nor \U$7785 ( \8162 , \8161 , \3147 );
not \U$7786 ( \8163 , \8162 );
not \U$7787 ( \8164 , \2011 );
not \U$7788 ( \8165 , RIae79610_148);
not \U$7789 ( \8166 , \994 );
or \U$7790 ( \8167 , \8165 , \8166 );
or \U$7791 ( \8168 , \992 , RIae79610_148);
nand \U$7792 ( \8169 , \8167 , \8168 );
not \U$7793 ( \8170 , \8169 );
not \U$7794 ( \8171 , \8170 );
or \U$7795 ( \8172 , \8164 , \8171 );
not \U$7796 ( \8173 , \7886 );
nand \U$7797 ( \8174 , \8173 , \2063 );
nand \U$7798 ( \8175 , \8172 , \8174 );
not \U$7799 ( \8176 , \8175 );
or \U$7800 ( \8177 , \8163 , \8176 );
or \U$7801 ( \8178 , \8175 , \8162 );
nand \U$7802 ( \8179 , \8177 , \8178 );
and \U$7803 ( \8180 , RIae79250_140, \1291 );
not \U$7804 ( \8181 , RIae79250_140);
and \U$7805 ( \8182 , \8181 , \1290 );
nor \U$7806 ( \8183 , \8180 , \8182 );
and \U$7807 ( \8184 , \8183 , \1501 );
and \U$7808 ( \8185 , \7876 , \1499 );
nor \U$7809 ( \8186 , \8184 , \8185 );
not \U$7810 ( \8187 , \8186 );
and \U$7811 ( \8188 , \8179 , \8187 );
not \U$7812 ( \8189 , \8179 );
and \U$7813 ( \8190 , \8189 , \8186 );
nor \U$7814 ( \8191 , \8188 , \8190 );
xor \U$7815 ( \8192 , \8160 , \8191 );
not \U$7816 ( \8193 , \1864 );
and \U$7817 ( \8194 , RIae793b8_143, \782 );
not \U$7818 ( \8195 , RIae793b8_143);
and \U$7819 ( \8196 , \8195 , \783 );
nor \U$7820 ( \8197 , \8194 , \8196 );
not \U$7821 ( \8198 , \8197 );
or \U$7822 ( \8199 , \8193 , \8198 );
or \U$7823 ( \8200 , \7858 , \6846 );
nand \U$7824 ( \8201 , \8199 , \8200 );
not \U$7825 ( \8202 , \868 );
and \U$7826 ( \8203 , RIae78b48_125, \1899 );
not \U$7827 ( \8204 , RIae78b48_125);
and \U$7828 ( \8205 , \8204 , \3785 );
nor \U$7829 ( \8206 , \8203 , \8205 );
not \U$7830 ( \8207 , \8206 );
or \U$7831 ( \8208 , \8202 , \8207 );
or \U$7832 ( \8209 , \7850 , \1976 );
nand \U$7833 ( \8210 , \8208 , \8209 );
and \U$7834 ( \8211 , \2231 , RIae78b48_125);
xor \U$7835 ( \8212 , \8210 , \8211 );
xor \U$7836 ( \8213 , \8201 , \8212 );
xor \U$7837 ( \8214 , \8192 , \8213 );
xor \U$7838 ( \8215 , \8130 , \8214 );
xnor \U$7839 ( \8216 , \8096 , \8215 );
not \U$7840 ( \8217 , \7936 );
or \U$7841 ( \8218 , \8217 , \7903 );
or \U$7842 ( \8219 , \7907 , \7932 );
nand \U$7843 ( \8220 , \8218 , \8219 );
xor \U$7844 ( \8221 , \8216 , \8220 );
not \U$7845 ( \8222 , \8221 );
or \U$7846 ( \8223 , \8044 , \8222 );
or \U$7847 ( \8224 , \8221 , \8043 );
nand \U$7848 ( \8225 , \8223 , \8224 );
not \U$7849 ( \8226 , \8225 );
not \U$7850 ( \8227 , \7939 );
nand \U$7851 ( \8228 , \8227 , \7963 );
nand \U$7852 ( \8229 , \7959 , \7951 );
nand \U$7853 ( \8230 , \8226 , \8228 , \8229 );
not \U$7854 ( \8231 , \8043 );
or \U$7855 ( \8232 , \8221 , \8231 );
not \U$7856 ( \8233 , \8214 );
not \U$7857 ( \8234 , \8130 );
or \U$7858 ( \8235 , \8233 , \8234 );
nand \U$7859 ( \8236 , \8118 , \8125 );
nand \U$7860 ( \8237 , \8235 , \8236 );
not \U$7861 ( \8238 , \8237 );
not \U$7862 ( \8239 , \8078 );
not \U$7863 ( \8240 , \8083 );
or \U$7864 ( \8241 , \8239 , \8240 );
not \U$7865 ( \8242 , \8067 );
nand \U$7866 ( \8243 , \8242 , \8074 );
nand \U$7867 ( \8244 , \8241 , \8243 );
not \U$7868 ( \8245 , \8244 );
not \U$7869 ( \8246 , \8245 );
not \U$7870 ( \8247 , \8099 );
not \U$7871 ( \8248 , \8114 );
or \U$7872 ( \8249 , \8247 , \8248 );
not \U$7873 ( \8250 , \8104 );
nand \U$7874 ( \8251 , \8250 , \8110 );
nand \U$7875 ( \8252 , \8249 , \8251 );
not \U$7876 ( \8253 , \7803 );
not \U$7877 ( \8254 , \8062 );
or \U$7878 ( \8255 , \8253 , \8254 );
not \U$7879 ( \8256 , \8052 );
nand \U$7880 ( \8257 , \8256 , \8063 );
nand \U$7881 ( \8258 , \8255 , \8257 );
not \U$7882 ( \8259 , \8258 );
not \U$7883 ( \8260 , \1074 );
and \U$7884 ( \8261 , RIae78e90_132, \1188 );
not \U$7885 ( \8262 , RIae78e90_132);
and \U$7886 ( \8263 , \8262 , \1187 );
nor \U$7887 ( \8264 , \8261 , \8263 );
not \U$7888 ( \8265 , \8264 );
or \U$7889 ( \8266 , \8260 , \8265 );
nand \U$7890 ( \8267 , \8135 , \1259 );
nand \U$7891 ( \8268 , \8266 , \8267 );
and \U$7892 ( \8269 , RIae78f80_134, \1473 );
not \U$7893 ( \8270 , RIae78f80_134);
and \U$7894 ( \8271 , \8270 , \1472 );
nor \U$7895 ( \8272 , \8269 , \8271 );
not \U$7896 ( \8273 , \8272 );
not \U$7897 ( \8274 , \8273 );
not \U$7898 ( \8275 , \1227 );
and \U$7899 ( \8276 , \8274 , \8275 );
and \U$7900 ( \8277 , \8049 , \797 );
nor \U$7901 ( \8278 , \8276 , \8277 );
xnor \U$7902 ( \8279 , \8268 , \8278 );
and \U$7903 ( \8280 , \1503 , \1146 );
not \U$7904 ( \8281 , \1503 );
and \U$7905 ( \8282 , \8281 , \1147 );
nor \U$7906 ( \8283 , \8280 , \8282 );
and \U$7907 ( \8284 , \8283 , \1501 );
and \U$7908 ( \8285 , \8183 , \1499 );
nor \U$7909 ( \8286 , \8284 , \8285 );
and \U$7910 ( \8287 , \8279 , \8286 );
not \U$7911 ( \8288 , \8279 );
not \U$7912 ( \8289 , \8286 );
and \U$7913 ( \8290 , \8288 , \8289 );
nor \U$7914 ( \8291 , \8287 , \8290 );
not \U$7915 ( \8292 , \8291 );
and \U$7916 ( \8293 , \8259 , \8292 );
and \U$7917 ( \8294 , \8258 , \8291 );
nor \U$7918 ( \8295 , \8293 , \8294 );
xnor \U$7919 ( \8296 , \8252 , \8295 );
not \U$7920 ( \8297 , \8296 );
or \U$7921 ( \8298 , \8246 , \8297 );
or \U$7922 ( \8299 , \8296 , \8245 );
nand \U$7923 ( \8300 , \8298 , \8299 );
not \U$7924 ( \8301 , \8300 );
not \U$7925 ( \8302 , \8301 );
or \U$7926 ( \8303 , \8238 , \8302 );
not \U$7927 ( \8304 , \8237 );
nand \U$7928 ( \8305 , \8304 , \8300 );
nand \U$7929 ( \8306 , \8303 , \8305 );
xor \U$7930 ( \8307 , \8139 , \8148 );
not \U$7931 ( \8308 , \8158 );
and \U$7932 ( \8309 , \8307 , \8308 );
and \U$7933 ( \8310 , \8139 , \8148 );
or \U$7934 ( \8311 , \8309 , \8310 );
not \U$7935 ( \8312 , \8311 );
not \U$7936 ( \8313 , \8162 );
not \U$7937 ( \8314 , \8313 );
not \U$7938 ( \8315 , \8175 );
or \U$7939 ( \8316 , \8314 , \8315 );
nand \U$7940 ( \8317 , \8179 , \8187 );
nand \U$7941 ( \8318 , \8316 , \8317 );
not \U$7942 ( \8319 , \8169 );
not \U$7943 ( \8320 , \2063 );
not \U$7944 ( \8321 , \8320 );
and \U$7945 ( \8322 , \8319 , \8321 );
and \U$7946 ( \8323 , \2011 , RIae79610_148);
nor \U$7947 ( \8324 , \8322 , \8323 );
not \U$7948 ( \8325 , \8324 );
and \U$7949 ( \8326 , \8318 , \8325 );
not \U$7950 ( \8327 , \8318 );
and \U$7951 ( \8328 , \8327 , \8324 );
or \U$7952 ( \8329 , \8326 , \8328 );
xnor \U$7953 ( \8330 , \8312 , \8329 );
xor \U$7954 ( \8331 , \8160 , \8191 );
and \U$7955 ( \8332 , \8331 , \8213 );
and \U$7956 ( \8333 , \8160 , \8191 );
or \U$7957 ( \8334 , \8332 , \8333 );
xor \U$7958 ( \8335 , \8330 , \8334 );
not \U$7959 ( \8336 , \1049 );
and \U$7960 ( \8337 , \1024 , \1039 );
not \U$7961 ( \8338 , \1024 );
and \U$7962 ( \8339 , \8338 , RIae79070_136);
nor \U$7963 ( \8340 , \8337 , \8339 );
not \U$7964 ( \8341 , \8340 );
or \U$7965 ( \8342 , \8336 , \8341 );
or \U$7966 ( \8343 , \8059 , \1249 );
nand \U$7967 ( \8344 , \8342 , \8343 );
and \U$7968 ( \8345 , \6665 , RIae78b48_125);
xnor \U$7969 ( \8346 , \8344 , \8345 );
xnor \U$7970 ( \8347 , \3431 , RIae793b8_143);
and \U$7971 ( \8348 , \8347 , \1864 );
and \U$7972 ( \8349 , \8197 , \1910 );
nor \U$7973 ( \8350 , \8348 , \8349 );
xnor \U$7974 ( \8351 , \8346 , \8350 );
not \U$7975 ( \8352 , \8351 );
and \U$7976 ( \8353 , \3443 , RIae79160_138);
not \U$7977 ( \8354 , \3443 );
and \U$7978 ( \8355 , \8354 , \997 );
nor \U$7979 ( \8356 , \8353 , \8355 );
not \U$7980 ( \8357 , \8356 );
not \U$7981 ( \8358 , \1013 );
not \U$7982 ( \8359 , \8358 );
and \U$7983 ( \8360 , \8357 , \8359 );
and \U$7984 ( \8361 , \8156 , \1430 );
nor \U$7985 ( \8362 , \8360 , \8361 );
not \U$7986 ( \8363 , \8143 );
not \U$7987 ( \8364 , \8146 );
and \U$7988 ( \8365 , \8363 , \8364 );
xnor \U$7989 ( \8366 , \2027 , RIae78bc0_126);
and \U$7990 ( \8367 , \8366 , \1027 );
nor \U$7991 ( \8368 , \8365 , \8367 );
xor \U$7992 ( \8369 , \8362 , \8368 );
xor \U$7993 ( \8370 , RIae78b48_125, \6855 );
and \U$7994 ( \8371 , \8370 , \868 );
and \U$7995 ( \8372 , \8206 , \1129 );
nor \U$7996 ( \8373 , \8371 , \8372 );
xor \U$7997 ( \8374 , \8369 , \8373 );
not \U$7998 ( \8375 , \8374 );
not \U$7999 ( \8376 , \8201 );
not \U$8000 ( \8377 , \8212 );
or \U$8001 ( \8378 , \8376 , \8377 );
nand \U$8002 ( \8379 , \8210 , \8211 );
nand \U$8003 ( \8380 , \8378 , \8379 );
not \U$8004 ( \8381 , \8380 );
or \U$8005 ( \8382 , \8375 , \8381 );
or \U$8006 ( \8383 , \8380 , \8374 );
nand \U$8007 ( \8384 , \8382 , \8383 );
not \U$8008 ( \8385 , \8384 );
or \U$8009 ( \8386 , \8352 , \8385 );
or \U$8010 ( \8387 , \8384 , \8351 );
nand \U$8011 ( \8388 , \8386 , \8387 );
xor \U$8012 ( \8389 , \8335 , \8388 );
and \U$8013 ( \8390 , \8306 , \8389 );
not \U$8014 ( \8391 , \8306 );
not \U$8015 ( \8392 , \8389 );
and \U$8016 ( \8393 , \8391 , \8392 );
nor \U$8017 ( \8394 , \8390 , \8393 );
buf \U$8018 ( \8395 , \8394 );
not \U$8019 ( \8396 , \8395 );
not \U$8020 ( \8397 , \8215 );
not \U$8021 ( \8398 , \8096 );
or \U$8022 ( \8399 , \8397 , \8398 );
nand \U$8023 ( \8400 , \8095 , \8084 );
nand \U$8024 ( \8401 , \8399 , \8400 );
not \U$8025 ( \8402 , \8401 );
not \U$8026 ( \8403 , \8402 );
and \U$8027 ( \8404 , \8396 , \8403 );
and \U$8028 ( \8405 , \8395 , \8402 );
nor \U$8029 ( \8406 , \8404 , \8405 );
not \U$8030 ( \8407 , \8216 );
nand \U$8031 ( \8408 , \8407 , \8220 );
nand \U$8032 ( \8409 , \8232 , \8406 , \8408 );
and \U$8033 ( \8410 , \7969 , \8038 , \8230 , \8409 );
not \U$8034 ( \8411 , \7340 );
not \U$8035 ( \8412 , \7292 );
not \U$8036 ( \8413 , \8412 );
and \U$8037 ( \8414 , \8411 , \8413 );
and \U$8038 ( \8415 , \7340 , \8412 );
nor \U$8039 ( \8416 , \8414 , \8415 );
not \U$8040 ( \8417 , \7304 );
not \U$8041 ( \8418 , \7334 );
not \U$8042 ( \8419 , \8418 );
or \U$8043 ( \8420 , \8417 , \8419 );
or \U$8044 ( \8421 , \8418 , \7304 );
nand \U$8045 ( \8422 , \8420 , \8421 );
not \U$8046 ( \8423 , \8422 );
not \U$8047 ( \8424 , \6638 );
or \U$8048 ( \8425 , \6659 , \6604 );
not \U$8049 ( \8426 , \8425 );
or \U$8050 ( \8427 , \8424 , \8426 );
nand \U$8051 ( \8428 , \6659 , \6604 );
nand \U$8052 ( \8429 , \8427 , \8428 );
not \U$8053 ( \8430 , \8429 );
or \U$8054 ( \8431 , \8423 , \8430 );
not \U$8055 ( \8432 , \8429 );
and \U$8056 ( \8433 , \8422 , \8432 );
not \U$8057 ( \8434 , \8422 );
and \U$8058 ( \8435 , \8434 , \8429 );
nor \U$8059 ( \8436 , \8433 , \8435 );
not \U$8060 ( \8437 , \8436 );
xor \U$8061 ( \8438 , \7269 , \7263 );
xnor \U$8062 ( \8439 , \8438 , \7283 );
nand \U$8063 ( \8440 , \8437 , \8439 );
nand \U$8064 ( \8441 , \8431 , \8440 );
not \U$8065 ( \8442 , \8441 );
xor \U$8066 ( \8443 , \8416 , \8442 );
not \U$8067 ( \8444 , \6730 );
not \U$8068 ( \8445 , \6694 );
not \U$8069 ( \8446 , \8445 );
and \U$8070 ( \8447 , \8444 , \8446 );
and \U$8071 ( \8448 , \6744 , \6734 );
nor \U$8072 ( \8449 , \8447 , \8448 );
not \U$8073 ( \8450 , \6811 );
not \U$8074 ( \8451 , \8450 );
not \U$8075 ( \8452 , \6818 );
and \U$8076 ( \8453 , \8451 , \8452 );
and \U$8077 ( \8454 , \6788 , \6810 );
nor \U$8078 ( \8455 , \8453 , \8454 );
xor \U$8079 ( \8456 , \8449 , \8455 );
xor \U$8080 ( \8457 , \8010 , \8005 );
xnor \U$8081 ( \8458 , \8457 , \8015 );
and \U$8082 ( \8459 , \8456 , \8458 );
and \U$8083 ( \8460 , \8449 , \8455 );
or \U$8084 ( \8461 , \8459 , \8460 );
and \U$8085 ( \8462 , \8443 , \8461 );
and \U$8086 ( \8463 , \8416 , \8442 );
or \U$8087 ( \8464 , \8462 , \8463 );
not \U$8088 ( \8465 , \8464 );
not \U$8089 ( \8466 , \7344 );
not \U$8090 ( \8467 , \8466 );
not \U$8091 ( \8468 , \7410 );
or \U$8092 ( \8469 , \8467 , \8468 );
or \U$8093 ( \8470 , \7410 , \8466 );
nand \U$8094 ( \8471 , \8469 , \8470 );
not \U$8095 ( \8472 , \8471 );
not \U$8096 ( \8473 , \8030 );
not \U$8097 ( \8474 , \8032 );
not \U$8098 ( \8475 , \7988 );
or \U$8099 ( \8476 , \8474 , \8475 );
nand \U$8100 ( \8477 , \7987 , \7985 );
nand \U$8101 ( \8478 , \8476 , \8477 );
not \U$8102 ( \8479 , \8478 );
or \U$8103 ( \8480 , \8473 , \8479 );
or \U$8104 ( \8481 , \8478 , \8030 );
nand \U$8105 ( \8482 , \8480 , \8481 );
not \U$8106 ( \8483 , \8482 );
or \U$8107 ( \8484 , \8472 , \8483 );
or \U$8108 ( \8485 , \8482 , \8471 );
nand \U$8109 ( \8486 , \8484 , \8485 );
not \U$8110 ( \8487 , \8486 );
not \U$8111 ( \8488 , \8487 );
or \U$8112 ( \8489 , \8465 , \8488 );
not \U$8113 ( \8490 , \8464 );
nand \U$8114 ( \8491 , \8490 , \8486 );
nand \U$8115 ( \8492 , \8489 , \8491 );
xor \U$8116 ( \8493 , \8002 , \8000 );
xor \U$8117 ( \8494 , \8493 , \8025 );
and \U$8118 ( \8495 , \6661 , \6745 );
and \U$8119 ( \8496 , \6599 , \6660 );
nor \U$8120 ( \8497 , \8495 , \8496 );
not \U$8121 ( \8498 , \8436 );
not \U$8122 ( \8499 , \8439 );
and \U$8123 ( \8500 , \8498 , \8499 );
and \U$8124 ( \8501 , \8436 , \8439 );
nor \U$8125 ( \8502 , \8500 , \8501 );
xor \U$8126 ( \8503 , \8497 , \8502 );
xor \U$8127 ( \8504 , \8449 , \8455 );
xor \U$8128 ( \8505 , \8504 , \8458 );
and \U$8129 ( \8506 , \8503 , \8505 );
and \U$8130 ( \8507 , \8497 , \8502 );
or \U$8131 ( \8508 , \8506 , \8507 );
xor \U$8132 ( \8509 , \8494 , \8508 );
xor \U$8133 ( \8510 , \8416 , \8442 );
xor \U$8134 ( \8511 , \8510 , \8461 );
and \U$8135 ( \8512 , \8509 , \8511 );
and \U$8136 ( \8513 , \8494 , \8508 );
or \U$8137 ( \8514 , \8512 , \8513 );
nand \U$8138 ( \8515 , \8492 , \8514 );
xor \U$8139 ( \8516 , \7975 , \8034 );
xnor \U$8140 ( \8517 , \8516 , \7979 );
not \U$8141 ( \8518 , \8464 );
not \U$8142 ( \8519 , \8486 );
or \U$8143 ( \8520 , \8518 , \8519 );
not \U$8144 ( \8521 , \8471 );
nand \U$8145 ( \8522 , \8521 , \8482 );
nand \U$8146 ( \8523 , \8520 , \8522 );
nand \U$8147 ( \8524 , \8517 , \8523 );
and \U$8148 ( \8525 , \8515 , \8524 );
not \U$8149 ( \8526 , \6758 );
not \U$8150 ( \8527 , \6819 );
or \U$8151 ( \8528 , \8526 , \8527 );
or \U$8152 ( \8529 , \6819 , \6758 );
not \U$8153 ( \8530 , \6767 );
nand \U$8154 ( \8531 , \8529 , \8530 );
nand \U$8155 ( \8532 , \8528 , \8531 );
xor \U$8156 ( \8533 , \6746 , \6750 );
and \U$8157 ( \8534 , \8533 , \6820 );
and \U$8158 ( \8535 , \6746 , \6750 );
or \U$8159 ( \8536 , \8534 , \8535 );
xor \U$8160 ( \8537 , \8532 , \8536 );
xor \U$8161 ( \8538 , \8497 , \8502 );
xor \U$8162 ( \8539 , \8538 , \8505 );
xnor \U$8163 ( \8540 , \8537 , \8539 );
xor \U$8164 ( \8541 , \6592 , \6587 );
or \U$8165 ( \8542 , \8541 , \6821 );
not \U$8166 ( \8543 , \6592 );
nand \U$8167 ( \8544 , \8543 , \6587 );
nand \U$8168 ( \8545 , \8542 , \8544 );
nand \U$8169 ( \8546 , \8540 , \8545 );
not \U$8170 ( \8547 , \8536 );
not \U$8171 ( \8548 , \8547 );
not \U$8172 ( \8549 , \8532 );
not \U$8173 ( \8550 , \8549 );
not \U$8174 ( \8551 , \8539 );
or \U$8175 ( \8552 , \8550 , \8551 );
or \U$8176 ( \8553 , \8539 , \8549 );
nand \U$8177 ( \8554 , \8552 , \8553 );
not \U$8178 ( \8555 , \8554 );
or \U$8179 ( \8556 , \8548 , \8555 );
nand \U$8180 ( \8557 , \8539 , \8532 );
nand \U$8181 ( \8558 , \8556 , \8557 );
xor \U$8182 ( \8559 , \8494 , \8508 );
xor \U$8183 ( \8560 , \8559 , \8511 );
nand \U$8184 ( \8561 , \8558 , \8560 );
buf \U$8185 ( \8562 , \8561 );
and \U$8186 ( \8563 , \8525 , \8546 , \8562 );
nand \U$8187 ( \8564 , \8410 , \8563 );
not \U$8188 ( \8565 , \8564 );
not \U$8189 ( \8566 , \8237 );
not \U$8190 ( \8567 , \8300 );
or \U$8191 ( \8568 , \8566 , \8567 );
not \U$8192 ( \8569 , \8245 );
nand \U$8193 ( \8570 , \8569 , \8296 );
nand \U$8194 ( \8571 , \8568 , \8570 );
not \U$8195 ( \8572 , \8571 );
not \U$8196 ( \8573 , \8324 );
not \U$8197 ( \8574 , \8318 );
or \U$8198 ( \8575 , \8573 , \8574 );
not \U$8199 ( \8576 , \8312 );
nand \U$8200 ( \8577 , \8576 , \8329 );
nand \U$8201 ( \8578 , \8575 , \8577 );
not \U$8202 ( \8579 , \8380 );
and \U$8203 ( \8580 , \8579 , \8351 );
nor \U$8204 ( \8581 , \8580 , \8374 );
nor \U$8205 ( \8582 , \8579 , \8351 );
nor \U$8206 ( \8583 , \8581 , \8582 );
xor \U$8207 ( \8584 , \8578 , \8583 );
not \U$8208 ( \8585 , \8346 );
not \U$8209 ( \8586 , \8350 );
and \U$8210 ( \8587 , \8585 , \8586 );
and \U$8211 ( \8588 , \8344 , \8345 );
nor \U$8212 ( \8589 , \8587 , \8588 );
not \U$8213 ( \8590 , \8589 );
not \U$8214 ( \8591 , \8289 );
not \U$8215 ( \8592 , \8279 );
or \U$8216 ( \8593 , \8591 , \8592 );
not \U$8217 ( \8594 , \8278 );
nand \U$8218 ( \8595 , \8594 , \8268 );
nand \U$8219 ( \8596 , \8593 , \8595 );
not \U$8220 ( \8597 , \8596 );
or \U$8221 ( \8598 , \8590 , \8597 );
or \U$8222 ( \8599 , \8596 , \8589 );
nand \U$8223 ( \8600 , \8598 , \8599 );
nand \U$8224 ( \8601 , \1899 , RIae78b48_125);
xor \U$8225 ( \8602 , \3814 , RIae79250_140);
not \U$8226 ( \8603 , \8602 );
not \U$8227 ( \8604 , \1502 );
and \U$8228 ( \8605 , \8603 , \8604 );
and \U$8229 ( \8606 , \8283 , \1499 );
nor \U$8230 ( \8607 , \8605 , \8606 );
xor \U$8231 ( \8608 , \8601 , \8607 );
xor \U$8232 ( \8609 , \880 , RIae78f80_134);
and \U$8233 ( \8610 , \8609 , \840 );
and \U$8234 ( \8611 , \8272 , \797 );
nor \U$8235 ( \8612 , \8610 , \8611 );
xor \U$8236 ( \8613 , \8608 , \8612 );
not \U$8237 ( \8614 , \8613 );
xnor \U$8238 ( \8615 , \8600 , \8614 );
xor \U$8239 ( \8616 , \8584 , \8615 );
not \U$8240 ( \8617 , \8616 );
not \U$8241 ( \8618 , \8388 );
not \U$8242 ( \8619 , \8335 );
or \U$8243 ( \8620 , \8618 , \8619 );
nand \U$8244 ( \8621 , \8330 , \8334 );
nand \U$8245 ( \8622 , \8620 , \8621 );
not \U$8246 ( \8623 , \8252 );
nor \U$8247 ( \8624 , \8623 , \8295 );
not \U$8248 ( \8625 , \8258 );
nor \U$8249 ( \8626 , \8625 , \8291 );
nor \U$8250 ( \8627 , \8624 , \8626 );
and \U$8251 ( \8628 , \2594 , RIae78b48_125);
and \U$8252 ( \8629 , \2595 , \860 );
nor \U$8253 ( \8630 , \8628 , \8629 );
not \U$8254 ( \8631 , \8630 );
not \U$8255 ( \8632 , \1603 );
and \U$8256 ( \8633 , \8631 , \8632 );
and \U$8257 ( \8634 , \8370 , \1129 );
nor \U$8258 ( \8635 , \8633 , \8634 );
not \U$8259 ( \8636 , \8635 );
and \U$8260 ( \8637 , \1286 , \3688 );
not \U$8261 ( \8638 , \1286 );
and \U$8262 ( \8639 , \8638 , \1406 );
nor \U$8263 ( \8640 , \8637 , \8639 );
and \U$8264 ( \8641 , \8640 , \1028 );
and \U$8265 ( \8642 , \8366 , \953 );
nor \U$8266 ( \8643 , \8641 , \8642 );
not \U$8267 ( \8644 , \8643 );
not \U$8268 ( \8645 , \1062 );
not \U$8269 ( \8646 , \8340 );
or \U$8270 ( \8647 , \8645 , \8646 );
and \U$8271 ( \8648 , \940 , RIae79070_136);
and \U$8272 ( \8649 , \939 , \1039 );
nor \U$8273 ( \8650 , \8648 , \8649 );
or \U$8274 ( \8651 , \8650 , \1203 );
nand \U$8275 ( \8652 , \8647 , \8651 );
not \U$8276 ( \8653 , \8652 );
or \U$8277 ( \8654 , \8644 , \8653 );
or \U$8278 ( \8655 , \8652 , \8643 );
nand \U$8279 ( \8656 , \8654 , \8655 );
not \U$8280 ( \8657 , \8656 );
or \U$8281 ( \8658 , \8636 , \8657 );
or \U$8282 ( \8659 , \8635 , \8656 );
nand \U$8283 ( \8660 , \8658 , \8659 );
not \U$8284 ( \8661 , \8660 );
xor \U$8285 ( \8662 , \1291 , RIae79160_138);
and \U$8286 ( \8663 , \8662 , \1013 );
not \U$8287 ( \8664 , \8356 );
and \U$8288 ( \8665 , \8664 , \1010 );
nor \U$8289 ( \8666 , \8663 , \8665 );
nand \U$8290 ( \8667 , RIae79598_147, RIae79688_149);
and \U$8291 ( \8668 , \8667 , RIae79610_148);
xor \U$8292 ( \8669 , \8666 , \8668 );
not \U$8293 ( \8670 , \1910 );
not \U$8294 ( \8671 , \8347 );
or \U$8295 ( \8672 , \8670 , \8671 );
and \U$8296 ( \8673 , \994 , RIae793b8_143);
not \U$8297 ( \8674 , \994 );
and \U$8298 ( \8675 , \8674 , \1884 );
nor \U$8299 ( \8676 , \8673 , \8675 );
nand \U$8300 ( \8677 , \1864 , \8676 );
nand \U$8301 ( \8678 , \8672 , \8677 );
not \U$8302 ( \8679 , \8678 );
xor \U$8303 ( \8680 , \8669 , \8679 );
not \U$8304 ( \8681 , \8680 );
or \U$8305 ( \8682 , \8661 , \8681 );
or \U$8306 ( \8683 , \8680 , \8660 );
nand \U$8307 ( \8684 , \8682 , \8683 );
xor \U$8308 ( \8685 , \8362 , \8368 );
and \U$8309 ( \8686 , \8685 , \8373 );
and \U$8310 ( \8687 , \8362 , \8368 );
nor \U$8311 ( \8688 , \8686 , \8687 );
xor \U$8312 ( \8689 , RIae78e90_132, \3718 );
and \U$8313 ( \8690 , \8689 , \1074 );
and \U$8314 ( \8691 , \8264 , \1087 );
nor \U$8315 ( \8692 , \8690 , \8691 );
and \U$8316 ( \8693 , \8692 , \8324 );
not \U$8317 ( \8694 , \8692 );
and \U$8318 ( \8695 , \8694 , \8325 );
nor \U$8319 ( \8696 , \8693 , \8695 );
xnor \U$8320 ( \8697 , \8688 , \8696 );
xnor \U$8321 ( \8698 , \8684 , \8697 );
not \U$8322 ( \8699 , \8698 );
and \U$8323 ( \8700 , \8627 , \8699 );
not \U$8324 ( \8701 , \8627 );
and \U$8325 ( \8702 , \8701 , \8698 );
nor \U$8326 ( \8703 , \8700 , \8702 );
not \U$8327 ( \8704 , \8703 );
and \U$8328 ( \8705 , \8622 , \8704 );
not \U$8329 ( \8706 , \8622 );
and \U$8330 ( \8707 , \8706 , \8703 );
nor \U$8331 ( \8708 , \8705 , \8707 );
not \U$8332 ( \8709 , \8708 );
or \U$8333 ( \8710 , \8617 , \8709 );
or \U$8334 ( \8711 , \8616 , \8708 );
nand \U$8335 ( \8712 , \8710 , \8711 );
not \U$8336 ( \8713 , \8712 );
or \U$8337 ( \8714 , \8572 , \8713 );
not \U$8338 ( \8715 , \8708 );
nand \U$8339 ( \8716 , \8715 , \8616 );
nand \U$8340 ( \8717 , \8714 , \8716 );
not \U$8341 ( \8718 , \8680 );
not \U$8342 ( \8719 , \8660 );
not \U$8343 ( \8720 , \8719 );
and \U$8344 ( \8721 , \8718 , \8720 );
not \U$8345 ( \8722 , \8697 );
and \U$8346 ( \8723 , \8684 , \8722 );
nor \U$8347 ( \8724 , \8721 , \8723 );
not \U$8348 ( \8725 , \929 );
xor \U$8349 ( \8726 , \1188 , RIae78bc0_126);
not \U$8350 ( \8727 , \8726 );
or \U$8351 ( \8728 , \8725 , \8727 );
nand \U$8352 ( \8729 , \8640 , \953 );
nand \U$8353 ( \8730 , \8728 , \8729 );
not \U$8354 ( \8731 , \8730 );
not \U$8355 ( \8732 , \1322 );
and \U$8356 ( \8733 , RIae78e90_132, \1120 );
not \U$8357 ( \8734 , RIae78e90_132);
and \U$8358 ( \8735 , \8734 , \1119 );
nor \U$8359 ( \8736 , \8733 , \8735 );
not \U$8360 ( \8737 , \8736 );
or \U$8361 ( \8738 , \8732 , \8737 );
nand \U$8362 ( \8739 , \8689 , \1087 );
nand \U$8363 ( \8740 , \8738 , \8739 );
not \U$8364 ( \8741 , \8740 );
not \U$8365 ( \8742 , \1910 );
not \U$8366 ( \8743 , \8676 );
or \U$8367 ( \8744 , \8742 , \8743 );
nand \U$8368 ( \8745 , \1864 , RIae793b8_143);
nand \U$8369 ( \8746 , \8744 , \8745 );
not \U$8370 ( \8747 , \8746 );
and \U$8371 ( \8748 , \8741 , \8747 );
and \U$8372 ( \8749 , \8746 , \8740 );
nor \U$8373 ( \8750 , \8748 , \8749 );
not \U$8374 ( \8751 , \8750 );
or \U$8375 ( \8752 , \8731 , \8751 );
or \U$8376 ( \8753 , \8750 , \8730 );
nand \U$8377 ( \8754 , \8752 , \8753 );
not \U$8378 ( \8755 , \1440 );
not \U$8379 ( \8756 , RIae79070_136);
and \U$8380 ( \8757 , \8755 , \8756 );
and \U$8381 ( \8758 , \1440 , RIae79070_136);
nor \U$8382 ( \8759 , \8757 , \8758 );
or \U$8383 ( \8760 , \8759 , \1203 );
or \U$8384 ( \8761 , \8650 , \1249 );
nand \U$8385 ( \8762 , \8760 , \8761 );
and \U$8386 ( \8763 , RIae78b48_125, \6855 );
xnor \U$8387 ( \8764 , \8762 , \8763 );
not \U$8388 ( \8765 , \860 );
not \U$8389 ( \8766 , \2374 );
or \U$8390 ( \8767 , \8765 , \8766 );
nand \U$8391 ( \8768 , \2031 , RIae78b48_125);
nand \U$8392 ( \8769 , \8767 , \8768 );
or \U$8393 ( \8770 , \8769 , \1959 );
or \U$8394 ( \8771 , \8630 , \1128 );
nand \U$8395 ( \8772 , \8770 , \8771 );
and \U$8396 ( \8773 , \8764 , \8772 );
not \U$8397 ( \8774 , \8764 );
not \U$8398 ( \8775 , \8772 );
and \U$8399 ( \8776 , \8774 , \8775 );
nor \U$8400 ( \8777 , \8773 , \8776 );
xor \U$8401 ( \8778 , \8754 , \8777 );
and \U$8402 ( \8779 , \997 , \1143 );
not \U$8403 ( \8780 , \997 );
and \U$8404 ( \8781 , \8780 , \1366 );
nor \U$8405 ( \8782 , \8779 , \8781 );
and \U$8406 ( \8783 , \8782 , \1209 );
and \U$8407 ( \8784 , \8662 , \1010 );
nor \U$8408 ( \8785 , \8783 , \8784 );
not \U$8409 ( \8786 , \8602 );
not \U$8410 ( \8787 , \1498 );
and \U$8411 ( \8788 , \8786 , \8787 );
not \U$8412 ( \8789 , RIae79250_140);
and \U$8413 ( \8790 , \8789 , \829 );
not \U$8414 ( \8791 , \8789 );
and \U$8415 ( \8792 , \8791 , \1424 );
nor \U$8416 ( \8793 , \8790 , \8792 );
and \U$8417 ( \8794 , \8793 , \1501 );
nor \U$8418 ( \8795 , \8788 , \8794 );
xor \U$8419 ( \8796 , \8785 , \8795 );
xor \U$8420 ( \8797 , \858 , RIae78f80_134);
and \U$8421 ( \8798 , \8797 , \840 );
and \U$8422 ( \8799 , \8609 , \797 );
nor \U$8423 ( \8800 , \8798 , \8799 );
xor \U$8424 ( \8801 , \8796 , \8800 );
xnor \U$8425 ( \8802 , \8778 , \8801 );
xor \U$8426 ( \8803 , \8724 , \8802 );
or \U$8427 ( \8804 , \8584 , \8615 );
not \U$8428 ( \8805 , \8583 );
nand \U$8429 ( \8806 , \8805 , \8578 );
nand \U$8430 ( \8807 , \8804 , \8806 );
xor \U$8431 ( \8808 , \8803 , \8807 );
and \U$8432 ( \8809 , \8688 , \8696 );
nor \U$8433 ( \8810 , \8692 , \8324 );
nor \U$8434 ( \8811 , \8809 , \8810 );
not \U$8435 ( \8812 , \8811 );
not \U$8436 ( \8813 , \8614 );
not \U$8437 ( \8814 , \8600 );
or \U$8438 ( \8815 , \8813 , \8814 );
not \U$8439 ( \8816 , \8589 );
nand \U$8440 ( \8817 , \8816 , \8596 );
nand \U$8441 ( \8818 , \8815 , \8817 );
not \U$8442 ( \8819 , \8818 );
or \U$8443 ( \8820 , \8812 , \8819 );
or \U$8444 ( \8821 , \8818 , \8811 );
nand \U$8445 ( \8822 , \8820 , \8821 );
xor \U$8446 ( \8823 , \8666 , \8668 );
not \U$8447 ( \8824 , \8678 );
and \U$8448 ( \8825 , \8823 , \8824 );
and \U$8449 ( \8826 , \8666 , \8668 );
or \U$8450 ( \8827 , \8825 , \8826 );
not \U$8451 ( \8828 , \8827 );
xor \U$8452 ( \8829 , \8601 , \8607 );
and \U$8453 ( \8830 , \8829 , \8612 );
and \U$8454 ( \8831 , \8601 , \8607 );
nor \U$8455 ( \8832 , \8830 , \8831 );
xor \U$8456 ( \8833 , \8828 , \8832 );
not \U$8457 ( \8834 , \8656 );
or \U$8458 ( \8835 , \8834 , \8635 );
not \U$8459 ( \8836 , \8652 );
or \U$8460 ( \8837 , \8836 , \8643 );
nand \U$8461 ( \8838 , \8835 , \8837 );
xor \U$8462 ( \8839 , \8833 , \8838 );
xor \U$8463 ( \8840 , \8822 , \8839 );
not \U$8464 ( \8841 , \8622 );
not \U$8465 ( \8842 , \8703 );
or \U$8466 ( \8843 , \8841 , \8842 );
not \U$8467 ( \8844 , \8627 );
nand \U$8468 ( \8845 , \8844 , \8698 );
nand \U$8469 ( \8846 , \8843 , \8845 );
xor \U$8470 ( \8847 , \8840 , \8846 );
not \U$8471 ( \8848 , \8847 );
and \U$8472 ( \8849 , \8808 , \8848 );
not \U$8473 ( \8850 , \8808 );
and \U$8474 ( \8851 , \8850 , \8847 );
or \U$8475 ( \8852 , \8849 , \8851 );
nor \U$8476 ( \8853 , \8717 , \8852 );
not \U$8477 ( \8854 , \8853 );
not \U$8478 ( \8855 , \8401 );
not \U$8479 ( \8856 , \8394 );
or \U$8480 ( \8857 , \8855 , \8856 );
nand \U$8481 ( \8858 , \8306 , \8389 );
nand \U$8482 ( \8859 , \8857 , \8858 );
not \U$8483 ( \8860 , \8571 );
not \U$8484 ( \8861 , \8712 );
not \U$8485 ( \8862 , \8861 );
or \U$8486 ( \8863 , \8860 , \8862 );
not \U$8487 ( \8864 , \8571 );
nand \U$8488 ( \8865 , \8864 , \8712 );
nand \U$8489 ( \8866 , \8863 , \8865 );
or \U$8490 ( \8867 , \8859 , \8866 );
nand \U$8491 ( \8868 , \8854 , \8867 );
and \U$8492 ( \8869 , \8847 , \8808 );
and \U$8493 ( \8870 , \8840 , \8846 );
nor \U$8494 ( \8871 , \8869 , \8870 );
not \U$8495 ( \8872 , \8764 );
not \U$8496 ( \8873 , \8775 );
and \U$8497 ( \8874 , \8872 , \8873 );
buf \U$8498 ( \8875 , \8762 );
and \U$8499 ( \8876 , \8875 , \8763 );
nor \U$8500 ( \8877 , \8874 , \8876 );
not \U$8501 ( \8878 , \8746 );
and \U$8502 ( \8879 , \8877 , \8878 );
not \U$8503 ( \8880 , \8877 );
and \U$8504 ( \8881 , \8880 , \8746 );
nor \U$8505 ( \8882 , \8879 , \8881 );
xor \U$8506 ( \8883 , \8785 , \8795 );
and \U$8507 ( \8884 , \8883 , \8800 );
and \U$8508 ( \8885 , \8785 , \8795 );
nor \U$8509 ( \8886 , \8884 , \8885 );
xnor \U$8510 ( \8887 , \8882 , \8886 );
nand \U$8511 ( \8888 , \2595 , RIae78b48_125);
not \U$8512 ( \8889 , \8888 );
not \U$8513 ( \8890 , \868 );
xor \U$8514 ( \8891 , RIae78b48_125, \1406 );
not \U$8515 ( \8892 , \8891 );
or \U$8516 ( \8893 , \8890 , \8892 );
not \U$8517 ( \8894 , \8769 );
nand \U$8518 ( \8895 , \8894 , \893 );
nand \U$8519 ( \8896 , \8893 , \8895 );
not \U$8520 ( \8897 , \8896 );
or \U$8521 ( \8898 , \8889 , \8897 );
or \U$8522 ( \8899 , \8896 , \8888 );
nand \U$8523 ( \8900 , \8898 , \8899 );
not \U$8524 ( \8901 , \8900 );
and \U$8525 ( \8902 , \940 , \1132 );
and \U$8526 ( \8903 , \1077 , RIae78f80_134);
nor \U$8527 ( \8904 , \8902 , \8903 );
and \U$8528 ( \8905 , \8904 , \840 );
and \U$8529 ( \8906 , \8797 , \797 );
nor \U$8530 ( \8907 , \8905 , \8906 );
not \U$8531 ( \8908 , \8907 );
and \U$8532 ( \8909 , \8901 , \8908 );
and \U$8533 ( \8910 , \8900 , \8907 );
nor \U$8534 ( \8911 , \8909 , \8910 );
xor \U$8535 ( \8912 , \8887 , \8911 );
xor \U$8536 ( \8913 , \8828 , \8832 );
and \U$8537 ( \8914 , \8913 , \8838 );
and \U$8538 ( \8915 , \8828 , \8832 );
nor \U$8539 ( \8916 , \8914 , \8915 );
xor \U$8540 ( \8917 , \8912 , \8916 );
not \U$8541 ( \8918 , \8917 );
not \U$8542 ( \8919 , \8839 );
not \U$8543 ( \8920 , \8822 );
or \U$8544 ( \8921 , \8919 , \8920 );
not \U$8545 ( \8922 , \8811 );
nand \U$8546 ( \8923 , \8922 , \8818 );
nand \U$8547 ( \8924 , \8921 , \8923 );
not \U$8548 ( \8925 , \8778 );
not \U$8549 ( \8926 , \8801 );
and \U$8550 ( \8927 , \8925 , \8926 );
buf \U$8551 ( \8928 , \8754 );
not \U$8552 ( \8929 , \8777 );
and \U$8553 ( \8930 , \8928 , \8929 );
nor \U$8554 ( \8931 , \8927 , \8930 );
nand \U$8555 ( \8932 , RIae79610_148, RIae799d0_156);
and \U$8556 ( \8933 , \8932 , RIae793b8_143);
not \U$8557 ( \8934 , \8933 );
not \U$8558 ( \8935 , \1062 );
not \U$8559 ( \8936 , \8759 );
not \U$8560 ( \8937 , \8936 );
or \U$8561 ( \8938 , \8935 , \8937 );
xor \U$8562 ( \8939 , RIae79070_136, \1162 );
not \U$8563 ( \8940 , \8939 );
nand \U$8564 ( \8941 , \8940 , \1049 );
nand \U$8565 ( \8942 , \8938 , \8941 );
not \U$8566 ( \8943 , \8942 );
or \U$8567 ( \8944 , \8934 , \8943 );
or \U$8568 ( \8945 , \8942 , \8933 );
nand \U$8569 ( \8946 , \8944 , \8945 );
not \U$8570 ( \8947 , \8946 );
and \U$8571 ( \8948 , \8793 , \1499 );
and \U$8572 ( \8949 , \1488 , \1501 );
nor \U$8573 ( \8950 , \8948 , \8949 );
not \U$8574 ( \8951 , \8950 );
and \U$8575 ( \8952 , \8947 , \8951 );
and \U$8576 ( \8953 , \8950 , \8946 );
nor \U$8577 ( \8954 , \8952 , \8953 );
not \U$8578 ( \8955 , \8954 );
not \U$8579 ( \8956 , \8730 );
not \U$8580 ( \8957 , \8750 );
not \U$8581 ( \8958 , \8957 );
or \U$8582 ( \8959 , \8956 , \8958 );
nand \U$8583 ( \8960 , \8740 , \8878 );
nand \U$8584 ( \8961 , \8959 , \8960 );
not \U$8585 ( \8962 , \8961 );
or \U$8586 ( \8963 , \8955 , \8962 );
or \U$8587 ( \8964 , \8961 , \8954 );
nand \U$8588 ( \8965 , \8963 , \8964 );
and \U$8589 ( \8966 , RIae78bc0_126, \7702 );
not \U$8590 ( \8967 , RIae78bc0_126);
and \U$8591 ( \8968 , \8967 , \8047 );
nor \U$8592 ( \8969 , \8966 , \8968 );
nand \U$8593 ( \8970 , \8969 , \929 );
nand \U$8594 ( \8971 , \8726 , \953 );
and \U$8595 ( \8972 , \8970 , \8971 );
and \U$8596 ( \8973 , \8736 , \1259 );
and \U$8597 ( \8974 , RIae78e90_132, \880 );
not \U$8598 ( \8975 , RIae78e90_132);
and \U$8599 ( \8976 , \8975 , \879 );
nor \U$8600 ( \8977 , \8974 , \8976 );
and \U$8601 ( \8978 , \8977 , \1322 );
nor \U$8602 ( \8979 , \8973 , \8978 );
xnor \U$8603 ( \8980 , \8972 , \8979 );
and \U$8604 ( \8981 , \6414 , \782 );
not \U$8605 ( \8982 , \6414 );
and \U$8606 ( \8983 , \8982 , \783 );
or \U$8607 ( \8984 , \8981 , \8983 );
and \U$8608 ( \8985 , \8984 , \1209 );
and \U$8609 ( \8986 , \8782 , \1430 );
nor \U$8610 ( \8987 , \8985 , \8986 );
xor \U$8611 ( \8988 , \8980 , \8987 );
and \U$8612 ( \8989 , \8965 , \8988 );
not \U$8613 ( \8990 , \8965 );
not \U$8614 ( \8991 , \8988 );
and \U$8615 ( \8992 , \8990 , \8991 );
nor \U$8616 ( \8993 , \8989 , \8992 );
and \U$8617 ( \8994 , \8931 , \8993 );
not \U$8618 ( \8995 , \8931 );
not \U$8619 ( \8996 , \8993 );
and \U$8620 ( \8997 , \8995 , \8996 );
nor \U$8621 ( \8998 , \8994 , \8997 );
xnor \U$8622 ( \8999 , \8924 , \8998 );
not \U$8623 ( \9000 , \8999 );
or \U$8624 ( \9001 , \8918 , \9000 );
or \U$8625 ( \9002 , \8999 , \8917 );
nand \U$8626 ( \9003 , \9001 , \9002 );
not \U$8627 ( \9004 , \9003 );
not \U$8628 ( \9005 , \8724 );
not \U$8629 ( \9006 , \8802 );
and \U$8630 ( \9007 , \9005 , \9006 );
and \U$8631 ( \9008 , \8803 , \8807 );
nor \U$8632 ( \9009 , \9007 , \9008 );
not \U$8633 ( \9010 , \9009 );
and \U$8634 ( \9011 , \9004 , \9010 );
and \U$8635 ( \9012 , \9003 , \9009 );
nor \U$8636 ( \9013 , \9011 , \9012 );
nand \U$8637 ( \9014 , \8871 , \9013 );
not \U$8638 ( \9015 , \9009 );
not \U$8639 ( \9016 , \9015 );
not \U$8640 ( \9017 , \9003 );
or \U$8641 ( \9018 , \9016 , \9017 );
not \U$8642 ( \9019 , \8917 );
nand \U$8643 ( \9020 , \9019 , \8999 );
nand \U$8644 ( \9021 , \9018 , \9020 );
not \U$8645 ( \9022 , \9021 );
xor \U$8646 ( \9023 , \8887 , \8911 );
and \U$8647 ( \9024 , \9023 , \8916 );
and \U$8648 ( \9025 , \8887 , \8911 );
or \U$8649 ( \9026 , \9024 , \9025 );
not \U$8650 ( \9027 , \9026 );
not \U$8651 ( \9028 , \8886 );
not \U$8652 ( \9029 , \8882 );
or \U$8653 ( \9030 , \9028 , \9029 );
or \U$8654 ( \9031 , \8877 , \8878 );
nand \U$8655 ( \9032 , \9030 , \9031 );
and \U$8656 ( \9033 , \1429 , \1013 );
and \U$8657 ( \9034 , \8984 , \1010 );
nor \U$8658 ( \9035 , \9033 , \9034 );
xor \U$8659 ( \9036 , \8768 , \9035 );
and \U$8660 ( \9037 , \1445 , \840 );
and \U$8661 ( \9038 , \8904 , \797 );
nor \U$8662 ( \9039 , \9037 , \9038 );
xor \U$8663 ( \9040 , \9036 , \9039 );
not \U$8664 ( \9041 , \8933 );
not \U$8665 ( \9042 , \9041 );
not \U$8666 ( \9043 , \8942 );
or \U$8667 ( \9044 , \9042 , \9043 );
not \U$8668 ( \9045 , \8950 );
nand \U$8669 ( \9046 , \9045 , \8946 );
nand \U$8670 ( \9047 , \9044 , \9046 );
not \U$8671 ( \9048 , \1129 );
not \U$8672 ( \9049 , \8891 );
or \U$8673 ( \9050 , \9048 , \9049 );
nand \U$8674 ( \9051 , \1512 , \868 );
nand \U$8675 ( \9052 , \9050 , \9051 );
not \U$8676 ( \9053 , \9052 );
not \U$8677 ( \9054 , \1506 );
and \U$8678 ( \9055 , \9053 , \9054 );
and \U$8679 ( \9056 , \9052 , \1506 );
nor \U$8680 ( \9057 , \9055 , \9056 );
xor \U$8681 ( \9058 , \9047 , \9057 );
xor \U$8682 ( \9059 , \9040 , \9058 );
xor \U$8683 ( \9060 , \9032 , \9059 );
not \U$8684 ( \9061 , \9060 );
not \U$8685 ( \9062 , \1412 );
not \U$8686 ( \9063 , \1646 );
and \U$8687 ( \9064 , \9062 , \9063 );
and \U$8688 ( \9065 , \8977 , \1259 );
nor \U$8689 ( \9066 , \9064 , \9065 );
not \U$8690 ( \9067 , \1394 );
or \U$8691 ( \9068 , \9067 , \1203 );
or \U$8692 ( \9069 , \8939 , \1249 );
nand \U$8693 ( \9070 , \9068 , \9069 );
and \U$8694 ( \9071 , \9066 , \9070 );
not \U$8695 ( \9072 , \9066 );
not \U$8696 ( \9073 , \9070 );
and \U$8697 ( \9074 , \9072 , \9073 );
nor \U$8698 ( \9075 , \9071 , \9074 );
and \U$8699 ( \9076 , \1477 , \929 );
and \U$8700 ( \9077 , \8969 , \953 );
nor \U$8701 ( \9078 , \9076 , \9077 );
xnor \U$8702 ( \9079 , \9075 , \9078 );
not \U$8703 ( \9080 , \9079 );
not \U$8704 ( \9081 , \8888 );
not \U$8705 ( \9082 , \9081 );
not \U$8706 ( \9083 , \8896 );
or \U$8707 ( \9084 , \9082 , \9083 );
not \U$8708 ( \9085 , \8907 );
nand \U$8709 ( \9086 , \9085 , \8900 );
nand \U$8710 ( \9087 , \9084 , \9086 );
or \U$8711 ( \9088 , \8980 , \8987 );
or \U$8712 ( \9089 , \8972 , \8979 );
nand \U$8713 ( \9090 , \9088 , \9089 );
xor \U$8714 ( \9091 , \9087 , \9090 );
not \U$8715 ( \9092 , \9091 );
or \U$8716 ( \9093 , \9080 , \9092 );
or \U$8717 ( \9094 , \9091 , \9079 );
nand \U$8718 ( \9095 , \9093 , \9094 );
not \U$8719 ( \9096 , \9095 );
and \U$8720 ( \9097 , \8965 , \8988 );
not \U$8721 ( \9098 , \8954 );
and \U$8722 ( \9099 , \8961 , \9098 );
nor \U$8723 ( \9100 , \9097 , \9099 );
not \U$8724 ( \9101 , \9100 );
or \U$8725 ( \9102 , \9096 , \9101 );
or \U$8726 ( \9103 , \9100 , \9095 );
nand \U$8727 ( \9104 , \9102 , \9103 );
not \U$8728 ( \9105 , \9104 );
not \U$8729 ( \9106 , \9105 );
or \U$8730 ( \9107 , \9061 , \9106 );
not \U$8731 ( \9108 , \9060 );
nand \U$8732 ( \9109 , \9108 , \9104 );
nand \U$8733 ( \9110 , \9107 , \9109 );
not \U$8734 ( \9111 , \9110 );
or \U$8735 ( \9112 , \9027 , \9111 );
or \U$8736 ( \9113 , \9110 , \9026 );
nand \U$8737 ( \9114 , \9112 , \9113 );
not \U$8738 ( \9115 , \8998 );
not \U$8739 ( \9116 , \9115 );
not \U$8740 ( \9117 , \8924 );
or \U$8741 ( \9118 , \9116 , \9117 );
or \U$8742 ( \9119 , \8996 , \8931 );
nand \U$8743 ( \9120 , \9118 , \9119 );
xnor \U$8744 ( \9121 , \9114 , \9120 );
nand \U$8745 ( \9122 , \9022 , \9121 );
nand \U$8746 ( \9123 , \9014 , \9122 );
nor \U$8747 ( \9124 , \8868 , \9123 );
not \U$8748 ( \9125 , \9120 );
not \U$8749 ( \9126 , \9114 );
or \U$8750 ( \9127 , \9125 , \9126 );
not \U$8751 ( \9128 , \9026 );
nand \U$8752 ( \9129 , \9128 , \9110 );
nand \U$8753 ( \9130 , \9127 , \9129 );
not \U$8754 ( \9131 , \9130 );
not \U$8755 ( \9132 , \9057 );
and \U$8756 ( \9133 , \9047 , \9132 );
and \U$8757 ( \9134 , \9052 , \1505 );
nor \U$8758 ( \9135 , \9133 , \9134 );
not \U$8759 ( \9136 , \9135 );
xnor \U$8760 ( \9137 , \1408 , \1415 );
xnor \U$8761 ( \9138 , \1510 , \1514 );
xor \U$8762 ( \9139 , \9137 , \9138 );
not \U$8763 ( \9140 , \9139 );
or \U$8764 ( \9141 , \9136 , \9140 );
or \U$8765 ( \9142 , \9139 , \9135 );
nand \U$8766 ( \9143 , \9141 , \9142 );
not \U$8767 ( \9144 , \9091 );
not \U$8768 ( \9145 , \9144 );
not \U$8769 ( \9146 , \9079 );
and \U$8770 ( \9147 , \9145 , \9146 );
and \U$8771 ( \9148 , \9090 , \9087 );
nor \U$8772 ( \9149 , \9147 , \9148 );
or \U$8773 ( \9150 , \9075 , \9078 );
or \U$8774 ( \9151 , \9066 , \9073 );
nand \U$8775 ( \9152 , \9150 , \9151 );
xor \U$8776 ( \9153 , \8768 , \9035 );
and \U$8777 ( \9154 , \9153 , \9039 );
and \U$8778 ( \9155 , \8768 , \9035 );
nor \U$8779 ( \9156 , \9154 , \9155 );
xor \U$8780 ( \9157 , \9152 , \9156 );
not \U$8781 ( \9158 , \1447 );
not \U$8782 ( \9159 , \1453 );
or \U$8783 ( \9160 , \9158 , \9159 );
or \U$8784 ( \9161 , \1453 , \1447 );
nand \U$8785 ( \9162 , \9160 , \9161 );
and \U$8786 ( \9163 , \9157 , \9162 );
not \U$8787 ( \9164 , \9157 );
not \U$8788 ( \9165 , \9162 );
and \U$8789 ( \9166 , \9164 , \9165 );
nor \U$8790 ( \9167 , \9163 , \9166 );
not \U$8791 ( \9168 , \9167 );
and \U$8792 ( \9169 , \9149 , \9168 );
not \U$8793 ( \9170 , \9149 );
and \U$8794 ( \9171 , \9170 , \9167 );
nor \U$8795 ( \9172 , \9169 , \9171 );
not \U$8796 ( \9173 , \9172 );
not \U$8797 ( \9174 , \9058 );
not \U$8798 ( \9175 , \9040 );
and \U$8799 ( \9176 , \9174 , \9175 );
and \U$8800 ( \9177 , \9059 , \9032 );
nor \U$8801 ( \9178 , \9176 , \9177 );
not \U$8802 ( \9179 , \9178 );
and \U$8803 ( \9180 , \9173 , \9179 );
and \U$8804 ( \9181 , \9172 , \9178 );
nor \U$8805 ( \9182 , \9180 , \9181 );
xnor \U$8806 ( \9183 , \9143 , \9182 );
not \U$8807 ( \9184 , \9183 );
not \U$8808 ( \9185 , \9100 );
not \U$8809 ( \9186 , \9095 );
not \U$8810 ( \9187 , \9186 );
and \U$8811 ( \9188 , \9185 , \9187 );
not \U$8812 ( \9189 , \9105 );
and \U$8813 ( \9190 , \9189 , \9060 );
nor \U$8814 ( \9191 , \9188 , \9190 );
not \U$8815 ( \9192 , \9191 );
and \U$8816 ( \9193 , \9184 , \9192 );
and \U$8817 ( \9194 , \9183 , \9191 );
nor \U$8818 ( \9195 , \9193 , \9194 );
nand \U$8819 ( \9196 , \9131 , \9195 );
not \U$8820 ( \9197 , \9172 );
or \U$8821 ( \9198 , \9197 , \9178 );
or \U$8822 ( \9199 , \9149 , \9168 );
nand \U$8823 ( \9200 , \9198 , \9199 );
xnor \U$8824 ( \9201 , \1519 , \1522 );
xnor \U$8825 ( \9202 , \1418 , \1459 );
not \U$8826 ( \9203 , \9202 );
nand \U$8827 ( \9204 , \9157 , \9162 );
nand \U$8828 ( \9205 , \9152 , \9156 );
and \U$8829 ( \9206 , \9204 , \9205 );
not \U$8830 ( \9207 , \9206 );
or \U$8831 ( \9208 , \9203 , \9207 );
or \U$8832 ( \9209 , \9206 , \9202 );
nand \U$8833 ( \9210 , \9208 , \9209 );
nor \U$8834 ( \9211 , \9201 , \9210 );
not \U$8835 ( \9212 , \9211 );
nand \U$8836 ( \9213 , \9210 , \9201 );
nand \U$8837 ( \9214 , \9212 , \9213 );
not \U$8838 ( \9215 , \9214 );
and \U$8839 ( \9216 , \9137 , \9138 );
or \U$8840 ( \9217 , \9135 , \9216 );
or \U$8841 ( \9218 , \9138 , \9137 );
nand \U$8842 ( \9219 , \9217 , \9218 );
not \U$8843 ( \9220 , \9219 );
not \U$8844 ( \9221 , \9220 );
and \U$8845 ( \9222 , \9215 , \9221 );
and \U$8846 ( \9223 , \9214 , \9220 );
nor \U$8847 ( \9224 , \9222 , \9223 );
xnor \U$8848 ( \9225 , \9200 , \9224 );
not \U$8849 ( \9226 , \9191 );
not \U$8850 ( \9227 , \9226 );
not \U$8851 ( \9228 , \9183 );
or \U$8852 ( \9229 , \9227 , \9228 );
not \U$8853 ( \9230 , \9182 );
nand \U$8854 ( \9231 , \9230 , \9143 );
nand \U$8855 ( \9232 , \9229 , \9231 );
nor \U$8856 ( \9233 , \9225 , \9232 );
not \U$8857 ( \9234 , \9233 );
not \U$8858 ( \9235 , \9200 );
not \U$8859 ( \9236 , \9224 );
not \U$8860 ( \9237 , \9236 );
or \U$8861 ( \9238 , \9235 , \9237 );
not \U$8862 ( \9239 , \9214 );
or \U$8863 ( \9240 , \9239 , \9220 );
nand \U$8864 ( \9241 , \9238 , \9240 );
and \U$8865 ( \9242 , \1471 , \1525 );
not \U$8866 ( \9243 , \1471 );
not \U$8867 ( \9244 , \1525 );
and \U$8868 ( \9245 , \9243 , \9244 );
nor \U$8869 ( \9246 , \9242 , \9245 );
xor \U$8870 ( \9247 , \1193 , \1221 );
xor \U$8871 ( \9248 , \9247 , \1239 );
xor \U$8872 ( \9249 , \9246 , \9248 );
not \U$8873 ( \9250 , \9201 );
not \U$8874 ( \9251 , \9250 );
not \U$8875 ( \9252 , \9210 );
or \U$8876 ( \9253 , \9251 , \9252 );
not \U$8877 ( \9254 , \9202 );
or \U$8878 ( \9255 , \9206 , \9254 );
nand \U$8879 ( \9256 , \9253 , \9255 );
xor \U$8880 ( \9257 , \9249 , \9256 );
or \U$8881 ( \9258 , \9241 , \9257 );
and \U$8882 ( \9259 , \9196 , \9234 , \9258 );
not \U$8883 ( \9260 , \1534 );
xor \U$8884 ( \9261 , \1527 , \1528 );
not \U$8885 ( \9262 , \9261 );
or \U$8886 ( \9263 , \9260 , \9262 );
or \U$8887 ( \9264 , \9261 , \1534 );
nand \U$8888 ( \9265 , \9263 , \9264 );
xor \U$8889 ( \9266 , \9246 , \9248 );
and \U$8890 ( \9267 , \9266 , \9256 );
and \U$8891 ( \9268 , \9246 , \9248 );
or \U$8892 ( \9269 , \9267 , \9268 );
or \U$8893 ( \9270 , \9265 , \9269 );
and \U$8894 ( \9271 , \9124 , \9259 , \9270 );
nand \U$8895 ( \9272 , \6825 , \8565 , \9271 );
not \U$8896 ( \9273 , \9272 );
not \U$8897 ( \9274 , \9273 );
not \U$8898 ( \9275 , \2249 );
not \U$8899 ( \9276 , \5722 );
not \U$8900 ( \9277 , RIae79ac0_158);
and \U$8901 ( \9278 , \9276 , \9277 );
buf \U$8902 ( \9279 , \5721 );
buf \U$8903 ( \9280 , \9279 );
and \U$8904 ( \9281 , \9280 , RIae79ac0_158);
nor \U$8905 ( \9282 , \9278 , \9281 );
not \U$8906 ( \9283 , \9282 );
or \U$8907 ( \9284 , \9275 , \9283 );
not \U$8908 ( \9285 , RIae79ac0_158);
not \U$8909 ( \9286 , \6345 );
not \U$8910 ( \9287 , \9286 );
or \U$8911 ( \9288 , \9285 , \9287 );
buf \U$8912 ( \9289 , \6344 );
buf \U$8913 ( \9290 , \9289 );
not \U$8914 ( \9291 , \9290 );
or \U$8915 ( \9292 , \9291 , RIae79ac0_158);
nand \U$8916 ( \9293 , \9288 , \9292 );
nand \U$8917 ( \9294 , \9293 , \2272 );
nand \U$8918 ( \9295 , \9284 , \9294 );
not \U$8919 ( \9296 , \1820 );
not \U$8920 ( \9297 , RIae79688_149);
buf \U$8921 ( \9298 , \6229 );
not \U$8922 ( \9299 , \9298 );
not \U$8923 ( \9300 , \9299 );
or \U$8924 ( \9301 , \9297 , \9300 );
nand \U$8925 ( \9302 , \6230 , \2970 );
nand \U$8926 ( \9303 , \9301 , \9302 );
not \U$8927 ( \9304 , \9303 );
or \U$8928 ( \9305 , \9296 , \9304 );
buf \U$8929 ( \9306 , \3183 );
not \U$8930 ( \9307 , \9306 );
nand \U$8931 ( \9308 , \6217 , \589 );
not \U$8932 ( \9309 , \9308 );
and \U$8933 ( \9310 , \9307 , \9309 );
and \U$8934 ( \9311 , \9306 , \9308 );
nor \U$8935 ( \9312 , \9310 , \9311 );
buf \U$8936 ( \9313 , \9312 );
and \U$8937 ( \9314 , RIae79688_149, \9313 );
not \U$8938 ( \9315 , RIae79688_149);
buf \U$8939 ( \9316 , \9312 );
not \U$8940 ( \9317 , \9316 );
and \U$8941 ( \9318 , \9315 , \9317 );
or \U$8942 ( \9319 , \9314 , \9318 );
buf \U$8943 ( \9320 , \1843 );
nand \U$8944 ( \9321 , \9319 , \9320 );
nand \U$8945 ( \9322 , \9305 , \9321 );
xor \U$8946 ( \9323 , \9295 , \9322 );
not \U$8947 ( \9324 , \2011 );
not \U$8948 ( \9325 , \512 );
not \U$8949 ( \9326 , \9325 );
buf \U$8950 ( \9327 , \510 );
not \U$8951 ( \9328 , \9327 );
not \U$8952 ( \9329 , \562 );
not \U$8953 ( \9330 , \3170 );
or \U$8954 ( \9331 , \9329 , \9330 );
nand \U$8955 ( \9332 , \9331 , \3178 );
not \U$8956 ( \9333 , \9332 );
or \U$8957 ( \9334 , \9328 , \9333 );
not \U$8958 ( \9335 , \575 );
nand \U$8959 ( \9336 , \9334 , \9335 );
not \U$8960 ( \9337 , \9336 );
or \U$8961 ( \9338 , \9326 , \9337 );
nand \U$8962 ( \9339 , \9338 , \578 );
not \U$8963 ( \9340 , \9339 );
not \U$8964 ( \9341 , \511 );
nand \U$8965 ( \9342 , \9341 , \580 );
not \U$8966 ( \9343 , \9342 );
and \U$8967 ( \9344 , \9340 , \9343 );
and \U$8968 ( \9345 , \9339 , \9342 );
nor \U$8969 ( \9346 , \9344 , \9345 );
buf \U$8970 ( \9347 , \9346 );
and \U$8971 ( \9348 , RIae79610_148, \9347 );
not \U$8972 ( \9349 , RIae79610_148);
not \U$8973 ( \9350 , \9347 );
and \U$8974 ( \9351 , \9349 , \9350 );
or \U$8975 ( \9352 , \9348 , \9351 );
not \U$8976 ( \9353 , \9352 );
or \U$8977 ( \9354 , \9324 , \9353 );
not \U$8978 ( \9355 , \9327 );
not \U$8979 ( \9356 , \9332 );
or \U$8980 ( \9357 , \9355 , \9356 );
nand \U$8981 ( \9358 , \9357 , \9335 );
nand \U$8982 ( \9359 , \9325 , \578 );
or \U$8983 ( \9360 , \9358 , \9359 );
nand \U$8984 ( \9361 , \9358 , \9359 );
nand \U$8985 ( \9362 , \9360 , \9361 );
buf \U$8986 ( \9363 , \9362 );
not \U$8987 ( \9364 , \9363 );
and \U$8988 ( \9365 , RIae79610_148, \9364 );
not \U$8989 ( \9366 , RIae79610_148);
buf \U$8990 ( \9367 , \9362 );
and \U$8991 ( \9368 , \9366 , \9367 );
or \U$8992 ( \9369 , \9365 , \9368 );
buf \U$8993 ( \9370 , \2063 );
nand \U$8994 ( \9371 , \9369 , \9370 );
nand \U$8995 ( \9372 , \9354 , \9371 );
xor \U$8996 ( \9373 , \9323 , \9372 );
not \U$8997 ( \9374 , \9373 );
not \U$8998 ( \9375 , \1501 );
not \U$8999 ( \9376 , \489 );
not \U$9000 ( \9377 , \9376 );
not \U$9001 ( \9378 , \496 );
buf \U$9002 ( \9379 , \3170 );
not \U$9003 ( \9380 , \9379 );
or \U$9004 ( \9381 , \9378 , \9380 );
not \U$9005 ( \9382 , \458 );
nand \U$9006 ( \9383 , \9381 , \9382 );
not \U$9007 ( \9384 , \9383 );
or \U$9008 ( \9385 , \9377 , \9384 );
buf \U$9009 ( \9386 , \459 );
nand \U$9010 ( \9387 , \9385 , \9386 );
not \U$9011 ( \9388 , \9387 );
or \U$9012 ( \9389 , \3174 , \490 );
not \U$9013 ( \9390 , \9389 );
and \U$9014 ( \9391 , \9388 , \9390 );
and \U$9015 ( \9392 , \9387 , \9389 );
nor \U$9016 ( \9393 , \9391 , \9392 );
not \U$9017 ( \9394 , \9393 );
buf \U$9018 ( \9395 , \9394 );
and \U$9019 ( \9396 , RIae79250_140, \9395 );
not \U$9020 ( \9397 , RIae79250_140);
not \U$9021 ( \9398 , \9395 );
and \U$9022 ( \9399 , \9397 , \9398 );
nor \U$9023 ( \9400 , \9396 , \9399 );
not \U$9024 ( \9401 , \9400 );
or \U$9025 ( \9402 , \9375 , \9401 );
not \U$9026 ( \9403 , \1498 );
not \U$9027 ( \9404 , RIae79250_140);
buf \U$9028 ( \9405 , \9383 );
not \U$9029 ( \9406 , \9405 );
nand \U$9030 ( \9407 , \9376 , \9386 );
not \U$9031 ( \9408 , \9407 );
and \U$9032 ( \9409 , \9406 , \9408 );
and \U$9033 ( \9410 , \9405 , \9407 );
nor \U$9034 ( \9411 , \9409 , \9410 );
buf \U$9035 ( \9412 , \9411 );
not \U$9036 ( \9413 , \9412 );
or \U$9037 ( \9414 , \9404 , \9413 );
not \U$9038 ( \9415 , \9411 );
buf \U$9039 ( \9416 , \9415 );
not \U$9040 ( \9417 , \9416 );
or \U$9041 ( \9418 , \9417 , RIae79250_140);
nand \U$9042 ( \9419 , \9414 , \9418 );
nand \U$9043 ( \9420 , \9403 , \9419 );
nand \U$9044 ( \9421 , \9402 , \9420 );
not \U$9045 ( \9422 , \9421 );
not \U$9046 ( \9423 , \1864 );
not \U$9047 ( \9424 , \1902 );
not \U$9048 ( \9425 , \509 );
not \U$9049 ( \9426 , \9425 );
not \U$9050 ( \9427 , \9332 );
or \U$9051 ( \9428 , \9426 , \9427 );
not \U$9052 ( \9429 , \569 );
buf \U$9053 ( \9430 , \9429 );
nand \U$9054 ( \9431 , \9428 , \9430 );
nand \U$9055 ( \9432 , \571 , \574 );
not \U$9056 ( \9433 , \9432 );
and \U$9057 ( \9434 , \9431 , \9433 );
not \U$9058 ( \9435 , \9431 );
and \U$9059 ( \9436 , \9435 , \9432 );
nor \U$9060 ( \9437 , \9434 , \9436 );
buf \U$9061 ( \9438 , \9437 );
not \U$9062 ( \9439 , \9438 );
or \U$9063 ( \9440 , \9424 , \9439 );
buf \U$9064 ( \9441 , \9437 );
not \U$9065 ( \9442 , \9441 );
nand \U$9066 ( \9443 , \9442 , RIae793b8_143);
nand \U$9067 ( \9444 , \9440 , \9443 );
not \U$9068 ( \9445 , \9444 );
or \U$9069 ( \9446 , \9423 , \9445 );
not \U$9070 ( \9447 , RIae793b8_143);
buf \U$9071 ( \9448 , \9332 );
nand \U$9072 ( \9449 , \9425 , \9429 );
not \U$9073 ( \9450 , \9449 );
and \U$9074 ( \9451 , \9448 , \9450 );
not \U$9075 ( \9452 , \9448 );
and \U$9076 ( \9453 , \9452 , \9449 );
nor \U$9077 ( \9454 , \9451 , \9453 );
buf \U$9078 ( \9455 , \9454 );
not \U$9079 ( \9456 , \9455 );
not \U$9080 ( \9457 , \9456 );
or \U$9081 ( \9458 , \9447 , \9457 );
buf \U$9082 ( \9459 , \9454 );
nand \U$9083 ( \9460 , \9459 , \1902 );
nand \U$9084 ( \9461 , \9458 , \9460 );
nand \U$9085 ( \9462 , \9461 , \1910 );
nand \U$9086 ( \9463 , \9446 , \9462 );
not \U$9087 ( \9464 , \9463 );
or \U$9088 ( \9465 , \9422 , \9464 );
or \U$9089 ( \9466 , \9421 , \9463 );
nand \U$9090 ( \9467 , \9465 , \9466 );
xor \U$9091 ( \9468 , RIae7a6f0_184, RIae7a858_187);
not \U$9092 ( \9469 , \9468 );
xor \U$9093 ( \9470 , RIae7a858_187, RIae7a8d0_188);
nor \U$9094 ( \9471 , \9469 , \9470 );
buf \U$9095 ( \9472 , \9471 );
buf \U$9096 ( \9473 , \9472 );
not \U$9097 ( \9474 , \9473 );
xor \U$9098 ( \9475 , RIae7a6f0_184, \991 );
not \U$9099 ( \9476 , \9475 );
or \U$9100 ( \9477 , \9474 , \9476 );
buf \U$9101 ( \9478 , \9470 );
nand \U$9102 ( \9479 , \9478 , RIae7a6f0_184);
nand \U$9103 ( \9480 , \9477 , \9479 );
xor \U$9104 ( \9481 , \9467 , \9480 );
not \U$9105 ( \9482 , \9481 );
not \U$9106 ( \9483 , \9482 );
or \U$9107 ( \9484 , \9374 , \9483 );
not \U$9108 ( \9485 , \9373 );
not \U$9109 ( \9486 , \9485 );
not \U$9110 ( \9487 , \9481 );
or \U$9111 ( \9488 , \9486 , \9487 );
and \U$9112 ( \9489 , RIae7a2b8_175, RIae7a678_183);
not \U$9113 ( \9490 , RIae7a2b8_175);
not \U$9114 ( \9491 , RIae7a678_183);
and \U$9115 ( \9492 , \9490 , \9491 );
nor \U$9116 ( \9493 , \9489 , \9492 );
not \U$9117 ( \9494 , \9493 );
and \U$9118 ( \9495 , RIae79fe8_169, RIae7a678_183);
not \U$9119 ( \9496 , RIae79fe8_169);
and \U$9120 ( \9497 , \9496 , \9491 );
nor \U$9121 ( \9498 , \9495 , \9497 );
and \U$9122 ( \9499 , \9494 , \9498 );
not \U$9123 ( \9500 , \9499 );
not \U$9124 ( \9501 , \3069 );
and \U$9125 ( \9502 , \9501 , RIae79fe8_169);
not \U$9126 ( \9503 , \9501 );
not \U$9127 ( \9504 , RIae79fe8_169);
and \U$9128 ( \9505 , \9503 , \9504 );
nor \U$9129 ( \9506 , \9502 , \9505 );
not \U$9130 ( \9507 , \9506 );
or \U$9131 ( \9508 , \9500 , \9507 );
not \U$9132 ( \9509 , \9504 );
not \U$9133 ( \9510 , \3765 );
or \U$9134 ( \9511 , \9509 , \9510 );
not \U$9135 ( \9512 , \2993 );
not \U$9136 ( \9513 , RIae79fe8_169);
or \U$9137 ( \9514 , \9512 , \9513 );
nand \U$9138 ( \9515 , \9511 , \9514 );
not \U$9139 ( \9516 , \9494 );
buf \U$9140 ( \9517 , \9516 );
buf \U$9141 ( \9518 , \9517 );
nand \U$9142 ( \9519 , \9515 , \9518 );
nand \U$9143 ( \9520 , \9508 , \9519 );
not \U$9144 ( \9521 , \9520 );
not \U$9145 ( \9522 , RIae7a768_185);
and \U$9146 ( \9523 , RIae7a6f0_184, \9522 );
not \U$9147 ( \9524 , RIae7a6f0_184);
and \U$9148 ( \9525 , \9524 , RIae7a768_185);
nor \U$9149 ( \9526 , \9523 , \9525 );
not \U$9150 ( \9527 , \9526 );
not \U$9151 ( \9528 , \9527 );
not \U$9152 ( \9529 , RIae7a7e0_186);
and \U$9153 ( \9530 , \9529 , \1993 );
not \U$9154 ( \9531 , \9529 );
not \U$9155 ( \9532 , \780 );
and \U$9156 ( \9533 , \9531 , \9532 );
nor \U$9157 ( \9534 , \9530 , \9533 );
not \U$9158 ( \9535 , \9534 );
or \U$9159 ( \9536 , \9528 , \9535 );
not \U$9160 ( \9537 , RIae7a7e0_186);
not \U$9161 ( \9538 , \9537 );
not \U$9162 ( \9539 , \2323 );
or \U$9163 ( \9540 , \9538 , \9539 );
not \U$9164 ( \9541 , RIae7a7e0_186);
or \U$9165 ( \9542 , \1141 , \9541 );
nand \U$9166 ( \9543 , \9540 , \9542 );
and \U$9167 ( \9544 , RIae7a7e0_186, RIae7a768_185);
not \U$9168 ( \9545 , RIae7a7e0_186);
and \U$9169 ( \9546 , \9545 , \9522 );
nor \U$9170 ( \9547 , \9544 , \9546 );
nand \U$9171 ( \9548 , \9526 , \9547 );
not \U$9172 ( \9549 , \9548 );
nand \U$9173 ( \9550 , \9543 , \9549 );
nand \U$9174 ( \9551 , \9536 , \9550 );
not \U$9175 ( \9552 , \6214 );
not \U$9176 ( \9553 , RIae79ef8_167);
not \U$9177 ( \9554 , \2954 );
or \U$9178 ( \9555 , \9553 , \9554 );
or \U$9179 ( \9556 , \2153 , RIae79ef8_167);
nand \U$9180 ( \9557 , \9555 , \9556 );
not \U$9181 ( \9558 , \9557 );
or \U$9182 ( \9559 , \9552 , \9558 );
not \U$9183 ( \9560 , RIae79ef8_167);
not \U$9184 ( \9561 , \9560 );
not \U$9185 ( \9562 , \2309 );
or \U$9186 ( \9563 , \9561 , \9562 );
nand \U$9187 ( \9564 , \2305 , RIae79ef8_167);
nand \U$9188 ( \9565 , \9563 , \9564 );
nand \U$9189 ( \9566 , \9565 , \6201 );
nand \U$9190 ( \9567 , \9559 , \9566 );
or \U$9191 ( \9568 , \9551 , \9567 );
not \U$9192 ( \9569 , \9568 );
or \U$9193 ( \9570 , \9521 , \9569 );
nand \U$9194 ( \9571 , \9551 , \9567 );
nand \U$9195 ( \9572 , \9570 , \9571 );
nand \U$9196 ( \9573 , \9488 , \9572 );
nand \U$9197 ( \9574 , \9484 , \9573 );
not \U$9198 ( \9575 , \9574 );
buf \U$9199 ( \9576 , \2431 );
not \U$9200 ( \9577 , \9576 );
not \U$9201 ( \9578 , RIae79778_151);
not \U$9202 ( \9579 , \4112 );
or \U$9203 ( \9580 , \9578 , \9579 );
nand \U$9204 ( \9581 , \5911 , \2504 );
nand \U$9205 ( \9582 , \9580 , \9581 );
not \U$9206 ( \9583 , \9582 );
or \U$9207 ( \9584 , \9577 , \9583 );
and \U$9208 ( \9585 , RIae79778_151, \5890 );
not \U$9209 ( \9586 , RIae79778_151);
and \U$9210 ( \9587 , \9586 , \2093 );
or \U$9211 ( \9588 , \9585 , \9587 );
nand \U$9212 ( \9589 , \9588 , \2450 );
nand \U$9213 ( \9590 , \9584 , \9589 );
not \U$9214 ( \9591 , \9590 );
not \U$9215 ( \9592 , \9403 );
not \U$9216 ( \9593 , \495 );
not \U$9217 ( \9594 , \9593 );
buf \U$9218 ( \9595 , \9379 );
not \U$9219 ( \9596 , \9595 );
or \U$9220 ( \9597 , \9594 , \9596 );
buf \U$9221 ( \9598 , \455 );
nand \U$9222 ( \9599 , \9597 , \9598 );
not \U$9223 ( \9600 , \454 );
nand \U$9224 ( \9601 , \9600 , \457 );
not \U$9225 ( \9602 , \9601 );
and \U$9226 ( \9603 , \9599 , \9602 );
not \U$9227 ( \9604 , \9599 );
and \U$9228 ( \9605 , \9604 , \9601 );
nor \U$9229 ( \9606 , \9603 , \9605 );
buf \U$9230 ( \9607 , \9606 );
not \U$9231 ( \9608 , \9607 );
not \U$9232 ( \9609 , \9608 );
and \U$9233 ( \9610 , \9609 , RIae79250_140);
not \U$9234 ( \9611 , \9609 );
and \U$9235 ( \9612 , \9611 , \1503 );
nor \U$9236 ( \9613 , \9610 , \9612 );
not \U$9237 ( \9614 , \9613 );
or \U$9238 ( \9615 , \9592 , \9614 );
nand \U$9239 ( \9616 , \1501 , \9419 );
nand \U$9240 ( \9617 , \9615 , \9616 );
not \U$9241 ( \9618 , \9617 );
not \U$9242 ( \9619 , \9618 );
xor \U$9243 ( \9620 , RIae7a510_180, RIae7a600_182);
buf \U$9244 ( \9621 , \9620 );
buf \U$9245 ( \9622 , \9621 );
not \U$9246 ( \9623 , \9622 );
not \U$9247 ( \9624 , \1404 );
not \U$9248 ( \9625 , \9624 );
and \U$9249 ( \9626 , RIae7a3a8_177, \9625 );
not \U$9250 ( \9627 , RIae7a3a8_177);
and \U$9251 ( \9628 , \9627 , \2849 );
nor \U$9252 ( \9629 , \9626 , \9628 );
not \U$9253 ( \9630 , \9629 );
or \U$9254 ( \9631 , \9623 , \9630 );
not \U$9255 ( \9632 , RIae7a3a8_177);
not \U$9256 ( \9633 , \5134 );
or \U$9257 ( \9634 , \9632 , \9633 );
or \U$9258 ( \9635 , \5134 , RIae7a3a8_177);
nand \U$9259 ( \9636 , \9634 , \9635 );
not \U$9260 ( \9637 , \9620 );
and \U$9261 ( \9638 , RIae7a3a8_177, RIae7a600_182);
not \U$9262 ( \9639 , RIae7a3a8_177);
not \U$9263 ( \9640 , RIae7a600_182);
and \U$9264 ( \9641 , \9639 , \9640 );
nor \U$9265 ( \9642 , \9638 , \9641 );
and \U$9266 ( \9643 , \9637 , \9642 );
buf \U$9267 ( \9644 , \9643 );
nand \U$9268 ( \9645 , \9636 , \9644 );
nand \U$9269 ( \9646 , \9631 , \9645 );
not \U$9270 ( \9647 , \9646 );
or \U$9271 ( \9648 , \9619 , \9647 );
or \U$9272 ( \9649 , \9646 , \9618 );
nand \U$9273 ( \9650 , \9648 , \9649 );
not \U$9274 ( \9651 , \9650 );
or \U$9275 ( \9652 , \9591 , \9651 );
nand \U$9276 ( \9653 , \9646 , \9617 );
nand \U$9277 ( \9654 , \9652 , \9653 );
not \U$9278 ( \9655 , \1988 );
not \U$9279 ( \9656 , RIae797f0_152);
buf \U$9280 ( \9657 , \1858 );
not \U$9281 ( \9658 , \9657 );
or \U$9282 ( \9659 , \9656 , \9658 );
or \U$9283 ( \9660 , \1859 , RIae797f0_152);
nand \U$9284 ( \9661 , \9659 , \9660 );
not \U$9285 ( \9662 , \9661 );
or \U$9286 ( \9663 , \9655 , \9662 );
not \U$9287 ( \9664 , RIae797f0_152);
not \U$9288 ( \9665 , \1969 );
or \U$9289 ( \9666 , \9664 , \9665 );
not \U$9290 ( \9667 , \1961 );
not \U$9291 ( \9668 , \1964 );
and \U$9292 ( \9669 , \9667 , \9668 );
and \U$9293 ( \9670 , \1961 , \1964 );
nor \U$9294 ( \9671 , \9669 , \9670 );
buf \U$9295 ( \9672 , \9671 );
not \U$9296 ( \9673 , \9672 );
nand \U$9297 ( \9674 , \9673 , \1991 );
nand \U$9298 ( \9675 , \9666 , \9674 );
nand \U$9299 ( \9676 , \9675 , \2007 );
nand \U$9300 ( \9677 , \9663 , \9676 );
not \U$9301 ( \9678 , \9677 );
not \U$9302 ( \9679 , RIae7a240_174);
not \U$9303 ( \9680 , RIae7a330_176);
and \U$9304 ( \9681 , \9679 , \9680 );
and \U$9305 ( \9682 , RIae7a240_174, RIae7a330_176);
and \U$9306 ( \9683 , RIae7a3a8_177, RIae7a330_176);
not \U$9307 ( \9684 , RIae7a3a8_177);
and \U$9308 ( \9685 , \9684 , \9680 );
nor \U$9309 ( \9686 , \9683 , \9685 );
nor \U$9310 ( \9687 , \9681 , \9682 , \9686 );
buf \U$9311 ( \9688 , \9687 );
not \U$9312 ( \9689 , \9688 );
xnor \U$9313 ( \9690 , RIae7a240_174, \1878 );
not \U$9314 ( \9691 , \9690 );
or \U$9315 ( \9692 , \9689 , \9691 );
not \U$9316 ( \9693 , RIae7a240_174);
not \U$9317 ( \9694 , \2047 );
or \U$9318 ( \9695 , \9693 , \9694 );
not \U$9319 ( \9696 , \3144 );
or \U$9320 ( \9697 , \9696 , RIae7a240_174);
nand \U$9321 ( \9698 , \9695 , \9697 );
buf \U$9322 ( \9699 , \9686 );
nand \U$9323 ( \9700 , \9698 , \9699 );
nand \U$9324 ( \9701 , \9692 , \9700 );
not \U$9325 ( \9702 , \9701 );
nand \U$9326 ( \9703 , \9678 , \9702 );
not \U$9327 ( \9704 , \9703 );
buf \U$9328 ( \9705 , \9478 );
not \U$9329 ( \9706 , \9705 );
not \U$9330 ( \9707 , \9475 );
or \U$9331 ( \9708 , \9706 , \9707 );
and \U$9332 ( \9709 , RIae7a6f0_184, \4413 );
not \U$9333 ( \9710 , RIae7a6f0_184);
buf \U$9334 ( \9711 , \833 );
and \U$9335 ( \9712 , \9710 , \9711 );
or \U$9336 ( \9713 , \9709 , \9712 );
nand \U$9337 ( \9714 , \9713 , \9473 );
nand \U$9338 ( \9715 , \9708 , \9714 );
not \U$9339 ( \9716 , \9715 );
or \U$9340 ( \9717 , \9704 , \9716 );
nand \U$9341 ( \9718 , \9701 , \9677 );
nand \U$9342 ( \9719 , \9717 , \9718 );
nor \U$9343 ( \9720 , \9654 , \9719 );
xor \U$9344 ( \9721 , RIae7a948_189, RIae7a7e0_186);
not \U$9345 ( \9722 , \9721 );
and \U$9346 ( \9723 , RIae7a060_170, RIae7a948_189);
not \U$9347 ( \9724 , RIae7a060_170);
not \U$9348 ( \9725 , RIae7a948_189);
and \U$9349 ( \9726 , \9724 , \9725 );
nor \U$9350 ( \9727 , \9723 , \9726 );
and \U$9351 ( \9728 , \9722 , \9727 );
buf \U$9352 ( \9729 , \9728 );
buf \U$9353 ( \9730 , \9729 );
not \U$9354 ( \9731 , \9730 );
not \U$9355 ( \9732 , RIae7a060_170);
not \U$9356 ( \9733 , \1439 );
or \U$9357 ( \9734 , \9732 , \9733 );
or \U$9358 ( \9735 , \3443 , RIae7a060_170);
nand \U$9359 ( \9736 , \9734 , \9735 );
not \U$9360 ( \9737 , \9736 );
or \U$9361 ( \9738 , \9731 , \9737 );
not \U$9362 ( \9739 , RIae7a060_170);
not \U$9363 ( \9740 , \1288 );
or \U$9364 ( \9741 , \9739 , \9740 );
or \U$9365 ( \9742 , \1288 , RIae7a060_170);
nand \U$9366 ( \9743 , \9741 , \9742 );
buf \U$9367 ( \9744 , \9721 );
buf \U$9368 ( \9745 , \9744 );
nand \U$9369 ( \9746 , \9743 , \9745 );
nand \U$9370 ( \9747 , \9738 , \9746 );
not \U$9371 ( \9748 , \9747 );
not \U$9372 ( \9749 , RIae7a060_170);
not \U$9373 ( \9750 , RIae7a150_172);
and \U$9374 ( \9751 , \9749 , \9750 );
not \U$9375 ( \9752 , RIae7a0d8_171);
and \U$9376 ( \9753 , \9752 , RIae7a060_170);
and \U$9377 ( \9754 , RIae7a0d8_171, RIae7a150_172);
nor \U$9378 ( \9755 , \9751 , \9753 , \9754 );
not \U$9379 ( \9756 , \9755 );
not \U$9380 ( \9757 , \9756 );
buf \U$9381 ( \9758 , \9757 );
not \U$9382 ( \9759 , \9758 );
not \U$9383 ( \9760 , \854 );
not \U$9384 ( \9761 , \9760 );
and \U$9385 ( \9762 , RIae7a150_172, \9761 );
not \U$9386 ( \9763 , RIae7a150_172);
and \U$9387 ( \9764 , \9763 , \2166 );
nor \U$9388 ( \9765 , \9762 , \9764 );
not \U$9389 ( \9766 , \9765 );
or \U$9390 ( \9767 , \9759 , \9766 );
and \U$9391 ( \9768 , RIae7a150_172, \3235 );
not \U$9392 ( \9769 , RIae7a150_172);
not \U$9393 ( \9770 , \936 );
and \U$9394 ( \9771 , \9769 , \9770 );
or \U$9395 ( \9772 , \9768 , \9771 );
nand \U$9396 ( \9773 , \9749 , \9752 );
nand \U$9397 ( \9774 , RIae7a060_170, RIae7a0d8_171);
and \U$9398 ( \9775 , \9773 , \9774 );
buf \U$9399 ( \9776 , \9775 );
buf \U$9400 ( \9777 , \9776 );
nand \U$9401 ( \9778 , \9772 , \9777 );
nand \U$9402 ( \9779 , \9767 , \9778 );
not \U$9403 ( \9780 , \9779 );
or \U$9404 ( \9781 , \9748 , \9780 );
not \U$9405 ( \9782 , RIae7a1c8_173);
and \U$9406 ( \9783 , RIae7a240_174, \9782 );
not \U$9407 ( \9784 , RIae7a240_174);
and \U$9408 ( \9785 , \9784 , RIae7a1c8_173);
nor \U$9409 ( \9786 , \9783 , \9785 );
and \U$9410 ( \9787 , RIae7a2b8_175, RIae7a1c8_173);
not \U$9411 ( \9788 , RIae7a2b8_175);
and \U$9412 ( \9789 , \9788 , \9782 );
nor \U$9413 ( \9790 , \9787 , \9789 );
and \U$9414 ( \9791 , \9786 , \9790 );
buf \U$9415 ( \9792 , \9791 );
not \U$9416 ( \9793 , \9792 );
not \U$9417 ( \9794 , RIae7a2b8_175);
not \U$9418 ( \9795 , \3051 );
or \U$9419 ( \9796 , \9794 , \9795 );
not \U$9420 ( \9797 , \2628 );
not \U$9421 ( \9798 , \9797 );
not \U$9422 ( \9799 , RIae7a2b8_175);
nand \U$9423 ( \9800 , \9798 , \9799 );
nand \U$9424 ( \9801 , \9796 , \9800 );
not \U$9425 ( \9802 , \9801 );
or \U$9426 ( \9803 , \9793 , \9802 );
not \U$9427 ( \9804 , RIae7a2b8_175);
not \U$9428 ( \9805 , \9804 );
not \U$9429 ( \9806 , \1898 );
not \U$9430 ( \9807 , \9806 );
not \U$9431 ( \9808 , \9807 );
or \U$9432 ( \9809 , \9805 , \9808 );
not \U$9433 ( \9810 , RIae7a2b8_175);
or \U$9434 ( \9811 , \1899 , \9810 );
nand \U$9435 ( \9812 , \9809 , \9811 );
not \U$9436 ( \9813 , \9786 );
buf \U$9437 ( \9814 , \9813 );
buf \U$9438 ( \9815 , \9814 );
nand \U$9439 ( \9816 , \9812 , \9815 );
nand \U$9440 ( \9817 , \9803 , \9816 );
not \U$9441 ( \9818 , \9817 );
nand \U$9442 ( \9819 , \9781 , \9818 );
or \U$9443 ( \9820 , \9779 , \9747 );
nand \U$9444 ( \9821 , \9819 , \9820 );
or \U$9445 ( \9822 , \9720 , \9821 );
nand \U$9446 ( \9823 , \9654 , \9719 );
nand \U$9447 ( \9824 , \9822 , \9823 );
not \U$9448 ( \9825 , \9824 );
or \U$9449 ( \9826 , \9575 , \9825 );
or \U$9450 ( \9827 , \9574 , \9824 );
buf \U$9451 ( \9828 , \1932 );
not \U$9452 ( \9829 , \9828 );
not \U$9453 ( \9830 , \4982 );
and \U$9454 ( \9831 , RIae794a8_145, \9830 );
not \U$9455 ( \9832 , RIae794a8_145);
and \U$9456 ( \9833 , \9832 , \3207 );
or \U$9457 ( \9834 , \9831 , \9833 );
not \U$9458 ( \9835 , \9834 );
or \U$9459 ( \9836 , \9829 , \9835 );
not \U$9460 ( \9837 , \3810 );
not \U$9461 ( \9838 , \5673 );
or \U$9462 ( \9839 , \9837 , \9838 );
nand \U$9463 ( \9840 , \2402 , RIae794a8_145);
nand \U$9464 ( \9841 , \9839 , \9840 );
nand \U$9465 ( \9842 , \9841 , \2467 );
nand \U$9466 ( \9843 , \9836 , \9842 );
not \U$9467 ( \9844 , \1086 );
not \U$9468 ( \9845 , \921 );
not \U$9469 ( \9846 , \429 );
not \U$9470 ( \9847 , \9846 );
not \U$9471 ( \9848 , \433 );
not \U$9472 ( \9849 , \539 );
not \U$9473 ( \9850 , \9849 );
not \U$9474 ( \9851 , \534 );
or \U$9475 ( \9852 , \9850 , \9851 );
not \U$9476 ( \9853 , \419 );
nand \U$9477 ( \9854 , \9852 , \9853 );
not \U$9478 ( \9855 , \9854 );
or \U$9479 ( \9856 , \9848 , \9855 );
not \U$9480 ( \9857 , \553 );
nand \U$9481 ( \9858 , \9856 , \9857 );
not \U$9482 ( \9859 , \9858 );
or \U$9483 ( \9860 , \9847 , \9859 );
nand \U$9484 ( \9861 , \9860 , \544 );
nand \U$9485 ( \9862 , \546 , \543 );
not \U$9486 ( \9863 , \9862 );
and \U$9487 ( \9864 , \9861 , \9863 );
not \U$9488 ( \9865 , \9861 );
and \U$9489 ( \9866 , \9865 , \9862 );
nor \U$9490 ( \9867 , \9864 , \9866 );
buf \U$9491 ( \9868 , \9867 );
not \U$9492 ( \9869 , \9868 );
or \U$9493 ( \9870 , \9845 , \9869 );
and \U$9494 ( \9871 , \9861 , \9863 );
not \U$9495 ( \9872 , \9861 );
and \U$9496 ( \9873 , \9872 , \9862 );
or \U$9497 ( \9874 , \9871 , \9873 );
buf \U$9498 ( \9875 , \9874 );
nand \U$9499 ( \9876 , \9875 , RIae78e90_132);
nand \U$9500 ( \9877 , \9870 , \9876 );
not \U$9501 ( \9878 , \9877 );
or \U$9502 ( \9879 , \9844 , \9878 );
not \U$9503 ( \9880 , \435 );
not \U$9504 ( \9881 , \9854 );
or \U$9505 ( \9882 , \9880 , \9881 );
not \U$9506 ( \9883 , \544 );
and \U$9507 ( \9884 , \546 , \9883 );
not \U$9508 ( \9885 , \543 );
nor \U$9509 ( \9886 , \9884 , \9885 );
and \U$9510 ( \9887 , \554 , \9886 );
nand \U$9511 ( \9888 , \9882 , \9887 );
buf \U$9512 ( \9889 , \9888 );
not \U$9513 ( \9890 , \420 );
nand \U$9514 ( \9891 , \9890 , \438 );
and \U$9515 ( \9892 , \9889 , \9891 );
not \U$9516 ( \9893 , \9889 );
not \U$9517 ( \9894 , \9891 );
and \U$9518 ( \9895 , \9893 , \9894 );
nor \U$9519 ( \9896 , \9892 , \9895 );
buf \U$9520 ( \9897 , \9896 );
and \U$9521 ( \9898 , RIae78e90_132, \9897 );
not \U$9522 ( \9899 , RIae78e90_132);
not \U$9523 ( \9900 , \9897 );
and \U$9524 ( \9901 , \9899 , \9900 );
or \U$9525 ( \9902 , \9898 , \9901 );
nand \U$9526 ( \9903 , \9902 , \1072 );
nand \U$9527 ( \9904 , \9879 , \9903 );
not \U$9528 ( \9905 , \1062 );
not \U$9529 ( \9906 , RIae79070_136);
or \U$9530 ( \9907 , RIae771f8_71, RIae77270_72);
not \U$9531 ( \9908 , \9907 );
nor \U$9532 ( \9909 , \420 , \421 );
not \U$9533 ( \9910 , \9909 );
not \U$9534 ( \9911 , \9888 );
or \U$9535 ( \9912 , \9910 , \9911 );
not \U$9536 ( \9913 , \441 );
nand \U$9537 ( \9914 , \9912 , \9913 );
not \U$9538 ( \9915 , \9914 );
or \U$9539 ( \9916 , \9908 , \9915 );
nand \U$9540 ( \9917 , \9916 , \447 );
not \U$9541 ( \9918 , \9917 );
or \U$9542 ( \9919 , \450 , \445 );
not \U$9543 ( \9920 , \9919 );
and \U$9544 ( \9921 , \9918 , \9920 );
and \U$9545 ( \9922 , \9917 , \9919 );
nor \U$9546 ( \9923 , \9921 , \9922 );
not \U$9547 ( \9924 , \9923 );
not \U$9548 ( \9925 , \9924 );
not \U$9549 ( \9926 , \9925 );
or \U$9550 ( \9927 , \9906 , \9926 );
not \U$9551 ( \9928 , \9925 );
nand \U$9552 ( \9929 , \9928 , \1039 );
nand \U$9553 ( \9930 , \9927 , \9929 );
not \U$9554 ( \9931 , \9930 );
or \U$9555 ( \9932 , \9905 , \9931 );
not \U$9556 ( \9933 , RIae79070_136);
nand \U$9557 ( \9934 , \9593 , \9598 );
and \U$9558 ( \9935 , \9595 , \9934 );
not \U$9559 ( \9936 , \9595 );
not \U$9560 ( \9937 , \9934 );
and \U$9561 ( \9938 , \9936 , \9937 );
nor \U$9562 ( \9939 , \9935 , \9938 );
not \U$9563 ( \9940 , \9939 );
not \U$9564 ( \9941 , \9940 );
not \U$9565 ( \9942 , \9941 );
or \U$9566 ( \9943 , \9933 , \9942 );
not \U$9567 ( \9944 , \9941 );
nand \U$9568 ( \9945 , \9944 , \1039 );
nand \U$9569 ( \9946 , \9943 , \9945 );
buf \U$9570 ( \9947 , \1049 );
nand \U$9571 ( \9948 , \9946 , \9947 );
nand \U$9572 ( \9949 , \9932 , \9948 );
xor \U$9573 ( \9950 , \9904 , \9949 );
xor \U$9574 ( \9951 , \9843 , \9950 );
not \U$9575 ( \9952 , \9295 );
not \U$9576 ( \9953 , \9372 );
or \U$9577 ( \9954 , \9952 , \9953 );
or \U$9578 ( \9955 , \9372 , \9295 );
nand \U$9579 ( \9956 , \9955 , \9322 );
nand \U$9580 ( \9957 , \9954 , \9956 );
and \U$9581 ( \9958 , \9951 , \9957 );
not \U$9582 ( \9959 , \9951 );
not \U$9583 ( \9960 , \9957 );
and \U$9584 ( \9961 , \9959 , \9960 );
or \U$9585 ( \9962 , \9958 , \9961 );
and \U$9586 ( \9963 , \9463 , \9421 );
or \U$9587 ( \9964 , \9480 , \9963 );
or \U$9588 ( \9965 , \9463 , \9421 );
nand \U$9589 ( \9966 , \9964 , \9965 );
not \U$9590 ( \9967 , \9966 );
not \U$9591 ( \9968 , \9967 );
and \U$9592 ( \9969 , \9962 , \9968 );
not \U$9593 ( \9970 , \9962 );
and \U$9594 ( \9971 , \9970 , \9967 );
nor \U$9595 ( \9972 , \9969 , \9971 );
nand \U$9596 ( \9973 , \9827 , \9972 );
nand \U$9597 ( \9974 , \9826 , \9973 );
not \U$9598 ( \9975 , \951 );
not \U$9599 ( \9976 , \431 );
not \U$9600 ( \9977 , \9976 );
buf \U$9601 ( \9978 , \9854 );
not \U$9602 ( \9979 , \9978 );
or \U$9603 ( \9980 , \9977 , \9979 );
nand \U$9604 ( \9981 , \9980 , \550 );
not \U$9605 ( \9982 , \549 );
nand \U$9606 ( \9983 , \9982 , \552 );
and \U$9607 ( \9984 , \9981 , \9983 );
not \U$9608 ( \9985 , \9981 );
not \U$9609 ( \9986 , \9983 );
and \U$9610 ( \9987 , \9985 , \9986 );
nor \U$9611 ( \9988 , \9984 , \9987 );
buf \U$9612 ( \9989 , \9988 );
xnor \U$9613 ( \9990 , \9989 , RIae78bc0_126);
not \U$9614 ( \9991 , \9990 );
or \U$9615 ( \9992 , \9975 , \9991 );
buf \U$9616 ( \9993 , \9858 );
nand \U$9617 ( \9994 , \9846 , \544 );
and \U$9618 ( \9995 , \9993 , \9994 );
not \U$9619 ( \9996 , \9993 );
not \U$9620 ( \9997 , \9994 );
and \U$9621 ( \9998 , \9996 , \9997 );
nor \U$9622 ( \9999 , \9995 , \9998 );
buf \U$9623 ( \10000 , \9999 );
and \U$9624 ( \10001 , RIae78bc0_126, \10000 );
not \U$9625 ( \10002 , RIae78bc0_126);
and \U$9626 ( \10003 , \9993 , \9997 );
not \U$9627 ( \10004 , \9993 );
and \U$9628 ( \10005 , \10004 , \9994 );
nor \U$9629 ( \10006 , \10003 , \10005 );
buf \U$9630 ( \10007 , \10006 );
and \U$9631 ( \10008 , \10002 , \10007 );
or \U$9632 ( \10009 , \10001 , \10008 );
nand \U$9633 ( \10010 , \10009 , \926 );
nand \U$9634 ( \10011 , \9992 , \10010 );
not \U$9635 ( \10012 , \867 );
not \U$9636 ( \10013 , \402 );
not \U$9637 ( \10014 , \10013 );
not \U$9638 ( \10015 , \538 );
buf \U$9639 ( \10016 , \534 );
not \U$9640 ( \10017 , \10016 );
or \U$9641 ( \10018 , \10015 , \10017 );
not \U$9642 ( \10019 , \410 );
nand \U$9643 ( \10020 , \10018 , \10019 );
not \U$9644 ( \10021 , \10020 );
or \U$9645 ( \10022 , \10014 , \10021 );
nand \U$9646 ( \10023 , \10022 , \414 );
not \U$9647 ( \10024 , \416 );
nor \U$9648 ( \10025 , \10024 , \413 );
and \U$9649 ( \10026 , \10023 , \10025 );
not \U$9650 ( \10027 , \10023 );
not \U$9651 ( \10028 , \10025 );
and \U$9652 ( \10029 , \10027 , \10028 );
nor \U$9653 ( \10030 , \10026 , \10029 );
buf \U$9654 ( \10031 , \10030 );
buf \U$9655 ( \10032 , \10031 );
and \U$9656 ( \10033 , \10032 , RIae78b48_125);
not \U$9657 ( \10034 , \10032 );
and \U$9658 ( \10035 , \10034 , \860 );
nor \U$9659 ( \10036 , \10033 , \10035 );
not \U$9660 ( \10037 , \10036 );
or \U$9661 ( \10038 , \10012 , \10037 );
not \U$9662 ( \10039 , \860 );
nand \U$9663 ( \10040 , \10013 , \414 );
xnor \U$9664 ( \10041 , \10020 , \10040 );
buf \U$9665 ( \10042 , \10041 );
buf \U$9666 ( \10043 , \10042 );
not \U$9667 ( \10044 , \10043 );
or \U$9668 ( \10045 , \10039 , \10044 );
not \U$9669 ( \10046 , \10042 );
not \U$9670 ( \10047 , \10046 );
or \U$9671 ( \10048 , \10047 , \860 );
nand \U$9672 ( \10049 , \10045 , \10048 );
nand \U$9673 ( \10050 , \10049 , \892 );
nand \U$9674 ( \10051 , \10038 , \10050 );
xor \U$9675 ( \10052 , \10011 , \10051 );
not \U$9676 ( \10053 , \797 );
not \U$9677 ( \10054 , \9890 );
not \U$9678 ( \10055 , \9888 );
or \U$9679 ( \10056 , \10054 , \10055 );
buf \U$9680 ( \10057 , \438 );
nand \U$9681 ( \10058 , \10056 , \10057 );
not \U$9682 ( \10059 , \440 );
nor \U$9683 ( \10060 , \10059 , \437 );
and \U$9684 ( \10061 , \10058 , \10060 );
not \U$9685 ( \10062 , \10058 );
not \U$9686 ( \10063 , \10060 );
and \U$9687 ( \10064 , \10062 , \10063 );
nor \U$9688 ( \10065 , \10061 , \10064 );
buf \U$9689 ( \10066 , \10065 );
not \U$9690 ( \10067 , \10066 );
and \U$9691 ( \10068 , RIae78f80_134, \10067 );
not \U$9692 ( \10069 , RIae78f80_134);
buf \U$9693 ( \10070 , \10065 );
not \U$9694 ( \10071 , \10070 );
not \U$9695 ( \10072 , \10071 );
and \U$9696 ( \10073 , \10069 , \10072 );
or \U$9697 ( \10074 , \10068 , \10073 );
not \U$9698 ( \10075 , \10074 );
or \U$9699 ( \10076 , \10053 , \10075 );
nand \U$9700 ( \10077 , \9907 , \447 );
and \U$9701 ( \10078 , \9914 , \10077 );
not \U$9702 ( \10079 , \9914 );
not \U$9703 ( \10080 , \10077 );
and \U$9704 ( \10081 , \10079 , \10080 );
nor \U$9705 ( \10082 , \10078 , \10081 );
buf \U$9706 ( \10083 , \10082 );
buf \U$9707 ( \10084 , \10083 );
and \U$9708 ( \10085 , RIae78f80_134, \10084 );
not \U$9709 ( \10086 , RIae78f80_134);
not \U$9710 ( \10087 , \10084 );
and \U$9711 ( \10088 , \10086 , \10087 );
or \U$9712 ( \10089 , \10085 , \10088 );
nand \U$9713 ( \10090 , \10089 , \838 );
nand \U$9714 ( \10091 , \10076 , \10090 );
and \U$9715 ( \10092 , \10052 , \10091 );
and \U$9716 ( \10093 , \10011 , \10051 );
nor \U$9717 ( \10094 , \10092 , \10093 );
not \U$9718 ( \10095 , \10094 );
not \U$9719 ( \10096 , \2007 );
not \U$9720 ( \10097 , RIae797f0_152);
not \U$9721 ( \10098 , \3417 );
or \U$9722 ( \10099 , \10097 , \10098 );
or \U$9723 ( \10100 , \2564 , RIae797f0_152);
nand \U$9724 ( \10101 , \10099 , \10100 );
not \U$9725 ( \10102 , \10101 );
or \U$9726 ( \10103 , \10096 , \10102 );
and \U$9727 ( \10104 , RIae797f0_152, \2785 );
not \U$9728 ( \10105 , RIae797f0_152);
and \U$9729 ( \10106 , \10105 , \2093 );
or \U$9730 ( \10107 , \10104 , \10106 );
nand \U$9731 ( \10108 , \10107 , \1988 );
nand \U$9732 ( \10109 , \10103 , \10108 );
not \U$9733 ( \10110 , \10109 );
and \U$9734 ( \10111 , \10095 , \10110 );
and \U$9735 ( \10112 , \10109 , \10094 );
nor \U$9736 ( \10113 , \10111 , \10112 );
not \U$9737 ( \10114 , \9950 );
not \U$9738 ( \10115 , \9843 );
or \U$9739 ( \10116 , \10114 , \10115 );
nand \U$9740 ( \10117 , \9949 , \9904 );
nand \U$9741 ( \10118 , \10116 , \10117 );
xor \U$9742 ( \10119 , \10113 , \10118 );
not \U$9743 ( \10120 , \10119 );
not \U$9744 ( \10121 , \9966 );
not \U$9745 ( \10122 , \9960 );
or \U$9746 ( \10123 , \10121 , \10122 );
nand \U$9747 ( \10124 , \10123 , \9951 );
nand \U$9748 ( \10125 , \9967 , \9957 );
nand \U$9749 ( \10126 , \10124 , \10125 );
not \U$9750 ( \10127 , \10126 );
or \U$9751 ( \10128 , \10120 , \10127 );
or \U$9752 ( \10129 , \10126 , \10119 );
nand \U$9753 ( \10130 , \10128 , \10129 );
not \U$9754 ( \10131 , \10130 );
not \U$9755 ( \10132 , \926 );
not \U$9756 ( \10133 , \9990 );
or \U$9757 ( \10134 , \10132 , \10133 );
buf \U$9758 ( \10135 , \9978 );
nand \U$9759 ( \10136 , \9976 , \550 );
not \U$9760 ( \10137 , \10136 );
and \U$9761 ( \10138 , \10135 , \10137 );
not \U$9762 ( \10139 , \10135 );
and \U$9763 ( \10140 , \10139 , \10136 );
nor \U$9764 ( \10141 , \10138 , \10140 );
buf \U$9765 ( \10142 , \10141 );
and \U$9766 ( \10143 , RIae78bc0_126, \10142 );
not \U$9767 ( \10144 , RIae78bc0_126);
and \U$9768 ( \10145 , \10135 , \10136 );
not \U$9769 ( \10146 , \10135 );
and \U$9770 ( \10147 , \10146 , \10137 );
nor \U$9771 ( \10148 , \10145 , \10147 );
buf \U$9772 ( \10149 , \10148 );
and \U$9773 ( \10150 , \10144 , \10149 );
nor \U$9774 ( \10151 , \10143 , \10150 );
nand \U$9775 ( \10152 , \10151 , \951 );
nand \U$9776 ( \10153 , \10134 , \10152 );
not \U$9777 ( \10154 , \1072 );
not \U$9778 ( \10155 , \9877 );
or \U$9779 ( \10156 , \10154 , \10155 );
and \U$9780 ( \10157 , RIae78e90_132, \10007 );
not \U$9781 ( \10158 , RIae78e90_132);
and \U$9782 ( \10159 , \10158 , \10000 );
nor \U$9783 ( \10160 , \10157 , \10159 );
nand \U$9784 ( \10161 , \10160 , \1086 );
nand \U$9785 ( \10162 , \10156 , \10161 );
or \U$9786 ( \10163 , \10153 , \10162 );
not \U$9787 ( \10164 , \839 );
not \U$9788 ( \10165 , \10074 );
or \U$9789 ( \10166 , \10164 , \10165 );
not \U$9790 ( \10167 , RIae78f80_134);
buf \U$9791 ( \10168 , \9896 );
not \U$9792 ( \10169 , \10168 );
or \U$9793 ( \10170 , \10167 , \10169 );
buf \U$9794 ( \10171 , \9897 );
or \U$9795 ( \10172 , \10171 , RIae78f80_134);
nand \U$9796 ( \10173 , \10170 , \10172 );
nand \U$9797 ( \10174 , \10173 , \797 );
nand \U$9798 ( \10175 , \10166 , \10174 );
nand \U$9799 ( \10176 , \10163 , \10175 );
nand \U$9800 ( \10177 , \10153 , \10162 );
nand \U$9801 ( \10178 , \10176 , \10177 );
not \U$9802 ( \10179 , \10178 );
buf \U$9803 ( \10180 , \536 );
not \U$9804 ( \10181 , \10180 );
not \U$9805 ( \10182 , \10181 );
not \U$9806 ( \10183 , \10016 );
or \U$9807 ( \10184 , \10182 , \10183 );
buf \U$9808 ( \10185 , \406 );
nand \U$9809 ( \10186 , \10184 , \10185 );
xor \U$9810 ( \10187 , RIae77978_87, RIae779f0_88);
and \U$9811 ( \10188 , \10186 , \10187 );
not \U$9812 ( \10189 , \10186 );
not \U$9813 ( \10190 , \10187 );
and \U$9814 ( \10191 , \10189 , \10190 );
nor \U$9815 ( \10192 , \10188 , \10191 );
buf \U$9816 ( \10193 , \10192 );
not \U$9817 ( \10194 , \10193 );
not \U$9818 ( \10195 , \10194 );
nand \U$9819 ( \10196 , \10195 , RIae78b48_125);
not \U$9820 ( \10197 , \10051 );
and \U$9821 ( \10198 , \10196 , \10197 );
not \U$9822 ( \10199 , \10196 );
and \U$9823 ( \10200 , \10199 , \10051 );
or \U$9824 ( \10201 , \10198 , \10200 );
not \U$9825 ( \10202 , \10201 );
not \U$9826 ( \10203 , \1049 );
not \U$9827 ( \10204 , \9930 );
or \U$9828 ( \10205 , \10203 , \10204 );
not \U$9829 ( \10206 , \1039 );
not \U$9830 ( \10207 , \10083 );
buf \U$9831 ( \10208 , \10207 );
not \U$9832 ( \10209 , \10208 );
or \U$9833 ( \10210 , \10206 , \10209 );
nand \U$9834 ( \10211 , \10084 , RIae79070_136);
nand \U$9835 ( \10212 , \10210 , \10211 );
nand \U$9836 ( \10213 , \10212 , \1062 );
nand \U$9837 ( \10214 , \10205 , \10213 );
not \U$9838 ( \10215 , \10214 );
or \U$9839 ( \10216 , \10202 , \10215 );
not \U$9840 ( \10217 , \10196 );
nand \U$9841 ( \10218 , \10217 , \10197 );
nand \U$9842 ( \10219 , \10216 , \10218 );
not \U$9843 ( \10220 , \10219 );
nand \U$9844 ( \10221 , \10179 , \10220 );
not \U$9845 ( \10222 , \10221 );
buf \U$9846 ( \10223 , \2162 );
not \U$9847 ( \10224 , \10223 );
not \U$9848 ( \10225 , \2183 );
buf \U$9849 ( \10226 , \4959 );
not \U$9850 ( \10227 , \10226 );
not \U$9851 ( \10228 , \10227 );
or \U$9852 ( \10229 , \10225 , \10228 );
nand \U$9853 ( \10230 , \4960 , RIae79520_146);
nand \U$9854 ( \10231 , \10229 , \10230 );
not \U$9855 ( \10232 , \10231 );
or \U$9856 ( \10233 , \10224 , \10232 );
not \U$9857 ( \10234 , \2183 );
not \U$9858 ( \10235 , \5109 );
or \U$9859 ( \10236 , \10234 , \10235 );
not \U$9860 ( \10237 , \6256 );
nand \U$9861 ( \10238 , \10237 , RIae79520_146);
nand \U$9862 ( \10239 , \10236 , \10238 );
nand \U$9863 ( \10240 , \10239 , \2602 );
nand \U$9864 ( \10241 , \10233 , \10240 );
buf \U$9865 ( \10242 , \518 );
nand \U$9866 ( \10243 , RIae775b8_79, RIae77630_80);
or \U$9867 ( \10244 , \10242 , \10243 );
nand \U$9868 ( \10245 , RIae774c8_77, RIae77540_78);
nand \U$9869 ( \10246 , \10244 , \10245 );
not \U$9870 ( \10247 , \10246 );
not \U$9871 ( \10248 , \519 );
not \U$9872 ( \10249 , \10248 );
or \U$9873 ( \10250 , \10247 , \10249 );
nand \U$9874 ( \10251 , RIae776a8_81, RIae77720_82);
nand \U$9875 ( \10252 , \10250 , \10251 );
xor \U$9876 ( \10253 , RIae773d8_75, RIae77450_76);
not \U$9877 ( \10254 , \10253 );
and \U$9878 ( \10255 , \10252 , \10254 );
not \U$9879 ( \10256 , \10252 );
and \U$9880 ( \10257 , \10256 , \10253 );
nor \U$9881 ( \10258 , \10255 , \10257 );
buf \U$9882 ( \10259 , \10258 );
or \U$9883 ( \10260 , \10259 , \860 );
not \U$9884 ( \10261 , \10260 );
not \U$9885 ( \10262 , \10185 );
nor \U$9886 ( \10263 , \10262 , \10180 );
not \U$9887 ( \10264 , \10263 );
not \U$9888 ( \10265 , \10016 );
not \U$9889 ( \10266 , \10265 );
or \U$9890 ( \10267 , \10264 , \10266 );
not \U$9891 ( \10268 , \10263 );
not \U$9892 ( \10269 , \10265 );
nand \U$9893 ( \10270 , \10268 , \10269 );
nand \U$9894 ( \10271 , \10267 , \10270 );
buf \U$9895 ( \10272 , \10271 );
nand \U$9896 ( \10273 , \10272 , RIae78b48_125);
xor \U$9897 ( \10274 , RIae7a9c0_190, RIae7aa38_191);
buf \U$9898 ( \10275 , \10274 );
not \U$9899 ( \10276 , \10275 );
not \U$9900 ( \10277 , \10276 );
and \U$9901 ( \10278 , RIae7a8d0_188, RIae7a9c0_190);
nor \U$9902 ( \10279 , RIae7a8d0_188, RIae7a9c0_190);
nor \U$9903 ( \10280 , \10278 , \10274 , \10279 );
not \U$9904 ( \10281 , \10280 );
not \U$9905 ( \10282 , \10281 );
or \U$9906 ( \10283 , \10277 , \10282 );
nand \U$9907 ( \10284 , \10283 , RIae7a8d0_188);
xor \U$9908 ( \10285 , \10273 , \10284 );
not \U$9909 ( \10286 , \10285 );
and \U$9910 ( \10287 , \10261 , \10286 );
not \U$9911 ( \10288 , \10273 );
and \U$9912 ( \10289 , \10288 , \10284 );
nor \U$9913 ( \10290 , \10287 , \10289 );
not \U$9914 ( \10291 , \10290 );
or \U$9915 ( \10292 , \10241 , \10291 );
not \U$9916 ( \10293 , \2467 );
not \U$9917 ( \10294 , \9834 );
or \U$9918 ( \10295 , \10293 , \10294 );
not \U$9919 ( \10296 , \3810 );
not \U$9920 ( \10297 , \4169 );
or \U$9921 ( \10298 , \10296 , \10297 );
nand \U$9922 ( \10299 , \6242 , RIae794a8_145);
nand \U$9923 ( \10300 , \10298 , \10299 );
nand \U$9924 ( \10301 , \10300 , \9828 );
nand \U$9925 ( \10302 , \10295 , \10301 );
nand \U$9926 ( \10303 , \10292 , \10302 );
nand \U$9927 ( \10304 , \10291 , \10241 );
nand \U$9928 ( \10305 , \10303 , \10304 );
not \U$9929 ( \10306 , \10305 );
or \U$9930 ( \10307 , \10222 , \10306 );
nand \U$9931 ( \10308 , \10219 , \10178 );
nand \U$9932 ( \10309 , \10307 , \10308 );
not \U$9933 ( \10310 , \10309 );
not \U$9934 ( \10311 , \10310 );
and \U$9935 ( \10312 , \10131 , \10311 );
and \U$9936 ( \10313 , \10130 , \10310 );
nor \U$9937 ( \10314 , \10312 , \10313 );
xor \U$9938 ( \10315 , \9974 , \10314 );
not \U$9939 ( \10316 , \5950 );
not \U$9940 ( \10317 , RIae79520_146);
not \U$9941 ( \10318 , \6242 );
or \U$9942 ( \10319 , \10317 , \10318 );
nand \U$9943 ( \10320 , \4653 , \4168 );
nand \U$9944 ( \10321 , \10319 , \10320 );
not \U$9945 ( \10322 , \10321 );
or \U$9946 ( \10323 , \10316 , \10322 );
not \U$9947 ( \10324 , \3153 );
not \U$9948 ( \10325 , \3202 );
or \U$9949 ( \10326 , \10324 , \10325 );
or \U$9950 ( \10327 , \3153 , \3202 );
nand \U$9951 ( \10328 , \10326 , \10327 );
and \U$9952 ( \10329 , RIae79520_146, \10328 );
not \U$9953 ( \10330 , RIae79520_146);
not \U$9954 ( \10331 , \10328 );
and \U$9955 ( \10332 , \10330 , \10331 );
nor \U$9956 ( \10333 , \10329 , \10332 );
nand \U$9957 ( \10334 , \10333 , \10223 );
nand \U$9958 ( \10335 , \10323 , \10334 );
not \U$9959 ( \10336 , \10335 );
not \U$9960 ( \10337 , \10031 );
not \U$9961 ( \10338 , \10337 );
nand \U$9962 ( \10339 , \10338 , RIae78b48_125);
not \U$9963 ( \10340 , \926 );
not \U$9964 ( \10341 , \1286 );
not \U$9965 ( \10342 , \9868 );
or \U$9966 ( \10343 , \10341 , \10342 );
nand \U$9967 ( \10344 , \9875 , RIae78bc0_126);
nand \U$9968 ( \10345 , \10343 , \10344 );
not \U$9969 ( \10346 , \10345 );
or \U$9970 ( \10347 , \10340 , \10346 );
nand \U$9971 ( \10348 , \10009 , \951 );
nand \U$9972 ( \10349 , \10347 , \10348 );
xor \U$9973 ( \10350 , \10339 , \10349 );
not \U$9974 ( \10351 , \10350 );
not \U$9975 ( \10352 , \10351 );
and \U$9976 ( \10353 , \10336 , \10352 );
and \U$9977 ( \10354 , \10335 , \10351 );
nor \U$9978 ( \10355 , \10353 , \10354 );
not \U$9979 ( \10356 , \10355 );
not \U$9980 ( \10357 , \10356 );
not \U$9981 ( \10358 , \9403 );
not \U$9982 ( \10359 , \9400 );
or \U$9983 ( \10360 , \10358 , \10359 );
not \U$9984 ( \10361 , \9455 );
and \U$9985 ( \10362 , RIae79250_140, \10361 );
not \U$9986 ( \10363 , RIae79250_140);
and \U$9987 ( \10364 , \10363 , \9459 );
or \U$9988 ( \10365 , \10362 , \10364 );
nand \U$9989 ( \10366 , \10365 , \1501 );
nand \U$9990 ( \10367 , \10360 , \10366 );
not \U$9991 ( \10368 , \10367 );
not \U$9992 ( \10369 , \10368 );
not \U$9993 ( \10370 , \1910 );
not \U$9994 ( \10371 , \9444 );
or \U$9995 ( \10372 , \10370 , \10371 );
and \U$9996 ( \10373 , RIae793b8_143, \9364 );
not \U$9997 ( \10374 , RIae793b8_143);
and \U$9998 ( \10375 , \10374 , \9367 );
or \U$9999 ( \10376 , \10373 , \10375 );
nand \U$10000 ( \10377 , \10376 , \1864 );
nand \U$10001 ( \10378 , \10372 , \10377 );
not \U$10002 ( \10379 , \10378 );
not \U$10003 ( \10380 , \10379 );
or \U$10004 ( \10381 , \10369 , \10380 );
not \U$10005 ( \10382 , \2063 );
not \U$10006 ( \10383 , \9352 );
or \U$10007 ( \10384 , \10382 , \10383 );
not \U$10008 ( \10385 , \2056 );
not \U$10009 ( \10386 , \9316 );
not \U$10010 ( \10387 , \10386 );
or \U$10011 ( \10388 , \10385 , \10387 );
nand \U$10012 ( \10389 , \9313 , RIae79610_148);
nand \U$10013 ( \10390 , \10388 , \10389 );
nand \U$10014 ( \10391 , \10390 , \2011 );
nand \U$10015 ( \10392 , \10384 , \10391 );
nand \U$10016 ( \10393 , \10381 , \10392 );
nand \U$10017 ( \10394 , \10378 , \10367 );
nand \U$10018 ( \10395 , \10393 , \10394 );
not \U$10019 ( \10396 , \10395 );
not \U$10020 ( \10397 , \10396 );
or \U$10021 ( \10398 , \10357 , \10397 );
nand \U$10022 ( \10399 , \10395 , \10355 );
nand \U$10023 ( \10400 , \10398 , \10399 );
buf \U$10024 ( \10401 , \1843 );
not \U$10025 ( \10402 , \10401 );
not \U$10026 ( \10403 , \9303 );
or \U$10027 ( \10404 , \10402 , \10403 );
not \U$10028 ( \10405 , RIae79688_149);
not \U$10029 ( \10406 , \9289 );
not \U$10030 ( \10407 , \10406 );
or \U$10031 ( \10408 , \10405 , \10407 );
not \U$10032 ( \10409 , \6345 );
or \U$10033 ( \10410 , \10409 , RIae79688_149);
nand \U$10034 ( \10411 , \10408 , \10410 );
nand \U$10035 ( \10412 , \10411 , \1820 );
nand \U$10036 ( \10413 , \10404 , \10412 );
not \U$10037 ( \10414 , \2250 );
not \U$10038 ( \10415 , \10414 );
not \U$10039 ( \10416 , RIae79ac0_158);
not \U$10040 ( \10417 , \6257 );
or \U$10041 ( \10418 , \10416 , \10417 );
not \U$10042 ( \10419 , RIae79ac0_158);
nand \U$10043 ( \10420 , \6256 , \10419 );
nand \U$10044 ( \10421 , \10418 , \10420 );
not \U$10045 ( \10422 , \10421 );
or \U$10046 ( \10423 , \10415 , \10422 );
nand \U$10047 ( \10424 , \9282 , \2272 );
nand \U$10048 ( \10425 , \10423 , \10424 );
xor \U$10049 ( \10426 , \10413 , \10425 );
not \U$10050 ( \10427 , \5950 );
not \U$10051 ( \10428 , \10231 );
or \U$10052 ( \10429 , \10427 , \10428 );
nand \U$10053 ( \10430 , \10321 , \10223 );
nand \U$10054 ( \10431 , \10429 , \10430 );
and \U$10055 ( \10432 , \10426 , \10431 );
and \U$10056 ( \10433 , \10413 , \10425 );
or \U$10057 ( \10434 , \10432 , \10433 );
not \U$10058 ( \10435 , \10434 );
and \U$10059 ( \10436 , \10400 , \10435 );
not \U$10060 ( \10437 , \10400 );
and \U$10061 ( \10438 , \10437 , \10434 );
nor \U$10062 ( \10439 , \10436 , \10438 );
not \U$10063 ( \10440 , \9687 );
not \U$10064 ( \10441 , \9698 );
or \U$10065 ( \10442 , \10440 , \10441 );
not \U$10066 ( \10443 , RIae7a240_174);
not \U$10067 ( \10444 , \2025 );
not \U$10068 ( \10445 , \10444 );
or \U$10069 ( \10446 , \10443 , \10445 );
or \U$10070 ( \10447 , \10444 , RIae7a240_174);
nand \U$10071 ( \10448 , \10446 , \10447 );
nand \U$10072 ( \10449 , \10448 , \9699 );
nand \U$10073 ( \10450 , \10442 , \10449 );
buf \U$10074 ( \10451 , \1012 );
not \U$10075 ( \10452 , \10451 );
not \U$10076 ( \10453 , \9607 );
and \U$10077 ( \10454 , \10453 , \997 );
not \U$10078 ( \10455 , \10453 );
and \U$10079 ( \10456 , \10455 , RIae79160_138);
nor \U$10080 ( \10457 , \10454 , \10456 );
not \U$10081 ( \10458 , \10457 );
or \U$10082 ( \10459 , \10452 , \10458 );
not \U$10083 ( \10460 , RIae79160_138);
buf \U$10084 ( \10461 , \9939 );
not \U$10085 ( \10462 , \10461 );
or \U$10086 ( \10463 , \10460 , \10462 );
not \U$10087 ( \10464 , \9940 );
not \U$10088 ( \10465 , \10464 );
nand \U$10089 ( \10466 , \10465 , \997 );
nand \U$10090 ( \10467 , \10463 , \10466 );
nand \U$10091 ( \10468 , \10467 , \1008 );
nand \U$10092 ( \10469 , \10459 , \10468 );
or \U$10093 ( \10470 , \10450 , \10469 );
not \U$10094 ( \10471 , \2007 );
xnor \U$10095 ( \10472 , RIae797f0_152, \1954 );
not \U$10096 ( \10473 , \10472 );
or \U$10097 ( \10474 , \10471 , \10473 );
nand \U$10098 ( \10475 , \9675 , \1989 );
nand \U$10099 ( \10476 , \10474 , \10475 );
nand \U$10100 ( \10477 , \10470 , \10476 );
nand \U$10101 ( \10478 , \10450 , \10469 );
nand \U$10102 ( \10479 , \10477 , \10478 );
xor \U$10103 ( \10480 , \10052 , \10091 );
or \U$10104 ( \10481 , \10479 , \10480 );
not \U$10105 ( \10482 , \10481 );
not \U$10106 ( \10483 , \2322 );
not \U$10107 ( \10484 , RIae798e0_154);
not \U$10108 ( \10485 , \9657 );
or \U$10109 ( \10486 , \10484 , \10485 );
or \U$10110 ( \10487 , \1859 , RIae798e0_154);
nand \U$10111 ( \10488 , \10486 , \10487 );
not \U$10112 ( \10489 , \10488 );
or \U$10113 ( \10490 , \10483 , \10489 );
not \U$10114 ( \10491 , RIae798e0_154);
not \U$10115 ( \10492 , \3269 );
not \U$10116 ( \10493 , \10492 );
or \U$10117 ( \10494 , \10491 , \10493 );
or \U$10118 ( \10495 , \3270 , RIae798e0_154);
nand \U$10119 ( \10496 , \10494 , \10495 );
nand \U$10120 ( \10497 , \10496 , \2340 );
nand \U$10121 ( \10498 , \10490 , \10497 );
not \U$10122 ( \10499 , \9814 );
not \U$10123 ( \10500 , RIae7a2b8_175);
not \U$10124 ( \10501 , \1878 );
or \U$10125 ( \10502 , \10500 , \10501 );
or \U$10126 ( \10503 , \1878 , RIae7a2b8_175);
nand \U$10127 ( \10504 , \10502 , \10503 );
not \U$10128 ( \10505 , \10504 );
or \U$10129 ( \10506 , \10499 , \10505 );
nand \U$10130 ( \10507 , \9812 , \9792 );
nand \U$10131 ( \10508 , \10506 , \10507 );
xor \U$10132 ( \10509 , \10498 , \10508 );
buf \U$10133 ( \10510 , \9549 );
not \U$10134 ( \10511 , \10510 );
not \U$10135 ( \10512 , \9534 );
or \U$10136 ( \10513 , \10511 , \10512 );
not \U$10137 ( \10514 , RIae7a7e0_186);
not \U$10138 ( \10515 , \4413 );
or \U$10139 ( \10516 , \10514 , \10515 );
or \U$10140 ( \10517 , \827 , RIae7a7e0_186);
nand \U$10141 ( \10518 , \10516 , \10517 );
buf \U$10142 ( \10519 , \9527 );
nand \U$10143 ( \10520 , \10518 , \10519 );
nand \U$10144 ( \10521 , \10513 , \10520 );
and \U$10145 ( \10522 , \10509 , \10521 );
and \U$10146 ( \10523 , \10498 , \10508 );
or \U$10147 ( \10524 , \10522 , \10523 );
not \U$10148 ( \10525 , \10524 );
or \U$10149 ( \10526 , \10482 , \10525 );
nand \U$10150 ( \10527 , \10479 , \10480 );
nand \U$10151 ( \10528 , \10526 , \10527 );
xor \U$10152 ( \10529 , \10439 , \10528 );
not \U$10153 ( \10530 , \6091 );
not \U$10154 ( \10531 , RIae79d90_164);
not \U$10155 ( \10532 , \2286 );
or \U$10156 ( \10533 , \10531 , \10532 );
buf \U$10157 ( \10534 , \2285 );
or \U$10158 ( \10535 , \10534 , RIae79d90_164);
nand \U$10159 ( \10536 , \10533 , \10535 );
not \U$10160 ( \10537 , \10536 );
or \U$10161 ( \10538 , \10530 , \10537 );
xor \U$10162 ( \10539 , \2308 , RIae79d90_164);
nand \U$10163 ( \10540 , \10539 , \5048 );
nand \U$10164 ( \10541 , \10538 , \10540 );
buf \U$10165 ( \10542 , \9744 );
not \U$10166 ( \10543 , \10542 );
and \U$10167 ( \10544 , \1137 , \1139 );
not \U$10168 ( \10545 , \1137 );
not \U$10169 ( \10546 , \1139 );
and \U$10170 ( \10547 , \10545 , \10546 );
nor \U$10171 ( \10548 , \10544 , \10547 );
and \U$10172 ( \10549 , RIae7a060_170, \10548 );
not \U$10173 ( \10550 , RIae7a060_170);
not \U$10174 ( \10551 , \10548 );
and \U$10175 ( \10552 , \10550 , \10551 );
or \U$10176 ( \10553 , \10549 , \10552 );
not \U$10177 ( \10554 , \10553 );
or \U$10178 ( \10555 , \10543 , \10554 );
nand \U$10179 ( \10556 , \9743 , \9729 );
nand \U$10180 ( \10557 , \10555 , \10556 );
xor \U$10181 ( \10558 , \10541 , \10557 );
not \U$10182 ( \10559 , \6201 );
not \U$10183 ( \10560 , \9557 );
or \U$10184 ( \10561 , \10559 , \10560 );
not \U$10185 ( \10562 , \2128 );
not \U$10186 ( \10563 , \2130 );
and \U$10187 ( \10564 , \10562 , \10563 );
and \U$10188 ( \10565 , \2128 , \2130 );
nor \U$10189 ( \10566 , \10564 , \10565 );
not \U$10190 ( \10567 , \10566 );
and \U$10191 ( \10568 , RIae79ef8_167, \10567 );
not \U$10192 ( \10569 , RIae79ef8_167);
buf \U$10193 ( \10570 , \10566 );
and \U$10194 ( \10571 , \10569 , \10570 );
nor \U$10195 ( \10572 , \10568 , \10571 );
not \U$10196 ( \10573 , \6213 );
nand \U$10197 ( \10574 , \10572 , \10573 );
nand \U$10198 ( \10575 , \10561 , \10574 );
and \U$10199 ( \10576 , \10558 , \10575 );
and \U$10200 ( \10577 , \10541 , \10557 );
or \U$10201 ( \10578 , \10576 , \10577 );
not \U$10202 ( \10579 , \2767 );
not \U$10203 ( \10580 , RIae79c28_161);
not \U$10204 ( \10581 , \1788 );
or \U$10205 ( \10582 , \10580 , \10581 );
not \U$10206 ( \10583 , \1788 );
not \U$10207 ( \10584 , RIae79c28_161);
nand \U$10208 ( \10585 , \10583 , \10584 );
nand \U$10209 ( \10586 , \10582 , \10585 );
not \U$10210 ( \10587 , \10586 );
or \U$10211 ( \10588 , \10579 , \10587 );
not \U$10212 ( \10589 , RIae79c28_161);
not \U$10213 ( \10590 , \2696 );
or \U$10214 ( \10591 , \10589 , \10590 );
or \U$10215 ( \10592 , \2696 , RIae79c28_161);
nand \U$10216 ( \10593 , \10591 , \10592 );
nand \U$10217 ( \10594 , \10593 , \2418 );
nand \U$10218 ( \10595 , \10588 , \10594 );
not \U$10219 ( \10596 , \10595 );
not \U$10220 ( \10597 , \10596 );
not \U$10221 ( \10598 , \4853 );
and \U$10222 ( \10599 , RIae79ca0_162, \3094 );
not \U$10223 ( \10600 , RIae79ca0_162);
and \U$10224 ( \10601 , \10600 , \3098 );
nor \U$10225 ( \10602 , \10599 , \10601 );
not \U$10226 ( \10603 , \10602 );
or \U$10227 ( \10604 , \10598 , \10603 );
buf \U$10228 ( \10605 , \4582 );
and \U$10229 ( \10606 , RIae79ca0_162, \10605 );
not \U$10230 ( \10607 , RIae79ca0_162);
not \U$10231 ( \10608 , \1753 );
and \U$10232 ( \10609 , \10607 , \10608 );
nor \U$10233 ( \10610 , \10606 , \10609 );
nand \U$10234 ( \10611 , \10610 , \4154 );
nand \U$10235 ( \10612 , \10604 , \10611 );
not \U$10236 ( \10613 , \10612 );
not \U$10237 ( \10614 , \10613 );
or \U$10238 ( \10615 , \10597 , \10614 );
not \U$10239 ( \10616 , \10595 );
not \U$10240 ( \10617 , \10612 );
or \U$10241 ( \10618 , \10616 , \10617 );
not \U$10242 ( \10619 , RIae7a510_180);
not \U$10243 ( \10620 , \2918 );
or \U$10244 ( \10621 , \10619 , \10620 );
or \U$10245 ( \10622 , \1472 , RIae7a510_180);
nand \U$10246 ( \10623 , \10621 , \10622 );
not \U$10247 ( \10624 , RIae7a588_181);
not \U$10248 ( \10625 , RIae7a498_179);
not \U$10249 ( \10626 , \10625 );
or \U$10250 ( \10627 , \10624 , \10626 );
not \U$10251 ( \10628 , RIae7a588_181);
nand \U$10252 ( \10629 , \10628 , RIae7a498_179);
nand \U$10253 ( \10630 , \10627 , \10629 );
buf \U$10254 ( \10631 , \10630 );
and \U$10255 ( \10632 , \10623 , \10631 );
not \U$10256 ( \10633 , RIae7a510_180);
or \U$10257 ( \10634 , \10633 , \10628 );
or \U$10258 ( \10635 , RIae7a498_179, RIae7a510_180);
nand \U$10259 ( \10636 , \10634 , \10635 , \10629 );
not \U$10260 ( \10637 , \10636 );
buf \U$10261 ( \10638 , \10637 );
not \U$10262 ( \10639 , \10638 );
not \U$10263 ( \10640 , \968 );
not \U$10264 ( \10641 , \970 );
and \U$10265 ( \10642 , \10640 , \10641 );
and \U$10266 ( \10643 , \968 , \970 );
nor \U$10267 ( \10644 , \10642 , \10643 );
not \U$10268 ( \10645 , \10644 );
not \U$10269 ( \10646 , RIae7a510_180);
and \U$10270 ( \10647 , \10645 , \10646 );
not \U$10271 ( \10648 , \10645 );
and \U$10272 ( \10649 , \10648 , RIae7a510_180);
nor \U$10273 ( \10650 , \10647 , \10649 );
nor \U$10274 ( \10651 , \10639 , \10650 );
nor \U$10275 ( \10652 , \10632 , \10651 );
nand \U$10276 ( \10653 , \10618 , \10652 );
nand \U$10277 ( \10654 , \10615 , \10653 );
not \U$10278 ( \10655 , \10654 );
or \U$10279 ( \10656 , \10578 , \10655 );
not \U$10280 ( \10657 , \9776 );
not \U$10281 ( \10658 , RIae7a150_172);
not \U$10282 ( \10659 , \10658 );
not \U$10283 ( \10660 , \917 );
or \U$10284 ( \10661 , \10659 , \10660 );
not \U$10285 ( \10662 , \917 );
nand \U$10286 ( \10663 , \10662 , RIae7a150_172);
nand \U$10287 ( \10664 , \10661 , \10663 );
not \U$10288 ( \10665 , \10664 );
or \U$10289 ( \10666 , \10657 , \10665 );
buf \U$10290 ( \10667 , \9757 );
nand \U$10291 ( \10668 , \9772 , \10667 );
nand \U$10292 ( \10669 , \10666 , \10668 );
not \U$10293 ( \10670 , RIae7a420_178);
and \U$10294 ( \10671 , \10670 , RIae7a150_172);
not \U$10295 ( \10672 , RIae7a150_172);
and \U$10296 ( \10673 , \10672 , RIae7a420_178);
nor \U$10297 ( \10674 , \10671 , \10673 );
not \U$10298 ( \10675 , \10674 );
buf \U$10299 ( \10676 , \10675 );
buf \U$10300 ( \10677 , \10676 );
not \U$10301 ( \10678 , \10677 );
and \U$10302 ( \10679 , RIae7a498_179, \854 );
not \U$10303 ( \10680 , RIae7a498_179);
and \U$10304 ( \10681 , \10680 , \855 );
nor \U$10305 ( \10682 , \10679 , \10681 );
not \U$10306 ( \10683 , \10682 );
or \U$10307 ( \10684 , \10678 , \10683 );
not \U$10308 ( \10685 , \10625 );
not \U$10309 ( \10686 , \883 );
or \U$10310 ( \10687 , \10685 , \10686 );
not \U$10311 ( \10688 , \2175 );
or \U$10312 ( \10689 , \10688 , \10625 );
nand \U$10313 ( \10690 , \10687 , \10689 );
and \U$10314 ( \10691 , RIae7a498_179, RIae7a420_178);
not \U$10315 ( \10692 , RIae7a498_179);
and \U$10316 ( \10693 , \10692 , \10670 );
nor \U$10317 ( \10694 , \10691 , \10693 );
and \U$10318 ( \10695 , \10674 , \10694 );
buf \U$10319 ( \10696 , \10695 );
nand \U$10320 ( \10697 , \10690 , \10696 );
nand \U$10321 ( \10698 , \10684 , \10697 );
xor \U$10322 ( \10699 , \10669 , \10698 );
buf \U$10323 ( \10700 , \9517 );
not \U$10324 ( \10701 , \10700 );
not \U$10325 ( \10702 , RIae79fe8_169);
not \U$10326 ( \10703 , \2629 );
or \U$10327 ( \10704 , \10702 , \10703 );
or \U$10328 ( \10705 , \4064 , RIae79fe8_169);
nand \U$10329 ( \10706 , \10704 , \10705 );
not \U$10330 ( \10707 , \10706 );
or \U$10331 ( \10708 , \10701 , \10707 );
buf \U$10332 ( \10709 , \9499 );
nand \U$10333 ( \10710 , \9515 , \10709 );
nand \U$10334 ( \10711 , \10708 , \10710 );
and \U$10335 ( \10712 , \10699 , \10711 );
and \U$10336 ( \10713 , \10669 , \10698 );
or \U$10337 ( \10714 , \10712 , \10713 );
nand \U$10338 ( \10715 , \10656 , \10714 );
nand \U$10339 ( \10716 , \10578 , \10655 );
nand \U$10340 ( \10717 , \10715 , \10716 );
buf \U$10341 ( \10718 , \10717 );
xor \U$10342 ( \10719 , \10529 , \10718 );
xnor \U$10343 ( \10720 , \10315 , \10719 );
not \U$10344 ( \10721 , \10720 );
not \U$10345 ( \10722 , \1008 );
not \U$10346 ( \10723 , RIae79160_138);
buf \U$10347 ( \10724 , \9923 );
buf \U$10348 ( \10725 , \10724 );
not \U$10349 ( \10726 , \10725 );
or \U$10350 ( \10727 , \10723 , \10726 );
not \U$10351 ( \10728 , \10724 );
not \U$10352 ( \10729 , \10728 );
or \U$10353 ( \10730 , \10729 , RIae79160_138);
nand \U$10354 ( \10731 , \10727 , \10730 );
not \U$10355 ( \10732 , \10731 );
or \U$10356 ( \10733 , \10722 , \10732 );
nand \U$10357 ( \10734 , \10467 , \1012 );
nand \U$10358 ( \10735 , \10733 , \10734 );
not \U$10359 ( \10736 , \10735 );
not \U$10360 ( \10737 , \1320 );
not \U$10361 ( \10738 , \10160 );
or \U$10362 ( \10739 , \10737 , \10738 );
buf \U$10363 ( \10740 , \9988 );
and \U$10364 ( \10741 , RIae78e90_132, \10740 );
not \U$10365 ( \10742 , RIae78e90_132);
not \U$10366 ( \10743 , \10740 );
and \U$10367 ( \10744 , \10742 , \10743 );
or \U$10368 ( \10745 , \10741 , \10744 );
nand \U$10369 ( \10746 , \10745 , \1086 );
nand \U$10370 ( \10747 , \10739 , \10746 );
not \U$10371 ( \10748 , \796 );
buf \U$10372 ( \10749 , \9874 );
buf \U$10373 ( \10750 , \10749 );
and \U$10374 ( \10751 , RIae78f80_134, \10750 );
not \U$10375 ( \10752 , RIae78f80_134);
and \U$10376 ( \10753 , \10752 , \9868 );
or \U$10377 ( \10754 , \10751 , \10753 );
not \U$10378 ( \10755 , \10754 );
or \U$10379 ( \10756 , \10748 , \10755 );
nand \U$10380 ( \10757 , \10173 , \838 );
nand \U$10381 ( \10758 , \10756 , \10757 );
xor \U$10382 ( \10759 , \10747 , \10758 );
not \U$10383 ( \10760 , \10759 );
or \U$10384 ( \10761 , \10736 , \10760 );
nand \U$10385 ( \10762 , \10758 , \10747 );
nand \U$10386 ( \10763 , \10761 , \10762 );
not \U$10387 ( \10764 , \2272 );
not \U$10388 ( \10765 , RIae79ac0_158);
not \U$10389 ( \10766 , \9299 );
or \U$10390 ( \10767 , \10765 , \10766 );
or \U$10391 ( \10768 , \9299 , RIae79ac0_158);
nand \U$10392 ( \10769 , \10767 , \10768 );
not \U$10393 ( \10770 , \10769 );
or \U$10394 ( \10771 , \10764 , \10770 );
nand \U$10395 ( \10772 , \9293 , \10414 );
nand \U$10396 ( \10773 , \10771 , \10772 );
not \U$10397 ( \10774 , \10773 );
not \U$10398 ( \10775 , \10401 );
not \U$10399 ( \10776 , \2970 );
not \U$10400 ( \10777 , \9347 );
not \U$10401 ( \10778 , \10777 );
or \U$10402 ( \10779 , \10776 , \10778 );
not \U$10403 ( \10780 , \9347 );
not \U$10404 ( \10781 , RIae79688_149);
or \U$10405 ( \10782 , \10780 , \10781 );
nand \U$10406 ( \10783 , \10779 , \10782 );
not \U$10407 ( \10784 , \10783 );
or \U$10408 ( \10785 , \10775 , \10784 );
nand \U$10409 ( \10786 , \9319 , \1820 );
nand \U$10410 ( \10787 , \10785 , \10786 );
not \U$10411 ( \10788 , \10787 );
or \U$10412 ( \10789 , \10774 , \10788 );
not \U$10413 ( \10790 , \10223 );
not \U$10414 ( \10791 , \10239 );
or \U$10415 ( \10792 , \10790 , \10791 );
not \U$10416 ( \10793 , \5722 );
and \U$10417 ( \10794 , RIae79520_146, \10793 );
not \U$10418 ( \10795 , RIae79520_146);
and \U$10419 ( \10796 , \10795 , \5722 );
or \U$10420 ( \10797 , \10794 , \10796 );
nand \U$10421 ( \10798 , \10797 , \5950 );
nand \U$10422 ( \10799 , \10792 , \10798 );
not \U$10423 ( \10800 , \10799 );
nand \U$10424 ( \10801 , \10789 , \10800 );
not \U$10425 ( \10802 , \10773 );
not \U$10426 ( \10803 , \10787 );
nand \U$10427 ( \10804 , \10802 , \10803 );
and \U$10428 ( \10805 , \10801 , \10804 );
xor \U$10429 ( \10806 , \10763 , \10805 );
buf \U$10430 ( \10807 , \2339 );
not \U$10431 ( \10808 , \10807 );
not \U$10432 ( \10809 , \4982 );
and \U$10433 ( \10810 , RIae798e0_154, \10809 );
not \U$10434 ( \10811 , RIae798e0_154);
not \U$10435 ( \10812 , \9830 );
and \U$10436 ( \10813 , \10811 , \10812 );
or \U$10437 ( \10814 , \10810 , \10813 );
not \U$10438 ( \10815 , \10814 );
or \U$10439 ( \10816 , \10808 , \10815 );
nand \U$10440 ( \10817 , \2322 , \10496 );
nand \U$10441 ( \10818 , \10816 , \10817 );
not \U$10442 ( \10819 , \10818 );
not \U$10443 ( \10820 , \1919 );
not \U$10444 ( \10821 , \10300 );
or \U$10445 ( \10822 , \10820 , \10821 );
not \U$10446 ( \10823 , RIae794a8_145);
not \U$10447 ( \10824 , \4953 );
not \U$10448 ( \10825 , \4955 );
and \U$10449 ( \10826 , \10824 , \10825 );
and \U$10450 ( \10827 , \4953 , \4955 );
nor \U$10451 ( \10828 , \10826 , \10827 );
buf \U$10452 ( \10829 , \10828 );
not \U$10453 ( \10830 , \10829 );
or \U$10454 ( \10831 , \10823 , \10830 );
or \U$10455 ( \10832 , \10226 , RIae794a8_145);
nand \U$10456 ( \10833 , \10831 , \10832 );
nand \U$10457 ( \10834 , \10833 , \1933 );
nand \U$10458 ( \10835 , \10822 , \10834 );
or \U$10459 ( \10836 , \10243 , \10242 );
nand \U$10460 ( \10837 , \10836 , \10245 );
not \U$10461 ( \10838 , \10837 );
nand \U$10462 ( \10839 , \10248 , \10251 );
not \U$10463 ( \10840 , \10839 );
and \U$10464 ( \10841 , \10838 , \10840 );
and \U$10465 ( \10842 , \10837 , \10839 );
nor \U$10466 ( \10843 , \10841 , \10842 );
buf \U$10467 ( \10844 , \10843 );
not \U$10468 ( \10845 , \10844 );
and \U$10469 ( \10846 , RIae78b48_125, \10845 );
not \U$10470 ( \10847 , \10846 );
nand \U$10471 ( \10848 , \10847 , RIae7aa38_191);
and \U$10472 ( \10849 , \10848 , \10260 );
not \U$10473 ( \10850 , \10848 );
not \U$10474 ( \10851 , \10260 );
and \U$10475 ( \10852 , \10850 , \10851 );
nor \U$10476 ( \10853 , \10849 , \10852 );
not \U$10477 ( \10854 , \10853 );
not \U$10478 ( \10855 , \926 );
buf \U$10479 ( \10856 , \10031 );
not \U$10480 ( \10857 , \10856 );
and \U$10481 ( \10858 , RIae78bc0_126, \10857 );
not \U$10482 ( \10859 , RIae78bc0_126);
and \U$10483 ( \10860 , \10859 , \10856 );
or \U$10484 ( \10861 , \10858 , \10860 );
not \U$10485 ( \10862 , \10861 );
or \U$10486 ( \10863 , \10855 , \10862 );
not \U$10487 ( \10864 , \10042 );
not \U$10488 ( \10865 , \1286 );
or \U$10489 ( \10866 , \10864 , \10865 );
or \U$10490 ( \10867 , \10047 , \1286 );
nand \U$10491 ( \10868 , \10866 , \10867 );
nand \U$10492 ( \10869 , \10868 , \951 );
nand \U$10493 ( \10870 , \10863 , \10869 );
not \U$10494 ( \10871 , \10870 );
or \U$10495 ( \10872 , \10854 , \10871 );
nand \U$10496 ( \10873 , \10260 , \10848 );
nand \U$10497 ( \10874 , \10872 , \10873 );
xor \U$10498 ( \10875 , \10835 , \10874 );
not \U$10499 ( \10876 , \10875 );
or \U$10500 ( \10877 , \10819 , \10876 );
nand \U$10501 ( \10878 , \10835 , \10874 );
nand \U$10502 ( \10879 , \10877 , \10878 );
xor \U$10503 ( \10880 , \10806 , \10879 );
not \U$10504 ( \10881 , \10880 );
not \U$10505 ( \10882 , \4853 );
not \U$10506 ( \10883 , \1808 );
not \U$10507 ( \10884 , \10883 );
xor \U$10508 ( \10885 , \10884 , RIae79ca0_162);
not \U$10509 ( \10886 , \10885 );
or \U$10510 ( \10887 , \10882 , \10886 );
not \U$10511 ( \10888 , RIae79ca0_162);
not \U$10512 ( \10889 , \2577 );
or \U$10513 ( \10890 , \10888 , \10889 );
not \U$10514 ( \10891 , \1788 );
not \U$10515 ( \10892 , RIae79ca0_162);
nand \U$10516 ( \10893 , \10891 , \10892 );
nand \U$10517 ( \10894 , \10890 , \10893 );
nand \U$10518 ( \10895 , \10894 , \6276 );
nand \U$10519 ( \10896 , \10887 , \10895 );
not \U$10520 ( \10897 , \5049 );
and \U$10521 ( \10898 , \1740 , RIae79d90_164);
not \U$10522 ( \10899 , \1740 );
not \U$10523 ( \10900 , RIae79d90_164);
and \U$10524 ( \10901 , \10899 , \10900 );
nor \U$10525 ( \10902 , \10898 , \10901 );
not \U$10526 ( \10903 , \10902 );
or \U$10527 ( \10904 , \10897 , \10903 );
not \U$10528 ( \10905 , \4582 );
and \U$10529 ( \10906 , RIae79d90_164, \10905 );
not \U$10530 ( \10907 , RIae79d90_164);
not \U$10531 ( \10908 , \10905 );
and \U$10532 ( \10909 , \10907 , \10908 );
or \U$10533 ( \10910 , \10906 , \10909 );
nand \U$10534 ( \10911 , \10910 , \6091 );
nand \U$10535 ( \10912 , \10904 , \10911 );
or \U$10536 ( \10913 , \10896 , \10912 );
not \U$10537 ( \10914 , \10913 );
not \U$10538 ( \10915 , \10631 );
not \U$10539 ( \10916 , \1186 );
and \U$10540 ( \10917 , RIae7a510_180, \10916 );
not \U$10541 ( \10918 , RIae7a510_180);
and \U$10542 ( \10919 , \10918 , \1186 );
nor \U$10543 ( \10920 , \10917 , \10919 );
not \U$10544 ( \10921 , \10920 );
or \U$10545 ( \10922 , \10915 , \10921 );
and \U$10546 ( \10923 , RIae7a510_180, \1834 );
not \U$10547 ( \10924 , RIae7a510_180);
and \U$10548 ( \10925 , \10924 , \2850 );
or \U$10549 ( \10926 , \10923 , \10925 );
buf \U$10550 ( \10927 , \10637 );
nand \U$10551 ( \10928 , \10926 , \10927 );
nand \U$10552 ( \10929 , \10922 , \10928 );
not \U$10553 ( \10930 , \10929 );
or \U$10554 ( \10931 , \10914 , \10930 );
nand \U$10555 ( \10932 , \10896 , \10912 );
nand \U$10556 ( \10933 , \10931 , \10932 );
not \U$10557 ( \10934 , \10933 );
not \U$10558 ( \10935 , \1910 );
buf \U$10559 ( \10936 , \9394 );
not \U$10560 ( \10937 , \10936 );
not \U$10561 ( \10938 , \10937 );
xor \U$10562 ( \10939 , \10938 , RIae793b8_143);
not \U$10563 ( \10940 , \10939 );
or \U$10564 ( \10941 , \10935 , \10940 );
nand \U$10565 ( \10942 , \9461 , \1864 );
nand \U$10566 ( \10943 , \10941 , \10942 );
not \U$10567 ( \10944 , \10943 );
not \U$10568 ( \10945 , \10944 );
and \U$10569 ( \10946 , \10285 , \10851 );
not \U$10570 ( \10947 , \10285 );
and \U$10571 ( \10948 , \10947 , \10260 );
or \U$10572 ( \10949 , \10946 , \10948 );
not \U$10573 ( \10950 , \10949 );
not \U$10574 ( \10951 , \2011 );
not \U$10575 ( \10952 , \9369 );
or \U$10576 ( \10953 , \10951 , \10952 );
not \U$10577 ( \10954 , \2056 );
not \U$10578 ( \10955 , \9441 );
or \U$10579 ( \10956 , \10954 , \10955 );
not \U$10580 ( \10957 , RIae79610_148);
or \U$10581 ( \10958 , \9441 , \10957 );
nand \U$10582 ( \10959 , \10956 , \10958 );
nand \U$10583 ( \10960 , \10959 , \2063 );
nand \U$10584 ( \10961 , \10953 , \10960 );
not \U$10585 ( \10962 , \10961 );
not \U$10586 ( \10963 , \10962 );
or \U$10587 ( \10964 , \10950 , \10963 );
or \U$10588 ( \10965 , \10962 , \10949 );
nand \U$10589 ( \10966 , \10964 , \10965 );
not \U$10590 ( \10967 , \10966 );
or \U$10591 ( \10968 , \10945 , \10967 );
or \U$10592 ( \10969 , \10944 , \10966 );
nand \U$10593 ( \10970 , \10968 , \10969 );
not \U$10594 ( \10971 , \10970 );
not \U$10595 ( \10972 , \10773 );
not \U$10596 ( \10973 , \10803 );
or \U$10597 ( \10974 , \10972 , \10973 );
or \U$10598 ( \10975 , \10803 , \10773 );
nand \U$10599 ( \10976 , \10974 , \10975 );
not \U$10600 ( \10977 , \10976 );
not \U$10601 ( \10978 , \10800 );
and \U$10602 ( \10979 , \10977 , \10978 );
and \U$10603 ( \10980 , \10976 , \10800 );
nor \U$10604 ( \10981 , \10979 , \10980 );
not \U$10605 ( \10982 , \10981 );
or \U$10606 ( \10983 , \10971 , \10982 );
or \U$10607 ( \10984 , \10970 , \10981 );
nand \U$10608 ( \10985 , \10983 , \10984 );
not \U$10609 ( \10986 , \10985 );
or \U$10610 ( \10987 , \10934 , \10986 );
not \U$10611 ( \10988 , \10981 );
nand \U$10612 ( \10989 , \10988 , \10970 );
nand \U$10613 ( \10990 , \10987 , \10989 );
not \U$10614 ( \10991 , \10990 );
xnor \U$10615 ( \10992 , \10214 , \10201 );
xor \U$10616 ( \10993 , \10153 , \10175 );
xnor \U$10617 ( \10994 , \10993 , \10162 );
not \U$10618 ( \10995 , \10994 );
xor \U$10619 ( \10996 , \10992 , \10995 );
not \U$10620 ( \10997 , \10943 );
not \U$10621 ( \10998 , \10966 );
or \U$10622 ( \10999 , \10997 , \10998 );
not \U$10623 ( \11000 , \10962 );
nand \U$10624 ( \11001 , \11000 , \10949 );
nand \U$10625 ( \11002 , \10999 , \11001 );
buf \U$10626 ( \11003 , \11002 );
xor \U$10627 ( \11004 , \10996 , \11003 );
nand \U$10628 ( \11005 , \10991 , \11004 );
not \U$10629 ( \11006 , \11005 );
or \U$10630 ( \11007 , \10881 , \11006 );
not \U$10631 ( \11008 , \11004 );
nand \U$10632 ( \11009 , \11008 , \10990 );
nand \U$10633 ( \11010 , \11007 , \11009 );
not \U$10634 ( \11011 , \11010 );
not \U$10635 ( \11012 , \11011 );
buf \U$10636 ( \11013 , \9643 );
buf \U$10637 ( \11014 , \11013 );
not \U$10638 ( \11015 , \11014 );
and \U$10639 ( \11016 , RIae7a3a8_177, \2593 );
not \U$10640 ( \11017 , RIae7a3a8_177);
and \U$10641 ( \11018 , \11017 , \3146 );
or \U$10642 ( \11019 , \11016 , \11018 );
not \U$10643 ( \11020 , \11019 );
or \U$10644 ( \11021 , \11015 , \11020 );
nand \U$10645 ( \11022 , \9636 , \9622 );
nand \U$10646 ( \11023 , \11021 , \11022 );
not \U$10647 ( \11024 , \2007 );
not \U$10648 ( \11025 , \9661 );
or \U$10649 ( \11026 , \11024 , \11025 );
and \U$10650 ( \11027 , \2403 , \1997 );
not \U$10651 ( \11028 , \2403 );
and \U$10652 ( \11029 , \11028 , RIae797f0_152);
nor \U$10653 ( \11030 , \11027 , \11029 );
nand \U$10654 ( \11031 , \11030 , \1988 );
nand \U$10655 ( \11032 , \11026 , \11031 );
or \U$10656 ( \11033 , \11023 , \11032 );
not \U$10657 ( \11034 , \11032 );
not \U$10658 ( \11035 , \11023 );
or \U$10659 ( \11036 , \11034 , \11035 );
buf \U$10660 ( \11037 , \2450 );
not \U$10661 ( \11038 , \11037 );
not \U$10662 ( \11039 , \9582 );
or \U$10663 ( \11040 , \11038 , \11039 );
not \U$10664 ( \11041 , RIae79778_151);
not \U$10665 ( \11042 , \3216 );
or \U$10666 ( \11043 , \11041 , \11042 );
or \U$10667 ( \11044 , \1969 , RIae79778_151);
nand \U$10668 ( \11045 , \11043 , \11044 );
nand \U$10669 ( \11046 , \11045 , \2545 );
nand \U$10670 ( \11047 , \11040 , \11046 );
not \U$10671 ( \11048 , \11047 );
nand \U$10672 ( \11049 , \11036 , \11048 );
and \U$10673 ( \11050 , \11033 , \11049 );
not \U$10674 ( \11051 , \11050 );
not \U$10675 ( \11052 , \11051 );
not \U$10676 ( \11053 , \9792 );
not \U$10677 ( \11054 , RIae7a2b8_175);
not \U$10678 ( \11055 , \11054 );
not \U$10679 ( \11056 , \2230 );
not \U$10680 ( \11057 , \11056 );
or \U$10681 ( \11058 , \11055 , \11057 );
nand \U$10682 ( \11059 , \2993 , RIae7a2b8_175);
nand \U$10683 ( \11060 , \11058 , \11059 );
not \U$10684 ( \11061 , \11060 );
or \U$10685 ( \11062 , \11053 , \11061 );
nand \U$10686 ( \11063 , \9801 , \9815 );
nand \U$10687 ( \11064 , \11062 , \11063 );
not \U$10688 ( \11065 , \11064 );
not \U$10689 ( \11066 , \10700 );
not \U$10690 ( \11067 , \9506 );
or \U$10691 ( \11068 , \11066 , \11067 );
not \U$10692 ( \11069 , RIae79fe8_169);
not \U$10693 ( \11070 , \11069 );
not \U$10694 ( \11071 , \2153 );
not \U$10695 ( \11072 , \11071 );
or \U$10696 ( \11073 , \11070 , \11072 );
nand \U$10697 ( \11074 , \2153 , RIae79fe8_169);
nand \U$10698 ( \11075 , \11073 , \11074 );
nand \U$10699 ( \11076 , \11075 , \10709 );
nand \U$10700 ( \11077 , \11068 , \11076 );
not \U$10701 ( \11078 , \11077 );
or \U$10702 ( \11079 , \11065 , \11078 );
not \U$10703 ( \11080 , \9777 );
not \U$10704 ( \11081 , \9765 );
or \U$10705 ( \11082 , \11080 , \11081 );
and \U$10706 ( \11083 , RIae7a150_172, \2175 );
not \U$10707 ( \11084 , RIae7a150_172);
and \U$10708 ( \11085 , \11084 , \10688 );
or \U$10709 ( \11086 , \11083 , \11085 );
buf \U$10710 ( \11087 , \9758 );
nand \U$10711 ( \11088 , \11086 , \11087 );
nand \U$10712 ( \11089 , \11082 , \11088 );
not \U$10713 ( \11090 , \11089 );
nand \U$10714 ( \11091 , \11079 , \11090 );
not \U$10715 ( \11092 , \11064 );
not \U$10716 ( \11093 , \11077 );
nand \U$10717 ( \11094 , \11092 , \11093 );
nand \U$10718 ( \11095 , \11091 , \11094 );
not \U$10719 ( \11096 , \11095 );
or \U$10720 ( \11097 , \11052 , \11096 );
buf \U$10721 ( \11098 , \10542 );
not \U$10722 ( \11099 , \11098 );
not \U$10723 ( \11100 , \9736 );
or \U$10724 ( \11101 , \11099 , \11100 );
not \U$10725 ( \11102 , RIae7a060_170);
not \U$10726 ( \11103 , \11102 );
not \U$10727 ( \11104 , \939 );
or \U$10728 ( \11105 , \11103 , \11104 );
or \U$10729 ( \11106 , \939 , \11102 );
nand \U$10730 ( \11107 , \11105 , \11106 );
nand \U$10731 ( \11108 , \11107 , \9730 );
nand \U$10732 ( \11109 , \11101 , \11108 );
not \U$10733 ( \11110 , \11109 );
not \U$10734 ( \11111 , \9699 );
not \U$10735 ( \11112 , \9690 );
or \U$10736 ( \11113 , \11111 , \11112 );
not \U$10737 ( \11114 , RIae7a240_174);
not \U$10738 ( \11115 , \11114 );
not \U$10739 ( \11116 , \3294 );
or \U$10740 ( \11117 , \11115 , \11116 );
or \U$10741 ( \11118 , \9807 , \11114 );
nand \U$10742 ( \11119 , \11117 , \11118 );
nand \U$10743 ( \11120 , \11119 , \9687 );
nand \U$10744 ( \11121 , \11113 , \11120 );
not \U$10745 ( \11122 , \9473 );
and \U$10746 ( \11123 , RIae7a6f0_184, \781 );
not \U$10747 ( \11124 , RIae7a6f0_184);
and \U$10748 ( \11125 , \11124 , \1993 );
nor \U$10749 ( \11126 , \11123 , \11125 );
not \U$10750 ( \11127 , \11126 );
or \U$10751 ( \11128 , \11122 , \11127 );
nand \U$10752 ( \11129 , \9713 , \9705 );
nand \U$10753 ( \11130 , \11128 , \11129 );
and \U$10754 ( \11131 , \11121 , \11130 );
not \U$10755 ( \11132 , \11121 );
not \U$10756 ( \11133 , \11130 );
and \U$10757 ( \11134 , \11132 , \11133 );
nor \U$10758 ( \11135 , \11131 , \11134 );
not \U$10759 ( \11136 , \11135 );
or \U$10760 ( \11137 , \11110 , \11136 );
nand \U$10761 ( \11138 , \11130 , \11121 );
nand \U$10762 ( \11139 , \11137 , \11138 );
nand \U$10763 ( \11140 , \11097 , \11139 );
nand \U$10764 ( \11141 , \11050 , \11094 , \11091 );
nand \U$10765 ( \11142 , \11140 , \11141 );
not \U$10766 ( \11143 , \11142 );
not \U$10767 ( \11144 , \2011 );
not \U$10768 ( \11145 , \10959 );
or \U$10769 ( \11146 , \11144 , \11145 );
not \U$10770 ( \11147 , \2056 );
not \U$10771 ( \11148 , \9455 );
or \U$10772 ( \11149 , \11147 , \11148 );
not \U$10773 ( \11150 , RIae79610_148);
or \U$10774 ( \11151 , \9459 , \11150 );
nand \U$10775 ( \11152 , \11149 , \11151 );
nand \U$10776 ( \11153 , \11152 , \2063 );
nand \U$10777 ( \11154 , \11146 , \11153 );
not \U$10778 ( \11155 , \1820 );
not \U$10779 ( \11156 , \10783 );
or \U$10780 ( \11157 , \11155 , \11156 );
xor \U$10781 ( \11158 , RIae79688_149, \9363 );
nand \U$10782 ( \11159 , \11158 , \1843 );
nand \U$10783 ( \11160 , \11157 , \11159 );
and \U$10784 ( \11161 , \11154 , \11160 );
not \U$10785 ( \11162 , \11154 );
not \U$10786 ( \11163 , \11160 );
and \U$10787 ( \11164 , \11162 , \11163 );
nor \U$10788 ( \11165 , \11161 , \11164 );
not \U$10789 ( \11166 , \2251 );
not \U$10790 ( \11167 , \10769 );
or \U$10791 ( \11168 , \11166 , \11167 );
and \U$10792 ( \11169 , \9313 , \2268 );
not \U$10793 ( \11170 , \9313 );
and \U$10794 ( \11171 , \11170 , RIae79ac0_158);
nor \U$10795 ( \11172 , \11169 , \11171 );
nand \U$10796 ( \11173 , \2272 , \11172 );
nand \U$10797 ( \11174 , \11168 , \11173 );
nand \U$10798 ( \11175 , \11165 , \11174 );
nand \U$10799 ( \11176 , \11160 , \11154 );
nand \U$10800 ( \11177 , \11175 , \11176 );
xor \U$10801 ( \11178 , \10735 , \10759 );
xor \U$10802 ( \11179 , \11177 , \11178 );
not \U$10803 ( \11180 , \11179 );
not \U$10804 ( \11181 , \1501 );
not \U$10805 ( \11182 , \9613 );
or \U$10806 ( \11183 , \11181 , \11182 );
and \U$10807 ( \11184 , RIae79250_140, \10465 );
not \U$10808 ( \11185 , RIae79250_140);
buf \U$10809 ( \11186 , \9940 );
not \U$10810 ( \11187 , \11186 );
and \U$10811 ( \11188 , \11185 , \11187 );
nor \U$10812 ( \11189 , \11184 , \11188 );
nand \U$10813 ( \11190 , \11189 , \1499 );
nand \U$10814 ( \11191 , \11183 , \11190 );
not \U$10815 ( \11192 , \1863 );
not \U$10816 ( \11193 , \10939 );
or \U$10817 ( \11194 , \11192 , \11193 );
buf \U$10818 ( \11195 , \9412 );
and \U$10819 ( \11196 , RIae793b8_143, \11195 );
not \U$10820 ( \11197 , RIae793b8_143);
not \U$10821 ( \11198 , \9412 );
and \U$10822 ( \11199 , \11197 , \11198 );
or \U$10823 ( \11200 , \11196 , \11199 );
nand \U$10824 ( \11201 , \1910 , \11200 );
nand \U$10825 ( \11202 , \11194 , \11201 );
xor \U$10826 ( \11203 , \11191 , \11202 );
buf \U$10827 ( \11204 , \10280 );
buf \U$10828 ( \11205 , \11204 );
not \U$10829 ( \11206 , \11205 );
not \U$10830 ( \11207 , RIae7a8d0_188);
not \U$10831 ( \11208 , \11207 );
not \U$10832 ( \11209 , \991 );
or \U$10833 ( \11210 , \11208 , \11209 );
or \U$10834 ( \11211 , \2444 , \11207 );
nand \U$10835 ( \11212 , \11210 , \11211 );
not \U$10836 ( \11213 , \11212 );
or \U$10837 ( \11214 , \11206 , \11213 );
nand \U$10838 ( \11215 , \10275 , RIae7a8d0_188);
nand \U$10839 ( \11216 , \11214 , \11215 );
and \U$10840 ( \11217 , \11203 , \11216 );
and \U$10841 ( \11218 , \11191 , \11202 );
or \U$10842 ( \11219 , \11217 , \11218 );
not \U$10843 ( \11220 , \11219 );
or \U$10844 ( \11221 , \11180 , \11220 );
not \U$10845 ( \11222 , \11176 );
not \U$10846 ( \11223 , \11175 );
or \U$10847 ( \11224 , \11222 , \11223 );
nand \U$10848 ( \11225 , \11224 , \11178 );
nand \U$10849 ( \11226 , \11221 , \11225 );
not \U$10850 ( \11227 , \9947 );
not \U$10851 ( \11228 , \10212 );
or \U$10852 ( \11229 , \11227 , \11228 );
not \U$10853 ( \11230 , \10070 );
and \U$10854 ( \11231 , RIae79070_136, \11230 );
not \U$10855 ( \11232 , RIae79070_136);
and \U$10856 ( \11233 , \11232 , \10072 );
or \U$10857 ( \11234 , \11231 , \11233 );
nand \U$10858 ( \11235 , \11234 , \1062 );
nand \U$10859 ( \11236 , \11229 , \11235 );
not \U$10860 ( \11237 , \867 );
not \U$10861 ( \11238 , \10049 );
or \U$10862 ( \11239 , \11237 , \11238 );
not \U$10863 ( \11240 , \10193 );
and \U$10864 ( \11241 , RIae78b48_125, \11240 );
not \U$10865 ( \11242 , RIae78b48_125);
and \U$10866 ( \11243 , \11242 , \10195 );
or \U$10867 ( \11244 , \11241 , \11243 );
nand \U$10868 ( \11245 , \11244 , \1129 );
nand \U$10869 ( \11246 , \11239 , \11245 );
nand \U$10870 ( \11247 , \10861 , \951 );
nand \U$10871 ( \11248 , \10151 , \926 );
and \U$10872 ( \11249 , \11247 , \11248 );
and \U$10873 ( \11250 , \11246 , \11249 );
not \U$10874 ( \11251 , \11246 );
nand \U$10875 ( \11252 , \11248 , \11247 );
and \U$10876 ( \11253 , \11251 , \11252 );
or \U$10877 ( \11254 , \11250 , \11253 );
xor \U$10878 ( \11255 , \11236 , \11254 );
not \U$10879 ( \11256 , \838 );
not \U$10880 ( \11257 , \10754 );
or \U$10881 ( \11258 , \11256 , \11257 );
not \U$10882 ( \11259 , \9999 );
not \U$10883 ( \11260 , \11259 );
and \U$10884 ( \11261 , RIae78f80_134, \11260 );
not \U$10885 ( \11262 , RIae78f80_134);
and \U$10886 ( \11263 , \11262 , \10007 );
or \U$10887 ( \11264 , \11261 , \11263 );
nand \U$10888 ( \11265 , \11264 , \797 );
nand \U$10889 ( \11266 , \11258 , \11265 );
not \U$10890 ( \11267 , \1049 );
not \U$10891 ( \11268 , \11234 );
or \U$10892 ( \11269 , \11267 , \11268 );
and \U$10893 ( \11270 , RIae79070_136, \10168 );
not \U$10894 ( \11271 , RIae79070_136);
not \U$10895 ( \11272 , \9897 );
and \U$10896 ( \11273 , \11271 , \11272 );
or \U$10897 ( \11274 , \11270 , \11273 );
nand \U$10898 ( \11275 , \11274 , \1062 );
nand \U$10899 ( \11276 , \11269 , \11275 );
and \U$10900 ( \11277 , \11266 , \11276 );
not \U$10901 ( \11278 , \11266 );
not \U$10902 ( \11279 , \11276 );
and \U$10903 ( \11280 , \11278 , \11279 );
nor \U$10904 ( \11281 , \11277 , \11280 );
not \U$10905 ( \11282 , \11281 );
not \U$10906 ( \11283 , \1919 );
not \U$10907 ( \11284 , \10833 );
or \U$10908 ( \11285 , \11283 , \11284 );
not \U$10909 ( \11286 , RIae794a8_145);
not \U$10910 ( \11287 , \10237 );
or \U$10911 ( \11288 , \11286 , \11287 );
or \U$10912 ( \11289 , \10237 , RIae794a8_145);
nand \U$10913 ( \11290 , \11288 , \11289 );
nand \U$10914 ( \11291 , \11290 , \2457 );
nand \U$10915 ( \11292 , \11285 , \11291 );
not \U$10916 ( \11293 , \11292 );
or \U$10917 ( \11294 , \11282 , \11293 );
nand \U$10918 ( \11295 , \11276 , \11266 );
nand \U$10919 ( \11296 , \11294 , \11295 );
xor \U$10920 ( \11297 , \11255 , \11296 );
not \U$10921 ( \11298 , \2322 );
not \U$10922 ( \11299 , \10814 );
or \U$10923 ( \11300 , \11298 , \11299 );
and \U$10924 ( \11301 , RIae798e0_154, \6238 );
not \U$10925 ( \11302 , RIae798e0_154);
and \U$10926 ( \11303 , \11302 , \4169 );
or \U$10927 ( \11304 , \11301 , \11303 );
nand \U$10928 ( \11305 , \11304 , \10807 );
nand \U$10929 ( \11306 , \11300 , \11305 );
not \U$10930 ( \11307 , \11306 );
not \U$10931 ( \11308 , \892 );
not \U$10932 ( \11309 , \10259 );
and \U$10933 ( \11310 , RIae78b48_125, \11309 );
not \U$10934 ( \11311 , RIae78b48_125);
and \U$10935 ( \11312 , \11311 , \10259 );
nor \U$10936 ( \11313 , \11310 , \11312 );
not \U$10937 ( \11314 , \11313 );
or \U$10938 ( \11315 , \11308 , \11314 );
not \U$10939 ( \11316 , \860 );
buf \U$10940 ( \11317 , \10271 );
buf \U$10941 ( \11318 , \11317 );
not \U$10942 ( \11319 , \11318 );
or \U$10943 ( \11320 , \11316 , \11319 );
buf \U$10944 ( \11321 , \11317 );
or \U$10945 ( \11322 , \11321 , \860 );
nand \U$10946 ( \11323 , \11320 , \11322 );
nand \U$10947 ( \11324 , \11323 , \867 );
nand \U$10948 ( \11325 , \11315 , \11324 );
not \U$10949 ( \11326 , RIae7aa38_191);
not \U$10950 ( \11327 , \11326 );
not \U$10951 ( \11328 , \10846 );
or \U$10952 ( \11329 , \11327 , \11328 );
nand \U$10953 ( \11330 , \11329 , \10848 );
and \U$10954 ( \11331 , \11325 , \11330 );
not \U$10955 ( \11332 , \5950 );
and \U$10956 ( \11333 , RIae79520_146, \10409 );
not \U$10957 ( \11334 , RIae79520_146);
and \U$10958 ( \11335 , \11334 , \6345 );
or \U$10959 ( \11336 , \11333 , \11335 );
not \U$10960 ( \11337 , \11336 );
or \U$10961 ( \11338 , \11332 , \11337 );
nand \U$10962 ( \11339 , \10797 , \10223 );
nand \U$10963 ( \11340 , \11338 , \11339 );
xor \U$10964 ( \11341 , \11331 , \11340 );
not \U$10965 ( \11342 , \11341 );
or \U$10966 ( \11343 , \11307 , \11342 );
nand \U$10967 ( \11344 , \11340 , \11331 );
nand \U$10968 ( \11345 , \11343 , \11344 );
and \U$10969 ( \11346 , \11297 , \11345 );
and \U$10970 ( \11347 , \11255 , \11296 );
or \U$10971 ( \11348 , \11346 , \11347 );
or \U$10972 ( \11349 , \11226 , \11348 );
not \U$10973 ( \11350 , \11349 );
or \U$10974 ( \11351 , \11143 , \11350 );
nand \U$10975 ( \11352 , \11226 , \11348 );
nand \U$10976 ( \11353 , \11351 , \11352 );
not \U$10977 ( \11354 , \11353 );
not \U$10978 ( \11355 , \11354 );
or \U$10979 ( \11356 , \11012 , \11355 );
not \U$10980 ( \11357 , \2767 );
and \U$10981 ( \11358 , \6413 , RIae79c28_161);
not \U$10982 ( \11359 , \6413 );
and \U$10983 ( \11360 , \11359 , \10584 );
nor \U$10984 ( \11361 , \11358 , \11360 );
not \U$10985 ( \11362 , \11361 );
or \U$10986 ( \11363 , \11357 , \11362 );
not \U$10987 ( \11364 , \2410 );
nand \U$10988 ( \11365 , \10586 , \11364 );
nand \U$10989 ( \11366 , \11363 , \11365 );
not \U$10990 ( \11367 , \867 );
not \U$10991 ( \11368 , \11244 );
or \U$10992 ( \11369 , \11367 , \11368 );
nand \U$10993 ( \11370 , \11323 , \892 );
nand \U$10994 ( \11371 , \11369 , \11370 );
not \U$10995 ( \11372 , \1072 );
not \U$10996 ( \11373 , \10745 );
or \U$10997 ( \11374 , \11372 , \11373 );
and \U$10998 ( \11375 , RIae78e90_132, \10149 );
not \U$10999 ( \11376 , RIae78e90_132);
and \U$11000 ( \11377 , \11376 , \10142 );
or \U$11001 ( \11378 , \11375 , \11377 );
nand \U$11002 ( \11379 , \11378 , \1086 );
nand \U$11003 ( \11380 , \11374 , \11379 );
xor \U$11004 ( \11381 , \11371 , \11380 );
not \U$11005 ( \11382 , \11381 );
not \U$11006 ( \11383 , \1012 );
not \U$11007 ( \11384 , \10731 );
or \U$11008 ( \11385 , \11383 , \11384 );
not \U$11009 ( \11386 , \10083 );
not \U$11010 ( \11387 , \11386 );
and \U$11011 ( \11388 , RIae79160_138, \11387 );
not \U$11012 ( \11389 , RIae79160_138);
and \U$11013 ( \11390 , \11389 , \10208 );
or \U$11014 ( \11391 , \11388 , \11390 );
nand \U$11015 ( \11392 , \11391 , \1008 );
nand \U$11016 ( \11393 , \11385 , \11392 );
not \U$11017 ( \11394 , \11393 );
or \U$11018 ( \11395 , \11382 , \11394 );
nand \U$11019 ( \11396 , \11380 , \11371 );
nand \U$11020 ( \11397 , \11395 , \11396 );
not \U$11021 ( \11398 , \11397 );
xor \U$11022 ( \11399 , \11366 , \11398 );
not \U$11023 ( \11400 , \10636 );
not \U$11024 ( \11401 , \11400 );
not \U$11025 ( \11402 , \10920 );
or \U$11026 ( \11403 , \11401 , \11402 );
not \U$11027 ( \11404 , \10650 );
nand \U$11028 ( \11405 , \11404 , \10631 );
nand \U$11029 ( \11406 , \11403 , \11405 );
xnor \U$11030 ( \11407 , \11399 , \11406 );
not \U$11031 ( \11408 , \11407 );
buf \U$11032 ( \11409 , \6201 );
not \U$11033 ( \11410 , \11409 );
not \U$11034 ( \11411 , RIae79ef8_167);
not \U$11035 ( \11412 , \2287 );
or \U$11036 ( \11413 , \11411 , \11412 );
or \U$11037 ( \11414 , \2287 , RIae79ef8_167);
nand \U$11038 ( \11415 , \11413 , \11414 );
not \U$11039 ( \11416 , \11415 );
or \U$11040 ( \11417 , \11410 , \11416 );
nand \U$11041 ( \11418 , \9565 , \6214 );
nand \U$11042 ( \11419 , \11417 , \11418 );
not \U$11043 ( \11420 , \11419 );
not \U$11044 ( \11421 , \10675 );
not \U$11045 ( \11422 , \11421 );
not \U$11046 ( \11423 , \11422 );
xor \U$11047 ( \11424 , RIae7a498_179, \1118 );
not \U$11048 ( \11425 , \11424 );
or \U$11049 ( \11426 , \11423 , \11425 );
not \U$11050 ( \11427 , RIae7a498_179);
not \U$11051 ( \11428 , \11427 );
not \U$11052 ( \11429 , \10644 );
not \U$11053 ( \11430 , \11429 );
or \U$11054 ( \11431 , \11428 , \11430 );
or \U$11055 ( \11432 , \10645 , \10625 );
nand \U$11056 ( \11433 , \11431 , \11432 );
buf \U$11057 ( \11434 , \10695 );
nand \U$11058 ( \11435 , \11433 , \11434 );
nand \U$11059 ( \11436 , \11426 , \11435 );
not \U$11060 ( \11437 , \11436 );
and \U$11061 ( \11438 , \9543 , \9527 );
buf \U$11062 ( \11439 , \9549 );
not \U$11063 ( \11440 , \11439 );
not \U$11064 ( \11441 , \1157 );
not \U$11065 ( \11442 , \11441 );
not \U$11066 ( \11443 , RIae7a7e0_186);
and \U$11067 ( \11444 , \11442 , \11443 );
and \U$11068 ( \11445 , \1288 , RIae7a7e0_186);
nor \U$11069 ( \11446 , \11444 , \11445 );
nor \U$11070 ( \11447 , \11440 , \11446 );
nor \U$11071 ( \11448 , \11438 , \11447 );
not \U$11072 ( \11449 , \11448 );
or \U$11073 ( \11450 , \11437 , \11449 );
or \U$11074 ( \11451 , \11436 , \11448 );
nand \U$11075 ( \11452 , \11450 , \11451 );
not \U$11076 ( \11453 , \11452 );
or \U$11077 ( \11454 , \11420 , \11453 );
not \U$11078 ( \11455 , \11448 );
nand \U$11079 ( \11456 , \11455 , \11436 );
nand \U$11080 ( \11457 , \11454 , \11456 );
xor \U$11081 ( \11458 , \10818 , \10875 );
xor \U$11082 ( \11459 , \11457 , \11458 );
not \U$11083 ( \11460 , \11459 );
or \U$11084 ( \11461 , \11408 , \11460 );
nand \U$11085 ( \11462 , \11458 , \11457 );
nand \U$11086 ( \11463 , \11461 , \11462 );
xor \U$11087 ( \11464 , \9373 , \9481 );
xnor \U$11088 ( \11465 , \11464 , \9572 );
nand \U$11089 ( \11466 , \11463 , \11465 );
and \U$11090 ( \11467 , \9821 , \9719 );
not \U$11091 ( \11468 , \9821 );
not \U$11092 ( \11469 , \9719 );
and \U$11093 ( \11470 , \11468 , \11469 );
nor \U$11094 ( \11471 , \11467 , \11470 );
xor \U$11095 ( \11472 , \11471 , \9654 );
and \U$11096 ( \11473 , \11466 , \11472 );
nor \U$11097 ( \11474 , \11463 , \11465 );
nor \U$11098 ( \11475 , \11473 , \11474 );
nand \U$11099 ( \11476 , \11356 , \11475 );
nand \U$11100 ( \11477 , \11353 , \11010 );
nand \U$11101 ( \11478 , \11476 , \11477 );
not \U$11102 ( \11479 , \11478 );
xor \U$11103 ( \11480 , \10721 , \11479 );
xor \U$11104 ( \11481 , \9972 , \9574 );
not \U$11105 ( \11482 , \9824 );
xnor \U$11106 ( \11483 , \11481 , \11482 );
xor \U$11107 ( \11484 , \10290 , \10302 );
xor \U$11108 ( \11485 , \11484 , \10241 );
not \U$11109 ( \11486 , \11485 );
not \U$11110 ( \11487 , \11434 );
not \U$11111 ( \11488 , \11424 );
or \U$11112 ( \11489 , \11487 , \11488 );
nand \U$11113 ( \11490 , \10690 , \10676 );
nand \U$11114 ( \11491 , \11489 , \11490 );
not \U$11115 ( \11492 , \5039 );
not \U$11116 ( \11493 , \10902 );
or \U$11117 ( \11494 , \11492 , \11493 );
nand \U$11118 ( \11495 , \10536 , \5049 );
nand \U$11119 ( \11496 , \11494 , \11495 );
nor \U$11120 ( \11497 , \11491 , \11496 );
not \U$11121 ( \11498 , \6276 );
not \U$11122 ( \11499 , \10885 );
or \U$11123 ( \11500 , \11498 , \11499 );
nand \U$11124 ( \11501 , \4853 , \10610 );
nand \U$11125 ( \11502 , \11500 , \11501 );
not \U$11126 ( \11503 , \11502 );
or \U$11127 ( \11504 , \11497 , \11503 );
nand \U$11128 ( \11505 , \11491 , \11496 );
nand \U$11129 ( \11506 , \11504 , \11505 );
nand \U$11130 ( \11507 , \11486 , \11506 );
not \U$11131 ( \11508 , \11506 );
nand \U$11132 ( \11509 , \11485 , \11508 );
nand \U$11133 ( \11510 , \11507 , \11509 );
not \U$11134 ( \11511 , \2450 );
not \U$11135 ( \11512 , \2563 );
and \U$11136 ( \11513 , RIae79778_151, \11512 );
not \U$11137 ( \11514 , RIae79778_151);
and \U$11138 ( \11515 , \11514 , \2676 );
nor \U$11139 ( \11516 , \11513 , \11515 );
not \U$11140 ( \11517 , \11516 );
or \U$11141 ( \11518 , \11511 , \11517 );
nand \U$11142 ( \11519 , \9588 , \9576 );
nand \U$11143 ( \11520 , \11518 , \11519 );
not \U$11144 ( \11521 , \11236 );
not \U$11145 ( \11522 , \11254 );
or \U$11146 ( \11523 , \11521 , \11522 );
not \U$11147 ( \11524 , \11249 );
nand \U$11148 ( \11525 , \11524 , \11246 );
nand \U$11149 ( \11526 , \11523 , \11525 );
xor \U$11150 ( \11527 , \11520 , \11526 );
not \U$11151 ( \11528 , \9622 );
not \U$11152 ( \11529 , RIae7a3a8_177);
not \U$11153 ( \11530 , \1178 );
not \U$11154 ( \11531 , \1180 );
and \U$11155 ( \11532 , \11530 , \11531 );
and \U$11156 ( \11533 , \1178 , \1180 );
nor \U$11157 ( \11534 , \11532 , \11533 );
not \U$11158 ( \11535 , \11534 );
or \U$11159 ( \11536 , \11529 , \11535 );
not \U$11160 ( \11537 , \11534 );
not \U$11161 ( \11538 , \11537 );
or \U$11162 ( \11539 , \11538 , RIae7a3a8_177);
nand \U$11163 ( \11540 , \11536 , \11539 );
not \U$11164 ( \11541 , \11540 );
or \U$11165 ( \11542 , \11528 , \11541 );
nand \U$11166 ( \11543 , \9629 , \9644 );
nand \U$11167 ( \11544 , \11542 , \11543 );
xnor \U$11168 ( \11545 , \11527 , \11544 );
not \U$11169 ( \11546 , \11545 );
and \U$11170 ( \11547 , \11510 , \11546 );
not \U$11171 ( \11548 , \11510 );
and \U$11172 ( \11549 , \11548 , \11545 );
nor \U$11173 ( \11550 , \11547 , \11549 );
not \U$11174 ( \11551 , \11364 );
not \U$11175 ( \11552 , \11361 );
or \U$11176 ( \11553 , \11551 , \11552 );
and \U$11177 ( \11554 , RIae79c28_161, \2786 );
not \U$11178 ( \11555 , RIae79c28_161);
and \U$11179 ( \11556 , \11555 , \2093 );
or \U$11180 ( \11557 , \11554 , \11556 );
nand \U$11181 ( \11558 , \11557 , \2767 );
nand \U$11182 ( \11559 , \11553 , \11558 );
not \U$11183 ( \11560 , \11559 );
not \U$11184 ( \11561 , \1008 );
not \U$11185 ( \11562 , \10066 );
and \U$11186 ( \11563 , RIae79160_138, \11562 );
not \U$11187 ( \11564 , RIae79160_138);
and \U$11188 ( \11565 , \11564 , \10070 );
or \U$11189 ( \11566 , \11563 , \11565 );
not \U$11190 ( \11567 , \11566 );
or \U$11191 ( \11568 , \11561 , \11567 );
nand \U$11192 ( \11569 , \11391 , \1012 );
nand \U$11193 ( \11570 , \11568 , \11569 );
not \U$11194 ( \11571 , \11570 );
not \U$11195 ( \11572 , \926 );
not \U$11196 ( \11573 , \10868 );
or \U$11197 ( \11574 , \11572 , \11573 );
not \U$11198 ( \11575 , \1286 );
buf \U$11199 ( \11576 , \10192 );
not \U$11200 ( \11577 , \11576 );
not \U$11201 ( \11578 , \11577 );
not \U$11202 ( \11579 , \11578 );
or \U$11203 ( \11580 , \11575 , \11579 );
not \U$11204 ( \11581 , \11576 );
nand \U$11205 ( \11582 , \11581 , RIae78bc0_126);
nand \U$11206 ( \11583 , \11580 , \11582 );
nand \U$11207 ( \11584 , \11583 , \951 );
nand \U$11208 ( \11585 , \11574 , \11584 );
not \U$11209 ( \11586 , \1086 );
and \U$11210 ( \11587 , RIae78e90_132, \10338 );
not \U$11211 ( \11588 , RIae78e90_132);
not \U$11212 ( \11589 , \10031 );
and \U$11213 ( \11590 , \11588 , \11589 );
nor \U$11214 ( \11591 , \11587 , \11590 );
not \U$11215 ( \11592 , \11591 );
or \U$11216 ( \11593 , \11586 , \11592 );
nand \U$11217 ( \11594 , \11378 , \1072 );
nand \U$11218 ( \11595 , \11593 , \11594 );
xor \U$11219 ( \11596 , \11585 , \11595 );
not \U$11220 ( \11597 , \11596 );
or \U$11221 ( \11598 , \11571 , \11597 );
nand \U$11222 ( \11599 , \11595 , \11585 );
nand \U$11223 ( \11600 , \11598 , \11599 );
not \U$11224 ( \11601 , \11600 );
and \U$11225 ( \11602 , \10870 , \10853 );
not \U$11226 ( \11603 , \10870 );
not \U$11227 ( \11604 , \10853 );
and \U$11228 ( \11605 , \11603 , \11604 );
nor \U$11229 ( \11606 , \11602 , \11605 );
not \U$11230 ( \11607 , \11606 );
and \U$11231 ( \11608 , \11601 , \11607 );
not \U$11232 ( \11609 , \11601 );
and \U$11233 ( \11610 , \11609 , \11606 );
nor \U$11234 ( \11611 , \11608 , \11610 );
not \U$11235 ( \11612 , \11611 );
or \U$11236 ( \11613 , \11560 , \11612 );
nand \U$11237 ( \11614 , \11600 , \11606 );
nand \U$11238 ( \11615 , \11613 , \11614 );
not \U$11239 ( \11616 , \11615 );
xor \U$11240 ( \11617 , \9677 , \9702 );
xnor \U$11241 ( \11618 , \11617 , \9715 );
not \U$11242 ( \11619 , \11618 );
or \U$11243 ( \11620 , \11616 , \11619 );
not \U$11244 ( \11621 , \9747 );
not \U$11245 ( \11622 , \9779 );
or \U$11246 ( \11623 , \11621 , \11622 );
or \U$11247 ( \11624 , \9779 , \9747 );
nand \U$11248 ( \11625 , \11623 , \11624 );
and \U$11249 ( \11626 , \11625 , \9817 );
not \U$11250 ( \11627 , \11625 );
and \U$11251 ( \11628 , \11627 , \9818 );
nor \U$11252 ( \11629 , \11626 , \11628 );
nand \U$11253 ( \11630 , \11620 , \11629 );
not \U$11254 ( \11631 , \11618 );
not \U$11255 ( \11632 , \11615 );
nand \U$11256 ( \11633 , \11631 , \11632 );
buf \U$11257 ( \11634 , \11633 );
nand \U$11258 ( \11635 , \11630 , \11634 );
and \U$11259 ( \11636 , \11550 , \11635 );
xor \U$11260 ( \11637 , \9590 , \9617 );
xnor \U$11261 ( \11638 , \11637 , \9646 );
xor \U$11262 ( \11639 , \11496 , \11491 );
xor \U$11263 ( \11640 , \11639 , \11503 );
xor \U$11264 ( \11641 , \11638 , \11640 );
xor \U$11265 ( \11642 , \9551 , \9567 );
xnor \U$11266 ( \11643 , \11642 , \9520 );
and \U$11267 ( \11644 , \11641 , \11643 );
and \U$11268 ( \11645 , \11638 , \11640 );
or \U$11269 ( \11646 , \11644 , \11645 );
or \U$11270 ( \11647 , \11636 , \11646 );
or \U$11271 ( \11648 , \11550 , \11635 );
nand \U$11272 ( \11649 , \11647 , \11648 );
xor \U$11273 ( \11650 , \11483 , \11649 );
not \U$11274 ( \11651 , \11507 );
not \U$11275 ( \11652 , \11545 );
or \U$11276 ( \11653 , \11651 , \11652 );
buf \U$11277 ( \11654 , \11509 );
nand \U$11278 ( \11655 , \11653 , \11654 );
not \U$11279 ( \11656 , \892 );
not \U$11280 ( \11657 , \10036 );
or \U$11281 ( \11658 , \11656 , \11657 );
and \U$11282 ( \11659 , RIae78b48_125, \10149 );
not \U$11283 ( \11660 , RIae78b48_125);
and \U$11284 ( \11661 , \11660 , \10142 );
or \U$11285 ( \11662 , \11659 , \11661 );
nand \U$11286 ( \11663 , \11662 , \867 );
nand \U$11287 ( \11664 , \11658 , \11663 );
buf \U$11288 ( \11665 , \10042 );
and \U$11289 ( \11666 , \11665 , RIae78b48_125);
nand \U$11290 ( \11667 , RIae7a858_187, RIae7a8d0_188);
and \U$11291 ( \11668 , \11667 , RIae7a6f0_184);
not \U$11292 ( \11669 , \11668 );
and \U$11293 ( \11670 , \11666 , \11669 );
not \U$11294 ( \11671 , \11666 );
and \U$11295 ( \11672 , \11671 , \11668 );
nor \U$11296 ( \11673 , \11670 , \11672 );
xor \U$11297 ( \11674 , \11664 , \11673 );
not \U$11298 ( \11675 , \2432 );
not \U$11299 ( \11676 , \11516 );
or \U$11300 ( \11677 , \11675 , \11676 );
and \U$11301 ( \11678 , RIae79778_151, \10583 );
not \U$11302 ( \11679 , RIae79778_151);
not \U$11303 ( \11680 , \1788 );
not \U$11304 ( \11681 , \11680 );
and \U$11305 ( \11682 , \11679 , \11681 );
nor \U$11306 ( \11683 , \11678 , \11682 );
nand \U$11307 ( \11684 , \11683 , \2450 );
nand \U$11308 ( \11685 , \11677 , \11684 );
xor \U$11309 ( \11686 , \11674 , \11685 );
not \U$11310 ( \11687 , \11540 );
not \U$11311 ( \11688 , \9644 );
or \U$11312 ( \11689 , \11687 , \11688 );
not \U$11313 ( \11690 , RIae7a3a8_177);
not \U$11314 ( \11691 , \11690 );
not \U$11315 ( \11692 , \11429 );
or \U$11316 ( \11693 , \11691 , \11692 );
not \U$11317 ( \11694 , \974 );
not \U$11318 ( \11695 , RIae7a3a8_177);
or \U$11319 ( \11696 , \11694 , \11695 );
nand \U$11320 ( \11697 , \11693 , \11696 );
nand \U$11321 ( \11698 , \11697 , \9622 );
nand \U$11322 ( \11699 , \11689 , \11698 );
xor \U$11323 ( \11700 , \11686 , \11699 );
not \U$11324 ( \11701 , \11700 );
not \U$11325 ( \11702 , \10367 );
not \U$11326 ( \11703 , \10379 );
or \U$11327 ( \11704 , \11702 , \11703 );
nand \U$11328 ( \11705 , \10368 , \10378 );
nand \U$11329 ( \11706 , \11704 , \11705 );
xnor \U$11330 ( \11707 , \11706 , \10392 );
not \U$11331 ( \11708 , \11707 );
xor \U$11332 ( \11709 , \10413 , \10425 );
xor \U$11333 ( \11710 , \11709 , \10431 );
not \U$11334 ( \11711 , \11710 );
or \U$11335 ( \11712 , \11708 , \11711 );
or \U$11336 ( \11713 , \11707 , \11710 );
nand \U$11337 ( \11714 , \11712 , \11713 );
not \U$11338 ( \11715 , \11714 );
or \U$11339 ( \11716 , \11701 , \11715 );
or \U$11340 ( \11717 , \11714 , \11700 );
nand \U$11341 ( \11718 , \11716 , \11717 );
xor \U$11342 ( \11719 , \11655 , \11718 );
xor \U$11343 ( \11720 , \10498 , \10508 );
xor \U$11344 ( \11721 , \11720 , \10521 );
not \U$11345 ( \11722 , \11721 );
not \U$11346 ( \11723 , \10612 );
not \U$11347 ( \11724 , \10596 );
or \U$11348 ( \11725 , \11723 , \11724 );
nand \U$11349 ( \11726 , \10595 , \10613 );
nand \U$11350 ( \11727 , \11725 , \11726 );
and \U$11351 ( \11728 , \11727 , \10652 );
not \U$11352 ( \11729 , \11727 );
not \U$11353 ( \11730 , \10652 );
and \U$11354 ( \11731 , \11729 , \11730 );
nor \U$11355 ( \11732 , \11728 , \11731 );
xor \U$11356 ( \11733 , \10450 , \10469 );
not \U$11357 ( \11734 , \10476 );
xor \U$11358 ( \11735 , \11733 , \11734 );
or \U$11359 ( \11736 , \11732 , \11735 );
and \U$11360 ( \11737 , \11722 , \11736 );
and \U$11361 ( \11738 , \11735 , \11732 );
nor \U$11362 ( \11739 , \11737 , \11738 );
xor \U$11363 ( \11740 , \11719 , \11739 );
and \U$11364 ( \11741 , \11650 , \11740 );
and \U$11365 ( \11742 , \11483 , \11649 );
or \U$11366 ( \11743 , \11741 , \11742 );
buf \U$11367 ( \11744 , \11743 );
and \U$11368 ( \11745 , \11480 , \11744 );
not \U$11369 ( \11746 , \11480 );
not \U$11370 ( \11747 , \11744 );
and \U$11371 ( \11748 , \11746 , \11747 );
nor \U$11372 ( \11749 , \11745 , \11748 );
not \U$11373 ( \11750 , \11749 );
not \U$11374 ( \11751 , \4853 );
not \U$11375 ( \11752 , RIae79ca0_162);
not \U$11376 ( \11753 , \10534 );
or \U$11377 ( \11754 , \11752 , \11753 );
not \U$11378 ( \11755 , RIae79ca0_162);
nand \U$11379 ( \11756 , \3747 , \11755 );
nand \U$11380 ( \11757 , \11754 , \11756 );
not \U$11381 ( \11758 , \11757 );
or \U$11382 ( \11759 , \11751 , \11758 );
not \U$11383 ( \11760 , \4154 );
not \U$11384 ( \11761 , \11760 );
buf \U$11385 ( \11762 , \11761 );
nand \U$11386 ( \11763 , \10602 , \11762 );
nand \U$11387 ( \11764 , \11759 , \11763 );
not \U$11388 ( \11765 , \11764 );
not \U$11389 ( \11766 , \2767 );
not \U$11390 ( \11767 , \10593 );
or \U$11391 ( \11768 , \11766 , \11767 );
and \U$11392 ( \11769 , RIae79c28_161, \10608 );
not \U$11393 ( \11770 , RIae79c28_161);
and \U$11394 ( \11771 , \11770 , \10605 );
or \U$11395 ( \11772 , \11769 , \11771 );
nand \U$11396 ( \11773 , \11772 , \2776 );
nand \U$11397 ( \11774 , \11768 , \11773 );
not \U$11398 ( \11775 , \11774 );
or \U$11399 ( \11776 , \11765 , \11775 );
or \U$11400 ( \11777 , \11774 , \11764 );
nand \U$11401 ( \11778 , \11776 , \11777 );
not \U$11402 ( \11779 , \10927 );
not \U$11403 ( \11780 , \10623 );
or \U$11404 ( \11781 , \11779 , \11780 );
not \U$11405 ( \11782 , \10633 );
not \U$11406 ( \11783 , \2178 );
or \U$11407 ( \11784 , \11782 , \11783 );
or \U$11408 ( \11785 , \5351 , \10633 );
nand \U$11409 ( \11786 , \11784 , \11785 );
nand \U$11410 ( \11787 , \11786 , \10631 );
nand \U$11411 ( \11788 , \11781 , \11787 );
xor \U$11412 ( \11789 , \11778 , \11788 );
not \U$11413 ( \11790 , \9699 );
and \U$11414 ( \11791 , RIae7a240_174, \2848 );
not \U$11415 ( \11792 , RIae7a240_174);
and \U$11416 ( \11793 , \11792 , \2847 );
nor \U$11417 ( \11794 , \11791 , \11793 );
not \U$11418 ( \11795 , \11794 );
or \U$11419 ( \11796 , \11790 , \11795 );
nand \U$11420 ( \11797 , \10448 , \9688 );
nand \U$11421 ( \11798 , \11796 , \11797 );
not \U$11422 ( \11799 , \1008 );
not \U$11423 ( \11800 , \10457 );
or \U$11424 ( \11801 , \11799 , \11800 );
not \U$11425 ( \11802 , RIae79160_138);
buf \U$11426 ( \11803 , \9415 );
not \U$11427 ( \11804 , \11803 );
not \U$11428 ( \11805 , \11804 );
or \U$11429 ( \11806 , \11802 , \11805 );
or \U$11430 ( \11807 , \11804 , RIae79160_138);
nand \U$11431 ( \11808 , \11806 , \11807 );
nand \U$11432 ( \11809 , \11808 , \10451 );
nand \U$11433 ( \11810 , \11801 , \11809 );
xnor \U$11434 ( \11811 , \11798 , \11810 );
not \U$11435 ( \11812 , \1988 );
not \U$11436 ( \11813 , \10472 );
or \U$11437 ( \11814 , \11812 , \11813 );
nand \U$11438 ( \11815 , \10107 , \2007 );
nand \U$11439 ( \11816 , \11814 , \11815 );
xor \U$11440 ( \11817 , \11811 , \11816 );
nand \U$11441 ( \11818 , \11789 , \11817 );
or \U$11442 ( \11819 , \11789 , \11817 );
nand \U$11443 ( \11820 , \11818 , \11819 );
not \U$11444 ( \11821 , \11520 );
or \U$11445 ( \11822 , \11544 , \11526 );
not \U$11446 ( \11823 , \11822 );
or \U$11447 ( \11824 , \11821 , \11823 );
nand \U$11448 ( \11825 , \11544 , \11526 );
nand \U$11449 ( \11826 , \11824 , \11825 );
buf \U$11450 ( \11827 , \11826 );
xor \U$11451 ( \11828 , \11820 , \11827 );
not \U$11452 ( \11829 , \11828 );
not \U$11453 ( \11830 , \2339 );
not \U$11454 ( \11831 , \10488 );
or \U$11455 ( \11832 , \11830 , \11831 );
not \U$11456 ( \11833 , RIae798e0_154);
not \U$11457 ( \11834 , \9672 );
or \U$11458 ( \11835 , \11833 , \11834 );
or \U$11459 ( \11836 , \9672 , RIae798e0_154);
nand \U$11460 ( \11837 , \11835 , \11836 );
nand \U$11461 ( \11838 , \2322 , \11837 );
nand \U$11462 ( \11839 , \11832 , \11838 );
not \U$11463 ( \11840 , \9814 );
not \U$11464 ( \11841 , RIae7a2b8_175);
not \U$11465 ( \11842 , \9696 );
or \U$11466 ( \11843 , \11841 , \11842 );
or \U$11467 ( \11844 , \3145 , RIae7a2b8_175);
nand \U$11468 ( \11845 , \11843 , \11844 );
not \U$11469 ( \11846 , \11845 );
or \U$11470 ( \11847 , \11840 , \11846 );
nand \U$11471 ( \11848 , \10504 , \9792 );
nand \U$11472 ( \11849 , \11847 , \11848 );
xor \U$11473 ( \11850 , \11839 , \11849 );
buf \U$11474 ( \11851 , \11439 );
not \U$11475 ( \11852 , \11851 );
not \U$11476 ( \11853 , \10518 );
or \U$11477 ( \11854 , \11852 , \11853 );
not \U$11478 ( \11855 , \818 );
not \U$11479 ( \11856 , \987 );
or \U$11480 ( \11857 , \11855 , \11856 );
nand \U$11481 ( \11858 , \11857 , \819 );
xor \U$11482 ( \11859 , RIae7a7e0_186, \11858 );
nand \U$11483 ( \11860 , \11859 , \9527 );
nand \U$11484 ( \11861 , \11854 , \11860 );
xor \U$11485 ( \11862 , \11850 , \11861 );
not \U$11486 ( \11863 , \5048 );
not \U$11487 ( \11864 , \4968 );
not \U$11488 ( \11865 , \2154 );
or \U$11489 ( \11866 , \11864 , \11865 );
nand \U$11490 ( \11867 , \2954 , RIae79d90_164);
nand \U$11491 ( \11868 , \11866 , \11867 );
not \U$11492 ( \11869 , \11868 );
or \U$11493 ( \11870 , \11863 , \11869 );
nand \U$11494 ( \11871 , \10539 , \6091 );
nand \U$11495 ( \11872 , \11870 , \11871 );
not \U$11496 ( \11873 , \9730 );
not \U$11497 ( \11874 , \10553 );
or \U$11498 ( \11875 , \11873 , \11874 );
and \U$11499 ( \11876 , RIae7a060_170, \6086 );
not \U$11500 ( \11877 , RIae7a060_170);
and \U$11501 ( \11878 , \11877 , \780 );
nor \U$11502 ( \11879 , \11876 , \11878 );
nand \U$11503 ( \11880 , \11879 , \9745 );
nand \U$11504 ( \11881 , \11875 , \11880 );
xor \U$11505 ( \11882 , \11872 , \11881 );
not \U$11506 ( \11883 , \6214 );
not \U$11507 ( \11884 , \6203 );
not \U$11508 ( \11885 , \2230 );
not \U$11509 ( \11886 , \11885 );
or \U$11510 ( \11887 , \11884 , \11886 );
not \U$11511 ( \11888 , \2230 );
or \U$11512 ( \11889 , \11888 , \6203 );
nand \U$11513 ( \11890 , \11887 , \11889 );
not \U$11514 ( \11891 , \11890 );
or \U$11515 ( \11892 , \11883 , \11891 );
nand \U$11516 ( \11893 , \10572 , \6201 );
nand \U$11517 ( \11894 , \11892 , \11893 );
xor \U$11518 ( \11895 , \11882 , \11894 );
xor \U$11519 ( \11896 , \11862 , \11895 );
and \U$11520 ( \11897 , \10664 , \9758 );
not \U$11521 ( \11898 , \9777 );
not \U$11522 ( \11899 , \2330 );
and \U$11523 ( \11900 , RIae7a150_172, \11899 );
not \U$11524 ( \11901 , RIae7a150_172);
and \U$11525 ( \11902 , \11901 , \2330 );
nor \U$11526 ( \11903 , \11900 , \11902 );
nor \U$11527 ( \11904 , \11898 , \11903 );
nor \U$11528 ( \11905 , \11897 , \11904 );
not \U$11529 ( \11906 , \10696 );
not \U$11530 ( \11907 , \10682 );
or \U$11531 ( \11908 , \11906 , \11907 );
xor \U$11532 ( \11909 , \9770 , RIae7a498_179);
nand \U$11533 ( \11910 , \11909 , \10675 );
nand \U$11534 ( \11911 , \11908 , \11910 );
xnor \U$11535 ( \11912 , \11905 , \11911 );
buf \U$11536 ( \11913 , \9499 );
buf \U$11537 ( \11914 , \11913 );
not \U$11538 ( \11915 , \11914 );
not \U$11539 ( \11916 , \10706 );
or \U$11540 ( \11917 , \11915 , \11916 );
not \U$11541 ( \11918 , RIae79fe8_169);
or \U$11542 ( \11919 , \1899 , \11918 );
nand \U$11543 ( \11920 , \11918 , \1899 );
nand \U$11544 ( \11921 , \11919 , \11920 );
nand \U$11545 ( \11922 , \9518 , \11921 );
nand \U$11546 ( \11923 , \11917 , \11922 );
xnor \U$11547 ( \11924 , \11912 , \11923 );
xor \U$11548 ( \11925 , \11896 , \11924 );
not \U$11549 ( \11926 , \11925 );
not \U$11550 ( \11927 , \11926 );
or \U$11551 ( \11928 , \11829 , \11927 );
not \U$11552 ( \11929 , \11828 );
nand \U$11553 ( \11930 , \11925 , \11929 );
nand \U$11554 ( \11931 , \11928 , \11930 );
nand \U$11555 ( \11932 , \10994 , \10992 );
not \U$11556 ( \11933 , \11932 );
not \U$11557 ( \11934 , \11002 );
or \U$11558 ( \11935 , \11933 , \11934 );
not \U$11559 ( \11936 , \10992 );
nand \U$11560 ( \11937 , \11936 , \10995 );
nand \U$11561 ( \11938 , \11935 , \11937 );
not \U$11562 ( \11939 , \10305 );
not \U$11563 ( \11940 , \10178 );
not \U$11564 ( \11941 , \10220 );
or \U$11565 ( \11942 , \11940 , \11941 );
or \U$11566 ( \11943 , \10220 , \10178 );
nand \U$11567 ( \11944 , \11942 , \11943 );
not \U$11568 ( \11945 , \11944 );
and \U$11569 ( \11946 , \11939 , \11945 );
and \U$11570 ( \11947 , \10305 , \11944 );
nor \U$11571 ( \11948 , \11946 , \11947 );
xor \U$11572 ( \11949 , \11938 , \11948 );
xor \U$11573 ( \11950 , \10763 , \10805 );
and \U$11574 ( \11951 , \11950 , \10879 );
and \U$11575 ( \11952 , \10763 , \10805 );
or \U$11576 ( \11953 , \11951 , \11952 );
xor \U$11577 ( \11954 , \11949 , \11953 );
buf \U$11578 ( \11955 , \11954 );
and \U$11579 ( \11956 , \11931 , \11955 );
not \U$11580 ( \11957 , \11931 );
not \U$11581 ( \11958 , \11955 );
and \U$11582 ( \11959 , \11957 , \11958 );
nor \U$11583 ( \11960 , \11956 , \11959 );
not \U$11584 ( \11961 , \11960 );
xor \U$11585 ( \11962 , \10480 , \10479 );
not \U$11586 ( \11963 , \10524 );
xor \U$11587 ( \11964 , \11962 , \11963 );
not \U$11588 ( \11965 , \11964 );
not \U$11589 ( \11966 , \10714 );
not \U$11590 ( \11967 , \10655 );
not \U$11591 ( \11968 , \10578 );
or \U$11592 ( \11969 , \11967 , \11968 );
or \U$11593 ( \11970 , \10578 , \10655 );
nand \U$11594 ( \11971 , \11969 , \11970 );
not \U$11595 ( \11972 , \11971 );
or \U$11596 ( \11973 , \11966 , \11972 );
or \U$11597 ( \11974 , \11971 , \10714 );
nand \U$11598 ( \11975 , \11973 , \11974 );
not \U$11599 ( \11976 , \11975 );
or \U$11600 ( \11977 , \11965 , \11976 );
or \U$11601 ( \11978 , \11975 , \11964 );
nand \U$11602 ( \11979 , \11977 , \11978 );
not \U$11603 ( \11980 , \11979 );
xor \U$11604 ( \11981 , \10541 , \10557 );
xor \U$11605 ( \11982 , \11981 , \10575 );
xor \U$11606 ( \11983 , \10669 , \10698 );
xor \U$11607 ( \11984 , \11983 , \10711 );
xor \U$11608 ( \11985 , \11982 , \11984 );
not \U$11609 ( \11986 , \11366 );
and \U$11610 ( \11987 , \11406 , \11397 );
not \U$11611 ( \11988 , \11406 );
and \U$11612 ( \11989 , \11988 , \11398 );
nor \U$11613 ( \11990 , \11987 , \11989 );
not \U$11614 ( \11991 , \11990 );
or \U$11615 ( \11992 , \11986 , \11991 );
nand \U$11616 ( \11993 , \11406 , \11397 );
nand \U$11617 ( \11994 , \11992 , \11993 );
and \U$11618 ( \11995 , \11985 , \11994 );
and \U$11619 ( \11996 , \11982 , \11984 );
or \U$11620 ( \11997 , \11995 , \11996 );
not \U$11621 ( \11998 , \11997 );
not \U$11622 ( \11999 , \11998 );
and \U$11623 ( \12000 , \11980 , \11999 );
and \U$11624 ( \12001 , \11979 , \11998 );
nor \U$11625 ( \12002 , \12000 , \12001 );
not \U$11626 ( \12003 , \12002 );
xor \U$11627 ( \12004 , \11735 , \11732 );
and \U$11628 ( \12005 , \12004 , \11722 );
not \U$11629 ( \12006 , \12004 );
and \U$11630 ( \12007 , \12006 , \11721 );
nor \U$11631 ( \12008 , \12005 , \12007 );
not \U$11632 ( \12009 , \12008 );
not \U$11633 ( \12010 , \12009 );
xor \U$11634 ( \12011 , \11982 , \11984 );
xor \U$11635 ( \12012 , \12011 , \11994 );
not \U$11636 ( \12013 , \12012 );
or \U$11637 ( \12014 , \12010 , \12013 );
not \U$11638 ( \12015 , \12012 );
not \U$11639 ( \12016 , \12015 );
not \U$11640 ( \12017 , \12008 );
or \U$11641 ( \12018 , \12016 , \12017 );
not \U$11642 ( \12019 , \11226 );
xor \U$11643 ( \12020 , \11348 , \12019 );
xnor \U$11644 ( \12021 , \12020 , \11142 );
nand \U$11645 ( \12022 , \12018 , \12021 );
nand \U$11646 ( \12023 , \12014 , \12022 );
not \U$11647 ( \12024 , \12023 );
or \U$11648 ( \12025 , \12003 , \12024 );
or \U$11649 ( \12026 , \12002 , \12023 );
nand \U$11650 ( \12027 , \12025 , \12026 );
not \U$11651 ( \12028 , \12027 );
or \U$11652 ( \12029 , \11961 , \12028 );
not \U$11653 ( \12030 , \12002 );
buf \U$11654 ( \12031 , \12023 );
nand \U$11655 ( \12032 , \12030 , \12031 );
nand \U$11656 ( \12033 , \12029 , \12032 );
not \U$11657 ( \12034 , \12033 );
not \U$11658 ( \12035 , \11718 );
not \U$11659 ( \12036 , \11655 );
or \U$11660 ( \12037 , \12035 , \12036 );
nand \U$11661 ( \12038 , \12037 , \11739 );
or \U$11662 ( \12039 , \11655 , \11718 );
nand \U$11663 ( \12040 , \12038 , \12039 );
xor \U$11664 ( \12041 , \11674 , \11685 );
and \U$11665 ( \12042 , \12041 , \11699 );
and \U$11666 ( \12043 , \11674 , \11685 );
or \U$11667 ( \12044 , \12042 , \12043 );
not \U$11668 ( \12045 , \1501 );
and \U$11669 ( \12046 , RIae79250_140, \9442 );
not \U$11670 ( \12047 , RIae79250_140);
and \U$11671 ( \12048 , \12047 , \9441 );
or \U$11672 ( \12049 , \12046 , \12048 );
not \U$11673 ( \12050 , \12049 );
or \U$11674 ( \12051 , \12045 , \12050 );
nand \U$11675 ( \12052 , \10365 , \9403 );
nand \U$11676 ( \12053 , \12051 , \12052 );
not \U$11677 ( \12054 , \2011 );
not \U$11678 ( \12055 , RIae79610_148);
not \U$11679 ( \12056 , \6230 );
not \U$11680 ( \12057 , \12056 );
or \U$11681 ( \12058 , \12055 , \12057 );
nand \U$11682 ( \12059 , \6230 , \2056 );
nand \U$11683 ( \12060 , \12058 , \12059 );
not \U$11684 ( \12061 , \12060 );
or \U$11685 ( \12062 , \12054 , \12061 );
nand \U$11686 ( \12063 , \10390 , \2063 );
nand \U$11687 ( \12064 , \12062 , \12063 );
xor \U$11688 ( \12065 , \12053 , \12064 );
not \U$11689 ( \12066 , \1863 );
not \U$11690 ( \12067 , \9347 );
xor \U$11691 ( \12068 , RIae793b8_143, \12067 );
not \U$11692 ( \12069 , \12068 );
or \U$11693 ( \12070 , \12066 , \12069 );
nand \U$11694 ( \12071 , \10376 , \1910 );
nand \U$11695 ( \12072 , \12070 , \12071 );
xnor \U$11696 ( \12073 , \12065 , \12072 );
not \U$11697 ( \12074 , \12073 );
xor \U$11698 ( \12075 , \12044 , \12074 );
not \U$11699 ( \12076 , \1049 );
buf \U$11700 ( \12077 , \9607 );
and \U$11701 ( \12078 , \12077 , RIae79070_136);
not \U$11702 ( \12079 , \12077 );
and \U$11703 ( \12080 , \12079 , \1039 );
nor \U$11704 ( \12081 , \12078 , \12080 );
not \U$11705 ( \12082 , \12081 );
or \U$11706 ( \12083 , \12076 , \12082 );
nand \U$11707 ( \12084 , \9946 , \1062 );
nand \U$11708 ( \12085 , \12083 , \12084 );
not \U$11709 ( \12086 , \12085 );
not \U$11710 ( \12087 , \1013 );
buf \U$11711 ( \12088 , \9395 );
xor \U$11712 ( \12089 , \12088 , RIae79160_138);
not \U$11713 ( \12090 , \12089 );
or \U$11714 ( \12091 , \12087 , \12090 );
nand \U$11715 ( \12092 , \11808 , \1008 );
nand \U$11716 ( \12093 , \12091 , \12092 );
xor \U$11717 ( \12094 , \12086 , \12093 );
not \U$11718 ( \12095 , \11851 );
not \U$11719 ( \12096 , \11859 );
or \U$11720 ( \12097 , \12095 , \12096 );
nand \U$11721 ( \12098 , \10519 , RIae7a7e0_186);
nand \U$11722 ( \12099 , \12097 , \12098 );
xnor \U$11723 ( \12100 , \12094 , \12099 );
xor \U$11724 ( \12101 , \12075 , \12100 );
not \U$11725 ( \12102 , \11923 );
not \U$11726 ( \12103 , \11912 );
or \U$11727 ( \12104 , \12102 , \12103 );
not \U$11728 ( \12105 , \11905 );
nand \U$11729 ( \12106 , \12105 , \11911 );
nand \U$11730 ( \12107 , \12104 , \12106 );
not \U$11731 ( \12108 , \838 );
not \U$11732 ( \12109 , RIae78f80_134);
not \U$11733 ( \12110 , \10724 );
or \U$11734 ( \12111 , \12109 , \12110 );
or \U$11735 ( \12112 , \10724 , RIae78f80_134);
nand \U$11736 ( \12113 , \12111 , \12112 );
not \U$11737 ( \12114 , \12113 );
or \U$11738 ( \12115 , \12108 , \12114 );
nand \U$11739 ( \12116 , \10089 , \797 );
nand \U$11740 ( \12117 , \12115 , \12116 );
not \U$11741 ( \12118 , \867 );
xor \U$11742 ( \12119 , RIae78b48_125, \10743 );
not \U$11743 ( \12120 , \12119 );
or \U$11744 ( \12121 , \12118 , \12120 );
nand \U$11745 ( \12122 , \11662 , \892 );
nand \U$11746 ( \12123 , \12121 , \12122 );
not \U$11747 ( \12124 , \1072 );
xor \U$11748 ( \12125 , RIae78e90_132, \10070 );
not \U$11749 ( \12126 , \12125 );
or \U$11750 ( \12127 , \12124 , \12126 );
nand \U$11751 ( \12128 , \9902 , \1086 );
nand \U$11752 ( \12129 , \12127 , \12128 );
not \U$11753 ( \12130 , \12129 );
xnor \U$11754 ( \12131 , \12123 , \12130 );
xor \U$11755 ( \12132 , \12117 , \12131 );
not \U$11756 ( \12133 , \11810 );
not \U$11757 ( \12134 , \11816 );
or \U$11758 ( \12135 , \12133 , \12134 );
or \U$11759 ( \12136 , \11816 , \11810 );
nand \U$11760 ( \12137 , \12136 , \11798 );
nand \U$11761 ( \12138 , \12135 , \12137 );
and \U$11762 ( \12139 , \12132 , \12138 );
not \U$11763 ( \12140 , \12132 );
not \U$11764 ( \12141 , \12138 );
and \U$11765 ( \12142 , \12140 , \12141 );
nor \U$11766 ( \12143 , \12139 , \12142 );
xnor \U$11767 ( \12144 , \12107 , \12143 );
xor \U$11768 ( \12145 , \12101 , \12144 );
not \U$11769 ( \12146 , \11700 );
not \U$11770 ( \12147 , \11710 );
nand \U$11771 ( \12148 , \12147 , \11707 );
not \U$11772 ( \12149 , \12148 );
or \U$11773 ( \12150 , \12146 , \12149 );
or \U$11774 ( \12151 , \11707 , \12147 );
nand \U$11775 ( \12152 , \12150 , \12151 );
xor \U$11776 ( \12153 , \12145 , \12152 );
xor \U$11777 ( \12154 , \12040 , \12153 );
not \U$11778 ( \12155 , \11997 );
not \U$11779 ( \12156 , \11979 );
or \U$11780 ( \12157 , \12155 , \12156 );
not \U$11781 ( \12158 , \11964 );
nand \U$11782 ( \12159 , \12158 , \11975 );
nand \U$11783 ( \12160 , \12157 , \12159 );
not \U$11784 ( \12161 , \12160 );
xnor \U$11785 ( \12162 , \12154 , \12161 );
not \U$11786 ( \12163 , \12162 );
or \U$11787 ( \12164 , \12034 , \12163 );
not \U$11788 ( \12165 , \12033 );
xor \U$11789 ( \12166 , \12040 , \12153 );
xor \U$11790 ( \12167 , \12166 , \12161 );
nand \U$11791 ( \12168 , \12165 , \12167 );
nand \U$11792 ( \12169 , \12164 , \12168 );
not \U$11793 ( \12170 , \1919 );
not \U$11794 ( \12171 , RIae794a8_145);
not \U$11795 ( \12172 , \1859 );
or \U$11796 ( \12173 , \12171 , \12172 );
or \U$11797 ( \12174 , \1859 , RIae794a8_145);
nand \U$11798 ( \12175 , \12173 , \12174 );
not \U$11799 ( \12176 , \12175 );
or \U$11800 ( \12177 , \12170 , \12176 );
nand \U$11801 ( \12178 , \9841 , \2457 );
nand \U$11802 ( \12179 , \12177 , \12178 );
not \U$11803 ( \12180 , \9792 );
not \U$11804 ( \12181 , \11845 );
or \U$11805 ( \12182 , \12180 , \12181 );
not \U$11806 ( \12183 , \2025 );
not \U$11807 ( \12184 , RIae7a2b8_175);
and \U$11808 ( \12185 , \12183 , \12184 );
not \U$11809 ( \12186 , \12183 );
and \U$11810 ( \12187 , \12186 , RIae7a2b8_175);
nor \U$11811 ( \12188 , \12185 , \12187 );
nand \U$11812 ( \12189 , \12188 , \9814 );
nand \U$11813 ( \12190 , \12182 , \12189 );
xor \U$11814 ( \12191 , \12179 , \12190 );
not \U$11815 ( \12192 , \2322 );
and \U$11816 ( \12193 , \5912 , RIae798e0_154);
not \U$11817 ( \12194 , \5912 );
and \U$11818 ( \12195 , \12194 , \2334 );
nor \U$11819 ( \12196 , \12193 , \12195 );
not \U$11820 ( \12197 , \12196 );
or \U$11821 ( \12198 , \12192 , \12197 );
nand \U$11822 ( \12199 , \10807 , \11837 );
nand \U$11823 ( \12200 , \12198 , \12199 );
xor \U$11824 ( \12201 , \12191 , \12200 );
not \U$11825 ( \12202 , \6214 );
not \U$11826 ( \12203 , RIae79ef8_167);
not \U$11827 ( \12204 , \2629 );
or \U$11828 ( \12205 , \12203 , \12204 );
buf \U$11829 ( \12206 , \2206 );
not \U$11830 ( \12207 , \12206 );
not \U$11831 ( \12208 , \12207 );
not \U$11832 ( \12209 , RIae79ef8_167);
nand \U$11833 ( \12210 , \12208 , \12209 );
nand \U$11834 ( \12211 , \12205 , \12210 );
not \U$11835 ( \12212 , \12211 );
or \U$11836 ( \12213 , \12202 , \12212 );
nand \U$11837 ( \12214 , \11890 , \6201 );
nand \U$11838 ( \12215 , \12213 , \12214 );
not \U$11839 ( \12216 , \12215 );
not \U$11840 ( \12217 , \5048 );
not \U$11841 ( \12218 , \6084 );
not \U$11842 ( \12219 , \9501 );
or \U$11843 ( \12220 , \12218 , \12219 );
nand \U$11844 ( \12221 , \2140 , RIae79d90_164);
nand \U$11845 ( \12222 , \12220 , \12221 );
not \U$11846 ( \12223 , \12222 );
or \U$11847 ( \12224 , \12217 , \12223 );
nand \U$11848 ( \12225 , \11868 , \6091 );
nand \U$11849 ( \12226 , \12224 , \12225 );
not \U$11850 ( \12227 , \12226 );
not \U$11851 ( \12228 , \12227 );
or \U$11852 ( \12229 , \12216 , \12228 );
or \U$11853 ( \12230 , \12227 , \12215 );
nand \U$11854 ( \12231 , \12229 , \12230 );
not \U$11855 ( \12232 , \10631 );
not \U$11856 ( \12233 , \12232 );
not \U$11857 ( \12234 , \12233 );
and \U$11858 ( \12235 , \9761 , RIae7a510_180);
not \U$11859 ( \12236 , \9761 );
and \U$11860 ( \12237 , \12236 , \10633 );
nor \U$11861 ( \12238 , \12235 , \12237 );
not \U$11862 ( \12239 , \12238 );
or \U$11863 ( \12240 , \12234 , \12239 );
nand \U$11864 ( \12241 , \11786 , \11400 );
nand \U$11865 ( \12242 , \12240 , \12241 );
and \U$11866 ( \12243 , \12231 , \12242 );
not \U$11867 ( \12244 , \12231 );
not \U$11868 ( \12245 , \12242 );
and \U$11869 ( \12246 , \12244 , \12245 );
nor \U$11870 ( \12247 , \12243 , \12246 );
xor \U$11871 ( \12248 , \12201 , \12247 );
not \U$11872 ( \12249 , \4853 );
not \U$11873 ( \12250 , \2406 );
not \U$11874 ( \12251 , \2310 );
or \U$11875 ( \12252 , \12250 , \12251 );
or \U$11876 ( \12253 , \2310 , \6270 );
nand \U$11877 ( \12254 , \12252 , \12253 );
not \U$11878 ( \12255 , \12254 );
or \U$11879 ( \12256 , \12249 , \12255 );
nand \U$11880 ( \12257 , \11757 , \6276 );
nand \U$11881 ( \12258 , \12256 , \12257 );
not \U$11882 ( \12259 , RIae7a150_172);
not \U$11883 ( \12260 , \3999 );
or \U$11884 ( \12261 , \12259 , \12260 );
buf \U$11885 ( \12262 , \2323 );
nand \U$11886 ( \12263 , \12262 , \10672 );
nand \U$11887 ( \12264 , \12261 , \12263 );
not \U$11888 ( \12265 , \12264 );
not \U$11889 ( \12266 , \9777 );
or \U$11890 ( \12267 , \12265 , \12266 );
not \U$11891 ( \12268 , \11903 );
nand \U$11892 ( \12269 , \12268 , \11087 );
nand \U$11893 ( \12270 , \12267 , \12269 );
xor \U$11894 ( \12271 , \12258 , \12270 );
xnor \U$11895 ( \12272 , RIae7a3a8_177, \1119 );
not \U$11896 ( \12273 , \12272 );
not \U$11897 ( \12274 , \9621 );
or \U$11898 ( \12275 , \12273 , \12274 );
nand \U$11899 ( \12276 , \11697 , \11014 );
nand \U$11900 ( \12277 , \12275 , \12276 );
xor \U$11901 ( \12278 , \12271 , \12277 );
xor \U$11902 ( \12279 , \12248 , \12278 );
not \U$11903 ( \12280 , \11938 );
not \U$11904 ( \12281 , \11948 );
nand \U$11905 ( \12282 , \12280 , \12281 );
not \U$11906 ( \12283 , \12282 );
not \U$11907 ( \12284 , \11953 );
or \U$11908 ( \12285 , \12283 , \12284 );
nand \U$11909 ( \12286 , \11948 , \11938 );
nand \U$11910 ( \12287 , \12285 , \12286 );
not \U$11911 ( \12288 , \12287 );
not \U$11912 ( \12289 , \2776 );
not \U$11913 ( \12290 , RIae79c28_161);
not \U$11914 ( \12291 , \1741 );
or \U$11915 ( \12292 , \12290 , \12291 );
nand \U$11916 ( \12293 , \4431 , \10584 );
nand \U$11917 ( \12294 , \12292 , \12293 );
not \U$11918 ( \12295 , \12294 );
or \U$11919 ( \12296 , \12289 , \12295 );
nand \U$11920 ( \12297 , \11772 , \2767 );
nand \U$11921 ( \12298 , \12296 , \12297 );
not \U$11922 ( \12299 , \2432 );
not \U$11923 ( \12300 , \11683 );
or \U$11924 ( \12301 , \12299 , \12300 );
and \U$11925 ( \12302 , RIae79778_151, \10883 );
not \U$11926 ( \12303 , RIae79778_151);
and \U$11927 ( \12304 , \12303 , \3529 );
or \U$11928 ( \12305 , \12302 , \12304 );
nand \U$11929 ( \12306 , \12305 , \11037 );
nand \U$11930 ( \12307 , \12301 , \12306 );
not \U$11931 ( \12308 , \12307 );
not \U$11932 ( \12309 , \11114 );
not \U$11933 ( \12310 , \11537 );
or \U$11934 ( \12311 , \12309 , \12310 );
not \U$11935 ( \12312 , RIae7a240_174);
or \U$11936 ( \12313 , \11537 , \12312 );
nand \U$11937 ( \12314 , \12311 , \12313 );
nand \U$11938 ( \12315 , \12314 , \9699 );
nand \U$11939 ( \12316 , \11794 , \9688 );
nand \U$11940 ( \12317 , \12315 , \12316 );
not \U$11941 ( \12318 , \12317 );
not \U$11942 ( \12319 , \12318 );
or \U$11943 ( \12320 , \12308 , \12319 );
not \U$11944 ( \12321 , \12316 );
not \U$11945 ( \12322 , \12315 );
or \U$11946 ( \12323 , \12321 , \12322 );
not \U$11947 ( \12324 , \12307 );
nand \U$11948 ( \12325 , \12323 , \12324 );
nand \U$11949 ( \12326 , \12320 , \12325 );
xor \U$11950 ( \12327 , \12298 , \12326 );
not \U$11951 ( \12328 , \11673 );
not \U$11952 ( \12329 , \11664 );
or \U$11953 ( \12330 , \12328 , \12329 );
nand \U$11954 ( \12331 , \11666 , \11669 );
nand \U$11955 ( \12332 , \12330 , \12331 );
not \U$11956 ( \12333 , \12332 );
not \U$11957 ( \12334 , \9279 );
and \U$11958 ( \12335 , RIae79688_149, \12334 );
not \U$11959 ( \12336 , RIae79688_149);
and \U$11960 ( \12337 , \12336 , \5722 );
or \U$11961 ( \12338 , \12335 , \12337 );
and \U$11962 ( \12339 , \12338 , \1820 );
and \U$11963 ( \12340 , \10411 , \9320 );
nor \U$11964 ( \12341 , \12339 , \12340 );
not \U$11965 ( \12342 , \12341 );
or \U$11966 ( \12343 , \12333 , \12342 );
not \U$11967 ( \12344 , \12340 );
not \U$11968 ( \12345 , \12344 );
nand \U$11969 ( \12346 , \12338 , \1820 );
not \U$11970 ( \12347 , \12346 );
or \U$11971 ( \12348 , \12345 , \12347 );
not \U$11972 ( \12349 , \12332 );
nand \U$11973 ( \12350 , \12348 , \12349 );
nand \U$11974 ( \12351 , \12343 , \12350 );
not \U$11975 ( \12352 , \10414 );
not \U$11976 ( \12353 , RIae79ac0_158);
xor \U$11977 ( \12354 , \10226 , \12353 );
not \U$11978 ( \12355 , \12354 );
or \U$11979 ( \12356 , \12352 , \12355 );
nand \U$11980 ( \12357 , \10421 , \2272 );
nand \U$11981 ( \12358 , \12356 , \12357 );
xnor \U$11982 ( \12359 , \12351 , \12358 );
xnor \U$11983 ( \12360 , \12327 , \12359 );
buf \U$11984 ( \12361 , \12360 );
not \U$11985 ( \12362 , \9517 );
and \U$11986 ( \12363 , \5944 , RIae79fe8_169);
not \U$11987 ( \12364 , \5944 );
and \U$11988 ( \12365 , \12364 , \9504 );
nor \U$11989 ( \12366 , \12363 , \12365 );
not \U$11990 ( \12367 , \12366 );
or \U$11991 ( \12368 , \12362 , \12367 );
nand \U$11992 ( \12369 , \11921 , \10709 );
nand \U$11993 ( \12370 , \12368 , \12369 );
buf \U$11994 ( \12371 , \10676 );
not \U$11995 ( \12372 , \12371 );
not \U$11996 ( \12373 , \10625 );
not \U$11997 ( \12374 , \5957 );
or \U$11998 ( \12375 , \12373 , \12374 );
or \U$11999 ( \12376 , \918 , \10625 );
nand \U$12000 ( \12377 , \12375 , \12376 );
not \U$12001 ( \12378 , \12377 );
or \U$12002 ( \12379 , \12372 , \12378 );
nand \U$12003 ( \12380 , \11909 , \10696 );
nand \U$12004 ( \12381 , \12379 , \12380 );
xor \U$12005 ( \12382 , \12370 , \12381 );
not \U$12006 ( \12383 , \9730 );
not \U$12007 ( \12384 , \11879 );
or \U$12008 ( \12385 , \12383 , \12384 );
and \U$12009 ( \12386 , RIae7a060_170, \833 );
not \U$12010 ( \12387 , RIae7a060_170);
and \U$12011 ( \12388 , \12387 , \827 );
nor \U$12012 ( \12389 , \12386 , \12388 );
nand \U$12013 ( \12390 , \12389 , \9745 );
nand \U$12014 ( \12391 , \12385 , \12390 );
xor \U$12015 ( \12392 , \12382 , \12391 );
not \U$12016 ( \12393 , \12392 );
and \U$12017 ( \12394 , \12361 , \12393 );
not \U$12018 ( \12395 , \12361 );
not \U$12019 ( \12396 , \12393 );
and \U$12020 ( \12397 , \12395 , \12396 );
nor \U$12021 ( \12398 , \12394 , \12397 );
not \U$12022 ( \12399 , \12398 );
and \U$12023 ( \12400 , \12288 , \12399 );
and \U$12024 ( \12401 , \12287 , \12398 );
nor \U$12025 ( \12402 , \12400 , \12401 );
xnor \U$12026 ( \12403 , \12279 , \12402 );
not \U$12027 ( \12404 , \11828 );
not \U$12028 ( \12405 , \11925 );
or \U$12029 ( \12406 , \12404 , \12405 );
nand \U$12030 ( \12407 , \12406 , \11954 );
nand \U$12031 ( \12408 , \11926 , \11929 );
nand \U$12032 ( \12409 , \12407 , \12408 );
not \U$12033 ( \12410 , \12409 );
not \U$12034 ( \12411 , \11818 );
not \U$12035 ( \12412 , \11826 );
or \U$12036 ( \12413 , \12411 , \12412 );
nand \U$12037 ( \12414 , \12413 , \11819 );
not \U$12038 ( \12415 , \12414 );
xor \U$12039 ( \12416 , \11839 , \11849 );
and \U$12040 ( \12417 , \12416 , \11861 );
and \U$12041 ( \12418 , \11839 , \11849 );
or \U$12042 ( \12419 , \12417 , \12418 );
not \U$12043 ( \12420 , \11788 );
not \U$12044 ( \12421 , \11774 );
not \U$12045 ( \12422 , \11764 );
nand \U$12046 ( \12423 , \12421 , \12422 );
not \U$12047 ( \12424 , \12423 );
or \U$12048 ( \12425 , \12420 , \12424 );
nand \U$12049 ( \12426 , \11774 , \11764 );
nand \U$12050 ( \12427 , \12425 , \12426 );
not \U$12051 ( \12428 , \12427 );
xor \U$12052 ( \12429 , \12419 , \12428 );
not \U$12053 ( \12430 , \11872 );
not \U$12054 ( \12431 , \11894 );
or \U$12055 ( \12432 , \12430 , \12431 );
or \U$12056 ( \12433 , \11894 , \11872 );
nand \U$12057 ( \12434 , \12433 , \11881 );
nand \U$12058 ( \12435 , \12432 , \12434 );
xor \U$12059 ( \12436 , \12429 , \12435 );
not \U$12060 ( \12437 , \12436 );
or \U$12061 ( \12438 , \12415 , \12437 );
or \U$12062 ( \12439 , \12414 , \12436 );
nand \U$12063 ( \12440 , \12438 , \12439 );
not \U$12064 ( \12441 , \12440 );
nor \U$12065 ( \12442 , \11895 , \11862 );
or \U$12066 ( \12443 , \12442 , \11924 );
nand \U$12067 ( \12444 , \11895 , \11862 );
nand \U$12068 ( \12445 , \12443 , \12444 );
not \U$12069 ( \12446 , \12445 );
not \U$12070 ( \12447 , \12446 );
and \U$12071 ( \12448 , \12441 , \12447 );
and \U$12072 ( \12449 , \12440 , \12446 );
nor \U$12073 ( \12450 , \12448 , \12449 );
not \U$12074 ( \12451 , \12450 );
or \U$12075 ( \12452 , \12410 , \12451 );
or \U$12076 ( \12453 , \12450 , \12409 );
nand \U$12077 ( \12454 , \12452 , \12453 );
xor \U$12078 ( \12455 , \12403 , \12454 );
and \U$12079 ( \12456 , \12169 , \12455 );
not \U$12080 ( \12457 , \12169 );
not \U$12081 ( \12458 , \12455 );
and \U$12082 ( \12459 , \12457 , \12458 );
nor \U$12083 ( \12460 , \12456 , \12459 );
or \U$12084 ( \12461 , \11750 , \12460 );
not \U$12085 ( \12462 , \10631 );
not \U$12086 ( \12463 , \10926 );
or \U$12087 ( \12464 , \12462 , \12463 );
xnor \U$12088 ( \12465 , \10444 , RIae7a510_180);
nand \U$12089 ( \12466 , \12465 , \10927 );
nand \U$12090 ( \12467 , \12464 , \12466 );
not \U$12091 ( \12468 , \12467 );
not \U$12092 ( \12469 , \2767 );
and \U$12093 ( \12470 , RIae79c28_161, \4112 );
not \U$12094 ( \12471 , RIae79c28_161);
and \U$12095 ( \12472 , \12471 , \5911 );
or \U$12096 ( \12473 , \12470 , \12472 );
not \U$12097 ( \12474 , \12473 );
or \U$12098 ( \12475 , \12469 , \12474 );
nand \U$12099 ( \12476 , \11557 , \2776 );
nand \U$12100 ( \12477 , \12475 , \12476 );
not \U$12101 ( \12478 , \1864 );
not \U$12102 ( \12479 , \11200 );
or \U$12103 ( \12480 , \12478 , \12479 );
not \U$12104 ( \12481 , \1902 );
buf \U$12105 ( \12482 , \9606 );
not \U$12106 ( \12483 , \12482 );
not \U$12107 ( \12484 , \12483 );
not \U$12108 ( \12485 , \12484 );
or \U$12109 ( \12486 , \12481 , \12485 );
nand \U$12110 ( \12487 , \10453 , RIae793b8_143);
nand \U$12111 ( \12488 , \12486 , \12487 );
nand \U$12112 ( \12489 , \12488 , \1910 );
nand \U$12113 ( \12490 , \12480 , \12489 );
nand \U$12114 ( \12491 , \12477 , \12490 );
nand \U$12115 ( \12492 , \12468 , \12491 );
not \U$12116 ( \12493 , \12477 );
not \U$12117 ( \12494 , \12490 );
nand \U$12118 ( \12495 , \12493 , \12494 );
nand \U$12119 ( \12496 , \12492 , \12495 );
not \U$12120 ( \12497 , \2450 );
not \U$12121 ( \12498 , \11045 );
or \U$12122 ( \12499 , \12497 , \12498 );
and \U$12123 ( \12500 , RIae79778_151, \9657 );
not \U$12124 ( \12501 , RIae79778_151);
not \U$12125 ( \12502 , \9657 );
and \U$12126 ( \12503 , \12501 , \12502 );
or \U$12127 ( \12504 , \12500 , \12503 );
nand \U$12128 ( \12505 , \12504 , \9576 );
nand \U$12129 ( \12506 , \12499 , \12505 );
not \U$12130 ( \12507 , \9622 );
not \U$12131 ( \12508 , \11019 );
or \U$12132 ( \12509 , \12507 , \12508 );
not \U$12133 ( \12510 , RIae7a3a8_177);
not \U$12134 ( \12511 , \4199 );
or \U$12135 ( \12512 , \12510 , \12511 );
or \U$12136 ( \12513 , \1880 , RIae7a3a8_177);
nand \U$12137 ( \12514 , \12512 , \12513 );
buf \U$12138 ( \12515 , \11014 );
nand \U$12139 ( \12516 , \12514 , \12515 );
nand \U$12140 ( \12517 , \12509 , \12516 );
xor \U$12141 ( \12518 , \12506 , \12517 );
not \U$12142 ( \12519 , \11205 );
and \U$12143 ( \12520 , RIae7a8d0_188, \834 );
not \U$12144 ( \12521 , RIae7a8d0_188);
not \U$12145 ( \12522 , \4413 );
and \U$12146 ( \12523 , \12521 , \12522 );
or \U$12147 ( \12524 , \12520 , \12523 );
not \U$12148 ( \12525 , \12524 );
or \U$12149 ( \12526 , \12519 , \12525 );
nand \U$12150 ( \12527 , \11212 , \10275 );
nand \U$12151 ( \12528 , \12526 , \12527 );
and \U$12152 ( \12529 , \12518 , \12528 );
and \U$12153 ( \12530 , \12506 , \12517 );
or \U$12154 ( \12531 , \12529 , \12530 );
and \U$12155 ( \12532 , \12496 , \12531 );
not \U$12156 ( \12533 , \12496 );
not \U$12157 ( \12534 , \12531 );
and \U$12158 ( \12535 , \12533 , \12534 );
or \U$12159 ( \12536 , \12532 , \12535 );
not \U$12160 ( \12537 , \12536 );
and \U$12161 ( \12538 , \11075 , \10700 );
not \U$12162 ( \12539 , \2309 );
not \U$12163 ( \12540 , RIae79fe8_169);
and \U$12164 ( \12541 , \12539 , \12540 );
and \U$12165 ( \12542 , \2309 , RIae79fe8_169);
nor \U$12166 ( \12543 , \12541 , \12542 );
and \U$12167 ( \12544 , \12543 , \9499 );
nor \U$12168 ( \12545 , \12538 , \12544 );
not \U$12169 ( \12546 , \12545 );
not \U$12170 ( \12547 , \9473 );
not \U$12171 ( \12548 , \2324 );
not \U$12172 ( \12549 , \12548 );
not \U$12173 ( \12550 , RIae7a6f0_184);
and \U$12174 ( \12551 , \12549 , \12550 );
not \U$12175 ( \12552 , \1142 );
and \U$12176 ( \12553 , \12552 , RIae7a6f0_184);
nor \U$12177 ( \12554 , \12551 , \12553 );
not \U$12178 ( \12555 , \12554 );
or \U$12179 ( \12556 , \12547 , \12555 );
nand \U$12180 ( \12557 , \11126 , \9478 );
nand \U$12181 ( \12558 , \12556 , \12557 );
not \U$12182 ( \12559 , \12558 );
not \U$12183 ( \12560 , \12559 );
not \U$12184 ( \12561 , \9792 );
and \U$12185 ( \12562 , RIae7a2b8_175, \4080 );
not \U$12186 ( \12563 , RIae7a2b8_175);
not \U$12187 ( \12564 , \9501 );
and \U$12188 ( \12565 , \12563 , \12564 );
nor \U$12189 ( \12566 , \12562 , \12565 );
not \U$12190 ( \12567 , \12566 );
or \U$12191 ( \12568 , \12561 , \12567 );
nand \U$12192 ( \12569 , \11060 , \9814 );
nand \U$12193 ( \12570 , \12568 , \12569 );
not \U$12194 ( \12571 , \12570 );
or \U$12195 ( \12572 , \12560 , \12571 );
or \U$12196 ( \12573 , \12570 , \12559 );
nand \U$12197 ( \12574 , \12572 , \12573 );
not \U$12198 ( \12575 , \12574 );
or \U$12199 ( \12576 , \12546 , \12575 );
not \U$12200 ( \12577 , \12570 );
nand \U$12201 ( \12578 , \12577 , \12559 );
nand \U$12202 ( \12579 , \12576 , \12578 );
not \U$12203 ( \12580 , \12579 );
or \U$12204 ( \12581 , \12537 , \12580 );
nand \U$12205 ( \12582 , \12534 , \12496 );
nand \U$12206 ( \12583 , \12581 , \12582 );
xor \U$12207 ( \12584 , \11179 , \11219 );
xor \U$12208 ( \12585 , \11255 , \11296 );
xor \U$12209 ( \12586 , \12585 , \11345 );
nor \U$12210 ( \12587 , \12584 , \12586 );
or \U$12211 ( \12588 , \12583 , \12587 );
nand \U$12212 ( \12589 , \12584 , \12586 );
nand \U$12213 ( \12590 , \12588 , \12589 );
and \U$12214 ( \12591 , \11393 , \11381 );
not \U$12215 ( \12592 , \11393 );
not \U$12216 ( \12593 , \11381 );
and \U$12217 ( \12594 , \12592 , \12593 );
nor \U$12218 ( \12595 , \12591 , \12594 );
not \U$12219 ( \12596 , \12595 );
not \U$12220 ( \12597 , \12596 );
not \U$12221 ( \12598 , \9370 );
not \U$12222 ( \12599 , \2056 );
buf \U$12223 ( \12600 , \9394 );
not \U$12224 ( \12601 , \12600 );
or \U$12225 ( \12602 , \12599 , \12601 );
not \U$12226 ( \12603 , \12600 );
nand \U$12227 ( \12604 , \12603 , RIae79610_148);
nand \U$12228 ( \12605 , \12602 , \12604 );
not \U$12229 ( \12606 , \12605 );
or \U$12230 ( \12607 , \12598 , \12606 );
nand \U$12231 ( \12608 , \11152 , \2011 );
nand \U$12232 ( \12609 , \12607 , \12608 );
not \U$12233 ( \12610 , \12609 );
xnor \U$12234 ( \12611 , \11330 , \11325 );
not \U$12235 ( \12612 , \12611 );
not \U$12236 ( \12613 , \9320 );
buf \U$12237 ( \12614 , \9441 );
not \U$12238 ( \12615 , \12614 );
and \U$12239 ( \12616 , RIae79688_149, \12615 );
not \U$12240 ( \12617 , RIae79688_149);
and \U$12241 ( \12618 , \12617 , \9438 );
or \U$12242 ( \12619 , \12616 , \12618 );
not \U$12243 ( \12620 , \12619 );
or \U$12244 ( \12621 , \12613 , \12620 );
nand \U$12245 ( \12622 , \11158 , \1820 );
nand \U$12246 ( \12623 , \12621 , \12622 );
not \U$12247 ( \12624 , \12623 );
or \U$12248 ( \12625 , \12612 , \12624 );
or \U$12249 ( \12626 , \12611 , \12623 );
nand \U$12250 ( \12627 , \12625 , \12626 );
not \U$12251 ( \12628 , \12627 );
or \U$12252 ( \12629 , \12610 , \12628 );
not \U$12253 ( \12630 , \12611 );
nand \U$12254 ( \12631 , \12630 , \12623 );
nand \U$12255 ( \12632 , \12629 , \12631 );
not \U$12256 ( \12633 , \12632 );
not \U$12257 ( \12634 , \12633 );
or \U$12258 ( \12635 , \12597 , \12634 );
not \U$12259 ( \12636 , \12595 );
not \U$12260 ( \12637 , \12632 );
or \U$12261 ( \12638 , \12636 , \12637 );
xnor \U$12262 ( \12639 , \11292 , \11281 );
nand \U$12263 ( \12640 , \12638 , \12639 );
nand \U$12264 ( \12641 , \12635 , \12640 );
not \U$12265 ( \12642 , \12641 );
not \U$12266 ( \12643 , \1499 );
buf \U$12267 ( \12644 , \9924 );
and \U$12268 ( \12645 , \12644 , RIae79250_140);
not \U$12269 ( \12646 , \12644 );
not \U$12270 ( \12647 , RIae79250_140);
and \U$12271 ( \12648 , \12646 , \12647 );
nor \U$12272 ( \12649 , \12645 , \12648 );
not \U$12273 ( \12650 , \12649 );
or \U$12274 ( \12651 , \12643 , \12650 );
nand \U$12275 ( \12652 , \11189 , \1501 );
nand \U$12276 ( \12653 , \12651 , \12652 );
not \U$12277 ( \12654 , \12653 );
not \U$12278 ( \12655 , \1062 );
not \U$12279 ( \12656 , \1039 );
not \U$12280 ( \12657 , \9868 );
or \U$12281 ( \12658 , \12656 , \12657 );
nand \U$12282 ( \12659 , \10749 , RIae79070_136);
nand \U$12283 ( \12660 , \12658 , \12659 );
not \U$12284 ( \12661 , \12660 );
or \U$12285 ( \12662 , \12655 , \12661 );
nand \U$12286 ( \12663 , \11274 , \1049 );
nand \U$12287 ( \12664 , \12662 , \12663 );
not \U$12288 ( \12665 , \797 );
and \U$12289 ( \12666 , \10740 , \1132 );
not \U$12290 ( \12667 , \10740 );
and \U$12291 ( \12668 , \12667 , RIae78f80_134);
nor \U$12292 ( \12669 , \12666 , \12668 );
not \U$12293 ( \12670 , \12669 );
or \U$12294 ( \12671 , \12665 , \12670 );
nand \U$12295 ( \12672 , \11264 , \838 );
nand \U$12296 ( \12673 , \12671 , \12672 );
nor \U$12297 ( \12674 , \12664 , \12673 );
not \U$12298 ( \12675 , \12674 );
not \U$12299 ( \12676 , \12675 );
or \U$12300 ( \12677 , \12654 , \12676 );
nand \U$12301 ( \12678 , \12664 , \12673 );
nand \U$12302 ( \12679 , \12677 , \12678 );
buf \U$12303 ( \12680 , \2188 );
not \U$12304 ( \12681 , \12680 );
not \U$12305 ( \12682 , RIae79520_146);
not \U$12306 ( \12683 , \9298 );
buf \U$12307 ( \12684 , \12683 );
not \U$12308 ( \12685 , \12684 );
or \U$12309 ( \12686 , \12682 , \12685 );
not \U$12310 ( \12687 , \9298 );
or \U$12311 ( \12688 , \12687 , RIae79520_146);
nand \U$12312 ( \12689 , \12686 , \12688 );
not \U$12313 ( \12690 , \12689 );
or \U$12314 ( \12691 , \12681 , \12690 );
nand \U$12315 ( \12692 , \11336 , \2163 );
nand \U$12316 ( \12693 , \12691 , \12692 );
not \U$12317 ( \12694 , \2467 );
not \U$12318 ( \12695 , \11290 );
or \U$12319 ( \12696 , \12694 , \12695 );
not \U$12320 ( \12697 , \3039 );
not \U$12321 ( \12698 , \9280 );
or \U$12322 ( \12699 , \12697 , \12698 );
not \U$12323 ( \12700 , \5722 );
nand \U$12324 ( \12701 , \12700 , RIae794a8_145);
nand \U$12325 ( \12702 , \12699 , \12701 );
nand \U$12326 ( \12703 , \12702 , \9828 );
nand \U$12327 ( \12704 , \12696 , \12703 );
xor \U$12328 ( \12705 , \12693 , \12704 );
not \U$12329 ( \12706 , \2272 );
buf \U$12330 ( \12707 , \9347 );
and \U$12331 ( \12708 , RIae79ac0_158, \12707 );
not \U$12332 ( \12709 , RIae79ac0_158);
not \U$12333 ( \12710 , \12707 );
and \U$12334 ( \12711 , \12709 , \12710 );
or \U$12335 ( \12712 , \12708 , \12711 );
not \U$12336 ( \12713 , \12712 );
or \U$12337 ( \12714 , \12706 , \12713 );
nand \U$12338 ( \12715 , \11172 , \2252 );
nand \U$12339 ( \12716 , \12714 , \12715 );
and \U$12340 ( \12717 , \12705 , \12716 );
and \U$12341 ( \12718 , \12693 , \12704 );
or \U$12342 ( \12719 , \12717 , \12718 );
xor \U$12343 ( \12720 , \12679 , \12719 );
not \U$12344 ( \12721 , \2340 );
and \U$12345 ( \12722 , RIae798e0_154, \10226 );
not \U$12346 ( \12723 , RIae798e0_154);
not \U$12347 ( \12724 , \4960 );
and \U$12348 ( \12725 , \12723 , \12724 );
or \U$12349 ( \12726 , \12722 , \12725 );
not \U$12350 ( \12727 , \12726 );
or \U$12351 ( \12728 , \12721 , \12727 );
nand \U$12352 ( \12729 , \11304 , \2322 );
nand \U$12353 ( \12730 , \12728 , \12729 );
not \U$12354 ( \12731 , \1989 );
not \U$12355 ( \12732 , RIae797f0_152);
not \U$12356 ( \12733 , \5860 );
or \U$12357 ( \12734 , \12732 , \12733 );
nand \U$12358 ( \12735 , \4982 , \2521 );
nand \U$12359 ( \12736 , \12734 , \12735 );
not \U$12360 ( \12737 , \12736 );
or \U$12361 ( \12738 , \12731 , \12737 );
nand \U$12362 ( \12739 , \11030 , \2519 );
nand \U$12363 ( \12740 , \12738 , \12739 );
xor \U$12364 ( \12741 , \12730 , \12740 );
not \U$12365 ( \12742 , \867 );
not \U$12366 ( \12743 , \11313 );
or \U$12367 ( \12744 , \12742 , \12743 );
xor \U$12368 ( \12745 , RIae78b48_125, \10845 );
nand \U$12369 ( \12746 , \12745 , \892 );
nand \U$12370 ( \12747 , \12744 , \12746 );
xor \U$12371 ( \12748 , RIae774c8_77, RIae77540_78);
xor \U$12372 ( \12749 , \10243 , \12748 );
buf \U$12373 ( \12750 , \12749 );
not \U$12374 ( \12751 , \12750 );
nand \U$12375 ( \12752 , \12751 , RIae78b48_125);
xor \U$12376 ( \12753 , \12747 , \12752 );
not \U$12377 ( \12754 , \12753 );
not \U$12378 ( \12755 , \1072 );
not \U$12379 ( \12756 , \11591 );
or \U$12380 ( \12757 , \12755 , \12756 );
not \U$12381 ( \12758 , \10042 );
not \U$12382 ( \12759 , \1066 );
or \U$12383 ( \12760 , \12758 , \12759 );
or \U$12384 ( \12761 , \10042 , \921 );
nand \U$12385 ( \12762 , \12760 , \12761 );
nand \U$12386 ( \12763 , \1086 , \12762 );
nand \U$12387 ( \12764 , \12757 , \12763 );
nand \U$12388 ( \12765 , \12754 , \12764 );
not \U$12389 ( \12766 , \12752 );
nand \U$12390 ( \12767 , \12766 , \12747 );
and \U$12391 ( \12768 , \12765 , \12767 );
not \U$12392 ( \12769 , \12768 );
and \U$12393 ( \12770 , \12741 , \12769 );
and \U$12394 ( \12771 , \12730 , \12740 );
or \U$12395 ( \12772 , \12770 , \12771 );
and \U$12396 ( \12773 , \12720 , \12772 );
and \U$12397 ( \12774 , \12679 , \12719 );
or \U$12398 ( \12775 , \12773 , \12774 );
xor \U$12399 ( \12776 , \12642 , \12775 );
xor \U$12400 ( \12777 , \11154 , \11174 );
xor \U$12401 ( \12778 , \12777 , \11160 );
not \U$12402 ( \12779 , \10573 );
not \U$12403 ( \12780 , \11415 );
or \U$12404 ( \12781 , \12779 , \12780 );
not \U$12405 ( \12782 , \4023 );
not \U$12406 ( \12783 , RIae79ef8_167);
and \U$12407 ( \12784 , \12782 , \12783 );
and \U$12408 ( \12785 , \2858 , RIae79ef8_167);
nor \U$12409 ( \12786 , \12784 , \12785 );
nand \U$12410 ( \12787 , \12786 , \6201 );
nand \U$12411 ( \12788 , \12781 , \12787 );
not \U$12412 ( \12789 , \6091 );
and \U$12413 ( \12790 , RIae79d90_164, \3524 );
not \U$12414 ( \12791 , RIae79d90_164);
and \U$12415 ( \12792 , \12791 , \10884 );
or \U$12416 ( \12793 , \12790 , \12792 );
not \U$12417 ( \12794 , \12793 );
or \U$12418 ( \12795 , \12789 , \12794 );
nand \U$12419 ( \12796 , \10910 , \5049 );
nand \U$12420 ( \12797 , \12795 , \12796 );
xor \U$12421 ( \12798 , \12788 , \12797 );
not \U$12422 ( \12799 , \10667 );
not \U$12423 ( \12800 , \1117 );
not \U$12424 ( \12801 , \12800 );
and \U$12425 ( \12802 , RIae7a150_172, \12801 );
not \U$12426 ( \12803 , RIae7a150_172);
and \U$12427 ( \12804 , \12803 , \12800 );
nor \U$12428 ( \12805 , \12802 , \12804 );
not \U$12429 ( \12806 , \12805 );
or \U$12430 ( \12807 , \12799 , \12806 );
nand \U$12431 ( \12808 , \11086 , \9777 );
nand \U$12432 ( \12809 , \12807 , \12808 );
and \U$12433 ( \12810 , \12798 , \12809 );
and \U$12434 ( \12811 , \12788 , \12797 );
or \U$12435 ( \12812 , \12810 , \12811 );
xor \U$12436 ( \12813 , \12778 , \12812 );
xor \U$12437 ( \12814 , \11191 , \11202 );
xor \U$12438 ( \12815 , \12814 , \11216 );
and \U$12439 ( \12816 , \12813 , \12815 );
and \U$12440 ( \12817 , \12778 , \12812 );
or \U$12441 ( \12818 , \12816 , \12817 );
and \U$12442 ( \12819 , \12776 , \12818 );
and \U$12443 ( \12820 , \12642 , \12775 );
or \U$12444 ( \12821 , \12819 , \12820 );
xor \U$12445 ( \12822 , \12590 , \12821 );
buf \U$12446 ( \12823 , \10985 );
not \U$12447 ( \12824 , \12823 );
not \U$12448 ( \12825 , \10933 );
not \U$12449 ( \12826 , \12825 );
and \U$12450 ( \12827 , \12824 , \12826 );
and \U$12451 ( \12828 , \12823 , \12825 );
nor \U$12452 ( \12829 , \12827 , \12828 );
not \U$12453 ( \12830 , \12829 );
not \U$12454 ( \12831 , \12830 );
xor \U$12455 ( \12832 , \11032 , \11023 );
xnor \U$12456 ( \12833 , \12832 , \11047 );
xor \U$12457 ( \12834 , \11121 , \11109 );
xor \U$12458 ( \12835 , \12834 , \11133 );
xor \U$12459 ( \12836 , \12833 , \12835 );
not \U$12460 ( \12837 , \926 );
not \U$12461 ( \12838 , RIae78bc0_126);
not \U$12462 ( \12839 , \12838 );
not \U$12463 ( \12840 , \11321 );
or \U$12464 ( \12841 , \12839 , \12840 );
buf \U$12465 ( \12842 , \11317 );
not \U$12466 ( \12843 , RIae78bc0_126);
or \U$12467 ( \12844 , \12842 , \12843 );
nand \U$12468 ( \12845 , \12841 , \12844 );
not \U$12469 ( \12846 , \12845 );
or \U$12470 ( \12847 , \12837 , \12846 );
not \U$12471 ( \12848 , RIae78bc0_126);
not \U$12472 ( \12849 , \10259 );
or \U$12473 ( \12850 , \12848 , \12849 );
or \U$12474 ( \12851 , \10259 , RIae78bc0_126);
nand \U$12475 ( \12852 , \12850 , \12851 );
nand \U$12476 ( \12853 , \12852 , \949 );
nand \U$12477 ( \12854 , \12847 , \12853 );
not \U$12478 ( \12855 , \12854 );
xor \U$12479 ( \12856 , RIae775b8_79, RIae77630_80);
buf \U$12480 ( \12857 , \12856 );
buf \U$12481 ( \12858 , \12857 );
and \U$12482 ( \12859 , RIae78b48_125, \12858 );
not \U$12483 ( \12860 , \867 );
not \U$12484 ( \12861 , \12745 );
or \U$12485 ( \12862 , \12860 , \12861 );
nand \U$12486 ( \12863 , \12750 , \860 );
nand \U$12487 ( \12864 , \12752 , \12863 , \892 );
nand \U$12488 ( \12865 , \12862 , \12864 );
xor \U$12489 ( \12866 , \12859 , \12865 );
not \U$12490 ( \12867 , \12866 );
or \U$12491 ( \12868 , \12855 , \12867 );
nand \U$12492 ( \12869 , \12865 , \12859 );
nand \U$12493 ( \12870 , \12868 , \12869 );
not \U$12494 ( \12871 , \926 );
not \U$12495 ( \12872 , \11583 );
or \U$12496 ( \12873 , \12871 , \12872 );
nand \U$12497 ( \12874 , \12845 , \951 );
nand \U$12498 ( \12875 , \12873 , \12874 );
not \U$12499 ( \12876 , \12875 );
and \U$12500 ( \12877 , \12870 , \12876 );
not \U$12501 ( \12878 , \12870 );
and \U$12502 ( \12879 , \12878 , \12875 );
nor \U$12503 ( \12880 , \12877 , \12879 );
not \U$12504 ( \12881 , \12880 );
not \U$12505 ( \12882 , \12881 );
not \U$12506 ( \12883 , \1501 );
not \U$12507 ( \12884 , \12649 );
or \U$12508 ( \12885 , \12883 , \12884 );
not \U$12509 ( \12886 , RIae79250_140);
not \U$12510 ( \12887 , \10084 );
or \U$12511 ( \12888 , \12886 , \12887 );
or \U$12512 ( \12889 , \10084 , RIae79250_140);
nand \U$12513 ( \12890 , \12888 , \12889 );
nand \U$12514 ( \12891 , \12890 , \9403 );
nand \U$12515 ( \12892 , \12885 , \12891 );
not \U$12516 ( \12893 , \12892 );
or \U$12517 ( \12894 , \12882 , \12893 );
not \U$12518 ( \12895 , \12876 );
nand \U$12519 ( \12896 , \12895 , \12870 );
nand \U$12520 ( \12897 , \12894 , \12896 );
not \U$12521 ( \12898 , \10696 );
xor \U$12522 ( \12899 , RIae7a498_179, \1826 );
not \U$12523 ( \12900 , \12899 );
or \U$12524 ( \12901 , \12898 , \12900 );
nand \U$12525 ( \12902 , \11433 , \10677 );
nand \U$12526 ( \12903 , \12901 , \12902 );
xor \U$12527 ( \12904 , \12897 , \12903 );
nand \U$12528 ( \12905 , \10894 , \4853 );
and \U$12529 ( \12906 , RIae79ca0_162, \2564 );
not \U$12530 ( \12907 , RIae79ca0_162);
and \U$12531 ( \12908 , \12907 , \4837 );
or \U$12532 ( \12909 , \12906 , \12908 );
nand \U$12533 ( \12910 , \12909 , \11761 );
and \U$12534 ( \12911 , \12905 , \12910 );
not \U$12535 ( \12912 , \12911 );
and \U$12536 ( \12913 , \12904 , \12912 );
and \U$12537 ( \12914 , \12897 , \12903 );
nor \U$12538 ( \12915 , \12913 , \12914 );
and \U$12539 ( \12916 , \12836 , \12915 );
and \U$12540 ( \12917 , \12833 , \12835 );
or \U$12541 ( \12918 , \12916 , \12917 );
not \U$12542 ( \12919 , \12918 );
not \U$12543 ( \12920 , \12919 );
or \U$12544 ( \12921 , \12831 , \12920 );
not \U$12545 ( \12922 , \12829 );
not \U$12546 ( \12923 , \12918 );
or \U$12547 ( \12924 , \12922 , \12923 );
xor \U$12548 ( \12925 , \10912 , \10896 );
xnor \U$12549 ( \12926 , \12925 , \10929 );
not \U$12550 ( \12927 , \11452 );
not \U$12551 ( \12928 , \11419 );
not \U$12552 ( \12929 , \12928 );
and \U$12553 ( \12930 , \12927 , \12929 );
and \U$12554 ( \12931 , \11452 , \12928 );
nor \U$12555 ( \12932 , \12930 , \12931 );
xor \U$12556 ( \12933 , \12926 , \12932 );
not \U$12557 ( \12934 , \11089 );
not \U$12558 ( \12935 , \11093 );
or \U$12559 ( \12936 , \12934 , \12935 );
nand \U$12560 ( \12937 , \11090 , \11077 );
nand \U$12561 ( \12938 , \12936 , \12937 );
and \U$12562 ( \12939 , \12938 , \11092 );
not \U$12563 ( \12940 , \12938 );
not \U$12564 ( \12941 , \11092 );
and \U$12565 ( \12942 , \12940 , \12941 );
nor \U$12566 ( \12943 , \12939 , \12942 );
and \U$12567 ( \12944 , \12933 , \12943 );
and \U$12568 ( \12945 , \12926 , \12932 );
or \U$12569 ( \12946 , \12944 , \12945 );
not \U$12570 ( \12947 , \12946 );
nand \U$12571 ( \12948 , \12924 , \12947 );
nand \U$12572 ( \12949 , \12921 , \12948 );
and \U$12573 ( \12950 , \12822 , \12949 );
and \U$12574 ( \12951 , \12590 , \12821 );
or \U$12575 ( \12952 , \12950 , \12951 );
not \U$12576 ( \12953 , \11010 );
not \U$12577 ( \12954 , \11354 );
or \U$12578 ( \12955 , \12953 , \12954 );
nand \U$12579 ( \12956 , \11353 , \11011 );
nand \U$12580 ( \12957 , \12955 , \12956 );
not \U$12581 ( \12958 , \12957 );
not \U$12582 ( \12959 , \11475 );
and \U$12583 ( \12960 , \12958 , \12959 );
and \U$12584 ( \12961 , \12957 , \11475 );
nor \U$12585 ( \12962 , \12960 , \12961 );
xor \U$12586 ( \12963 , \12952 , \12962 );
xor \U$12587 ( \12964 , \11483 , \11649 );
xor \U$12588 ( \12965 , \12964 , \11740 );
and \U$12589 ( \12966 , \12963 , \12965 );
and \U$12590 ( \12967 , \12952 , \12962 );
or \U$12591 ( \12968 , \12966 , \12967 );
nand \U$12592 ( \12969 , \12461 , \12968 );
nand \U$12593 ( \12970 , \12460 , \11750 );
nand \U$12594 ( \12971 , \12969 , \12970 );
not \U$12595 ( \12972 , \12971 );
not \U$12596 ( \12973 , \12454 );
not \U$12597 ( \12974 , \12403 );
or \U$12598 ( \12975 , \12973 , \12974 );
not \U$12599 ( \12976 , \12450 );
nand \U$12600 ( \12977 , \12976 , \12409 );
nand \U$12601 ( \12978 , \12975 , \12977 );
not \U$12602 ( \12979 , \12978 );
not \U$12603 ( \12980 , \12153 );
not \U$12604 ( \12981 , \12980 );
xnor \U$12605 ( \12982 , \12040 , \12161 );
not \U$12606 ( \12983 , \12982 );
or \U$12607 ( \12984 , \12981 , \12983 );
nand \U$12608 ( \12985 , \12160 , \12040 );
nand \U$12609 ( \12986 , \12984 , \12985 );
not \U$12610 ( \12987 , \12986 );
not \U$12611 ( \12988 , \12987 );
or \U$12612 ( \12989 , \12979 , \12988 );
not \U$12613 ( \12990 , \12978 );
nand \U$12614 ( \12991 , \12990 , \12986 );
nand \U$12615 ( \12992 , \12989 , \12991 );
not \U$12616 ( \12993 , \9828 );
not \U$12617 ( \12994 , \12175 );
or \U$12618 ( \12995 , \12993 , \12994 );
not \U$12619 ( \12996 , \1968 );
not \U$12620 ( \12997 , \12996 );
and \U$12621 ( \12998 , \12997 , \3810 );
not \U$12622 ( \12999 , \12997 );
and \U$12623 ( \13000 , \12999 , RIae794a8_145);
nor \U$12624 ( \13001 , \12998 , \13000 );
nand \U$12625 ( \13002 , \13001 , \2467 );
nand \U$12626 ( \13003 , \12995 , \13002 );
not \U$12627 ( \13004 , \2340 );
not \U$12628 ( \13005 , \12196 );
or \U$12629 ( \13006 , \13004 , \13005 );
not \U$12630 ( \13007 , RIae798e0_154);
not \U$12631 ( \13008 , \2093 );
not \U$12632 ( \13009 , \13008 );
or \U$12633 ( \13010 , \13007 , \13009 );
or \U$12634 ( \13011 , \2785 , RIae798e0_154);
nand \U$12635 ( \13012 , \13010 , \13011 );
nand \U$12636 ( \13013 , \13012 , \2322 );
nand \U$12637 ( \13014 , \13006 , \13013 );
xor \U$12638 ( \13015 , \13003 , \13014 );
not \U$12639 ( \13016 , \9814 );
and \U$12640 ( \13017 , RIae7a2b8_175, \1834 );
not \U$12641 ( \13018 , RIae7a2b8_175);
and \U$12642 ( \13019 , \13018 , \6148 );
or \U$12643 ( \13020 , \13017 , \13019 );
not \U$12644 ( \13021 , \13020 );
or \U$12645 ( \13022 , \13016 , \13021 );
nand \U$12646 ( \13023 , \12188 , \9792 );
nand \U$12647 ( \13024 , \13022 , \13023 );
xnor \U$12648 ( \13025 , \13015 , \13024 );
not \U$12649 ( \13026 , \10709 );
not \U$12650 ( \13027 , \12366 );
or \U$12651 ( \13028 , \13026 , \13027 );
not \U$12652 ( \13029 , RIae79fe8_169);
not \U$12653 ( \13030 , \2593 );
or \U$12654 ( \13031 , \13029 , \13030 );
not \U$12655 ( \13032 , \2047 );
not \U$12656 ( \13033 , \13032 );
or \U$12657 ( \13034 , \13033 , RIae79fe8_169);
nand \U$12658 ( \13035 , \13031 , \13034 );
nand \U$12659 ( \13036 , \13035 , \9517 );
nand \U$12660 ( \13037 , \13028 , \13036 );
not \U$12661 ( \13038 , RIae7a498_179);
not \U$12662 ( \13039 , \1158 );
or \U$12663 ( \13040 , \13038 , \13039 );
or \U$12664 ( \13041 , \3326 , RIae7a498_179);
nand \U$12665 ( \13042 , \13040 , \13041 );
and \U$12666 ( \13043 , \13042 , \10677 );
and \U$12667 ( \13044 , \12377 , \11434 );
nor \U$12668 ( \13045 , \13043 , \13044 );
not \U$12669 ( \13046 , \13045 );
xor \U$12670 ( \13047 , \13037 , \13046 );
not \U$12671 ( \13048 , \10542 );
xor \U$12672 ( \13049 , RIae7a060_170, \11858 );
not \U$12673 ( \13050 , \13049 );
or \U$12674 ( \13051 , \13048 , \13050 );
nand \U$12675 ( \13052 , \12389 , \9730 );
nand \U$12676 ( \13053 , \13051 , \13052 );
xnor \U$12677 ( \13054 , \13047 , \13053 );
xor \U$12678 ( \13055 , \13025 , \13054 );
not \U$12679 ( \13056 , \5040 );
not \U$12680 ( \13057 , \12222 );
or \U$12681 ( \13058 , \13056 , \13057 );
not \U$12682 ( \13059 , RIae79d90_164);
not \U$12683 ( \13060 , \13059 );
not \U$12684 ( \13061 , \2230 );
not \U$12685 ( \13062 , \13061 );
or \U$12686 ( \13063 , \13060 , \13062 );
nand \U$12687 ( \13064 , \2230 , RIae79d90_164);
nand \U$12688 ( \13065 , \13063 , \13064 );
nand \U$12689 ( \13066 , \13065 , \6080 );
nand \U$12690 ( \13067 , \13058 , \13066 );
not \U$12691 ( \13068 , \10638 );
not \U$12692 ( \13069 , \12238 );
or \U$12693 ( \13070 , \13068 , \13069 );
and \U$12694 ( \13071 , RIae7a510_180, \938 );
not \U$12695 ( \13072 , RIae7a510_180);
and \U$12696 ( \13073 , \13072 , \939 );
or \U$12697 ( \13074 , \13071 , \13073 );
nand \U$12698 ( \13075 , \13074 , \10631 );
nand \U$12699 ( \13076 , \13070 , \13075 );
and \U$12700 ( \13077 , \13067 , \13076 );
not \U$12701 ( \13078 , \13067 );
not \U$12702 ( \13079 , \13076 );
and \U$12703 ( \13080 , \13078 , \13079 );
nor \U$12704 ( \13081 , \13077 , \13080 );
not \U$12705 ( \13082 , \11409 );
not \U$12706 ( \13083 , \12211 );
or \U$12707 ( \13084 , \13082 , \13083 );
not \U$12708 ( \13085 , \6203 );
not \U$12709 ( \13086 , \1897 );
not \U$12710 ( \13087 , \13086 );
not \U$12711 ( \13088 , \13087 );
or \U$12712 ( \13089 , \13085 , \13088 );
or \U$12713 ( \13090 , \1899 , \9560 );
nand \U$12714 ( \13091 , \13089 , \13090 );
nand \U$12715 ( \13092 , \13091 , \6214 );
nand \U$12716 ( \13093 , \13084 , \13092 );
not \U$12717 ( \13094 , \13093 );
and \U$12718 ( \13095 , \13081 , \13094 );
not \U$12719 ( \13096 , \13081 );
and \U$12720 ( \13097 , \13096 , \13093 );
nor \U$12721 ( \13098 , \13095 , \13097 );
xor \U$12722 ( \13099 , \13055 , \13098 );
not \U$12723 ( \13100 , \13099 );
not \U$12724 ( \13101 , \2433 );
not \U$12725 ( \13102 , \12305 );
or \U$12726 ( \13103 , \13101 , \13102 );
and \U$12727 ( \13104 , RIae79778_151, \1760 );
not \U$12728 ( \13105 , RIae79778_151);
and \U$12729 ( \13106 , \13105 , \10605 );
or \U$12730 ( \13107 , \13104 , \13106 );
nand \U$12731 ( \13108 , \13107 , \2450 );
nand \U$12732 ( \13109 , \13103 , \13108 );
not \U$12733 ( \13110 , \2776 );
not \U$12734 ( \13111 , RIae79c28_161);
not \U$12735 ( \13112 , \2287 );
or \U$12736 ( \13113 , \13111 , \13112 );
or \U$12737 ( \13114 , \10534 , RIae79c28_161);
nand \U$12738 ( \13115 , \13113 , \13114 );
not \U$12739 ( \13116 , \13115 );
or \U$12740 ( \13117 , \13110 , \13116 );
nand \U$12741 ( \13118 , \12294 , \2767 );
nand \U$12742 ( \13119 , \13117 , \13118 );
xor \U$12743 ( \13120 , \13109 , \13119 );
buf \U$12744 ( \13121 , \9699 );
not \U$12745 ( \13122 , \13121 );
not \U$12746 ( \13123 , RIae7a240_174);
not \U$12747 ( \13124 , \977 );
or \U$12748 ( \13125 , \13123 , \13124 );
nand \U$12749 ( \13126 , \5082 , \9679 );
nand \U$12750 ( \13127 , \13125 , \13126 );
not \U$12751 ( \13128 , \13127 );
or \U$12752 ( \13129 , \13122 , \13128 );
buf \U$12753 ( \13130 , \9688 );
nand \U$12754 ( \13131 , \12314 , \13130 );
nand \U$12755 ( \13132 , \13129 , \13131 );
xor \U$12756 ( \13133 , \13120 , \13132 );
not \U$12757 ( \13134 , \12245 );
not \U$12758 ( \13135 , \12227 );
or \U$12759 ( \13136 , \13134 , \13135 );
nand \U$12760 ( \13137 , \13136 , \12215 );
nand \U$12761 ( \13138 , \12226 , \12242 );
nand \U$12762 ( \13139 , \13137 , \13138 );
xor \U$12763 ( \13140 , \13133 , \13139 );
not \U$12764 ( \13141 , \4853 );
not \U$12765 ( \13142 , \5631 );
and \U$12766 ( \13143 , RIae79ca0_162, \13142 );
not \U$12767 ( \13144 , RIae79ca0_162);
and \U$12768 ( \13145 , \13144 , \2955 );
or \U$12769 ( \13146 , \13143 , \13145 );
not \U$12770 ( \13147 , \13146 );
or \U$12771 ( \13148 , \13141 , \13147 );
nand \U$12772 ( \13149 , \12254 , \6276 );
nand \U$12773 ( \13150 , \13148 , \13149 );
not \U$12774 ( \13151 , \9777 );
and \U$12775 ( \13152 , \10658 , \780 );
not \U$12776 ( \13153 , \10658 );
and \U$12777 ( \13154 , \13153 , \781 );
nor \U$12778 ( \13155 , \13152 , \13154 );
not \U$12779 ( \13156 , \13155 );
or \U$12780 ( \13157 , \13151 , \13156 );
buf \U$12781 ( \13158 , \9758 );
nand \U$12782 ( \13159 , \12264 , \13158 );
nand \U$12783 ( \13160 , \13157 , \13159 );
xor \U$12784 ( \13161 , \13150 , \13160 );
not \U$12785 ( \13162 , \12515 );
not \U$12786 ( \13163 , \12272 );
or \U$12787 ( \13164 , \13162 , \13163 );
not \U$12788 ( \13165 , RIae7a3a8_177);
not \U$12789 ( \13166 , \13165 );
not \U$12790 ( \13167 , \5351 );
or \U$12791 ( \13168 , \13166 , \13167 );
nand \U$12792 ( \13169 , \2175 , RIae7a3a8_177);
nand \U$12793 ( \13170 , \13168 , \13169 );
nand \U$12794 ( \13171 , \13170 , \9621 );
nand \U$12795 ( \13172 , \13164 , \13171 );
xnor \U$12796 ( \13173 , \13161 , \13172 );
xnor \U$12797 ( \13174 , \13140 , \13173 );
not \U$12798 ( \13175 , \13174 );
or \U$12799 ( \13176 , \13100 , \13175 );
or \U$12800 ( \13177 , \13174 , \13099 );
nand \U$12801 ( \13178 , \13176 , \13177 );
not \U$12802 ( \13179 , \10309 );
not \U$12803 ( \13180 , \10130 );
or \U$12804 ( \13181 , \13179 , \13180 );
not \U$12805 ( \13182 , \10119 );
nand \U$12806 ( \13183 , \13182 , \10126 );
nand \U$12807 ( \13184 , \13181 , \13183 );
not \U$12808 ( \13185 , \13184 );
and \U$12809 ( \13186 , \13178 , \13185 );
not \U$12810 ( \13187 , \13178 );
and \U$12811 ( \13188 , \13187 , \13184 );
nor \U$12812 ( \13189 , \13186 , \13188 );
not \U$12813 ( \13190 , \13189 );
not \U$12814 ( \13191 , \12279 );
not \U$12815 ( \13192 , \13191 );
not \U$12816 ( \13193 , \12398 );
or \U$12817 ( \13194 , \13192 , \13193 );
not \U$12818 ( \13195 , \12398 );
not \U$12819 ( \13196 , \13195 );
not \U$12820 ( \13197 , \12279 );
or \U$12821 ( \13198 , \13196 , \13197 );
not \U$12822 ( \13199 , \12287 );
nand \U$12823 ( \13200 , \13198 , \13199 );
nand \U$12824 ( \13201 , \13194 , \13200 );
not \U$12825 ( \13202 , \13201 );
nand \U$12826 ( \13203 , \13190 , \13202 );
nand \U$12827 ( \13204 , \13189 , \13201 );
nand \U$12828 ( \13205 , \13203 , \13204 );
not \U$12829 ( \13206 , \12298 );
not \U$12830 ( \13207 , \12326 );
not \U$12831 ( \13208 , \13207 );
not \U$12832 ( \13209 , \13208 );
or \U$12833 ( \13210 , \13206 , \13209 );
nand \U$12834 ( \13211 , \12317 , \12307 );
nand \U$12835 ( \13212 , \13210 , \13211 );
xor \U$12836 ( \13213 , \12258 , \12270 );
and \U$12837 ( \13214 , \13213 , \12277 );
and \U$12838 ( \13215 , \12258 , \12270 );
or \U$12839 ( \13216 , \13214 , \13215 );
not \U$12840 ( \13217 , \13216 );
not \U$12841 ( \13218 , \12370 );
and \U$12842 ( \13219 , \12391 , \12381 );
not \U$12843 ( \13220 , \12391 );
not \U$12844 ( \13221 , \12381 );
and \U$12845 ( \13222 , \13220 , \13221 );
nor \U$12846 ( \13223 , \13219 , \13222 );
not \U$12847 ( \13224 , \13223 );
or \U$12848 ( \13225 , \13218 , \13224 );
nand \U$12849 ( \13226 , \12391 , \12381 );
nand \U$12850 ( \13227 , \13225 , \13226 );
not \U$12851 ( \13228 , \13227 );
not \U$12852 ( \13229 , \13228 );
or \U$12853 ( \13230 , \13217 , \13229 );
or \U$12854 ( \13231 , \13228 , \13216 );
nand \U$12855 ( \13232 , \13230 , \13231 );
xor \U$12856 ( \13233 , \13212 , \13232 );
not \U$12857 ( \13234 , \12392 );
not \U$12858 ( \13235 , \12360 );
or \U$12859 ( \13236 , \13234 , \13235 );
not \U$12860 ( \13237 , \12298 );
nand \U$12861 ( \13238 , \13237 , \12326 );
not \U$12862 ( \13239 , \13238 );
nand \U$12863 ( \13240 , \13207 , \12298 );
not \U$12864 ( \13241 , \13240 );
or \U$12865 ( \13242 , \13239 , \13241 );
not \U$12866 ( \13243 , \12359 );
nand \U$12867 ( \13244 , \13242 , \13243 );
nand \U$12868 ( \13245 , \13236 , \13244 );
not \U$12869 ( \13246 , \13245 );
not \U$12870 ( \13247 , \1820 );
not \U$12871 ( \13248 , \5107 );
xnor \U$12872 ( \13249 , RIae79688_149, \13248 );
not \U$12873 ( \13250 , \13249 );
or \U$12874 ( \13251 , \13247 , \13250 );
nand \U$12875 ( \13252 , \12338 , \10401 );
nand \U$12876 ( \13253 , \13251 , \13252 );
not \U$12877 ( \13254 , \2063 );
not \U$12878 ( \13255 , \12060 );
or \U$12879 ( \13256 , \13254 , \13255 );
not \U$12880 ( \13257 , \9286 );
xor \U$12881 ( \13258 , RIae79610_148, \13257 );
nand \U$12882 ( \13259 , \13258 , \2011 );
nand \U$12883 ( \13260 , \13256 , \13259 );
not \U$12884 ( \13261 , \13260 );
and \U$12885 ( \13262 , \13253 , \13261 );
not \U$12886 ( \13263 , \13253 );
and \U$12887 ( \13264 , \13263 , \13260 );
nor \U$12888 ( \13265 , \13262 , \13264 );
not \U$12889 ( \13266 , \1910 );
not \U$12890 ( \13267 , \12068 );
or \U$12891 ( \13268 , \13266 , \13267 );
and \U$12892 ( \13269 , \9317 , RIae793b8_143);
not \U$12893 ( \13270 , \9317 );
and \U$12894 ( \13271 , \13270 , \1884 );
nor \U$12895 ( \13272 , \13269 , \13271 );
nand \U$12896 ( \13273 , \13272 , \1863 );
nand \U$12897 ( \13274 , \13268 , \13273 );
not \U$12898 ( \13275 , \13274 );
and \U$12899 ( \13276 , \13265 , \13275 );
not \U$12900 ( \13277 , \13265 );
and \U$12901 ( \13278 , \13277 , \13274 );
nor \U$12902 ( \13279 , \13276 , \13278 );
not \U$12903 ( \13280 , \1062 );
not \U$12904 ( \13281 , \12081 );
or \U$12905 ( \13282 , \13280 , \13281 );
xor \U$12906 ( \13283 , \9416 , RIae79070_136);
nand \U$12907 ( \13284 , \13283 , \9947 );
nand \U$12908 ( \13285 , \13282 , \13284 );
not \U$12909 ( \13286 , \1501 );
not \U$12910 ( \13287 , \9367 );
and \U$12911 ( \13288 , RIae79250_140, \13287 );
not \U$12912 ( \13289 , RIae79250_140);
buf \U$12913 ( \13290 , \9367 );
and \U$12914 ( \13291 , \13289 , \13290 );
or \U$12915 ( \13292 , \13288 , \13291 );
not \U$12916 ( \13293 , \13292 );
or \U$12917 ( \13294 , \13286 , \13293 );
nand \U$12918 ( \13295 , \12049 , \1499 );
nand \U$12919 ( \13296 , \13294 , \13295 );
xor \U$12920 ( \13297 , \13285 , \13296 );
not \U$12921 ( \13298 , \2157 );
not \U$12922 ( \13299 , \12089 );
or \U$12923 ( \13300 , \13298 , \13299 );
not \U$12924 ( \13301 , \9455 );
buf \U$12925 ( \13302 , \13301 );
and \U$12926 ( \13303 , RIae79160_138, \13302 );
not \U$12927 ( \13304 , RIae79160_138);
and \U$12928 ( \13305 , \13304 , \9459 );
or \U$12929 ( \13306 , \13303 , \13305 );
nand \U$12930 ( \13307 , \13306 , \1209 );
nand \U$12931 ( \13308 , \13300 , \13307 );
xnor \U$12932 ( \13309 , \13297 , \13308 );
not \U$12933 ( \13310 , \13309 );
xor \U$12934 ( \13311 , \13279 , \13310 );
not \U$12935 ( \13312 , \2272 );
not \U$12936 ( \13313 , \12354 );
or \U$12937 ( \13314 , \13312 , \13313 );
not \U$12938 ( \13315 , RIae79ac0_158);
not \U$12939 ( \13316 , \6242 );
or \U$12940 ( \13317 , \13315 , \13316 );
or \U$12941 ( \13318 , \6242 , RIae79ac0_158);
nand \U$12942 ( \13319 , \13317 , \13318 );
nand \U$12943 ( \13320 , \13319 , \10414 );
nand \U$12944 ( \13321 , \13314 , \13320 );
not \U$12945 ( \13322 , \10339 );
not \U$12946 ( \13323 , \13322 );
not \U$12947 ( \13324 , \12680 );
not \U$12948 ( \13325 , \10333 );
or \U$12949 ( \13326 , \13324 , \13325 );
and \U$12950 ( \13327 , RIae79520_146, \5673 );
not \U$12951 ( \13328 , RIae79520_146);
and \U$12952 ( \13329 , \13328 , \10492 );
nor \U$12953 ( \13330 , \13327 , \13329 );
nand \U$12954 ( \13331 , \13330 , \3440 );
nand \U$12955 ( \13332 , \13326 , \13331 );
not \U$12956 ( \13333 , \13332 );
not \U$12957 ( \13334 , \13333 );
or \U$12958 ( \13335 , \13323 , \13334 );
nand \U$12959 ( \13336 , \13332 , \10339 );
nand \U$12960 ( \13337 , \13335 , \13336 );
xor \U$12961 ( \13338 , \13321 , \13337 );
buf \U$12962 ( \13339 , \13338 );
xnor \U$12963 ( \13340 , \13311 , \13339 );
not \U$12964 ( \13341 , \13340 );
or \U$12965 ( \13342 , \13246 , \13341 );
or \U$12966 ( \13343 , \13245 , \13340 );
nand \U$12967 ( \13344 , \13342 , \13343 );
buf \U$12968 ( \13345 , \13344 );
xor \U$12969 ( \13346 , \13233 , \13345 );
not \U$12970 ( \13347 , \13346 );
and \U$12971 ( \13348 , \13205 , \13347 );
not \U$12972 ( \13349 , \13205 );
and \U$12973 ( \13350 , \13349 , \13346 );
nor \U$12974 ( \13351 , \13348 , \13350 );
and \U$12975 ( \13352 , \12992 , \13351 );
not \U$12976 ( \13353 , \12992 );
not \U$12977 ( \13354 , \13351 );
and \U$12978 ( \13355 , \13353 , \13354 );
nor \U$12979 ( \13356 , \13352 , \13355 );
not \U$12980 ( \13357 , \13356 );
or \U$12981 ( \13358 , \12455 , \12033 );
nand \U$12982 ( \13359 , \13358 , \12167 );
nand \U$12983 ( \13360 , \12033 , \12455 );
nand \U$12984 ( \13361 , \13359 , \13360 );
not \U$12985 ( \13362 , \13361 );
not \U$12986 ( \13363 , \13362 );
not \U$12987 ( \13364 , \10721 );
not \U$12988 ( \13365 , \11478 );
or \U$12989 ( \13366 , \13364 , \13365 );
not \U$12990 ( \13367 , \10720 );
not \U$12991 ( \13368 , \11479 );
or \U$12992 ( \13369 , \13367 , \13368 );
nand \U$12993 ( \13370 , \13369 , \11743 );
nand \U$12994 ( \13371 , \13366 , \13370 );
not \U$12995 ( \13372 , \13371 );
not \U$12996 ( \13373 , \9974 );
and \U$12997 ( \13374 , \10314 , \13373 );
or \U$12998 ( \13375 , \13374 , \10719 );
or \U$12999 ( \13376 , \13373 , \10314 );
nand \U$13000 ( \13377 , \13375 , \13376 );
not \U$13001 ( \13378 , \13377 );
not \U$13002 ( \13379 , \12144 );
not \U$13003 ( \13380 , \13379 );
not \U$13004 ( \13381 , \12101 );
or \U$13005 ( \13382 , \13380 , \13381 );
or \U$13006 ( \13383 , \12101 , \13379 );
nand \U$13007 ( \13384 , \13383 , \12152 );
nand \U$13008 ( \13385 , \13382 , \13384 );
not \U$13009 ( \13386 , \13385 );
not \U$13010 ( \13387 , \10528 );
not \U$13011 ( \13388 , \10717 );
or \U$13012 ( \13389 , \13387 , \13388 );
or \U$13013 ( \13390 , \10717 , \10528 );
not \U$13014 ( \13391 , \10439 );
nand \U$13015 ( \13392 , \13390 , \13391 );
nand \U$13016 ( \13393 , \13389 , \13392 );
not \U$13017 ( \13394 , \13393 );
not \U$13018 ( \13395 , \2007 );
and \U$13019 ( \13396 , RIae797f0_152, \1789 );
not \U$13020 ( \13397 , RIae797f0_152);
not \U$13021 ( \13398 , \1789 );
and \U$13022 ( \13399 , \13397 , \13398 );
or \U$13023 ( \13400 , \13396 , \13399 );
not \U$13024 ( \13401 , \13400 );
or \U$13025 ( \13402 , \13395 , \13401 );
nand \U$13026 ( \13403 , \10101 , \1988 );
nand \U$13027 ( \13404 , \13402 , \13403 );
not \U$13028 ( \13405 , \12123 );
not \U$13029 ( \13406 , \13405 );
not \U$13030 ( \13407 , \12130 );
or \U$13031 ( \13408 , \13406 , \13407 );
nand \U$13032 ( \13409 , \13408 , \12117 );
nand \U$13033 ( \13410 , \12129 , \12123 );
nand \U$13034 ( \13411 , \13409 , \13410 );
not \U$13035 ( \13412 , RIae7a768_185);
not \U$13036 ( \13413 , RIae7a6f0_184);
or \U$13037 ( \13414 , \13412 , \13413 );
nand \U$13038 ( \13415 , \13414 , RIae7a7e0_186);
not \U$13039 ( \13416 , \13415 );
nand \U$13040 ( \13417 , \10142 , RIae78b48_125);
not \U$13041 ( \13418 , \13417 );
or \U$13042 ( \13419 , \13416 , \13418 );
not \U$13043 ( \13420 , \13415 );
nand \U$13044 ( \13421 , \13420 , \10142 , RIae78b48_125);
nand \U$13045 ( \13422 , \13419 , \13421 );
not \U$13046 ( \13423 , \13422 );
not \U$13047 ( \13424 , \1072 );
not \U$13048 ( \13425 , \921 );
not \U$13049 ( \13426 , \11386 );
or \U$13050 ( \13427 , \13425 , \13426 );
nand \U$13051 ( \13428 , \10084 , RIae78e90_132);
nand \U$13052 ( \13429 , \13427 , \13428 );
not \U$13053 ( \13430 , \13429 );
or \U$13054 ( \13431 , \13424 , \13430 );
nand \U$13055 ( \13432 , \12125 , \1086 );
nand \U$13056 ( \13433 , \13431 , \13432 );
not \U$13057 ( \13434 , \13433 );
not \U$13058 ( \13435 , \13434 );
or \U$13059 ( \13436 , \13423 , \13435 );
or \U$13060 ( \13437 , \13434 , \13422 );
nand \U$13061 ( \13438 , \13436 , \13437 );
xor \U$13062 ( \13439 , \13411 , \13438 );
xor \U$13063 ( \13440 , \13404 , \13439 );
not \U$13064 ( \13441 , \13440 );
not \U$13065 ( \13442 , \13441 );
not \U$13066 ( \13443 , \10118 );
or \U$13067 ( \13444 , \13443 , \10113 );
not \U$13068 ( \13445 , \10109 );
or \U$13069 ( \13446 , \13445 , \10094 );
nand \U$13070 ( \13447 , \13444 , \13446 );
not \U$13071 ( \13448 , \13447 );
or \U$13072 ( \13449 , \13442 , \13448 );
or \U$13073 ( \13450 , \13447 , \13441 );
nand \U$13074 ( \13451 , \13449 , \13450 );
not \U$13075 ( \13452 , \13451 );
not \U$13076 ( \13453 , \10356 );
not \U$13077 ( \13454 , \10395 );
or \U$13078 ( \13455 , \13453 , \13454 );
not \U$13079 ( \13456 , \10355 );
not \U$13080 ( \13457 , \10396 );
or \U$13081 ( \13458 , \13456 , \13457 );
nand \U$13082 ( \13459 , \13458 , \10434 );
nand \U$13083 ( \13460 , \13455 , \13459 );
not \U$13084 ( \13461 , \13460 );
not \U$13085 ( \13462 , \13461 );
and \U$13086 ( \13463 , \13452 , \13462 );
and \U$13087 ( \13464 , \13451 , \13461 );
nor \U$13088 ( \13465 , \13463 , \13464 );
not \U$13089 ( \13466 , \13465 );
or \U$13090 ( \13467 , \13394 , \13466 );
or \U$13091 ( \13468 , \13393 , \13465 );
nand \U$13092 ( \13469 , \13467 , \13468 );
not \U$13093 ( \13470 , \13469 );
or \U$13094 ( \13471 , \13386 , \13470 );
or \U$13095 ( \13472 , \13385 , \13469 );
nand \U$13096 ( \13473 , \13471 , \13472 );
not \U$13097 ( \13474 , \13473 );
or \U$13098 ( \13475 , \13378 , \13474 );
or \U$13099 ( \13476 , \13473 , \13377 );
nand \U$13100 ( \13477 , \13475 , \13476 );
not \U$13101 ( \13478 , \13477 );
or \U$13102 ( \13479 , \12247 , \12201 );
nand \U$13103 ( \13480 , \13479 , \12278 );
nand \U$13104 ( \13481 , \12247 , \12201 );
nand \U$13105 ( \13482 , \13480 , \13481 );
not \U$13106 ( \13483 , \12107 );
not \U$13107 ( \13484 , \12143 );
or \U$13108 ( \13485 , \13483 , \13484 );
not \U$13109 ( \13486 , \12141 );
nand \U$13110 ( \13487 , \13486 , \12132 );
nand \U$13111 ( \13488 , \13485 , \13487 );
not \U$13112 ( \13489 , \13488 );
nand \U$13113 ( \13490 , \12435 , \12427 );
nand \U$13114 ( \13491 , \12435 , \12419 );
nand \U$13115 ( \13492 , \12427 , \12419 );
and \U$13116 ( \13493 , \13490 , \13491 , \13492 );
not \U$13117 ( \13494 , \13493 );
or \U$13118 ( \13495 , \13489 , \13494 );
or \U$13119 ( \13496 , \13493 , \13488 );
nand \U$13120 ( \13497 , \13495 , \13496 );
xor \U$13121 ( \13498 , \13482 , \13497 );
not \U$13122 ( \13499 , \13498 );
or \U$13123 ( \13500 , \12072 , \12053 );
nand \U$13124 ( \13501 , \13500 , \12064 );
nand \U$13125 ( \13502 , \12072 , \12053 );
nand \U$13126 ( \13503 , \13501 , \13502 );
not \U$13127 ( \13504 , \10350 );
not \U$13128 ( \13505 , \10335 );
or \U$13129 ( \13506 , \13504 , \13505 );
nand \U$13130 ( \13507 , \10349 , \10339 );
nand \U$13131 ( \13508 , \13506 , \13507 );
xor \U$13132 ( \13509 , \13503 , \13508 );
not \U$13133 ( \13510 , \12358 );
not \U$13134 ( \13511 , \12351 );
or \U$13135 ( \13512 , \13510 , \13511 );
not \U$13136 ( \13513 , \12344 );
not \U$13137 ( \13514 , \12346 );
or \U$13138 ( \13515 , \13513 , \13514 );
nand \U$13139 ( \13516 , \13515 , \12332 );
nand \U$13140 ( \13517 , \13512 , \13516 );
xor \U$13141 ( \13518 , \13509 , \13517 );
not \U$13142 ( \13519 , \13518 );
not \U$13143 ( \13520 , \12100 );
not \U$13144 ( \13521 , \12044 );
nand \U$13145 ( \13522 , \13521 , \12073 );
not \U$13146 ( \13523 , \13522 );
or \U$13147 ( \13524 , \13520 , \13523 );
nand \U$13148 ( \13525 , \12074 , \12044 );
nand \U$13149 ( \13526 , \13524 , \13525 );
not \U$13150 ( \13527 , \13526 );
not \U$13151 ( \13528 , \13527 );
or \U$13152 ( \13529 , \13519 , \13528 );
not \U$13153 ( \13530 , \13518 );
nand \U$13154 ( \13531 , \13530 , \13526 );
nand \U$13155 ( \13532 , \13529 , \13531 );
not \U$13156 ( \13533 , \867 );
xor \U$13157 ( \13534 , RIae78b48_125, \10007 );
not \U$13158 ( \13535 , \13534 );
or \U$13159 ( \13536 , \13533 , \13535 );
nand \U$13160 ( \13537 , \12119 , \892 );
nand \U$13161 ( \13538 , \13536 , \13537 );
not \U$13162 ( \13539 , \951 );
not \U$13163 ( \13540 , \10345 );
or \U$13164 ( \13541 , \13539 , \13540 );
and \U$13165 ( \13542 , \1286 , \9897 );
not \U$13166 ( \13543 , \1286 );
not \U$13167 ( \13544 , \10168 );
and \U$13168 ( \13545 , \13543 , \13544 );
nor \U$13169 ( \13546 , \13542 , \13545 );
nand \U$13170 ( \13547 , \13546 , \926 );
nand \U$13171 ( \13548 , \13541 , \13547 );
xor \U$13172 ( \13549 , \13538 , \13548 );
not \U$13173 ( \13550 , \796 );
xnor \U$13174 ( \13551 , RIae78f80_134, \10724 );
not \U$13175 ( \13552 , \13551 );
or \U$13176 ( \13553 , \13550 , \13552 );
and \U$13177 ( \13554 , RIae78f80_134, \10465 );
not \U$13178 ( \13555 , RIae78f80_134);
and \U$13179 ( \13556 , \13555 , \10461 );
nor \U$13180 ( \13557 , \13554 , \13556 );
nand \U$13181 ( \13558 , \13557 , \838 );
nand \U$13182 ( \13559 , \13553 , \13558 );
xor \U$13183 ( \13560 , \13549 , \13559 );
xor \U$13184 ( \13561 , \12179 , \12190 );
not \U$13185 ( \13562 , \13561 );
not \U$13186 ( \13563 , \12200 );
or \U$13187 ( \13564 , \13562 , \13563 );
nand \U$13188 ( \13565 , \12190 , \12179 );
nand \U$13189 ( \13566 , \13564 , \13565 );
xor \U$13190 ( \13567 , \13560 , \13566 );
not \U$13191 ( \13568 , \12093 );
not \U$13192 ( \13569 , \12086 );
not \U$13193 ( \13570 , \12099 );
or \U$13194 ( \13571 , \13569 , \13570 );
or \U$13195 ( \13572 , \12099 , \12086 );
nand \U$13196 ( \13573 , \13571 , \13572 );
not \U$13197 ( \13574 , \13573 );
or \U$13198 ( \13575 , \13568 , \13574 );
nand \U$13199 ( \13576 , \12099 , \12085 );
nand \U$13200 ( \13577 , \13575 , \13576 );
xor \U$13201 ( \13578 , \13567 , \13577 );
xnor \U$13202 ( \13579 , \13532 , \13578 );
not \U$13203 ( \13580 , \13579 );
or \U$13204 ( \13581 , \13499 , \13580 );
or \U$13205 ( \13582 , \13498 , \13579 );
nand \U$13206 ( \13583 , \13581 , \13582 );
not \U$13207 ( \13584 , \12445 );
not \U$13208 ( \13585 , \12440 );
or \U$13209 ( \13586 , \13584 , \13585 );
not \U$13210 ( \13587 , \12436 );
nand \U$13211 ( \13588 , \13587 , \12414 );
nand \U$13212 ( \13589 , \13586 , \13588 );
not \U$13213 ( \13590 , \13589 );
and \U$13214 ( \13591 , \13583 , \13590 );
not \U$13215 ( \13592 , \13583 );
and \U$13216 ( \13593 , \13592 , \13589 );
nor \U$13217 ( \13594 , \13591 , \13593 );
not \U$13218 ( \13595 , \13594 );
or \U$13219 ( \13596 , \13478 , \13595 );
or \U$13220 ( \13597 , \13594 , \13477 );
nand \U$13221 ( \13598 , \13596 , \13597 );
not \U$13222 ( \13599 , \13598 );
not \U$13223 ( \13600 , \13599 );
or \U$13224 ( \13601 , \13372 , \13600 );
not \U$13225 ( \13602 , \13371 );
nand \U$13226 ( \13603 , \13602 , \13598 );
nand \U$13227 ( \13604 , \13601 , \13603 );
not \U$13228 ( \13605 , \13604 );
and \U$13229 ( \13606 , \13363 , \13605 );
and \U$13230 ( \13607 , \13362 , \13604 );
nor \U$13231 ( \13608 , \13606 , \13607 );
not \U$13232 ( \13609 , \13608 );
or \U$13233 ( \13610 , \13357 , \13609 );
or \U$13234 ( \13611 , \13608 , \13356 );
nand \U$13235 ( \13612 , \13610 , \13611 );
not \U$13236 ( \13613 , \13612 );
or \U$13237 ( \13614 , \12972 , \13613 );
not \U$13238 ( \13615 , \13608 );
nand \U$13239 ( \13616 , \13615 , \13356 );
nand \U$13240 ( \13617 , \13614 , \13616 );
not \U$13241 ( \13618 , \13351 );
not \U$13242 ( \13619 , \12992 );
or \U$13243 ( \13620 , \13618 , \13619 );
nand \U$13244 ( \13621 , \12986 , \12978 );
nand \U$13245 ( \13622 , \13620 , \13621 );
buf \U$13246 ( \13623 , \13377 );
not \U$13247 ( \13624 , \13623 );
buf \U$13248 ( \13625 , \13473 );
nand \U$13249 ( \13626 , \13624 , \13625 );
not \U$13250 ( \13627 , \13626 );
not \U$13251 ( \13628 , \13594 );
not \U$13252 ( \13629 , \13628 );
or \U$13253 ( \13630 , \13627 , \13629 );
not \U$13254 ( \13631 , \13625 );
nand \U$13255 ( \13632 , \13631 , \13623 );
nand \U$13256 ( \13633 , \13630 , \13632 );
buf \U$13257 ( \13634 , \13385 );
not \U$13258 ( \13635 , \13465 );
or \U$13259 ( \13636 , \13634 , \13635 );
buf \U$13260 ( \13637 , \13393 );
nand \U$13261 ( \13638 , \13636 , \13637 );
nand \U$13262 ( \13639 , \13634 , \13635 );
nand \U$13263 ( \13640 , \13638 , \13639 );
not \U$13264 ( \13641 , \13233 );
not \U$13265 ( \13642 , \13344 );
or \U$13266 ( \13643 , \13641 , \13642 );
not \U$13267 ( \13644 , \13340 );
buf \U$13268 ( \13645 , \13245 );
nand \U$13269 ( \13646 , \13644 , \13645 );
nand \U$13270 ( \13647 , \13643 , \13646 );
not \U$13271 ( \13648 , \13647 );
not \U$13272 ( \13649 , \13578 );
not \U$13273 ( \13650 , \13532 );
or \U$13274 ( \13651 , \13649 , \13650 );
buf \U$13275 ( \13652 , \13526 );
nand \U$13276 ( \13653 , \13652 , \13518 );
nand \U$13277 ( \13654 , \13651 , \13653 );
not \U$13278 ( \13655 , \1320 );
not \U$13279 ( \13656 , RIae78e90_132);
not \U$13280 ( \13657 , \12644 );
not \U$13281 ( \13658 , \13657 );
or \U$13282 ( \13659 , \13656 , \13658 );
buf \U$13283 ( \13660 , \9925 );
not \U$13284 ( \13661 , \13660 );
nand \U$13285 ( \13662 , \13661 , \921 );
nand \U$13286 ( \13663 , \13659 , \13662 );
not \U$13287 ( \13664 , \13663 );
or \U$13288 ( \13665 , \13655 , \13664 );
nand \U$13289 ( \13666 , \13429 , \1086 );
nand \U$13290 ( \13667 , \13665 , \13666 );
not \U$13291 ( \13668 , \2450 );
and \U$13292 ( \13669 , RIae79778_151, \3098 );
not \U$13293 ( \13670 , RIae79778_151);
not \U$13294 ( \13671 , \3098 );
and \U$13295 ( \13672 , \13670 , \13671 );
or \U$13296 ( \13673 , \13669 , \13672 );
not \U$13297 ( \13674 , \13673 );
or \U$13298 ( \13675 , \13668 , \13674 );
nand \U$13299 ( \13676 , \13107 , \2432 );
nand \U$13300 ( \13677 , \13675 , \13676 );
xor \U$13301 ( \13678 , \13667 , \13677 );
not \U$13302 ( \13679 , \1989 );
not \U$13303 ( \13680 , \13400 );
or \U$13304 ( \13681 , \13679 , \13680 );
and \U$13305 ( \13682 , RIae797f0_152, \2697 );
not \U$13306 ( \13683 , RIae797f0_152);
and \U$13307 ( \13684 , \13683 , \3529 );
or \U$13308 ( \13685 , \13682 , \13684 );
nand \U$13309 ( \13686 , \13685 , \2007 );
nand \U$13310 ( \13687 , \13681 , \13686 );
xnor \U$13311 ( \13688 , \13678 , \13687 );
not \U$13312 ( \13689 , \10677 );
not \U$13313 ( \13690 , RIae7a498_179);
not \U$13314 ( \13691 , \2324 );
or \U$13315 ( \13692 , \13690 , \13691 );
or \U$13316 ( \13693 , \1146 , RIae7a498_179);
nand \U$13317 ( \13694 , \13692 , \13693 );
not \U$13318 ( \13695 , \13694 );
or \U$13319 ( \13696 , \13689 , \13695 );
nand \U$13320 ( \13697 , \13042 , \11434 );
nand \U$13321 ( \13698 , \13696 , \13697 );
not \U$13322 ( \13699 , \2767 );
not \U$13323 ( \13700 , \13115 );
or \U$13324 ( \13701 , \13699 , \13700 );
not \U$13325 ( \13702 , \10584 );
not \U$13326 ( \13703 , \2309 );
or \U$13327 ( \13704 , \13702 , \13703 );
or \U$13328 ( \13705 , \2309 , \10584 );
nand \U$13329 ( \13706 , \13704 , \13705 );
nand \U$13330 ( \13707 , \13706 , \11364 );
nand \U$13331 ( \13708 , \13701 , \13707 );
nor \U$13332 ( \13709 , \13698 , \13708 );
not \U$13333 ( \13710 , \13709 );
nand \U$13334 ( \13711 , \13698 , \13708 );
nand \U$13335 ( \13712 , \13710 , \13711 );
not \U$13336 ( \13713 , \9699 );
and \U$13337 ( \13714 , RIae7a240_174, \1119 );
not \U$13338 ( \13715 , RIae7a240_174);
and \U$13339 ( \13716 , \13715 , \2917 );
or \U$13340 ( \13717 , \13714 , \13716 );
not \U$13341 ( \13718 , \13717 );
or \U$13342 ( \13719 , \13713 , \13718 );
buf \U$13343 ( \13720 , \9687 );
nand \U$13344 ( \13721 , \13127 , \13720 );
nand \U$13345 ( \13722 , \13719 , \13721 );
and \U$13346 ( \13723 , \13712 , \13722 );
not \U$13347 ( \13724 , \13712 );
not \U$13348 ( \13725 , \13722 );
and \U$13349 ( \13726 , \13724 , \13725 );
nor \U$13350 ( \13727 , \13723 , \13726 );
xor \U$13351 ( \13728 , \13688 , \13727 );
not \U$13352 ( \13729 , \6214 );
not \U$13353 ( \13730 , \6207 );
not \U$13354 ( \13731 , \1879 );
or \U$13355 ( \13732 , \13730 , \13731 );
not \U$13356 ( \13733 , RIae79ef8_167);
or \U$13357 ( \13734 , \1879 , \13733 );
nand \U$13358 ( \13735 , \13732 , \13734 );
not \U$13359 ( \13736 , \13735 );
or \U$13360 ( \13737 , \13729 , \13736 );
nand \U$13361 ( \13738 , \11409 , \13091 );
nand \U$13362 ( \13739 , \13737 , \13738 );
not \U$13363 ( \13740 , \10631 );
not \U$13364 ( \13741 , RIae7a510_180);
not \U$13365 ( \13742 , \1438 );
or \U$13366 ( \13743 , \13741 , \13742 );
or \U$13367 ( \13744 , \10662 , RIae7a510_180);
nand \U$13368 ( \13745 , \13743 , \13744 );
not \U$13369 ( \13746 , \13745 );
or \U$13370 ( \13747 , \13740 , \13746 );
nand \U$13371 ( \13748 , \13074 , \10638 );
nand \U$13372 ( \13749 , \13747 , \13748 );
xor \U$13373 ( \13750 , \13739 , \13749 );
not \U$13374 ( \13751 , \9777 );
and \U$13375 ( \13752 , RIae7a150_172, \12522 );
not \U$13376 ( \13753 , RIae7a150_172);
and \U$13377 ( \13754 , \13753 , \834 );
nor \U$13378 ( \13755 , \13752 , \13754 );
not \U$13379 ( \13756 , \13755 );
or \U$13380 ( \13757 , \13751 , \13756 );
nand \U$13381 ( \13758 , \13155 , \10667 );
nand \U$13382 ( \13759 , \13757 , \13758 );
xor \U$13383 ( \13760 , \13750 , \13759 );
xor \U$13384 ( \13761 , \13728 , \13760 );
xor \U$13385 ( \13762 , \13654 , \13761 );
not \U$13386 ( \13763 , \13762 );
or \U$13387 ( \13764 , \13648 , \13763 );
not \U$13388 ( \13765 , \13647 );
nand \U$13389 ( \13766 , \13532 , \13578 );
and \U$13390 ( \13767 , \13766 , \13653 );
and \U$13391 ( \13768 , \13767 , \13761 );
not \U$13392 ( \13769 , \13767 );
not \U$13393 ( \13770 , \13761 );
and \U$13394 ( \13771 , \13769 , \13770 );
nor \U$13395 ( \13772 , \13768 , \13771 );
nand \U$13396 ( \13773 , \13765 , \13772 );
nand \U$13397 ( \13774 , \13764 , \13773 );
xor \U$13398 ( \13775 , \13640 , \13774 );
not \U$13399 ( \13776 , \13589 );
not \U$13400 ( \13777 , \13583 );
or \U$13401 ( \13778 , \13776 , \13777 );
not \U$13402 ( \13779 , \13579 );
nand \U$13403 ( \13780 , \13779 , \13498 );
nand \U$13404 ( \13781 , \13778 , \13780 );
xor \U$13405 ( \13782 , \13775 , \13781 );
xor \U$13406 ( \13783 , \13633 , \13782 );
xor \U$13407 ( \13784 , \13622 , \13783 );
not \U$13408 ( \13785 , \13784 );
not \U$13409 ( \13786 , \13785 );
not \U$13410 ( \13787 , \13204 );
not \U$13411 ( \13788 , \13346 );
or \U$13412 ( \13789 , \13787 , \13788 );
nand \U$13413 ( \13790 , \13789 , \13203 );
not \U$13414 ( \13791 , \13482 );
not \U$13415 ( \13792 , \13497 );
or \U$13416 ( \13793 , \13791 , \13792 );
not \U$13417 ( \13794 , \13493 );
nand \U$13418 ( \13795 , \13794 , \13488 );
nand \U$13419 ( \13796 , \13793 , \13795 );
not \U$13420 ( \13797 , \13796 );
not \U$13421 ( \13798 , \13797 );
xnor \U$13422 ( \13799 , \13309 , \13338 );
not \U$13423 ( \13800 , \13799 );
not \U$13424 ( \13801 , \13279 );
or \U$13425 ( \13802 , \13800 , \13801 );
nand \U$13426 ( \13803 , \13339 , \13310 );
nand \U$13427 ( \13804 , \13802 , \13803 );
xor \U$13428 ( \13805 , \13560 , \13566 );
and \U$13429 ( \13806 , \13805 , \13577 );
and \U$13430 ( \13807 , \13560 , \13566 );
or \U$13431 ( \13808 , \13806 , \13807 );
and \U$13432 ( \13809 , \13804 , \13808 );
not \U$13433 ( \13810 , \13804 );
not \U$13434 ( \13811 , \13808 );
and \U$13435 ( \13812 , \13810 , \13811 );
nor \U$13436 ( \13813 , \13809 , \13812 );
not \U$13437 ( \13814 , \13003 );
not \U$13438 ( \13815 , \13024 );
or \U$13439 ( \13816 , \13814 , \13815 );
or \U$13440 ( \13817 , \13024 , \13003 );
nand \U$13441 ( \13818 , \13817 , \13014 );
nand \U$13442 ( \13819 , \13816 , \13818 );
not \U$13443 ( \13820 , \13037 );
not \U$13444 ( \13821 , \13045 );
not \U$13445 ( \13822 , \13053 );
or \U$13446 ( \13823 , \13821 , \13822 );
or \U$13447 ( \13824 , \13053 , \13045 );
nand \U$13448 ( \13825 , \13823 , \13824 );
not \U$13449 ( \13826 , \13825 );
or \U$13450 ( \13827 , \13820 , \13826 );
nand \U$13451 ( \13828 , \13053 , \13046 );
nand \U$13452 ( \13829 , \13827 , \13828 );
and \U$13453 ( \13830 , \13819 , \13829 );
not \U$13454 ( \13831 , \13819 );
not \U$13455 ( \13832 , \13829 );
and \U$13456 ( \13833 , \13831 , \13832 );
nor \U$13457 ( \13834 , \13830 , \13833 );
not \U$13458 ( \13835 , \13093 );
not \U$13459 ( \13836 , \13081 );
or \U$13460 ( \13837 , \13835 , \13836 );
nand \U$13461 ( \13838 , \13076 , \13067 );
nand \U$13462 ( \13839 , \13837 , \13838 );
not \U$13463 ( \13840 , \13839 );
and \U$13464 ( \13841 , \13834 , \13840 );
not \U$13465 ( \13842 , \13834 );
and \U$13466 ( \13843 , \13842 , \13839 );
nor \U$13467 ( \13844 , \13841 , \13843 );
and \U$13468 ( \13845 , \13813 , \13844 );
not \U$13469 ( \13846 , \13813 );
not \U$13470 ( \13847 , \13844 );
and \U$13471 ( \13848 , \13846 , \13847 );
nor \U$13472 ( \13849 , \13845 , \13848 );
not \U$13473 ( \13850 , \13849 );
not \U$13474 ( \13851 , \13850 );
not \U$13475 ( \13852 , \13851 );
or \U$13476 ( \13853 , \13798 , \13852 );
nand \U$13477 ( \13854 , \13850 , \13796 );
nand \U$13478 ( \13855 , \13853 , \13854 );
not \U$13479 ( \13856 , \13212 );
not \U$13480 ( \13857 , \13232 );
or \U$13481 ( \13858 , \13856 , \13857 );
nand \U$13482 ( \13859 , \13227 , \13216 );
nand \U$13483 ( \13860 , \13858 , \13859 );
not \U$13484 ( \13861 , \13860 );
or \U$13485 ( \13862 , \13274 , \13260 );
nand \U$13486 ( \13863 , \13862 , \13253 );
nand \U$13487 ( \13864 , \13274 , \13260 );
nand \U$13488 ( \13865 , \13863 , \13864 );
not \U$13489 ( \13866 , \13422 );
not \U$13490 ( \13867 , \13433 );
or \U$13491 ( \13868 , \13866 , \13867 );
not \U$13492 ( \13869 , \13417 );
nand \U$13493 ( \13870 , \13869 , \13415 );
nand \U$13494 ( \13871 , \13868 , \13870 );
xor \U$13495 ( \13872 , \13865 , \13871 );
buf \U$13496 ( \13873 , \13872 );
not \U$13497 ( \13874 , \13321 );
not \U$13498 ( \13875 , \13337 );
or \U$13499 ( \13876 , \13874 , \13875 );
nand \U$13500 ( \13877 , \13332 , \13322 );
nand \U$13501 ( \13878 , \13876 , \13877 );
not \U$13502 ( \13879 , \13878 );
and \U$13503 ( \13880 , \13873 , \13879 );
not \U$13504 ( \13881 , \13873 );
and \U$13505 ( \13882 , \13881 , \13878 );
nor \U$13506 ( \13883 , \13880 , \13882 );
not \U$13507 ( \13884 , \13883 );
nor \U$13508 ( \13885 , \13172 , \13160 );
not \U$13509 ( \13886 , \13150 );
or \U$13510 ( \13887 , \13885 , \13886 );
nand \U$13511 ( \13888 , \13172 , \13160 );
nand \U$13512 ( \13889 , \13887 , \13888 );
not \U$13513 ( \13890 , \13889 );
and \U$13514 ( \13891 , RIae78b48_125, \10743 );
not \U$13515 ( \13892 , \867 );
not \U$13516 ( \13893 , \860 );
not \U$13517 ( \13894 , \9868 );
or \U$13518 ( \13895 , \13893 , \13894 );
buf \U$13519 ( \13896 , \10749 );
nand \U$13520 ( \13897 , \13896 , RIae78b48_125);
nand \U$13521 ( \13898 , \13895 , \13897 );
not \U$13522 ( \13899 , \13898 );
or \U$13523 ( \13900 , \13892 , \13899 );
nand \U$13524 ( \13901 , \13534 , \1129 );
nand \U$13525 ( \13902 , \13900 , \13901 );
xor \U$13526 ( \13903 , \13891 , \13902 );
not \U$13527 ( \13904 , \927 );
not \U$13528 ( \13905 , \11230 );
xor \U$13529 ( \13906 , \13905 , RIae78bc0_126);
not \U$13530 ( \13907 , \13906 );
or \U$13531 ( \13908 , \13904 , \13907 );
nand \U$13532 ( \13909 , \951 , \13546 );
nand \U$13533 ( \13910 , \13908 , \13909 );
xor \U$13534 ( \13911 , \13903 , \13910 );
and \U$13535 ( \13912 , \13297 , \13308 );
and \U$13536 ( \13913 , \13285 , \13296 );
nor \U$13537 ( \13914 , \13912 , \13913 );
xor \U$13538 ( \13915 , \13911 , \13914 );
not \U$13539 ( \13916 , \13915 );
or \U$13540 ( \13917 , \13890 , \13916 );
or \U$13541 ( \13918 , \13889 , \13915 );
nand \U$13542 ( \13919 , \13917 , \13918 );
not \U$13543 ( \13920 , \13919 );
and \U$13544 ( \13921 , \13884 , \13920 );
and \U$13545 ( \13922 , \13919 , \13883 );
nor \U$13546 ( \13923 , \13921 , \13922 );
not \U$13547 ( \13924 , \13923 );
or \U$13548 ( \13925 , \13861 , \13924 );
or \U$13549 ( \13926 , \13860 , \13923 );
nand \U$13550 ( \13927 , \13925 , \13926 );
buf \U$13551 ( \13928 , \13927 );
not \U$13552 ( \13929 , \13928 );
and \U$13553 ( \13930 , \13855 , \13929 );
not \U$13554 ( \13931 , \13855 );
and \U$13555 ( \13932 , \13931 , \13928 );
nor \U$13556 ( \13933 , \13930 , \13932 );
xor \U$13557 ( \13934 , \13790 , \13933 );
xor \U$13558 ( \13935 , \13538 , \13548 );
and \U$13559 ( \13936 , \13935 , \13559 );
and \U$13560 ( \13937 , \13538 , \13548 );
or \U$13561 ( \13938 , \13936 , \13937 );
not \U$13562 ( \13939 , \2322 );
and \U$13563 ( \13940 , RIae798e0_154, \6413 );
not \U$13564 ( \13941 , RIae798e0_154);
not \U$13565 ( \13942 , \11512 );
and \U$13566 ( \13943 , \13941 , \13942 );
nor \U$13567 ( \13944 , \13940 , \13943 );
not \U$13568 ( \13945 , \13944 );
or \U$13569 ( \13946 , \13939 , \13945 );
nand \U$13570 ( \13947 , \13012 , \10807 );
nand \U$13571 ( \13948 , \13946 , \13947 );
xor \U$13572 ( \13949 , \13938 , \13948 );
not \U$13573 ( \13950 , \9815 );
not \U$13574 ( \13951 , RIae7a2b8_175);
not \U$13575 ( \13952 , \1186 );
or \U$13576 ( \13953 , \13951 , \13952 );
or \U$13577 ( \13954 , \1186 , RIae7a2b8_175);
nand \U$13578 ( \13955 , \13953 , \13954 );
not \U$13579 ( \13956 , \13955 );
or \U$13580 ( \13957 , \13950 , \13956 );
nand \U$13581 ( \13958 , \13020 , \9792 );
nand \U$13582 ( \13959 , \13957 , \13958 );
xor \U$13583 ( \13960 , \13949 , \13959 );
not \U$13584 ( \13961 , \13960 );
not \U$13585 ( \13962 , \13404 );
not \U$13586 ( \13963 , \13439 );
or \U$13587 ( \13964 , \13962 , \13963 );
not \U$13588 ( \13965 , \13410 );
not \U$13589 ( \13966 , \13409 );
or \U$13590 ( \13967 , \13965 , \13966 );
nand \U$13591 ( \13968 , \13967 , \13438 );
nand \U$13592 ( \13969 , \13964 , \13968 );
not \U$13593 ( \13970 , \2063 );
not \U$13594 ( \13971 , \13258 );
or \U$13595 ( \13972 , \13970 , \13971 );
not \U$13596 ( \13973 , \6674 );
not \U$13597 ( \13974 , \5722 );
or \U$13598 ( \13975 , \13973 , \13974 );
not \U$13599 ( \13976 , \5722 );
nand \U$13600 ( \13977 , \13976 , RIae79610_148);
nand \U$13601 ( \13978 , \13975 , \13977 );
nand \U$13602 ( \13979 , \13978 , \2011 );
nand \U$13603 ( \13980 , \13972 , \13979 );
not \U$13604 ( \13981 , \1820 );
not \U$13605 ( \13982 , RIae79688_149);
not \U$13606 ( \13983 , \10226 );
or \U$13607 ( \13984 , \13982 , \13983 );
not \U$13608 ( \13985 , \10829 );
not \U$13609 ( \13986 , RIae79688_149);
nand \U$13610 ( \13987 , \13985 , \13986 );
nand \U$13611 ( \13988 , \13984 , \13987 );
not \U$13612 ( \13989 , \13988 );
or \U$13613 ( \13990 , \13981 , \13989 );
nand \U$13614 ( \13991 , \13249 , \9320 );
nand \U$13615 ( \13992 , \13990 , \13991 );
xor \U$13616 ( \13993 , \13980 , \13992 );
not \U$13617 ( \13994 , \2272 );
not \U$13618 ( \13995 , \13319 );
or \U$13619 ( \13996 , \13994 , \13995 );
and \U$13620 ( \13997 , RIae79ac0_158, \4982 );
not \U$13621 ( \13998 , RIae79ac0_158);
not \U$13622 ( \13999 , \3207 );
and \U$13623 ( \14000 , \13998 , \13999 );
nor \U$13624 ( \14001 , \13997 , \14000 );
nand \U$13625 ( \14002 , \10414 , \14001 );
nand \U$13626 ( \14003 , \13996 , \14002 );
xor \U$13627 ( \14004 , \13993 , \14003 );
and \U$13628 ( \14005 , \13969 , \14004 );
not \U$13629 ( \14006 , \13969 );
not \U$13630 ( \14007 , \14004 );
and \U$13631 ( \14008 , \14006 , \14007 );
nor \U$13632 ( \14009 , \14005 , \14008 );
not \U$13633 ( \14010 , \14009 );
not \U$13634 ( \14011 , \14010 );
or \U$13635 ( \14012 , \13961 , \14011 );
or \U$13636 ( \14013 , \13960 , \14010 );
nand \U$13637 ( \14014 , \14012 , \14013 );
not \U$13638 ( \14015 , \13460 );
not \U$13639 ( \14016 , \13451 );
or \U$13640 ( \14017 , \14015 , \14016 );
nand \U$13641 ( \14018 , \13447 , \13440 );
nand \U$13642 ( \14019 , \14017 , \14018 );
xor \U$13643 ( \14020 , \14014 , \14019 );
not \U$13644 ( \14021 , \4853 );
not \U$13645 ( \14022 , \11755 );
not \U$13646 ( \14023 , \3069 );
not \U$13647 ( \14024 , \14023 );
or \U$13648 ( \14025 , \14022 , \14024 );
nand \U$13649 ( \14026 , \10570 , RIae79ca0_162);
nand \U$13650 ( \14027 , \14025 , \14026 );
not \U$13651 ( \14028 , \14027 );
or \U$13652 ( \14029 , \14021 , \14028 );
nand \U$13653 ( \14030 , \13146 , \6276 );
nand \U$13654 ( \14031 , \14029 , \14030 );
not \U$13655 ( \14032 , \6091 );
not \U$13656 ( \14033 , \13065 );
or \U$13657 ( \14034 , \14032 , \14033 );
not \U$13658 ( \14035 , \4968 );
not \U$13659 ( \14036 , \12206 );
or \U$13660 ( \14037 , \14035 , \14036 );
or \U$13661 ( \14038 , \12206 , \4968 );
nand \U$13662 ( \14039 , \14037 , \14038 );
nand \U$13663 ( \14040 , \5049 , \14039 );
nand \U$13664 ( \14041 , \14034 , \14040 );
not \U$13665 ( \14042 , \14041 );
and \U$13666 ( \14043 , \14031 , \14042 );
not \U$13667 ( \14044 , \14031 );
and \U$13668 ( \14045 , \14044 , \14041 );
or \U$13669 ( \14046 , \14043 , \14045 );
not \U$13670 ( \14047 , \9622 );
and \U$13671 ( \14048 , \854 , RIae7a3a8_177);
not \U$13672 ( \14049 , \854 );
and \U$13673 ( \14050 , \14049 , \11690 );
nor \U$13674 ( \14051 , \14048 , \14050 );
not \U$13675 ( \14052 , \14051 );
or \U$13676 ( \14053 , \14047 , \14052 );
nand \U$13677 ( \14054 , \13170 , \11014 );
nand \U$13678 ( \14055 , \14053 , \14054 );
not \U$13679 ( \14056 , \14055 );
xnor \U$13680 ( \14057 , \14046 , \14056 );
not \U$13681 ( \14058 , \3440 );
not \U$13682 ( \14059 , RIae79520_146);
not \U$13683 ( \14060 , \1859 );
or \U$13684 ( \14061 , \14059 , \14060 );
or \U$13685 ( \14062 , \1859 , RIae79520_146);
nand \U$13686 ( \14063 , \14061 , \14062 );
not \U$13687 ( \14064 , \14063 );
or \U$13688 ( \14065 , \14058 , \14064 );
nand \U$13689 ( \14066 , \13330 , \12680 );
nand \U$13690 ( \14067 , \14065 , \14066 );
not \U$13691 ( \14068 , \9499 );
not \U$13692 ( \14069 , \13035 );
or \U$13693 ( \14070 , \14068 , \14069 );
buf \U$13694 ( \14071 , \2025 );
and \U$13695 ( \14072 , RIae79fe8_169, \14071 );
not \U$13696 ( \14073 , RIae79fe8_169);
and \U$13697 ( \14074 , \14073 , \2026 );
nor \U$13698 ( \14075 , \14072 , \14074 );
nand \U$13699 ( \14076 , \14075 , \10700 );
nand \U$13700 ( \14077 , \14070 , \14076 );
xor \U$13701 ( \14078 , \14067 , \14077 );
not \U$13702 ( \14079 , \2467 );
and \U$13703 ( \14080 , \4112 , \3810 );
not \U$13704 ( \14081 , \4112 );
and \U$13705 ( \14082 , \14081 , RIae794a8_145);
nor \U$13706 ( \14083 , \14080 , \14082 );
not \U$13707 ( \14084 , \14083 );
or \U$13708 ( \14085 , \14079 , \14084 );
nand \U$13709 ( \14086 , \13001 , \2458 );
nand \U$13710 ( \14087 , \14085 , \14086 );
xor \U$13711 ( \14088 , \14078 , \14087 );
nand \U$13712 ( \14089 , \14057 , \14088 );
not \U$13713 ( \14090 , \14057 );
not \U$13714 ( \14091 , \14088 );
nand \U$13715 ( \14092 , \14090 , \14091 );
nand \U$13716 ( \14093 , \14089 , \14092 );
not \U$13717 ( \14094 , \13517 );
not \U$13718 ( \14095 , \13509 );
or \U$13719 ( \14096 , \14094 , \14095 );
not \U$13720 ( \14097 , \13502 );
not \U$13721 ( \14098 , \13501 );
or \U$13722 ( \14099 , \14097 , \14098 );
nand \U$13723 ( \14100 , \14099 , \13508 );
nand \U$13724 ( \14101 , \14096 , \14100 );
not \U$13725 ( \14102 , \14101 );
and \U$13726 ( \14103 , \14093 , \14102 );
not \U$13727 ( \14104 , \14093 );
and \U$13728 ( \14105 , \14104 , \14101 );
nor \U$13729 ( \14106 , \14103 , \14105 );
xnor \U$13730 ( \14107 , \14020 , \14106 );
not \U$13731 ( \14108 , \10451 );
not \U$13732 ( \14109 , \997 );
buf \U$13733 ( \14110 , \9438 );
not \U$13734 ( \14111 , \14110 );
or \U$13735 ( \14112 , \14109 , \14111 );
or \U$13736 ( \14113 , \12614 , \6414 );
nand \U$13737 ( \14114 , \14112 , \14113 );
not \U$13738 ( \14115 , \14114 );
or \U$13739 ( \14116 , \14108 , \14115 );
nand \U$13740 ( \14117 , \13306 , \1008 );
nand \U$13741 ( \14118 , \14116 , \14117 );
not \U$13742 ( \14119 , \1863 );
not \U$13743 ( \14120 , \6230 );
and \U$13744 ( \14121 , \14120 , \1902 );
not \U$13745 ( \14122 , \14120 );
and \U$13746 ( \14123 , \14122 , RIae793b8_143);
nor \U$13747 ( \14124 , \14121 , \14123 );
not \U$13748 ( \14125 , \14124 );
or \U$13749 ( \14126 , \14119 , \14125 );
nand \U$13750 ( \14127 , \13272 , \1910 );
nand \U$13751 ( \14128 , \14126 , \14127 );
xor \U$13752 ( \14129 , \14118 , \14128 );
not \U$13753 ( \14130 , \1501 );
and \U$13754 ( \14131 , RIae79250_140, \12710 );
not \U$13755 ( \14132 , RIae79250_140);
and \U$13756 ( \14133 , \14132 , \12707 );
nor \U$13757 ( \14134 , \14131 , \14133 );
not \U$13758 ( \14135 , \14134 );
or \U$13759 ( \14136 , \14130 , \14135 );
nand \U$13760 ( \14137 , \13292 , \2650 );
nand \U$13761 ( \14138 , \14136 , \14137 );
xor \U$13762 ( \14139 , \14129 , \14138 );
xor \U$13763 ( \14140 , \13109 , \13119 );
and \U$13764 ( \14141 , \14140 , \13132 );
and \U$13765 ( \14142 , \13109 , \13119 );
or \U$13766 ( \14143 , \14141 , \14142 );
xor \U$13767 ( \14144 , \14139 , \14143 );
not \U$13768 ( \14145 , \839 );
and \U$13769 ( \14146 , RIae78f80_134, \10453 );
not \U$13770 ( \14147 , RIae78f80_134);
not \U$13771 ( \14148 , \10453 );
and \U$13772 ( \14149 , \14147 , \14148 );
or \U$13773 ( \14150 , \14146 , \14149 );
not \U$13774 ( \14151 , \14150 );
or \U$13775 ( \14152 , \14145 , \14151 );
nand \U$13776 ( \14153 , \13557 , \797 );
nand \U$13777 ( \14154 , \14152 , \14153 );
not \U$13778 ( \14155 , \1049 );
not \U$13779 ( \14156 , \10936 );
and \U$13780 ( \14157 , RIae79070_136, \14156 );
not \U$13781 ( \14158 , RIae79070_136);
and \U$13782 ( \14159 , \14158 , \9395 );
or \U$13783 ( \14160 , \14157 , \14159 );
not \U$13784 ( \14161 , \14160 );
or \U$13785 ( \14162 , \14155 , \14161 );
nand \U$13786 ( \14163 , \13283 , \1062 );
nand \U$13787 ( \14164 , \14162 , \14163 );
xor \U$13788 ( \14165 , \14154 , \14164 );
not \U$13789 ( \14166 , \9730 );
not \U$13790 ( \14167 , \13049 );
or \U$13791 ( \14168 , \14166 , \14167 );
nand \U$13792 ( \14169 , \10542 , RIae7a060_170);
nand \U$13793 ( \14170 , \14168 , \14169 );
xor \U$13794 ( \14171 , \14165 , \14170 );
xnor \U$13795 ( \14172 , \14144 , \14171 );
not \U$13796 ( \14173 , \13133 );
not \U$13797 ( \14174 , \13139 );
or \U$13798 ( \14175 , \14173 , \14174 );
nand \U$13799 ( \14176 , \14175 , \13173 );
not \U$13800 ( \14177 , \13133 );
nand \U$13801 ( \14178 , \14177 , \13137 , \13138 );
and \U$13802 ( \14179 , \14176 , \14178 );
xor \U$13803 ( \14180 , \14172 , \14179 );
xor \U$13804 ( \14181 , \13025 , \13054 );
and \U$13805 ( \14182 , \14181 , \13098 );
and \U$13806 ( \14183 , \13025 , \13054 );
or \U$13807 ( \14184 , \14182 , \14183 );
not \U$13808 ( \14185 , \14184 );
xor \U$13809 ( \14186 , \14180 , \14185 );
nand \U$13810 ( \14187 , \14107 , \14186 );
not \U$13811 ( \14188 , \14107 );
not \U$13812 ( \14189 , \14186 );
nand \U$13813 ( \14190 , \14188 , \14189 );
nand \U$13814 ( \14191 , \14187 , \14190 );
not \U$13815 ( \14192 , \13099 );
not \U$13816 ( \14193 , \13185 );
or \U$13817 ( \14194 , \14192 , \14193 );
nand \U$13818 ( \14195 , \14194 , \13174 );
not \U$13819 ( \14196 , \13099 );
nand \U$13820 ( \14197 , \14196 , \13184 );
nand \U$13821 ( \14198 , \14195 , \14197 );
not \U$13822 ( \14199 , \14198 );
and \U$13823 ( \14200 , \14191 , \14199 );
not \U$13824 ( \14201 , \14191 );
and \U$13825 ( \14202 , \14201 , \14198 );
nor \U$13826 ( \14203 , \14200 , \14202 );
xor \U$13827 ( \14204 , \13934 , \14203 );
not \U$13828 ( \14205 , \13361 );
not \U$13829 ( \14206 , \13604 );
or \U$13830 ( \14207 , \14205 , \14206 );
nand \U$13831 ( \14208 , \13598 , \13371 );
nand \U$13832 ( \14209 , \14207 , \14208 );
and \U$13833 ( \14210 , \14204 , \14209 );
not \U$13834 ( \14211 , \14204 );
not \U$13835 ( \14212 , \14209 );
and \U$13836 ( \14213 , \14211 , \14212 );
nor \U$13837 ( \14214 , \14210 , \14213 );
not \U$13838 ( \14215 , \14214 );
or \U$13839 ( \14216 , \13786 , \14215 );
not \U$13840 ( \14217 , \14214 );
nand \U$13841 ( \14218 , \14217 , \13784 );
nand \U$13842 ( \14219 , \14216 , \14218 );
nor \U$13843 ( \14220 , \13617 , \14219 );
xor \U$13844 ( \14221 , \13356 , \13608 );
xnor \U$13845 ( \14222 , \14221 , \12971 );
xor \U$13846 ( \14223 , \12027 , \11960 );
not \U$13847 ( \14224 , \14223 );
xor \U$13848 ( \14225 , \11638 , \11640 );
xor \U$13849 ( \14226 , \14225 , \11643 );
not \U$13850 ( \14227 , \14226 );
nand \U$13851 ( \14228 , \11618 , \11615 );
nand \U$13852 ( \14229 , \11633 , \14228 );
and \U$13853 ( \14230 , \14229 , \11629 );
not \U$13854 ( \14231 , \14229 );
not \U$13855 ( \14232 , \11629 );
and \U$13856 ( \14233 , \14231 , \14232 );
nor \U$13857 ( \14234 , \14230 , \14233 );
not \U$13858 ( \14235 , \14234 );
not \U$13859 ( \14236 , \14235 );
or \U$13860 ( \14237 , \14227 , \14236 );
xor \U$13861 ( \14238 , \12642 , \12775 );
xor \U$13862 ( \14239 , \14238 , \12818 );
nand \U$13863 ( \14240 , \14237 , \14239 );
not \U$13864 ( \14241 , \14226 );
nand \U$13865 ( \14242 , \14241 , \14234 );
nand \U$13866 ( \14243 , \14240 , \14242 );
not \U$13867 ( \14244 , \14243 );
xor \U$13868 ( \14245 , \12008 , \12012 );
xnor \U$13869 ( \14246 , \14245 , \12021 );
not \U$13870 ( \14247 , \14246 );
or \U$13871 ( \14248 , \14244 , \14247 );
or \U$13872 ( \14249 , \14246 , \14243 );
not \U$13873 ( \14250 , \11635 );
not \U$13874 ( \14251 , \11550 );
or \U$13875 ( \14252 , \14250 , \14251 );
or \U$13876 ( \14253 , \11550 , \11635 );
nand \U$13877 ( \14254 , \14252 , \14253 );
not \U$13878 ( \14255 , \11646 );
and \U$13879 ( \14256 , \14254 , \14255 );
not \U$13880 ( \14257 , \14254 );
and \U$13881 ( \14258 , \14257 , \11646 );
nor \U$13882 ( \14259 , \14256 , \14258 );
not \U$13883 ( \14260 , \14259 );
nand \U$13884 ( \14261 , \14249 , \14260 );
nand \U$13885 ( \14262 , \14248 , \14261 );
buf \U$13886 ( \14263 , \14262 );
not \U$13887 ( \14264 , \14263 );
xor \U$13888 ( \14265 , \11465 , \11472 );
xnor \U$13889 ( \14266 , \14265 , \11463 );
not \U$13890 ( \14267 , \14266 );
xor \U$13891 ( \14268 , \11004 , \10991 );
xnor \U$13892 ( \14269 , \14268 , \10880 );
xor \U$13893 ( \14270 , \11050 , \11095 );
xnor \U$13894 ( \14271 , \14270 , \11139 );
not \U$13895 ( \14272 , \14271 );
xor \U$13896 ( \14273 , \11559 , \11611 );
not \U$13897 ( \14274 , \14273 );
xor \U$13898 ( \14275 , \11306 , \11341 );
not \U$13899 ( \14276 , \13720 );
xor \U$13900 ( \14277 , RIae7a240_174, \2207 );
not \U$13901 ( \14278 , \14277 );
or \U$13902 ( \14279 , \14276 , \14278 );
nand \U$13903 ( \14280 , \11119 , \13121 );
nand \U$13904 ( \14281 , \14279 , \14280 );
not \U$13905 ( \14282 , \14281 );
not \U$13906 ( \14283 , \9730 );
and \U$13907 ( \14284 , RIae7a060_170, \854 );
not \U$13908 ( \14285 , RIae7a060_170);
and \U$13909 ( \14286 , \14285 , \1022 );
nor \U$13910 ( \14287 , \14284 , \14286 );
not \U$13911 ( \14288 , \14287 );
or \U$13912 ( \14289 , \14283 , \14288 );
nand \U$13913 ( \14290 , \11107 , \10542 );
nand \U$13914 ( \14291 , \14289 , \14290 );
not \U$13915 ( \14292 , \14291 );
or \U$13916 ( \14293 , \14282 , \14292 );
or \U$13917 ( \14294 , \14291 , \14281 );
not \U$13918 ( \14295 , \10510 );
not \U$13919 ( \14296 , RIae7a7e0_186);
not \U$13920 ( \14297 , \1439 );
or \U$13921 ( \14298 , \14296 , \14297 );
or \U$13922 ( \14299 , \3443 , RIae7a7e0_186);
nand \U$13923 ( \14300 , \14298 , \14299 );
not \U$13924 ( \14301 , \14300 );
or \U$13925 ( \14302 , \14295 , \14301 );
not \U$13926 ( \14303 , \11446 );
nand \U$13927 ( \14304 , \14303 , \10519 );
nand \U$13928 ( \14305 , \14302 , \14304 );
nand \U$13929 ( \14306 , \14294 , \14305 );
nand \U$13930 ( \14307 , \14293 , \14306 );
xor \U$13931 ( \14308 , \14275 , \14307 );
not \U$13932 ( \14309 , \14308 );
or \U$13933 ( \14310 , \14274 , \14309 );
nand \U$13934 ( \14311 , \14307 , \14275 );
nand \U$13935 ( \14312 , \14310 , \14311 );
not \U$13936 ( \14313 , \14312 );
not \U$13937 ( \14314 , \14313 );
xor \U$13938 ( \14315 , \11407 , \11459 );
not \U$13939 ( \14316 , \14315 );
or \U$13940 ( \14317 , \14314 , \14316 );
or \U$13941 ( \14318 , \14315 , \14313 );
nand \U$13942 ( \14319 , \14317 , \14318 );
not \U$13943 ( \14320 , \14319 );
or \U$13944 ( \14321 , \14272 , \14320 );
not \U$13945 ( \14322 , \14313 );
nand \U$13946 ( \14323 , \14322 , \14315 );
nand \U$13947 ( \14324 , \14321 , \14323 );
xnor \U$13948 ( \14325 , \14269 , \14324 );
not \U$13949 ( \14326 , \14325 );
or \U$13950 ( \14327 , \14267 , \14326 );
not \U$13951 ( \14328 , \14269 );
nand \U$13952 ( \14329 , \14328 , \14324 );
nand \U$13953 ( \14330 , \14327 , \14329 );
not \U$13954 ( \14331 , \14330 );
not \U$13955 ( \14332 , \14331 );
or \U$13956 ( \14333 , \14264 , \14332 );
or \U$13957 ( \14334 , \14331 , \14263 );
nand \U$13958 ( \14335 , \14333 , \14334 );
not \U$13959 ( \14336 , \14335 );
or \U$13960 ( \14337 , \14224 , \14336 );
nand \U$13961 ( \14338 , \14330 , \14263 );
nand \U$13962 ( \14339 , \14337 , \14338 );
not \U$13963 ( \14340 , \14339 );
not \U$13964 ( \14341 , \14340 );
not \U$13965 ( \14342 , \12968 );
not \U$13966 ( \14343 , \11749 );
or \U$13967 ( \14344 , \14342 , \14343 );
or \U$13968 ( \14345 , \12968 , \11749 );
nand \U$13969 ( \14346 , \14344 , \14345 );
xnor \U$13970 ( \14347 , \14346 , \12460 );
not \U$13971 ( \14348 , \14347 );
or \U$13972 ( \14349 , \14341 , \14348 );
xor \U$13973 ( \14350 , \12778 , \12812 );
xor \U$13974 ( \14351 , \14350 , \12815 );
not \U$13975 ( \14352 , \14351 );
not \U$13976 ( \14353 , \14352 );
xor \U$13977 ( \14354 , \12579 , \12536 );
not \U$13978 ( \14355 , \14354 );
or \U$13979 ( \14356 , \14353 , \14355 );
xor \U$13980 ( \14357 , \12679 , \12719 );
xor \U$13981 ( \14358 , \14357 , \12772 );
nand \U$13982 ( \14359 , \14356 , \14358 );
not \U$13983 ( \14360 , \14354 );
nand \U$13984 ( \14361 , \14360 , \14351 );
nand \U$13985 ( \14362 , \14359 , \14361 );
not \U$13986 ( \14363 , \14362 );
xor \U$13987 ( \14364 , \12595 , \12639 );
xnor \U$13988 ( \14365 , \14364 , \12632 );
not \U$13989 ( \14366 , \14365 );
not \U$13990 ( \14367 , \9527 );
not \U$13991 ( \14368 , \14300 );
or \U$13992 ( \14369 , \14367 , \14368 );
not \U$13993 ( \14370 , \9770 );
not \U$13994 ( \14371 , RIae7a7e0_186);
and \U$13995 ( \14372 , \14370 , \14371 );
and \U$13996 ( \14373 , \3236 , RIae7a7e0_186);
nor \U$13997 ( \14374 , \14372 , \14373 );
nand \U$13998 ( \14375 , \14374 , \10510 );
nand \U$13999 ( \14376 , \14369 , \14375 );
not \U$14000 ( \14377 , \9622 );
not \U$14001 ( \14378 , \12514 );
or \U$14002 ( \14379 , \14377 , \14378 );
not \U$14003 ( \14380 , \11690 );
not \U$14004 ( \14381 , \1899 );
or \U$14005 ( \14382 , \14380 , \14381 );
or \U$14006 ( \14383 , \1899 , \13165 );
nand \U$14007 ( \14384 , \14382 , \14383 );
nand \U$14008 ( \14385 , \14384 , \9644 );
nand \U$14009 ( \14386 , \14379 , \14385 );
xor \U$14010 ( \14387 , \14376 , \14386 );
not \U$14011 ( \14388 , \9687 );
xor \U$14012 ( \14389 , RIae7a240_174, \9512 );
not \U$14013 ( \14390 , \14389 );
or \U$14014 ( \14391 , \14388 , \14390 );
nand \U$14015 ( \14392 , \14277 , \13121 );
nand \U$14016 ( \14393 , \14391 , \14392 );
and \U$14017 ( \14394 , \14387 , \14393 );
and \U$14018 ( \14395 , \14376 , \14386 );
nor \U$14019 ( \14396 , \14394 , \14395 );
not \U$14020 ( \14397 , \14396 );
not \U$14021 ( \14398 , \1863 );
not \U$14022 ( \14399 , \12488 );
or \U$14023 ( \14400 , \14398 , \14399 );
and \U$14024 ( \14401 , RIae793b8_143, \11187 );
not \U$14025 ( \14402 , RIae793b8_143);
and \U$14026 ( \14403 , \14402 , \10465 );
or \U$14027 ( \14404 , \14401 , \14403 );
nand \U$14028 ( \14405 , \14404 , \1910 );
nand \U$14029 ( \14406 , \14400 , \14405 );
not \U$14030 ( \14407 , \2011 );
not \U$14031 ( \14408 , \12605 );
or \U$14032 ( \14409 , \14407 , \14408 );
and \U$14033 ( \14410 , RIae79610_148, \9412 );
not \U$14034 ( \14411 , RIae79610_148);
and \U$14035 ( \14412 , \14411 , \11198 );
or \U$14036 ( \14413 , \14410 , \14412 );
nand \U$14037 ( \14414 , \14413 , \2063 );
nand \U$14038 ( \14415 , \14409 , \14414 );
xor \U$14039 ( \14416 , \14406 , \14415 );
buf \U$14040 ( \14417 , \14416 );
not \U$14041 ( \14418 , \2776 );
not \U$14042 ( \14419 , \12473 );
or \U$14043 ( \14420 , \14418 , \14419 );
not \U$14044 ( \14421 , \10584 );
not \U$14045 ( \14422 , \1969 );
not \U$14046 ( \14423 , \14422 );
or \U$14047 ( \14424 , \14421 , \14423 );
nand \U$14048 ( \14425 , \3216 , RIae79c28_161);
nand \U$14049 ( \14426 , \14424 , \14425 );
nand \U$14050 ( \14427 , \14426 , \2767 );
nand \U$14051 ( \14428 , \14420 , \14427 );
and \U$14052 ( \14429 , \14417 , \14428 );
and \U$14053 ( \14430 , \14406 , \14415 );
nor \U$14054 ( \14431 , \14429 , \14430 );
not \U$14055 ( \14432 , \14431 );
not \U$14056 ( \14433 , \4853 );
not \U$14057 ( \14434 , \12909 );
or \U$14058 ( \14435 , \14433 , \14434 );
not \U$14059 ( \14436 , RIae79ca0_162);
not \U$14060 ( \14437 , \13008 );
or \U$14061 ( \14438 , \14436 , \14437 );
not \U$14062 ( \14439 , \2093 );
or \U$14063 ( \14440 , \14439 , RIae79ca0_162);
nand \U$14064 ( \14441 , \14438 , \14440 );
nand \U$14065 ( \14442 , \14441 , \11761 );
nand \U$14066 ( \14443 , \14435 , \14442 );
not \U$14067 ( \14444 , \14443 );
not \U$14068 ( \14445 , \14444 );
not \U$14069 ( \14446 , RIae79d90_164);
not \U$14070 ( \14447 , \1789 );
or \U$14071 ( \14448 , \14446 , \14447 );
nand \U$14072 ( \14449 , \11680 , \6084 );
nand \U$14073 ( \14450 , \14448 , \14449 );
not \U$14074 ( \14451 , \14450 );
not \U$14075 ( \14452 , \6091 );
or \U$14076 ( \14453 , \14451 , \14452 );
nand \U$14077 ( \14454 , \12793 , \5049 );
nand \U$14078 ( \14455 , \14453 , \14454 );
not \U$14079 ( \14456 , \14455 );
not \U$14080 ( \14457 , \14456 );
or \U$14081 ( \14458 , \14445 , \14457 );
not \U$14082 ( \14459 , \10677 );
not \U$14083 ( \14460 , \12899 );
or \U$14084 ( \14461 , \14459 , \14460 );
not \U$14085 ( \14462 , RIae7a498_179);
not \U$14086 ( \14463 , \2101 );
or \U$14087 ( \14464 , \14462 , \14463 );
or \U$14088 ( \14465 , \6147 , RIae7a498_179);
nand \U$14089 ( \14466 , \14464 , \14465 );
nand \U$14090 ( \14467 , \14466 , \10696 );
nand \U$14091 ( \14468 , \14461 , \14467 );
nand \U$14092 ( \14469 , \14458 , \14468 );
not \U$14093 ( \14470 , \14456 );
nand \U$14094 ( \14471 , \14470 , \14443 );
nand \U$14095 ( \14472 , \14469 , \14471 );
nand \U$14096 ( \14473 , \14432 , \14472 );
not \U$14097 ( \14474 , \14473 );
or \U$14098 ( \14475 , \14397 , \14474 );
and \U$14099 ( \14476 , \14469 , \14431 , \14471 );
not \U$14100 ( \14477 , \14476 );
nand \U$14101 ( \14478 , \14475 , \14477 );
not \U$14102 ( \14479 , \14478 );
not \U$14103 ( \14480 , \14479 );
or \U$14104 ( \14481 , \14366 , \14480 );
not \U$14105 ( \14482 , \14365 );
not \U$14106 ( \14483 , \14482 );
not \U$14107 ( \14484 , \14478 );
or \U$14108 ( \14485 , \14483 , \14484 );
not \U$14109 ( \14486 , \11037 );
not \U$14110 ( \14487 , \12504 );
or \U$14111 ( \14488 , \14486 , \14487 );
xnor \U$14112 ( \14489 , \2402 , RIae79778_151);
nand \U$14113 ( \14490 , \14489 , \9576 );
nand \U$14114 ( \14491 , \14488 , \14490 );
not \U$14115 ( \14492 , \10927 );
and \U$14116 ( \14493 , RIae7a510_180, \13032 );
not \U$14117 ( \14494 , RIae7a510_180);
and \U$14118 ( \14495 , \14494 , \2047 );
nor \U$14119 ( \14496 , \14493 , \14495 );
not \U$14120 ( \14497 , \14496 );
or \U$14121 ( \14498 , \14492 , \14497 );
nand \U$14122 ( \14499 , \12465 , \10631 );
nand \U$14123 ( \14500 , \14498 , \14499 );
xor \U$14124 ( \14501 , \14491 , \14500 );
not \U$14125 ( \14502 , \10275 );
not \U$14126 ( \14503 , \12524 );
or \U$14127 ( \14504 , \14502 , \14503 );
not \U$14128 ( \14505 , RIae7a8d0_188);
not \U$14129 ( \14506 , \1993 );
or \U$14130 ( \14507 , \14505 , \14506 );
or \U$14131 ( \14508 , \1993 , RIae7a8d0_188);
nand \U$14132 ( \14509 , \14507 , \14508 );
buf \U$14133 ( \14510 , \11204 );
nand \U$14134 ( \14511 , \14509 , \14510 );
nand \U$14135 ( \14512 , \14504 , \14511 );
and \U$14136 ( \14513 , \14501 , \14512 );
and \U$14137 ( \14514 , \14491 , \14500 );
or \U$14138 ( \14515 , \14513 , \14514 );
xor \U$14139 ( \14516 , \12693 , \12704 );
xor \U$14140 ( \14517 , \14516 , \12716 );
or \U$14141 ( \14518 , \14515 , \14517 );
xor \U$14142 ( \14519 , \12768 , \12730 );
xnor \U$14143 ( \14520 , \14519 , \12740 );
nand \U$14144 ( \14521 , \14518 , \14520 );
nand \U$14145 ( \14522 , \14517 , \14515 );
nand \U$14146 ( \14523 , \14521 , \14522 );
nand \U$14147 ( \14524 , \14485 , \14523 );
nand \U$14148 ( \14525 , \14481 , \14524 );
xor \U$14149 ( \14526 , \11570 , \11596 );
not \U$14150 ( \14527 , \838 );
not \U$14151 ( \14528 , \12669 );
or \U$14152 ( \14529 , \14527 , \14528 );
and \U$14153 ( \14530 , RIae78f80_134, \10149 );
not \U$14154 ( \14531 , RIae78f80_134);
and \U$14155 ( \14532 , \14531 , \10142 );
or \U$14156 ( \14533 , \14530 , \14532 );
nand \U$14157 ( \14534 , \14533 , \796 );
nand \U$14158 ( \14535 , \14529 , \14534 );
not \U$14159 ( \14536 , \1049 );
not \U$14160 ( \14537 , \12660 );
or \U$14161 ( \14538 , \14536 , \14537 );
xor \U$14162 ( \14539 , RIae79070_136, \10007 );
nand \U$14163 ( \14540 , \14539 , \1062 );
nand \U$14164 ( \14541 , \14538 , \14540 );
or \U$14165 ( \14542 , \14535 , \14541 );
not \U$14166 ( \14543 , \10451 );
not \U$14167 ( \14544 , \11566 );
or \U$14168 ( \14545 , \14543 , \14544 );
not \U$14169 ( \14546 , \9897 );
xor \U$14170 ( \14547 , RIae79160_138, \14546 );
nand \U$14171 ( \14548 , \14547 , \1008 );
nand \U$14172 ( \14549 , \14545 , \14548 );
nand \U$14173 ( \14550 , \14542 , \14549 );
nand \U$14174 ( \14551 , \14541 , \14535 );
nand \U$14175 ( \14552 , \14550 , \14551 );
or \U$14176 ( \14553 , \14526 , \14552 );
not \U$14177 ( \14554 , \14553 );
not \U$14178 ( \14555 , \2007 );
not \U$14179 ( \14556 , \12736 );
or \U$14180 ( \14557 , \14555 , \14556 );
and \U$14181 ( \14558 , \2521 , \6238 );
not \U$14182 ( \14559 , \2521 );
and \U$14183 ( \14560 , \14559 , \4169 );
nor \U$14184 ( \14561 , \14558 , \14560 );
nand \U$14185 ( \14562 , \14561 , \1988 );
nand \U$14186 ( \14563 , \14557 , \14562 );
not \U$14187 ( \14564 , \12764 );
not \U$14188 ( \14565 , \12753 );
and \U$14189 ( \14566 , \14564 , \14565 );
and \U$14190 ( \14567 , \12764 , \12753 );
nor \U$14191 ( \14568 , \14566 , \14567 );
not \U$14192 ( \14569 , \14568 );
or \U$14193 ( \14570 , \14563 , \14569 );
not \U$14194 ( \14571 , \2322 );
not \U$14195 ( \14572 , \12726 );
or \U$14196 ( \14573 , \14571 , \14572 );
not \U$14197 ( \14574 , RIae798e0_154);
not \U$14198 ( \14575 , \13248 );
or \U$14199 ( \14576 , \14574 , \14575 );
not \U$14200 ( \14577 , \10237 );
nand \U$14201 ( \14578 , \14577 , \2334 );
nand \U$14202 ( \14579 , \14576 , \14578 );
buf \U$14203 ( \14580 , \2339 );
nand \U$14204 ( \14581 , \14579 , \14580 );
nand \U$14205 ( \14582 , \14573 , \14581 );
nand \U$14206 ( \14583 , \14570 , \14582 );
nand \U$14207 ( \14584 , \14563 , \14569 );
nand \U$14208 ( \14585 , \14583 , \14584 );
not \U$14209 ( \14586 , \14585 );
or \U$14210 ( \14587 , \14554 , \14586 );
nand \U$14211 ( \14588 , \14526 , \14552 );
nand \U$14212 ( \14589 , \14587 , \14588 );
not \U$14213 ( \14590 , \14589 );
not \U$14214 ( \14591 , \12674 );
nand \U$14215 ( \14592 , \14591 , \12678 );
xor \U$14216 ( \14593 , \12653 , \14592 );
not \U$14217 ( \14594 , \797 );
xor \U$14218 ( \14595 , RIae78f80_134, \10032 );
not \U$14219 ( \14596 , \14595 );
or \U$14220 ( \14597 , \14594 , \14596 );
nand \U$14221 ( \14598 , \14533 , \838 );
nand \U$14222 ( \14599 , \14597 , \14598 );
not \U$14223 ( \14600 , \14599 );
not \U$14224 ( \14601 , \12857 );
or \U$14225 ( \14602 , \14601 , \865 );
nand \U$14226 ( \14603 , \14602 , \863 , RIae78b48_125);
not \U$14227 ( \14604 , \14603 );
not \U$14228 ( \14605 , \892 );
xor \U$14229 ( \14606 , RIae78b48_125, \12858 );
not \U$14230 ( \14607 , \14606 );
or \U$14231 ( \14608 , \14605 , \14607 );
nand \U$14232 ( \14609 , \12752 , \12863 , \867 );
nand \U$14233 ( \14610 , \14608 , \14609 );
nand \U$14234 ( \14611 , \14604 , \14610 );
not \U$14235 ( \14612 , \1072 );
not \U$14236 ( \14613 , \12762 );
or \U$14237 ( \14614 , \14612 , \14613 );
and \U$14238 ( \14615 , \10193 , RIae78e90_132);
not \U$14239 ( \14616 , \10193 );
and \U$14240 ( \14617 , \14616 , \1066 );
nor \U$14241 ( \14618 , \14615 , \14617 );
nand \U$14242 ( \14619 , \14618 , \1086 );
nand \U$14243 ( \14620 , \14614 , \14619 );
xnor \U$14244 ( \14621 , \14611 , \14620 );
not \U$14245 ( \14622 , \14621 );
or \U$14246 ( \14623 , \14600 , \14622 );
not \U$14247 ( \14624 , \14611 );
nand \U$14248 ( \14625 , \14624 , \14620 );
nand \U$14249 ( \14626 , \14623 , \14625 );
not \U$14250 ( \14627 , \1933 );
and \U$14251 ( \14628 , RIae794a8_145, \9286 );
not \U$14252 ( \14629 , RIae794a8_145);
not \U$14253 ( \14630 , \9290 );
not \U$14254 ( \14631 , \14630 );
and \U$14255 ( \14632 , \14629 , \14631 );
or \U$14256 ( \14633 , \14628 , \14632 );
not \U$14257 ( \14634 , \14633 );
or \U$14258 ( \14635 , \14627 , \14634 );
nand \U$14259 ( \14636 , \12702 , \2467 );
nand \U$14260 ( \14637 , \14635 , \14636 );
xor \U$14261 ( \14638 , \14626 , \14637 );
not \U$14262 ( \14639 , \10223 );
not \U$14263 ( \14640 , \12689 );
or \U$14264 ( \14641 , \14639 , \14640 );
and \U$14265 ( \14642 , RIae79520_146, \9313 );
not \U$14266 ( \14643 , RIae79520_146);
not \U$14267 ( \14644 , \9313 );
and \U$14268 ( \14645 , \14643 , \14644 );
or \U$14269 ( \14646 , \14642 , \14645 );
nand \U$14270 ( \14647 , \14646 , \2189 );
nand \U$14271 ( \14648 , \14641 , \14647 );
and \U$14272 ( \14649 , \14638 , \14648 );
and \U$14273 ( \14650 , \14626 , \14637 );
nor \U$14274 ( \14651 , \14649 , \14650 );
xor \U$14275 ( \14652 , \14593 , \14651 );
not \U$14276 ( \14653 , \1820 );
not \U$14277 ( \14654 , \12619 );
or \U$14278 ( \14655 , \14653 , \14654 );
not \U$14279 ( \14656 , RIae79688_149);
not \U$14280 ( \14657 , \9459 );
not \U$14281 ( \14658 , \14657 );
or \U$14282 ( \14659 , \14656 , \14658 );
or \U$14283 ( \14660 , \13302 , RIae79688_149);
nand \U$14284 ( \14661 , \14659 , \14660 );
nand \U$14285 ( \14662 , \14661 , \9320 );
nand \U$14286 ( \14663 , \14655 , \14662 );
not \U$14287 ( \14664 , \14663 );
not \U$14288 ( \14665 , \14664 );
not \U$14289 ( \14666 , RIae7aab0_192);
and \U$14290 ( \14667 , \14666 , RIae7aa38_191);
buf \U$14291 ( \14668 , \14667 );
buf \U$14292 ( \14669 , \14668 );
not \U$14293 ( \14670 , \14669 );
not \U$14294 ( \14671 , RIae7aa38_191);
not \U$14295 ( \14672 , \14671 );
not \U$14296 ( \14673 , \991 );
or \U$14297 ( \14674 , \14672 , \14673 );
or \U$14298 ( \14675 , \991 , \14671 );
nand \U$14299 ( \14676 , \14674 , \14675 );
not \U$14300 ( \14677 , \14676 );
or \U$14301 ( \14678 , \14670 , \14677 );
nand \U$14302 ( \14679 , RIae7aa38_191, RIae7aab0_192);
nand \U$14303 ( \14680 , \14678 , \14679 );
not \U$14304 ( \14681 , \14680 );
not \U$14305 ( \14682 , \14681 );
or \U$14306 ( \14683 , \14665 , \14682 );
not \U$14307 ( \14684 , \14663 );
not \U$14308 ( \14685 , \14680 );
or \U$14309 ( \14686 , \14684 , \14685 );
not \U$14310 ( \14687 , \3014 );
not \U$14311 ( \14688 , \12712 );
or \U$14312 ( \14689 , \14687 , \14688 );
not \U$14313 ( \14690 , \2268 );
buf \U$14314 ( \14691 , \9363 );
not \U$14315 ( \14692 , \14691 );
or \U$14316 ( \14693 , \14690 , \14692 );
or \U$14317 ( \14694 , \14691 , \2268 );
nand \U$14318 ( \14695 , \14693 , \14694 );
nand \U$14319 ( \14696 , \2272 , \14695 );
nand \U$14320 ( \14697 , \14689 , \14696 );
not \U$14321 ( \14698 , \14697 );
nand \U$14322 ( \14699 , \14686 , \14698 );
nand \U$14323 ( \14700 , \14683 , \14699 );
and \U$14324 ( \14701 , \14652 , \14700 );
and \U$14325 ( \14702 , \14593 , \14651 );
or \U$14326 ( \14703 , \14701 , \14702 );
nand \U$14327 ( \14704 , \14590 , \14703 );
not \U$14328 ( \14705 , \14704 );
not \U$14329 ( \14706 , \9815 );
not \U$14330 ( \14707 , \12566 );
or \U$14331 ( \14708 , \14706 , \14707 );
not \U$14332 ( \14709 , RIae7a2b8_175);
not \U$14333 ( \14710 , \2954 );
or \U$14334 ( \14711 , \14709 , \14710 );
not \U$14335 ( \14712 , \5631 );
or \U$14336 ( \14713 , \14712 , RIae7a2b8_175);
nand \U$14337 ( \14714 , \14711 , \14713 );
nand \U$14338 ( \14715 , \14714 , \9792 );
nand \U$14339 ( \14716 , \14708 , \14715 );
not \U$14340 ( \14717 , \14716 );
not \U$14341 ( \14718 , \9745 );
not \U$14342 ( \14719 , \14287 );
or \U$14343 ( \14720 , \14718 , \14719 );
not \U$14344 ( \14721 , RIae7a060_170);
not \U$14345 ( \14722 , \14721 );
not \U$14346 ( \14723 , \5351 );
or \U$14347 ( \14724 , \14722 , \14723 );
or \U$14348 ( \14725 , \883 , \14721 );
nand \U$14349 ( \14726 , \14724 , \14725 );
nand \U$14350 ( \14727 , \14726 , \9730 );
nand \U$14351 ( \14728 , \14720 , \14727 );
not \U$14352 ( \14729 , \14728 );
nand \U$14353 ( \14730 , \14717 , \14729 );
not \U$14354 ( \14731 , \9705 );
not \U$14355 ( \14732 , \12554 );
or \U$14356 ( \14733 , \14731 , \14732 );
not \U$14357 ( \14734 , RIae7a6f0_184);
not \U$14358 ( \14735 , \2510 );
or \U$14359 ( \14736 , \14734 , \14735 );
or \U$14360 ( \14737 , \2331 , RIae7a6f0_184);
nand \U$14361 ( \14738 , \14736 , \14737 );
nand \U$14362 ( \14739 , \14738 , \9473 );
nand \U$14363 ( \14740 , \14733 , \14739 );
and \U$14364 ( \14741 , \14730 , \14740 );
and \U$14365 ( \14742 , \14728 , \14716 );
nor \U$14366 ( \14743 , \14741 , \14742 );
not \U$14367 ( \14744 , \14743 );
xor \U$14368 ( \14745 , \12611 , \12609 );
xnor \U$14369 ( \14746 , \14745 , \12623 );
not \U$14370 ( \14747 , \14746 );
not \U$14371 ( \14748 , \9517 );
not \U$14372 ( \14749 , \12543 );
or \U$14373 ( \14750 , \14748 , \14749 );
not \U$14374 ( \14751 , RIae79fe8_169);
not \U$14375 ( \14752 , \10534 );
or \U$14376 ( \14753 , \14751 , \14752 );
or \U$14377 ( \14754 , \2287 , RIae79fe8_169);
nand \U$14378 ( \14755 , \14753 , \14754 );
nand \U$14379 ( \14756 , \14755 , \11914 );
nand \U$14380 ( \14757 , \14750 , \14756 );
not \U$14381 ( \14758 , \14757 );
not \U$14382 ( \14759 , \14758 );
not \U$14383 ( \14760 , \6214 );
not \U$14384 ( \14761 , \12786 );
or \U$14385 ( \14762 , \14760 , \14761 );
not \U$14386 ( \14763 , \1759 );
not \U$14387 ( \14764 , RIae79ef8_167);
and \U$14388 ( \14765 , \14763 , \14764 );
and \U$14389 ( \14766 , \1755 , RIae79ef8_167);
nor \U$14390 ( \14767 , \14765 , \14766 );
buf \U$14391 ( \14768 , \6201 );
nand \U$14392 ( \14769 , \14767 , \14768 );
nand \U$14393 ( \14770 , \14762 , \14769 );
not \U$14394 ( \14771 , \14770 );
not \U$14395 ( \14772 , \14771 );
or \U$14396 ( \14773 , \14759 , \14772 );
not \U$14397 ( \14774 , \9777 );
not \U$14398 ( \14775 , \12805 );
or \U$14399 ( \14776 , \14774 , \14775 );
not \U$14400 ( \14777 , RIae7a150_172);
not \U$14401 ( \14778 , \11694 );
not \U$14402 ( \14779 , \14778 );
or \U$14403 ( \14780 , \14777 , \14779 );
or \U$14404 ( \14781 , \5081 , RIae7a150_172);
nand \U$14405 ( \14782 , \14780 , \14781 );
nand \U$14406 ( \14783 , \14782 , \11087 );
nand \U$14407 ( \14784 , \14776 , \14783 );
nand \U$14408 ( \14785 , \14773 , \14784 );
not \U$14409 ( \14786 , \14758 );
nand \U$14410 ( \14787 , \14786 , \14770 );
and \U$14411 ( \14788 , \14785 , \14787 );
nand \U$14412 ( \14789 , \14747 , \14788 );
nand \U$14413 ( \14790 , \14744 , \14789 );
not \U$14414 ( \14791 , \14788 );
nand \U$14415 ( \14792 , \14791 , \14746 );
nand \U$14416 ( \14793 , \14790 , \14792 );
not \U$14417 ( \14794 , \14793 );
or \U$14418 ( \14795 , \14705 , \14794 );
not \U$14419 ( \14796 , \14703 );
nand \U$14420 ( \14797 , \14796 , \14589 );
nand \U$14421 ( \14798 , \14795 , \14797 );
xor \U$14422 ( \14799 , \14525 , \14798 );
not \U$14423 ( \14800 , \14799 );
or \U$14424 ( \14801 , \14363 , \14800 );
nand \U$14425 ( \14802 , \14798 , \14525 );
nand \U$14426 ( \14803 , \14801 , \14802 );
not \U$14427 ( \14804 , \14803 );
xor \U$14428 ( \14805 , \12590 , \12821 );
xor \U$14429 ( \14806 , \14805 , \12949 );
not \U$14430 ( \14807 , \14806 );
or \U$14431 ( \14808 , \14804 , \14807 );
not \U$14432 ( \14809 , \14803 );
not \U$14433 ( \14810 , \14809 );
not \U$14434 ( \14811 , \14806 );
not \U$14435 ( \14812 , \14811 );
or \U$14436 ( \14813 , \14810 , \14812 );
and \U$14437 ( \14814 , \12947 , \12829 );
not \U$14438 ( \14815 , \12947 );
and \U$14439 ( \14816 , \14815 , \12830 );
nor \U$14440 ( \14817 , \14814 , \14816 );
xnor \U$14441 ( \14818 , \12919 , \14817 );
not \U$14442 ( \14819 , \14818 );
xor \U$14443 ( \14820 , \12584 , \12586 );
xor \U$14444 ( \14821 , \14820 , \12583 );
xor \U$14445 ( \14822 , \14305 , \14281 );
xor \U$14446 ( \14823 , \14291 , \14822 );
not \U$14447 ( \14824 , \14823 );
xor \U$14448 ( \14825 , \12545 , \12559 );
xnor \U$14449 ( \14826 , \14825 , \12577 );
not \U$14450 ( \14827 , \14826 );
or \U$14451 ( \14828 , \14824 , \14827 );
or \U$14452 ( \14829 , \14826 , \14823 );
xor \U$14453 ( \14830 , \12506 , \12517 );
xor \U$14454 ( \14831 , \14830 , \12528 );
nand \U$14455 ( \14832 , \14829 , \14831 );
nand \U$14456 ( \14833 , \14828 , \14832 );
not \U$14457 ( \14834 , \14833 );
not \U$14458 ( \14835 , \14273 );
and \U$14459 ( \14836 , \14308 , \14835 );
not \U$14460 ( \14837 , \14308 );
and \U$14461 ( \14838 , \14837 , \14273 );
nor \U$14462 ( \14839 , \14836 , \14838 );
not \U$14463 ( \14840 , \14839 );
xor \U$14464 ( \14841 , \12897 , \12911 );
xnor \U$14465 ( \14842 , \14841 , \12903 );
not \U$14466 ( \14843 , \14842 );
xor \U$14467 ( \14844 , \12494 , \12477 );
xnor \U$14468 ( \14845 , \14844 , \12467 );
not \U$14469 ( \14846 , \14845 );
or \U$14470 ( \14847 , \14843 , \14846 );
or \U$14471 ( \14848 , \14842 , \14845 );
xor \U$14472 ( \14849 , \12788 , \12797 );
xor \U$14473 ( \14850 , \14849 , \12809 );
nand \U$14474 ( \14851 , \14848 , \14850 );
nand \U$14475 ( \14852 , \14847 , \14851 );
not \U$14476 ( \14853 , \14852 );
or \U$14477 ( \14854 , \14840 , \14853 );
or \U$14478 ( \14855 , \14839 , \14852 );
nand \U$14479 ( \14856 , \14854 , \14855 );
not \U$14480 ( \14857 , \14856 );
or \U$14481 ( \14858 , \14834 , \14857 );
not \U$14482 ( \14859 , \14839 );
nand \U$14483 ( \14860 , \14859 , \14852 );
nand \U$14484 ( \14861 , \14858 , \14860 );
xnor \U$14485 ( \14862 , \14821 , \14861 );
not \U$14486 ( \14863 , \14862 );
or \U$14487 ( \14864 , \14819 , \14863 );
not \U$14488 ( \14865 , \14821 );
nand \U$14489 ( \14866 , \14865 , \14861 );
nand \U$14490 ( \14867 , \14864 , \14866 );
nand \U$14491 ( \14868 , \14813 , \14867 );
nand \U$14492 ( \14869 , \14808 , \14868 );
xor \U$14493 ( \14870 , \12952 , \12962 );
xor \U$14494 ( \14871 , \14870 , \12965 );
or \U$14495 ( \14872 , \14869 , \14871 );
not \U$14496 ( \14873 , \14872 );
xor \U$14497 ( \14874 , \14262 , \14223 );
xnor \U$14498 ( \14875 , \14874 , \14331 );
not \U$14499 ( \14876 , \14875 );
or \U$14500 ( \14877 , \14873 , \14876 );
nand \U$14501 ( \14878 , \14871 , \14869 );
nand \U$14502 ( \14879 , \14877 , \14878 );
nand \U$14503 ( \14880 , \14349 , \14879 );
or \U$14504 ( \14881 , \14340 , \14347 );
nand \U$14505 ( \14882 , \14880 , \14881 );
nor \U$14506 ( \14883 , \14222 , \14882 );
nor \U$14507 ( \14884 , \14220 , \14883 );
not \U$14508 ( \14885 , \14102 );
not \U$14509 ( \14886 , \14089 );
or \U$14510 ( \14887 , \14885 , \14886 );
nand \U$14511 ( \14888 , \14887 , \14092 );
not \U$14512 ( \14889 , \796 );
and \U$14513 ( \14890 , RIae78f80_134, \14148 );
not \U$14514 ( \14891 , RIae78f80_134);
and \U$14515 ( \14892 , \14891 , \10453 );
nor \U$14516 ( \14893 , \14890 , \14892 );
not \U$14517 ( \14894 , \14893 );
or \U$14518 ( \14895 , \14889 , \14894 );
and \U$14519 ( \14896 , \9412 , \1132 );
not \U$14520 ( \14897 , \9412 );
and \U$14521 ( \14898 , \14897 , RIae78f80_134);
nor \U$14522 ( \14899 , \14896 , \14898 );
nand \U$14523 ( \14900 , \14899 , \839 );
nand \U$14524 ( \14901 , \14895 , \14900 );
not \U$14525 ( \14902 , \9828 );
not \U$14526 ( \14903 , \14083 );
or \U$14527 ( \14904 , \14902 , \14903 );
and \U$14528 ( \14905 , RIae794a8_145, \5890 );
not \U$14529 ( \14906 , RIae794a8_145);
not \U$14530 ( \14907 , \2785 );
and \U$14531 ( \14908 , \14906 , \14907 );
or \U$14532 ( \14909 , \14905 , \14908 );
nand \U$14533 ( \14910 , \14909 , \1919 );
nand \U$14534 ( \14911 , \14904 , \14910 );
xor \U$14535 ( \14912 , \14901 , \14911 );
not \U$14536 ( \14913 , \9517 );
not \U$14537 ( \14914 , RIae79fe8_169);
not \U$14538 ( \14915 , \9624 );
or \U$14539 ( \14916 , \14914 , \14915 );
or \U$14540 ( \14917 , \2849 , RIae79fe8_169);
nand \U$14541 ( \14918 , \14916 , \14917 );
not \U$14542 ( \14919 , \14918 );
or \U$14543 ( \14920 , \14913 , \14919 );
nand \U$14544 ( \14921 , \14075 , \9499 );
nand \U$14545 ( \14922 , \14920 , \14921 );
xor \U$14546 ( \14923 , \14912 , \14922 );
not \U$14547 ( \14924 , \14923 );
not \U$14548 ( \14925 , \10637 );
not \U$14549 ( \14926 , \13745 );
or \U$14550 ( \14927 , \14925 , \14926 );
not \U$14551 ( \14928 , \10633 );
not \U$14552 ( \14929 , \1289 );
or \U$14553 ( \14930 , \14928 , \14929 );
not \U$14554 ( \14931 , RIae7a510_180);
or \U$14555 ( \14932 , \1289 , \14931 );
nand \U$14556 ( \14933 , \14930 , \14932 );
nand \U$14557 ( \14934 , \14933 , \10631 );
nand \U$14558 ( \14935 , \14927 , \14934 );
not \U$14559 ( \14936 , \6091 );
not \U$14560 ( \14937 , \14039 );
or \U$14561 ( \14938 , \14936 , \14937 );
xor \U$14562 ( \14939 , RIae79d90_164, \1897 );
buf \U$14563 ( \14940 , \5048 );
nand \U$14564 ( \14941 , \14939 , \14940 );
nand \U$14565 ( \14942 , \14938 , \14941 );
xor \U$14566 ( \14943 , \14935 , \14942 );
not \U$14567 ( \14944 , \11014 );
not \U$14568 ( \14945 , \14051 );
or \U$14569 ( \14946 , \14944 , \14945 );
and \U$14570 ( \14947 , RIae7a3a8_177, \936 );
not \U$14571 ( \14948 , RIae7a3a8_177);
and \U$14572 ( \14949 , \14948 , \937 );
or \U$14573 ( \14950 , \14947 , \14949 );
nand \U$14574 ( \14951 , \14950 , \9622 );
nand \U$14575 ( \14952 , \14946 , \14951 );
not \U$14576 ( \14953 , \14952 );
and \U$14577 ( \14954 , \14943 , \14953 );
not \U$14578 ( \14955 , \14943 );
and \U$14579 ( \14956 , \14955 , \14952 );
nor \U$14580 ( \14957 , \14954 , \14956 );
not \U$14581 ( \14958 , \14957 );
or \U$14582 ( \14959 , \14924 , \14958 );
or \U$14583 ( \14960 , \14923 , \14957 );
nand \U$14584 ( \14961 , \14959 , \14960 );
not \U$14585 ( \14962 , \13878 );
not \U$14586 ( \14963 , \13872 );
or \U$14587 ( \14964 , \14962 , \14963 );
nand \U$14588 ( \14965 , \13865 , \13871 );
nand \U$14589 ( \14966 , \14964 , \14965 );
xor \U$14590 ( \14967 , \14961 , \14966 );
xor \U$14591 ( \14968 , \14888 , \14967 );
not \U$14592 ( \14969 , \12680 );
not \U$14593 ( \14970 , \14063 );
or \U$14594 ( \14971 , \14969 , \14970 );
not \U$14595 ( \14972 , \12996 );
not \U$14596 ( \14973 , RIae79520_146);
and \U$14597 ( \14974 , \14972 , \14973 );
and \U$14598 ( \14975 , \14422 , RIae79520_146);
nor \U$14599 ( \14976 , \14974 , \14975 );
nand \U$14600 ( \14977 , \14976 , \10223 );
nand \U$14601 ( \14978 , \14971 , \14977 );
not \U$14602 ( \14979 , \14768 );
not \U$14603 ( \14980 , \13735 );
or \U$14604 ( \14981 , \14979 , \14980 );
not \U$14605 ( \14982 , RIae79ef8_167);
not \U$14606 ( \14983 , \3145 );
or \U$14607 ( \14984 , \14982 , \14983 );
or \U$14608 ( \14985 , \2047 , RIae79ef8_167);
nand \U$14609 ( \14986 , \14984 , \14985 );
nand \U$14610 ( \14987 , \14986 , \6214 );
nand \U$14611 ( \14988 , \14981 , \14987 );
xor \U$14612 ( \14989 , \14978 , \14988 );
not \U$14613 ( \14990 , \11087 );
not \U$14614 ( \14991 , \13755 );
or \U$14615 ( \14992 , \14990 , \14991 );
xor \U$14616 ( \14993 , RIae7a150_172, \11858 );
nand \U$14617 ( \14994 , \14993 , \9776 );
nand \U$14618 ( \14995 , \14992 , \14994 );
xor \U$14619 ( \14996 , \14989 , \14995 );
not \U$14620 ( \14997 , \2433 );
not \U$14621 ( \14998 , \13673 );
or \U$14622 ( \14999 , \14997 , \14998 );
not \U$14623 ( \15000 , RIae79778_151);
not \U$14624 ( \15001 , \2835 );
or \U$14625 ( \15002 , \15000 , \15001 );
or \U$14626 ( \15003 , \10534 , RIae79778_151);
nand \U$14627 ( \15004 , \15002 , \15003 );
nand \U$14628 ( \15005 , \15004 , \2450 );
nand \U$14629 ( \15006 , \14999 , \15005 );
not \U$14630 ( \15007 , \1989 );
not \U$14631 ( \15008 , \13685 );
or \U$14632 ( \15009 , \15007 , \15008 );
not \U$14633 ( \15010 , \1982 );
not \U$14634 ( \15011 , \1759 );
or \U$14635 ( \15012 , \15010 , \15011 );
nand \U$14636 ( \15013 , \1754 , RIae797f0_152);
nand \U$14637 ( \15014 , \15012 , \15013 );
nand \U$14638 ( \15015 , \15014 , \2519 );
nand \U$14639 ( \15016 , \15009 , \15015 );
xor \U$14640 ( \15017 , \15006 , \15016 );
not \U$14641 ( \15018 , \13130 );
not \U$14642 ( \15019 , \13717 );
or \U$14643 ( \15020 , \15018 , \15019 );
not \U$14644 ( \15021 , RIae7a240_174);
not \U$14645 ( \15022 , \2175 );
or \U$14646 ( \15023 , \15021 , \15022 );
or \U$14647 ( \15024 , \878 , RIae7a240_174);
nand \U$14648 ( \15025 , \15023 , \15024 );
nand \U$14649 ( \15026 , \15025 , \13121 );
nand \U$14650 ( \15027 , \15020 , \15026 );
xor \U$14651 ( \15028 , \15017 , \15027 );
xor \U$14652 ( \15029 , \14996 , \15028 );
not \U$14653 ( \15030 , \11364 );
and \U$14654 ( \15031 , RIae79c28_161, \2153 );
not \U$14655 ( \15032 , RIae79c28_161);
not \U$14656 ( \15033 , \2153 );
and \U$14657 ( \15034 , \15032 , \15033 );
or \U$14658 ( \15035 , \15031 , \15034 );
not \U$14659 ( \15036 , \15035 );
or \U$14660 ( \15037 , \15030 , \15036 );
nand \U$14661 ( \15038 , \13706 , \2767 );
nand \U$14662 ( \15039 , \15037 , \15038 );
not \U$14663 ( \15040 , \10696 );
not \U$14664 ( \15041 , \13694 );
or \U$14665 ( \15042 , \15040 , \15041 );
not \U$14666 ( \15043 , RIae7a498_179);
not \U$14667 ( \15044 , \780 );
or \U$14668 ( \15045 , \15043 , \15044 );
or \U$14669 ( \15046 , \1993 , RIae7a498_179);
nand \U$14670 ( \15047 , \15045 , \15046 );
nand \U$14671 ( \15048 , \15047 , \12371 );
nand \U$14672 ( \15049 , \15042 , \15048 );
xor \U$14673 ( \15050 , \15039 , \15049 );
not \U$14674 ( \15051 , \11761 );
not \U$14675 ( \15052 , \14027 );
or \U$14676 ( \15053 , \15051 , \15052 );
and \U$14677 ( \15054 , RIae79ca0_162, \9512 );
not \U$14678 ( \15055 , RIae79ca0_162);
and \U$14679 ( \15056 , \15055 , \2993 );
nor \U$14680 ( \15057 , \15054 , \15056 );
nand \U$14681 ( \15058 , \15057 , \4853 );
nand \U$14682 ( \15059 , \15053 , \15058 );
xor \U$14683 ( \15060 , \15050 , \15059 );
xnor \U$14684 ( \15061 , \15029 , \15060 );
xnor \U$14685 ( \15062 , \14968 , \15061 );
not \U$14686 ( \15063 , \13960 );
not \U$14687 ( \15064 , \14009 );
or \U$14688 ( \15065 , \15063 , \15064 );
not \U$14689 ( \15066 , \14007 );
nand \U$14690 ( \15067 , \15066 , \13969 );
nand \U$14691 ( \15068 , \15065 , \15067 );
not \U$14692 ( \15069 , \13688 );
not \U$14693 ( \15070 , \13760 );
or \U$14694 ( \15071 , \15069 , \15070 );
nand \U$14695 ( \15072 , \15071 , \13727 );
or \U$14696 ( \15073 , \13688 , \13760 );
and \U$14697 ( \15074 , \15072 , \15073 );
xor \U$14698 ( \15075 , \15068 , \15074 );
not \U$14699 ( \15076 , \1062 );
not \U$14700 ( \15077 , \14160 );
or \U$14701 ( \15078 , \15076 , \15077 );
not \U$14702 ( \15079 , RIae79070_136);
not \U$14703 ( \15080 , \14657 );
or \U$14704 ( \15081 , \15079 , \15080 );
or \U$14705 ( \15082 , \9456 , RIae79070_136);
nand \U$14706 ( \15083 , \15081 , \15082 );
nand \U$14707 ( \15084 , \15083 , \9947 );
nand \U$14708 ( \15085 , \15078 , \15084 );
not \U$14709 ( \15086 , \10451 );
not \U$14710 ( \15087 , \6414 );
not \U$14711 ( \15088 , \13287 );
not \U$14712 ( \15089 , \15088 );
or \U$14713 ( \15090 , \15087 , \15089 );
buf \U$14714 ( \15091 , \9367 );
or \U$14715 ( \15092 , \15091 , \6414 );
nand \U$14716 ( \15093 , \15090 , \15092 );
not \U$14717 ( \15094 , \15093 );
or \U$14718 ( \15095 , \15086 , \15094 );
nand \U$14719 ( \15096 , \1008 , \14114 );
nand \U$14720 ( \15097 , \15095 , \15096 );
xor \U$14721 ( \15098 , \15085 , \15097 );
not \U$14722 ( \15099 , \9403 );
not \U$14723 ( \15100 , \14134 );
or \U$14724 ( \15101 , \15099 , \15100 );
not \U$14725 ( \15102 , \9313 );
and \U$14726 ( \15103 , RIae79250_140, \15102 );
not \U$14727 ( \15104 , RIae79250_140);
and \U$14728 ( \15105 , \15104 , \9316 );
or \U$14729 ( \15106 , \15103 , \15105 );
not \U$14730 ( \15107 , \15106 );
nand \U$14731 ( \15108 , \15107 , \1501 );
nand \U$14732 ( \15109 , \15101 , \15108 );
xor \U$14733 ( \15110 , \15098 , \15109 );
or \U$14734 ( \15111 , \13725 , \13709 );
nand \U$14735 ( \15112 , \15111 , \13711 );
xor \U$14736 ( \15113 , \15110 , \15112 );
not \U$14737 ( \15114 , \1910 );
not \U$14738 ( \15115 , \14124 );
or \U$14739 ( \15116 , \15114 , \15115 );
not \U$14740 ( \15117 , \6345 );
and \U$14741 ( \15118 , \15117 , \1902 );
not \U$14742 ( \15119 , \15117 );
and \U$14743 ( \15120 , \15119 , RIae793b8_143);
nor \U$14744 ( \15121 , \15118 , \15120 );
nand \U$14745 ( \15122 , \15121 , \1864 );
nand \U$14746 ( \15123 , \15116 , \15122 );
not \U$14747 ( \15124 , \2011 );
not \U$14748 ( \15125 , RIae79610_148);
not \U$14749 ( \15126 , \10237 );
or \U$14750 ( \15127 , \15125 , \15126 );
not \U$14751 ( \15128 , \6256 );
or \U$14752 ( \15129 , \15128 , RIae79610_148);
nand \U$14753 ( \15130 , \15127 , \15129 );
not \U$14754 ( \15131 , \15130 );
or \U$14755 ( \15132 , \15124 , \15131 );
nand \U$14756 ( \15133 , \13978 , \2063 );
nand \U$14757 ( \15134 , \15132 , \15133 );
xor \U$14758 ( \15135 , \15123 , \15134 );
not \U$14759 ( \15136 , \1843 );
not \U$14760 ( \15137 , \13988 );
or \U$14761 ( \15138 , \15136 , \15137 );
not \U$14762 ( \15139 , RIae79688_149);
not \U$14763 ( \15140 , \6242 );
or \U$14764 ( \15141 , \15139 , \15140 );
not \U$14765 ( \15142 , RIae79688_149);
nand \U$14766 ( \15143 , \15142 , \4169 );
nand \U$14767 ( \15144 , \15141 , \15143 );
nand \U$14768 ( \15145 , \15144 , \1821 );
nand \U$14769 ( \15146 , \15138 , \15145 );
xor \U$14770 ( \15147 , \15135 , \15146 );
xor \U$14771 ( \15148 , \15113 , \15147 );
xor \U$14772 ( \15149 , \15075 , \15148 );
not \U$14773 ( \15150 , \14019 );
not \U$14774 ( \15151 , \14014 );
nand \U$14775 ( \15152 , \15150 , \15151 );
not \U$14776 ( \15153 , \15152 );
not \U$14777 ( \15154 , \14106 );
or \U$14778 ( \15155 , \15153 , \15154 );
not \U$14779 ( \15156 , \15151 );
nand \U$14780 ( \15157 , \15156 , \14019 );
nand \U$14781 ( \15158 , \15155 , \15157 );
nor \U$14782 ( \15159 , \15149 , \15158 );
or \U$14783 ( \15160 , \15062 , \15159 );
nand \U$14784 ( \15161 , \15149 , \15158 );
nand \U$14785 ( \15162 , \15160 , \15161 );
not \U$14786 ( \15163 , \14042 );
not \U$14787 ( \15164 , \14031 );
not \U$14788 ( \15165 , \15164 );
or \U$14789 ( \15166 , \15163 , \15165 );
not \U$14790 ( \15167 , \14041 );
not \U$14791 ( \15168 , \14031 );
or \U$14792 ( \15169 , \15167 , \15168 );
nand \U$14793 ( \15170 , \15169 , \14056 );
nand \U$14794 ( \15171 , \15166 , \15170 );
not \U$14795 ( \15172 , \15171 );
not \U$14796 ( \15173 , \15172 );
xor \U$14797 ( \15174 , \14067 , \14077 );
and \U$14798 ( \15175 , \15174 , \14087 );
and \U$14799 ( \15176 , \14067 , \14077 );
or \U$14800 ( \15177 , \15175 , \15176 );
not \U$14801 ( \15178 , \15177 );
or \U$14802 ( \15179 , \15173 , \15178 );
not \U$14803 ( \15180 , \15177 );
not \U$14804 ( \15181 , \15180 );
not \U$14805 ( \15182 , \15171 );
or \U$14806 ( \15183 , \15181 , \15182 );
xor \U$14807 ( \15184 , \13739 , \13749 );
and \U$14808 ( \15185 , \15184 , \13759 );
and \U$14809 ( \15186 , \13739 , \13749 );
or \U$14810 ( \15187 , \15185 , \15186 );
nand \U$14811 ( \15188 , \15183 , \15187 );
nand \U$14812 ( \15189 , \15179 , \15188 );
xor \U$14813 ( \15190 , \15110 , \15112 );
and \U$14814 ( \15191 , \15190 , \15147 );
and \U$14815 ( \15192 , \15110 , \15112 );
or \U$14816 ( \15193 , \15191 , \15192 );
xor \U$14817 ( \15194 , \15189 , \15193 );
xor \U$14818 ( \15195 , \14978 , \14988 );
and \U$14819 ( \15196 , \15195 , \14995 );
and \U$14820 ( \15197 , \14978 , \14988 );
or \U$14821 ( \15198 , \15196 , \15197 );
xor \U$14822 ( \15199 , \14901 , \14911 );
and \U$14823 ( \15200 , \15199 , \14922 );
and \U$14824 ( \15201 , \14901 , \14911 );
or \U$14825 ( \15202 , \15200 , \15201 );
xor \U$14826 ( \15203 , \15198 , \15202 );
not \U$14827 ( \15204 , \1910 );
not \U$14828 ( \15205 , \15121 );
or \U$14829 ( \15206 , \15204 , \15205 );
not \U$14830 ( \15207 , \5722 );
and \U$14831 ( \15208 , RIae793b8_143, \15207 );
not \U$14832 ( \15209 , RIae793b8_143);
and \U$14833 ( \15210 , \15209 , \5722 );
or \U$14834 ( \15211 , \15208 , \15210 );
nand \U$14835 ( \15212 , \15211 , \1864 );
nand \U$14836 ( \15213 , \15206 , \15212 );
not \U$14837 ( \15214 , \15106 );
not \U$14838 ( \15215 , \1498 );
and \U$14839 ( \15216 , \15214 , \15215 );
buf \U$14840 ( \15217 , \12056 );
and \U$14841 ( \15218 , RIae79250_140, \15217 );
not \U$14842 ( \15219 , RIae79250_140);
not \U$14843 ( \15220 , \12687 );
and \U$14844 ( \15221 , \15219 , \15220 );
or \U$14845 ( \15222 , \15218 , \15221 );
and \U$14846 ( \15223 , \15222 , \1501 );
nor \U$14847 ( \15224 , \15216 , \15223 );
not \U$14848 ( \15225 , \15224 );
xor \U$14849 ( \15226 , \15213 , \15225 );
not \U$14850 ( \15227 , \2011 );
not \U$14851 ( \15228 , RIae79610_148);
not \U$14852 ( \15229 , \10829 );
or \U$14853 ( \15230 , \15228 , \15229 );
or \U$14854 ( \15231 , \10829 , RIae79610_148);
nand \U$14855 ( \15232 , \15230 , \15231 );
not \U$14856 ( \15233 , \15232 );
or \U$14857 ( \15234 , \15227 , \15233 );
nand \U$14858 ( \15235 , \15130 , \2063 );
nand \U$14859 ( \15236 , \15234 , \15235 );
xor \U$14860 ( \15237 , \15226 , \15236 );
xor \U$14861 ( \15238 , \15203 , \15237 );
xor \U$14862 ( \15239 , \15194 , \15238 );
xor \U$14863 ( \15240 , \15068 , \15074 );
and \U$14864 ( \15241 , \15240 , \15148 );
and \U$14865 ( \15242 , \15068 , \15074 );
or \U$14866 ( \15243 , \15241 , \15242 );
xor \U$14867 ( \15244 , \15239 , \15243 );
not \U$14868 ( \15245 , \15187 );
xor \U$14869 ( \15246 , \15172 , \15180 );
not \U$14870 ( \15247 , \15246 );
or \U$14871 ( \15248 , \15245 , \15247 );
not \U$14872 ( \15249 , \15246 );
not \U$14873 ( \15250 , \15187 );
nand \U$14874 ( \15251 , \15249 , \15250 );
nand \U$14875 ( \15252 , \15248 , \15251 );
not \U$14876 ( \15253 , \15252 );
not \U$14877 ( \15254 , \13915 );
not \U$14878 ( \15255 , \15254 );
not \U$14879 ( \15256 , \13889 );
or \U$14880 ( \15257 , \15255 , \15256 );
not \U$14881 ( \15258 , \13914 );
nand \U$14882 ( \15259 , \15258 , \13911 );
nand \U$14883 ( \15260 , \15257 , \15259 );
not \U$14884 ( \15261 , \13819 );
not \U$14885 ( \15262 , \13839 );
or \U$14886 ( \15263 , \15261 , \15262 );
or \U$14887 ( \15264 , \13819 , \13839 );
not \U$14888 ( \15265 , \13037 );
not \U$14889 ( \15266 , \13825 );
or \U$14890 ( \15267 , \15265 , \15266 );
nand \U$14891 ( \15268 , \15267 , \13828 );
nand \U$14892 ( \15269 , \15264 , \15268 );
nand \U$14893 ( \15270 , \15263 , \15269 );
xor \U$14894 ( \15271 , \15260 , \15270 );
not \U$14895 ( \15272 , \15271 );
or \U$14896 ( \15273 , \15253 , \15272 );
buf \U$14897 ( \15274 , \15270 );
nand \U$14898 ( \15275 , \15274 , \15260 );
nand \U$14899 ( \15276 , \15273 , \15275 );
xor \U$14900 ( \15277 , \15244 , \15276 );
xor \U$14901 ( \15278 , \15162 , \15277 );
xor \U$14902 ( \15279 , \15039 , \15049 );
and \U$14903 ( \15280 , \15279 , \15059 );
and \U$14904 ( \15281 , \15039 , \15049 );
or \U$14905 ( \15282 , \15280 , \15281 );
xor \U$14906 ( \15283 , \15006 , \15016 );
and \U$14907 ( \15284 , \15283 , \15027 );
and \U$14908 ( \15285 , \15006 , \15016 );
or \U$14909 ( \15286 , \15284 , \15285 );
not \U$14910 ( \15287 , \15286 );
and \U$14911 ( \15288 , \15282 , \15287 );
not \U$14912 ( \15289 , \15282 );
and \U$14913 ( \15290 , \15289 , \15286 );
nor \U$14914 ( \15291 , \15288 , \15290 );
not \U$14915 ( \15292 , \14942 );
not \U$14916 ( \15293 , \15292 );
not \U$14917 ( \15294 , \14953 );
or \U$14918 ( \15295 , \15293 , \15294 );
not \U$14919 ( \15296 , \14942 );
not \U$14920 ( \15297 , \14952 );
or \U$14921 ( \15298 , \15296 , \15297 );
not \U$14922 ( \15299 , \14935 );
nand \U$14923 ( \15300 , \15298 , \15299 );
nand \U$14924 ( \15301 , \15295 , \15300 );
and \U$14925 ( \15302 , \15291 , \15301 );
not \U$14926 ( \15303 , \15291 );
not \U$14927 ( \15304 , \15301 );
and \U$14928 ( \15305 , \15303 , \15304 );
nor \U$14929 ( \15306 , \15302 , \15305 );
not \U$14930 ( \15307 , \14966 );
not \U$14931 ( \15308 , \14961 );
or \U$14932 ( \15309 , \15307 , \15308 );
not \U$14933 ( \15310 , \14957 );
nand \U$14934 ( \15311 , \15310 , \14923 );
nand \U$14935 ( \15312 , \15309 , \15311 );
and \U$14936 ( \15313 , \15306 , \15312 );
not \U$14937 ( \15314 , \15306 );
not \U$14938 ( \15315 , \15312 );
and \U$14939 ( \15316 , \15314 , \15315 );
nor \U$14940 ( \15317 , \15313 , \15316 );
not \U$14941 ( \15318 , \9814 );
xor \U$14942 ( \15319 , RIae7a2b8_175, \2917 );
not \U$14943 ( \15320 , \15319 );
or \U$14944 ( \15321 , \15318 , \15320 );
not \U$14945 ( \15322 , RIae7a2b8_175);
not \U$14946 ( \15323 , \975 );
or \U$14947 ( \15324 , \15322 , \15323 );
or \U$14948 ( \15325 , \14778 , RIae7a2b8_175);
nand \U$14949 ( \15326 , \15324 , \15325 );
nand \U$14950 ( \15327 , \15326 , \9792 );
nand \U$14951 ( \15328 , \15321 , \15327 );
not \U$14952 ( \15329 , \2432 );
not \U$14953 ( \15330 , \15004 );
or \U$14954 ( \15331 , \15329 , \15330 );
not \U$14955 ( \15332 , \2447 );
not \U$14956 ( \15333 , \2309 );
or \U$14957 ( \15334 , \15332 , \15333 );
or \U$14958 ( \15335 , \2309 , \2447 );
nand \U$14959 ( \15336 , \15334 , \15335 );
buf \U$14960 ( \15337 , \2450 );
nand \U$14961 ( \15338 , \15336 , \15337 );
nand \U$14962 ( \15339 , \15331 , \15338 );
not \U$14963 ( \15340 , \15339 );
not \U$14964 ( \15341 , \2007 );
not \U$14965 ( \15342 , \2521 );
not \U$14966 ( \15343 , \6171 );
or \U$14967 ( \15344 , \15342 , \15343 );
nand \U$14968 ( \15345 , \2857 , RIae797f0_152);
nand \U$14969 ( \15346 , \15344 , \15345 );
not \U$14970 ( \15347 , \15346 );
or \U$14971 ( \15348 , \15341 , \15347 );
nand \U$14972 ( \15349 , \15014 , \1988 );
nand \U$14973 ( \15350 , \15348 , \15349 );
not \U$14974 ( \15351 , \15350 );
not \U$14975 ( \15352 , \15351 );
or \U$14976 ( \15353 , \15340 , \15352 );
or \U$14977 ( \15354 , \15351 , \15339 );
nand \U$14978 ( \15355 , \15353 , \15354 );
xor \U$14979 ( \15356 , \15328 , \15355 );
not \U$14980 ( \15357 , \3014 );
not \U$14981 ( \15358 , RIae79ac0_158);
not \U$14982 ( \15359 , \1859 );
or \U$14983 ( \15360 , \15358 , \15359 );
or \U$14984 ( \15361 , \1859 , RIae79ac0_158);
nand \U$14985 ( \15362 , \15360 , \15361 );
not \U$14986 ( \15363 , \15362 );
or \U$14987 ( \15364 , \15357 , \15363 );
and \U$14988 ( \15365 , RIae79ac0_158, \2402 );
not \U$14989 ( \15366 , RIae79ac0_158);
and \U$14990 ( \15367 , \15366 , \3273 );
or \U$14991 ( \15368 , \15365 , \15367 );
nand \U$14992 ( \15369 , \15368 , \2272 );
nand \U$14993 ( \15370 , \15364 , \15369 );
not \U$14994 ( \15371 , \2163 );
not \U$14995 ( \15372 , RIae79520_146);
not \U$14996 ( \15373 , \2357 );
or \U$14997 ( \15374 , \15372 , \15373 );
or \U$14998 ( \15375 , \4112 , RIae79520_146);
nand \U$14999 ( \15376 , \15374 , \15375 );
not \U$15000 ( \15377 , \15376 );
or \U$15001 ( \15378 , \15371 , \15377 );
nand \U$15002 ( \15379 , \5950 , \14976 );
nand \U$15003 ( \15380 , \15378 , \15379 );
xor \U$15004 ( \15381 , \15370 , \15380 );
buf \U$15005 ( \15382 , \10696 );
not \U$15006 ( \15383 , \15382 );
not \U$15007 ( \15384 , \15047 );
or \U$15008 ( \15385 , \15383 , \15384 );
and \U$15009 ( \15386 , RIae7a498_179, \12522 );
not \U$15010 ( \15387 , RIae7a498_179);
and \U$15011 ( \15388 , \15387 , \827 );
nor \U$15012 ( \15389 , \15386 , \15388 );
nand \U$15013 ( \15390 , \15389 , \12371 );
nand \U$15014 ( \15391 , \15385 , \15390 );
xor \U$15015 ( \15392 , \15381 , \15391 );
xor \U$15016 ( \15393 , \15356 , \15392 );
not \U$15017 ( \15394 , \11364 );
not \U$15018 ( \15395 , RIae79c28_161);
not \U$15019 ( \15396 , \10570 );
or \U$15020 ( \15397 , \15395 , \15396 );
nand \U$15021 ( \15398 , \10567 , \10584 );
nand \U$15022 ( \15399 , \15397 , \15398 );
not \U$15023 ( \15400 , \15399 );
or \U$15024 ( \15401 , \15394 , \15400 );
nand \U$15025 ( \15402 , \15035 , \2767 );
nand \U$15026 ( \15403 , \15401 , \15402 );
not \U$15027 ( \15404 , \10631 );
xor \U$15028 ( \15405 , RIae7a510_180, \2323 );
not \U$15029 ( \15406 , \15405 );
or \U$15030 ( \15407 , \15404 , \15406 );
nand \U$15031 ( \15408 , \14933 , \10927 );
nand \U$15032 ( \15409 , \15407 , \15408 );
and \U$15033 ( \15410 , \15403 , \15409 );
not \U$15034 ( \15411 , \15403 );
not \U$15035 ( \15412 , \15409 );
and \U$15036 ( \15413 , \15411 , \15412 );
nor \U$15037 ( \15414 , \15410 , \15413 );
not \U$15038 ( \15415 , \13121 );
xor \U$15039 ( \15416 , \854 , RIae7a240_174);
not \U$15040 ( \15417 , \15416 );
or \U$15041 ( \15418 , \15415 , \15417 );
nand \U$15042 ( \15419 , \15025 , \13130 );
nand \U$15043 ( \15420 , \15418 , \15419 );
xor \U$15044 ( \15421 , \15414 , \15420 );
xor \U$15045 ( \15422 , \15393 , \15421 );
xnor \U$15046 ( \15423 , \15317 , \15422 );
not \U$15047 ( \15424 , \15423 );
not \U$15048 ( \15425 , \14888 );
nor \U$15049 ( \15426 , \15425 , \14967 );
or \U$15050 ( \15427 , \15426 , \15061 );
nand \U$15051 ( \15428 , \15425 , \14967 );
nand \U$15052 ( \15429 , \15427 , \15428 );
not \U$15053 ( \15430 , \15429 );
not \U$15054 ( \15431 , \13677 );
nand \U$15055 ( \15432 , \15431 , \13667 );
and \U$15056 ( \15433 , \15432 , \13687 );
not \U$15057 ( \15434 , \13667 );
and \U$15058 ( \15435 , \13677 , \15434 );
nor \U$15059 ( \15436 , \15433 , \15435 );
xor \U$15060 ( \15437 , \13938 , \13948 );
and \U$15061 ( \15438 , \15437 , \13959 );
and \U$15062 ( \15439 , \13938 , \13948 );
or \U$15063 ( \15440 , \15438 , \15439 );
not \U$15064 ( \15441 , \15440 );
xor \U$15065 ( \15442 , \15436 , \15441 );
not \U$15066 ( \15443 , \9792 );
not \U$15067 ( \15444 , \13955 );
or \U$15068 ( \15445 , \15443 , \15444 );
nand \U$15069 ( \15446 , \15326 , \9814 );
nand \U$15070 ( \15447 , \15445 , \15446 );
not \U$15071 ( \15448 , \2322 );
not \U$15072 ( \15449 , RIae798e0_154);
not \U$15073 ( \15450 , \11681 );
or \U$15074 ( \15451 , \15449 , \15450 );
or \U$15075 ( \15452 , \1789 , RIae798e0_154);
nand \U$15076 ( \15453 , \15451 , \15452 );
not \U$15077 ( \15454 , \15453 );
or \U$15078 ( \15455 , \15448 , \15454 );
nand \U$15079 ( \15456 , \13944 , \14580 );
nand \U$15080 ( \15457 , \15455 , \15456 );
and \U$15081 ( \15458 , \15457 , \13667 );
not \U$15082 ( \15459 , \15457 );
and \U$15083 ( \15460 , \15459 , \15434 );
nor \U$15084 ( \15461 , \15458 , \15460 );
xnor \U$15085 ( \15462 , \15447 , \15461 );
and \U$15086 ( \15463 , \15442 , \15462 );
and \U$15087 ( \15464 , \15436 , \15441 );
or \U$15088 ( \15465 , \15463 , \15464 );
not \U$15089 ( \15466 , \15465 );
not \U$15090 ( \15467 , \14996 );
not \U$15091 ( \15468 , \15060 );
or \U$15092 ( \15469 , \15467 , \15468 );
or \U$15093 ( \15470 , \15060 , \14996 );
nand \U$15094 ( \15471 , \15470 , \15028 );
nand \U$15095 ( \15472 , \15469 , \15471 );
not \U$15096 ( \15473 , \15472 );
or \U$15097 ( \15474 , \15466 , \15473 );
or \U$15098 ( \15475 , \15472 , \15465 );
nand \U$15099 ( \15476 , \15474 , \15475 );
not \U$15100 ( \15477 , \10573 );
not \U$15101 ( \15478 , RIae79ef8_167);
not \U$15102 ( \15479 , \12183 );
or \U$15103 ( \15480 , \15478 , \15479 );
nand \U$15104 ( \15481 , \2031 , \12209 );
nand \U$15105 ( \15482 , \15480 , \15481 );
not \U$15106 ( \15483 , \15482 );
or \U$15107 ( \15484 , \15477 , \15483 );
nand \U$15108 ( \15485 , \14986 , \6201 );
nand \U$15109 ( \15486 , \15484 , \15485 );
not \U$15110 ( \15487 , \839 );
not \U$15111 ( \15488 , \10936 );
and \U$15112 ( \15489 , \15488 , \1132 );
not \U$15113 ( \15490 , \15488 );
and \U$15114 ( \15491 , \15490 , RIae78f80_134);
nor \U$15115 ( \15492 , \15489 , \15491 );
not \U$15116 ( \15493 , \15492 );
or \U$15117 ( \15494 , \15487 , \15493 );
nand \U$15118 ( \15495 , \14899 , \796 );
nand \U$15119 ( \15496 , \15494 , \15495 );
not \U$15120 ( \15497 , \1072 );
xor \U$15121 ( \15498 , RIae78e90_132, \12482 );
not \U$15122 ( \15499 , \15498 );
or \U$15123 ( \15500 , \15497 , \15499 );
buf \U$15124 ( \15501 , \9941 );
and \U$15125 ( \15502 , \921 , \15501 );
not \U$15126 ( \15503 , \921 );
not \U$15127 ( \15504 , \10461 );
and \U$15128 ( \15505 , \15503 , \15504 );
nor \U$15129 ( \15506 , \15502 , \15505 );
nand \U$15130 ( \15507 , \15506 , \5858 );
nand \U$15131 ( \15508 , \15500 , \15507 );
xor \U$15132 ( \15509 , \15496 , \15508 );
xor \U$15133 ( \15510 , \15486 , \15509 );
not \U$15134 ( \15511 , \15510 );
xor \U$15135 ( \15512 , RIae79070_136, \9438 );
not \U$15136 ( \15513 , \15512 );
not \U$15137 ( \15514 , \1049 );
or \U$15138 ( \15515 , \15513 , \15514 );
nand \U$15139 ( \15516 , \15083 , \1062 );
nand \U$15140 ( \15517 , \15515 , \15516 );
not \U$15141 ( \15518 , \1209 );
not \U$15142 ( \15519 , \9347 );
not \U$15143 ( \15520 , \15519 );
and \U$15144 ( \15521 , \15520 , \997 );
not \U$15145 ( \15522 , \15520 );
and \U$15146 ( \15523 , \15522 , RIae79160_138);
nor \U$15147 ( \15524 , \15521 , \15523 );
not \U$15148 ( \15525 , \15524 );
or \U$15149 ( \15526 , \15518 , \15525 );
nand \U$15150 ( \15527 , \15093 , \1008 );
nand \U$15151 ( \15528 , \15526 , \15527 );
xor \U$15152 ( \15529 , \15517 , \15528 );
not \U$15153 ( \15530 , \10667 );
not \U$15154 ( \15531 , \14993 );
or \U$15155 ( \15532 , \15530 , \15531 );
nand \U$15156 ( \15533 , \9776 , RIae7a150_172);
nand \U$15157 ( \15534 , \15532 , \15533 );
buf \U$15158 ( \15535 , \15534 );
xnor \U$15159 ( \15536 , \15529 , \15535 );
not \U$15160 ( \15537 , \15536 );
or \U$15161 ( \15538 , \15511 , \15537 );
or \U$15162 ( \15539 , \15536 , \15510 );
nand \U$15163 ( \15540 , \15538 , \15539 );
not \U$15164 ( \15541 , \15447 );
not \U$15165 ( \15542 , \15461 );
or \U$15166 ( \15543 , \15541 , \15542 );
nand \U$15167 ( \15544 , \15457 , \13667 );
nand \U$15168 ( \15545 , \15543 , \15544 );
xnor \U$15169 ( \15546 , \15540 , \15545 );
not \U$15170 ( \15547 , \15546 );
xnor \U$15171 ( \15548 , \15476 , \15547 );
not \U$15172 ( \15549 , \15548 );
or \U$15173 ( \15550 , \15430 , \15549 );
or \U$15174 ( \15551 , \15429 , \15548 );
nand \U$15175 ( \15552 , \15550 , \15551 );
not \U$15176 ( \15553 , \15552 );
or \U$15177 ( \15554 , \15424 , \15553 );
or \U$15178 ( \15555 , \15423 , \15552 );
nand \U$15179 ( \15556 , \15554 , \15555 );
xor \U$15180 ( \15557 , \15278 , \15556 );
xor \U$15181 ( \15558 , \13790 , \13933 );
and \U$15182 ( \15559 , \15558 , \14203 );
and \U$15183 ( \15560 , \13790 , \13933 );
or \U$15184 ( \15561 , \15559 , \15560 );
not \U$15185 ( \15562 , \15561 );
not \U$15186 ( \15563 , \13781 );
and \U$15187 ( \15564 , \13774 , \13640 );
not \U$15188 ( \15565 , \13774 );
not \U$15189 ( \15566 , \13640 );
and \U$15190 ( \15567 , \15565 , \15566 );
nor \U$15191 ( \15568 , \15564 , \15567 );
not \U$15192 ( \15569 , \15568 );
or \U$15193 ( \15570 , \15563 , \15569 );
nand \U$15194 ( \15571 , \13640 , \13774 );
nand \U$15195 ( \15572 , \15570 , \15571 );
not \U$15196 ( \15573 , \15572 );
xor \U$15197 ( \15574 , \15436 , \15441 );
xor \U$15198 ( \15575 , \15574 , \15462 );
not \U$15199 ( \15576 , \14172 );
not \U$15200 ( \15577 , \15576 );
not \U$15201 ( \15578 , \14185 );
or \U$15202 ( \15579 , \15577 , \15578 );
or \U$15203 ( \15580 , \14185 , \15576 );
nand \U$15204 ( \15581 , \15580 , \14179 );
nand \U$15205 ( \15582 , \15579 , \15581 );
xor \U$15206 ( \15583 , \15575 , \15582 );
not \U$15207 ( \15584 , \13923 );
not \U$15208 ( \15585 , \15584 );
not \U$15209 ( \15586 , \13860 );
or \U$15210 ( \15587 , \15585 , \15586 );
not \U$15211 ( \15588 , \13883 );
nand \U$15212 ( \15589 , \15588 , \13919 );
nand \U$15213 ( \15590 , \15587 , \15589 );
xor \U$15214 ( \15591 , \15583 , \15590 );
not \U$15215 ( \15592 , \15591 );
not \U$15216 ( \15593 , \13797 );
not \U$15217 ( \15594 , \13849 );
or \U$15218 ( \15595 , \15593 , \15594 );
nand \U$15219 ( \15596 , \15595 , \13927 );
nand \U$15220 ( \15597 , \15596 , \13854 );
nand \U$15221 ( \15598 , \13772 , \13647 );
not \U$15222 ( \15599 , \13653 );
not \U$15223 ( \15600 , \13766 );
or \U$15224 ( \15601 , \15599 , \15600 );
nand \U$15225 ( \15602 , \15601 , \13770 );
nand \U$15226 ( \15603 , \15598 , \15602 );
xor \U$15227 ( \15604 , \15597 , \15603 );
not \U$15228 ( \15605 , \15604 );
or \U$15229 ( \15606 , \15592 , \15605 );
or \U$15230 ( \15607 , \15591 , \15604 );
nand \U$15231 ( \15608 , \15606 , \15607 );
not \U$15232 ( \15609 , \15608 );
not \U$15233 ( \15610 , \15609 );
or \U$15234 ( \15611 , \15573 , \15610 );
not \U$15235 ( \15612 , \15572 );
nand \U$15236 ( \15613 , \15612 , \15608 );
nand \U$15237 ( \15614 , \15611 , \15613 );
not \U$15238 ( \15615 , \15614 );
or \U$15239 ( \15616 , \15562 , \15615 );
not \U$15240 ( \15617 , \15609 );
buf \U$15241 ( \15618 , \15572 );
nand \U$15242 ( \15619 , \15617 , \15618 );
nand \U$15243 ( \15620 , \15616 , \15619 );
xor \U$15244 ( \15621 , \15557 , \15620 );
not \U$15245 ( \15622 , \9518 );
not \U$15246 ( \15623 , RIae79fe8_169);
not \U$15247 ( \15624 , \1186 );
or \U$15248 ( \15625 , \15623 , \15624 );
or \U$15249 ( \15626 , \11538 , RIae79fe8_169);
nand \U$15250 ( \15627 , \15625 , \15626 );
not \U$15251 ( \15628 , \15627 );
or \U$15252 ( \15629 , \15622 , \15628 );
nand \U$15253 ( \15630 , \14918 , \9499 );
nand \U$15254 ( \15631 , \15629 , \15630 );
not \U$15255 ( \15632 , \2322 );
and \U$15256 ( \15633 , RIae798e0_154, \1809 );
not \U$15257 ( \15634 , RIae798e0_154);
and \U$15258 ( \15635 , \15634 , \3529 );
or \U$15259 ( \15636 , \15633 , \15635 );
not \U$15260 ( \15637 , \15636 );
or \U$15261 ( \15638 , \15632 , \15637 );
nand \U$15262 ( \15639 , \15453 , \2340 );
nand \U$15263 ( \15640 , \15638 , \15639 );
not \U$15264 ( \15641 , \927 );
not \U$15265 ( \15642 , RIae78bc0_126);
not \U$15266 ( \15643 , \13657 );
or \U$15267 ( \15644 , \15642 , \15643 );
nand \U$15268 ( \15645 , \12644 , \1286 );
nand \U$15269 ( \15646 , \15644 , \15645 );
not \U$15270 ( \15647 , \15646 );
or \U$15271 ( \15648 , \15641 , \15647 );
not \U$15272 ( \15649 , \1286 );
not \U$15273 ( \15650 , \10084 );
not \U$15274 ( \15651 , \15650 );
or \U$15275 ( \15652 , \15649 , \15651 );
not \U$15276 ( \15653 , \10207 );
nand \U$15277 ( \15654 , \15653 , RIae78bc0_126);
nand \U$15278 ( \15655 , \15652 , \15654 );
nand \U$15279 ( \15656 , \15655 , \951 );
nand \U$15280 ( \15657 , \15648 , \15656 );
and \U$15281 ( \15658 , \15640 , \15657 );
not \U$15282 ( \15659 , \15640 );
not \U$15283 ( \15660 , \15657 );
and \U$15284 ( \15661 , \15659 , \15660 );
or \U$15285 ( \15662 , \15658 , \15661 );
xor \U$15286 ( \15663 , \15631 , \15662 );
not \U$15287 ( \15664 , \5048 );
not \U$15288 ( \15665 , \1878 );
xor \U$15289 ( \15666 , RIae79d90_164, \15665 );
not \U$15290 ( \15667 , \15666 );
or \U$15291 ( \15668 , \15664 , \15667 );
nand \U$15292 ( \15669 , \14939 , \6091 );
nand \U$15293 ( \15670 , \15668 , \15669 );
not \U$15294 ( \15671 , \9622 );
and \U$15295 ( \15672 , \911 , \913 );
not \U$15296 ( \15673 , \911 );
and \U$15297 ( \15674 , \15673 , \912 );
nor \U$15298 ( \15675 , \15672 , \15674 );
and \U$15299 ( \15676 , RIae7a3a8_177, \15675 );
not \U$15300 ( \15677 , RIae7a3a8_177);
and \U$15301 ( \15678 , \15677 , \10662 );
nor \U$15302 ( \15679 , \15676 , \15678 );
not \U$15303 ( \15680 , \15679 );
or \U$15304 ( \15681 , \15671 , \15680 );
nand \U$15305 ( \15682 , \14950 , \9644 );
nand \U$15306 ( \15683 , \15681 , \15682 );
xor \U$15307 ( \15684 , \15670 , \15683 );
not \U$15308 ( \15685 , \4853 );
xnor \U$15309 ( \15686 , \12207 , RIae79ca0_162);
not \U$15310 ( \15687 , \15686 );
or \U$15311 ( \15688 , \15685 , \15687 );
nand \U$15312 ( \15689 , \15057 , \4842 );
nand \U$15313 ( \15690 , \15688 , \15689 );
xor \U$15314 ( \15691 , \15684 , \15690 );
xor \U$15315 ( \15692 , \15663 , \15691 );
xor \U$15316 ( \15693 , \14118 , \14128 );
and \U$15317 ( \15694 , \15693 , \14138 );
and \U$15318 ( \15695 , \14118 , \14128 );
or \U$15319 ( \15696 , \15694 , \15695 );
not \U$15320 ( \15697 , \15696 );
xor \U$15321 ( \15698 , \13891 , \13902 );
and \U$15322 ( \15699 , \15698 , \13910 );
and \U$15323 ( \15700 , \13891 , \13902 );
nor \U$15324 ( \15701 , \15699 , \15700 );
not \U$15325 ( \15702 , \15701 );
xor \U$15326 ( \15703 , \13980 , \13992 );
and \U$15327 ( \15704 , \15703 , \14003 );
and \U$15328 ( \15705 , \13980 , \13992 );
or \U$15329 ( \15706 , \15704 , \15705 );
not \U$15330 ( \15707 , \15706 );
or \U$15331 ( \15708 , \15702 , \15707 );
or \U$15332 ( \15709 , \15706 , \15701 );
nand \U$15333 ( \15710 , \15708 , \15709 );
not \U$15334 ( \15711 , \15710 );
or \U$15335 ( \15712 , \15697 , \15711 );
not \U$15336 ( \15713 , \15701 );
nand \U$15337 ( \15714 , \15713 , \15706 );
nand \U$15338 ( \15715 , \15712 , \15714 );
xor \U$15339 ( \15716 , \15692 , \15715 );
xor \U$15340 ( \15717 , \15701 , \15706 );
xnor \U$15341 ( \15718 , \15717 , \15696 );
not \U$15342 ( \15719 , \15718 );
or \U$15343 ( \15720 , \14171 , \14139 );
buf \U$15344 ( \15721 , \14143 );
nand \U$15345 ( \15722 , \15720 , \15721 );
nand \U$15346 ( \15723 , \14171 , \14139 );
nand \U$15347 ( \15724 , \15722 , \15723 );
not \U$15348 ( \15725 , \15724 );
or \U$15349 ( \15726 , \15719 , \15725 );
or \U$15350 ( \15727 , \15724 , \15718 );
not \U$15351 ( \15728 , RIae7a948_189);
not \U$15352 ( \15729 , RIae7a7e0_186);
or \U$15353 ( \15730 , \15728 , \15729 );
nand \U$15354 ( \15731 , \15730 , RIae7a060_170);
not \U$15355 ( \15732 , \951 );
not \U$15356 ( \15733 , \13906 );
or \U$15357 ( \15734 , \15732 , \15733 );
nand \U$15358 ( \15735 , \15655 , \926 );
nand \U$15359 ( \15736 , \15734 , \15735 );
xor \U$15360 ( \15737 , \15731 , \15736 );
not \U$15361 ( \15738 , \5858 );
not \U$15362 ( \15739 , \13663 );
or \U$15363 ( \15740 , \15738 , \15739 );
nand \U$15364 ( \15741 , \15506 , \1320 );
nand \U$15365 ( \15742 , \15740 , \15741 );
xor \U$15366 ( \15743 , \15737 , \15742 );
and \U$15367 ( \15744 , RIae78b48_125, \10007 );
not \U$15368 ( \15745 , \1129 );
not \U$15369 ( \15746 , \13898 );
or \U$15370 ( \15747 , \15745 , \15746 );
and \U$15371 ( \15748 , RIae78b48_125, \10171 );
not \U$15372 ( \15749 , RIae78b48_125);
and \U$15373 ( \15750 , \15749 , \13544 );
or \U$15374 ( \15751 , \15748 , \15750 );
nand \U$15375 ( \15752 , \15751 , \867 );
nand \U$15376 ( \15753 , \15747 , \15752 );
xor \U$15377 ( \15754 , \15744 , \15753 );
not \U$15378 ( \15755 , \2272 );
not \U$15379 ( \15756 , \14001 );
or \U$15380 ( \15757 , \15755 , \15756 );
nand \U$15381 ( \15758 , \15368 , \10414 );
nand \U$15382 ( \15759 , \15757 , \15758 );
xor \U$15383 ( \15760 , \15754 , \15759 );
xor \U$15384 ( \15761 , \15743 , \15760 );
xor \U$15385 ( \15762 , \14154 , \14164 );
and \U$15386 ( \15763 , \15762 , \14170 );
and \U$15387 ( \15764 , \14154 , \14164 );
or \U$15388 ( \15765 , \15763 , \15764 );
xor \U$15389 ( \15766 , \15761 , \15765 );
nand \U$15390 ( \15767 , \15727 , \15766 );
nand \U$15391 ( \15768 , \15726 , \15767 );
xor \U$15392 ( \15769 , \15716 , \15768 );
xor \U$15393 ( \15770 , \15743 , \15760 );
and \U$15394 ( \15771 , \15770 , \15765 );
and \U$15395 ( \15772 , \15743 , \15760 );
or \U$15396 ( \15773 , \15771 , \15772 );
not \U$15397 ( \15774 , \15773 );
xor \U$15398 ( \15775 , \15731 , \15736 );
and \U$15399 ( \15776 , \15775 , \15742 );
and \U$15400 ( \15777 , \15731 , \15736 );
nor \U$15401 ( \15778 , \15776 , \15777 );
not \U$15402 ( \15779 , \15778 );
not \U$15403 ( \15780 , \1919 );
not \U$15404 ( \15781 , \3039 );
buf \U$15405 ( \15782 , \2675 );
not \U$15406 ( \15783 , \15782 );
or \U$15407 ( \15784 , \15781 , \15783 );
nand \U$15408 ( \15785 , \2676 , RIae794a8_145);
nand \U$15409 ( \15786 , \15784 , \15785 );
not \U$15410 ( \15787 , \15786 );
or \U$15411 ( \15788 , \15780 , \15787 );
nand \U$15412 ( \15789 , \14909 , \1933 );
nand \U$15413 ( \15790 , \15788 , \15789 );
not \U$15414 ( \15791 , \15790 );
or \U$15415 ( \15792 , \15779 , \15791 );
or \U$15416 ( \15793 , \15790 , \15778 );
nand \U$15417 ( \15794 , \15792 , \15793 );
not \U$15418 ( \15795 , \15134 );
xor \U$15419 ( \15796 , \15123 , \15146 );
not \U$15420 ( \15797 , \15796 );
or \U$15421 ( \15798 , \15795 , \15797 );
nand \U$15422 ( \15799 , \15146 , \15123 );
nand \U$15423 ( \15800 , \15798 , \15799 );
xor \U$15424 ( \15801 , \15794 , \15800 );
xor \U$15425 ( \15802 , \15774 , \15801 );
xor \U$15426 ( \15803 , \15744 , \15753 );
and \U$15427 ( \15804 , \15803 , \15759 );
and \U$15428 ( \15805 , \15744 , \15753 );
or \U$15429 ( \15806 , \15804 , \15805 );
xor \U$15430 ( \15807 , \15085 , \15097 );
and \U$15431 ( \15808 , \15807 , \15109 );
and \U$15432 ( \15809 , \15085 , \15097 );
or \U$15433 ( \15810 , \15808 , \15809 );
xor \U$15434 ( \15811 , \15806 , \15810 );
nand \U$15435 ( \15812 , \9868 , RIae78b48_125);
not \U$15436 ( \15813 , \867 );
and \U$15437 ( \15814 , RIae78b48_125, \10067 );
not \U$15438 ( \15815 , RIae78b48_125);
and \U$15439 ( \15816 , \15815 , \10070 );
or \U$15440 ( \15817 , \15814 , \15816 );
not \U$15441 ( \15818 , \15817 );
or \U$15442 ( \15819 , \15813 , \15818 );
nand \U$15443 ( \15820 , \15751 , \1129 );
nand \U$15444 ( \15821 , \15819 , \15820 );
xor \U$15445 ( \15822 , \15812 , \15821 );
not \U$15446 ( \15823 , \1820 );
not \U$15447 ( \15824 , RIae79688_149);
not \U$15448 ( \15825 , \9830 );
or \U$15449 ( \15826 , \15824 , \15825 );
nand \U$15450 ( \15827 , \4982 , \3147 );
nand \U$15451 ( \15828 , \15826 , \15827 );
not \U$15452 ( \15829 , \15828 );
or \U$15453 ( \15830 , \15823 , \15829 );
nand \U$15454 ( \15831 , \15144 , \9320 );
nand \U$15455 ( \15832 , \15830 , \15831 );
xnor \U$15456 ( \15833 , \15822 , \15832 );
xor \U$15457 ( \15834 , \15811 , \15833 );
buf \U$15458 ( \15835 , \15834 );
xnor \U$15459 ( \15836 , \15802 , \15835 );
xor \U$15460 ( \15837 , \15769 , \15836 );
not \U$15461 ( \15838 , \15575 );
nand \U$15462 ( \15839 , \15590 , \15838 );
not \U$15463 ( \15840 , \15582 );
and \U$15464 ( \15841 , \15839 , \15840 );
nor \U$15465 ( \15842 , \15590 , \15838 );
nor \U$15466 ( \15843 , \15841 , \15842 );
xor \U$15467 ( \15844 , \15837 , \15843 );
xor \U$15468 ( \15845 , \15260 , \15252 );
xor \U$15469 ( \15846 , \15845 , \15274 );
not \U$15470 ( \15847 , \15846 );
xor \U$15471 ( \15848 , \15766 , \15718 );
xnor \U$15472 ( \15849 , \15848 , \15724 );
not \U$15473 ( \15850 , \13811 );
nand \U$15474 ( \15851 , \15850 , \13847 );
not \U$15475 ( \15852 , \13811 );
not \U$15476 ( \15853 , \13844 );
or \U$15477 ( \15854 , \15852 , \15853 );
buf \U$15478 ( \15855 , \13804 );
nand \U$15479 ( \15856 , \15854 , \15855 );
and \U$15480 ( \15857 , \15851 , \15856 );
and \U$15481 ( \15858 , \15849 , \15857 );
not \U$15482 ( \15859 , \15849 );
nand \U$15483 ( \15860 , \15856 , \15851 );
and \U$15484 ( \15861 , \15859 , \15860 );
nor \U$15485 ( \15862 , \15858 , \15861 );
not \U$15486 ( \15863 , \15862 );
or \U$15487 ( \15864 , \15847 , \15863 );
not \U$15488 ( \15865 , \15851 );
not \U$15489 ( \15866 , \15856 );
or \U$15490 ( \15867 , \15865 , \15866 );
not \U$15491 ( \15868 , \15849 );
nand \U$15492 ( \15869 , \15867 , \15868 );
nand \U$15493 ( \15870 , \15864 , \15869 );
xor \U$15494 ( \15871 , \15844 , \15870 );
xor \U$15495 ( \15872 , \15158 , \15149 );
not \U$15496 ( \15873 , \15872 );
xor \U$15497 ( \15874 , \15062 , \15873 );
not \U$15498 ( \15875 , \15874 );
nand \U$15499 ( \15876 , \14187 , \14198 );
nand \U$15500 ( \15877 , \14190 , \15876 );
not \U$15501 ( \15878 , \15877 );
not \U$15502 ( \15879 , \15846 );
and \U$15503 ( \15880 , \15862 , \15879 );
not \U$15504 ( \15881 , \15862 );
and \U$15505 ( \15882 , \15881 , \15846 );
nor \U$15506 ( \15883 , \15880 , \15882 );
not \U$15507 ( \15884 , \15883 );
or \U$15508 ( \15885 , \15878 , \15884 );
or \U$15509 ( \15886 , \15877 , \15883 );
nand \U$15510 ( \15887 , \15885 , \15886 );
not \U$15511 ( \15888 , \15887 );
or \U$15512 ( \15889 , \15875 , \15888 );
not \U$15513 ( \15890 , \15883 );
nand \U$15514 ( \15891 , \15890 , \15877 );
nand \U$15515 ( \15892 , \15889 , \15891 );
not \U$15516 ( \15893 , \15892 );
xor \U$15517 ( \15894 , \15871 , \15893 );
not \U$15518 ( \15895 , \15591 );
not \U$15519 ( \15896 , \15895 );
not \U$15520 ( \15897 , \15604 );
or \U$15521 ( \15898 , \15896 , \15897 );
not \U$15522 ( \15899 , \15602 );
not \U$15523 ( \15900 , \15598 );
or \U$15524 ( \15901 , \15899 , \15900 );
nand \U$15525 ( \15902 , \15901 , \15597 );
nand \U$15526 ( \15903 , \15898 , \15902 );
xnor \U$15527 ( \15904 , \15894 , \15903 );
xnor \U$15528 ( \15905 , \15621 , \15904 );
xnor \U$15529 ( \15906 , \15874 , \15887 );
not \U$15530 ( \15907 , \15561 );
and \U$15531 ( \15908 , \15614 , \15907 );
not \U$15532 ( \15909 , \15614 );
and \U$15533 ( \15910 , \15909 , \15561 );
nor \U$15534 ( \15911 , \15908 , \15910 );
xor \U$15535 ( \15912 , \15906 , \15911 );
and \U$15536 ( \15913 , \13783 , \13622 );
and \U$15537 ( \15914 , \13633 , \13782 );
nor \U$15538 ( \15915 , \15913 , \15914 );
and \U$15539 ( \15916 , \15912 , \15915 );
and \U$15540 ( \15917 , \15906 , \15911 );
or \U$15541 ( \15918 , \15916 , \15917 );
nand \U$15542 ( \15919 , \15905 , \15918 );
not \U$15543 ( \15920 , \13784 );
not \U$15544 ( \15921 , \14214 );
or \U$15545 ( \15922 , \15920 , \15921 );
not \U$15546 ( \15923 , \14212 );
nand \U$15547 ( \15924 , \15923 , \14204 );
nand \U$15548 ( \15925 , \15922 , \15924 );
not \U$15549 ( \15926 , \15925 );
xor \U$15550 ( \15927 , \15906 , \15911 );
xor \U$15551 ( \15928 , \15927 , \15915 );
nand \U$15552 ( \15929 , \15926 , \15928 );
nand \U$15553 ( \15930 , \14884 , \15919 , \15929 );
not \U$15554 ( \15931 , \15930 );
not \U$15555 ( \15932 , \1820 );
not \U$15556 ( \15933 , RIae79688_149);
not \U$15557 ( \15934 , \12603 );
or \U$15558 ( \15935 , \15933 , \15934 );
or \U$15559 ( \15936 , \14156 , RIae79688_149);
nand \U$15560 ( \15937 , \15935 , \15936 );
not \U$15561 ( \15938 , \15937 );
or \U$15562 ( \15939 , \15932 , \15938 );
not \U$15563 ( \15940 , \9405 );
not \U$15564 ( \15941 , \9407 );
and \U$15565 ( \15942 , \15940 , \15941 );
and \U$15566 ( \15943 , \9405 , \9407 );
nor \U$15567 ( \15944 , \15942 , \15943 );
and \U$15568 ( \15945 , RIae79688_149, \15944 );
not \U$15569 ( \15946 , RIae79688_149);
not \U$15570 ( \15947 , \15944 );
and \U$15571 ( \15948 , \15946 , \15947 );
or \U$15572 ( \15949 , \15945 , \15948 );
nand \U$15573 ( \15950 , \15949 , \10401 );
nand \U$15574 ( \15951 , \15939 , \15950 );
not \U$15575 ( \15952 , \2011 );
xor \U$15576 ( \15953 , RIae79610_148, \12482 );
not \U$15577 ( \15954 , \15953 );
or \U$15578 ( \15955 , \15952 , \15954 );
not \U$15579 ( \15956 , RIae79610_148);
not \U$15580 ( \15957 , \10464 );
or \U$15581 ( \15958 , \15956 , \15957 );
or \U$15582 ( \15959 , \10461 , RIae79610_148);
nand \U$15583 ( \15960 , \15958 , \15959 );
nand \U$15584 ( \15961 , \15960 , \2063 );
nand \U$15585 ( \15962 , \15955 , \15961 );
and \U$15586 ( \15963 , \15951 , \15962 );
not \U$15587 ( \15964 , \15951 );
not \U$15588 ( \15965 , \15962 );
and \U$15589 ( \15966 , \15964 , \15965 );
nor \U$15590 ( \15967 , \15963 , \15966 );
not \U$15591 ( \15968 , \15967 );
not \U$15592 ( \15969 , \11037 );
and \U$15593 ( \15970 , RIae79778_151, \3207 );
not \U$15594 ( \15971 , RIae79778_151);
and \U$15595 ( \15972 , \15971 , \10809 );
nor \U$15596 ( \15973 , \15970 , \15972 );
not \U$15597 ( \15974 , \15973 );
or \U$15598 ( \15975 , \15969 , \15974 );
not \U$15599 ( \15976 , RIae79778_151);
not \U$15600 ( \15977 , \6242 );
or \U$15601 ( \15978 , \15976 , \15977 );
or \U$15602 ( \15979 , \6242 , RIae79778_151);
nand \U$15603 ( \15980 , \15978 , \15979 );
nand \U$15604 ( \15981 , \15980 , \9576 );
nand \U$15605 ( \15982 , \15975 , \15981 );
not \U$15606 ( \15983 , \15982 );
and \U$15607 ( \15984 , \15968 , \15983 );
and \U$15608 ( \15985 , \15982 , \15967 );
nor \U$15609 ( \15986 , \15984 , \15985 );
not \U$15610 ( \15987 , \15986 );
not \U$15611 ( \15988 , \15987 );
buf \U$15612 ( \15989 , \6200 );
not \U$15613 ( \15990 , \15989 );
xnor \U$15614 ( \15991 , RIae79ef8_167, \3416 );
not \U$15615 ( \15992 , \15991 );
or \U$15616 ( \15993 , \15990 , \15992 );
xnor \U$15617 ( \15994 , RIae79ef8_167, \1788 );
nand \U$15618 ( \15995 , \15994 , \10573 );
nand \U$15619 ( \15996 , \15993 , \15995 );
not \U$15620 ( \15997 , \15996 );
nand \U$15621 ( \15998 , \1066 , \922 );
not \U$15622 ( \15999 , \15998 );
not \U$15623 ( \16000 , \12857 );
or \U$15624 ( \16001 , \15999 , \16000 );
nand \U$15625 ( \16002 , \16001 , \1706 );
not \U$15626 ( \16003 , \16002 );
not \U$15627 ( \16004 , \926 );
buf \U$15628 ( \16005 , \12749 );
buf \U$15629 ( \16006 , \16005 );
and \U$15630 ( \16007 , \1286 , \16006 );
not \U$15631 ( \16008 , \1286 );
not \U$15632 ( \16009 , \16006 );
and \U$15633 ( \16010 , \16008 , \16009 );
nor \U$15634 ( \16011 , \16007 , \16010 );
not \U$15635 ( \16012 , \16011 );
or \U$15636 ( \16013 , \16004 , \16012 );
not \U$15637 ( \16014 , \1286 );
not \U$15638 ( \16015 , \12857 );
or \U$15639 ( \16016 , \16014 , \16015 );
or \U$15640 ( \16017 , \12857 , \1286 );
nand \U$15641 ( \16018 , \16016 , \16017 );
nand \U$15642 ( \16019 , \16018 , \949 );
nand \U$15643 ( \16020 , \16013 , \16019 );
nand \U$15644 ( \16021 , \16003 , \16020 );
not \U$15645 ( \16022 , \16021 );
not \U$15646 ( \16023 , \838 );
not \U$15647 ( \16024 , \10042 );
not \U$15648 ( \16025 , \3105 );
or \U$15649 ( \16026 , \16024 , \16025 );
or \U$15650 ( \16027 , \10042 , \3105 );
nand \U$15651 ( \16028 , \16026 , \16027 );
not \U$15652 ( \16029 , \16028 );
or \U$15653 ( \16030 , \16023 , \16029 );
not \U$15654 ( \16031 , RIae78f80_134);
and \U$15655 ( \16032 , \10186 , \10187 );
not \U$15656 ( \16033 , \10186 );
and \U$15657 ( \16034 , \16033 , \10190 );
nor \U$15658 ( \16035 , \16032 , \16034 );
not \U$15659 ( \16036 , \16035 );
not \U$15660 ( \16037 , \16036 );
or \U$15661 ( \16038 , \16031 , \16037 );
or \U$15662 ( \16039 , \11581 , RIae78f80_134);
nand \U$15663 ( \16040 , \16038 , \16039 );
nand \U$15664 ( \16041 , \16040 , \796 );
nand \U$15665 ( \16042 , \16030 , \16041 );
not \U$15666 ( \16043 , \16042 );
or \U$15667 ( \16044 , \16022 , \16043 );
or \U$15668 ( \16045 , \16042 , \16021 );
nand \U$15669 ( \16046 , \16044 , \16045 );
buf \U$15670 ( \16047 , \16046 );
not \U$15671 ( \16048 , \16047 );
not \U$15672 ( \16049 , \1062 );
not \U$15673 ( \16050 , \1039 );
not \U$15674 ( \16051 , \10031 );
or \U$15675 ( \16052 , \16050 , \16051 );
or \U$15676 ( \16053 , \10032 , \1039 );
nand \U$15677 ( \16054 , \16052 , \16053 );
not \U$15678 ( \16055 , \16054 );
or \U$15679 ( \16056 , \16049 , \16055 );
not \U$15680 ( \16057 , \1039 );
not \U$15681 ( \16058 , \10141 );
or \U$15682 ( \16059 , \16057 , \16058 );
nand \U$15683 ( \16060 , \10149 , RIae79070_136);
nand \U$15684 ( \16061 , \16059 , \16060 );
nand \U$15685 ( \16062 , \16061 , \1049 );
nand \U$15686 ( \16063 , \16056 , \16062 );
not \U$15687 ( \16064 , \16063 );
not \U$15688 ( \16065 , \16064 );
and \U$15689 ( \16066 , \16048 , \16065 );
and \U$15690 ( \16067 , \16047 , \16064 );
nor \U$15691 ( \16068 , \16066 , \16067 );
not \U$15692 ( \16069 , \16068 );
not \U$15693 ( \16070 , \16069 );
or \U$15694 ( \16071 , \15997 , \16070 );
not \U$15695 ( \16072 , \16068 );
not \U$15696 ( \16073 , \15996 );
not \U$15697 ( \16074 , \16073 );
or \U$15698 ( \16075 , \16072 , \16074 );
not \U$15699 ( \16076 , \9776 );
and \U$15700 ( \16077 , RIae7a150_172, \1404 );
not \U$15701 ( \16078 , RIae7a150_172);
and \U$15702 ( \16079 , \16078 , \9624 );
nor \U$15703 ( \16080 , \16077 , \16079 );
not \U$15704 ( \16081 , \16080 );
or \U$15705 ( \16082 , \16076 , \16081 );
not \U$15706 ( \16083 , RIae7a150_172);
not \U$15707 ( \16084 , \5134 );
or \U$15708 ( \16085 , \16083 , \16084 );
not \U$15709 ( \16086 , \14071 );
or \U$15710 ( \16087 , \16086 , RIae7a150_172);
nand \U$15711 ( \16088 , \16085 , \16087 );
nand \U$15712 ( \16089 , \16088 , \13158 );
nand \U$15713 ( \16090 , \16082 , \16089 );
nand \U$15714 ( \16091 , \16075 , \16090 );
nand \U$15715 ( \16092 , \16071 , \16091 );
not \U$15716 ( \16093 , \16092 );
not \U$15717 ( \16094 , \16093 );
or \U$15718 ( \16095 , \15988 , \16094 );
nand \U$15719 ( \16096 , \15986 , \16092 );
nand \U$15720 ( \16097 , \16095 , \16096 );
not \U$15721 ( \16098 , \16097 );
not \U$15722 ( \16099 , \9473 );
not \U$15723 ( \16100 , \854 );
not \U$15724 ( \16101 , RIae7a6f0_184);
not \U$15725 ( \16102 , \16101 );
or \U$15726 ( \16103 , \16100 , \16102 );
not \U$15727 ( \16104 , RIae7a6f0_184);
or \U$15728 ( \16105 , \854 , \16104 );
nand \U$15729 ( \16106 , \16103 , \16105 );
not \U$15730 ( \16107 , \16106 );
or \U$15731 ( \16108 , \16099 , \16107 );
and \U$15732 ( \16109 , RIae7a6f0_184, \9770 );
not \U$15733 ( \16110 , RIae7a6f0_184);
and \U$15734 ( \16111 , \16110 , \3235 );
nor \U$15735 ( \16112 , \16109 , \16111 );
nand \U$15736 ( \16113 , \16112 , \9705 );
nand \U$15737 ( \16114 , \16108 , \16113 );
not \U$15738 ( \16115 , \10709 );
xor \U$15739 ( \16116 , RIae79fe8_169, \1808 );
not \U$15740 ( \16117 , \16116 );
or \U$15741 ( \16118 , \16115 , \16117 );
and \U$15742 ( \16119 , RIae79fe8_169, \1758 );
not \U$15743 ( \16120 , RIae79fe8_169);
and \U$15744 ( \16121 , \16120 , \4582 );
or \U$15745 ( \16122 , \16119 , \16121 );
nand \U$15746 ( \16123 , \16122 , \9518 );
nand \U$15747 ( \16124 , \16118 , \16123 );
not \U$15748 ( \16125 , \16124 );
not \U$15749 ( \16126 , \9792 );
xor \U$15750 ( \16127 , RIae7a2b8_175, \3093 );
not \U$15751 ( \16128 , \16127 );
or \U$15752 ( \16129 , \16126 , \16128 );
not \U$15753 ( \16130 , RIae7a2b8_175);
not \U$15754 ( \16131 , \2835 );
or \U$15755 ( \16132 , \16130 , \16131 );
nand \U$15756 ( \16133 , \3747 , \9804 );
nand \U$15757 ( \16134 , \16132 , \16133 );
buf \U$15758 ( \16135 , \9813 );
nand \U$15759 ( \16136 , \16134 , \16135 );
nand \U$15760 ( \16137 , \16129 , \16136 );
not \U$15761 ( \16138 , \16137 );
nor \U$15762 ( \16139 , \16125 , \16138 );
or \U$15763 ( \16140 , \16114 , \16139 );
not \U$15764 ( \16141 , \16124 );
nand \U$15765 ( \16142 , \16141 , \16138 );
nand \U$15766 ( \16143 , \16140 , \16142 );
not \U$15767 ( \16144 , \16143 );
not \U$15768 ( \16145 , \16144 );
and \U$15769 ( \16146 , \16098 , \16145 );
and \U$15770 ( \16147 , \16097 , \16144 );
nor \U$15771 ( \16148 , \16146 , \16147 );
not \U$15772 ( \16149 , \16148 );
not \U$15773 ( \16150 , \16149 );
not \U$15774 ( \16151 , \9403 );
xor \U$15775 ( \16152 , RIae79250_140, \9868 );
not \U$15776 ( \16153 , \16152 );
or \U$15777 ( \16154 , \16151 , \16153 );
not \U$15778 ( \16155 , \8789 );
not \U$15779 ( \16156 , \13544 );
or \U$15780 ( \16157 , \16155 , \16156 );
or \U$15781 ( \16158 , \9900 , \1503 );
nand \U$15782 ( \16159 , \16157 , \16158 );
nand \U$15783 ( \16160 , \16159 , \1501 );
nand \U$15784 ( \16161 , \16154 , \16160 );
and \U$15785 ( \16162 , \12857 , \867 );
not \U$15786 ( \16163 , \926 );
not \U$15787 ( \16164 , \10844 );
not \U$15788 ( \16165 , \16164 );
buf \U$15789 ( \16166 , \16165 );
and \U$15790 ( \16167 , \16166 , \1286 );
not \U$15791 ( \16168 , \16166 );
and \U$15792 ( \16169 , \16168 , RIae78bc0_126);
nor \U$15793 ( \16170 , \16167 , \16169 );
not \U$15794 ( \16171 , \16170 );
or \U$15795 ( \16172 , \16163 , \16171 );
nand \U$15796 ( \16173 , \16011 , \949 );
nand \U$15797 ( \16174 , \16172 , \16173 );
xor \U$15798 ( \16175 , \16162 , \16174 );
not \U$15799 ( \16176 , \1072 );
not \U$15800 ( \16177 , \1066 );
not \U$15801 ( \16178 , \10272 );
or \U$15802 ( \16179 , \16177 , \16178 );
or \U$15803 ( \16180 , \11318 , \921 );
nand \U$15804 ( \16181 , \16179 , \16180 );
not \U$15805 ( \16182 , \16181 );
or \U$15806 ( \16183 , \16176 , \16182 );
and \U$15807 ( \16184 , RIae78e90_132, \10259 );
not \U$15808 ( \16185 , RIae78e90_132);
and \U$15809 ( \16186 , \16185 , \11309 );
or \U$15810 ( \16187 , \16184 , \16186 );
nand \U$15811 ( \16188 , \16187 , \1086 );
nand \U$15812 ( \16189 , \16183 , \16188 );
xor \U$15813 ( \16190 , \16175 , \16189 );
xor \U$15814 ( \16191 , \16161 , \16190 );
not \U$15815 ( \16192 , \1008 );
buf \U$15816 ( \16193 , \9988 );
not \U$15817 ( \16194 , \16193 );
and \U$15818 ( \16195 , \16194 , RIae79160_138);
not \U$15819 ( \16196 , \16194 );
and \U$15820 ( \16197 , \16196 , \997 );
nor \U$15821 ( \16198 , \16195 , \16197 );
not \U$15822 ( \16199 , \16198 );
or \U$15823 ( \16200 , \16192 , \16199 );
and \U$15824 ( \16201 , RIae79160_138, \11260 );
not \U$15825 ( \16202 , RIae79160_138);
and \U$15826 ( \16203 , \16202 , \10007 );
or \U$15827 ( \16204 , \16201 , \16203 );
nand \U$15828 ( \16205 , \16204 , \1012 );
nand \U$15829 ( \16206 , \16200 , \16205 );
and \U$15830 ( \16207 , \16191 , \16206 );
and \U$15831 ( \16208 , \16161 , \16190 );
nor \U$15832 ( \16209 , \16207 , \16208 );
not \U$15833 ( \16210 , \16209 );
not \U$15834 ( \16211 , \10675 );
and \U$15835 ( \16212 , RIae7a498_179, \2025 );
not \U$15836 ( \16213 , RIae7a498_179);
and \U$15837 ( \16214 , \16213 , \2030 );
nor \U$15838 ( \16215 , \16212 , \16214 );
not \U$15839 ( \16216 , \16215 );
or \U$15840 ( \16217 , \16211 , \16216 );
not \U$15841 ( \16218 , RIae7a498_179);
not \U$15842 ( \16219 , \3145 );
or \U$15843 ( \16220 , \16218 , \16219 );
or \U$15844 ( \16221 , \9696 , RIae7a498_179);
nand \U$15845 ( \16222 , \16220 , \16221 );
nand \U$15846 ( \16223 , \16222 , \10696 );
nand \U$15847 ( \16224 , \16217 , \16223 );
not \U$15848 ( \16225 , \16224 );
or \U$15849 ( \16226 , \16210 , \16225 );
or \U$15850 ( \16227 , \16224 , \16209 );
nand \U$15851 ( \16228 , \16226 , \16227 );
not \U$15852 ( \16229 , \5048 );
and \U$15853 ( \16230 , \2676 , \4968 );
not \U$15854 ( \16231 , \2676 );
and \U$15855 ( \16232 , \16231 , RIae79d90_164);
nor \U$15856 ( \16233 , \16230 , \16232 );
not \U$15857 ( \16234 , \16233 );
or \U$15858 ( \16235 , \16229 , \16234 );
and \U$15859 ( \16236 , RIae79d90_164, \2089 );
not \U$15860 ( \16237 , RIae79d90_164);
and \U$15861 ( \16238 , \16237 , \2785 );
nor \U$15862 ( \16239 , \16236 , \16238 );
nand \U$15863 ( \16240 , \16239 , \6091 );
nand \U$15864 ( \16241 , \16235 , \16240 );
xnor \U$15865 ( \16242 , \16228 , \16241 );
not \U$15866 ( \16243 , \16242 );
not \U$15867 ( \16244 , \3440 );
not \U$15868 ( \16245 , RIae79520_146);
not \U$15869 ( \16246 , \12707 );
or \U$15870 ( \16247 , \16245 , \16246 );
nand \U$15871 ( \16248 , \15519 , \4653 );
nand \U$15872 ( \16249 , \16247 , \16248 );
not \U$15873 ( \16250 , \16249 );
or \U$15874 ( \16251 , \16244 , \16250 );
and \U$15875 ( \16252 , RIae79520_146, \9367 );
not \U$15876 ( \16253 , RIae79520_146);
not \U$15877 ( \16254 , \9363 );
and \U$15878 ( \16255 , \16253 , \16254 );
nor \U$15879 ( \16256 , \16252 , \16255 );
nand \U$15880 ( \16257 , \16256 , \12680 );
nand \U$15881 ( \16258 , \16251 , \16257 );
not \U$15882 ( \16259 , \1919 );
not \U$15883 ( \16260 , \9298 );
and \U$15884 ( \16261 , RIae794a8_145, \16260 );
not \U$15885 ( \16262 , RIae794a8_145);
and \U$15886 ( \16263 , \16262 , \6230 );
or \U$15887 ( \16264 , \16261 , \16263 );
not \U$15888 ( \16265 , \16264 );
or \U$15889 ( \16266 , \16259 , \16265 );
not \U$15890 ( \16267 , \9306 );
not \U$15891 ( \16268 , \9308 );
and \U$15892 ( \16269 , \16267 , \16268 );
and \U$15893 ( \16270 , \9306 , \9308 );
nor \U$15894 ( \16271 , \16269 , \16270 );
and \U$15895 ( \16272 , RIae794a8_145, \16271 );
not \U$15896 ( \16273 , RIae794a8_145);
not \U$15897 ( \16274 , \16271 );
and \U$15898 ( \16275 , \16273 , \16274 );
or \U$15899 ( \16276 , \16272 , \16275 );
nand \U$15900 ( \16277 , \16276 , \2457 );
nand \U$15901 ( \16278 , \16266 , \16277 );
not \U$15902 ( \16279 , \2251 );
not \U$15903 ( \16280 , \2268 );
not \U$15904 ( \16281 , \9441 );
or \U$15905 ( \16282 , \16280 , \16281 );
or \U$15906 ( \16283 , \9441 , \2268 );
nand \U$15907 ( \16284 , \16282 , \16283 );
not \U$15908 ( \16285 , \16284 );
or \U$15909 ( \16286 , \16279 , \16285 );
and \U$15910 ( \16287 , RIae79ac0_158, \9455 );
not \U$15911 ( \16288 , RIae79ac0_158);
and \U$15912 ( \16289 , \16288 , \13301 );
nor \U$15913 ( \16290 , \16287 , \16289 );
nand \U$15914 ( \16291 , \16290 , \2272 );
nand \U$15915 ( \16292 , \16286 , \16291 );
and \U$15916 ( \16293 , \16278 , \16292 );
not \U$15917 ( \16294 , \16278 );
not \U$15918 ( \16295 , \16292 );
and \U$15919 ( \16296 , \16294 , \16295 );
nor \U$15920 ( \16297 , \16293 , \16296 );
xor \U$15921 ( \16298 , \16258 , \16297 );
not \U$15922 ( \16299 , \16298 );
not \U$15923 ( \16300 , \16299 );
not \U$15924 ( \16301 , \2007 );
not \U$15925 ( \16302 , RIae797f0_152);
not \U$15926 ( \16303 , \10829 );
or \U$15927 ( \16304 , \16302 , \16303 );
or \U$15928 ( \16305 , \10829 , RIae797f0_152);
nand \U$15929 ( \16306 , \16304 , \16305 );
not \U$15930 ( \16307 , \16306 );
or \U$15931 ( \16308 , \16301 , \16307 );
not \U$15932 ( \16309 , \2521 );
not \U$15933 ( \16310 , \5107 );
not \U$15934 ( \16311 , \16310 );
not \U$15935 ( \16312 , \16311 );
or \U$15936 ( \16313 , \16309 , \16312 );
nand \U$15937 ( \16314 , \13248 , RIae797f0_152);
nand \U$15938 ( \16315 , \16313 , \16314 );
nand \U$15939 ( \16316 , \16315 , \1988 );
nand \U$15940 ( \16317 , \16308 , \16316 );
not \U$15941 ( \16318 , \16063 );
not \U$15942 ( \16319 , \16046 );
or \U$15943 ( \16320 , \16318 , \16319 );
not \U$15944 ( \16321 , \16021 );
nand \U$15945 ( \16322 , \16321 , \16042 );
nand \U$15946 ( \16323 , \16320 , \16322 );
not \U$15947 ( \16324 , \16323 );
not \U$15948 ( \16325 , \2339 );
xor \U$15949 ( \16326 , RIae798e0_154, \9289 );
not \U$15950 ( \16327 , \16326 );
or \U$15951 ( \16328 , \16325 , \16327 );
and \U$15952 ( \16329 , RIae798e0_154, \5722 );
not \U$15953 ( \16330 , RIae798e0_154);
and \U$15954 ( \16331 , \16330 , \10793 );
nor \U$15955 ( \16332 , \16329 , \16331 );
nand \U$15956 ( \16333 , \16332 , \2321 );
nand \U$15957 ( \16334 , \16328 , \16333 );
not \U$15958 ( \16335 , \16334 );
not \U$15959 ( \16336 , \16335 );
or \U$15960 ( \16337 , \16324 , \16336 );
or \U$15961 ( \16338 , \16335 , \16323 );
nand \U$15962 ( \16339 , \16337 , \16338 );
xnor \U$15963 ( \16340 , \16317 , \16339 );
not \U$15964 ( \16341 , \16340 );
not \U$15965 ( \16342 , \16341 );
or \U$15966 ( \16343 , \16300 , \16342 );
nand \U$15967 ( \16344 , \16340 , \16298 );
nand \U$15968 ( \16345 , \16343 , \16344 );
not \U$15969 ( \16346 , \16345 );
or \U$15970 ( \16347 , \16243 , \16346 );
or \U$15971 ( \16348 , \16345 , \16242 );
nand \U$15972 ( \16349 , \16347 , \16348 );
not \U$15973 ( \16350 , \16349 );
not \U$15974 ( \16351 , \16350 );
or \U$15975 ( \16352 , \16150 , \16351 );
nand \U$15976 ( \16353 , \16349 , \16148 );
nand \U$15977 ( \16354 , \16352 , \16353 );
not \U$15978 ( \16355 , \1878 );
xor \U$15979 ( \16356 , RIae7a510_180, \16355 );
not \U$15980 ( \16357 , \16356 );
not \U$15981 ( \16358 , \12232 );
not \U$15982 ( \16359 , \16358 );
or \U$15983 ( \16360 , \16357 , \16359 );
not \U$15984 ( \16361 , \10633 );
not \U$15985 ( \16362 , \1897 );
or \U$15986 ( \16363 , \16361 , \16362 );
or \U$15987 ( \16364 , \1898 , \14931 );
nand \U$15988 ( \16365 , \16363 , \16364 );
nand \U$15989 ( \16366 , \16365 , \10638 );
nand \U$15990 ( \16367 , \16360 , \16366 );
not \U$15991 ( \16368 , \16367 );
not \U$15992 ( \16369 , RIae79ca0_162);
not \U$15993 ( \16370 , \2357 );
or \U$15994 ( \16371 , \16369 , \16370 );
or \U$15995 ( \16372 , \2357 , RIae79ca0_162);
nand \U$15996 ( \16373 , \16371 , \16372 );
and \U$15997 ( \16374 , \4853 , \16373 );
xnor \U$15998 ( \16375 , \1969 , RIae79ca0_162);
and \U$15999 ( \16376 , \16375 , \4154 );
nor \U$16000 ( \16377 , \16374 , \16376 );
not \U$16001 ( \16378 , \16377 );
or \U$16002 ( \16379 , \16368 , \16378 );
or \U$16003 ( \16380 , \16377 , \16367 );
nand \U$16004 ( \16381 , \16379 , \16380 );
not \U$16005 ( \16382 , \16381 );
buf \U$16006 ( \16383 , \14667 );
not \U$16007 ( \16384 , \16383 );
not \U$16008 ( \16385 , \1994 );
not \U$16009 ( \16386 , RIae7aa38_191);
and \U$16010 ( \16387 , \16385 , \16386 );
and \U$16011 ( \16388 , \781 , RIae7aa38_191);
nor \U$16012 ( \16389 , \16387 , \16388 );
not \U$16013 ( \16390 , \16389 );
or \U$16014 ( \16391 , \16384 , \16390 );
not \U$16015 ( \16392 , RIae7aa38_191);
not \U$16016 ( \16393 , \834 );
or \U$16017 ( \16394 , \16392 , \16393 );
not \U$16018 ( \16395 , \9711 );
or \U$16019 ( \16396 , \16395 , RIae7aa38_191);
nand \U$16020 ( \16397 , \16394 , \16396 );
nand \U$16021 ( \16398 , \16397 , RIae7aab0_192);
nand \U$16022 ( \16399 , \16391 , \16398 );
not \U$16023 ( \16400 , \16399 );
and \U$16024 ( \16401 , \16382 , \16400 );
and \U$16025 ( \16402 , \16399 , \16381 );
nor \U$16026 ( \16403 , \16401 , \16402 );
not \U$16027 ( \16404 , \9777 );
not \U$16028 ( \16405 , RIae7a150_172);
not \U$16029 ( \16406 , \1186 );
or \U$16030 ( \16407 , \16405 , \16406 );
or \U$16031 ( \16408 , \1186 , RIae7a150_172);
nand \U$16032 ( \16409 , \16407 , \16408 );
not \U$16033 ( \16410 , \16409 );
or \U$16034 ( \16411 , \16404 , \16410 );
nand \U$16035 ( \16412 , \16080 , \13158 );
nand \U$16036 ( \16413 , \16411 , \16412 );
not \U$16037 ( \16414 , \16413 );
not \U$16038 ( \16415 , \10573 );
not \U$16039 ( \16416 , RIae79ef8_167);
not \U$16040 ( \16417 , \10883 );
or \U$16041 ( \16418 , \16416 , \16417 );
or \U$16042 ( \16419 , \3528 , RIae79ef8_167);
nand \U$16043 ( \16420 , \16418 , \16419 );
not \U$16044 ( \16421 , \16420 );
or \U$16045 ( \16422 , \16415 , \16421 );
nand \U$16046 ( \16423 , \15994 , \11409 );
nand \U$16047 ( \16424 , \16422 , \16423 );
not \U$16048 ( \16425 , \9517 );
and \U$16049 ( \16426 , RIae79fe8_169, \6171 );
not \U$16050 ( \16427 , RIae79fe8_169);
and \U$16051 ( \16428 , \16427 , \4024 );
nor \U$16052 ( \16429 , \16426 , \16428 );
not \U$16053 ( \16430 , \16429 );
or \U$16054 ( \16431 , \16425 , \16430 );
nand \U$16055 ( \16432 , \16122 , \10709 );
nand \U$16056 ( \16433 , \16431 , \16432 );
not \U$16057 ( \16434 , \16433 );
xor \U$16058 ( \16435 , \16424 , \16434 );
not \U$16059 ( \16436 , \16435 );
or \U$16060 ( \16437 , \16414 , \16436 );
or \U$16061 ( \16438 , \16413 , \16435 );
nand \U$16062 ( \16439 , \16437 , \16438 );
xor \U$16063 ( \16440 , \16403 , \16439 );
not \U$16064 ( \16441 , \10275 );
and \U$16065 ( \16442 , RIae7a8d0_188, \12262 );
not \U$16066 ( \16443 , RIae7a8d0_188);
and \U$16067 ( \16444 , \16443 , \3999 );
nor \U$16068 ( \16445 , \16442 , \16444 );
not \U$16069 ( \16446 , \16445 );
or \U$16070 ( \16447 , \16441 , \16446 );
not \U$16071 ( \16448 , RIae7a8d0_188);
not \U$16072 ( \16449 , \1288 );
or \U$16073 ( \16450 , \16448 , \16449 );
or \U$16074 ( \16451 , \1158 , RIae7a8d0_188);
nand \U$16075 ( \16452 , \16450 , \16451 );
nand \U$16076 ( \16453 , \16452 , \11205 );
nand \U$16077 ( \16454 , \16447 , \16453 );
not \U$16078 ( \16455 , \13121 );
xor \U$16079 ( \16456 , RIae7a240_174, \10567 );
not \U$16080 ( \16457 , \16456 );
or \U$16081 ( \16458 , \16455 , \16457 );
not \U$16082 ( \16459 , \2153 );
not \U$16083 ( \16460 , RIae7a240_174);
and \U$16084 ( \16461 , \16459 , \16460 );
and \U$16085 ( \16462 , \2954 , RIae7a240_174);
nor \U$16086 ( \16463 , \16461 , \16462 );
not \U$16087 ( \16464 , \16463 );
nand \U$16088 ( \16465 , \16464 , \13720 );
nand \U$16089 ( \16466 , \16458 , \16465 );
xor \U$16090 ( \16467 , \16454 , \16466 );
not \U$16091 ( \16468 , \9621 );
not \U$16092 ( \16469 , RIae7a3a8_177);
and \U$16093 ( \16470 , \3051 , \16469 );
not \U$16094 ( \16471 , \3051 );
and \U$16095 ( \16472 , \16471 , RIae7a3a8_177);
nor \U$16096 ( \16473 , \16470 , \16472 );
not \U$16097 ( \16474 , \16473 );
or \U$16098 ( \16475 , \16468 , \16474 );
not \U$16099 ( \16476 , RIae7a3a8_177);
not \U$16100 ( \16477 , \2230 );
or \U$16101 ( \16478 , \16476 , \16477 );
or \U$16102 ( \16479 , \2230 , RIae7a3a8_177);
nand \U$16103 ( \16480 , \16478 , \16479 );
nand \U$16104 ( \16481 , \16480 , \11014 );
nand \U$16105 ( \16482 , \16475 , \16481 );
xor \U$16106 ( \16483 , \16467 , \16482 );
xor \U$16107 ( \16484 , \16440 , \16483 );
and \U$16108 ( \16485 , \16354 , \16484 );
not \U$16109 ( \16486 , \16354 );
not \U$16110 ( \16487 , \16484 );
and \U$16111 ( \16488 , \16486 , \16487 );
nor \U$16112 ( \16489 , \16485 , \16488 );
xor \U$16113 ( \16490 , \16137 , \16124 );
xor \U$16114 ( \16491 , \16490 , \16114 );
not \U$16115 ( \16492 , \16073 );
xor \U$16116 ( \16493 , \16068 , \16492 );
xnor \U$16117 ( \16494 , \16493 , \16090 );
xor \U$16118 ( \16495 , \16491 , \16494 );
not \U$16119 ( \16496 , \11114 );
not \U$16120 ( \16497 , \2309 );
or \U$16121 ( \16498 , \16496 , \16497 );
or \U$16122 ( \16499 , \2309 , \11114 );
nand \U$16123 ( \16500 , \16498 , \16499 );
not \U$16124 ( \16501 , \16500 );
not \U$16125 ( \16502 , \9688 );
or \U$16126 ( \16503 , \16501 , \16502 );
not \U$16127 ( \16504 , \13121 );
or \U$16128 ( \16505 , \16463 , \16504 );
nand \U$16129 ( \16506 , \16503 , \16505 );
not \U$16130 ( \16507 , \10542 );
and \U$16131 ( \16508 , RIae7a060_170, \10645 );
not \U$16132 ( \16509 , RIae7a060_170);
not \U$16133 ( \16510 , \11694 );
and \U$16134 ( \16511 , \16509 , \16510 );
nor \U$16135 ( \16512 , \16508 , \16511 );
not \U$16136 ( \16513 , \16512 );
or \U$16137 ( \16514 , \16507 , \16513 );
not \U$16138 ( \16515 , \9749 );
not \U$16139 ( \16516 , \11537 );
or \U$16140 ( \16517 , \16515 , \16516 );
or \U$16141 ( \16518 , \3538 , \11102 );
nand \U$16142 ( \16519 , \16517 , \16518 );
nand \U$16143 ( \16520 , \16519 , \9728 );
nand \U$16144 ( \16521 , \16514 , \16520 );
xor \U$16145 ( \16522 , \16506 , \16521 );
not \U$16146 ( \16523 , RIae7aab0_192);
not \U$16147 ( \16524 , \16389 );
or \U$16148 ( \16525 , \16523 , \16524 );
not \U$16149 ( \16526 , \14671 );
not \U$16150 ( \16527 , \2323 );
or \U$16151 ( \16528 , \16526 , \16527 );
or \U$16152 ( \16529 , \1141 , \14671 );
nand \U$16153 ( \16530 , \16528 , \16529 );
nand \U$16154 ( \16531 , \16530 , \14668 );
nand \U$16155 ( \16532 , \16525 , \16531 );
xor \U$16156 ( \16533 , \16522 , \16532 );
and \U$16157 ( \16534 , \16495 , \16533 );
and \U$16158 ( \16535 , \16491 , \16494 );
or \U$16159 ( \16536 , \16534 , \16535 );
not \U$16160 ( \16537 , \6091 );
and \U$16161 ( \16538 , RIae79d90_164, \5911 );
not \U$16162 ( \16539 , RIae79d90_164);
and \U$16163 ( \16540 , \16539 , \4112 );
nor \U$16164 ( \16541 , \16538 , \16540 );
not \U$16165 ( \16542 , \16541 );
or \U$16166 ( \16543 , \16537 , \16542 );
nand \U$16167 ( \16544 , \16239 , \14940 );
nand \U$16168 ( \16545 , \16543 , \16544 );
not \U$16169 ( \16546 , \4842 );
not \U$16170 ( \16547 , RIae79ca0_162);
not \U$16171 ( \16548 , \1859 );
or \U$16172 ( \16549 , \16547 , \16548 );
or \U$16173 ( \16550 , \9657 , RIae79ca0_162);
nand \U$16174 ( \16551 , \16549 , \16550 );
not \U$16175 ( \16552 , \16551 );
or \U$16176 ( \16553 , \16546 , \16552 );
nand \U$16177 ( \16554 , \16375 , \4853 );
nand \U$16178 ( \16555 , \16553 , \16554 );
nor \U$16179 ( \16556 , \16545 , \16555 );
and \U$16180 ( \16557 , \16222 , \10675 );
not \U$16181 ( \16558 , RIae7a498_179);
not \U$16182 ( \16559 , \5945 );
or \U$16183 ( \16560 , \16558 , \16559 );
not \U$16184 ( \16561 , \4194 );
or \U$16185 ( \16562 , \16561 , RIae7a498_179);
nand \U$16186 ( \16563 , \16560 , \16562 );
buf \U$16187 ( \16564 , \10695 );
and \U$16188 ( \16565 , \16563 , \16564 );
nor \U$16189 ( \16566 , \16557 , \16565 );
or \U$16190 ( \16567 , \16556 , \16566 );
nand \U$16191 ( \16568 , \16545 , \16555 );
nand \U$16192 ( \16569 , \16567 , \16568 );
xor \U$16193 ( \16570 , \16506 , \16521 );
and \U$16194 ( \16571 , \16570 , \16532 );
and \U$16195 ( \16572 , \16506 , \16521 );
or \U$16196 ( \16573 , \16571 , \16572 );
xor \U$16197 ( \16574 , \16569 , \16573 );
not \U$16198 ( \16575 , \12515 );
not \U$16199 ( \16576 , RIae7a3a8_177);
not \U$16200 ( \16577 , \10570 );
or \U$16201 ( \16578 , \16576 , \16577 );
or \U$16202 ( \16579 , \10570 , RIae7a3a8_177);
nand \U$16203 ( \16580 , \16578 , \16579 );
not \U$16204 ( \16581 , \16580 );
or \U$16205 ( \16582 , \16575 , \16581 );
nand \U$16206 ( \16583 , \16480 , \9621 );
nand \U$16207 ( \16584 , \16582 , \16583 );
not \U$16208 ( \16585 , \10275 );
not \U$16209 ( \16586 , \16452 );
or \U$16210 ( \16587 , \16585 , \16586 );
not \U$16211 ( \16588 , RIae7a8d0_188);
not \U$16212 ( \16589 , \15675 );
not \U$16213 ( \16590 , \16589 );
or \U$16214 ( \16591 , \16588 , \16590 );
or \U$16215 ( \16592 , \16589 , RIae7a8d0_188);
nand \U$16216 ( \16593 , \16591 , \16592 );
buf \U$16217 ( \16594 , \11204 );
nand \U$16218 ( \16595 , \16593 , \16594 );
nand \U$16219 ( \16596 , \16587 , \16595 );
nor \U$16220 ( \16597 , \16584 , \16596 );
not \U$16221 ( \16598 , \10510 );
not \U$16222 ( \16599 , \9529 );
not \U$16223 ( \16600 , \2917 );
or \U$16224 ( \16601 , \16599 , \16600 );
or \U$16225 ( \16602 , \1118 , \9529 );
nand \U$16226 ( \16603 , \16601 , \16602 );
not \U$16227 ( \16604 , \16603 );
or \U$16228 ( \16605 , \16598 , \16604 );
not \U$16229 ( \16606 , RIae7a7e0_186);
not \U$16230 ( \16607 , \2175 );
or \U$16231 ( \16608 , \16606 , \16607 );
or \U$16232 ( \16609 , \2175 , RIae7a7e0_186);
nand \U$16233 ( \16610 , \16608 , \16609 );
nand \U$16234 ( \16611 , \16610 , \10519 );
nand \U$16235 ( \16612 , \16605 , \16611 );
not \U$16236 ( \16613 , \16612 );
or \U$16237 ( \16614 , \16597 , \16613 );
nand \U$16238 ( \16615 , \16584 , \16596 );
nand \U$16239 ( \16616 , \16614 , \16615 );
xor \U$16240 ( \16617 , \16574 , \16616 );
xor \U$16241 ( \16618 , \16536 , \16617 );
xor \U$16242 ( \16619 , \16545 , \16555 );
xnor \U$16243 ( \16620 , \16619 , \16566 );
not \U$16244 ( \16621 , \16620 );
not \U$16245 ( \16622 , \2011 );
and \U$16246 ( \16623 , RIae79610_148, \11387 );
not \U$16247 ( \16624 , RIae79610_148);
and \U$16248 ( \16625 , \16624 , \15650 );
or \U$16249 ( \16626 , \16623 , \16625 );
not \U$16250 ( \16627 , \16626 );
or \U$16251 ( \16628 , \16622 , \16627 );
xor \U$16252 ( \16629 , RIae79610_148, \10066 );
nand \U$16253 ( \16630 , \16629 , \2063 );
nand \U$16254 ( \16631 , \16628 , \16630 );
not \U$16255 ( \16632 , \16631 );
not \U$16256 ( \16633 , RIae793b8_143);
not \U$16257 ( \16634 , \10749 );
or \U$16258 ( \16635 , \16633 , \16634 );
or \U$16259 ( \16636 , \10749 , RIae793b8_143);
nand \U$16260 ( \16637 , \16635 , \16636 );
nand \U$16261 ( \16638 , \16637 , \1910 );
and \U$16262 ( \16639 , RIae793b8_143, \10168 );
not \U$16263 ( \16640 , RIae793b8_143);
and \U$16264 ( \16641 , \16640 , \9900 );
or \U$16265 ( \16642 , \16639 , \16641 );
nand \U$16266 ( \16643 , \16642 , \1864 );
nand \U$16267 ( \16644 , \16638 , \16643 );
nand \U$16268 ( \16645 , \12857 , \926 );
not \U$16269 ( \16646 , \16645 );
not \U$16270 ( \16647 , \1072 );
not \U$16271 ( \16648 , \16164 );
not \U$16272 ( \16649 , RIae78e90_132);
and \U$16273 ( \16650 , \16648 , \16649 );
buf \U$16274 ( \16651 , \10844 );
not \U$16275 ( \16652 , \16651 );
and \U$16276 ( \16653 , \16652 , RIae78e90_132);
nor \U$16277 ( \16654 , \16650 , \16653 );
not \U$16278 ( \16655 , \16654 );
or \U$16279 ( \16656 , \16647 , \16655 );
and \U$16280 ( \16657 , \16006 , RIae78e90_132);
not \U$16281 ( \16658 , \16006 );
and \U$16282 ( \16659 , \16658 , \1066 );
or \U$16283 ( \16660 , \16657 , \16659 );
nand \U$16284 ( \16661 , \16660 , \1086 );
nand \U$16285 ( \16662 , \16656 , \16661 );
not \U$16286 ( \16663 , \16662 );
or \U$16287 ( \16664 , \16646 , \16663 );
or \U$16288 ( \16665 , \16662 , \16645 );
nand \U$16289 ( \16666 , \16664 , \16665 );
not \U$16290 ( \16667 , \838 );
not \U$16291 ( \16668 , \10272 );
not \U$16292 ( \16669 , RIae78f80_134);
and \U$16293 ( \16670 , \16668 , \16669 );
and \U$16294 ( \16671 , \11318 , RIae78f80_134);
nor \U$16295 ( \16672 , \16670 , \16671 );
not \U$16296 ( \16673 , \16672 );
or \U$16297 ( \16674 , \16667 , \16673 );
and \U$16298 ( \16675 , RIae78f80_134, \10259 );
not \U$16299 ( \16676 , RIae78f80_134);
and \U$16300 ( \16677 , \16676 , \11309 );
or \U$16301 ( \16678 , \16675 , \16677 );
nand \U$16302 ( \16679 , \16678 , \796 );
nand \U$16303 ( \16680 , \16674 , \16679 );
xor \U$16304 ( \16681 , \16666 , \16680 );
xor \U$16305 ( \16682 , \16644 , \16681 );
not \U$16306 ( \16683 , \16682 );
or \U$16307 ( \16684 , \16632 , \16683 );
not \U$16308 ( \16685 , \16643 );
not \U$16309 ( \16686 , \16638 );
or \U$16310 ( \16687 , \16685 , \16686 );
nand \U$16311 ( \16688 , \16687 , \16681 );
nand \U$16312 ( \16689 , \16684 , \16688 );
not \U$16313 ( \16690 , \4853 );
not \U$16314 ( \16691 , \16551 );
or \U$16315 ( \16692 , \16690 , \16691 );
not \U$16316 ( \16693 , RIae79ca0_162);
not \U$16317 ( \16694 , \2402 );
or \U$16318 ( \16695 , \16693 , \16694 );
or \U$16319 ( \16696 , \2402 , RIae79ca0_162);
nand \U$16320 ( \16697 , \16695 , \16696 );
nand \U$16321 ( \16698 , \16697 , \4154 );
nand \U$16322 ( \16699 , \16692 , \16698 );
not \U$16323 ( \16700 , \838 );
and \U$16324 ( \16701 , RIae78f80_134, \16036 );
not \U$16325 ( \16702 , RIae78f80_134);
and \U$16326 ( \16703 , \16702 , \11576 );
or \U$16327 ( \16704 , \16701 , \16703 );
not \U$16328 ( \16705 , \16704 );
or \U$16329 ( \16706 , \16700 , \16705 );
nand \U$16330 ( \16707 , \16672 , \796 );
nand \U$16331 ( \16708 , \16706 , \16707 );
not \U$16332 ( \16709 , \16680 );
not \U$16333 ( \16710 , \16666 );
or \U$16334 ( \16711 , \16709 , \16710 );
not \U$16335 ( \16712 , \16645 );
nand \U$16336 ( \16713 , \16712 , \16662 );
nand \U$16337 ( \16714 , \16711 , \16713 );
xor \U$16338 ( \16715 , \16708 , \16714 );
not \U$16339 ( \16716 , \1501 );
not \U$16340 ( \16717 , \16152 );
or \U$16341 ( \16718 , \16716 , \16717 );
not \U$16342 ( \16719 , \11259 );
and \U$16343 ( \16720 , \16719 , \1503 );
not \U$16344 ( \16721 , \16719 );
and \U$16345 ( \16722 , \16721 , RIae79250_140);
nor \U$16346 ( \16723 , \16720 , \16722 );
nand \U$16347 ( \16724 , \16723 , \9403 );
nand \U$16348 ( \16725 , \16718 , \16724 );
not \U$16349 ( \16726 , \16725 );
and \U$16350 ( \16727 , \16715 , \16726 );
not \U$16351 ( \16728 , \16715 );
and \U$16352 ( \16729 , \16728 , \16725 );
nor \U$16353 ( \16730 , \16727 , \16729 );
xnor \U$16354 ( \16731 , \16699 , \16730 );
and \U$16355 ( \16732 , \16689 , \16731 );
not \U$16356 ( \16733 , \16699 );
nor \U$16357 ( \16734 , \16733 , \16730 );
nor \U$16358 ( \16735 , \16732 , \16734 );
xor \U$16359 ( \16736 , \16596 , \16735 );
xor \U$16360 ( \16737 , \16584 , \16612 );
xnor \U$16361 ( \16738 , \16736 , \16737 );
not \U$16362 ( \16739 , \16738 );
or \U$16363 ( \16740 , \16621 , \16739 );
buf \U$16364 ( \16741 , \16735 );
not \U$16365 ( \16742 , \16741 );
xor \U$16366 ( \16743 , \16737 , \16596 );
nand \U$16367 ( \16744 , \16742 , \16743 );
nand \U$16368 ( \16745 , \16740 , \16744 );
xor \U$16369 ( \16746 , \16618 , \16745 );
xor \U$16370 ( \16747 , \16489 , \16746 );
not \U$16371 ( \16748 , \2251 );
not \U$16372 ( \16749 , \2268 );
not \U$16373 ( \16750 , \9609 );
or \U$16374 ( \16751 , \16749 , \16750 );
buf \U$16375 ( \16752 , \12482 );
or \U$16376 ( \16753 , \16752 , \2268 );
nand \U$16377 ( \16754 , \16751 , \16753 );
not \U$16378 ( \16755 , \16754 );
or \U$16379 ( \16756 , \16748 , \16755 );
and \U$16380 ( \16757 , \10465 , RIae79ac0_158);
not \U$16381 ( \16758 , \10465 );
and \U$16382 ( \16759 , \16758 , \2268 );
nor \U$16383 ( \16760 , \16757 , \16759 );
nand \U$16384 ( \16761 , \16760 , \2272 );
nand \U$16385 ( \16762 , \16756 , \16761 );
not \U$16386 ( \16763 , \10223 );
and \U$16387 ( \16764 , RIae79520_146, \9395 );
not \U$16388 ( \16765 , RIae79520_146);
not \U$16389 ( \16766 , \12600 );
and \U$16390 ( \16767 , \16765 , \16766 );
nor \U$16391 ( \16768 , \16764 , \16767 );
not \U$16392 ( \16769 , \16768 );
or \U$16393 ( \16770 , \16763 , \16769 );
and \U$16394 ( \16771 , RIae79520_146, \9412 );
not \U$16395 ( \16772 , RIae79520_146);
and \U$16396 ( \16773 , \16772 , \11803 );
or \U$16397 ( \16774 , \16771 , \16773 );
nand \U$16398 ( \16775 , \16774 , \12680 );
nand \U$16399 ( \16776 , \16770 , \16775 );
xor \U$16400 ( \16777 , \16762 , \16776 );
not \U$16401 ( \16778 , \1919 );
not \U$16402 ( \16779 , \3810 );
not \U$16403 ( \16780 , \12614 );
or \U$16404 ( \16781 , \16779 , \16780 );
or \U$16405 ( \16782 , \12614 , \3039 );
nand \U$16406 ( \16783 , \16781 , \16782 );
not \U$16407 ( \16784 , \16783 );
or \U$16408 ( \16785 , \16778 , \16784 );
not \U$16409 ( \16786 , \9456 );
and \U$16410 ( \16787 , \16786 , RIae794a8_145);
not \U$16411 ( \16788 , \16786 );
and \U$16412 ( \16789 , \16788 , \3039 );
nor \U$16413 ( \16790 , \16787 , \16789 );
nand \U$16414 ( \16791 , \16790 , \2457 );
nand \U$16415 ( \16792 , \16785 , \16791 );
and \U$16416 ( \16793 , \16777 , \16792 );
and \U$16417 ( \16794 , \16762 , \16776 );
nor \U$16418 ( \16795 , \16793 , \16794 );
not \U$16419 ( \16796 , \16795 );
not \U$16420 ( \16797 , \16796 );
not \U$16421 ( \16798 , \16631 );
and \U$16422 ( \16799 , \16682 , \16798 );
not \U$16423 ( \16800 , \16682 );
and \U$16424 ( \16801 , \16800 , \16631 );
nor \U$16425 ( \16802 , \16799 , \16801 );
not \U$16426 ( \16803 , \16802 );
buf \U$16427 ( \16804 , \11761 );
not \U$16428 ( \16805 , \16804 );
and \U$16429 ( \16806 , \3207 , RIae79ca0_162);
not \U$16430 ( \16807 , \3207 );
and \U$16431 ( \16808 , \16807 , \4844 );
nor \U$16432 ( \16809 , \16806 , \16808 );
not \U$16433 ( \16810 , \16809 );
or \U$16434 ( \16811 , \16805 , \16810 );
nand \U$16435 ( \16812 , \16697 , \4853 );
nand \U$16436 ( \16813 , \16811 , \16812 );
not \U$16437 ( \16814 , \1501 );
not \U$16438 ( \16815 , \16723 );
or \U$16439 ( \16816 , \16814 , \16815 );
and \U$16440 ( \16817 , RIae79250_140, \16193 );
not \U$16441 ( \16818 , RIae79250_140);
and \U$16442 ( \16819 , \16818 , \10743 );
or \U$16443 ( \16820 , \16817 , \16819 );
nand \U$16444 ( \16821 , \16820 , \1499 );
nand \U$16445 ( \16822 , \16816 , \16821 );
not \U$16446 ( \16823 , \16822 );
not \U$16447 ( \16824 , \1843 );
not \U$16448 ( \16825 , RIae79688_149);
not \U$16449 ( \16826 , \9924 );
not \U$16450 ( \16827 , \16826 );
or \U$16451 ( \16828 , \16825 , \16827 );
not \U$16452 ( \16829 , \10724 );
nand \U$16453 ( \16830 , \16829 , \5229 );
nand \U$16454 ( \16831 , \16828 , \16830 );
not \U$16455 ( \16832 , \16831 );
or \U$16456 ( \16833 , \16824 , \16832 );
not \U$16457 ( \16834 , RIae79688_149);
not \U$16458 ( \16835 , \9941 );
or \U$16459 ( \16836 , \16834 , \16835 );
not \U$16460 ( \16837 , \10461 );
nand \U$16461 ( \16838 , \16837 , \2970 );
nand \U$16462 ( \16839 , \16836 , \16838 );
nand \U$16463 ( \16840 , \16839 , \1820 );
nand \U$16464 ( \16841 , \16833 , \16840 );
not \U$16465 ( \16842 , \16841 );
not \U$16466 ( \16843 , \16842 );
or \U$16467 ( \16844 , \16823 , \16843 );
or \U$16468 ( \16845 , \16842 , \16822 );
nand \U$16469 ( \16846 , \16844 , \16845 );
and \U$16470 ( \16847 , \16813 , \16846 );
not \U$16471 ( \16848 , \16813 );
not \U$16472 ( \16849 , \16846 );
and \U$16473 ( \16850 , \16848 , \16849 );
nor \U$16474 ( \16851 , \16847 , \16850 );
not \U$16475 ( \16852 , \16851 );
or \U$16476 ( \16853 , \16803 , \16852 );
or \U$16477 ( \16854 , \16851 , \16802 );
nand \U$16478 ( \16855 , \16853 , \16854 );
not \U$16479 ( \16856 , \16855 );
or \U$16480 ( \16857 , \16797 , \16856 );
not \U$16481 ( \16858 , \16802 );
nand \U$16482 ( \16859 , \16858 , \16851 );
nand \U$16483 ( \16860 , \16857 , \16859 );
not \U$16484 ( \16861 , \16860 );
not \U$16485 ( \16862 , \4853 );
not \U$16486 ( \16863 , \16809 );
or \U$16487 ( \16864 , \16862 , \16863 );
not \U$16488 ( \16865 , RIae79ca0_162);
not \U$16489 ( \16866 , \6242 );
or \U$16490 ( \16867 , \16865 , \16866 );
or \U$16491 ( \16868 , \6238 , RIae79ca0_162);
nand \U$16492 ( \16869 , \16867 , \16868 );
nand \U$16493 ( \16870 , \16869 , \6276 );
nand \U$16494 ( \16871 , \16864 , \16870 );
not \U$16495 ( \16872 , \2450 );
not \U$16496 ( \16873 , \2447 );
not \U$16497 ( \16874 , \5722 );
or \U$16498 ( \16875 , \16873 , \16874 );
or \U$16499 ( \16876 , \9279 , \2447 );
nand \U$16500 ( \16877 , \16875 , \16876 );
not \U$16501 ( \16878 , \16877 );
or \U$16502 ( \16879 , \16872 , \16878 );
xor \U$16503 ( \16880 , RIae79778_151, \6345 );
nand \U$16504 ( \16881 , \16880 , \9576 );
nand \U$16505 ( \16882 , \16879 , \16881 );
not \U$16506 ( \16883 , \838 );
and \U$16507 ( \16884 , RIae78f80_134, \12751 );
not \U$16508 ( \16885 , RIae78f80_134);
and \U$16509 ( \16886 , \16885 , \12750 );
nor \U$16510 ( \16887 , \16884 , \16886 );
not \U$16511 ( \16888 , \16887 );
or \U$16512 ( \16889 , \16883 , \16888 );
not \U$16513 ( \16890 , \12857 );
and \U$16514 ( \16891 , \16890 , RIae78f80_134);
and \U$16515 ( \16892 , \12858 , \1132 );
nor \U$16516 ( \16893 , \16891 , \16892 );
not \U$16517 ( \16894 , \796 );
or \U$16518 ( \16895 , \16893 , \16894 );
nand \U$16519 ( \16896 , \16889 , \16895 );
not \U$16520 ( \16897 , \16896 );
not \U$16521 ( \16898 , \788 );
nand \U$16522 ( \16899 , \16898 , \12857 );
nand \U$16523 ( \16900 , \16899 , \786 , RIae78f80_134);
nor \U$16524 ( \16901 , \16897 , \16900 );
not \U$16525 ( \16902 , \1008 );
and \U$16526 ( \16903 , RIae79160_138, \10195 );
not \U$16527 ( \16904 , RIae79160_138);
and \U$16528 ( \16905 , \16904 , \10194 );
nor \U$16529 ( \16906 , \16903 , \16905 );
not \U$16530 ( \16907 , \16906 );
or \U$16531 ( \16908 , \16902 , \16907 );
not \U$16532 ( \16909 , \10042 );
and \U$16533 ( \16910 , RIae79160_138, \16909 );
not \U$16534 ( \16911 , RIae79160_138);
buf \U$16535 ( \16912 , \10042 );
and \U$16536 ( \16913 , \16911 , \16912 );
or \U$16537 ( \16914 , \16910 , \16913 );
nand \U$16538 ( \16915 , \16914 , \1012 );
nand \U$16539 ( \16916 , \16908 , \16915 );
xor \U$16540 ( \16917 , \16901 , \16916 );
not \U$16541 ( \16918 , \9403 );
not \U$16542 ( \16919 , RIae79250_140);
not \U$16543 ( \16920 , \10857 );
or \U$16544 ( \16921 , \16919 , \16920 );
not \U$16545 ( \16922 , \10856 );
or \U$16546 ( \16923 , \16922 , RIae79250_140);
nand \U$16547 ( \16924 , \16921 , \16923 );
not \U$16548 ( \16925 , \16924 );
or \U$16549 ( \16926 , \16918 , \16925 );
xor \U$16550 ( \16927 , \10142 , RIae79250_140);
nand \U$16551 ( \16928 , \16927 , \1501 );
nand \U$16552 ( \16929 , \16926 , \16928 );
and \U$16553 ( \16930 , \16917 , \16929 );
and \U$16554 ( \16931 , \16901 , \16916 );
or \U$16555 ( \16932 , \16930 , \16931 );
xor \U$16556 ( \16933 , \16882 , \16932 );
and \U$16557 ( \16934 , \16871 , \16933 );
and \U$16558 ( \16935 , \16882 , \16932 );
nor \U$16559 ( \16936 , \16934 , \16935 );
not \U$16560 ( \16937 , \16936 );
not \U$16561 ( \16938 , \16937 );
not \U$16562 ( \16939 , \1820 );
not \U$16563 ( \16940 , \16831 );
or \U$16564 ( \16941 , \16939 , \16940 );
and \U$16565 ( \16942 , \15650 , RIae79688_149);
not \U$16566 ( \16943 , \15650 );
and \U$16567 ( \16944 , \16943 , \2970 );
nor \U$16568 ( \16945 , \16942 , \16944 );
nand \U$16569 ( \16946 , \16945 , \10401 );
nand \U$16570 ( \16947 , \16941 , \16946 );
not \U$16571 ( \16948 , \16947 );
not \U$16572 ( \16949 , \1863 );
not \U$16573 ( \16950 , \16637 );
or \U$16574 ( \16951 , \16949 , \16950 );
and \U$16575 ( \16952 , RIae793b8_143, \11260 );
not \U$16576 ( \16953 , RIae793b8_143);
and \U$16577 ( \16954 , \16953 , \10007 );
or \U$16578 ( \16955 , \16952 , \16954 );
nand \U$16579 ( \16956 , \16955 , \1910 );
nand \U$16580 ( \16957 , \16951 , \16956 );
not \U$16581 ( \16958 , \16820 );
not \U$16582 ( \16959 , \16958 );
not \U$16583 ( \16960 , \1502 );
and \U$16584 ( \16961 , \16959 , \16960 );
and \U$16585 ( \16962 , \16927 , \1499 );
nor \U$16586 ( \16963 , \16961 , \16962 );
and \U$16587 ( \16964 , \16957 , \16963 );
not \U$16588 ( \16965 , \16957 );
not \U$16589 ( \16966 , \16963 );
and \U$16590 ( \16967 , \16965 , \16966 );
or \U$16591 ( \16968 , \16964 , \16967 );
not \U$16592 ( \16969 , \16968 );
or \U$16593 ( \16970 , \16948 , \16969 );
nand \U$16594 ( \16971 , \16957 , \16966 );
nand \U$16595 ( \16972 , \16970 , \16971 );
not \U$16596 ( \16973 , \16972 );
not \U$16597 ( \16974 , \16973 );
not \U$16598 ( \16975 , \2322 );
not \U$16599 ( \16976 , RIae798e0_154);
not \U$16600 ( \16977 , \12067 );
not \U$16601 ( \16978 , \16977 );
or \U$16602 ( \16979 , \16976 , \16978 );
or \U$16603 ( \16980 , \12707 , RIae798e0_154);
nand \U$16604 ( \16981 , \16979 , \16980 );
not \U$16605 ( \16982 , \16981 );
or \U$16606 ( \16983 , \16975 , \16982 );
and \U$16607 ( \16984 , \15091 , RIae798e0_154);
not \U$16608 ( \16985 , \15091 );
and \U$16609 ( \16986 , \16985 , \2981 );
nor \U$16610 ( \16987 , \16984 , \16986 );
nand \U$16611 ( \16988 , \16987 , \10807 );
nand \U$16612 ( \16989 , \16983 , \16988 );
not \U$16613 ( \16990 , \16989 );
not \U$16614 ( \16991 , \2007 );
and \U$16615 ( \16992 , RIae797f0_152, \14120 );
not \U$16616 ( \16993 , RIae797f0_152);
and \U$16617 ( \16994 , \16993 , \15220 );
or \U$16618 ( \16995 , \16992 , \16994 );
not \U$16619 ( \16996 , \16995 );
or \U$16620 ( \16997 , \16991 , \16996 );
not \U$16621 ( \16998 , RIae797f0_152);
not \U$16622 ( \16999 , \9316 );
or \U$16623 ( \17000 , \16998 , \16999 );
or \U$16624 ( \17001 , \9316 , RIae797f0_152);
nand \U$16625 ( \17002 , \17000 , \17001 );
nand \U$16626 ( \17003 , \17002 , \1988 );
nand \U$16627 ( \17004 , \16997 , \17003 );
not \U$16628 ( \17005 , \17004 );
nand \U$16629 ( \17006 , \16990 , \17005 );
not \U$16630 ( \17007 , \17006 );
not \U$16631 ( \17008 , \5324 );
not \U$16632 ( \17009 , \10226 );
not \U$16633 ( \17010 , \17009 );
and \U$16634 ( \17011 , RIae79c28_161, \17010 );
not \U$16635 ( \17012 , RIae79c28_161);
and \U$16636 ( \17013 , \17012 , \12724 );
or \U$16637 ( \17014 , \17011 , \17013 );
not \U$16638 ( \17015 , \17014 );
or \U$16639 ( \17016 , \17008 , \17015 );
and \U$16640 ( \17017 , RIae79c28_161, \13248 );
not \U$16641 ( \17018 , RIae79c28_161);
and \U$16642 ( \17019 , \17018 , \5109 );
nor \U$16643 ( \17020 , \17017 , \17019 );
not \U$16644 ( \17021 , \17020 );
nand \U$16645 ( \17022 , \17021 , \2767 );
nand \U$16646 ( \17023 , \17016 , \17022 );
not \U$16647 ( \17024 , \17023 );
or \U$16648 ( \17025 , \17007 , \17024 );
not \U$16649 ( \17026 , \17005 );
buf \U$16650 ( \17027 , \16989 );
nand \U$16651 ( \17028 , \17026 , \17027 );
nand \U$16652 ( \17029 , \17025 , \17028 );
not \U$16653 ( \17030 , \17029 );
or \U$16654 ( \17031 , \16974 , \17030 );
or \U$16655 ( \17032 , \17029 , \16973 );
nand \U$16656 ( \17033 , \17031 , \17032 );
not \U$16657 ( \17034 , \17033 );
or \U$16658 ( \17035 , \16938 , \17034 );
not \U$16659 ( \17036 , \16973 );
not \U$16660 ( \17037 , \17029 );
not \U$16661 ( \17038 , \17037 );
nand \U$16662 ( \17039 , \17036 , \17038 );
nand \U$16663 ( \17040 , \17035 , \17039 );
xor \U$16664 ( \17041 , \16731 , \16689 );
xor \U$16665 ( \17042 , \17040 , \17041 );
not \U$16666 ( \17043 , \17042 );
or \U$16667 ( \17044 , \16861 , \17043 );
buf \U$16668 ( \17045 , \17040 );
nand \U$16669 ( \17046 , \17045 , \17041 );
nand \U$16670 ( \17047 , \17044 , \17046 );
not \U$16671 ( \17048 , \17047 );
not \U$16672 ( \17049 , \14940 );
not \U$16673 ( \17050 , \16541 );
or \U$16674 ( \17051 , \17049 , \17050 );
not \U$16675 ( \17052 , \9671 );
and \U$16676 ( \17053 , RIae79d90_164, \17052 );
not \U$16677 ( \17054 , RIae79d90_164);
and \U$16678 ( \17055 , \17054 , \1969 );
nor \U$16679 ( \17056 , \17053 , \17055 );
nand \U$16680 ( \17057 , \17056 , \6091 );
nand \U$16681 ( \17058 , \17051 , \17057 );
not \U$16682 ( \17059 , \9776 );
not \U$16683 ( \17060 , \16088 );
or \U$16684 ( \17061 , \17059 , \17060 );
and \U$16685 ( \17062 , RIae7a150_172, \2047 );
not \U$16686 ( \17063 , RIae7a150_172);
and \U$16687 ( \17064 , \2040 , \2041 );
not \U$16688 ( \17065 , \2040 );
and \U$16689 ( \17066 , \17065 , \2044 );
nor \U$16690 ( \17067 , \17064 , \17066 );
not \U$16691 ( \17068 , \17067 );
and \U$16692 ( \17069 , \17063 , \17068 );
or \U$16693 ( \17070 , \17062 , \17069 );
nand \U$16694 ( \17071 , \17070 , \11087 );
nand \U$16695 ( \17072 , \17061 , \17071 );
xor \U$16696 ( \17073 , \17058 , \17072 );
not \U$16697 ( \17074 , \6214 );
not \U$16698 ( \17075 , \15991 );
or \U$16699 ( \17076 , \17074 , \17075 );
not \U$16700 ( \17077 , RIae79ef8_167);
not \U$16701 ( \17078 , \14439 );
or \U$16702 ( \17079 , \17077 , \17078 );
or \U$16703 ( \17080 , \5890 , RIae79ef8_167);
nand \U$16704 ( \17081 , \17079 , \17080 );
nand \U$16705 ( \17082 , \17081 , \15989 );
nand \U$16706 ( \17083 , \17076 , \17082 );
xor \U$16707 ( \17084 , \17073 , \17083 );
not \U$16708 ( \17085 , \17084 );
not \U$16709 ( \17086 , \10676 );
not \U$16710 ( \17087 , \16563 );
or \U$16711 ( \17088 , \17086 , \17087 );
and \U$16712 ( \17089 , RIae7a498_179, \1898 );
not \U$16713 ( \17090 , RIae7a498_179);
and \U$16714 ( \17091 , \17090 , \13086 );
nor \U$16715 ( \17092 , \17089 , \17091 );
nand \U$16716 ( \17093 , \17092 , \16564 );
nand \U$16717 ( \17094 , \17088 , \17093 );
not \U$16718 ( \17095 , \9622 );
not \U$16719 ( \17096 , \16580 );
or \U$16720 ( \17097 , \17095 , \17096 );
not \U$16721 ( \17098 , RIae7a3a8_177);
not \U$16722 ( \17099 , \2153 );
or \U$16723 ( \17100 , \17098 , \17099 );
or \U$16724 ( \17101 , \14712 , RIae7a3a8_177);
nand \U$16725 ( \17102 , \17100 , \17101 );
nand \U$16726 ( \17103 , \17102 , \9644 );
nand \U$16727 ( \17104 , \17097 , \17103 );
xor \U$16728 ( \17105 , \17094 , \17104 );
not \U$16729 ( \17106 , \10519 );
not \U$16730 ( \17107 , \16603 );
or \U$16731 ( \17108 , \17106 , \17107 );
not \U$16732 ( \17109 , \9529 );
not \U$16733 ( \17110 , \1124 );
or \U$16734 ( \17111 , \17109 , \17110 );
not \U$16735 ( \17112 , RIae7a7e0_186);
or \U$16736 ( \17113 , \1124 , \17112 );
nand \U$16737 ( \17114 , \17111 , \17113 );
nand \U$16738 ( \17115 , \17114 , \11851 );
nand \U$16739 ( \17116 , \17108 , \17115 );
not \U$16740 ( \17117 , \17116 );
xnor \U$16741 ( \17118 , \17105 , \17117 );
not \U$16742 ( \17119 , \11434 );
xor \U$16743 ( \17120 , RIae7a498_179, \2628 );
not \U$16744 ( \17121 , \17120 );
or \U$16745 ( \17122 , \17119 , \17121 );
nand \U$16746 ( \17123 , \17092 , \10676 );
nand \U$16747 ( \17124 , \17122 , \17123 );
xor \U$16748 ( \17125 , \1100 , RIae7a6f0_184);
xnor \U$16749 ( \17126 , \17125 , \1112 );
not \U$16750 ( \17127 , \17126 );
not \U$16751 ( \17128 , \9473 );
or \U$16752 ( \17129 , \17127 , \17128 );
not \U$16753 ( \17130 , \877 );
xor \U$16754 ( \17131 , RIae7a6f0_184, \17130 );
nand \U$16755 ( \17132 , \17131 , \9705 );
nand \U$16756 ( \17133 , \17129 , \17132 );
xor \U$16757 ( \17134 , \17124 , \17133 );
not \U$16758 ( \17135 , \1049 );
and \U$16759 ( \17136 , RIae79070_136, \16035 );
not \U$16760 ( \17137 , RIae79070_136);
and \U$16761 ( \17138 , \17137 , \16036 );
nor \U$16762 ( \17139 , \17136 , \17138 );
not \U$16763 ( \17140 , \17139 );
or \U$16764 ( \17141 , \17135 , \17140 );
xor \U$16765 ( \17142 , RIae79070_136, \10272 );
nand \U$16766 ( \17143 , \17142 , \1062 );
nand \U$16767 ( \17144 , \17141 , \17143 );
not \U$16768 ( \17145 , \1049 );
not \U$16769 ( \17146 , \17142 );
or \U$16770 ( \17147 , \17145 , \17146 );
not \U$16771 ( \17148 , \10259 );
not \U$16772 ( \17149 , RIae79070_136);
or \U$16773 ( \17150 , \17148 , \17149 );
not \U$16774 ( \17151 , \10252 );
and \U$16775 ( \17152 , \10254 , \17151 );
not \U$16776 ( \17153 , \10254 );
and \U$16777 ( \17154 , \17153 , \10252 );
or \U$16778 ( \17155 , \17152 , \17154 );
or \U$16779 ( \17156 , \17155 , RIae79070_136);
nand \U$16780 ( \17157 , \17150 , \17156 );
nand \U$16781 ( \17158 , \17157 , \1061 );
nand \U$16782 ( \17159 , \17147 , \17158 );
not \U$16783 ( \17160 , \17159 );
and \U$16784 ( \17161 , \12857 , \1072 );
not \U$16785 ( \17162 , \838 );
not \U$16786 ( \17163 , \16165 );
not \U$16787 ( \17164 , \3105 );
and \U$16788 ( \17165 , \17163 , \17164 );
not \U$16789 ( \17166 , \10845 );
and \U$16790 ( \17167 , \17166 , \1132 );
nor \U$16791 ( \17168 , \17165 , \17167 );
not \U$16792 ( \17169 , \17168 );
or \U$16793 ( \17170 , \17162 , \17169 );
nand \U$16794 ( \17171 , \16887 , \796 );
nand \U$16795 ( \17172 , \17170 , \17171 );
xor \U$16796 ( \17173 , \17161 , \17172 );
not \U$16797 ( \17174 , \17173 );
or \U$16798 ( \17175 , \17160 , \17174 );
nand \U$16799 ( \17176 , \17172 , \17161 );
nand \U$16800 ( \17177 , \17175 , \17176 );
xor \U$16801 ( \17178 , \17144 , \17177 );
not \U$16802 ( \17179 , \2011 );
not \U$16803 ( \17180 , \16629 );
or \U$16804 ( \17181 , \17179 , \17180 );
not \U$16805 ( \17182 , \2056 );
not \U$16806 ( \17183 , \13544 );
or \U$16807 ( \17184 , \17182 , \17183 );
not \U$16808 ( \17185 , \10168 );
or \U$16809 ( \17186 , \17185 , \11150 );
nand \U$16810 ( \17187 , \17184 , \17186 );
nand \U$16811 ( \17188 , \17187 , \2063 );
nand \U$16812 ( \17189 , \17181 , \17188 );
and \U$16813 ( \17190 , \17178 , \17189 );
and \U$16814 ( \17191 , \17144 , \17177 );
nor \U$16815 ( \17192 , \17190 , \17191 );
not \U$16816 ( \17193 , \17192 );
and \U$16817 ( \17194 , \17134 , \17193 );
and \U$16818 ( \17195 , \17124 , \17133 );
or \U$16819 ( \17196 , \17194 , \17195 );
and \U$16820 ( \17197 , \17118 , \17196 );
not \U$16821 ( \17198 , \17118 );
not \U$16822 ( \17199 , \17196 );
and \U$16823 ( \17200 , \17198 , \17199 );
nor \U$16824 ( \17201 , \17197 , \17200 );
not \U$16825 ( \17202 , \17201 );
or \U$16826 ( \17203 , \17085 , \17202 );
buf \U$16827 ( \17204 , \17118 );
not \U$16828 ( \17205 , \17199 );
nand \U$16829 ( \17206 , \17204 , \17205 );
nand \U$16830 ( \17207 , \17203 , \17206 );
not \U$16831 ( \17208 , \17207 );
not \U$16832 ( \17209 , \16002 );
not \U$16833 ( \17210 , \16020 );
or \U$16834 ( \17211 , \17209 , \17210 );
or \U$16835 ( \17212 , \16020 , \16002 );
nand \U$16836 ( \17213 , \17211 , \17212 );
not \U$16837 ( \17214 , \17213 );
not \U$16838 ( \17215 , \1072 );
not \U$16839 ( \17216 , \16187 );
or \U$16840 ( \17217 , \17215 , \17216 );
nand \U$16841 ( \17218 , \16654 , \1086 );
nand \U$16842 ( \17219 , \17217 , \17218 );
not \U$16843 ( \17220 , \17219 );
not \U$16844 ( \17221 , \17220 );
or \U$16845 ( \17222 , \17214 , \17221 );
or \U$16846 ( \17223 , \17220 , \17213 );
nand \U$16847 ( \17224 , \17222 , \17223 );
not \U$16848 ( \17225 , \17224 );
not \U$16849 ( \17226 , \1049 );
not \U$16850 ( \17227 , \16054 );
or \U$16851 ( \17228 , \17226 , \17227 );
and \U$16852 ( \17229 , RIae79070_136, \10046 );
not \U$16853 ( \17230 , RIae79070_136);
and \U$16854 ( \17231 , \17230 , \10042 );
nor \U$16855 ( \17232 , \17229 , \17231 );
not \U$16856 ( \17233 , \17232 );
nand \U$16857 ( \17234 , \17233 , \1062 );
nand \U$16858 ( \17235 , \17228 , \17234 );
not \U$16859 ( \17236 , \17235 );
or \U$16860 ( \17237 , \17225 , \17236 );
nand \U$16861 ( \17238 , \17219 , \17213 );
nand \U$16862 ( \17239 , \17237 , \17238 );
not \U$16863 ( \17240 , \2339 );
not \U$16864 ( \17241 , RIae798e0_154);
not \U$16865 ( \17242 , \6230 );
not \U$16866 ( \17243 , \17242 );
or \U$16867 ( \17244 , \17241 , \17243 );
not \U$16868 ( \17245 , \9298 );
or \U$16869 ( \17246 , \17245 , RIae798e0_154);
nand \U$16870 ( \17247 , \17244 , \17246 );
not \U$16871 ( \17248 , \17247 );
or \U$16872 ( \17249 , \17240 , \17248 );
nand \U$16873 ( \17250 , \16326 , \2321 );
nand \U$16874 ( \17251 , \17249 , \17250 );
xor \U$16875 ( \17252 , \17239 , \17251 );
not \U$16876 ( \17253 , \2007 );
not \U$16877 ( \17254 , \16315 );
or \U$16878 ( \17255 , \17253 , \17254 );
not \U$16879 ( \17256 , \2521 );
not \U$16880 ( \17257 , \9279 );
or \U$16881 ( \17258 , \17256 , \17257 );
or \U$16882 ( \17259 , \9279 , \1991 );
nand \U$16883 ( \17260 , \17258 , \17259 );
nand \U$16884 ( \17261 , \17260 , \1988 );
nand \U$16885 ( \17262 , \17255 , \17261 );
xor \U$16886 ( \17263 , \17252 , \17262 );
xor \U$16887 ( \17264 , \17058 , \17072 );
and \U$16888 ( \17265 , \17264 , \17083 );
and \U$16889 ( \17266 , \17058 , \17072 );
or \U$16890 ( \17267 , \17265 , \17266 );
not \U$16891 ( \17268 , \17267 );
xor \U$16892 ( \17269 , \17263 , \17268 );
not \U$16893 ( \17270 , RIae7aab0_192);
not \U$16894 ( \17271 , \16530 );
or \U$16895 ( \17272 , \17270 , \17271 );
and \U$16896 ( \17273 , RIae7aa38_191, \2330 );
not \U$16897 ( \17274 , RIae7aa38_191);
and \U$16898 ( \17275 , \17274 , \1158 );
nor \U$16899 ( \17276 , \17273 , \17275 );
nand \U$16900 ( \17277 , \17276 , \14667 );
nand \U$16901 ( \17278 , \17272 , \17277 );
not \U$16902 ( \17279 , \9699 );
not \U$16903 ( \17280 , \16500 );
or \U$16904 ( \17281 , \17279 , \17280 );
and \U$16905 ( \17282 , RIae7a240_174, \2286 );
not \U$16906 ( \17283 , RIae7a240_174);
and \U$16907 ( \17284 , \17283 , \3747 );
or \U$16908 ( \17285 , \17282 , \17284 );
nand \U$16909 ( \17286 , \17285 , \9688 );
nand \U$16910 ( \17287 , \17281 , \17286 );
or \U$16911 ( \17288 , \17278 , \17287 );
not \U$16912 ( \17289 , \9745 );
not \U$16913 ( \17290 , \16519 );
or \U$16914 ( \17291 , \17289 , \17290 );
and \U$16915 ( \17292 , RIae7a060_170, \1405 );
not \U$16916 ( \17293 , RIae7a060_170);
and \U$16917 ( \17294 , \17293 , \9625 );
or \U$16918 ( \17295 , \17292 , \17294 );
nand \U$16919 ( \17296 , \17295 , \9730 );
nand \U$16920 ( \17297 , \17291 , \17296 );
nand \U$16921 ( \17298 , \17288 , \17297 );
nand \U$16922 ( \17299 , \17278 , \17287 );
nand \U$16923 ( \17300 , \17298 , \17299 );
xor \U$16924 ( \17301 , \17269 , \17300 );
nand \U$16925 ( \17302 , \17208 , \17301 );
not \U$16926 ( \17303 , \17302 );
or \U$16927 ( \17304 , \17048 , \17303 );
buf \U$16928 ( \17305 , \17207 );
not \U$16929 ( \17306 , \17301 );
nand \U$16930 ( \17307 , \17305 , \17306 );
nand \U$16931 ( \17308 , \17304 , \17307 );
and \U$16932 ( \17309 , \16747 , \17308 );
and \U$16933 ( \17310 , \16489 , \16746 );
or \U$16934 ( \17311 , \17309 , \17310 );
not \U$16935 ( \17312 , \10401 );
and \U$16936 ( \17313 , \9608 , \2970 );
not \U$16937 ( \17314 , \9608 );
and \U$16938 ( \17315 , \17314 , RIae79688_149);
nor \U$16939 ( \17316 , \17313 , \17315 );
not \U$16940 ( \17317 , \17316 );
or \U$16941 ( \17318 , \17312 , \17317 );
nand \U$16942 ( \17319 , \15949 , \1820 );
nand \U$16943 ( \17320 , \17318 , \17319 );
not \U$16944 ( \17321 , \17320 );
not \U$16945 ( \17322 , \17321 );
not \U$16946 ( \17323 , \10927 );
not \U$16947 ( \17324 , RIae7a510_180);
not \U$16948 ( \17325 , \17324 );
not \U$16949 ( \17326 , \12206 );
or \U$16950 ( \17327 , \17325 , \17326 );
or \U$16951 ( \17328 , \12206 , \14931 );
nand \U$16952 ( \17329 , \17327 , \17328 );
not \U$16953 ( \17330 , \17329 );
or \U$16954 ( \17331 , \17323 , \17330 );
nand \U$16955 ( \17332 , \16365 , \10631 );
nand \U$16956 ( \17333 , \17331 , \17332 );
not \U$16957 ( \17334 , \17333 );
not \U$16958 ( \17335 , \17334 );
or \U$16959 ( \17336 , \17322 , \17335 );
not \U$16960 ( \17337 , \2417 );
not \U$16961 ( \17338 , \10331 );
not \U$16962 ( \17339 , \17338 );
not \U$16963 ( \17340 , RIae79c28_161);
and \U$16964 ( \17341 , \17339 , \17340 );
and \U$16965 ( \17342 , \4982 , RIae79c28_161);
nor \U$16966 ( \17343 , \17341 , \17342 );
not \U$16967 ( \17344 , \17343 );
or \U$16968 ( \17345 , \17337 , \17344 );
and \U$16969 ( \17346 , \10584 , \10492 );
not \U$16970 ( \17347 , \10584 );
and \U$16971 ( \17348 , \17347 , \3269 );
nor \U$16972 ( \17349 , \17346 , \17348 );
nand \U$16973 ( \17350 , \17349 , \2776 );
nand \U$16974 ( \17351 , \17345 , \17350 );
nand \U$16975 ( \17352 , \17336 , \17351 );
nand \U$16976 ( \17353 , \17333 , \17320 );
nand \U$16977 ( \17354 , \17352 , \17353 );
not \U$16978 ( \17355 , \17354 );
not \U$16979 ( \17356 , \2272 );
and \U$16980 ( \17357 , RIae79ac0_158, \12603 );
not \U$16981 ( \17358 , RIae79ac0_158);
and \U$16982 ( \17359 , \17358 , \12600 );
or \U$16983 ( \17360 , \17357 , \17359 );
not \U$16984 ( \17361 , \17360 );
or \U$16985 ( \17362 , \17356 , \17361 );
nand \U$16986 ( \17363 , \16290 , \10414 );
nand \U$16987 ( \17364 , \17362 , \17363 );
not \U$16988 ( \17365 , \17364 );
not \U$16989 ( \17366 , \10223 );
not \U$16990 ( \17367 , \16256 );
or \U$16991 ( \17368 , \17366 , \17367 );
not \U$16992 ( \17369 , \2183 );
not \U$16993 ( \17370 , \9438 );
or \U$16994 ( \17371 , \17369 , \17370 );
or \U$16995 ( \17372 , \9441 , \2183 );
nand \U$16996 ( \17373 , \17371 , \17372 );
nand \U$16997 ( \17374 , \17373 , \2602 );
nand \U$16998 ( \17375 , \17368 , \17374 );
not \U$16999 ( \17376 , \17375 );
or \U$17000 ( \17377 , \17365 , \17376 );
not \U$17001 ( \17378 , \17375 );
not \U$17002 ( \17379 , \17378 );
not \U$17003 ( \17380 , \17364 );
not \U$17004 ( \17381 , \17380 );
or \U$17005 ( \17382 , \17379 , \17381 );
not \U$17006 ( \17383 , \2457 );
not \U$17007 ( \17384 , RIae794a8_145);
not \U$17008 ( \17385 , \16977 );
or \U$17009 ( \17386 , \17384 , \17385 );
buf \U$17010 ( \17387 , \9347 );
or \U$17011 ( \17388 , \17387 , RIae794a8_145);
nand \U$17012 ( \17389 , \17386 , \17388 );
not \U$17013 ( \17390 , \17389 );
or \U$17014 ( \17391 , \17383 , \17390 );
nand \U$17015 ( \17392 , \16276 , \2467 );
nand \U$17016 ( \17393 , \17391 , \17392 );
nand \U$17017 ( \17394 , \17382 , \17393 );
nand \U$17018 ( \17395 , \17377 , \17394 );
not \U$17019 ( \17396 , \17395 );
not \U$17020 ( \17397 , \1864 );
and \U$17021 ( \17398 , RIae793b8_143, \12644 );
not \U$17022 ( \17399 , RIae793b8_143);
buf \U$17023 ( \17400 , \16826 );
and \U$17024 ( \17401 , \17399 , \17400 );
nor \U$17025 ( \17402 , \17398 , \17401 );
not \U$17026 ( \17403 , \17402 );
or \U$17027 ( \17404 , \17397 , \17403 );
not \U$17028 ( \17405 , RIae793b8_143);
not \U$17029 ( \17406 , \10208 );
not \U$17030 ( \17407 , \17406 );
or \U$17031 ( \17408 , \17405 , \17407 );
nand \U$17032 ( \17409 , \10208 , \1902 );
nand \U$17033 ( \17410 , \17408 , \17409 );
nand \U$17034 ( \17411 , \17410 , \1910 );
nand \U$17035 ( \17412 , \17404 , \17411 );
not \U$17036 ( \17413 , \1501 );
and \U$17037 ( \17414 , RIae79250_140, \10066 );
not \U$17038 ( \17415 , RIae79250_140);
and \U$17039 ( \17416 , \17415 , \11562 );
nor \U$17040 ( \17417 , \17414 , \17416 );
not \U$17041 ( \17418 , \17417 );
or \U$17042 ( \17419 , \17413 , \17418 );
nand \U$17043 ( \17420 , \16159 , \1497 );
nand \U$17044 ( \17421 , \17419 , \17420 );
not \U$17045 ( \17422 , \9947 );
not \U$17046 ( \17423 , \9989 );
and \U$17047 ( \17424 , RIae79070_136, \17423 );
not \U$17048 ( \17425 , RIae79070_136);
and \U$17049 ( \17426 , \17425 , \16193 );
nor \U$17050 ( \17427 , \17424 , \17426 );
not \U$17051 ( \17428 , \17427 );
or \U$17052 ( \17429 , \17422 , \17428 );
not \U$17053 ( \17430 , \1249 );
nand \U$17054 ( \17431 , \17430 , \16061 );
nand \U$17055 ( \17432 , \17429 , \17431 );
xor \U$17056 ( \17433 , \17421 , \17432 );
xnor \U$17057 ( \17434 , \17412 , \17433 );
not \U$17058 ( \17435 , \17434 );
and \U$17059 ( \17436 , \17396 , \17435 );
and \U$17060 ( \17437 , \17395 , \17434 );
nor \U$17061 ( \17438 , \17436 , \17437 );
not \U$17062 ( \17439 , \17438 );
not \U$17063 ( \17440 , \17439 );
or \U$17064 ( \17441 , \17355 , \17440 );
not \U$17065 ( \17442 , \17434 );
nand \U$17066 ( \17443 , \17442 , \17395 );
nand \U$17067 ( \17444 , \17441 , \17443 );
not \U$17068 ( \17445 , \17444 );
not \U$17069 ( \17446 , \16317 );
not \U$17070 ( \17447 , \16339 );
or \U$17071 ( \17448 , \17446 , \17447 );
nand \U$17072 ( \17449 , \16334 , \16323 );
nand \U$17073 ( \17450 , \17448 , \17449 );
not \U$17074 ( \17451 , \16258 );
not \U$17075 ( \17452 , \16297 );
or \U$17076 ( \17453 , \17451 , \17452 );
nand \U$17077 ( \17454 , \16292 , \16278 );
nand \U$17078 ( \17455 , \17453 , \17454 );
xor \U$17079 ( \17456 , \17450 , \17455 );
buf \U$17080 ( \17457 , \15951 );
not \U$17081 ( \17458 , \17457 );
nand \U$17082 ( \17459 , \17458 , \15965 );
not \U$17083 ( \17460 , \17459 );
not \U$17084 ( \17461 , \15982 );
or \U$17085 ( \17462 , \17460 , \17461 );
not \U$17086 ( \17463 , \15965 );
nand \U$17087 ( \17464 , \17463 , \17457 );
nand \U$17088 ( \17465 , \17462 , \17464 );
not \U$17089 ( \17466 , \17465 );
and \U$17090 ( \17467 , \17456 , \17466 );
not \U$17091 ( \17468 , \17456 );
and \U$17092 ( \17469 , \17468 , \17465 );
nor \U$17093 ( \17470 , \17467 , \17469 );
not \U$17094 ( \17471 , \17470 );
or \U$17095 ( \17472 , \17445 , \17471 );
or \U$17096 ( \17473 , \17470 , \17444 );
nand \U$17097 ( \17474 , \17472 , \17473 );
not \U$17098 ( \17475 , \16424 );
nand \U$17099 ( \17476 , \17475 , \16434 );
not \U$17100 ( \17477 , \17476 );
not \U$17101 ( \17478 , \16413 );
or \U$17102 ( \17479 , \17477 , \17478 );
not \U$17103 ( \17480 , \17475 );
nand \U$17104 ( \17481 , \17480 , \16433 );
nand \U$17105 ( \17482 , \17479 , \17481 );
not \U$17106 ( \17483 , \16135 );
not \U$17107 ( \17484 , \9804 );
not \U$17108 ( \17485 , \2309 );
or \U$17109 ( \17486 , \17484 , \17485 );
or \U$17110 ( \17487 , \2309 , \9799 );
nand \U$17111 ( \17488 , \17486 , \17487 );
not \U$17112 ( \17489 , \17488 );
or \U$17113 ( \17490 , \17483 , \17489 );
nand \U$17114 ( \17491 , \16134 , \9792 );
nand \U$17115 ( \17492 , \17490 , \17491 );
not \U$17116 ( \17493 , \17492 );
not \U$17117 ( \17494 , \17493 );
not \U$17118 ( \17495 , \9745 );
xor \U$17119 ( \17496 , RIae7a060_170, \2917 );
not \U$17120 ( \17497 , \17496 );
or \U$17121 ( \17498 , \17495 , \17497 );
nand \U$17122 ( \17499 , \16512 , \9730 );
nand \U$17123 ( \17500 , \17498 , \17499 );
not \U$17124 ( \17501 , \17500 );
not \U$17125 ( \17502 , \17501 );
or \U$17126 ( \17503 , \17494 , \17502 );
not \U$17127 ( \17504 , \17492 );
not \U$17128 ( \17505 , \17500 );
or \U$17129 ( \17506 , \17504 , \17505 );
buf \U$17130 ( \17507 , \9705 );
not \U$17131 ( \17508 , \17507 );
not \U$17132 ( \17509 , RIae7a6f0_184);
not \U$17133 ( \17510 , \1439 );
or \U$17134 ( \17511 , \17509 , \17510 );
or \U$17135 ( \17512 , \919 , RIae7a6f0_184);
nand \U$17136 ( \17513 , \17511 , \17512 );
not \U$17137 ( \17514 , \17513 );
or \U$17138 ( \17515 , \17508 , \17514 );
nand \U$17139 ( \17516 , \16112 , \9473 );
nand \U$17140 ( \17517 , \17515 , \17516 );
not \U$17141 ( \17518 , \17517 );
nand \U$17142 ( \17519 , \17506 , \17518 );
nand \U$17143 ( \17520 , \17503 , \17519 );
not \U$17144 ( \17521 , \17520 );
xor \U$17145 ( \17522 , \17482 , \17521 );
not \U$17146 ( \17523 , \16367 );
not \U$17147 ( \17524 , \17523 );
not \U$17148 ( \17525 , \16399 );
not \U$17149 ( \17526 , \17525 );
or \U$17150 ( \17527 , \17524 , \17526 );
not \U$17151 ( \17528 , \16367 );
not \U$17152 ( \17529 , \16399 );
or \U$17153 ( \17530 , \17528 , \17529 );
nand \U$17154 ( \17531 , \17530 , \16377 );
nand \U$17155 ( \17532 , \17527 , \17531 );
not \U$17156 ( \17533 , \17532 );
and \U$17157 ( \17534 , \17522 , \17533 );
not \U$17158 ( \17535 , \17522 );
and \U$17159 ( \17536 , \17535 , \17532 );
nor \U$17160 ( \17537 , \17534 , \17536 );
and \U$17161 ( \17538 , \17474 , \17537 );
not \U$17162 ( \17539 , \17474 );
not \U$17163 ( \17540 , \17537 );
and \U$17164 ( \17541 , \17539 , \17540 );
nor \U$17165 ( \17542 , \17538 , \17541 );
xor \U$17166 ( \17543 , \16536 , \16617 );
and \U$17167 ( \17544 , \17543 , \16745 );
and \U$17168 ( \17545 , \16536 , \16617 );
or \U$17169 ( \17546 , \17544 , \17545 );
xor \U$17170 ( \17547 , \17542 , \17546 );
xor \U$17171 ( \17548 , \16569 , \16573 );
and \U$17172 ( \17549 , \17548 , \16616 );
and \U$17173 ( \17550 , \16569 , \16573 );
or \U$17174 ( \17551 , \17549 , \17550 );
not \U$17175 ( \17552 , \17551 );
not \U$17176 ( \17553 , \16143 );
not \U$17177 ( \17554 , \16093 );
or \U$17178 ( \17555 , \17553 , \17554 );
nand \U$17179 ( \17556 , \17555 , \15986 );
not \U$17180 ( \17557 , \16093 );
nand \U$17181 ( \17558 , \17557 , \16144 );
nand \U$17182 ( \17559 , \17556 , \17558 );
buf \U$17183 ( \17560 , \17559 );
not \U$17184 ( \17561 , \17560 );
not \U$17185 ( \17562 , \1062 );
not \U$17186 ( \17563 , \17427 );
or \U$17187 ( \17564 , \17562 , \17563 );
nand \U$17188 ( \17565 , \14539 , \1049 );
nand \U$17189 ( \17566 , \17564 , \17565 );
xor \U$17190 ( \17567 , \12866 , \12854 );
xor \U$17191 ( \17568 , \17566 , \17567 );
not \U$17192 ( \17569 , \1008 );
and \U$17193 ( \17570 , \9875 , \997 );
not \U$17194 ( \17571 , \9875 );
and \U$17195 ( \17572 , \17571 , RIae79160_138);
nor \U$17196 ( \17573 , \17570 , \17572 );
not \U$17197 ( \17574 , \17573 );
or \U$17198 ( \17575 , \17569 , \17574 );
nand \U$17199 ( \17576 , \14547 , \1012 );
nand \U$17200 ( \17577 , \17575 , \17576 );
xnor \U$17201 ( \17578 , \17568 , \17577 );
not \U$17202 ( \17579 , \1910 );
not \U$17203 ( \17580 , \17402 );
or \U$17204 ( \17581 , \17579 , \17580 );
nand \U$17205 ( \17582 , \14404 , \1863 );
nand \U$17206 ( \17583 , \17581 , \17582 );
and \U$17207 ( \17584 , \12890 , \1501 );
and \U$17208 ( \17585 , \17417 , \1499 );
nor \U$17209 ( \17586 , \17584 , \17585 );
xnor \U$17210 ( \17587 , \17583 , \17586 );
xor \U$17211 ( \17588 , \17578 , \17587 );
not \U$17212 ( \17589 , \2322 );
not \U$17213 ( \17590 , \14579 );
or \U$17214 ( \17591 , \17589 , \17590 );
nand \U$17215 ( \17592 , \16332 , \14580 );
nand \U$17216 ( \17593 , \17591 , \17592 );
xnor \U$17217 ( \17594 , \17588 , \17593 );
not \U$17218 ( \17595 , \10584 );
not \U$17219 ( \17596 , \1859 );
not \U$17220 ( \17597 , \17596 );
or \U$17221 ( \17598 , \17595 , \17597 );
nand \U$17222 ( \17599 , \9657 , RIae79c28_161);
nand \U$17223 ( \17600 , \17598 , \17599 );
nand \U$17224 ( \17601 , \17600 , \2776 );
not \U$17225 ( \17602 , \838 );
not \U$17226 ( \17603 , \14595 );
or \U$17227 ( \17604 , \17602 , \17603 );
nand \U$17228 ( \17605 , \16028 , \797 );
nand \U$17229 ( \17606 , \17604 , \17605 );
not \U$17230 ( \17607 , \14603 );
not \U$17231 ( \17608 , \14610 );
or \U$17232 ( \17609 , \17607 , \17608 );
or \U$17233 ( \17610 , \14610 , \14603 );
nand \U$17234 ( \17611 , \17609 , \17610 );
not \U$17235 ( \17612 , \12852 );
not \U$17236 ( \17613 , \926 );
or \U$17237 ( \17614 , \17612 , \17613 );
not \U$17238 ( \17615 , \16170 );
or \U$17239 ( \17616 , \17615 , \950 );
nand \U$17240 ( \17617 , \17614 , \17616 );
xor \U$17241 ( \17618 , \17611 , \17617 );
xnor \U$17242 ( \17619 , \17606 , \17618 );
nand \U$17243 ( \17620 , \17349 , \2767 );
nand \U$17244 ( \17621 , \17601 , \17619 , \17620 );
not \U$17245 ( \17622 , \17621 );
not \U$17246 ( \17623 , \9527 );
xor \U$17247 ( \17624 , RIae7a7e0_186, \854 );
not \U$17248 ( \17625 , \17624 );
or \U$17249 ( \17626 , \17623 , \17625 );
nand \U$17250 ( \17627 , \16610 , \11439 );
nand \U$17251 ( \17628 , \17626 , \17627 );
not \U$17252 ( \17629 , \17628 );
or \U$17253 ( \17630 , \17622 , \17629 );
not \U$17254 ( \17631 , \17620 );
not \U$17255 ( \17632 , \17601 );
or \U$17256 ( \17633 , \17631 , \17632 );
not \U$17257 ( \17634 , \17619 );
nand \U$17258 ( \17635 , \17633 , \17634 );
nand \U$17259 ( \17636 , \17630 , \17635 );
not \U$17260 ( \17637 , \17636 );
and \U$17261 ( \17638 , \17594 , \17637 );
not \U$17262 ( \17639 , \17594 );
and \U$17263 ( \17640 , \17639 , \17636 );
nor \U$17264 ( \17641 , \17638 , \17640 );
not \U$17265 ( \17642 , \17641 );
not \U$17266 ( \17643 , \17642 );
or \U$17267 ( \17644 , \17561 , \17643 );
or \U$17268 ( \17645 , \17560 , \17642 );
nand \U$17269 ( \17646 , \17644 , \17645 );
not \U$17270 ( \17647 , \17646 );
or \U$17271 ( \17648 , \17552 , \17647 );
or \U$17272 ( \17649 , \17551 , \17646 );
nand \U$17273 ( \17650 , \17648 , \17649 );
xor \U$17274 ( \17651 , \17547 , \17650 );
xor \U$17275 ( \17652 , \17311 , \17651 );
and \U$17276 ( \17653 , \17635 , \17621 );
xor \U$17277 ( \17654 , \17653 , \17628 );
xor \U$17278 ( \17655 , \17493 , \17518 );
xnor \U$17279 ( \17656 , \17655 , \17501 );
xor \U$17280 ( \17657 , \17654 , \17656 );
not \U$17281 ( \17658 , \2163 );
not \U$17282 ( \17659 , \17373 );
or \U$17283 ( \17660 , \17658 , \17659 );
and \U$17284 ( \17661 , RIae79520_146, \10361 );
not \U$17285 ( \17662 , RIae79520_146);
and \U$17286 ( \17663 , \17662 , \9459 );
or \U$17287 ( \17664 , \17661 , \17663 );
nand \U$17288 ( \17665 , \17664 , \12680 );
nand \U$17289 ( \17666 , \17660 , \17665 );
not \U$17290 ( \17667 , \2322 );
not \U$17291 ( \17668 , \17247 );
or \U$17292 ( \17669 , \17667 , \17668 );
not \U$17293 ( \17670 , RIae798e0_154);
not \U$17294 ( \17671 , \16271 );
or \U$17295 ( \17672 , \17670 , \17671 );
or \U$17296 ( \17673 , \9316 , RIae798e0_154);
nand \U$17297 ( \17674 , \17672 , \17673 );
nand \U$17298 ( \17675 , \17674 , \2339 );
nand \U$17299 ( \17676 , \17669 , \17675 );
xor \U$17300 ( \17677 , \17666 , \17676 );
not \U$17301 ( \17678 , \1919 );
not \U$17302 ( \17679 , \17389 );
or \U$17303 ( \17680 , \17678 , \17679 );
not \U$17304 ( \17681 , \9367 );
not \U$17305 ( \17682 , \3810 );
or \U$17306 ( \17683 , \17681 , \17682 );
or \U$17307 ( \17684 , \15091 , \3810 );
nand \U$17308 ( \17685 , \17683 , \17684 );
nand \U$17309 ( \17686 , \17685 , \1933 );
nand \U$17310 ( \17687 , \17680 , \17686 );
and \U$17311 ( \17688 , \17677 , \17687 );
and \U$17312 ( \17689 , \17666 , \17676 );
or \U$17313 ( \17690 , \17688 , \17689 );
not \U$17314 ( \17691 , \1820 );
not \U$17315 ( \17692 , \17316 );
or \U$17316 ( \17693 , \17691 , \17692 );
nand \U$17317 ( \17694 , \16839 , \1843 );
nand \U$17318 ( \17695 , \17693 , \17694 );
not \U$17319 ( \17696 , \17695 );
not \U$17320 ( \17697 , \2251 );
not \U$17321 ( \17698 , \17360 );
or \U$17322 ( \17699 , \17697 , \17698 );
not \U$17323 ( \17700 , RIae79ac0_158);
not \U$17324 ( \17701 , \9417 );
or \U$17325 ( \17702 , \17700 , \17701 );
or \U$17326 ( \17703 , \11195 , RIae79ac0_158);
nand \U$17327 ( \17704 , \17702 , \17703 );
nand \U$17328 ( \17705 , \17704 , \2272 );
nand \U$17329 ( \17706 , \17699 , \17705 );
not \U$17330 ( \17707 , \17706 );
nand \U$17331 ( \17708 , \17696 , \17707 );
not \U$17332 ( \17709 , \17708 );
not \U$17333 ( \17710 , \2767 );
not \U$17334 ( \17711 , \6238 );
not \U$17335 ( \17712 , RIae79c28_161);
and \U$17336 ( \17713 , \17711 , \17712 );
and \U$17337 ( \17714 , \6238 , RIae79c28_161);
nor \U$17338 ( \17715 , \17713 , \17714 );
not \U$17339 ( \17716 , \17715 );
not \U$17340 ( \17717 , \17716 );
or \U$17341 ( \17718 , \17710 , \17717 );
nand \U$17342 ( \17719 , \17343 , \5324 );
nand \U$17343 ( \17720 , \17718 , \17719 );
not \U$17344 ( \17721 , \17720 );
or \U$17345 ( \17722 , \17709 , \17721 );
nand \U$17346 ( \17723 , \17706 , \17695 );
nand \U$17347 ( \17724 , \17722 , \17723 );
xor \U$17348 ( \17725 , \17690 , \17724 );
not \U$17349 ( \17726 , \1910 );
and \U$17350 ( \17727 , RIae793b8_143, \11230 );
not \U$17351 ( \17728 , RIae793b8_143);
and \U$17352 ( \17729 , \17728 , \10066 );
or \U$17353 ( \17730 , \17727 , \17729 );
not \U$17354 ( \17731 , \17730 );
or \U$17355 ( \17732 , \17726 , \17731 );
nand \U$17356 ( \17733 , \17410 , \1863 );
nand \U$17357 ( \17734 , \17732 , \17733 );
not \U$17358 ( \17735 , \2063 );
and \U$17359 ( \17736 , RIae79610_148, \12644 );
not \U$17360 ( \17737 , RIae79610_148);
and \U$17361 ( \17738 , \17737 , \10725 );
nor \U$17362 ( \17739 , \17736 , \17738 );
not \U$17363 ( \17740 , \17739 );
or \U$17364 ( \17741 , \17735 , \17740 );
nand \U$17365 ( \17742 , \15960 , \2011 );
nand \U$17366 ( \17743 , \17741 , \17742 );
xor \U$17367 ( \17744 , \17734 , \17743 );
not \U$17368 ( \17745 , \2450 );
not \U$17369 ( \17746 , \15980 );
or \U$17370 ( \17747 , \17745 , \17746 );
not \U$17371 ( \17748 , RIae79778_151);
not \U$17372 ( \17749 , \10829 );
or \U$17373 ( \17750 , \17748 , \17749 );
or \U$17374 ( \17751 , \10829 , RIae79778_151);
nand \U$17375 ( \17752 , \17750 , \17751 );
nand \U$17376 ( \17753 , \17752 , \2545 );
nand \U$17377 ( \17754 , \17747 , \17753 );
xor \U$17378 ( \17755 , \17744 , \17754 );
and \U$17379 ( \17756 , \17725 , \17755 );
and \U$17380 ( \17757 , \17690 , \17724 );
or \U$17381 ( \17758 , \17756 , \17757 );
and \U$17382 ( \17759 , \17657 , \17758 );
and \U$17383 ( \17760 , \17654 , \17656 );
or \U$17384 ( \17761 , \17759 , \17760 );
not \U$17385 ( \17762 , \16228 );
not \U$17386 ( \17763 , \16241 );
or \U$17387 ( \17764 , \17762 , \17763 );
not \U$17388 ( \17765 , \16209 );
nand \U$17389 ( \17766 , \17765 , \16224 );
nand \U$17390 ( \17767 , \17764 , \17766 );
not \U$17391 ( \17768 , \10638 );
not \U$17392 ( \17769 , \16356 );
or \U$17393 ( \17770 , \17768 , \17769 );
nand \U$17394 ( \17771 , \14496 , \16358 );
nand \U$17395 ( \17772 , \17770 , \17771 );
not \U$17396 ( \17773 , \11851 );
not \U$17397 ( \17774 , \17624 );
or \U$17398 ( \17775 , \17773 , \17774 );
nand \U$17399 ( \17776 , \14374 , \10519 );
nand \U$17400 ( \17777 , \17775 , \17776 );
xor \U$17401 ( \17778 , \17772 , \17777 );
not \U$17402 ( \17779 , \14667 );
not \U$17403 ( \17780 , \16397 );
or \U$17404 ( \17781 , \17779 , \17780 );
nand \U$17405 ( \17782 , \14676 , RIae7aab0_192);
nand \U$17406 ( \17783 , \17781 , \17782 );
xor \U$17407 ( \17784 , \17778 , \17783 );
xor \U$17408 ( \17785 , \17767 , \17784 );
not \U$17409 ( \17786 , \9814 );
not \U$17410 ( \17787 , \14714 );
or \U$17411 ( \17788 , \17786 , \17787 );
nand \U$17412 ( \17789 , \17488 , \9792 );
nand \U$17413 ( \17790 , \17788 , \17789 );
not \U$17414 ( \17791 , \9473 );
not \U$17415 ( \17792 , \17513 );
or \U$17416 ( \17793 , \17791 , \17792 );
nand \U$17417 ( \17794 , \14738 , \9478 );
nand \U$17418 ( \17795 , \17793 , \17794 );
xor \U$17419 ( \17796 , \17790 , \17795 );
buf \U$17420 ( \17797 , \9730 );
not \U$17421 ( \17798 , \17797 );
not \U$17422 ( \17799 , \17496 );
or \U$17423 ( \17800 , \17798 , \17799 );
nand \U$17424 ( \17801 , \14726 , \11098 );
nand \U$17425 ( \17802 , \17800 , \17801 );
xor \U$17426 ( \17803 , \17796 , \17802 );
xnor \U$17427 ( \17804 , \17785 , \17803 );
and \U$17428 ( \17805 , \17761 , \17804 );
not \U$17429 ( \17806 , \17761 );
not \U$17430 ( \17807 , \17804 );
and \U$17431 ( \17808 , \17806 , \17807 );
or \U$17432 ( \17809 , \17805 , \17808 );
not \U$17433 ( \17810 , \16804 );
not \U$17434 ( \17811 , \16373 );
or \U$17435 ( \17812 , \17810 , \17811 );
nand \U$17436 ( \17813 , \14441 , \4853 );
nand \U$17437 ( \17814 , \17812 , \17813 );
not \U$17438 ( \17815 , \6091 );
not \U$17439 ( \17816 , \16233 );
or \U$17440 ( \17817 , \17815 , \17816 );
nand \U$17441 ( \17818 , \14450 , \5048 );
nand \U$17442 ( \17819 , \17817 , \17818 );
xor \U$17443 ( \17820 , \17814 , \17819 );
not \U$17444 ( \17821 , \12371 );
not \U$17445 ( \17822 , \14466 );
or \U$17446 ( \17823 , \17821 , \17822 );
nand \U$17447 ( \17824 , \16215 , \16564 );
nand \U$17448 ( \17825 , \17823 , \17824 );
xor \U$17449 ( \17826 , \17820 , \17825 );
not \U$17450 ( \17827 , \16466 );
not \U$17451 ( \17828 , \16454 );
or \U$17452 ( \17829 , \17827 , \17828 );
or \U$17453 ( \17830 , \16466 , \16454 );
nand \U$17454 ( \17831 , \17830 , \16482 );
nand \U$17455 ( \17832 , \17829 , \17831 );
and \U$17456 ( \17833 , \17826 , \17832 );
not \U$17457 ( \17834 , \17826 );
not \U$17458 ( \17835 , \17832 );
and \U$17459 ( \17836 , \17834 , \17835 );
or \U$17460 ( \17837 , \17833 , \17836 );
not \U$17461 ( \17838 , \11014 );
not \U$17462 ( \17839 , \16473 );
or \U$17463 ( \17840 , \17838 , \17839 );
nand \U$17464 ( \17841 , \14384 , \9621 );
nand \U$17465 ( \17842 , \17840 , \17841 );
not \U$17466 ( \17843 , \17842 );
not \U$17467 ( \17844 , \10275 );
not \U$17468 ( \17845 , \14509 );
or \U$17469 ( \17846 , \17844 , \17845 );
buf \U$17470 ( \17847 , \11204 );
nand \U$17471 ( \17848 , \16445 , \17847 );
nand \U$17472 ( \17849 , \17846 , \17848 );
not \U$17473 ( \17850 , \13121 );
not \U$17474 ( \17851 , \14389 );
or \U$17475 ( \17852 , \17850 , \17851 );
nand \U$17476 ( \17853 , \16456 , \13720 );
nand \U$17477 ( \17854 , \17852 , \17853 );
and \U$17478 ( \17855 , \17849 , \17854 );
not \U$17479 ( \17856 , \17849 );
not \U$17480 ( \17857 , \17854 );
and \U$17481 ( \17858 , \17856 , \17857 );
nor \U$17482 ( \17859 , \17855 , \17858 );
not \U$17483 ( \17860 , \17859 );
not \U$17484 ( \17861 , \17860 );
or \U$17485 ( \17862 , \17843 , \17861 );
not \U$17486 ( \17863 , \17842 );
nand \U$17487 ( \17864 , \17863 , \17859 );
nand \U$17488 ( \17865 , \17862 , \17864 );
xor \U$17489 ( \17866 , \17837 , \17865 );
and \U$17490 ( \17867 , \17809 , \17866 );
not \U$17491 ( \17868 , \17809 );
not \U$17492 ( \17869 , \17866 );
and \U$17493 ( \17870 , \17868 , \17869 );
nor \U$17494 ( \17871 , \17867 , \17870 );
not \U$17495 ( \17872 , \16345 );
not \U$17496 ( \17873 , \16242 );
not \U$17497 ( \17874 , \17873 );
or \U$17498 ( \17875 , \17872 , \17874 );
nand \U$17499 ( \17876 , \16298 , \16341 );
nand \U$17500 ( \17877 , \17875 , \17876 );
xor \U$17501 ( \17878 , \16403 , \16439 );
and \U$17502 ( \17879 , \17878 , \16483 );
and \U$17503 ( \17880 , \16403 , \16439 );
or \U$17504 ( \17881 , \17879 , \17880 );
xor \U$17505 ( \17882 , \17877 , \17881 );
not \U$17506 ( \17883 , \10414 );
not \U$17507 ( \17884 , \14695 );
or \U$17508 ( \17885 , \17883 , \17884 );
nand \U$17509 ( \17886 , \16284 , \2272 );
nand \U$17510 ( \17887 , \17885 , \17886 );
not \U$17511 ( \17888 , \10401 );
not \U$17512 ( \17889 , \15937 );
or \U$17513 ( \17890 , \17888 , \17889 );
nand \U$17514 ( \17891 , \14661 , \1820 );
nand \U$17515 ( \17892 , \17890 , \17891 );
not \U$17516 ( \17893 , \17892 );
xor \U$17517 ( \17894 , \17887 , \17893 );
not \U$17518 ( \17895 , \5950 );
not \U$17519 ( \17896 , \16249 );
or \U$17520 ( \17897 , \17895 , \17896 );
nand \U$17521 ( \17898 , \14646 , \3440 );
nand \U$17522 ( \17899 , \17897 , \17898 );
xnor \U$17523 ( \17900 , \17894 , \17899 );
and \U$17524 ( \17901 , \17606 , \17618 );
and \U$17525 ( \17902 , \17611 , \17617 );
nor \U$17526 ( \17903 , \17901 , \17902 );
not \U$17527 ( \17904 , \1919 );
not \U$17528 ( \17905 , \14633 );
or \U$17529 ( \17906 , \17904 , \17905 );
nand \U$17530 ( \17907 , \16264 , \9828 );
nand \U$17531 ( \17908 , \17906 , \17907 );
xor \U$17532 ( \17909 , \17903 , \17908 );
not \U$17533 ( \17910 , \1988 );
not \U$17534 ( \17911 , \16306 );
or \U$17535 ( \17912 , \17910 , \17911 );
nand \U$17536 ( \17913 , \14561 , \2007 );
nand \U$17537 ( \17914 , \17912 , \17913 );
xnor \U$17538 ( \17915 , \17909 , \17914 );
xor \U$17539 ( \17916 , \17900 , \17915 );
not \U$17540 ( \17917 , \2011 );
not \U$17541 ( \17918 , \14413 );
or \U$17542 ( \17919 , \17917 , \17918 );
nand \U$17543 ( \17920 , \15953 , \9370 );
nand \U$17544 ( \17921 , \17919 , \17920 );
not \U$17545 ( \17922 , \2418 );
not \U$17546 ( \17923 , \14426 );
or \U$17547 ( \17924 , \17922 , \17923 );
nand \U$17548 ( \17925 , \17600 , \2767 );
nand \U$17549 ( \17926 , \17924 , \17925 );
not \U$17550 ( \17927 , \17926 );
xor \U$17551 ( \17928 , \17921 , \17927 );
not \U$17552 ( \17929 , \9576 );
not \U$17553 ( \17930 , \15973 );
or \U$17554 ( \17931 , \17929 , \17930 );
nand \U$17555 ( \17932 , \14489 , \2450 );
nand \U$17556 ( \17933 , \17931 , \17932 );
not \U$17557 ( \17934 , \17933 );
xnor \U$17558 ( \17935 , \17928 , \17934 );
xnor \U$17559 ( \17936 , \17916 , \17935 );
xor \U$17560 ( \17937 , \17882 , \17936 );
not \U$17561 ( \17938 , \16484 );
not \U$17562 ( \17939 , \16354 );
or \U$17563 ( \17940 , \17938 , \17939 );
or \U$17564 ( \17941 , \16350 , \16148 );
nand \U$17565 ( \17942 , \17940 , \17941 );
and \U$17566 ( \17943 , \17937 , \17942 );
not \U$17567 ( \17944 , \17937 );
not \U$17568 ( \17945 , \17942 );
and \U$17569 ( \17946 , \17944 , \17945 );
nor \U$17570 ( \17947 , \17943 , \17946 );
not \U$17571 ( \17948 , \17947 );
xor \U$17572 ( \17949 , \17871 , \17948 );
xor \U$17573 ( \17950 , \17652 , \17949 );
not \U$17574 ( \17951 , \1007 );
not \U$17575 ( \17952 , \997 );
not \U$17576 ( \17953 , \10338 );
or \U$17577 ( \17954 , \17952 , \17953 );
not \U$17578 ( \17955 , \10032 );
nand \U$17579 ( \17956 , \17955 , RIae79160_138);
nand \U$17580 ( \17957 , \17954 , \17956 );
not \U$17581 ( \17958 , \17957 );
or \U$17582 ( \17959 , \17951 , \17958 );
and \U$17583 ( \17960 , RIae79160_138, \10149 );
not \U$17584 ( \17961 , RIae79160_138);
and \U$17585 ( \17962 , \17961 , \10142 );
or \U$17586 ( \17963 , \17960 , \17962 );
nand \U$17587 ( \17964 , \17963 , \1012 );
nand \U$17588 ( \17965 , \17959 , \17964 );
not \U$17589 ( \17966 , \1072 );
not \U$17590 ( \17967 , \16660 );
or \U$17591 ( \17968 , \17966 , \17967 );
and \U$17592 ( \17969 , RIae78e90_132, \12857 );
not \U$17593 ( \17970 , RIae78e90_132);
not \U$17594 ( \17971 , \12857 );
and \U$17595 ( \17972 , \17970 , \17971 );
nor \U$17596 ( \17973 , \17969 , \17972 );
nand \U$17597 ( \17974 , \17973 , \1086 );
nand \U$17598 ( \17975 , \17968 , \17974 );
or \U$17599 ( \17976 , \3105 , \1083 );
or \U$17600 ( \17977 , RIae78f08_133, RIae78f80_134);
nand \U$17601 ( \17978 , \17977 , \12857 );
nand \U$17602 ( \17979 , \17976 , \17978 , RIae78e90_132);
not \U$17603 ( \17980 , \17979 );
and \U$17604 ( \17981 , \17975 , \17980 );
not \U$17605 ( \17982 , \17981 );
nor \U$17606 ( \17983 , \17232 , \1203 );
and \U$17607 ( \17984 , \17139 , \1061 );
nor \U$17608 ( \17985 , \17983 , \17984 );
not \U$17609 ( \17986 , \17985 );
or \U$17610 ( \17987 , \17982 , \17986 );
not \U$17611 ( \17988 , \17984 );
not \U$17612 ( \17989 , \17988 );
not \U$17613 ( \17990 , \17232 );
nand \U$17614 ( \17991 , \17990 , \1049 );
not \U$17615 ( \17992 , \17991 );
or \U$17616 ( \17993 , \17989 , \17992 );
not \U$17617 ( \17994 , \17981 );
nand \U$17618 ( \17995 , \17993 , \17994 );
nand \U$17619 ( \17996 , \17987 , \17995 );
xor \U$17620 ( \17997 , \17965 , \17996 );
not \U$17621 ( \17998 , \6091 );
not \U$17622 ( \17999 , RIae79d90_164);
not \U$17623 ( \18000 , \9657 );
or \U$17624 ( \18001 , \17999 , \18000 );
or \U$17625 ( \18002 , \1859 , RIae79d90_164);
nand \U$17626 ( \18003 , \18001 , \18002 );
not \U$17627 ( \18004 , \18003 );
or \U$17628 ( \18005 , \17998 , \18004 );
nand \U$17629 ( \18006 , \17056 , \5048 );
nand \U$17630 ( \18007 , \18005 , \18006 );
xor \U$17631 ( \18008 , \17997 , \18007 );
not \U$17632 ( \18009 , \6201 );
not \U$17633 ( \18010 , RIae79ef8_167);
not \U$17634 ( \18011 , \4112 );
or \U$17635 ( \18012 , \18010 , \18011 );
or \U$17636 ( \18013 , \4112 , RIae79ef8_167);
nand \U$17637 ( \18014 , \18012 , \18013 );
not \U$17638 ( \18015 , \18014 );
or \U$17639 ( \18016 , \18009 , \18015 );
nand \U$17640 ( \18017 , \17081 , \6214 );
nand \U$17641 ( \18018 , \18016 , \18017 );
xor \U$17642 ( \18019 , \18008 , \18018 );
not \U$17643 ( \18020 , \9776 );
not \U$17644 ( \18021 , \17070 );
or \U$17645 ( \18022 , \18020 , \18021 );
xor \U$17646 ( \18023 , RIae7a150_172, \5944 );
nand \U$17647 ( \18024 , \18023 , \10667 );
nand \U$17648 ( \18025 , \18022 , \18024 );
not \U$17649 ( \18026 , \10700 );
not \U$17650 ( \18027 , RIae79fe8_169);
not \U$17651 ( \18028 , \18027 );
not \U$17652 ( \18029 , \1788 );
not \U$17653 ( \18030 , \18029 );
or \U$17654 ( \18031 , \18028 , \18030 );
or \U$17655 ( \18032 , \11680 , \11069 );
nand \U$17656 ( \18033 , \18031 , \18032 );
not \U$17657 ( \18034 , \18033 );
or \U$17658 ( \18035 , \18026 , \18034 );
not \U$17659 ( \18036 , \9504 );
not \U$17660 ( \18037 , \11512 );
or \U$17661 ( \18038 , \18036 , \18037 );
or \U$17662 ( \18039 , \2675 , \11069 );
nand \U$17663 ( \18040 , \18038 , \18039 );
nand \U$17664 ( \18041 , \18040 , \11913 );
nand \U$17665 ( \18042 , \18035 , \18041 );
xor \U$17666 ( \18043 , \18025 , \18042 );
not \U$17667 ( \18044 , \17276 );
not \U$17668 ( \18045 , RIae7aab0_192);
or \U$17669 ( \18046 , \18044 , \18045 );
not \U$17670 ( \18047 , RIae7aa38_191);
not \U$17671 ( \18048 , \1439 );
or \U$17672 ( \18049 , \18047 , \18048 );
or \U$17673 ( \18050 , \1439 , RIae7aa38_191);
nand \U$17674 ( \18051 , \18049 , \18050 );
not \U$17675 ( \18052 , \18051 );
not \U$17676 ( \18053 , \14667 );
or \U$17677 ( \18054 , \18052 , \18053 );
nand \U$17678 ( \18055 , \18046 , \18054 );
xor \U$17679 ( \18056 , \18043 , \18055 );
xor \U$17680 ( \18057 , \18019 , \18056 );
not \U$17681 ( \18058 , \9621 );
not \U$17682 ( \18059 , \17102 );
or \U$17683 ( \18060 , \18058 , \18059 );
not \U$17684 ( \18061 , \11690 );
not \U$17685 ( \18062 , \2309 );
or \U$17686 ( \18063 , \18061 , \18062 );
or \U$17687 ( \18064 , \2309 , \13165 );
nand \U$17688 ( \18065 , \18063 , \18064 );
nand \U$17689 ( \18066 , \18065 , \12515 );
nand \U$17690 ( \18067 , \18060 , \18066 );
not \U$17691 ( \18068 , \11439 );
not \U$17692 ( \18069 , RIae7a7e0_186);
not \U$17693 ( \18070 , \11538 );
or \U$17694 ( \18071 , \18069 , \18070 );
or \U$17695 ( \18072 , \11538 , RIae7a7e0_186);
nand \U$17696 ( \18073 , \18071 , \18072 );
not \U$17697 ( \18074 , \18073 );
or \U$17698 ( \18075 , \18068 , \18074 );
nand \U$17699 ( \18076 , \17114 , \10519 );
nand \U$17700 ( \18077 , \18075 , \18076 );
not \U$17701 ( \18078 , \14510 );
and \U$17702 ( \18079 , RIae7a8d0_188, \9761 );
not \U$17703 ( \18080 , RIae7a8d0_188);
and \U$17704 ( \18081 , \18080 , \1022 );
nor \U$17705 ( \18082 , \18079 , \18081 );
not \U$17706 ( \18083 , \18082 );
or \U$17707 ( \18084 , \18078 , \18083 );
not \U$17708 ( \18085 , \11207 );
not \U$17709 ( \18086 , \937 );
or \U$17710 ( \18087 , \18085 , \18086 );
not \U$17711 ( \18088 , RIae7a8d0_188);
or \U$17712 ( \18089 , \9770 , \18088 );
nand \U$17713 ( \18090 , \18087 , \18089 );
nand \U$17714 ( \18091 , \18090 , \10275 );
nand \U$17715 ( \18092 , \18084 , \18091 );
xor \U$17716 ( \18093 , \18077 , \18092 );
xor \U$17717 ( \18094 , \18067 , \18093 );
and \U$17718 ( \18095 , \18057 , \18094 );
and \U$17719 ( \18096 , \18019 , \18056 );
or \U$17720 ( \18097 , \18095 , \18096 );
not \U$17721 ( \18098 , \18097 );
not \U$17722 ( \18099 , \2450 );
not \U$17723 ( \18100 , \17752 );
or \U$17724 ( \18101 , \18099 , \18100 );
and \U$17725 ( \18102 , RIae79778_151, \16310 );
not \U$17726 ( \18103 , RIae79778_151);
and \U$17727 ( \18104 , \18103 , \6256 );
nor \U$17728 ( \18105 , \18102 , \18104 );
not \U$17729 ( \18106 , \18105 );
nand \U$17730 ( \18107 , \18106 , \2432 );
nand \U$17731 ( \18108 , \18101 , \18107 );
not \U$17732 ( \18109 , \9289 );
not \U$17733 ( \18110 , RIae797f0_152);
and \U$17734 ( \18111 , \18109 , \18110 );
and \U$17735 ( \18112 , \6345 , RIae797f0_152);
nor \U$17736 ( \18113 , \18111 , \18112 );
nand \U$17737 ( \18114 , \18113 , \1988 );
nand \U$17738 ( \18115 , \17260 , \2007 );
nand \U$17739 ( \18116 , \18114 , \18115 );
not \U$17740 ( \18117 , \17965 );
not \U$17741 ( \18118 , \17996 );
or \U$17742 ( \18119 , \18117 , \18118 );
not \U$17743 ( \18120 , \17988 );
not \U$17744 ( \18121 , \17991 );
or \U$17745 ( \18122 , \18120 , \18121 );
nand \U$17746 ( \18123 , \18122 , \17981 );
nand \U$17747 ( \18124 , \18119 , \18123 );
xor \U$17748 ( \18125 , \18116 , \18124 );
xor \U$17749 ( \18126 , \18108 , \18125 );
not \U$17750 ( \18127 , \2457 );
not \U$17751 ( \18128 , \16783 );
or \U$17752 ( \18129 , \18127 , \18128 );
nand \U$17753 ( \18130 , \17685 , \2467 );
nand \U$17754 ( \18131 , \18129 , \18130 );
not \U$17755 ( \18132 , \2272 );
not \U$17756 ( \18133 , \16754 );
or \U$17757 ( \18134 , \18132 , \18133 );
nand \U$17758 ( \18135 , \17704 , \2249 );
nand \U$17759 ( \18136 , \18134 , \18135 );
or \U$17760 ( \18137 , \18131 , \18136 );
not \U$17761 ( \18138 , \18137 );
not \U$17762 ( \18139 , \10927 );
not \U$17763 ( \18140 , RIae7a510_180);
not \U$17764 ( \18141 , \2140 );
or \U$17765 ( \18142 , \18140 , \18141 );
or \U$17766 ( \18143 , \2136 , RIae7a510_180);
nand \U$17767 ( \18144 , \18142 , \18143 );
not \U$17768 ( \18145 , \18144 );
or \U$17769 ( \18146 , \18139 , \18145 );
and \U$17770 ( \18147 , \2230 , \10646 );
not \U$17771 ( \18148 , \2230 );
and \U$17772 ( \18149 , \18148 , RIae7a510_180);
nor \U$17773 ( \18150 , \18147 , \18149 );
nand \U$17774 ( \18151 , \18150 , \10631 );
nand \U$17775 ( \18152 , \18146 , \18151 );
not \U$17776 ( \18153 , \18152 );
or \U$17777 ( \18154 , \18138 , \18153 );
nand \U$17778 ( \18155 , \18131 , \18136 );
nand \U$17779 ( \18156 , \18154 , \18155 );
xor \U$17780 ( \18157 , \18126 , \18156 );
xor \U$17781 ( \18158 , \17695 , \17707 );
xnor \U$17782 ( \18159 , \18158 , \17720 );
xor \U$17783 ( \18160 , \18157 , \18159 );
and \U$17784 ( \18161 , \1012 , \16198 );
and \U$17785 ( \18162 , \17963 , \1007 );
nor \U$17786 ( \18163 , \18161 , \18162 );
and \U$17787 ( \18164 , \17730 , \1864 );
not \U$17788 ( \18165 , \16642 );
nor \U$17789 ( \18166 , \18165 , \6846 );
nor \U$17790 ( \18167 , \18164 , \18166 );
xor \U$17791 ( \18168 , \18163 , \18167 );
and \U$17792 ( \18169 , \2011 , \17739 );
and \U$17793 ( \18170 , \16626 , \2063 );
nor \U$17794 ( \18171 , \18169 , \18170 );
xor \U$17795 ( \18172 , \18168 , \18171 );
xor \U$17796 ( \18173 , \17997 , \18007 );
and \U$17797 ( \18174 , \18173 , \18018 );
and \U$17798 ( \18175 , \17997 , \18007 );
or \U$17799 ( \18176 , \18174 , \18175 );
xor \U$17800 ( \18177 , \18172 , \18176 );
xor \U$17801 ( \18178 , \17666 , \17676 );
xor \U$17802 ( \18179 , \18178 , \17687 );
xnor \U$17803 ( \18180 , \18177 , \18179 );
or \U$17804 ( \18181 , \18160 , \18180 );
not \U$17805 ( \18182 , \18181 );
or \U$17806 ( \18183 , \18098 , \18182 );
nand \U$17807 ( \18184 , \18160 , \18180 );
nand \U$17808 ( \18185 , \18183 , \18184 );
not \U$17809 ( \18186 , \18185 );
xor \U$17810 ( \18187 , \18126 , \18156 );
and \U$17811 ( \18188 , \18187 , \18159 );
and \U$17812 ( \18189 , \18126 , \18156 );
or \U$17813 ( \18190 , \18188 , \18189 );
not \U$17814 ( \18191 , \18190 );
xor \U$17815 ( \18192 , \17690 , \17724 );
xor \U$17816 ( \18193 , \18192 , \17755 );
not \U$17817 ( \18194 , \18193 );
not \U$17818 ( \18195 , \18194 );
or \U$17819 ( \18196 , \18191 , \18195 );
not \U$17820 ( \18197 , \18190 );
nand \U$17821 ( \18198 , \18197 , \18193 );
nand \U$17822 ( \18199 , \18196 , \18198 );
xor \U$17823 ( \18200 , \18025 , \18042 );
and \U$17824 ( \18201 , \18200 , \18055 );
and \U$17825 ( \18202 , \18025 , \18042 );
or \U$17826 ( \18203 , \18201 , \18202 );
not \U$17827 ( \18204 , \13720 );
and \U$17828 ( \18205 , RIae7a240_174, \1741 );
not \U$17829 ( \18206 , RIae7a240_174);
and \U$17830 ( \18207 , \18206 , \3099 );
or \U$17831 ( \18208 , \18205 , \18207 );
not \U$17832 ( \18209 , \18208 );
or \U$17833 ( \18210 , \18204 , \18209 );
nand \U$17834 ( \18211 , \17285 , \13121 );
nand \U$17835 ( \18212 , \18210 , \18211 );
not \U$17836 ( \18213 , \18212 );
xor \U$17837 ( \18214 , RIae7a2b8_175, \1808 );
not \U$17838 ( \18215 , \18214 );
not \U$17839 ( \18216 , \9792 );
or \U$17840 ( \18217 , \18215 , \18216 );
not \U$17841 ( \18218 , \9799 );
not \U$17842 ( \18219 , \1753 );
or \U$17843 ( \18220 , \18218 , \18219 );
nand \U$17844 ( \18221 , \1758 , RIae7a2b8_175);
nand \U$17845 ( \18222 , \18220 , \18221 );
nand \U$17846 ( \18223 , \18222 , \9814 );
nand \U$17847 ( \18224 , \18217 , \18223 );
not \U$17848 ( \18225 , \18224 );
or \U$17849 ( \18226 , \18213 , \18225 );
or \U$17850 ( \18227 , \18224 , \18212 );
not \U$17851 ( \18228 , \9745 );
not \U$17852 ( \18229 , \17295 );
or \U$17853 ( \18230 , \18228 , \18229 );
xor \U$17854 ( \18231 , RIae7a060_170, \2025 );
nand \U$17855 ( \18232 , \18231 , \9730 );
nand \U$17856 ( \18233 , \18230 , \18232 );
nand \U$17857 ( \18234 , \18227 , \18233 );
nand \U$17858 ( \18235 , \18226 , \18234 );
nand \U$17859 ( \18236 , \18203 , \18235 );
not \U$17860 ( \18237 , \18236 );
nand \U$17861 ( \18238 , \18093 , \18067 );
nand \U$17862 ( \18239 , \18092 , \18077 );
and \U$17863 ( \18240 , \18238 , \18239 );
not \U$17864 ( \18241 , \18240 );
or \U$17865 ( \18242 , \18237 , \18241 );
not \U$17866 ( \18243 , \18235 );
not \U$17867 ( \18244 , \18203 );
nand \U$17868 ( \18245 , \18243 , \18244 );
nand \U$17869 ( \18246 , \18242 , \18245 );
not \U$17870 ( \18247 , \18246 );
and \U$17871 ( \18248 , \18199 , \18247 );
not \U$17872 ( \18249 , \18199 );
and \U$17873 ( \18250 , \18249 , \18246 );
nor \U$17874 ( \18251 , \18248 , \18250 );
not \U$17875 ( \18252 , \18251 );
not \U$17876 ( \18253 , \16846 );
not \U$17877 ( \18254 , \16813 );
or \U$17878 ( \18255 , \18253 , \18254 );
not \U$17879 ( \18256 , \16842 );
nand \U$17880 ( \18257 , \18256 , \16822 );
nand \U$17881 ( \18258 , \18255 , \18257 );
not \U$17882 ( \18259 , \17715 );
not \U$17883 ( \18260 , \5323 );
and \U$17884 ( \18261 , \18259 , \18260 );
and \U$17885 ( \18262 , \17014 , \2767 );
nor \U$17886 ( \18263 , \18261 , \18262 );
not \U$17887 ( \18264 , \18263 );
not \U$17888 ( \18265 , \14580 );
not \U$17889 ( \18266 , \16981 );
or \U$17890 ( \18267 , \18265 , \18266 );
nand \U$17891 ( \18268 , \17674 , \2322 );
nand \U$17892 ( \18269 , \18267 , \18268 );
not \U$17893 ( \18270 , \12680 );
not \U$17894 ( \18271 , \16768 );
or \U$17895 ( \18272 , \18270 , \18271 );
nand \U$17896 ( \18273 , \17664 , \3440 );
nand \U$17897 ( \18274 , \18272 , \18273 );
nand \U$17898 ( \18275 , \18269 , \18274 );
not \U$17899 ( \18276 , \18275 );
or \U$17900 ( \18277 , \18264 , \18276 );
or \U$17901 ( \18278 , \18269 , \18274 );
nand \U$17902 ( \18279 , \18277 , \18278 );
xor \U$17903 ( \18280 , \18258 , \18279 );
not \U$17904 ( \18281 , \1988 );
not \U$17905 ( \18282 , \16995 );
or \U$17906 ( \18283 , \18281 , \18282 );
nand \U$17907 ( \18284 , \18113 , \2007 );
nand \U$17908 ( \18285 , \18283 , \18284 );
not \U$17909 ( \18286 , \18285 );
not \U$17910 ( \18287 , \17975 );
not \U$17911 ( \18288 , \17979 );
and \U$17912 ( \18289 , \18287 , \18288 );
and \U$17913 ( \18290 , \17975 , \17979 );
nor \U$17914 ( \18291 , \18289 , \18290 );
not \U$17915 ( \18292 , \18291 );
not \U$17916 ( \18293 , \838 );
not \U$17917 ( \18294 , \16678 );
or \U$17918 ( \18295 , \18293 , \18294 );
nand \U$17919 ( \18296 , \17168 , \796 );
nand \U$17920 ( \18297 , \18295 , \18296 );
not \U$17921 ( \18298 , \18297 );
or \U$17922 ( \18299 , \18292 , \18298 );
or \U$17923 ( \18300 , \18297 , \18291 );
nand \U$17924 ( \18301 , \18299 , \18300 );
not \U$17925 ( \18302 , \18301 );
not \U$17926 ( \18303 , \1012 );
not \U$17927 ( \18304 , \17957 );
or \U$17928 ( \18305 , \18303 , \18304 );
nand \U$17929 ( \18306 , \16914 , \1008 );
nand \U$17930 ( \18307 , \18305 , \18306 );
not \U$17931 ( \18308 , \18307 );
or \U$17932 ( \18309 , \18302 , \18308 );
not \U$17933 ( \18310 , \18291 );
nand \U$17934 ( \18311 , \18310 , \18297 );
nand \U$17935 ( \18312 , \18309 , \18311 );
not \U$17936 ( \18313 , \18312 );
not \U$17937 ( \18314 , \2450 );
nor \U$17938 ( \18315 , \18105 , \18314 );
and \U$17939 ( \18316 , \16877 , \2432 );
nor \U$17940 ( \18317 , \18315 , \18316 );
not \U$17941 ( \18318 , \18317 );
or \U$17942 ( \18319 , \18313 , \18318 );
not \U$17943 ( \18320 , \18316 );
not \U$17944 ( \18321 , \18320 );
not \U$17945 ( \18322 , \18315 );
not \U$17946 ( \18323 , \18322 );
or \U$17947 ( \18324 , \18321 , \18323 );
not \U$17948 ( \18325 , \18312 );
nand \U$17949 ( \18326 , \18324 , \18325 );
nand \U$17950 ( \18327 , \18319 , \18326 );
not \U$17951 ( \18328 , \18327 );
or \U$17952 ( \18329 , \18286 , \18328 );
not \U$17953 ( \18330 , \18320 );
not \U$17954 ( \18331 , \18322 );
or \U$17955 ( \18332 , \18330 , \18331 );
nand \U$17956 ( \18333 , \18332 , \18312 );
nand \U$17957 ( \18334 , \18329 , \18333 );
not \U$17958 ( \18335 , \18334 );
xor \U$17959 ( \18336 , \18280 , \18335 );
not \U$17960 ( \18337 , \9644 );
not \U$17961 ( \18338 , RIae7a3a8_177);
not \U$17962 ( \18339 , \2287 );
or \U$17963 ( \18340 , \18338 , \18339 );
or \U$17964 ( \18341 , \2287 , RIae7a3a8_177);
nand \U$17965 ( \18342 , \18340 , \18341 );
not \U$17966 ( \18343 , \18342 );
or \U$17967 ( \18344 , \18337 , \18343 );
nand \U$17968 ( \18345 , \18065 , \9621 );
nand \U$17969 ( \18346 , \18344 , \18345 );
not \U$17970 ( \18347 , \9699 );
not \U$17971 ( \18348 , \18208 );
or \U$17972 ( \18349 , \18347 , \18348 );
not \U$17973 ( \18350 , RIae7a240_174);
not \U$17974 ( \18351 , \1758 );
or \U$17975 ( \18352 , \18350 , \18351 );
or \U$17976 ( \18353 , \10608 , RIae7a240_174);
nand \U$17977 ( \18354 , \18352 , \18353 );
nand \U$17978 ( \18355 , \18354 , \9688 );
nand \U$17979 ( \18356 , \18349 , \18355 );
or \U$17980 ( \18357 , \18346 , \18356 );
not \U$17981 ( \18358 , \9527 );
not \U$17982 ( \18359 , \18073 );
or \U$17983 ( \18360 , \18358 , \18359 );
and \U$17984 ( \18361 , RIae7a7e0_186, \1404 );
not \U$17985 ( \18362 , RIae7a7e0_186);
and \U$17986 ( \18363 , \18362 , \3688 );
nor \U$17987 ( \18364 , \18361 , \18363 );
nand \U$17988 ( \18365 , \9549 , \18364 );
nand \U$17989 ( \18366 , \18360 , \18365 );
nand \U$17990 ( \18367 , \18357 , \18366 );
nand \U$17991 ( \18368 , \18346 , \18356 );
nand \U$17992 ( \18369 , \18367 , \18368 );
not \U$17993 ( \18370 , \5048 );
not \U$17994 ( \18371 , \18003 );
or \U$17995 ( \18372 , \18370 , \18371 );
and \U$17996 ( \18373 , RIae79d90_164, \3270 );
not \U$17997 ( \18374 , RIae79d90_164);
and \U$17998 ( \18375 , \18374 , \2404 );
or \U$17999 ( \18376 , \18373 , \18375 );
nand \U$18000 ( \18377 , \18376 , \6091 );
nand \U$18001 ( \18378 , \18372 , \18377 );
not \U$18002 ( \18379 , \18378 );
not \U$18003 ( \18380 , \15382 );
not \U$18004 ( \18381 , RIae7a498_179);
not \U$18005 ( \18382 , \3244 );
or \U$18006 ( \18383 , \18381 , \18382 );
not \U$18007 ( \18384 , \2230 );
not \U$18008 ( \18385 , \18384 );
or \U$18009 ( \18386 , \18385 , RIae7a498_179);
nand \U$18010 ( \18387 , \18383 , \18386 );
not \U$18011 ( \18388 , \18387 );
or \U$18012 ( \18389 , \18380 , \18388 );
nand \U$18013 ( \18390 , \17120 , \12371 );
nand \U$18014 ( \18391 , \18389 , \18390 );
not \U$18015 ( \18392 , \18391 );
or \U$18016 ( \18393 , \18379 , \18392 );
or \U$18017 ( \18394 , \18391 , \18378 );
not \U$18018 ( \18395 , \9473 );
not \U$18019 ( \18396 , RIae7a6f0_184);
not \U$18020 ( \18397 , \5081 );
or \U$18021 ( \18398 , \18396 , \18397 );
or \U$18022 ( \18399 , \1125 , RIae7a6f0_184);
nand \U$18023 ( \18400 , \18398 , \18399 );
not \U$18024 ( \18401 , \18400 );
or \U$18025 ( \18402 , \18395 , \18401 );
nand \U$18026 ( \18403 , \17126 , \9705 );
nand \U$18027 ( \18404 , \18402 , \18403 );
nand \U$18028 ( \18405 , \18394 , \18404 );
nand \U$18029 ( \18406 , \18393 , \18405 );
xor \U$18030 ( \18407 , \18369 , \18406 );
not \U$18031 ( \18408 , RIae7aab0_192);
not \U$18032 ( \18409 , \18051 );
or \U$18033 ( \18410 , \18408 , \18409 );
and \U$18034 ( \18411 , RIae7aa38_191, \938 );
not \U$18035 ( \18412 , RIae7aa38_191);
not \U$18036 ( \18413 , \9770 );
not \U$18037 ( \18414 , \18413 );
and \U$18038 ( \18415 , \18412 , \18414 );
or \U$18039 ( \18416 , \18411 , \18415 );
nand \U$18040 ( \18417 , \18416 , \16383 );
nand \U$18041 ( \18418 , \18410 , \18417 );
not \U$18042 ( \18419 , \18418 );
not \U$18043 ( \18420 , \9792 );
not \U$18044 ( \18421 , \11054 );
not \U$18045 ( \18422 , \18029 );
or \U$18046 ( \18423 , \18421 , \18422 );
or \U$18047 ( \18424 , \10583 , \9804 );
nand \U$18048 ( \18425 , \18423 , \18424 );
not \U$18049 ( \18426 , \18425 );
or \U$18050 ( \18427 , \18420 , \18426 );
nand \U$18051 ( \18428 , \18214 , \9814 );
nand \U$18052 ( \18429 , \18427 , \18428 );
not \U$18053 ( \18430 , \9728 );
and \U$18054 ( \18431 , RIae7a060_170, \17068 );
not \U$18055 ( \18432 , RIae7a060_170);
and \U$18056 ( \18433 , \18432 , \17067 );
nor \U$18057 ( \18434 , \18431 , \18433 );
not \U$18058 ( \18435 , \18434 );
or \U$18059 ( \18436 , \18430 , \18435 );
nand \U$18060 ( \18437 , \18231 , \10542 );
nand \U$18061 ( \18438 , \18436 , \18437 );
xor \U$18062 ( \18439 , \18429 , \18438 );
not \U$18063 ( \18440 , \18439 );
or \U$18064 ( \18441 , \18419 , \18440 );
nand \U$18065 ( \18442 , \18429 , \18438 );
nand \U$18066 ( \18443 , \18441 , \18442 );
and \U$18067 ( \18444 , \18407 , \18443 );
and \U$18068 ( \18445 , \18369 , \18406 );
or \U$18069 ( \18446 , \18444 , \18445 );
xor \U$18070 ( \18447 , \18336 , \18446 );
xor \U$18071 ( \18448 , \18274 , \18269 );
xnor \U$18072 ( \18449 , \18448 , \18263 );
not \U$18073 ( \18450 , \18152 );
not \U$18074 ( \18451 , \18131 );
not \U$18075 ( \18452 , \18136 );
and \U$18076 ( \18453 , \18451 , \18452 );
and \U$18077 ( \18454 , \18131 , \18136 );
nor \U$18078 ( \18455 , \18453 , \18454 );
not \U$18079 ( \18456 , \18455 );
and \U$18080 ( \18457 , \18450 , \18456 );
and \U$18081 ( \18458 , \18152 , \18455 );
nor \U$18082 ( \18459 , \18457 , \18458 );
or \U$18083 ( \18460 , \18449 , \18459 );
not \U$18084 ( \18461 , \9517 );
not \U$18085 ( \18462 , \18040 );
or \U$18086 ( \18463 , \18461 , \18462 );
and \U$18087 ( \18464 , RIae79fe8_169, \2093 );
not \U$18088 ( \18465 , RIae79fe8_169);
and \U$18089 ( \18466 , \18465 , \13008 );
nor \U$18090 ( \18467 , \18464 , \18466 );
nand \U$18091 ( \18468 , \18467 , \11914 );
nand \U$18092 ( \18469 , \18463 , \18468 );
not \U$18093 ( \18470 , \18469 );
not \U$18094 ( \18471 , \6214 );
not \U$18095 ( \18472 , \18014 );
or \U$18096 ( \18473 , \18471 , \18472 );
and \U$18097 ( \18474 , RIae79ef8_167, \3216 );
not \U$18098 ( \18475 , RIae79ef8_167);
and \U$18099 ( \18476 , \18475 , \12996 );
or \U$18100 ( \18477 , \18474 , \18476 );
nand \U$18101 ( \18478 , \18477 , \6201 );
nand \U$18102 ( \18479 , \18473 , \18478 );
not \U$18103 ( \18480 , \18479 );
or \U$18104 ( \18481 , \18470 , \18480 );
or \U$18105 ( \18482 , \18469 , \18479 );
not \U$18106 ( \18483 , \9758 );
not \U$18107 ( \18484 , \10658 );
not \U$18108 ( \18485 , \1898 );
or \U$18109 ( \18486 , \18484 , \18485 );
or \U$18110 ( \18487 , \1898 , \10658 );
nand \U$18111 ( \18488 , \18486 , \18487 );
not \U$18112 ( \18489 , \18488 );
or \U$18113 ( \18490 , \18483 , \18489 );
nand \U$18114 ( \18491 , \18023 , \9777 );
nand \U$18115 ( \18492 , \18490 , \18491 );
nand \U$18116 ( \18493 , \18482 , \18492 );
nand \U$18117 ( \18494 , \18481 , \18493 );
nand \U$18118 ( \18495 , \18460 , \18494 );
nand \U$18119 ( \18496 , \18449 , \18459 );
nand \U$18120 ( \18497 , \18495 , \18496 );
and \U$18121 ( \18498 , \18447 , \18497 );
and \U$18122 ( \18499 , \18336 , \18446 );
or \U$18123 ( \18500 , \18498 , \18499 );
not \U$18124 ( \18501 , \18500 );
nand \U$18125 ( \18502 , \18252 , \18501 );
not \U$18126 ( \18503 , \18502 );
or \U$18127 ( \18504 , \18186 , \18503 );
nand \U$18128 ( \18505 , \18251 , \18500 );
nand \U$18129 ( \18506 , \18504 , \18505 );
not \U$18130 ( \18507 , \18506 );
xor \U$18131 ( \18508 , \16620 , \16741 );
xnor \U$18132 ( \18509 , \18508 , \16743 );
xor \U$18133 ( \18510 , \16491 , \16494 );
xor \U$18134 ( \18511 , \18510 , \16533 );
xor \U$18135 ( \18512 , \18509 , \18511 );
xor \U$18136 ( \18513 , \18163 , \18167 );
and \U$18137 ( \18514 , \18513 , \18171 );
and \U$18138 ( \18515 , \18163 , \18167 );
or \U$18139 ( \18516 , \18514 , \18515 );
and \U$18140 ( \18517 , \16715 , \16725 );
and \U$18141 ( \18518 , \16708 , \16714 );
nor \U$18142 ( \18519 , \18517 , \18518 );
nor \U$18143 ( \18520 , \18516 , \18519 );
not \U$18144 ( \18521 , \18520 );
nand \U$18145 ( \18522 , \18516 , \18519 );
nand \U$18146 ( \18523 , \18521 , \18522 );
not \U$18147 ( \18524 , \18108 );
not \U$18148 ( \18525 , \18125 );
or \U$18149 ( \18526 , \18524 , \18525 );
not \U$18150 ( \18527 , \18115 );
not \U$18151 ( \18528 , \18114 );
or \U$18152 ( \18529 , \18527 , \18528 );
nand \U$18153 ( \18530 , \18529 , \18124 );
nand \U$18154 ( \18531 , \18526 , \18530 );
xor \U$18155 ( \18532 , \18523 , \18531 );
nand \U$18156 ( \18533 , \18334 , \18258 );
not \U$18157 ( \18534 , \18335 );
not \U$18158 ( \18535 , \18258 );
not \U$18159 ( \18536 , \18535 );
or \U$18160 ( \18537 , \18534 , \18536 );
not \U$18161 ( \18538 , \18279 );
nand \U$18162 ( \18539 , \18537 , \18538 );
and \U$18163 ( \18540 , \18533 , \18539 );
and \U$18164 ( \18541 , \18532 , \18540 );
not \U$18165 ( \18542 , \18532 );
nand \U$18166 ( \18543 , \18539 , \18533 );
and \U$18167 ( \18544 , \18542 , \18543 );
nor \U$18168 ( \18545 , \18541 , \18544 );
not \U$18169 ( \18546 , \18172 );
not \U$18170 ( \18547 , \18546 );
not \U$18171 ( \18548 , \18179 );
or \U$18172 ( \18549 , \18547 , \18548 );
not \U$18173 ( \18550 , \18176 );
nand \U$18174 ( \18551 , \18549 , \18550 );
not \U$18175 ( \18552 , \18179 );
nand \U$18176 ( \18553 , \18552 , \18172 );
nand \U$18177 ( \18554 , \18551 , \18553 );
not \U$18178 ( \18555 , \18554 );
and \U$18179 ( \18556 , \18545 , \18555 );
not \U$18180 ( \18557 , \18545 );
and \U$18181 ( \18558 , \18557 , \18554 );
nor \U$18182 ( \18559 , \18556 , \18558 );
nand \U$18183 ( \18560 , \18512 , \18559 );
not \U$18184 ( \18561 , \18555 );
not \U$18185 ( \18562 , \18532 );
not \U$18186 ( \18563 , \18562 );
or \U$18187 ( \18564 , \18561 , \18563 );
not \U$18188 ( \18565 , \18554 );
not \U$18189 ( \18566 , \18532 );
or \U$18190 ( \18567 , \18565 , \18566 );
nand \U$18191 ( \18568 , \18567 , \18543 );
nand \U$18192 ( \18569 , \18564 , \18568 );
not \U$18193 ( \18570 , \18569 );
xor \U$18194 ( \18571 , \17654 , \17656 );
xor \U$18195 ( \18572 , \18571 , \17758 );
not \U$18196 ( \18573 , \18572 );
nand \U$18197 ( \18574 , \18570 , \18573 );
nand \U$18198 ( \18575 , \18572 , \18569 );
nand \U$18199 ( \18576 , \18574 , \18575 );
not \U$18200 ( \18577 , \18193 );
not \U$18201 ( \18578 , \18247 );
or \U$18202 ( \18579 , \18577 , \18578 );
not \U$18203 ( \18580 , \18194 );
not \U$18204 ( \18581 , \18246 );
or \U$18205 ( \18582 , \18580 , \18581 );
buf \U$18206 ( \18583 , \18190 );
nand \U$18207 ( \18584 , \18582 , \18583 );
nand \U$18208 ( \18585 , \18579 , \18584 );
and \U$18209 ( \18586 , \18576 , \18585 );
not \U$18210 ( \18587 , \18576 );
not \U$18211 ( \18588 , \18585 );
and \U$18212 ( \18589 , \18587 , \18588 );
nor \U$18213 ( \18590 , \18586 , \18589 );
nand \U$18214 ( \18591 , \18509 , \18511 );
and \U$18215 ( \18592 , \18560 , \18590 , \18591 );
or \U$18216 ( \18593 , \18507 , \18592 );
not \U$18217 ( \18594 , \18591 );
not \U$18218 ( \18595 , \18560 );
or \U$18219 ( \18596 , \18594 , \18595 );
not \U$18220 ( \18597 , \18590 );
nand \U$18221 ( \18598 , \18596 , \18597 );
nand \U$18222 ( \18599 , \18593 , \18598 );
not \U$18223 ( \18600 , \18574 );
not \U$18224 ( \18601 , \18585 );
or \U$18225 ( \18602 , \18600 , \18601 );
nand \U$18226 ( \18603 , \18602 , \18575 );
not \U$18227 ( \18604 , \18522 );
not \U$18228 ( \18605 , \18531 );
or \U$18229 ( \18606 , \18604 , \18605 );
not \U$18230 ( \18607 , \18520 );
nand \U$18231 ( \18608 , \18606 , \18607 );
not \U$18232 ( \18609 , \9814 );
not \U$18233 ( \18610 , \16127 );
or \U$18234 ( \18611 , \18609 , \18610 );
nand \U$18235 ( \18612 , \18222 , \9792 );
nand \U$18236 ( \18613 , \18611 , \18612 );
not \U$18237 ( \18614 , \18613 );
not \U$18238 ( \18615 , \9499 );
not \U$18239 ( \18616 , \18033 );
or \U$18240 ( \18617 , \18615 , \18616 );
nand \U$18241 ( \18618 , \16116 , \9518 );
nand \U$18242 ( \18619 , \18617 , \18618 );
not \U$18243 ( \18620 , \18619 );
or \U$18244 ( \18621 , \18614 , \18620 );
or \U$18245 ( \18622 , \18613 , \18619 );
not \U$18246 ( \18623 , \9478 );
not \U$18247 ( \18624 , \16106 );
or \U$18248 ( \18625 , \18623 , \18624 );
nand \U$18249 ( \18626 , \17131 , \9473 );
nand \U$18250 ( \18627 , \18625 , \18626 );
nand \U$18251 ( \18628 , \18622 , \18627 );
nand \U$18252 ( \18629 , \18621 , \18628 );
and \U$18253 ( \18630 , \17380 , \17378 );
not \U$18254 ( \18631 , \17380 );
and \U$18255 ( \18632 , \18631 , \17375 );
nor \U$18256 ( \18633 , \18630 , \18632 );
xor \U$18257 ( \18634 , \17393 , \18633 );
nand \U$18258 ( \18635 , \18629 , \18634 );
not \U$18259 ( \18636 , \18635 );
not \U$18260 ( \18637 , \17321 );
not \U$18261 ( \18638 , \17351 );
or \U$18262 ( \18639 , \18637 , \18638 );
or \U$18263 ( \18640 , \17351 , \17321 );
nand \U$18264 ( \18641 , \18639 , \18640 );
buf \U$18265 ( \18642 , \17333 );
not \U$18266 ( \18643 , \18642 );
and \U$18267 ( \18644 , \18641 , \18643 );
not \U$18268 ( \18645 , \18641 );
and \U$18269 ( \18646 , \18645 , \18642 );
nor \U$18270 ( \18647 , \18644 , \18646 );
not \U$18271 ( \18648 , \18647 );
or \U$18272 ( \18649 , \18636 , \18648 );
not \U$18273 ( \18650 , \18629 );
not \U$18274 ( \18651 , \18634 );
nand \U$18275 ( \18652 , \18650 , \18651 );
nand \U$18276 ( \18653 , \18649 , \18652 );
not \U$18277 ( \18654 , \18653 );
xor \U$18278 ( \18655 , \18608 , \18654 );
nor \U$18279 ( \18656 , \17300 , \17263 );
or \U$18280 ( \18657 , \18656 , \17268 );
nand \U$18281 ( \18658 , \17300 , \17263 );
nand \U$18282 ( \18659 , \18657 , \18658 );
and \U$18283 ( \18660 , \18655 , \18659 );
and \U$18284 ( \18661 , \18608 , \18654 );
or \U$18285 ( \18662 , \18660 , \18661 );
xor \U$18286 ( \18663 , \14599 , \14621 );
not \U$18287 ( \18664 , \1072 );
not \U$18288 ( \18665 , \14618 );
or \U$18289 ( \18666 , \18664 , \18665 );
nand \U$18290 ( \18667 , \16181 , \1086 );
nand \U$18291 ( \18668 , \18666 , \18667 );
xor \U$18292 ( \18669 , \16162 , \16174 );
and \U$18293 ( \18670 , \18669 , \16189 );
and \U$18294 ( \18671 , \16162 , \16174 );
or \U$18295 ( \18672 , \18670 , \18671 );
xor \U$18296 ( \18673 , \18668 , \18672 );
not \U$18297 ( \18674 , \1012 );
not \U$18298 ( \18675 , \17573 );
or \U$18299 ( \18676 , \18674 , \18675 );
nand \U$18300 ( \18677 , \16204 , \1008 );
nand \U$18301 ( \18678 , \18676 , \18677 );
and \U$18302 ( \18679 , \18673 , \18678 );
and \U$18303 ( \18680 , \18668 , \18672 );
or \U$18304 ( \18681 , \18679 , \18680 );
xor \U$18305 ( \18682 , \18663 , \18681 );
not \U$18306 ( \18683 , \17412 );
not \U$18307 ( \18684 , \17433 );
or \U$18308 ( \18685 , \18683 , \18684 );
nand \U$18309 ( \18686 , \17421 , \17432 );
nand \U$18310 ( \18687 , \18685 , \18686 );
xnor \U$18311 ( \18688 , \18682 , \18687 );
not \U$18312 ( \18689 , \14768 );
not \U$18313 ( \18690 , \16420 );
or \U$18314 ( \18691 , \18689 , \18690 );
nand \U$18315 ( \18692 , \14767 , \6214 );
nand \U$18316 ( \18693 , \18691 , \18692 );
not \U$18317 ( \18694 , \18693 );
not \U$18318 ( \18695 , \11914 );
not \U$18319 ( \18696 , \16429 );
or \U$18320 ( \18697 , \18695 , \18696 );
nand \U$18321 ( \18698 , \14755 , \9517 );
nand \U$18322 ( \18699 , \18697 , \18698 );
not \U$18323 ( \18700 , \18699 );
xor \U$18324 ( \18701 , \18694 , \18700 );
not \U$18325 ( \18702 , \13158 );
not \U$18326 ( \18703 , \16409 );
or \U$18327 ( \18704 , \18702 , \18703 );
nand \U$18328 ( \18705 , \14782 , \9776 );
nand \U$18329 ( \18706 , \18704 , \18705 );
xor \U$18330 ( \18707 , \18701 , \18706 );
xor \U$18331 ( \18708 , \18688 , \18707 );
xor \U$18332 ( \18709 , \17734 , \17743 );
and \U$18333 ( \18710 , \18709 , \17754 );
and \U$18334 ( \18711 , \17734 , \17743 );
or \U$18335 ( \18712 , \18710 , \18711 );
xor \U$18336 ( \18713 , \18668 , \18672 );
xor \U$18337 ( \18714 , \18713 , \18678 );
or \U$18338 ( \18715 , \18712 , \18714 );
not \U$18339 ( \18716 , \17239 );
not \U$18340 ( \18717 , \17251 );
or \U$18341 ( \18718 , \18716 , \18717 );
nand \U$18342 ( \18719 , \17252 , \17262 );
nand \U$18343 ( \18720 , \18718 , \18719 );
nand \U$18344 ( \18721 , \18715 , \18720 );
nand \U$18345 ( \18722 , \18712 , \18714 );
nand \U$18346 ( \18723 , \18721 , \18722 );
buf \U$18347 ( \18724 , \18723 );
xnor \U$18348 ( \18725 , \18708 , \18724 );
xor \U$18349 ( \18726 , \18662 , \18725 );
not \U$18350 ( \18727 , \17354 );
not \U$18351 ( \18728 , \17438 );
or \U$18352 ( \18729 , \18727 , \18728 );
or \U$18353 ( \18730 , \17354 , \17438 );
nand \U$18354 ( \18731 , \18729 , \18730 );
not \U$18355 ( \18732 , \18731 );
xor \U$18356 ( \18733 , \18714 , \18720 );
xnor \U$18357 ( \18734 , \18733 , \18712 );
not \U$18358 ( \18735 , \18734 );
not \U$18359 ( \18736 , \18735 );
or \U$18360 ( \18737 , \18732 , \18736 );
not \U$18361 ( \18738 , \18734 );
not \U$18362 ( \18739 , \18731 );
not \U$18363 ( \18740 , \18739 );
or \U$18364 ( \18741 , \18738 , \18740 );
xor \U$18365 ( \18742 , \16191 , \16206 );
not \U$18366 ( \18743 , \18742 );
xor \U$18367 ( \18744 , \17224 , \17235 );
not \U$18368 ( \18745 , \10275 );
not \U$18369 ( \18746 , \16593 );
or \U$18370 ( \18747 , \18745 , \18746 );
nand \U$18371 ( \18748 , \18090 , \11205 );
nand \U$18372 ( \18749 , \18747 , \18748 );
not \U$18373 ( \18750 , \18749 );
and \U$18374 ( \18751 , \18744 , \18750 );
not \U$18375 ( \18752 , \18744 );
not \U$18376 ( \18753 , \10275 );
not \U$18377 ( \18754 , \16593 );
or \U$18378 ( \18755 , \18753 , \18754 );
nand \U$18379 ( \18756 , \18755 , \18748 );
and \U$18380 ( \18757 , \18752 , \18756 );
or \U$18381 ( \18758 , \18751 , \18757 );
not \U$18382 ( \18759 , \10631 );
not \U$18383 ( \18760 , \17329 );
or \U$18384 ( \18761 , \18759 , \18760 );
nand \U$18385 ( \18762 , \18150 , \11400 );
nand \U$18386 ( \18763 , \18761 , \18762 );
and \U$18387 ( \18764 , \18758 , \18763 );
and \U$18388 ( \18765 , \18749 , \18744 );
nor \U$18389 ( \18766 , \18764 , \18765 );
nand \U$18390 ( \18767 , \18743 , \18766 );
not \U$18391 ( \18768 , \18767 );
not \U$18392 ( \18769 , \17094 );
and \U$18393 ( \18770 , \17104 , \17116 );
not \U$18394 ( \18771 , \17104 );
and \U$18395 ( \18772 , \18771 , \17117 );
nor \U$18396 ( \18773 , \18770 , \18772 );
not \U$18397 ( \18774 , \18773 );
or \U$18398 ( \18775 , \18769 , \18774 );
nand \U$18399 ( \18776 , \17116 , \17104 );
nand \U$18400 ( \18777 , \18775 , \18776 );
not \U$18401 ( \18778 , \18777 );
or \U$18402 ( \18779 , \18768 , \18778 );
not \U$18403 ( \18780 , \18766 );
nand \U$18404 ( \18781 , \18780 , \18742 );
nand \U$18405 ( \18782 , \18779 , \18781 );
nand \U$18406 ( \18783 , \18741 , \18782 );
nand \U$18407 ( \18784 , \18737 , \18783 );
xor \U$18408 ( \18785 , \18726 , \18784 );
xor \U$18409 ( \18786 , \18603 , \18785 );
xor \U$18410 ( \18787 , \18608 , \18654 );
xor \U$18411 ( \18788 , \18787 , \18659 );
not \U$18412 ( \18789 , \18788 );
not \U$18413 ( \18790 , \18735 );
not \U$18414 ( \18791 , \18739 );
or \U$18415 ( \18792 , \18790 , \18791 );
nand \U$18416 ( \18793 , \18734 , \18731 );
nand \U$18417 ( \18794 , \18792 , \18793 );
not \U$18418 ( \18795 , \18782 );
and \U$18419 ( \18796 , \18794 , \18795 );
not \U$18420 ( \18797 , \18794 );
and \U$18421 ( \18798 , \18797 , \18782 );
nor \U$18422 ( \18799 , \18796 , \18798 );
nand \U$18423 ( \18800 , \18789 , \18799 );
not \U$18424 ( \18801 , \18800 );
xor \U$18425 ( \18802 , \18742 , \18766 );
xnor \U$18426 ( \18803 , \18802 , \18777 );
not \U$18427 ( \18804 , \18803 );
buf \U$18428 ( \18805 , \18629 );
xor \U$18429 ( \18806 , \18634 , \18805 );
xnor \U$18430 ( \18807 , \18806 , \18647 );
xor \U$18431 ( \18808 , \18613 , \18619 );
xnor \U$18432 ( \18809 , \18808 , \18627 );
not \U$18433 ( \18810 , \18809 );
and \U$18434 ( \18811 , \18758 , \18763 );
not \U$18435 ( \18812 , \18758 );
not \U$18436 ( \18813 , \18763 );
and \U$18437 ( \18814 , \18812 , \18813 );
nor \U$18438 ( \18815 , \18811 , \18814 );
not \U$18439 ( \18816 , \18815 );
not \U$18440 ( \18817 , \18816 );
or \U$18441 ( \18818 , \18810 , \18817 );
xor \U$18442 ( \18819 , \17287 , \17278 );
xor \U$18443 ( \18820 , \18819 , \17297 );
nand \U$18444 ( \18821 , \18818 , \18820 );
not \U$18445 ( \18822 , \18809 );
nand \U$18446 ( \18823 , \18822 , \18815 );
nand \U$18447 ( \18824 , \18821 , \18823 );
and \U$18448 ( \18825 , \18807 , \18824 );
not \U$18449 ( \18826 , \18807 );
not \U$18450 ( \18827 , \18824 );
and \U$18451 ( \18828 , \18826 , \18827 );
nor \U$18452 ( \18829 , \18825 , \18828 );
not \U$18453 ( \18830 , \18829 );
or \U$18454 ( \18831 , \18804 , \18830 );
nand \U$18455 ( \18832 , \18807 , \18824 );
nand \U$18456 ( \18833 , \18831 , \18832 );
not \U$18457 ( \18834 , \18833 );
or \U$18458 ( \18835 , \18801 , \18834 );
not \U$18459 ( \18836 , \18799 );
nand \U$18460 ( \18837 , \18836 , \18788 );
nand \U$18461 ( \18838 , \18835 , \18837 );
xor \U$18462 ( \18839 , \18786 , \18838 );
xor \U$18463 ( \18840 , \18599 , \18839 );
xnor \U$18464 ( \18841 , \18788 , \18799 );
xor \U$18465 ( \18842 , \18833 , \18841 );
xor \U$18466 ( \18843 , \16489 , \16746 );
xor \U$18467 ( \18844 , \18843 , \17308 );
xor \U$18468 ( \18845 , \18842 , \18844 );
buf \U$18469 ( \18846 , \17047 );
not \U$18470 ( \18847 , \17306 );
not \U$18471 ( \18848 , \17305 );
or \U$18472 ( \18849 , \18847 , \18848 );
or \U$18473 ( \18850 , \17305 , \17306 );
nand \U$18474 ( \18851 , \18849 , \18850 );
xor \U$18475 ( \18852 , \18846 , \18851 );
xnor \U$18476 ( \18853 , \18829 , \18803 );
not \U$18477 ( \18854 , \18853 );
not \U$18478 ( \18855 , \18816 );
not \U$18479 ( \18856 , \18822 );
or \U$18480 ( \18857 , \18855 , \18856 );
nand \U$18481 ( \18858 , \18815 , \18809 );
nand \U$18482 ( \18859 , \18857 , \18858 );
and \U$18483 ( \18860 , \18859 , \18820 );
not \U$18484 ( \18861 , \18859 );
not \U$18485 ( \18862 , \18820 );
and \U$18486 ( \18863 , \18861 , \18862 );
nor \U$18487 ( \18864 , \18860 , \18863 );
not \U$18488 ( \18865 , \18235 );
not \U$18489 ( \18866 , \18244 );
or \U$18490 ( \18867 , \18865 , \18866 );
or \U$18491 ( \18868 , \18244 , \18235 );
nand \U$18492 ( \18869 , \18867 , \18868 );
and \U$18493 ( \18870 , \18869 , \18240 );
not \U$18494 ( \18871 , \18869 );
nand \U$18495 ( \18872 , \18239 , \18238 );
and \U$18496 ( \18873 , \18871 , \18872 );
or \U$18497 ( \18874 , \18870 , \18873 );
xor \U$18498 ( \18875 , \18864 , \18874 );
not \U$18499 ( \18876 , \10631 );
not \U$18500 ( \18877 , \18144 );
or \U$18501 ( \18878 , \18876 , \18877 );
not \U$18502 ( \18879 , RIae7a510_180);
not \U$18503 ( \18880 , \2954 );
or \U$18504 ( \18881 , \18879 , \18880 );
or \U$18505 ( \18882 , \2954 , RIae7a510_180);
nand \U$18506 ( \18883 , \18881 , \18882 );
nand \U$18507 ( \18884 , \18883 , \10927 );
nand \U$18508 ( \18885 , \18878 , \18884 );
not \U$18509 ( \18886 , \18885 );
xor \U$18510 ( \18887 , \18307 , \18301 );
not \U$18511 ( \18888 , \10275 );
not \U$18512 ( \18889 , \18082 );
or \U$18513 ( \18890 , \18888 , \18889 );
not \U$18514 ( \18891 , \18088 );
not \U$18515 ( \18892 , \883 );
or \U$18516 ( \18893 , \18891 , \18892 );
nand \U$18517 ( \18894 , \877 , RIae7a8d0_188);
nand \U$18518 ( \18895 , \18893 , \18894 );
nand \U$18519 ( \18896 , \18895 , \16594 );
nand \U$18520 ( \18897 , \18890 , \18896 );
xor \U$18521 ( \18898 , \18887 , \18897 );
not \U$18522 ( \18899 , \18898 );
or \U$18523 ( \18900 , \18886 , \18899 );
nand \U$18524 ( \18901 , \18897 , \18887 );
nand \U$18525 ( \18902 , \18900 , \18901 );
not \U$18526 ( \18903 , \18902 );
xor \U$18527 ( \18904 , \17192 , \17133 );
xnor \U$18528 ( \18905 , \18904 , \17124 );
not \U$18529 ( \18906 , \18285 );
not \U$18530 ( \18907 , \18906 );
not \U$18531 ( \18908 , \18327 );
and \U$18532 ( \18909 , \18907 , \18908 );
and \U$18533 ( \18910 , \18327 , \18906 );
nor \U$18534 ( \18911 , \18909 , \18910 );
and \U$18535 ( \18912 , \18905 , \18911 );
not \U$18536 ( \18913 , \18905 );
not \U$18537 ( \18914 , \18911 );
and \U$18538 ( \18915 , \18913 , \18914 );
or \U$18539 ( \18916 , \18912 , \18915 );
not \U$18540 ( \18917 , \18916 );
or \U$18541 ( \18918 , \18903 , \18917 );
nand \U$18542 ( \18919 , \18905 , \18914 );
nand \U$18543 ( \18920 , \18918 , \18919 );
and \U$18544 ( \18921 , \18875 , \18920 );
and \U$18545 ( \18922 , \18864 , \18874 );
or \U$18546 ( \18923 , \18921 , \18922 );
nand \U$18547 ( \18924 , \18854 , \18923 );
and \U$18548 ( \18925 , \18852 , \18924 );
not \U$18549 ( \18926 , \18923 );
and \U$18550 ( \18927 , \18926 , \18853 );
nor \U$18551 ( \18928 , \18925 , \18927 );
and \U$18552 ( \18929 , \18845 , \18928 );
and \U$18553 ( \18930 , \18842 , \18844 );
or \U$18554 ( \18931 , \18929 , \18930 );
xor \U$18555 ( \18932 , \18840 , \18931 );
xor \U$18556 ( \18933 , \17950 , \18932 );
not \U$18557 ( \18934 , \18592 );
nand \U$18558 ( \18935 , \18934 , \18598 );
and \U$18559 ( \18936 , \18935 , \18506 );
not \U$18560 ( \18937 , \18935 );
and \U$18561 ( \18938 , \18937 , \18507 );
nor \U$18562 ( \18939 , \18936 , \18938 );
not \U$18563 ( \18940 , \18939 );
not \U$18564 ( \18941 , \18940 );
not \U$18565 ( \18942 , \18391 );
xnor \U$18566 ( \18943 , \18404 , \18378 );
not \U$18567 ( \18944 , \18943 );
or \U$18568 ( \18945 , \18942 , \18944 );
or \U$18569 ( \18946 , \18943 , \18391 );
nand \U$18570 ( \18947 , \18945 , \18946 );
not \U$18571 ( \18948 , \18947 );
not \U$18572 ( \18949 , \1820 );
not \U$18573 ( \18950 , RIae79688_149);
not \U$18574 ( \18951 , \11562 );
or \U$18575 ( \18952 , \18950 , \18951 );
or \U$18576 ( \18953 , \10067 , RIae79688_149);
nand \U$18577 ( \18954 , \18952 , \18953 );
not \U$18578 ( \18955 , \18954 );
or \U$18579 ( \18956 , \18949 , \18955 );
xor \U$18580 ( \18957 , \11272 , RIae79688_149);
nand \U$18581 ( \18958 , \18957 , \9320 );
nand \U$18582 ( \18959 , \18956 , \18958 );
not \U$18583 ( \18960 , \18959 );
not \U$18584 ( \18961 , \1012 );
not \U$18585 ( \18962 , \997 );
not \U$18586 ( \18963 , \10272 );
or \U$18587 ( \18964 , \18962 , \18963 );
or \U$18588 ( \18965 , \11321 , \6414 );
nand \U$18589 ( \18966 , \18964 , \18965 );
not \U$18590 ( \18967 , \18966 );
or \U$18591 ( \18968 , \18961 , \18967 );
and \U$18592 ( \18969 , \997 , \10259 );
not \U$18593 ( \18970 , \997 );
not \U$18594 ( \18971 , \10259 );
and \U$18595 ( \18972 , \18970 , \18971 );
nor \U$18596 ( \18973 , \18969 , \18972 );
nand \U$18597 ( \18974 , \18973 , \1007 );
nand \U$18598 ( \18975 , \18968 , \18974 );
not \U$18599 ( \18976 , \18975 );
and \U$18600 ( \18977 , \12857 , \838 );
not \U$18601 ( \18978 , \1049 );
and \U$18602 ( \18979 , RIae79070_136, \10844 );
not \U$18603 ( \18980 , RIae79070_136);
and \U$18604 ( \18981 , \18980 , \16164 );
or \U$18605 ( \18982 , \18979 , \18981 );
not \U$18606 ( \18983 , \18982 );
or \U$18607 ( \18984 , \18978 , \18983 );
not \U$18608 ( \18985 , \16005 );
not \U$18609 ( \18986 , \18985 );
and \U$18610 ( \18987 , \1039 , \18986 );
not \U$18611 ( \18988 , \1039 );
not \U$18612 ( \18989 , \16005 );
and \U$18613 ( \18990 , \18988 , \18989 );
nor \U$18614 ( \18991 , \18987 , \18990 );
nand \U$18615 ( \18992 , \18991 , \1061 );
nand \U$18616 ( \18993 , \18984 , \18992 );
xor \U$18617 ( \18994 , \18977 , \18993 );
not \U$18618 ( \18995 , \18994 );
or \U$18619 ( \18996 , \18976 , \18995 );
nand \U$18620 ( \18997 , \18993 , \18977 );
nand \U$18621 ( \18998 , \18996 , \18997 );
not \U$18622 ( \18999 , \1501 );
not \U$18623 ( \19000 , \16924 );
or \U$18624 ( \19001 , \18999 , \19000 );
not \U$18625 ( \19002 , \1503 );
not \U$18626 ( \19003 , \10042 );
or \U$18627 ( \19004 , \19002 , \19003 );
or \U$18628 ( \19005 , \10042 , \1503 );
nand \U$18629 ( \19006 , \19004 , \19005 );
nand \U$18630 ( \19007 , \19006 , \9403 );
nand \U$18631 ( \19008 , \19001 , \19007 );
xor \U$18632 ( \19009 , \18998 , \19008 );
not \U$18633 ( \19010 , \19009 );
or \U$18634 ( \19011 , \18960 , \19010 );
nand \U$18635 ( \19012 , \19008 , \18998 );
nand \U$18636 ( \19013 , \19011 , \19012 );
not \U$18637 ( \19014 , \2251 );
not \U$18638 ( \19015 , \12644 );
and \U$18639 ( \19016 , RIae79ac0_158, \19015 );
not \U$18640 ( \19017 , RIae79ac0_158);
and \U$18641 ( \19018 , \19017 , \10728 );
or \U$18642 ( \19019 , \19016 , \19018 );
not \U$18643 ( \19020 , \19019 );
or \U$18644 ( \19021 , \19014 , \19020 );
not \U$18645 ( \19022 , RIae79ac0_158);
not \U$18646 ( \19023 , \10084 );
or \U$18647 ( \19024 , \19022 , \19023 );
not \U$18648 ( \19025 , \10084 );
nand \U$18649 ( \19026 , \19025 , \2268 );
nand \U$18650 ( \19027 , \19024 , \19026 );
nand \U$18651 ( \19028 , \19027 , \2272 );
nand \U$18652 ( \19029 , \19021 , \19028 );
not \U$18653 ( \19030 , \19029 );
not \U$18654 ( \19031 , \1863 );
not \U$18655 ( \19032 , RIae793b8_143);
not \U$18656 ( \19033 , \16193 );
or \U$18657 ( \19034 , \19032 , \19033 );
buf \U$18658 ( \19035 , \9989 );
or \U$18659 ( \19036 , \19035 , RIae793b8_143);
nand \U$18660 ( \19037 , \19034 , \19036 );
not \U$18661 ( \19038 , \19037 );
or \U$18662 ( \19039 , \19031 , \19038 );
xnor \U$18663 ( \19040 , \10149 , RIae793b8_143);
nand \U$18664 ( \19041 , \19040 , \1910 );
nand \U$18665 ( \19042 , \19039 , \19041 );
not \U$18666 ( \19043 , \2011 );
not \U$18667 ( \19044 , RIae79610_148);
not \U$18668 ( \19045 , \10749 );
or \U$18669 ( \19046 , \19044 , \19045 );
or \U$18670 ( \19047 , \10749 , RIae79610_148);
nand \U$18671 ( \19048 , \19046 , \19047 );
not \U$18672 ( \19049 , \19048 );
or \U$18673 ( \19050 , \19043 , \19049 );
not \U$18674 ( \19051 , RIae79610_148);
not \U$18675 ( \19052 , \11260 );
or \U$18676 ( \19053 , \19051 , \19052 );
or \U$18677 ( \19054 , \16719 , RIae79610_148);
nand \U$18678 ( \19055 , \19053 , \19054 );
nand \U$18679 ( \19056 , \19055 , \2063 );
nand \U$18680 ( \19057 , \19050 , \19056 );
xor \U$18681 ( \19058 , \19042 , \19057 );
not \U$18682 ( \19059 , \19058 );
or \U$18683 ( \19060 , \19030 , \19059 );
nand \U$18684 ( \19061 , \19057 , \19042 );
nand \U$18685 ( \19062 , \19060 , \19061 );
xor \U$18686 ( \19063 , \19013 , \19062 );
not \U$18687 ( \19064 , \19063 );
not \U$18688 ( \19065 , \9473 );
xor \U$18689 ( \19066 , \3538 , RIae7a6f0_184);
not \U$18690 ( \19067 , \19066 );
or \U$18691 ( \19068 , \19065 , \19067 );
nand \U$18692 ( \19069 , \18400 , \9705 );
nand \U$18693 ( \19070 , \19068 , \19069 );
not \U$18694 ( \19071 , \19070 );
or \U$18695 ( \19072 , \19064 , \19071 );
nand \U$18696 ( \19073 , \19062 , \19013 );
nand \U$18697 ( \19074 , \19072 , \19073 );
not \U$18698 ( \19075 , \19074 );
not \U$18699 ( \19076 , \18885 );
and \U$18700 ( \19077 , \18898 , \19076 );
not \U$18701 ( \19078 , \18898 );
and \U$18702 ( \19079 , \19078 , \18885 );
nor \U$18703 ( \19080 , \19077 , \19079 );
not \U$18704 ( \19081 , \19080 );
or \U$18705 ( \19082 , \19075 , \19081 );
or \U$18706 ( \19083 , \19080 , \19074 );
nand \U$18707 ( \19084 , \19082 , \19083 );
not \U$18708 ( \19085 , \19084 );
or \U$18709 ( \19086 , \18948 , \19085 );
not \U$18710 ( \19087 , \19080 );
nand \U$18711 ( \19088 , \19087 , \19074 );
nand \U$18712 ( \19089 , \19086 , \19088 );
not \U$18713 ( \19090 , \19089 );
xor \U$18714 ( \19091 , \18459 , \18449 );
xnor \U$18715 ( \19092 , \19091 , \18494 );
not \U$18716 ( \19093 , \19092 );
xor \U$18717 ( \19094 , \18369 , \18406 );
xor \U$18718 ( \19095 , \19094 , \18443 );
not \U$18719 ( \19096 , \19095 );
or \U$18720 ( \19097 , \19093 , \19096 );
or \U$18721 ( \19098 , \19095 , \19092 );
nand \U$18722 ( \19099 , \19097 , \19098 );
not \U$18723 ( \19100 , \19099 );
or \U$18724 ( \19101 , \19090 , \19100 );
not \U$18725 ( \19102 , \19092 );
nand \U$18726 ( \19103 , \19102 , \19095 );
nand \U$18727 ( \19104 , \19101 , \19103 );
not \U$18728 ( \19105 , \19104 );
xor \U$18729 ( \19106 , \18346 , \18356 );
buf \U$18730 ( \19107 , \18366 );
xor \U$18731 ( \19108 , \19106 , \19107 );
not \U$18732 ( \19109 , \19108 );
not \U$18733 ( \19110 , \12515 );
not \U$18734 ( \19111 , RIae7a3a8_177);
not \U$18735 ( \19112 , \4024 );
or \U$18736 ( \19113 , \19111 , \19112 );
or \U$18737 ( \19114 , \1741 , RIae7a3a8_177);
nand \U$18738 ( \19115 , \19113 , \19114 );
not \U$18739 ( \19116 , \19115 );
or \U$18740 ( \19117 , \19110 , \19116 );
nand \U$18741 ( \19118 , \18342 , \9622 );
nand \U$18742 ( \19119 , \19117 , \19118 );
not \U$18743 ( \19120 , \19119 );
not \U$18744 ( \19121 , \12233 );
not \U$18745 ( \19122 , \18883 );
or \U$18746 ( \19123 , \19121 , \19122 );
not \U$18747 ( \19124 , \17324 );
not \U$18748 ( \19125 , \2309 );
or \U$18749 ( \19126 , \19124 , \19125 );
not \U$18750 ( \19127 , \14931 );
nand \U$18751 ( \19128 , \19127 , \2305 );
nand \U$18752 ( \19129 , \19126 , \19128 );
nand \U$18753 ( \19130 , \19129 , \10638 );
nand \U$18754 ( \19131 , \19123 , \19130 );
not \U$18755 ( \19132 , \19131 );
not \U$18756 ( \19133 , \9527 );
not \U$18757 ( \19134 , \18364 );
or \U$18758 ( \19135 , \19133 , \19134 );
not \U$18759 ( \19136 , RIae7a7e0_186);
not \U$18760 ( \19137 , \12183 );
or \U$18761 ( \19138 , \19136 , \19137 );
or \U$18762 ( \19139 , \5134 , RIae7a7e0_186);
nand \U$18763 ( \19140 , \19138 , \19139 );
nand \U$18764 ( \19141 , \19140 , \10510 );
nand \U$18765 ( \19142 , \19135 , \19141 );
not \U$18766 ( \19143 , \19142 );
not \U$18767 ( \19144 , \19143 );
or \U$18768 ( \19145 , \19132 , \19144 );
not \U$18769 ( \19146 , \19131 );
nand \U$18770 ( \19147 , \19146 , \19142 );
nand \U$18771 ( \19148 , \19145 , \19147 );
not \U$18772 ( \19149 , \19148 );
or \U$18773 ( \19150 , \19120 , \19149 );
nand \U$18774 ( \19151 , \19142 , \19131 );
nand \U$18775 ( \19152 , \19150 , \19151 );
not \U$18776 ( \19153 , \19152 );
xor \U$18777 ( \19154 , \17005 , \17027 );
xor \U$18778 ( \19155 , \19154 , \17023 );
not \U$18779 ( \19156 , \19155 );
or \U$18780 ( \19157 , \19153 , \19156 );
or \U$18781 ( \19158 , \19152 , \19155 );
nand \U$18782 ( \19159 , \19157 , \19158 );
not \U$18783 ( \19160 , \19159 );
or \U$18784 ( \19161 , \19109 , \19160 );
not \U$18785 ( \19162 , \19155 );
nand \U$18786 ( \19163 , \19162 , \19152 );
nand \U$18787 ( \19164 , \19161 , \19163 );
not \U$18788 ( \19165 , \19164 );
xor \U$18789 ( \19166 , \16973 , \16936 );
xnor \U$18790 ( \19167 , \19166 , \17037 );
not \U$18791 ( \19168 , \19167 );
not \U$18792 ( \19169 , \19168 );
xor \U$18793 ( \19170 , \18916 , \18902 );
not \U$18794 ( \19171 , \19170 );
or \U$18795 ( \19172 , \19169 , \19171 );
or \U$18796 ( \19173 , \19168 , \19170 );
nand \U$18797 ( \19174 , \19172 , \19173 );
not \U$18798 ( \19175 , \19174 );
or \U$18799 ( \19176 , \19165 , \19175 );
nand \U$18800 ( \19177 , \19170 , \19167 );
nand \U$18801 ( \19178 , \19176 , \19177 );
not \U$18802 ( \19179 , \19178 );
xor \U$18803 ( \19180 , \17041 , \16860 );
xor \U$18804 ( \19181 , \19180 , \17045 );
not \U$18805 ( \19182 , \19181 );
and \U$18806 ( \19183 , \19179 , \19182 );
not \U$18807 ( \19184 , \19179 );
and \U$18808 ( \19185 , \19184 , \19181 );
nor \U$18809 ( \19186 , \19183 , \19185 );
not \U$18810 ( \19187 , \19186 );
or \U$18811 ( \19188 , \19105 , \19187 );
nand \U$18812 ( \19189 , \19178 , \19181 );
nand \U$18813 ( \19190 , \19188 , \19189 );
not \U$18814 ( \19191 , \19190 );
xor \U$18815 ( \19192 , \18511 , \18559 );
xnor \U$18816 ( \19193 , \19192 , \18509 );
xor \U$18817 ( \19194 , \18212 , \18224 );
xor \U$18818 ( \19195 , \19194 , \18233 );
xor \U$18819 ( \19196 , \17173 , \17159 );
not \U$18820 ( \19197 , \1843 );
not \U$18821 ( \19198 , \18954 );
or \U$18822 ( \19199 , \19197 , \19198 );
nand \U$18823 ( \19200 , \16945 , \1820 );
nand \U$18824 ( \19201 , \19199 , \19200 );
xor \U$18825 ( \19202 , \19196 , \19201 );
not \U$18826 ( \19203 , \2272 );
not \U$18827 ( \19204 , \19019 );
or \U$18828 ( \19205 , \19203 , \19204 );
nand \U$18829 ( \19206 , \16760 , \2249 );
nand \U$18830 ( \19207 , \19205 , \19206 );
and \U$18831 ( \19208 , \19202 , \19207 );
and \U$18832 ( \19209 , \19196 , \19201 );
nor \U$18833 ( \19210 , \19208 , \19209 );
not \U$18834 ( \19211 , \19210 );
not \U$18835 ( \19212 , \19211 );
xnor \U$18836 ( \19213 , \17178 , \17189 );
not \U$18837 ( \19214 , \19213 );
not \U$18838 ( \19215 , \2431 );
xor \U$18839 ( \19216 , RIae79778_151, \9298 );
not \U$18840 ( \19217 , \19216 );
or \U$18841 ( \19218 , \19215 , \19217 );
nand \U$18842 ( \19219 , \16880 , \2450 );
nand \U$18843 ( \19220 , \19218 , \19219 );
not \U$18844 ( \19221 , \19220 );
not \U$18845 ( \19222 , \2063 );
not \U$18846 ( \19223 , \19048 );
or \U$18847 ( \19224 , \19222 , \19223 );
nand \U$18848 ( \19225 , \17187 , \2011 );
nand \U$18849 ( \19226 , \19224 , \19225 );
not \U$18850 ( \19227 , \19226 );
not \U$18851 ( \19228 , \1910 );
not \U$18852 ( \19229 , \19037 );
or \U$18853 ( \19230 , \19228 , \19229 );
nand \U$18854 ( \19231 , \16955 , \1863 );
nand \U$18855 ( \19232 , \19230 , \19231 );
not \U$18856 ( \19233 , \19232 );
nand \U$18857 ( \19234 , \19227 , \19233 );
not \U$18858 ( \19235 , \19234 );
or \U$18859 ( \19236 , \19221 , \19235 );
nand \U$18860 ( \19237 , \19226 , \19232 );
nand \U$18861 ( \19238 , \19236 , \19237 );
not \U$18862 ( \19239 , \19238 );
or \U$18863 ( \19240 , \19214 , \19239 );
or \U$18864 ( \19241 , \19238 , \19213 );
nand \U$18865 ( \19242 , \19240 , \19241 );
not \U$18866 ( \19243 , \19242 );
or \U$18867 ( \19244 , \19212 , \19243 );
not \U$18868 ( \19245 , \19213 );
nand \U$18869 ( \19246 , \19245 , \19238 );
nand \U$18870 ( \19247 , \19244 , \19246 );
xor \U$18871 ( \19248 , \19195 , \19247 );
not \U$18872 ( \19249 , \2322 );
not \U$18873 ( \19250 , \16987 );
or \U$18874 ( \19251 , \19249 , \19250 );
not \U$18875 ( \19252 , \5344 );
not \U$18876 ( \19253 , \14110 );
or \U$18877 ( \19254 , \19252 , \19253 );
not \U$18878 ( \19255 , RIae798e0_154);
or \U$18879 ( \19256 , \9438 , \19255 );
nand \U$18880 ( \19257 , \19254 , \19256 );
nand \U$18881 ( \19258 , \19257 , \14580 );
nand \U$18882 ( \19259 , \19251 , \19258 );
not \U$18883 ( \19260 , \19259 );
not \U$18884 ( \19261 , \1062 );
not \U$18885 ( \19262 , \18982 );
or \U$18886 ( \19263 , \19261 , \19262 );
nand \U$18887 ( \19264 , \17157 , \1049 );
nand \U$18888 ( \19265 , \19263 , \19264 );
not \U$18889 ( \19266 , \16896 );
not \U$18890 ( \19267 , \16900 );
and \U$18891 ( \19268 , \19266 , \19267 );
and \U$18892 ( \19269 , \16896 , \16900 );
nor \U$18893 ( \19270 , \19268 , \19269 );
xor \U$18894 ( \19271 , \19265 , \19270 );
not \U$18895 ( \19272 , \19271 );
not \U$18896 ( \19273 , \1012 );
not \U$18897 ( \19274 , \16906 );
or \U$18898 ( \19275 , \19273 , \19274 );
nand \U$18899 ( \19276 , \18966 , \1007 );
nand \U$18900 ( \19277 , \19275 , \19276 );
and \U$18901 ( \19278 , \19272 , \19277 );
not \U$18902 ( \19279 , \19270 );
and \U$18903 ( \19280 , \19265 , \19279 );
nor \U$18904 ( \19281 , \19278 , \19280 );
not \U$18905 ( \19282 , \1988 );
and \U$18906 ( \19283 , \12707 , \1991 );
not \U$18907 ( \19284 , \12707 );
and \U$18908 ( \19285 , \19284 , RIae797f0_152);
nor \U$18909 ( \19286 , \19283 , \19285 );
not \U$18910 ( \19287 , \19286 );
or \U$18911 ( \19288 , \19282 , \19287 );
nand \U$18912 ( \19289 , \17002 , \2519 );
nand \U$18913 ( \19290 , \19288 , \19289 );
xnor \U$18914 ( \19291 , \19281 , \19290 );
not \U$18915 ( \19292 , \19291 );
or \U$18916 ( \19293 , \19260 , \19292 );
not \U$18917 ( \19294 , \19281 );
nand \U$18918 ( \19295 , \19294 , \19290 );
nand \U$18919 ( \19296 , \19293 , \19295 );
not \U$18920 ( \19297 , \19296 );
xnor \U$18921 ( \19298 , \16968 , \16947 );
not \U$18922 ( \19299 , \19298 );
not \U$18923 ( \19300 , \2163 );
not \U$18924 ( \19301 , \16774 );
or \U$18925 ( \19302 , \19300 , \19301 );
not \U$18926 ( \19303 , RIae79520_146);
not \U$18927 ( \19304 , \10453 );
or \U$18928 ( \19305 , \19303 , \19304 );
not \U$18929 ( \19306 , \16752 );
or \U$18930 ( \19307 , \19306 , RIae79520_146);
nand \U$18931 ( \19308 , \19305 , \19307 );
nand \U$18932 ( \19309 , \19308 , \12680 );
nand \U$18933 ( \19310 , \19302 , \19309 );
not \U$18934 ( \19311 , RIae79c28_161);
not \U$18935 ( \19312 , \13976 );
or \U$18936 ( \19313 , \19311 , \19312 );
or \U$18937 ( \19314 , \15207 , RIae79c28_161);
nand \U$18938 ( \19315 , \19313 , \19314 );
not \U$18939 ( \19316 , \19315 );
not \U$18940 ( \19317 , \2767 );
or \U$18941 ( \19318 , \19316 , \19317 );
or \U$18942 ( \19319 , \17020 , \5323 );
nand \U$18943 ( \19320 , \19318 , \19319 );
xor \U$18944 ( \19321 , \19310 , \19320 );
not \U$18945 ( \19322 , \5049 );
not \U$18946 ( \19323 , \18376 );
or \U$18947 ( \19324 , \19322 , \19323 );
not \U$18948 ( \19325 , \4982 );
and \U$18949 ( \19326 , RIae79d90_164, \19325 );
not \U$18950 ( \19327 , RIae79d90_164);
and \U$18951 ( \19328 , \19327 , \3208 );
nor \U$18952 ( \19329 , \19326 , \19328 );
not \U$18953 ( \19330 , \6091 );
or \U$18954 ( \19331 , \19329 , \19330 );
nand \U$18955 ( \19332 , \19324 , \19331 );
and \U$18956 ( \19333 , \19321 , \19332 );
and \U$18957 ( \19334 , \19310 , \19320 );
or \U$18958 ( \19335 , \19333 , \19334 );
not \U$18959 ( \19336 , \19335 );
or \U$18960 ( \19337 , \19299 , \19336 );
or \U$18961 ( \19338 , \19335 , \19298 );
nand \U$18962 ( \19339 , \19337 , \19338 );
not \U$18963 ( \19340 , \19339 );
or \U$18964 ( \19341 , \19297 , \19340 );
not \U$18965 ( \19342 , \19298 );
nand \U$18966 ( \19343 , \19342 , \19335 );
nand \U$18967 ( \19344 , \19341 , \19343 );
and \U$18968 ( \19345 , \19248 , \19344 );
and \U$18969 ( \19346 , \19195 , \19247 );
or \U$18970 ( \19347 , \19345 , \19346 );
not \U$18971 ( \19348 , \16795 );
not \U$18972 ( \19349 , \16855 );
or \U$18973 ( \19350 , \19348 , \19349 );
or \U$18974 ( \19351 , \16855 , \16795 );
nand \U$18975 ( \19352 , \19350 , \19351 );
xor \U$18976 ( \19353 , \16762 , \16776 );
xor \U$18977 ( \19354 , \19353 , \16792 );
not \U$18978 ( \19355 , \6214 );
not \U$18979 ( \19356 , \18477 );
or \U$18980 ( \19357 , \19355 , \19356 );
and \U$18981 ( \19358 , RIae79ef8_167, \1859 );
not \U$18982 ( \19359 , RIae79ef8_167);
and \U$18983 ( \19360 , \19359 , \17596 );
or \U$18984 ( \19361 , \19358 , \19360 );
buf \U$18985 ( \19362 , \6199 );
nand \U$18986 ( \19363 , \19361 , \19362 );
nand \U$18987 ( \19364 , \19357 , \19363 );
not \U$18988 ( \19365 , \11914 );
xnor \U$18989 ( \19366 , \4112 , RIae79fe8_169);
not \U$18990 ( \19367 , \19366 );
or \U$18991 ( \19368 , \19365 , \19367 );
nand \U$18992 ( \19369 , \18467 , \9517 );
nand \U$18993 ( \19370 , \19368 , \19369 );
xor \U$18994 ( \19371 , \19364 , \19370 );
not \U$18995 ( \19372 , \10667 );
not \U$18996 ( \19373 , \2207 );
and \U$18997 ( \19374 , RIae7a150_172, \19373 );
not \U$18998 ( \19375 , RIae7a150_172);
and \U$18999 ( \19376 , \19375 , \2207 );
or \U$19000 ( \19377 , \19374 , \19376 );
not \U$19001 ( \19378 , \19377 );
or \U$19002 ( \19379 , \19372 , \19378 );
nand \U$19003 ( \19380 , \18488 , \9776 );
nand \U$19004 ( \19381 , \19379 , \19380 );
and \U$19005 ( \19382 , \19371 , \19381 );
and \U$19006 ( \19383 , \19364 , \19370 );
or \U$19007 ( \19384 , \19382 , \19383 );
xor \U$19008 ( \19385 , \19354 , \19384 );
xor \U$19009 ( \19386 , \16901 , \16916 );
xor \U$19010 ( \19387 , \19386 , \16929 );
not \U$19011 ( \19388 , \16383 );
and \U$19012 ( \19389 , RIae7aa38_191, \9761 );
not \U$19013 ( \19390 , RIae7aa38_191);
and \U$19014 ( \19391 , \19390 , \1022 );
nor \U$19015 ( \19392 , \19389 , \19391 );
not \U$19016 ( \19393 , \19392 );
or \U$19017 ( \19394 , \19388 , \19393 );
nand \U$19018 ( \19395 , \18416 , RIae7aab0_192);
nand \U$19019 ( \19396 , \19394 , \19395 );
xor \U$19020 ( \19397 , \19387 , \19396 );
not \U$19021 ( \19398 , \16564 );
not \U$19022 ( \19399 , RIae7a498_179);
not \U$19023 ( \19400 , \10567 );
not \U$19024 ( \19401 , \19400 );
or \U$19025 ( \19402 , \19399 , \19401 );
not \U$19026 ( \19403 , \14023 );
or \U$19027 ( \19404 , \19403 , RIae7a498_179);
nand \U$19028 ( \19405 , \19402 , \19404 );
not \U$19029 ( \19406 , \19405 );
or \U$19030 ( \19407 , \19398 , \19406 );
nand \U$19031 ( \19408 , \18387 , \10677 );
nand \U$19032 ( \19409 , \19407 , \19408 );
and \U$19033 ( \19410 , \19397 , \19409 );
and \U$19034 ( \19411 , \19387 , \19396 );
or \U$19035 ( \19412 , \19410 , \19411 );
and \U$19036 ( \19413 , \19385 , \19412 );
and \U$19037 ( \19414 , \19354 , \19384 );
or \U$19038 ( \19415 , \19413 , \19414 );
xor \U$19039 ( \19416 , \19352 , \19415 );
xor \U$19040 ( \19417 , \16871 , \16933 );
not \U$19041 ( \19418 , \9828 );
not \U$19042 ( \19419 , RIae794a8_145);
not \U$19043 ( \19420 , \15488 );
or \U$19044 ( \19421 , \19419 , \19420 );
buf \U$19045 ( \19422 , \14156 );
or \U$19046 ( \19423 , \19422 , RIae794a8_145);
nand \U$19047 ( \19424 , \19421 , \19423 );
not \U$19048 ( \19425 , \19424 );
or \U$19049 ( \19426 , \19418 , \19425 );
nand \U$19050 ( \19427 , \16790 , \1919 );
nand \U$19051 ( \19428 , \19426 , \19427 );
not \U$19052 ( \19429 , \11762 );
not \U$19053 ( \19430 , RIae79ca0_162);
not \U$19054 ( \19431 , \4960 );
or \U$19055 ( \19432 , \19430 , \19431 );
or \U$19056 ( \19433 , \4960 , RIae79ca0_162);
nand \U$19057 ( \19434 , \19432 , \19433 );
not \U$19058 ( \19435 , \19434 );
or \U$19059 ( \19436 , \19429 , \19435 );
nand \U$19060 ( \19437 , \16869 , \4853 );
nand \U$19061 ( \19438 , \19436 , \19437 );
xor \U$19062 ( \19439 , \19428 , \19438 );
not \U$19063 ( \19440 , \14510 );
not \U$19064 ( \19441 , \11207 );
not \U$19065 ( \19442 , \1118 );
or \U$19066 ( \19443 , \19441 , \19442 );
or \U$19067 ( \19444 , \12801 , \18088 );
nand \U$19068 ( \19445 , \19443 , \19444 );
not \U$19069 ( \19446 , \19445 );
or \U$19070 ( \19447 , \19440 , \19446 );
nand \U$19071 ( \19448 , \18895 , \10275 );
nand \U$19072 ( \19449 , \19447 , \19448 );
and \U$19073 ( \19450 , \19439 , \19449 );
and \U$19074 ( \19451 , \19428 , \19438 );
or \U$19075 ( \19452 , \19450 , \19451 );
xor \U$19076 ( \19453 , \19417 , \19452 );
not \U$19077 ( \19454 , \9792 );
not \U$19078 ( \19455 , RIae7a2b8_175);
not \U$19079 ( \19456 , \6413 );
not \U$19080 ( \19457 , \19456 );
or \U$19081 ( \19458 , \19455 , \19457 );
nand \U$19082 ( \19459 , \15782 , \9799 );
nand \U$19083 ( \19460 , \19458 , \19459 );
not \U$19084 ( \19461 , \19460 );
or \U$19085 ( \19462 , \19454 , \19461 );
nand \U$19086 ( \19463 , \18425 , \9814 );
nand \U$19087 ( \19464 , \19462 , \19463 );
not \U$19088 ( \19465 , \19464 );
buf \U$19089 ( \19466 , \9687 );
not \U$19090 ( \19467 , \19466 );
not \U$19091 ( \19468 , RIae7a240_174);
not \U$19092 ( \19469 , \10883 );
or \U$19093 ( \19470 , \19468 , \19469 );
or \U$19094 ( \19471 , \10883 , RIae7a240_174);
nand \U$19095 ( \19472 , \19470 , \19471 );
not \U$19096 ( \19473 , \19472 );
or \U$19097 ( \19474 , \19467 , \19473 );
nand \U$19098 ( \19475 , \18354 , \9699 );
nand \U$19099 ( \19476 , \19474 , \19475 );
not \U$19100 ( \19477 , \9729 );
not \U$19101 ( \19478 , \1878 );
xor \U$19102 ( \19479 , RIae7a060_170, \19478 );
not \U$19103 ( \19480 , \19479 );
or \U$19104 ( \19481 , \19477 , \19480 );
nand \U$19105 ( \19482 , \18434 , \10542 );
nand \U$19106 ( \19483 , \19481 , \19482 );
xor \U$19107 ( \19484 , \19476 , \19483 );
not \U$19108 ( \19485 , \19484 );
or \U$19109 ( \19486 , \19465 , \19485 );
nand \U$19110 ( \19487 , \19476 , \19483 );
nand \U$19111 ( \19488 , \19486 , \19487 );
and \U$19112 ( \19489 , \19453 , \19488 );
and \U$19113 ( \19490 , \19417 , \19452 );
or \U$19114 ( \19491 , \19489 , \19490 );
and \U$19115 ( \19492 , \19416 , \19491 );
and \U$19116 ( \19493 , \19352 , \19415 );
or \U$19117 ( \19494 , \19492 , \19493 );
xor \U$19118 ( \19495 , \19347 , \19494 );
xor \U$19119 ( \19496 , \17084 , \17205 );
xor \U$19120 ( \19497 , \19496 , \17204 );
and \U$19121 ( \19498 , \19495 , \19497 );
and \U$19122 ( \19499 , \19347 , \19494 );
or \U$19123 ( \19500 , \19498 , \19499 );
not \U$19124 ( \19501 , \19500 );
nand \U$19125 ( \19502 , \19193 , \19501 );
not \U$19126 ( \19503 , \19502 );
or \U$19127 ( \19504 , \19191 , \19503 );
or \U$19128 ( \19505 , \19193 , \19501 );
nand \U$19129 ( \19506 , \19504 , \19505 );
not \U$19130 ( \19507 , \19506 );
or \U$19131 ( \19508 , \18941 , \19507 );
not \U$19132 ( \19509 , \19506 );
not \U$19133 ( \19510 , \19509 );
not \U$19134 ( \19511 , \18939 );
or \U$19135 ( \19512 , \19510 , \19511 );
not \U$19136 ( \19513 , \18852 );
xor \U$19137 ( \19514 , \18926 , \18853 );
not \U$19138 ( \19515 , \19514 );
or \U$19139 ( \19516 , \19513 , \19515 );
or \U$19140 ( \19517 , \18852 , \19514 );
nand \U$19141 ( \19518 , \19516 , \19517 );
not \U$19142 ( \19519 , \19518 );
xor \U$19143 ( \19520 , \18336 , \18446 );
xor \U$19144 ( \19521 , \19520 , \18497 );
xor \U$19145 ( \19522 , \18180 , \18160 );
xor \U$19146 ( \19523 , \19522 , \18097 );
xor \U$19147 ( \19524 , \19521 , \19523 );
xor \U$19148 ( \19525 , \18864 , \18874 );
xor \U$19149 ( \19526 , \19525 , \18920 );
and \U$19150 ( \19527 , \19524 , \19526 );
and \U$19151 ( \19528 , \19521 , \19523 );
or \U$19152 ( \19529 , \19527 , \19528 );
not \U$19153 ( \19530 , \19529 );
nand \U$19154 ( \19531 , \18505 , \18502 );
and \U$19155 ( \19532 , \19531 , \18185 );
not \U$19156 ( \19533 , \19531 );
not \U$19157 ( \19534 , \18185 );
and \U$19158 ( \19535 , \19533 , \19534 );
nor \U$19159 ( \19536 , \19532 , \19535 );
not \U$19160 ( \19537 , \19536 );
or \U$19161 ( \19538 , \19530 , \19537 );
or \U$19162 ( \19539 , \19529 , \19536 );
nand \U$19163 ( \19540 , \19538 , \19539 );
not \U$19164 ( \19541 , \19540 );
or \U$19165 ( \19542 , \19519 , \19541 );
not \U$19166 ( \19543 , \19536 );
nand \U$19167 ( \19544 , \19543 , \19529 );
nand \U$19168 ( \19545 , \19542 , \19544 );
nand \U$19169 ( \19546 , \19512 , \19545 );
nand \U$19170 ( \19547 , \19508 , \19546 );
not \U$19171 ( \19548 , \19547 );
xnor \U$19172 ( \19549 , \18933 , \19548 );
not \U$19173 ( \19550 , \18940 );
not \U$19174 ( \19551 , \19509 );
or \U$19175 ( \19552 , \19550 , \19551 );
nand \U$19176 ( \19553 , \19506 , \18939 );
nand \U$19177 ( \19554 , \19552 , \19553 );
not \U$19178 ( \19555 , \19545 );
and \U$19179 ( \19556 , \19554 , \19555 );
not \U$19180 ( \19557 , \19554 );
and \U$19181 ( \19558 , \19557 , \19545 );
nor \U$19182 ( \19559 , \19556 , \19558 );
not \U$19183 ( \19560 , \19559 );
not \U$19184 ( \19561 , \19560 );
xor \U$19185 ( \19562 , \18842 , \18844 );
xor \U$19186 ( \19563 , \19562 , \18928 );
not \U$19187 ( \19564 , \19563 );
or \U$19188 ( \19565 , \19561 , \19564 );
not \U$19189 ( \19566 , \19563 );
nand \U$19190 ( \19567 , \19566 , \19559 );
not \U$19191 ( \19568 , \19242 );
not \U$19192 ( \19569 , \19210 );
and \U$19193 ( \19570 , \19568 , \19569 );
and \U$19194 ( \19571 , \19242 , \19210 );
nor \U$19195 ( \19572 , \19570 , \19571 );
not \U$19196 ( \19573 , \19572 );
not \U$19197 ( \19574 , \19573 );
and \U$19198 ( \19575 , \18439 , \18418 );
not \U$19199 ( \19576 , \18439 );
not \U$19200 ( \19577 , \18418 );
and \U$19201 ( \19578 , \19576 , \19577 );
nor \U$19202 ( \19579 , \19575 , \19578 );
not \U$19203 ( \19580 , \19579 );
not \U$19204 ( \19581 , \19580 );
or \U$19205 ( \19582 , \19574 , \19581 );
nand \U$19206 ( \19583 , \19579 , \19572 );
nand \U$19207 ( \19584 , \19582 , \19583 );
xor \U$19208 ( \19585 , \18492 , \18469 );
xnor \U$19209 ( \19586 , \19585 , \18479 );
not \U$19210 ( \19587 , \19586 );
nand \U$19211 ( \19588 , \19584 , \19587 );
nand \U$19212 ( \19589 , \19579 , \19573 );
and \U$19213 ( \19590 , \19588 , \19589 );
xor \U$19214 ( \19591 , \18019 , \18056 );
xor \U$19215 ( \19592 , \19591 , \18094 );
not \U$19216 ( \19593 , \19592 );
and \U$19217 ( \19594 , \19590 , \19593 );
not \U$19218 ( \19595 , \19590 );
and \U$19219 ( \19596 , \19595 , \19592 );
nor \U$19220 ( \19597 , \19594 , \19596 );
not \U$19221 ( \19598 , \19597 );
not \U$19222 ( \19599 , \11851 );
not \U$19223 ( \19600 , RIae7a7e0_186);
not \U$19224 ( \19601 , \2049 );
or \U$19225 ( \19602 , \19600 , \19601 );
or \U$19226 ( \19603 , \13033 , RIae7a7e0_186);
nand \U$19227 ( \19604 , \19602 , \19603 );
not \U$19228 ( \19605 , \19604 );
or \U$19229 ( \19606 , \19599 , \19605 );
nand \U$19230 ( \19607 , \19140 , \10519 );
nand \U$19231 ( \19608 , \19606 , \19607 );
not \U$19232 ( \19609 , \9622 );
not \U$19233 ( \19610 , \19115 );
or \U$19234 ( \19611 , \19609 , \19610 );
not \U$19235 ( \19612 , \11690 );
not \U$19236 ( \19613 , \1753 );
or \U$19237 ( \19614 , \19612 , \19613 );
or \U$19238 ( \19615 , \1759 , \11690 );
nand \U$19239 ( \19616 , \19614 , \19615 );
nand \U$19240 ( \19617 , \19616 , \11014 );
nand \U$19241 ( \19618 , \19611 , \19617 );
xor \U$19242 ( \19619 , \19608 , \19618 );
not \U$19243 ( \19620 , \13720 );
and \U$19244 ( \19621 , \2757 , RIae7a240_174);
not \U$19245 ( \19622 , \2757 );
not \U$19246 ( \19623 , RIae7a240_174);
and \U$19247 ( \19624 , \19622 , \19623 );
nor \U$19248 ( \19625 , \19621 , \19624 );
not \U$19249 ( \19626 , \19625 );
or \U$19250 ( \19627 , \19620 , \19626 );
nand \U$19251 ( \19628 , \19472 , \9699 );
nand \U$19252 ( \19629 , \19627 , \19628 );
and \U$19253 ( \19630 , \19619 , \19629 );
and \U$19254 ( \19631 , \19608 , \19618 );
or \U$19255 ( \19632 , \19630 , \19631 );
not \U$19256 ( \19633 , \19632 );
xor \U$19257 ( \19634 , \19310 , \19320 );
xor \U$19258 ( \19635 , \19634 , \19332 );
not \U$19259 ( \19636 , \19635 );
not \U$19260 ( \19637 , \19636 );
xor \U$19261 ( \19638 , \19281 , \19259 );
xnor \U$19262 ( \19639 , \19638 , \19290 );
not \U$19263 ( \19640 , \19639 );
or \U$19264 ( \19641 , \19637 , \19640 );
or \U$19265 ( \19642 , \19639 , \19636 );
nand \U$19266 ( \19643 , \19641 , \19642 );
not \U$19267 ( \19644 , \19643 );
or \U$19268 ( \19645 , \19633 , \19644 );
nand \U$19269 ( \19646 , \19639 , \19635 );
nand \U$19270 ( \19647 , \19645 , \19646 );
not \U$19271 ( \19648 , \19647 );
not \U$19272 ( \19649 , \19339 );
not \U$19273 ( \19650 , \19296 );
not \U$19274 ( \19651 , \19650 );
or \U$19275 ( \19652 , \19649 , \19651 );
or \U$19276 ( \19653 , \19650 , \19339 );
nand \U$19277 ( \19654 , \19652 , \19653 );
not \U$19278 ( \19655 , \19654 );
not \U$19279 ( \19656 , \2450 );
not \U$19280 ( \19657 , \19216 );
or \U$19281 ( \19658 , \19656 , \19657 );
and \U$19282 ( \19659 , RIae79778_151, \16274 );
not \U$19283 ( \19660 , RIae79778_151);
buf \U$19284 ( \19661 , \16271 );
and \U$19285 ( \19662 , \19660 , \19661 );
nor \U$19286 ( \19663 , \19659 , \19662 );
nand \U$19287 ( \19664 , \19663 , \2431 );
nand \U$19288 ( \19665 , \19658 , \19664 );
not \U$19289 ( \19666 , \1910 );
xor \U$19290 ( \19667 , RIae793b8_143, \10031 );
not \U$19291 ( \19668 , \19667 );
or \U$19292 ( \19669 , \19666 , \19668 );
nand \U$19293 ( \19670 , \19040 , \1863 );
nand \U$19294 ( \19671 , \19669 , \19670 );
not \U$19295 ( \19672 , \19671 );
not \U$19296 ( \19673 , \1059 );
not \U$19297 ( \19674 , \12858 );
or \U$19298 ( \19675 , \19673 , \19674 );
nand \U$19299 ( \19676 , \19675 , \1297 );
not \U$19300 ( \19677 , \19676 );
not \U$19301 ( \19678 , \18991 );
or \U$19302 ( \19679 , \19678 , \1203 );
xnor \U$19303 ( \19680 , \12857 , RIae79070_136);
not \U$19304 ( \19681 , \1061 );
or \U$19305 ( \19682 , \19680 , \19681 );
nand \U$19306 ( \19683 , \19679 , \19682 );
nand \U$19307 ( \19684 , \19677 , \19683 );
not \U$19308 ( \19685 , \19684 );
not \U$19309 ( \19686 , \1501 );
not \U$19310 ( \19687 , \19006 );
or \U$19311 ( \19688 , \19686 , \19687 );
not \U$19312 ( \19689 , \11576 );
and \U$19313 ( \19690 , \19689 , \12647 );
not \U$19314 ( \19691 , \19689 );
and \U$19315 ( \19692 , \19691 , RIae79250_140);
nor \U$19316 ( \19693 , \19690 , \19692 );
nand \U$19317 ( \19694 , \19693 , \1497 );
nand \U$19318 ( \19695 , \19688 , \19694 );
not \U$19319 ( \19696 , \19695 );
or \U$19320 ( \19697 , \19685 , \19696 );
or \U$19321 ( \19698 , \19695 , \19684 );
nand \U$19322 ( \19699 , \19697 , \19698 );
not \U$19323 ( \19700 , \19699 );
or \U$19324 ( \19701 , \19672 , \19700 );
not \U$19325 ( \19702 , \19684 );
nand \U$19326 ( \19703 , \19702 , \19695 );
nand \U$19327 ( \19704 , \19701 , \19703 );
xor \U$19328 ( \19705 , \19665 , \19704 );
not \U$19329 ( \19706 , \19705 );
not \U$19330 ( \19707 , \2519 );
not \U$19331 ( \19708 , \19286 );
or \U$19332 ( \19709 , \19707 , \19708 );
not \U$19333 ( \19710 , \1991 );
not \U$19334 ( \19711 , \15091 );
or \U$19335 ( \19712 , \19710 , \19711 );
not \U$19336 ( \19713 , RIae797f0_152);
or \U$19337 ( \19714 , \14691 , \19713 );
nand \U$19338 ( \19715 , \19712 , \19714 );
nand \U$19339 ( \19716 , \19715 , \1989 );
nand \U$19340 ( \19717 , \19709 , \19716 );
not \U$19341 ( \19718 , \19717 );
or \U$19342 ( \19719 , \19706 , \19718 );
nand \U$19343 ( \19720 , \19704 , \19665 );
nand \U$19344 ( \19721 , \19719 , \19720 );
not \U$19345 ( \19722 , \3440 );
not \U$19346 ( \19723 , \19308 );
or \U$19347 ( \19724 , \19722 , \19723 );
not \U$19348 ( \19725 , RIae79520_146);
not \U$19349 ( \19726 , \10461 );
or \U$19350 ( \19727 , \19725 , \19726 );
or \U$19351 ( \19728 , \10461 , RIae79520_146);
nand \U$19352 ( \19729 , \19727 , \19728 );
nand \U$19353 ( \19730 , \19729 , \12680 );
nand \U$19354 ( \19731 , \19724 , \19730 );
not \U$19355 ( \19732 , \19731 );
nand \U$19356 ( \19733 , \19257 , \2322 );
and \U$19357 ( \19734 , RIae798e0_154, \14657 );
not \U$19358 ( \19735 , RIae798e0_154);
not \U$19359 ( \19736 , \13301 );
and \U$19360 ( \19737 , \19735 , \19736 );
or \U$19361 ( \19738 , \19734 , \19737 );
nand \U$19362 ( \19739 , \19738 , \10807 );
nand \U$19363 ( \19740 , \19732 , \19733 , \19739 );
not \U$19364 ( \19741 , \19740 );
not \U$19365 ( \19742 , \6091 );
and \U$19366 ( \19743 , \4169 , RIae79d90_164);
not \U$19367 ( \19744 , \4169 );
and \U$19368 ( \19745 , \19744 , \6084 );
nor \U$19369 ( \19746 , \19743 , \19745 );
not \U$19370 ( \19747 , \19746 );
or \U$19371 ( \19748 , \19742 , \19747 );
not \U$19372 ( \19749 , \19329 );
nand \U$19373 ( \19750 , \19749 , \14940 );
nand \U$19374 ( \19751 , \19748 , \19750 );
not \U$19375 ( \19752 , \19751 );
or \U$19376 ( \19753 , \19741 , \19752 );
nand \U$19377 ( \19754 , \19733 , \19739 );
nand \U$19378 ( \19755 , \19754 , \19731 );
nand \U$19379 ( \19756 , \19753 , \19755 );
xor \U$19380 ( \19757 , \19721 , \19756 );
not \U$19381 ( \19758 , \1919 );
not \U$19382 ( \19759 , \19424 );
or \U$19383 ( \19760 , \19758 , \19759 );
and \U$19384 ( \19761 , RIae794a8_145, \9412 );
not \U$19385 ( \19762 , RIae794a8_145);
and \U$19386 ( \19763 , \19762 , \11198 );
or \U$19387 ( \19764 , \19761 , \19763 );
nand \U$19388 ( \19765 , \19764 , \2457 );
nand \U$19389 ( \19766 , \19760 , \19765 );
not \U$19390 ( \19767 , \2776 );
not \U$19391 ( \19768 , \19315 );
or \U$19392 ( \19769 , \19767 , \19768 );
and \U$19393 ( \19770 , RIae79c28_161, \9290 );
not \U$19394 ( \19771 , RIae79c28_161);
and \U$19395 ( \19772 , \19771 , \9286 );
nor \U$19396 ( \19773 , \19770 , \19772 );
nand \U$19397 ( \19774 , \19773 , \2767 );
nand \U$19398 ( \19775 , \19769 , \19774 );
xor \U$19399 ( \19776 , \19766 , \19775 );
not \U$19400 ( \19777 , \4853 );
not \U$19401 ( \19778 , \19434 );
or \U$19402 ( \19779 , \19777 , \19778 );
not \U$19403 ( \19780 , \4844 );
not \U$19404 ( \19781 , \5109 );
or \U$19405 ( \19782 , \19780 , \19781 );
nand \U$19406 ( \19783 , \15128 , RIae79ca0_162);
nand \U$19407 ( \19784 , \19782 , \19783 );
nand \U$19408 ( \19785 , \19784 , \4842 );
nand \U$19409 ( \19786 , \19779 , \19785 );
and \U$19410 ( \19787 , \19776 , \19786 );
and \U$19411 ( \19788 , \19766 , \19775 );
or \U$19412 ( \19789 , \19787 , \19788 );
and \U$19413 ( \19790 , \19757 , \19789 );
and \U$19414 ( \19791 , \19721 , \19756 );
or \U$19415 ( \19792 , \19790 , \19791 );
not \U$19416 ( \19793 , \19792 );
nand \U$19417 ( \19794 , \19655 , \19793 );
not \U$19418 ( \19795 , \19794 );
or \U$19419 ( \19796 , \19648 , \19795 );
nand \U$19420 ( \19797 , \19654 , \19792 );
nand \U$19421 ( \19798 , \19796 , \19797 );
not \U$19422 ( \19799 , \19798 );
or \U$19423 ( \19800 , \19598 , \19799 );
not \U$19424 ( \19801 , \19590 );
nand \U$19425 ( \19802 , \19801 , \19592 );
nand \U$19426 ( \19803 , \19800 , \19802 );
xor \U$19427 ( \19804 , \19347 , \19494 );
xor \U$19428 ( \19805 , \19804 , \19497 );
xor \U$19429 ( \19806 , \19803 , \19805 );
xor \U$19430 ( \19807 , \19352 , \19415 );
xor \U$19431 ( \19808 , \19807 , \19491 );
xor \U$19432 ( \19809 , \19195 , \19247 );
xor \U$19433 ( \19810 , \19809 , \19344 );
or \U$19434 ( \19811 , \19808 , \19810 );
not \U$19435 ( \19812 , \19811 );
not \U$19436 ( \19813 , \9814 );
not \U$19437 ( \19814 , \19460 );
or \U$19438 ( \19815 , \19813 , \19814 );
and \U$19439 ( \19816 , \2089 , RIae7a2b8_175);
not \U$19440 ( \19817 , \2089 );
and \U$19441 ( \19818 , \19817 , \9810 );
nor \U$19442 ( \19819 , \19816 , \19818 );
nand \U$19443 ( \19820 , \19819 , \9792 );
nand \U$19444 ( \19821 , \19815 , \19820 );
not \U$19445 ( \19822 , \19821 );
not \U$19446 ( \19823 , \9745 );
not \U$19447 ( \19824 , \19479 );
or \U$19448 ( \19825 , \19823 , \19824 );
not \U$19449 ( \19826 , \11102 );
not \U$19450 ( \19827 , \3294 );
or \U$19451 ( \19828 , \19826 , \19827 );
or \U$19452 ( \19829 , \9807 , \14721 );
nand \U$19453 ( \19830 , \19828 , \19829 );
nand \U$19454 ( \19831 , \19830 , \9730 );
nand \U$19455 ( \19832 , \19825 , \19831 );
not \U$19456 ( \19833 , \19832 );
not \U$19457 ( \19834 , \19833 );
not \U$19458 ( \19835 , \9517 );
not \U$19459 ( \19836 , \19366 );
or \U$19460 ( \19837 , \19835 , \19836 );
and \U$19461 ( \19838 , RIae79fe8_169, \3216 );
not \U$19462 ( \19839 , RIae79fe8_169);
and \U$19463 ( \19840 , \19839 , \14422 );
or \U$19464 ( \19841 , \19838 , \19840 );
nand \U$19465 ( \19842 , \19841 , \9499 );
nand \U$19466 ( \19843 , \19837 , \19842 );
not \U$19467 ( \19844 , \19843 );
or \U$19468 ( \19845 , \19834 , \19844 );
or \U$19469 ( \19846 , \19843 , \19833 );
nand \U$19470 ( \19847 , \19845 , \19846 );
not \U$19471 ( \19848 , \19847 );
or \U$19472 ( \19849 , \19822 , \19848 );
nand \U$19473 ( \19850 , \19843 , \19832 );
nand \U$19474 ( \19851 , \19849 , \19850 );
not \U$19475 ( \19852 , \19851 );
nand \U$19476 ( \19853 , \19377 , \9777 );
not \U$19477 ( \19854 , \10672 );
not \U$19478 ( \19855 , \11885 );
or \U$19479 ( \19856 , \19854 , \19855 );
not \U$19480 ( \19857 , \2993 );
or \U$19481 ( \19858 , \19857 , \9750 );
nand \U$19482 ( \19859 , \19856 , \19858 );
nand \U$19483 ( \19860 , \19859 , \11087 );
and \U$19484 ( \19861 , \19361 , \10573 );
not \U$19485 ( \19862 , RIae79ef8_167);
not \U$19486 ( \19863 , \2402 );
or \U$19487 ( \19864 , \19862 , \19863 );
or \U$19488 ( \19865 , \10492 , RIae79ef8_167);
nand \U$19489 ( \19866 , \19864 , \19865 );
not \U$19490 ( \19867 , \19866 );
not \U$19491 ( \19868 , \19362 );
nor \U$19492 ( \19869 , \19867 , \19868 );
nor \U$19493 ( \19870 , \19861 , \19869 );
nand \U$19494 ( \19871 , \19853 , \19860 , \19870 );
not \U$19495 ( \19872 , \19871 );
not \U$19496 ( \19873 , \12371 );
not \U$19497 ( \19874 , \19405 );
or \U$19498 ( \19875 , \19873 , \19874 );
and \U$19499 ( \19876 , RIae7a498_179, \14712 );
not \U$19500 ( \19877 , RIae7a498_179);
and \U$19501 ( \19878 , \19877 , \5631 );
or \U$19502 ( \19879 , \19876 , \19878 );
nand \U$19503 ( \19880 , \19879 , \16564 );
nand \U$19504 ( \19881 , \19875 , \19880 );
not \U$19505 ( \19882 , \19881 );
or \U$19506 ( \19883 , \19872 , \19882 );
not \U$19507 ( \19884 , \19870 );
nand \U$19508 ( \19885 , \19853 , \19860 );
nand \U$19509 ( \19886 , \19884 , \19885 );
nand \U$19510 ( \19887 , \19883 , \19886 );
xor \U$19511 ( \19888 , \19428 , \19438 );
xor \U$19512 ( \19889 , \19888 , \19449 );
xor \U$19513 ( \19890 , \19887 , \19889 );
not \U$19514 ( \19891 , \19890 );
or \U$19515 ( \19892 , \19852 , \19891 );
nand \U$19516 ( \19893 , \19889 , \19887 );
nand \U$19517 ( \19894 , \19892 , \19893 );
not \U$19518 ( \19895 , \19894 );
xor \U$19519 ( \19896 , \19233 , \19226 );
xnor \U$19520 ( \19897 , \19896 , \19220 );
not \U$19521 ( \19898 , \19897 );
and \U$19522 ( \19899 , \19202 , \19207 );
not \U$19523 ( \19900 , \19202 );
not \U$19524 ( \19901 , \19207 );
and \U$19525 ( \19902 , \19900 , \19901 );
nor \U$19526 ( \19903 , \19899 , \19902 );
not \U$19527 ( \19904 , \19903 );
nand \U$19528 ( \19905 , \19898 , \19904 );
not \U$19529 ( \19906 , \19905 );
not \U$19530 ( \19907 , \10637 );
xor \U$19531 ( \19908 , RIae7a510_180, \3747 );
not \U$19532 ( \19909 , \19908 );
or \U$19533 ( \19910 , \19907 , \19909 );
nand \U$19534 ( \19911 , \19129 , \12233 );
nand \U$19535 ( \19912 , \19910 , \19911 );
not \U$19536 ( \19913 , \19912 );
not \U$19537 ( \19914 , \19277 );
not \U$19538 ( \19915 , \19271 );
and \U$19539 ( \19916 , \19914 , \19915 );
and \U$19540 ( \19917 , \19277 , \19271 );
nor \U$19541 ( \19918 , \19916 , \19917 );
not \U$19542 ( \19919 , \19918 );
and \U$19543 ( \19920 , \19913 , \19919 );
and \U$19544 ( \19921 , \19912 , \19918 );
nor \U$19545 ( \19922 , \19920 , \19921 );
not \U$19546 ( \19923 , \19922 );
not \U$19547 ( \19924 , \19923 );
not \U$19548 ( \19925 , \10275 );
not \U$19549 ( \19926 , \19445 );
or \U$19550 ( \19927 , \19925 , \19926 );
not \U$19551 ( \19928 , RIae7a8d0_188);
not \U$19552 ( \19929 , \5081 );
or \U$19553 ( \19930 , \19928 , \19929 );
or \U$19554 ( \19931 , \5081 , RIae7a8d0_188);
nand \U$19555 ( \19932 , \19930 , \19931 );
nand \U$19556 ( \19933 , \19932 , \11205 );
nand \U$19557 ( \19934 , \19927 , \19933 );
not \U$19558 ( \19935 , \19934 );
or \U$19559 ( \19936 , \19924 , \19935 );
not \U$19560 ( \19937 , \19918 );
nand \U$19561 ( \19938 , \19937 , \19912 );
nand \U$19562 ( \19939 , \19936 , \19938 );
not \U$19563 ( \19940 , \19939 );
or \U$19564 ( \19941 , \19906 , \19940 );
nand \U$19565 ( \19942 , \19903 , \19897 );
nand \U$19566 ( \19943 , \19941 , \19942 );
not \U$19567 ( \19944 , \19943 );
or \U$19568 ( \19945 , \19895 , \19944 );
xnor \U$19569 ( \19946 , \19159 , \19108 );
not \U$19570 ( \19947 , \19946 );
xor \U$19571 ( \19948 , \19943 , \19894 );
nand \U$19572 ( \19949 , \19947 , \19948 );
nand \U$19573 ( \19950 , \19945 , \19949 );
not \U$19574 ( \19951 , \19950 );
or \U$19575 ( \19952 , \19812 , \19951 );
nand \U$19576 ( \19953 , \19808 , \19810 );
nand \U$19577 ( \19954 , \19952 , \19953 );
and \U$19578 ( \19955 , \19806 , \19954 );
and \U$19579 ( \19956 , \19803 , \19805 );
or \U$19580 ( \19957 , \19955 , \19956 );
not \U$19581 ( \19958 , \19500 );
not \U$19582 ( \19959 , \19193 );
or \U$19583 ( \19960 , \19958 , \19959 );
or \U$19584 ( \19961 , \19193 , \19500 );
nand \U$19585 ( \19962 , \19960 , \19961 );
xor \U$19586 ( \19963 , \19190 , \19962 );
xor \U$19587 ( \19964 , \19957 , \19963 );
xor \U$19588 ( \19965 , \19518 , \19540 );
and \U$19589 ( \19966 , \19964 , \19965 );
and \U$19590 ( \19967 , \19957 , \19963 );
or \U$19591 ( \19968 , \19966 , \19967 );
nand \U$19592 ( \19969 , \19567 , \19968 );
nand \U$19593 ( \19970 , \19565 , \19969 );
or \U$19594 ( \19971 , \19549 , \19970 );
xor \U$19595 ( \19972 , \18603 , \18785 );
and \U$19596 ( \19973 , \19972 , \18838 );
and \U$19597 ( \19974 , \18603 , \18785 );
or \U$19598 ( \19975 , \19973 , \19974 );
xor \U$19599 ( \19976 , \17877 , \17881 );
and \U$19600 ( \19977 , \19976 , \17936 );
and \U$19601 ( \19978 , \17877 , \17881 );
or \U$19602 ( \19979 , \19977 , \19978 );
and \U$19603 ( \19980 , \14757 , \14771 );
not \U$19604 ( \19981 , \14757 );
and \U$19605 ( \19982 , \19981 , \14770 );
nor \U$19606 ( \19983 , \19980 , \19982 );
not \U$19607 ( \19984 , \19983 );
not \U$19608 ( \19985 , \14784 );
and \U$19609 ( \19986 , \19984 , \19985 );
and \U$19610 ( \19987 , \14784 , \19983 );
nor \U$19611 ( \19988 , \19986 , \19987 );
not \U$19612 ( \19989 , \19988 );
xor \U$19613 ( \19990 , \12880 , \12892 );
and \U$19614 ( \19991 , \17568 , \17577 );
and \U$19615 ( \19992 , \17566 , \17567 );
nor \U$19616 ( \19993 , \19991 , \19992 );
xor \U$19617 ( \19994 , \19990 , \19993 );
not \U$19618 ( \19995 , \17593 );
not \U$19619 ( \19996 , \17583 );
nand \U$19620 ( \19997 , \19996 , \17586 );
not \U$19621 ( \19998 , \19997 );
or \U$19622 ( \19999 , \19995 , \19998 );
or \U$19623 ( \20000 , \19996 , \17586 );
nand \U$19624 ( \20001 , \19999 , \20000 );
xor \U$19625 ( \20002 , \19994 , \20001 );
not \U$19626 ( \20003 , \20002 );
or \U$19627 ( \20004 , \19989 , \20003 );
or \U$19628 ( \20005 , \20002 , \19988 );
nand \U$19629 ( \20006 , \20004 , \20005 );
not \U$19630 ( \20007 , \17465 );
not \U$19631 ( \20008 , \17456 );
or \U$19632 ( \20009 , \20007 , \20008 );
nand \U$19633 ( \20010 , \17455 , \17450 );
nand \U$19634 ( \20011 , \20009 , \20010 );
xnor \U$19635 ( \20012 , \20006 , \20011 );
not \U$19636 ( \20013 , \20012 );
not \U$19637 ( \20014 , \17551 );
not \U$19638 ( \20015 , \17559 );
nand \U$19639 ( \20016 , \20015 , \17641 );
not \U$19640 ( \20017 , \20016 );
or \U$19641 ( \20018 , \20014 , \20017 );
nand \U$19642 ( \20019 , \17559 , \17642 );
nand \U$19643 ( \20020 , \20018 , \20019 );
not \U$19644 ( \20021 , \20020 );
or \U$19645 ( \20022 , \20013 , \20021 );
or \U$19646 ( \20023 , \20012 , \20020 );
nand \U$19647 ( \20024 , \20022 , \20023 );
xor \U$19648 ( \20025 , \19979 , \20024 );
xor \U$19649 ( \20026 , \18662 , \18725 );
and \U$19650 ( \20027 , \20026 , \18784 );
and \U$19651 ( \20028 , \18662 , \18725 );
or \U$19652 ( \20029 , \20027 , \20028 );
and \U$19653 ( \20030 , \20025 , \20029 );
not \U$19654 ( \20031 , \20025 );
not \U$19655 ( \20032 , \20029 );
and \U$19656 ( \20033 , \20031 , \20032 );
nor \U$19657 ( \20034 , \20030 , \20033 );
not \U$19658 ( \20035 , \20034 );
xor \U$19659 ( \20036 , \17542 , \17546 );
and \U$19660 ( \20037 , \20036 , \17650 );
and \U$19661 ( \20038 , \17542 , \17546 );
or \U$19662 ( \20039 , \20037 , \20038 );
not \U$19663 ( \20040 , \20039 );
not \U$19664 ( \20041 , \20040 );
and \U$19665 ( \20042 , \20035 , \20041 );
and \U$19666 ( \20043 , \20034 , \20040 );
nor \U$19667 ( \20044 , \20042 , \20043 );
not \U$19668 ( \20045 , \20044 );
xor \U$19669 ( \20046 , \19975 , \20045 );
xor \U$19670 ( \20047 , \17311 , \17651 );
and \U$19671 ( \20048 , \20047 , \17949 );
and \U$19672 ( \20049 , \17311 , \17651 );
or \U$19673 ( \20050 , \20048 , \20049 );
xnor \U$19674 ( \20051 , \20046 , \20050 );
not \U$19675 ( \20052 , \20051 );
not \U$19676 ( \20053 , \17474 );
not \U$19677 ( \20054 , \17537 );
or \U$19678 ( \20055 , \20053 , \20054 );
not \U$19679 ( \20056 , \17470 );
nand \U$19680 ( \20057 , \20056 , \17444 );
nand \U$19681 ( \20058 , \20055 , \20057 );
not \U$19682 ( \20059 , \20058 );
not \U$19683 ( \20060 , \20059 );
not \U$19684 ( \20061 , \17887 );
nand \U$19685 ( \20062 , \20061 , \17893 );
not \U$19686 ( \20063 , \20062 );
not \U$19687 ( \20064 , \17899 );
or \U$19688 ( \20065 , \20063 , \20064 );
nand \U$19689 ( \20066 , \17892 , \17887 );
nand \U$19690 ( \20067 , \20065 , \20066 );
xor \U$19691 ( \20068 , \14535 , \14549 );
xnor \U$19692 ( \20069 , \20068 , \14541 );
xnor \U$19693 ( \20070 , \20067 , \20069 );
not \U$19694 ( \20071 , \20070 );
not \U$19695 ( \20072 , \17903 );
xor \U$19696 ( \20073 , \20072 , \17914 );
and \U$19697 ( \20074 , \20073 , \17908 );
and \U$19698 ( \20075 , \20072 , \17914 );
nor \U$19699 ( \20076 , \20074 , \20075 );
not \U$19700 ( \20077 , \20076 );
and \U$19701 ( \20078 , \20071 , \20077 );
and \U$19702 ( \20079 , \20070 , \20076 );
nor \U$19703 ( \20080 , \20078 , \20079 );
not \U$19704 ( \20081 , \20080 );
not \U$19705 ( \20082 , \17578 );
not \U$19706 ( \20083 , \17637 );
or \U$19707 ( \20084 , \20082 , \20083 );
xor \U$19708 ( \20085 , \17593 , \17587 );
nand \U$19709 ( \20086 , \20084 , \20085 );
not \U$19710 ( \20087 , \17578 );
nand \U$19711 ( \20088 , \20087 , \17636 );
nand \U$19712 ( \20089 , \20086 , \20088 );
nand \U$19713 ( \20090 , \20081 , \20089 );
not \U$19714 ( \20091 , \20089 );
nand \U$19715 ( \20092 , \20091 , \20080 );
nand \U$19716 ( \20093 , \20090 , \20092 );
not \U$19717 ( \20094 , \17900 );
nor \U$19718 ( \20095 , \17935 , \20094 );
or \U$19719 ( \20096 , \20095 , \17915 );
nand \U$19720 ( \20097 , \17935 , \20094 );
nand \U$19721 ( \20098 , \20096 , \20097 );
buf \U$19722 ( \20099 , \20098 );
not \U$19723 ( \20100 , \20099 );
and \U$19724 ( \20101 , \20093 , \20100 );
not \U$19725 ( \20102 , \20093 );
and \U$19726 ( \20103 , \20102 , \20099 );
nor \U$19727 ( \20104 , \20101 , \20103 );
not \U$19728 ( \20105 , \20104 );
not \U$19729 ( \20106 , \20105 );
or \U$19730 ( \20107 , \20060 , \20106 );
nand \U$19731 ( \20108 , \20104 , \20058 );
nand \U$19732 ( \20109 , \20107 , \20108 );
not \U$19733 ( \20110 , \17803 );
xor \U$19734 ( \20111 , \17767 , \17784 );
not \U$19735 ( \20112 , \20111 );
or \U$19736 ( \20113 , \20110 , \20112 );
nand \U$19737 ( \20114 , \17784 , \17767 );
nand \U$19738 ( \20115 , \20113 , \20114 );
not \U$19739 ( \20116 , \20115 );
not \U$19740 ( \20117 , \20116 );
not \U$19741 ( \20118 , \17865 );
not \U$19742 ( \20119 , \17826 );
nand \U$19743 ( \20120 , \20119 , \17835 );
not \U$19744 ( \20121 , \20120 );
or \U$19745 ( \20122 , \20118 , \20121 );
nand \U$19746 ( \20123 , \17832 , \17826 );
nand \U$19747 ( \20124 , \20122 , \20123 );
and \U$19748 ( \20125 , \14638 , \14648 );
not \U$19749 ( \20126 , \14638 );
not \U$19750 ( \20127 , \14648 );
and \U$19751 ( \20128 , \20126 , \20127 );
nor \U$19752 ( \20129 , \20125 , \20128 );
xor \U$19753 ( \20130 , \14568 , \14563 );
xnor \U$19754 ( \20131 , \20130 , \14582 );
xor \U$19755 ( \20132 , \20129 , \20131 );
xor \U$19756 ( \20133 , \14663 , \14697 );
xnor \U$19757 ( \20134 , \20133 , \14681 );
xor \U$19758 ( \20135 , \20132 , \20134 );
xor \U$19759 ( \20136 , \20124 , \20135 );
not \U$19760 ( \20137 , \20136 );
or \U$19761 ( \20138 , \20117 , \20137 );
or \U$19762 ( \20139 , \20116 , \20136 );
nand \U$19763 ( \20140 , \20138 , \20139 );
xnor \U$19764 ( \20141 , \20109 , \20140 );
not \U$19765 ( \20142 , \20141 );
not \U$19766 ( \20143 , \17942 );
not \U$19767 ( \20144 , \17937 );
or \U$19768 ( \20145 , \20143 , \20144 );
not \U$19769 ( \20146 , \17871 );
nand \U$19770 ( \20147 , \20146 , \17947 );
nand \U$19771 ( \20148 , \20145 , \20147 );
not \U$19772 ( \20149 , \20148 );
or \U$19773 ( \20150 , \20142 , \20149 );
or \U$19774 ( \20151 , \20141 , \20148 );
nand \U$19775 ( \20152 , \20150 , \20151 );
not \U$19776 ( \20153 , \17533 );
not \U$19777 ( \20154 , \17482 );
or \U$19778 ( \20155 , \20153 , \20154 );
or \U$19779 ( \20156 , \17482 , \17533 );
nand \U$19780 ( \20157 , \20156 , \17521 );
nand \U$19781 ( \20158 , \20155 , \20157 );
xor \U$19782 ( \20159 , \14416 , \14428 );
nand \U$19783 ( \20160 , \18694 , \18700 );
not \U$19784 ( \20161 , \20160 );
not \U$19785 ( \20162 , \18706 );
or \U$19786 ( \20163 , \20161 , \20162 );
nand \U$19787 ( \20164 , \18693 , \18699 );
nand \U$19788 ( \20165 , \20163 , \20164 );
xor \U$19789 ( \20166 , \20159 , \20165 );
xor \U$19790 ( \20167 , \17814 , \17819 );
and \U$19791 ( \20168 , \20167 , \17825 );
and \U$19792 ( \20169 , \17814 , \17819 );
or \U$19793 ( \20170 , \20168 , \20169 );
xor \U$19794 ( \20171 , \20166 , \20170 );
xor \U$19795 ( \20172 , \20158 , \20171 );
not \U$19796 ( \20173 , \17921 );
nand \U$19797 ( \20174 , \20173 , \17927 );
not \U$19798 ( \20175 , \20174 );
not \U$19799 ( \20176 , \17933 );
or \U$19800 ( \20177 , \20175 , \20176 );
nand \U$19801 ( \20178 , \17926 , \17921 );
nand \U$19802 ( \20179 , \20177 , \20178 );
xor \U$19803 ( \20180 , \17772 , \17777 );
and \U$19804 ( \20181 , \20180 , \17783 );
and \U$19805 ( \20182 , \17772 , \17777 );
or \U$19806 ( \20183 , \20181 , \20182 );
xor \U$19807 ( \20184 , \20179 , \20183 );
xor \U$19808 ( \20185 , \17790 , \17795 );
and \U$19809 ( \20186 , \20185 , \17802 );
and \U$19810 ( \20187 , \17790 , \17795 );
or \U$19811 ( \20188 , \20186 , \20187 );
xor \U$19812 ( \20189 , \20184 , \20188 );
xor \U$19813 ( \20190 , \20172 , \20189 );
not \U$19814 ( \20191 , \17807 );
not \U$19815 ( \20192 , \17869 );
or \U$19816 ( \20193 , \20191 , \20192 );
not \U$19817 ( \20194 , \17866 );
not \U$19818 ( \20195 , \17804 );
or \U$19819 ( \20196 , \20194 , \20195 );
nand \U$19820 ( \20197 , \20196 , \17761 );
nand \U$19821 ( \20198 , \20193 , \20197 );
buf \U$19822 ( \20199 , \20198 );
xor \U$19823 ( \20200 , \20190 , \20199 );
xor \U$19824 ( \20201 , \14491 , \14500 );
xor \U$19825 ( \20202 , \20201 , \14512 );
not \U$19826 ( \20203 , \18687 );
not \U$19827 ( \20204 , \18682 );
or \U$19828 ( \20205 , \20203 , \20204 );
nand \U$19829 ( \20206 , \18663 , \18681 );
nand \U$19830 ( \20207 , \20205 , \20206 );
and \U$19831 ( \20208 , \20202 , \20207 );
not \U$19832 ( \20209 , \20202 );
not \U$19833 ( \20210 , \20207 );
and \U$19834 ( \20211 , \20209 , \20210 );
nor \U$19835 ( \20212 , \20208 , \20211 );
xor \U$19836 ( \20213 , \14728 , \14716 );
and \U$19837 ( \20214 , \20213 , \14740 );
not \U$19838 ( \20215 , \20213 );
not \U$19839 ( \20216 , \14740 );
and \U$19840 ( \20217 , \20215 , \20216 );
nor \U$19841 ( \20218 , \20214 , \20217 );
xor \U$19842 ( \20219 , \20212 , \20218 );
xnor \U$19843 ( \20220 , \18688 , \18723 );
not \U$19844 ( \20221 , \20220 );
not \U$19845 ( \20222 , \18707 );
or \U$19846 ( \20223 , \20221 , \20222 );
not \U$19847 ( \20224 , \18688 );
nand \U$19848 ( \20225 , \20224 , \18724 );
nand \U$19849 ( \20226 , \20223 , \20225 );
xor \U$19850 ( \20227 , \20219 , \20226 );
and \U$19851 ( \20228 , \14455 , \14443 );
not \U$19852 ( \20229 , \14455 );
and \U$19853 ( \20230 , \20229 , \14444 );
nor \U$19854 ( \20231 , \20228 , \20230 );
xnor \U$19855 ( \20232 , \20231 , \14468 );
xnor \U$19856 ( \20233 , \14387 , \14393 );
xor \U$19857 ( \20234 , \20232 , \20233 );
not \U$19858 ( \20235 , \17842 );
not \U$19859 ( \20236 , \17859 );
or \U$19860 ( \20237 , \20235 , \20236 );
nand \U$19861 ( \20238 , \17854 , \17849 );
nand \U$19862 ( \20239 , \20237 , \20238 );
not \U$19863 ( \20240 , \20239 );
xor \U$19864 ( \20241 , \20234 , \20240 );
xnor \U$19865 ( \20242 , \20227 , \20241 );
xnor \U$19866 ( \20243 , \20200 , \20242 );
xor \U$19867 ( \20244 , \20152 , \20243 );
not \U$19868 ( \20245 , \20244 );
xor \U$19869 ( \20246 , \18599 , \18839 );
and \U$19870 ( \20247 , \20246 , \18931 );
and \U$19871 ( \20248 , \18599 , \18839 );
or \U$19872 ( \20249 , \20247 , \20248 );
not \U$19873 ( \20250 , \20249 );
or \U$19874 ( \20251 , \20245 , \20250 );
or \U$19875 ( \20252 , \20249 , \20244 );
nand \U$19876 ( \20253 , \20251 , \20252 );
not \U$19877 ( \20254 , \20253 );
or \U$19878 ( \20255 , \20052 , \20254 );
or \U$19879 ( \20256 , \20253 , \20051 );
nand \U$19880 ( \20257 , \20255 , \20256 );
not \U$19881 ( \20258 , \18932 );
xor \U$19882 ( \20259 , \17950 , \19547 );
not \U$19883 ( \20260 , \20259 );
or \U$19884 ( \20261 , \20258 , \20260 );
not \U$19885 ( \20262 , \19548 );
nand \U$19886 ( \20263 , \20262 , \17950 );
nand \U$19887 ( \20264 , \20261 , \20263 );
nor \U$19888 ( \20265 , \20257 , \20264 );
not \U$19889 ( \20266 , \20265 );
xor \U$19890 ( \20267 , \12926 , \12932 );
xor \U$19891 ( \20268 , \20267 , \12943 );
xor \U$19892 ( \20269 , \12833 , \12835 );
xor \U$19893 ( \20270 , \20269 , \12915 );
xor \U$19894 ( \20271 , \20268 , \20270 );
nand \U$19895 ( \20272 , \14584 , \14583 );
not \U$19896 ( \20273 , \14526 );
not \U$19897 ( \20274 , \14552 );
and \U$19898 ( \20275 , \20273 , \20274 );
and \U$19899 ( \20276 , \14526 , \14552 );
nor \U$19900 ( \20277 , \20275 , \20276 );
xor \U$19901 ( \20278 , \20272 , \20277 );
not \U$19902 ( \20279 , \20278 );
not \U$19903 ( \20280 , \20279 );
not \U$19904 ( \20281 , \19994 );
not \U$19905 ( \20282 , \20001 );
or \U$19906 ( \20283 , \20281 , \20282 );
not \U$19907 ( \20284 , \19993 );
and \U$19908 ( \20285 , \12892 , \12881 );
not \U$19909 ( \20286 , \12892 );
and \U$19910 ( \20287 , \20286 , \12880 );
nor \U$19911 ( \20288 , \20285 , \20287 );
nand \U$19912 ( \20289 , \20284 , \20288 );
nand \U$19913 ( \20290 , \20283 , \20289 );
not \U$19914 ( \20291 , \20290 );
not \U$19915 ( \20292 , \20291 );
and \U$19916 ( \20293 , \20280 , \20292 );
not \U$19917 ( \20294 , \20278 );
not \U$19918 ( \20295 , \20291 );
or \U$19919 ( \20296 , \20294 , \20295 );
or \U$19920 ( \20297 , \20278 , \20291 );
nand \U$19921 ( \20298 , \20296 , \20297 );
not \U$19922 ( \20299 , \20070 );
not \U$19923 ( \20300 , \20076 );
not \U$19924 ( \20301 , \20300 );
or \U$19925 ( \20302 , \20299 , \20301 );
not \U$19926 ( \20303 , \20069 );
nand \U$19927 ( \20304 , \20303 , \20067 );
nand \U$19928 ( \20305 , \20302 , \20304 );
and \U$19929 ( \20306 , \20298 , \20305 );
nor \U$19930 ( \20307 , \20293 , \20306 );
xor \U$19931 ( \20308 , \20271 , \20307 );
not \U$19932 ( \20309 , \20308 );
not \U$19933 ( \20310 , \20309 );
xor \U$19934 ( \20311 , \14358 , \14351 );
xor \U$19935 ( \20312 , \20311 , \14354 );
not \U$19936 ( \20313 , \20312 );
xor \U$19937 ( \20314 , \14831 , \14823 );
xnor \U$19938 ( \20315 , \20314 , \14826 );
not \U$19939 ( \20316 , \20315 );
not \U$19940 ( \20317 , \20316 );
xor \U$19941 ( \20318 , \14850 , \14845 );
xnor \U$19942 ( \20319 , \20318 , \14842 );
not \U$19943 ( \20320 , \20319 );
not \U$19944 ( \20321 , \20320 );
or \U$19945 ( \20322 , \20317 , \20321 );
not \U$19946 ( \20323 , \20315 );
not \U$19947 ( \20324 , \20319 );
or \U$19948 ( \20325 , \20323 , \20324 );
not \U$19949 ( \20326 , \20011 );
not \U$19950 ( \20327 , \20006 );
or \U$19951 ( \20328 , \20326 , \20327 );
not \U$19952 ( \20329 , \19988 );
nand \U$19953 ( \20330 , \20329 , \20002 );
nand \U$19954 ( \20331 , \20328 , \20330 );
nand \U$19955 ( \20332 , \20325 , \20331 );
nand \U$19956 ( \20333 , \20322 , \20332 );
not \U$19957 ( \20334 , \20333 );
or \U$19958 ( \20335 , \20313 , \20334 );
or \U$19959 ( \20336 , \20333 , \20312 );
nand \U$19960 ( \20337 , \20335 , \20336 );
not \U$19961 ( \20338 , \20337 );
or \U$19962 ( \20339 , \20310 , \20338 );
or \U$19963 ( \20340 , \20309 , \20337 );
nand \U$19964 ( \20341 , \20339 , \20340 );
xor \U$19965 ( \20342 , \20331 , \20320 );
xor \U$19966 ( \20343 , \20342 , \20316 );
not \U$19967 ( \20344 , \20343 );
not \U$19968 ( \20345 , \20212 );
not \U$19969 ( \20346 , \20218 );
or \U$19970 ( \20347 , \20345 , \20346 );
nand \U$19971 ( \20348 , \20207 , \20202 );
nand \U$19972 ( \20349 , \20347 , \20348 );
xor \U$19973 ( \20350 , \14515 , \14517 );
xnor \U$19974 ( \20351 , \20350 , \14520 );
xor \U$19975 ( \20352 , \20349 , \20351 );
xor \U$19976 ( \20353 , \20232 , \20233 );
and \U$19977 ( \20354 , \20353 , \20240 );
and \U$19978 ( \20355 , \20232 , \20233 );
or \U$19979 ( \20356 , \20354 , \20355 );
xnor \U$19980 ( \20357 , \20352 , \20356 );
xor \U$19981 ( \20358 , \14593 , \14651 );
xor \U$19982 ( \20359 , \20358 , \14700 );
xor \U$19983 ( \20360 , \14746 , \14788 );
xnor \U$19984 ( \20361 , \20360 , \14743 );
xor \U$19985 ( \20362 , \20359 , \20361 );
not \U$19986 ( \20363 , \14476 );
nand \U$19987 ( \20364 , \20363 , \14473 );
buf \U$19988 ( \20365 , \14396 );
xnor \U$19989 ( \20366 , \20364 , \20365 );
xnor \U$19990 ( \20367 , \20362 , \20366 );
xnor \U$19991 ( \20368 , \20357 , \20367 );
not \U$19992 ( \20369 , \20368 );
or \U$19993 ( \20370 , \20344 , \20369 );
not \U$19994 ( \20371 , \20357 );
nand \U$19995 ( \20372 , \20371 , \20367 );
nand \U$19996 ( \20373 , \20370 , \20372 );
not \U$19997 ( \20374 , \20349 );
not \U$19998 ( \20375 , \20374 );
not \U$19999 ( \20376 , \20356 );
or \U$20000 ( \20377 , \20375 , \20376 );
not \U$20001 ( \20378 , \20351 );
nand \U$20002 ( \20379 , \20377 , \20378 );
not \U$20003 ( \20380 , \20356 );
not \U$20004 ( \20381 , \20374 );
nand \U$20005 ( \20382 , \20380 , \20381 );
nand \U$20006 ( \20383 , \20379 , \20382 );
buf \U$20007 ( \20384 , \20361 );
or \U$20008 ( \20385 , \20384 , \20359 );
nand \U$20009 ( \20386 , \20385 , \20366 );
nand \U$20010 ( \20387 , \20384 , \20359 );
and \U$20011 ( \20388 , \20386 , \20387 );
xor \U$20012 ( \20389 , \20383 , \20388 );
xor \U$20013 ( \20390 , \14833 , \14856 );
xor \U$20014 ( \20391 , \20389 , \20390 );
nor \U$20015 ( \20392 , \20373 , \20391 );
not \U$20016 ( \20393 , \20392 );
nand \U$20017 ( \20394 , \20373 , \20391 );
nand \U$20018 ( \20395 , \20393 , \20394 );
xnor \U$20019 ( \20396 , \20341 , \20395 );
not \U$20020 ( \20397 , \19979 );
not \U$20021 ( \20398 , \20024 );
or \U$20022 ( \20399 , \20397 , \20398 );
not \U$20023 ( \20400 , \20012 );
nand \U$20024 ( \20401 , \20400 , \20020 );
nand \U$20025 ( \20402 , \20399 , \20401 );
xor \U$20026 ( \20403 , \20158 , \20171 );
and \U$20027 ( \20404 , \20403 , \20189 );
and \U$20028 ( \20405 , \20158 , \20171 );
or \U$20029 ( \20406 , \20404 , \20405 );
not \U$20030 ( \20407 , \20406 );
not \U$20031 ( \20408 , \20098 );
nand \U$20032 ( \20409 , \20408 , \20092 );
nand \U$20033 ( \20410 , \20409 , \20090 );
not \U$20034 ( \20411 , \20305 );
not \U$20035 ( \20412 , \20298 );
not \U$20036 ( \20413 , \20412 );
or \U$20037 ( \20414 , \20411 , \20413 );
not \U$20038 ( \20415 , \20305 );
nand \U$20039 ( \20416 , \20415 , \20298 );
nand \U$20040 ( \20417 , \20414 , \20416 );
xor \U$20041 ( \20418 , \20410 , \20417 );
not \U$20042 ( \20419 , \20418 );
not \U$20043 ( \20420 , \20419 );
or \U$20044 ( \20421 , \20407 , \20420 );
not \U$20045 ( \20422 , \20406 );
nand \U$20046 ( \20423 , \20422 , \20418 );
nand \U$20047 ( \20424 , \20421 , \20423 );
xor \U$20048 ( \20425 , \20402 , \20424 );
not \U$20049 ( \20426 , \20140 );
not \U$20050 ( \20427 , \20109 );
or \U$20051 ( \20428 , \20426 , \20427 );
nand \U$20052 ( \20429 , \20105 , \20058 );
nand \U$20053 ( \20430 , \20428 , \20429 );
xor \U$20054 ( \20431 , \20425 , \20430 );
not \U$20055 ( \20432 , \20039 );
not \U$20056 ( \20433 , \20034 );
or \U$20057 ( \20434 , \20432 , \20433 );
not \U$20058 ( \20435 , \20032 );
nand \U$20059 ( \20436 , \20435 , \20025 );
nand \U$20060 ( \20437 , \20434 , \20436 );
nand \U$20061 ( \20438 , \20431 , \20437 );
not \U$20062 ( \20439 , \20438 );
not \U$20063 ( \20440 , \20141 );
not \U$20064 ( \20441 , \20440 );
not \U$20065 ( \20442 , \20243 );
not \U$20066 ( \20443 , \20442 );
or \U$20067 ( \20444 , \20441 , \20443 );
not \U$20068 ( \20445 , \20141 );
not \U$20069 ( \20446 , \20243 );
or \U$20070 ( \20447 , \20445 , \20446 );
nand \U$20071 ( \20448 , \20447 , \20148 );
nand \U$20072 ( \20449 , \20444 , \20448 );
not \U$20073 ( \20450 , \20449 );
not \U$20074 ( \20451 , \20450 );
or \U$20075 ( \20452 , \20439 , \20451 );
nor \U$20076 ( \20453 , \20431 , \20437 );
not \U$20077 ( \20454 , \20453 );
nand \U$20078 ( \20455 , \20452 , \20454 );
xor \U$20079 ( \20456 , \20396 , \20455 );
not \U$20080 ( \20457 , \20406 );
not \U$20081 ( \20458 , \20418 );
or \U$20082 ( \20459 , \20457 , \20458 );
nand \U$20083 ( \20460 , \20417 , \20410 );
nand \U$20084 ( \20461 , \20459 , \20460 );
xor \U$20085 ( \20462 , \20159 , \20165 );
and \U$20086 ( \20463 , \20462 , \20170 );
and \U$20087 ( \20464 , \20159 , \20165 );
or \U$20088 ( \20465 , \20463 , \20464 );
xor \U$20089 ( \20466 , \20179 , \20183 );
and \U$20090 ( \20467 , \20466 , \20188 );
and \U$20091 ( \20468 , \20179 , \20183 );
or \U$20092 ( \20469 , \20467 , \20468 );
xor \U$20093 ( \20470 , \20465 , \20469 );
xor \U$20094 ( \20471 , \20129 , \20131 );
and \U$20095 ( \20472 , \20471 , \20134 );
and \U$20096 ( \20473 , \20129 , \20131 );
or \U$20097 ( \20474 , \20472 , \20473 );
and \U$20098 ( \20475 , \20470 , \20474 );
and \U$20099 ( \20476 , \20465 , \20469 );
or \U$20100 ( \20477 , \20475 , \20476 );
xor \U$20101 ( \20478 , \14589 , \14703 );
xnor \U$20102 ( \20479 , \20478 , \14793 );
xor \U$20103 ( \20480 , \20477 , \20479 );
xor \U$20104 ( \20481 , \14365 , \14523 );
xor \U$20105 ( \20482 , \20481 , \14479 );
xor \U$20106 ( \20483 , \20480 , \20482 );
xor \U$20107 ( \20484 , \20461 , \20483 );
not \U$20108 ( \20485 , \20115 );
not \U$20109 ( \20486 , \20124 );
or \U$20110 ( \20487 , \20485 , \20486 );
or \U$20111 ( \20488 , \20115 , \20124 );
nand \U$20112 ( \20489 , \20488 , \20135 );
nand \U$20113 ( \20490 , \20487 , \20489 );
xor \U$20114 ( \20491 , \20465 , \20469 );
xor \U$20115 ( \20492 , \20491 , \20474 );
nand \U$20116 ( \20493 , \20490 , \20492 );
not \U$20117 ( \20494 , \20219 );
not \U$20118 ( \20495 , \20494 );
not \U$20119 ( \20496 , \20241 );
or \U$20120 ( \20497 , \20495 , \20496 );
nand \U$20121 ( \20498 , \20497 , \20226 );
or \U$20122 ( \20499 , \20241 , \20494 );
and \U$20123 ( \20500 , \20493 , \20498 , \20499 );
nor \U$20124 ( \20501 , \20490 , \20492 );
nor \U$20125 ( \20502 , \20500 , \20501 );
xor \U$20126 ( \20503 , \20484 , \20502 );
not \U$20127 ( \20504 , \20503 );
xor \U$20128 ( \20505 , \20402 , \20424 );
and \U$20129 ( \20506 , \20505 , \20430 );
and \U$20130 ( \20507 , \20402 , \20424 );
or \U$20131 ( \20508 , \20506 , \20507 );
not \U$20132 ( \20509 , \20508 );
nand \U$20133 ( \20510 , \20504 , \20509 );
nand \U$20134 ( \20511 , \20503 , \20508 );
nand \U$20135 ( \20512 , \20510 , \20511 );
and \U$20136 ( \20513 , \20368 , \20343 );
not \U$20137 ( \20514 , \20368 );
not \U$20138 ( \20515 , \20343 );
and \U$20139 ( \20516 , \20514 , \20515 );
nor \U$20140 ( \20517 , \20513 , \20516 );
not \U$20141 ( \20518 , \20517 );
not \U$20142 ( \20519 , \20190 );
not \U$20143 ( \20520 , \20199 );
or \U$20144 ( \20521 , \20519 , \20520 );
not \U$20145 ( \20522 , \20198 );
not \U$20146 ( \20523 , \20190 );
nand \U$20147 ( \20524 , \20522 , \20523 );
nand \U$20148 ( \20525 , \20242 , \20524 );
nand \U$20149 ( \20526 , \20521 , \20525 );
not \U$20150 ( \20527 , \20526 );
nand \U$20151 ( \20528 , \20498 , \20499 );
not \U$20152 ( \20529 , \20528 );
not \U$20153 ( \20530 , \20501 );
nand \U$20154 ( \20531 , \20530 , \20493 );
not \U$20155 ( \20532 , \20531 );
and \U$20156 ( \20533 , \20529 , \20532 );
and \U$20157 ( \20534 , \20528 , \20531 );
nor \U$20158 ( \20535 , \20533 , \20534 );
not \U$20159 ( \20536 , \20535 );
or \U$20160 ( \20537 , \20527 , \20536 );
or \U$20161 ( \20538 , \20535 , \20526 );
nand \U$20162 ( \20539 , \20537 , \20538 );
not \U$20163 ( \20540 , \20539 );
or \U$20164 ( \20541 , \20518 , \20540 );
not \U$20165 ( \20542 , \20535 );
nand \U$20166 ( \20543 , \20542 , \20526 );
nand \U$20167 ( \20544 , \20541 , \20543 );
xor \U$20168 ( \20545 , \20512 , \20544 );
xor \U$20169 ( \20546 , \20456 , \20545 );
not \U$20170 ( \20547 , \20449 );
not \U$20171 ( \20548 , \20453 );
nand \U$20172 ( \20549 , \20548 , \20438 );
not \U$20173 ( \20550 , \20549 );
or \U$20174 ( \20551 , \20547 , \20550 );
or \U$20175 ( \20552 , \20549 , \20449 );
nand \U$20176 ( \20553 , \20551 , \20552 );
not \U$20177 ( \20554 , \20553 );
not \U$20178 ( \20555 , \20045 );
not \U$20179 ( \20556 , \19975 );
or \U$20180 ( \20557 , \20555 , \20556 );
not \U$20181 ( \20558 , \19975 );
not \U$20182 ( \20559 , \20558 );
not \U$20183 ( \20560 , \20044 );
or \U$20184 ( \20561 , \20559 , \20560 );
nand \U$20185 ( \20562 , \20561 , \20050 );
nand \U$20186 ( \20563 , \20557 , \20562 );
xor \U$20187 ( \20564 , \20517 , \20539 );
nand \U$20188 ( \20565 , \20563 , \20564 );
nand \U$20189 ( \20566 , \20554 , \20565 );
or \U$20190 ( \20567 , \20563 , \20564 );
nand \U$20191 ( \20568 , \20566 , \20567 );
nand \U$20192 ( \20569 , \20546 , \20568 );
not \U$20193 ( \20570 , \20553 );
not \U$20194 ( \20571 , \20564 );
not \U$20195 ( \20572 , \20563 );
or \U$20196 ( \20573 , \20571 , \20572 );
or \U$20197 ( \20574 , \20564 , \20563 );
nand \U$20198 ( \20575 , \20573 , \20574 );
not \U$20199 ( \20576 , \20575 );
or \U$20200 ( \20577 , \20570 , \20576 );
or \U$20201 ( \20578 , \20553 , \20575 );
nand \U$20202 ( \20579 , \20577 , \20578 );
not \U$20203 ( \20580 , \20051 );
not \U$20204 ( \20581 , \20580 );
not \U$20205 ( \20582 , \20253 );
or \U$20206 ( \20583 , \20581 , \20582 );
not \U$20207 ( \20584 , \20244 );
nand \U$20208 ( \20585 , \20584 , \20249 );
nand \U$20209 ( \20586 , \20583 , \20585 );
nor \U$20210 ( \20587 , \20579 , \20586 );
not \U$20211 ( \20588 , \20587 );
and \U$20212 ( \20589 , \19971 , \20266 , \20569 , \20588 );
xor \U$20213 ( \20590 , \14339 , \14879 );
xor \U$20214 ( \20591 , \20590 , \14347 );
xor \U$20215 ( \20592 , \14312 , \14271 );
xor \U$20216 ( \20593 , \20592 , \14315 );
not \U$20217 ( \20594 , \20593 );
not \U$20218 ( \20595 , \20594 );
xor \U$20219 ( \20596 , \20268 , \20270 );
and \U$20220 ( \20597 , \20596 , \20307 );
and \U$20221 ( \20598 , \20268 , \20270 );
or \U$20222 ( \20599 , \20597 , \20598 );
not \U$20223 ( \20600 , \20599 );
or \U$20224 ( \20601 , \20595 , \20600 );
not \U$20225 ( \20602 , \14234 );
not \U$20226 ( \20603 , \14226 );
or \U$20227 ( \20604 , \20602 , \20603 );
or \U$20228 ( \20605 , \14234 , \14226 );
nand \U$20229 ( \20606 , \20604 , \20605 );
not \U$20230 ( \20607 , \14239 );
and \U$20231 ( \20608 , \20606 , \20607 );
not \U$20232 ( \20609 , \20606 );
and \U$20233 ( \20610 , \20609 , \14239 );
nor \U$20234 ( \20611 , \20608 , \20610 );
not \U$20235 ( \20612 , \20611 );
nand \U$20236 ( \20613 , \20601 , \20612 );
not \U$20237 ( \20614 , \20599 );
nand \U$20238 ( \20615 , \20614 , \20593 );
nand \U$20239 ( \20616 , \20613 , \20615 );
not \U$20240 ( \20617 , \20616 );
not \U$20241 ( \20618 , \14266 );
and \U$20242 ( \20619 , \14325 , \20618 );
not \U$20243 ( \20620 , \14325 );
and \U$20244 ( \20621 , \20620 , \14266 );
nor \U$20245 ( \20622 , \20619 , \20621 );
nand \U$20246 ( \20623 , \20617 , \20622 );
not \U$20247 ( \20624 , \14260 );
not \U$20248 ( \20625 , \14243 );
not \U$20249 ( \20626 , \20625 );
or \U$20250 ( \20627 , \20624 , \20626 );
nand \U$20251 ( \20628 , \14243 , \14259 );
nand \U$20252 ( \20629 , \20627 , \20628 );
not \U$20253 ( \20630 , \14246 );
and \U$20254 ( \20631 , \20629 , \20630 );
not \U$20255 ( \20632 , \20629 );
and \U$20256 ( \20633 , \20632 , \14246 );
nor \U$20257 ( \20634 , \20631 , \20633 );
not \U$20258 ( \20635 , \20634 );
and \U$20259 ( \20636 , \20623 , \20635 );
not \U$20260 ( \20637 , \20616 );
nor \U$20261 ( \20638 , \20637 , \20622 );
nor \U$20262 ( \20639 , \20636 , \20638 );
xor \U$20263 ( \20640 , \20477 , \20479 );
and \U$20264 ( \20641 , \20640 , \20482 );
and \U$20265 ( \20642 , \20477 , \20479 );
or \U$20266 ( \20643 , \20641 , \20642 );
not \U$20267 ( \20644 , \14798 );
xor \U$20268 ( \20645 , \14525 , \20644 );
xnor \U$20269 ( \20646 , \20645 , \14362 );
xor \U$20270 ( \20647 , \20643 , \20646 );
xor \U$20271 ( \20648 , \20383 , \20388 );
and \U$20272 ( \20649 , \20648 , \20390 );
and \U$20273 ( \20650 , \20383 , \20388 );
or \U$20274 ( \20651 , \20649 , \20650 );
and \U$20275 ( \20652 , \20647 , \20651 );
and \U$20276 ( \20653 , \20643 , \20646 );
or \U$20277 ( \20654 , \20652 , \20653 );
xor \U$20278 ( \20655 , \14803 , \14806 );
xor \U$20279 ( \20656 , \20655 , \14867 );
xor \U$20280 ( \20657 , \20654 , \20656 );
not \U$20281 ( \20658 , \20312 );
nand \U$20282 ( \20659 , \20658 , \20309 );
not \U$20283 ( \20660 , \20312 );
not \U$20284 ( \20661 , \20308 );
or \U$20285 ( \20662 , \20660 , \20661 );
nand \U$20286 ( \20663 , \20662 , \20333 );
nand \U$20287 ( \20664 , \20659 , \20663 );
and \U$20288 ( \20665 , \20611 , \20593 );
not \U$20289 ( \20666 , \20611 );
and \U$20290 ( \20667 , \20666 , \20594 );
or \U$20291 ( \20668 , \20665 , \20667 );
buf \U$20292 ( \20669 , \20599 );
not \U$20293 ( \20670 , \20669 );
and \U$20294 ( \20671 , \20668 , \20670 );
not \U$20295 ( \20672 , \20668 );
and \U$20296 ( \20673 , \20672 , \20669 );
nor \U$20297 ( \20674 , \20671 , \20673 );
xor \U$20298 ( \20675 , \20664 , \20674 );
xor \U$20299 ( \20676 , \14821 , \14818 );
xnor \U$20300 ( \20677 , \20676 , \14861 );
and \U$20301 ( \20678 , \20675 , \20677 );
and \U$20302 ( \20679 , \20664 , \20674 );
or \U$20303 ( \20680 , \20678 , \20679 );
and \U$20304 ( \20681 , \20657 , \20680 );
and \U$20305 ( \20682 , \20654 , \20656 );
or \U$20306 ( \20683 , \20681 , \20682 );
not \U$20307 ( \20684 , \20683 );
xor \U$20308 ( \20685 , \20639 , \20684 );
xor \U$20309 ( \20686 , \14871 , \14869 );
xnor \U$20310 ( \20687 , \20686 , \14875 );
and \U$20311 ( \20688 , \20685 , \20687 );
and \U$20312 ( \20689 , \20639 , \20684 );
or \U$20313 ( \20690 , \20688 , \20689 );
nand \U$20314 ( \20691 , \20591 , \20690 );
xor \U$20315 ( \20692 , \20461 , \20483 );
and \U$20316 ( \20693 , \20692 , \20502 );
and \U$20317 ( \20694 , \20461 , \20483 );
or \U$20318 ( \20695 , \20693 , \20694 );
not \U$20319 ( \20696 , \20695 );
not \U$20320 ( \20697 , \20696 );
xor \U$20321 ( \20698 , \20643 , \20646 );
xor \U$20322 ( \20699 , \20698 , \20651 );
not \U$20323 ( \20700 , \20699 );
or \U$20324 ( \20701 , \20697 , \20700 );
not \U$20325 ( \20702 , \20699 );
nand \U$20326 ( \20703 , \20702 , \20695 );
nand \U$20327 ( \20704 , \20701 , \20703 );
or \U$20328 ( \20705 , \20341 , \20392 );
nand \U$20329 ( \20706 , \20705 , \20394 );
buf \U$20330 ( \20707 , \20706 );
xor \U$20331 ( \20708 , \20704 , \20707 );
not \U$20332 ( \20709 , \20708 );
not \U$20333 ( \20710 , \20511 );
or \U$20334 ( \20711 , \20544 , \20710 );
nand \U$20335 ( \20712 , \20711 , \20510 );
not \U$20336 ( \20713 , \20712 );
xor \U$20337 ( \20714 , \20664 , \20674 );
xor \U$20338 ( \20715 , \20714 , \20677 );
not \U$20339 ( \20716 , \20715 );
or \U$20340 ( \20717 , \20713 , \20716 );
or \U$20341 ( \20718 , \20715 , \20712 );
nand \U$20342 ( \20719 , \20717 , \20718 );
not \U$20343 ( \20720 , \20719 );
or \U$20344 ( \20721 , \20709 , \20720 );
or \U$20345 ( \20722 , \20708 , \20719 );
nand \U$20346 ( \20723 , \20721 , \20722 );
xor \U$20347 ( \20724 , \20396 , \20455 );
and \U$20348 ( \20725 , \20724 , \20545 );
and \U$20349 ( \20726 , \20396 , \20455 );
or \U$20350 ( \20727 , \20725 , \20726 );
nand \U$20351 ( \20728 , \20723 , \20727 );
xor \U$20352 ( \20729 , \20654 , \20656 );
xor \U$20353 ( \20730 , \20729 , \20680 );
xnor \U$20354 ( \20731 , \20616 , \20634 );
not \U$20355 ( \20732 , \20731 );
not \U$20356 ( \20733 , \20622 );
or \U$20357 ( \20734 , \20732 , \20733 );
or \U$20358 ( \20735 , \20731 , \20622 );
nand \U$20359 ( \20736 , \20734 , \20735 );
not \U$20360 ( \20737 , \20736 );
not \U$20361 ( \20738 , \20702 );
not \U$20362 ( \20739 , \20696 );
or \U$20363 ( \20740 , \20738 , \20739 );
not \U$20364 ( \20741 , \20695 );
not \U$20365 ( \20742 , \20699 );
or \U$20366 ( \20743 , \20741 , \20742 );
not \U$20367 ( \20744 , \20706 );
nand \U$20368 ( \20745 , \20743 , \20744 );
nand \U$20369 ( \20746 , \20740 , \20745 );
not \U$20370 ( \20747 , \20746 );
or \U$20371 ( \20748 , \20737 , \20747 );
or \U$20372 ( \20749 , \20746 , \20736 );
nand \U$20373 ( \20750 , \20748 , \20749 );
xnor \U$20374 ( \20751 , \20730 , \20750 );
not \U$20375 ( \20752 , \20708 );
not \U$20376 ( \20753 , \20752 );
not \U$20377 ( \20754 , \20719 );
or \U$20378 ( \20755 , \20753 , \20754 );
not \U$20379 ( \20756 , \20715 );
nand \U$20380 ( \20757 , \20756 , \20712 );
nand \U$20381 ( \20758 , \20755 , \20757 );
nand \U$20382 ( \20759 , \20751 , \20758 );
nand \U$20383 ( \20760 , \20728 , \20759 );
not \U$20384 ( \20761 , \20760 );
xor \U$20385 ( \20762 , \20639 , \20684 );
xor \U$20386 ( \20763 , \20762 , \20687 );
not \U$20387 ( \20764 , \20750 );
not \U$20388 ( \20765 , \20730 );
not \U$20389 ( \20766 , \20765 );
or \U$20390 ( \20767 , \20764 , \20766 );
not \U$20391 ( \20768 , \20736 );
nand \U$20392 ( \20769 , \20768 , \20746 );
nand \U$20393 ( \20770 , \20767 , \20769 );
nand \U$20394 ( \20771 , \20763 , \20770 );
and \U$20395 ( \20772 , \20589 , \20691 , \20761 , \20771 );
not \U$20396 ( \20773 , \15557 );
not \U$20397 ( \20774 , \20773 );
not \U$20398 ( \20775 , \15620 );
not \U$20399 ( \20776 , \20775 );
or \U$20400 ( \20777 , \20774 , \20776 );
nand \U$20401 ( \20778 , \20777 , \15904 );
nand \U$20402 ( \20779 , \15620 , \15557 );
nand \U$20403 ( \20780 , \20778 , \20779 );
not \U$20404 ( \20781 , \20780 );
xor \U$20405 ( \20782 , \15162 , \15277 );
and \U$20406 ( \20783 , \20782 , \15556 );
and \U$20407 ( \20784 , \15162 , \15277 );
or \U$20408 ( \20785 , \20783 , \20784 );
xor \U$20409 ( \20786 , \15198 , \15202 );
and \U$20410 ( \20787 , \20786 , \15237 );
and \U$20411 ( \20788 , \15198 , \15202 );
or \U$20412 ( \20789 , \20787 , \20788 );
not \U$20413 ( \20790 , \15282 );
not \U$20414 ( \20791 , \15304 );
or \U$20415 ( \20792 , \20790 , \20791 );
not \U$20416 ( \20793 , \15282 );
not \U$20417 ( \20794 , \20793 );
not \U$20418 ( \20795 , \15301 );
or \U$20419 ( \20796 , \20794 , \20795 );
nand \U$20420 ( \20797 , \20796 , \15286 );
nand \U$20421 ( \20798 , \20792 , \20797 );
xor \U$20422 ( \20799 , \20789 , \20798 );
not \U$20423 ( \20800 , \15545 );
not \U$20424 ( \20801 , \15540 );
or \U$20425 ( \20802 , \20800 , \20801 );
not \U$20426 ( \20803 , \15536 );
nand \U$20427 ( \20804 , \20803 , \15510 );
nand \U$20428 ( \20805 , \20802 , \20804 );
xor \U$20429 ( \20806 , \20799 , \20805 );
not \U$20430 ( \20807 , \15465 );
not \U$20431 ( \20808 , \20807 );
not \U$20432 ( \20809 , \15547 );
or \U$20433 ( \20810 , \20808 , \20809 );
not \U$20434 ( \20811 , \15546 );
not \U$20435 ( \20812 , \15465 );
or \U$20436 ( \20813 , \20811 , \20812 );
nand \U$20437 ( \20814 , \20813 , \15472 );
nand \U$20438 ( \20815 , \20810 , \20814 );
xor \U$20439 ( \20816 , \20806 , \20815 );
xor \U$20440 ( \20817 , \15189 , \15193 );
and \U$20441 ( \20818 , \20817 , \15238 );
and \U$20442 ( \20819 , \15189 , \15193 );
or \U$20443 ( \20820 , \20818 , \20819 );
xor \U$20444 ( \20821 , \20816 , \20820 );
not \U$20445 ( \20822 , \15306 );
not \U$20446 ( \20823 , \20822 );
not \U$20447 ( \20824 , \15422 );
not \U$20448 ( \20825 , \20824 );
or \U$20449 ( \20826 , \20823 , \20825 );
not \U$20450 ( \20827 , \15422 );
not \U$20451 ( \20828 , \15306 );
or \U$20452 ( \20829 , \20827 , \20828 );
nand \U$20453 ( \20830 , \20829 , \15315 );
nand \U$20454 ( \20831 , \20826 , \20830 );
not \U$20455 ( \20832 , \15328 );
or \U$20456 ( \20833 , \15339 , \15350 );
not \U$20457 ( \20834 , \20833 );
or \U$20458 ( \20835 , \20832 , \20834 );
nand \U$20459 ( \20836 , \15350 , \15339 );
nand \U$20460 ( \20837 , \20835 , \20836 );
not \U$20461 ( \20838 , \15508 );
not \U$20462 ( \20839 , \15496 );
or \U$20463 ( \20840 , \20838 , \20839 );
nand \U$20464 ( \20841 , \15509 , \15486 );
nand \U$20465 ( \20842 , \20840 , \20841 );
xnor \U$20466 ( \20843 , \20837 , \20842 );
xor \U$20467 ( \20844 , \15370 , \15380 );
and \U$20468 ( \20845 , \20844 , \15391 );
and \U$20469 ( \20846 , \15370 , \15380 );
or \U$20470 ( \20847 , \20845 , \20846 );
not \U$20471 ( \20848 , \20847 );
and \U$20472 ( \20849 , \20843 , \20848 );
not \U$20473 ( \20850 , \20843 );
and \U$20474 ( \20851 , \20850 , \20847 );
nor \U$20475 ( \20852 , \20849 , \20851 );
xor \U$20476 ( \20853 , \15356 , \15392 );
and \U$20477 ( \20854 , \20853 , \15421 );
and \U$20478 ( \20855 , \15356 , \15392 );
or \U$20479 ( \20856 , \20854 , \20855 );
xor \U$20480 ( \20857 , \20852 , \20856 );
not \U$20481 ( \20858 , \1864 );
not \U$20482 ( \20859 , \6256 );
not \U$20483 ( \20860 , RIae793b8_143);
and \U$20484 ( \20861 , \20859 , \20860 );
and \U$20485 ( \20862 , \5109 , RIae793b8_143);
nor \U$20486 ( \20863 , \20861 , \20862 );
not \U$20487 ( \20864 , \20863 );
or \U$20488 ( \20865 , \20858 , \20864 );
nand \U$20489 ( \20866 , \15211 , \1910 );
nand \U$20490 ( \20867 , \20865 , \20866 );
not \U$20491 ( \20868 , \1499 );
not \U$20492 ( \20869 , \15222 );
or \U$20493 ( \20870 , \20868 , \20869 );
and \U$20494 ( \20871 , RIae79250_140, \15117 );
not \U$20495 ( \20872 , RIae79250_140);
and \U$20496 ( \20873 , \20872 , \14631 );
or \U$20497 ( \20874 , \20871 , \20873 );
nand \U$20498 ( \20875 , \20874 , \1501 );
nand \U$20499 ( \20876 , \20870 , \20875 );
xor \U$20500 ( \20877 , \20867 , \20876 );
not \U$20501 ( \20878 , \1008 );
not \U$20502 ( \20879 , \15524 );
or \U$20503 ( \20880 , \20878 , \20879 );
not \U$20504 ( \20881 , RIae79160_138);
not \U$20505 ( \20882 , \9313 );
or \U$20506 ( \20883 , \20881 , \20882 );
nand \U$20507 ( \20884 , \10386 , \6414 );
nand \U$20508 ( \20885 , \20883 , \20884 );
nand \U$20509 ( \20886 , \20885 , \10451 );
nand \U$20510 ( \20887 , \20880 , \20886 );
xnor \U$20511 ( \20888 , \20877 , \20887 );
not \U$20512 ( \20889 , \20888 );
not \U$20513 ( \20890 , \20889 );
not \U$20514 ( \20891 , \1844 );
not \U$20515 ( \20892 , \15828 );
or \U$20516 ( \20893 , \20891 , \20892 );
and \U$20517 ( \20894 , \2403 , \2970 );
not \U$20518 ( \20895 , \2403 );
and \U$20519 ( \20896 , \20895 , RIae79688_149);
nor \U$20520 ( \20897 , \20894 , \20896 );
nand \U$20521 ( \20898 , \20897 , \1821 );
nand \U$20522 ( \20899 , \20893 , \20898 );
not \U$20523 ( \20900 , \20899 );
not \U$20524 ( \20901 , \20900 );
nand \U$20525 ( \20902 , \13544 , RIae78b48_125);
not \U$20526 ( \20903 , \20902 );
not \U$20527 ( \20904 , \2011 );
and \U$20528 ( \20905 , RIae79610_148, \6242 );
not \U$20529 ( \20906 , RIae79610_148);
and \U$20530 ( \20907 , \20906 , \4927 );
or \U$20531 ( \20908 , \20905 , \20907 );
not \U$20532 ( \20909 , \20908 );
or \U$20533 ( \20910 , \20904 , \20909 );
nand \U$20534 ( \20911 , \15232 , \9370 );
nand \U$20535 ( \20912 , \20910 , \20911 );
not \U$20536 ( \20913 , \20912 );
or \U$20537 ( \20914 , \20903 , \20913 );
or \U$20538 ( \20915 , \20912 , \20902 );
nand \U$20539 ( \20916 , \20914 , \20915 );
not \U$20540 ( \20917 , \20916 );
or \U$20541 ( \20918 , \20901 , \20917 );
or \U$20542 ( \20919 , \20916 , \20900 );
nand \U$20543 ( \20920 , \20918 , \20919 );
not \U$20544 ( \20921 , \20920 );
not \U$20545 ( \20922 , \20921 );
or \U$20546 ( \20923 , \20890 , \20922 );
nand \U$20547 ( \20924 , \20920 , \20888 );
nand \U$20548 ( \20925 , \20923 , \20924 );
not \U$20549 ( \20926 , \15631 );
not \U$20550 ( \20927 , \15662 );
or \U$20551 ( \20928 , \20926 , \20927 );
nand \U$20552 ( \20929 , \15640 , \15660 );
nand \U$20553 ( \20930 , \20928 , \20929 );
xor \U$20554 ( \20931 , \20925 , \20930 );
xnor \U$20555 ( \20932 , \20857 , \20931 );
xor \U$20556 ( \20933 , \20831 , \20932 );
xor \U$20557 ( \20934 , RIae78e90_132, \15944 );
not \U$20558 ( \20935 , \20934 );
not \U$20559 ( \20936 , \1073 );
and \U$20560 ( \20937 , \20935 , \20936 );
and \U$20561 ( \20938 , \15498 , \1086 );
nor \U$20562 ( \20939 , \20937 , \20938 );
not \U$20563 ( \20940 , \1062 );
not \U$20564 ( \20941 , \9438 );
and \U$20565 ( \20942 , RIae79070_136, \20941 );
not \U$20566 ( \20943 , RIae79070_136);
and \U$20567 ( \20944 , \20943 , \9438 );
or \U$20568 ( \20945 , \20942 , \20944 );
not \U$20569 ( \20946 , \20945 );
or \U$20570 ( \20947 , \20940 , \20946 );
and \U$20571 ( \20948 , RIae79070_136, \9364 );
not \U$20572 ( \20949 , RIae79070_136);
and \U$20573 ( \20950 , \20949 , \9367 );
or \U$20574 ( \20951 , \20948 , \20950 );
nand \U$20575 ( \20952 , \20951 , \1049 );
nand \U$20576 ( \20953 , \20947 , \20952 );
xor \U$20577 ( \20954 , \20939 , \20953 );
not \U$20578 ( \20955 , \797 );
not \U$20579 ( \20956 , \15492 );
or \U$20580 ( \20957 , \20955 , \20956 );
and \U$20581 ( \20958 , RIae78f80_134, \14657 );
not \U$20582 ( \20959 , RIae78f80_134);
and \U$20583 ( \20960 , \20959 , \9455 );
or \U$20584 ( \20961 , \20958 , \20960 );
nand \U$20585 ( \20962 , \20961 , \838 );
nand \U$20586 ( \20963 , \20957 , \20962 );
xnor \U$20587 ( \20964 , \20954 , \20963 );
xor \U$20588 ( \20965 , \15670 , \15683 );
and \U$20589 ( \20966 , \20965 , \15690 );
and \U$20590 ( \20967 , \15670 , \15683 );
or \U$20591 ( \20968 , \20966 , \20967 );
xor \U$20592 ( \20969 , \20964 , \20968 );
nor \U$20593 ( \20970 , \15403 , \15420 );
or \U$20594 ( \20971 , \20970 , \15412 );
nand \U$20595 ( \20972 , \15403 , \15420 );
nand \U$20596 ( \20973 , \20971 , \20972 );
xor \U$20597 ( \20974 , \20969 , \20973 );
xor \U$20598 ( \20975 , \15663 , \15691 );
and \U$20599 ( \20976 , \20975 , \15715 );
and \U$20600 ( \20977 , \15663 , \15691 );
or \U$20601 ( \20978 , \20976 , \20977 );
xor \U$20602 ( \20979 , \20974 , \20978 );
not \U$20603 ( \20980 , \15810 );
not \U$20604 ( \20981 , \15806 );
not \U$20605 ( \20982 , \20981 );
not \U$20606 ( \20983 , \15833 );
or \U$20607 ( \20984 , \20982 , \20983 );
or \U$20608 ( \20985 , \15833 , \20981 );
nand \U$20609 ( \20986 , \20984 , \20985 );
not \U$20610 ( \20987 , \20986 );
or \U$20611 ( \20988 , \20980 , \20987 );
not \U$20612 ( \20989 , \20981 );
nand \U$20613 ( \20990 , \20989 , \15833 );
nand \U$20614 ( \20991 , \20988 , \20990 );
not \U$20615 ( \20992 , \5048 );
and \U$20616 ( \20993 , RIae79d90_164, \2047 );
not \U$20617 ( \20994 , RIae79d90_164);
and \U$20618 ( \20995 , \20994 , \2048 );
or \U$20619 ( \20996 , \20993 , \20995 );
not \U$20620 ( \20997 , \20996 );
or \U$20621 ( \20998 , \20992 , \20997 );
nand \U$20622 ( \20999 , \15666 , \5040 );
nand \U$20623 ( \21000 , \20998 , \20999 );
not \U$20624 ( \21001 , \11014 );
not \U$20625 ( \21002 , \15679 );
or \U$20626 ( \21003 , \21001 , \21002 );
and \U$20627 ( \21004 , RIae7a3a8_177, \3326 );
not \U$20628 ( \21005 , RIae7a3a8_177);
and \U$20629 ( \21006 , \21005 , \1289 );
or \U$20630 ( \21007 , \21004 , \21006 );
nand \U$20631 ( \21008 , \21007 , \9622 );
nand \U$20632 ( \21009 , \21003 , \21008 );
xor \U$20633 ( \21010 , \21000 , \21009 );
not \U$20634 ( \21011 , \12371 );
not \U$20635 ( \21012 , \11427 );
not \U$20636 ( \21013 , \991 );
or \U$20637 ( \21014 , \21012 , \21013 );
or \U$20638 ( \21015 , \991 , \10625 );
nand \U$20639 ( \21016 , \21014 , \21015 );
not \U$20640 ( \21017 , \21016 );
or \U$20641 ( \21018 , \21011 , \21017 );
nand \U$20642 ( \21019 , \10696 , \15389 );
nand \U$20643 ( \21020 , \21018 , \21019 );
xor \U$20644 ( \21021 , \21010 , \21020 );
not \U$20645 ( \21022 , \21021 );
not \U$20646 ( \21023 , \15346 );
not \U$20647 ( \21024 , \1988 );
or \U$20648 ( \21025 , \21023 , \21024 );
not \U$20649 ( \21026 , RIae797f0_152);
not \U$20650 ( \21027 , \2287 );
or \U$20651 ( \21028 , \21026 , \21027 );
or \U$20652 ( \21029 , \2287 , RIae797f0_152);
nand \U$20653 ( \21030 , \21028 , \21029 );
nand \U$20654 ( \21031 , \21030 , \2007 );
nand \U$20655 ( \21032 , \21025 , \21031 );
not \U$20656 ( \21033 , \14580 );
not \U$20657 ( \21034 , \15636 );
or \U$20658 ( \21035 , \21033 , \21034 );
not \U$20659 ( \21036 , RIae798e0_154);
not \U$20660 ( \21037 , \21036 );
not \U$20661 ( \21038 , \1759 );
or \U$20662 ( \21039 , \21037 , \21038 );
nand \U$20663 ( \21040 , \10905 , RIae798e0_154);
nand \U$20664 ( \21041 , \21039 , \21040 );
nand \U$20665 ( \21042 , \21041 , \2322 );
nand \U$20666 ( \21043 , \21035 , \21042 );
and \U$20667 ( \21044 , \21032 , \21043 );
not \U$20668 ( \21045 , \21032 );
not \U$20669 ( \21046 , \21043 );
and \U$20670 ( \21047 , \21045 , \21046 );
nor \U$20671 ( \21048 , \21044 , \21047 );
not \U$20672 ( \21049 , \21048 );
not \U$20673 ( \21050 , \10709 );
not \U$20674 ( \21051 , \15627 );
or \U$20675 ( \21052 , \21050 , \21051 );
not \U$20676 ( \21053 , RIae79fe8_169);
not \U$20677 ( \21054 , \5081 );
or \U$20678 ( \21055 , \21053 , \21054 );
nand \U$20679 ( \21056 , \1124 , \18027 );
nand \U$20680 ( \21057 , \21055 , \21056 );
nand \U$20681 ( \21058 , \21057 , \9517 );
nand \U$20682 ( \21059 , \21052 , \21058 );
not \U$20683 ( \21060 , \21059 );
not \U$20684 ( \21061 , \21060 );
and \U$20685 ( \21062 , \21049 , \21061 );
and \U$20686 ( \21063 , \21048 , \21060 );
nor \U$20687 ( \21064 , \21062 , \21063 );
not \U$20688 ( \21065 , \21064 );
or \U$20689 ( \21066 , \21022 , \21065 );
or \U$20690 ( \21067 , \21021 , \21064 );
nand \U$20691 ( \21068 , \21066 , \21067 );
xor \U$20692 ( \21069 , \20991 , \21068 );
xor \U$20693 ( \21070 , \20979 , \21069 );
buf \U$20694 ( \21071 , \21070 );
xor \U$20695 ( \21072 , \20933 , \21071 );
xor \U$20696 ( \21073 , \20821 , \21072 );
not \U$20697 ( \21074 , \15423 );
not \U$20698 ( \21075 , \21074 );
not \U$20699 ( \21076 , \15552 );
or \U$20700 ( \21077 , \21075 , \21076 );
not \U$20701 ( \21078 , \15548 );
nand \U$20702 ( \21079 , \21078 , \15429 );
nand \U$20703 ( \21080 , \21077 , \21079 );
xor \U$20704 ( \21081 , \21073 , \21080 );
xor \U$20705 ( \21082 , \20785 , \21081 );
xor \U$20706 ( \21083 , \15837 , \15843 );
and \U$20707 ( \21084 , \21083 , \15870 );
and \U$20708 ( \21085 , \15837 , \15843 );
or \U$20709 ( \21086 , \21084 , \21085 );
not \U$20710 ( \21087 , \21086 );
xor \U$20711 ( \21088 , \15239 , \15243 );
and \U$20712 ( \21089 , \21088 , \15276 );
and \U$20713 ( \21090 , \15239 , \15243 );
or \U$20714 ( \21091 , \21089 , \21090 );
not \U$20715 ( \21092 , \21091 );
not \U$20716 ( \21093 , \21092 );
or \U$20717 ( \21094 , \15768 , \15716 );
and \U$20718 ( \21095 , \21094 , \15836 );
and \U$20719 ( \21096 , \15768 , \15716 );
nor \U$20720 ( \21097 , \21095 , \21096 );
not \U$20721 ( \21098 , \21097 );
nand \U$20722 ( \21099 , \9774 , RIae7a150_172);
not \U$20723 ( \21100 , \893 );
not \U$20724 ( \21101 , \15817 );
or \U$20725 ( \21102 , \21100 , \21101 );
not \U$20726 ( \21103 , RIae78b48_125);
not \U$20727 ( \21104 , \10084 );
or \U$20728 ( \21105 , \21103 , \21104 );
not \U$20729 ( \21106 , \10084 );
nand \U$20730 ( \21107 , \21106 , \860 );
nand \U$20731 ( \21108 , \21105 , \21107 );
nand \U$20732 ( \21109 , \21108 , \867 );
nand \U$20733 ( \21110 , \21102 , \21109 );
xor \U$20734 ( \21111 , \21099 , \21110 );
not \U$20735 ( \21112 , \951 );
not \U$20736 ( \21113 , \15646 );
or \U$20737 ( \21114 , \21112 , \21113 );
not \U$20738 ( \21115 , RIae78bc0_126);
not \U$20739 ( \21116 , \9941 );
or \U$20740 ( \21117 , \21115 , \21116 );
nand \U$20741 ( \21118 , \15504 , \1286 );
nand \U$20742 ( \21119 , \21117 , \21118 );
nand \U$20743 ( \21120 , \21119 , \926 );
nand \U$20744 ( \21121 , \21114 , \21120 );
xor \U$20745 ( \21122 , \21111 , \21121 );
not \U$20746 ( \21123 , \15821 );
nand \U$20747 ( \21124 , \21123 , \15812 );
not \U$20748 ( \21125 , \21124 );
not \U$20749 ( \21126 , \15832 );
or \U$20750 ( \21127 , \21125 , \21126 );
not \U$20751 ( \21128 , \15812 );
nand \U$20752 ( \21129 , \21128 , \15821 );
nand \U$20753 ( \21130 , \21127 , \21129 );
not \U$20754 ( \21131 , \21130 );
xor \U$20755 ( \21132 , \21122 , \21131 );
not \U$20756 ( \21133 , \15224 );
not \U$20757 ( \21134 , \15236 );
or \U$20758 ( \21135 , \21133 , \21134 );
or \U$20759 ( \21136 , \15236 , \15224 );
nand \U$20760 ( \21137 , \21135 , \21136 );
not \U$20761 ( \21138 , \15213 );
and \U$20762 ( \21139 , \21137 , \21138 );
nor \U$20763 ( \21140 , \15236 , \15225 );
nor \U$20764 ( \21141 , \21139 , \21140 );
xnor \U$20765 ( \21142 , \21132 , \21141 );
not \U$20766 ( \21143 , \15794 );
not \U$20767 ( \21144 , \15800 );
or \U$20768 ( \21145 , \21143 , \21144 );
not \U$20769 ( \21146 , \15778 );
nand \U$20770 ( \21147 , \21146 , \15790 );
nand \U$20771 ( \21148 , \21145 , \21147 );
xnor \U$20772 ( \21149 , \21142 , \21148 );
not \U$20773 ( \21150 , \15528 );
xor \U$20774 ( \21151 , \15517 , \15534 );
not \U$20775 ( \21152 , \21151 );
or \U$20776 ( \21153 , \21150 , \21152 );
nand \U$20777 ( \21154 , \15535 , \15517 );
nand \U$20778 ( \21155 , \21153 , \21154 );
not \U$20779 ( \21156 , \5285 );
not \U$20780 ( \21157 , RIae794a8_145);
not \U$20781 ( \21158 , \1789 );
or \U$20782 ( \21159 , \21157 , \21158 );
nand \U$20783 ( \21160 , \2576 , \3810 );
nand \U$20784 ( \21161 , \21159 , \21160 );
not \U$20785 ( \21162 , \21161 );
or \U$20786 ( \21163 , \21156 , \21162 );
nand \U$20787 ( \21164 , \15786 , \1933 );
nand \U$20788 ( \21165 , \21163 , \21164 );
xor \U$20789 ( \21166 , \15657 , \21165 );
xor \U$20790 ( \21167 , \21155 , \21166 );
buf \U$20791 ( \21168 , \21167 );
not \U$20792 ( \21169 , \21168 );
and \U$20793 ( \21170 , \21149 , \21169 );
not \U$20794 ( \21171 , \21149 );
and \U$20795 ( \21172 , \21171 , \21168 );
nor \U$20796 ( \21173 , \21170 , \21172 );
not \U$20797 ( \21174 , \15834 );
not \U$20798 ( \21175 , \15801 );
or \U$20799 ( \21176 , \21174 , \21175 );
or \U$20800 ( \21177 , \15834 , \15801 );
nand \U$20801 ( \21178 , \21177 , \15773 );
nand \U$20802 ( \21179 , \21176 , \21178 );
not \U$20803 ( \21180 , \21179 );
not \U$20804 ( \21181 , \2272 );
not \U$20805 ( \21182 , \15362 );
or \U$20806 ( \21183 , \21181 , \21182 );
and \U$20807 ( \21184 , RIae79ac0_158, \12997 );
not \U$20808 ( \21185 , RIae79ac0_158);
and \U$20809 ( \21186 , \21185 , \14422 );
or \U$20810 ( \21187 , \21184 , \21186 );
nand \U$20811 ( \21188 , \21187 , \2251 );
nand \U$20812 ( \21189 , \21183 , \21188 );
not \U$20813 ( \21190 , \2602 );
not \U$20814 ( \21191 , \15376 );
or \U$20815 ( \21192 , \21190 , \21191 );
not \U$20816 ( \21193 , RIae79520_146);
not \U$20817 ( \21194 , \13008 );
or \U$20818 ( \21195 , \21193 , \21194 );
or \U$20819 ( \21196 , \14439 , RIae79520_146);
nand \U$20820 ( \21197 , \21195 , \21196 );
nand \U$20821 ( \21198 , \21197 , \3440 );
nand \U$20822 ( \21199 , \21192 , \21198 );
xor \U$20823 ( \21200 , \21189 , \21199 );
not \U$20824 ( \21201 , \6214 );
and \U$20825 ( \21202 , RIae79ef8_167, \6147 );
not \U$20826 ( \21203 , RIae79ef8_167);
and \U$20827 ( \21204 , \21203 , \9625 );
or \U$20828 ( \21205 , \21202 , \21204 );
not \U$20829 ( \21206 , \21205 );
or \U$20830 ( \21207 , \21201 , \21206 );
nand \U$20831 ( \21208 , \15482 , \15989 );
nand \U$20832 ( \21209 , \21207 , \21208 );
xnor \U$20833 ( \21210 , \21200 , \21209 );
not \U$20834 ( \21211 , \6276 );
not \U$20835 ( \21212 , \15686 );
or \U$20836 ( \21213 , \21211 , \21212 );
not \U$20837 ( \21214 , \4844 );
not \U$20838 ( \21215 , \3294 );
or \U$20839 ( \21216 , \21214 , \21215 );
or \U$20840 ( \21217 , \1898 , \10892 );
nand \U$20841 ( \21218 , \21216 , \21217 );
nand \U$20842 ( \21219 , \21218 , \4853 );
nand \U$20843 ( \21220 , \21213 , \21219 );
not \U$20844 ( \21221 , \13720 );
not \U$20845 ( \21222 , \15416 );
or \U$20846 ( \21223 , \21221 , \21222 );
and \U$20847 ( \21224 , RIae7a240_174, \3236 );
not \U$20848 ( \21225 , RIae7a240_174);
and \U$20849 ( \21226 , \21225 , \18413 );
nor \U$20850 ( \21227 , \21224 , \21226 );
nand \U$20851 ( \21228 , \21227 , \13121 );
nand \U$20852 ( \21229 , \21223 , \21228 );
xor \U$20853 ( \21230 , \21220 , \21229 );
not \U$20854 ( \21231 , \11364 );
and \U$20855 ( \21232 , RIae79c28_161, \3244 );
not \U$20856 ( \21233 , RIae79c28_161);
and \U$20857 ( \21234 , \21233 , \3765 );
or \U$20858 ( \21235 , \21232 , \21234 );
not \U$20859 ( \21236 , \21235 );
or \U$20860 ( \21237 , \21231 , \21236 );
nand \U$20861 ( \21238 , \15399 , \2767 );
nand \U$20862 ( \21239 , \21237 , \21238 );
xnor \U$20863 ( \21240 , \21230 , \21239 );
xor \U$20864 ( \21241 , \21210 , \21240 );
not \U$20865 ( \21242 , \11037 );
not \U$20866 ( \21243 , \2442 );
not \U$20867 ( \21244 , \2955 );
or \U$20868 ( \21245 , \21243 , \21244 );
nand \U$20869 ( \21246 , \13142 , RIae79778_151);
nand \U$20870 ( \21247 , \21245 , \21246 );
not \U$20871 ( \21248 , \21247 );
or \U$20872 ( \21249 , \21242 , \21248 );
nand \U$20873 ( \21250 , \15336 , \2545 );
nand \U$20874 ( \21251 , \21249 , \21250 );
not \U$20875 ( \21252 , \10638 );
not \U$20876 ( \21253 , \15405 );
or \U$20877 ( \21254 , \21252 , \21253 );
not \U$20878 ( \21255 , RIae7a510_180);
not \U$20879 ( \21256 , \780 );
or \U$20880 ( \21257 , \21255 , \21256 );
or \U$20881 ( \21258 , \1993 , RIae7a510_180);
nand \U$20882 ( \21259 , \21257 , \21258 );
nand \U$20883 ( \21260 , \21259 , \10631 );
nand \U$20884 ( \21261 , \21254 , \21260 );
xor \U$20885 ( \21262 , \21251 , \21261 );
not \U$20886 ( \21263 , \9792 );
not \U$20887 ( \21264 , \15319 );
or \U$20888 ( \21265 , \21263 , \21264 );
not \U$20889 ( \21266 , RIae7a2b8_175);
not \U$20890 ( \21267 , \878 );
or \U$20891 ( \21268 , \21266 , \21267 );
or \U$20892 ( \21269 , \878 , RIae7a2b8_175);
nand \U$20893 ( \21270 , \21268 , \21269 );
nand \U$20894 ( \21271 , \21270 , \9815 );
nand \U$20895 ( \21272 , \21265 , \21271 );
xnor \U$20896 ( \21273 , \21262 , \21272 );
xor \U$20897 ( \21274 , \21241 , \21273 );
not \U$20898 ( \21275 , \21274 );
or \U$20899 ( \21276 , \21180 , \21275 );
or \U$20900 ( \21277 , \21274 , \21179 );
nand \U$20901 ( \21278 , \21276 , \21277 );
xor \U$20902 ( \21279 , \21173 , \21278 );
not \U$20903 ( \21280 , \21279 );
or \U$20904 ( \21281 , \21098 , \21280 );
or \U$20905 ( \21282 , \21279 , \21097 );
nand \U$20906 ( \21283 , \21281 , \21282 );
not \U$20907 ( \21284 , \21283 );
or \U$20908 ( \21285 , \21093 , \21284 );
or \U$20909 ( \21286 , \21283 , \21092 );
nand \U$20910 ( \21287 , \21285 , \21286 );
not \U$20911 ( \21288 , \21287 );
not \U$20912 ( \21289 , \21288 );
or \U$20913 ( \21290 , \21087 , \21289 );
not \U$20914 ( \21291 , \21086 );
nand \U$20915 ( \21292 , \21291 , \21287 );
nand \U$20916 ( \21293 , \21290 , \21292 );
xnor \U$20917 ( \21294 , \21082 , \21293 );
xor \U$20918 ( \21295 , \15871 , \15903 );
not \U$20919 ( \21296 , \21295 );
not \U$20920 ( \21297 , \15892 );
or \U$20921 ( \21298 , \21296 , \21297 );
nand \U$20922 ( \21299 , \15903 , \15871 );
nand \U$20923 ( \21300 , \21298 , \21299 );
and \U$20924 ( \21301 , \21294 , \21300 );
not \U$20925 ( \21302 , \21294 );
not \U$20926 ( \21303 , \21300 );
and \U$20927 ( \21304 , \21302 , \21303 );
nor \U$20928 ( \21305 , \21301 , \21304 );
nand \U$20929 ( \21306 , \20781 , \21305 );
not \U$20930 ( \21307 , \9517 );
and \U$20931 ( \21308 , RIae79fe8_169, \1118 );
not \U$20932 ( \21309 , RIae79fe8_169);
and \U$20933 ( \21310 , \21309 , \12800 );
nor \U$20934 ( \21311 , \21308 , \21310 );
not \U$20935 ( \21312 , \21311 );
or \U$20936 ( \21313 , \21307 , \21312 );
nand \U$20937 ( \21314 , \21057 , \9499 );
nand \U$20938 ( \21315 , \21313 , \21314 );
not \U$20939 ( \21316 , \2322 );
not \U$20940 ( \21317 , \6171 );
and \U$20941 ( \21318 , RIae798e0_154, \21317 );
not \U$20942 ( \21319 , RIae798e0_154);
and \U$20943 ( \21320 , \21319 , \3094 );
or \U$20944 ( \21321 , \21318 , \21320 );
not \U$20945 ( \21322 , \21321 );
or \U$20946 ( \21323 , \21316 , \21322 );
nand \U$20947 ( \21324 , \21041 , \14580 );
nand \U$20948 ( \21325 , \21323 , \21324 );
not \U$20949 ( \21326 , \21325 );
not \U$20950 ( \21327 , \2096 );
and \U$20951 ( \21328 , \12644 , RIae78b48_125);
not \U$20952 ( \21329 , \12644 );
and \U$20953 ( \21330 , \21329 , \860 );
nor \U$20954 ( \21331 , \21328 , \21330 );
not \U$20955 ( \21332 , \21331 );
or \U$20956 ( \21333 , \21327 , \21332 );
nand \U$20957 ( \21334 , \21108 , \893 );
nand \U$20958 ( \21335 , \21333 , \21334 );
and \U$20959 ( \21336 , \21326 , \21335 );
not \U$20960 ( \21337 , \21326 );
not \U$20961 ( \21338 , \21335 );
and \U$20962 ( \21339 , \21337 , \21338 );
nor \U$20963 ( \21340 , \21336 , \21339 );
xor \U$20964 ( \21341 , \21315 , \21340 );
not \U$20965 ( \21342 , \2163 );
not \U$20966 ( \21343 , RIae79520_146);
not \U$20967 ( \21344 , \2564 );
or \U$20968 ( \21345 , \21343 , \21344 );
nand \U$20969 ( \21346 , \6413 , \4653 );
nand \U$20970 ( \21347 , \21345 , \21346 );
not \U$20971 ( \21348 , \21347 );
or \U$20972 ( \21349 , \21342 , \21348 );
nand \U$20973 ( \21350 , \21197 , \5950 );
nand \U$20974 ( \21351 , \21349 , \21350 );
not \U$20975 ( \21352 , \21351 );
not \U$20976 ( \21353 , \1919 );
and \U$20977 ( \21354 , RIae794a8_145, \1809 );
not \U$20978 ( \21355 , RIae794a8_145);
and \U$20979 ( \21356 , \21355 , \4036 );
or \U$20980 ( \21357 , \21354 , \21356 );
not \U$20981 ( \21358 , \21357 );
or \U$20982 ( \21359 , \21353 , \21358 );
nand \U$20983 ( \21360 , \21161 , \9828 );
nand \U$20984 ( \21361 , \21359 , \21360 );
not \U$20985 ( \21362 , \21361 );
not \U$20986 ( \21363 , \21362 );
or \U$20987 ( \21364 , \21352 , \21363 );
not \U$20988 ( \21365 , \21351 );
nand \U$20989 ( \21366 , \21361 , \21365 );
nand \U$20990 ( \21367 , \21364 , \21366 );
not \U$20991 ( \21368 , \6214 );
not \U$20992 ( \21369 , \9560 );
not \U$20993 ( \21370 , \10916 );
or \U$20994 ( \21371 , \21369 , \21370 );
nand \U$20995 ( \21372 , \1186 , RIae79ef8_167);
nand \U$20996 ( \21373 , \21371 , \21372 );
not \U$20997 ( \21374 , \21373 );
or \U$20998 ( \21375 , \21368 , \21374 );
nand \U$20999 ( \21376 , \21205 , \15989 );
nand \U$21000 ( \21377 , \21375 , \21376 );
and \U$21001 ( \21378 , \21367 , \21377 );
not \U$21002 ( \21379 , \21367 );
not \U$21003 ( \21380 , \21377 );
and \U$21004 ( \21381 , \21379 , \21380 );
nor \U$21005 ( \21382 , \21378 , \21381 );
xor \U$21006 ( \21383 , \21341 , \21382 );
not \U$21007 ( \21384 , \2767 );
not \U$21008 ( \21385 , \21235 );
or \U$21009 ( \21386 , \21384 , \21385 );
not \U$21010 ( \21387 , RIae79c28_161);
not \U$21011 ( \21388 , \2629 );
or \U$21012 ( \21389 , \21387 , \21388 );
nand \U$21013 ( \21390 , \2207 , \10584 );
nand \U$21014 ( \21391 , \21389 , \21390 );
nand \U$21015 ( \21392 , \21391 , \5324 );
nand \U$21016 ( \21393 , \21386 , \21392 );
not \U$21017 ( \21394 , \13121 );
and \U$21018 ( \21395 , RIae7a240_174, \15675 );
not \U$21019 ( \21396 , RIae7a240_174);
and \U$21020 ( \21397 , \21396 , \16589 );
nor \U$21021 ( \21398 , \21395 , \21397 );
not \U$21022 ( \21399 , \21398 );
or \U$21023 ( \21400 , \21394 , \21399 );
nand \U$21024 ( \21401 , \21227 , \13720 );
nand \U$21025 ( \21402 , \21400 , \21401 );
not \U$21026 ( \21403 , \9814 );
not \U$21027 ( \21404 , \11054 );
not \U$21028 ( \21405 , \853 );
or \U$21029 ( \21406 , \21404 , \21405 );
or \U$21030 ( \21407 , \9810 , \853 );
nand \U$21031 ( \21408 , \21406 , \21407 );
not \U$21032 ( \21409 , \21408 );
or \U$21033 ( \21410 , \21403 , \21409 );
nand \U$21034 ( \21411 , \9792 , \21270 );
nand \U$21035 ( \21412 , \21410 , \21411 );
xor \U$21036 ( \21413 , \21402 , \21412 );
xor \U$21037 ( \21414 , \21393 , \21413 );
xor \U$21038 ( \21415 , \21383 , \21414 );
not \U$21039 ( \21416 , \21032 );
nand \U$21040 ( \21417 , \21416 , \21046 );
not \U$21041 ( \21418 , \21417 );
not \U$21042 ( \21419 , \21059 );
or \U$21043 ( \21420 , \21418 , \21419 );
nand \U$21044 ( \21421 , \21032 , \21043 );
nand \U$21045 ( \21422 , \21420 , \21421 );
not \U$21046 ( \21423 , \21229 );
not \U$21047 ( \21424 , \21423 );
not \U$21048 ( \21425 , \21220 );
not \U$21049 ( \21426 , \21425 );
or \U$21050 ( \21427 , \21424 , \21426 );
nand \U$21051 ( \21428 , \21427 , \21239 );
not \U$21052 ( \21429 , \21425 );
nand \U$21053 ( \21430 , \21429 , \21229 );
nand \U$21054 ( \21431 , \21428 , \21430 );
xor \U$21055 ( \21432 , \21422 , \21431 );
not \U$21056 ( \21433 , \21251 );
xor \U$21057 ( \21434 , \21261 , \21272 );
not \U$21058 ( \21435 , \21434 );
or \U$21059 ( \21436 , \21433 , \21435 );
nand \U$21060 ( \21437 , \21272 , \21261 );
nand \U$21061 ( \21438 , \21436 , \21437 );
xor \U$21062 ( \21439 , \21432 , \21438 );
xor \U$21063 ( \21440 , \21415 , \21439 );
not \U$21064 ( \21441 , \1027 );
not \U$21065 ( \21442 , \1286 );
not \U$21066 ( \21443 , \12077 );
or \U$21067 ( \21444 , \21442 , \21443 );
or \U$21068 ( \21445 , \16752 , \12838 );
nand \U$21069 ( \21446 , \21444 , \21445 );
not \U$21070 ( \21447 , \21446 );
or \U$21071 ( \21448 , \21441 , \21447 );
nand \U$21072 ( \21449 , \21119 , \951 );
nand \U$21073 ( \21450 , \21448 , \21449 );
not \U$21074 ( \21451 , \6091 );
not \U$21075 ( \21452 , \20996 );
or \U$21076 ( \21453 , \21451 , \21452 );
not \U$21077 ( \21454 , RIae79d90_164);
not \U$21078 ( \21455 , \12183 );
or \U$21079 ( \21456 , \21454 , \21455 );
or \U$21080 ( \21457 , \5134 , RIae79d90_164);
nand \U$21081 ( \21458 , \21456 , \21457 );
nand \U$21082 ( \21459 , \21458 , \14940 );
nand \U$21083 ( \21460 , \21453 , \21459 );
xor \U$21084 ( \21461 , \21450 , \21460 );
not \U$21085 ( \21462 , \10414 );
not \U$21086 ( \21463 , RIae79ac0_158);
not \U$21087 ( \21464 , \4113 );
or \U$21088 ( \21465 , \21463 , \21464 );
or \U$21089 ( \21466 , \4113 , RIae79ac0_158);
nand \U$21090 ( \21467 , \21465 , \21466 );
not \U$21091 ( \21468 , \21467 );
or \U$21092 ( \21469 , \21462 , \21468 );
nand \U$21093 ( \21470 , \21187 , \2272 );
nand \U$21094 ( \21471 , \21469 , \21470 );
xor \U$21095 ( \21472 , \21461 , \21471 );
not \U$21096 ( \21473 , \1821 );
not \U$21097 ( \21474 , RIae79688_149);
and \U$21098 ( \21475 , \1859 , \21474 );
not \U$21099 ( \21476 , \1859 );
and \U$21100 ( \21477 , \21476 , RIae79688_149);
nor \U$21101 ( \21478 , \21475 , \21477 );
not \U$21102 ( \21479 , \21478 );
or \U$21103 ( \21480 , \21473 , \21479 );
nand \U$21104 ( \21481 , \20897 , \10401 );
nand \U$21105 ( \21482 , \21480 , \21481 );
not \U$21106 ( \21483 , \6276 );
not \U$21107 ( \21484 , \21218 );
or \U$21108 ( \21485 , \21483 , \21484 );
not \U$21109 ( \21486 , \4844 );
not \U$21110 ( \21487 , \4194 );
or \U$21111 ( \21488 , \21486 , \21487 );
or \U$21112 ( \21489 , \4198 , \2406 );
nand \U$21113 ( \21490 , \21488 , \21489 );
nand \U$21114 ( \21491 , \21490 , \4853 );
nand \U$21115 ( \21492 , \21485 , \21491 );
xor \U$21116 ( \21493 , \21482 , \21492 );
not \U$21117 ( \21494 , \10631 );
and \U$21118 ( \21495 , RIae7a510_180, \9711 );
not \U$21119 ( \21496 , RIae7a510_180);
and \U$21120 ( \21497 , \21496 , \828 );
nor \U$21121 ( \21498 , \21495 , \21497 );
not \U$21122 ( \21499 , \21498 );
or \U$21123 ( \21500 , \21494 , \21499 );
nand \U$21124 ( \21501 , \21259 , \11400 );
nand \U$21125 ( \21502 , \21500 , \21501 );
xor \U$21126 ( \21503 , \21493 , \21502 );
xor \U$21127 ( \21504 , \21472 , \21503 );
not \U$21128 ( \21505 , \1988 );
not \U$21129 ( \21506 , \21030 );
or \U$21130 ( \21507 , \21505 , \21506 );
not \U$21131 ( \21508 , \1991 );
not \U$21132 ( \21509 , \2309 );
or \U$21133 ( \21510 , \21508 , \21509 );
nand \U$21134 ( \21511 , \2305 , RIae797f0_152);
nand \U$21135 ( \21512 , \21510 , \21511 );
nand \U$21136 ( \21513 , \21512 , \2007 );
nand \U$21137 ( \21514 , \21507 , \21513 );
not \U$21138 ( \21515 , \12515 );
not \U$21139 ( \21516 , \21007 );
or \U$21140 ( \21517 , \21515 , \21516 );
not \U$21141 ( \21518 , \11690 );
not \U$21142 ( \21519 , \10551 );
or \U$21143 ( \21520 , \21518 , \21519 );
or \U$21144 ( \21521 , \10551 , \11695 );
nand \U$21145 ( \21522 , \21520 , \21521 );
nand \U$21146 ( \21523 , \21522 , \9622 );
nand \U$21147 ( \21524 , \21517 , \21523 );
xor \U$21148 ( \21525 , \21514 , \21524 );
not \U$21149 ( \21526 , \2450 );
not \U$21150 ( \21527 , \2504 );
not \U$21151 ( \21528 , \9501 );
or \U$21152 ( \21529 , \21527 , \21528 );
nand \U$21153 ( \21530 , \2140 , RIae79778_151);
nand \U$21154 ( \21531 , \21529 , \21530 );
not \U$21155 ( \21532 , \21531 );
or \U$21156 ( \21533 , \21526 , \21532 );
nand \U$21157 ( \21534 , \21247 , \2545 );
nand \U$21158 ( \21535 , \21533 , \21534 );
xor \U$21159 ( \21536 , \21525 , \21535 );
not \U$21160 ( \21537 , \21536 );
xnor \U$21161 ( \21538 , \21504 , \21537 );
xor \U$21162 ( \21539 , \21440 , \21538 );
not \U$21163 ( \21540 , \21142 );
not \U$21164 ( \21541 , \21167 );
or \U$21165 ( \21542 , \21540 , \21541 );
or \U$21166 ( \21543 , \21142 , \21167 );
nand \U$21167 ( \21544 , \21543 , \21148 );
nand \U$21168 ( \21545 , \21542 , \21544 );
not \U$21169 ( \21546 , \21021 );
nand \U$21170 ( \21547 , \21546 , \21064 );
not \U$21171 ( \21548 , \21547 );
not \U$21172 ( \21549 , \20991 );
or \U$21173 ( \21550 , \21548 , \21549 );
or \U$21174 ( \21551 , \21546 , \21064 );
nand \U$21175 ( \21552 , \21550 , \21551 );
and \U$21176 ( \21553 , \21545 , \21552 );
not \U$21177 ( \21554 , \21545 );
not \U$21178 ( \21555 , \21552 );
and \U$21179 ( \21556 , \21554 , \21555 );
nor \U$21180 ( \21557 , \21553 , \21556 );
xor \U$21181 ( \21558 , \21099 , \21110 );
and \U$21182 ( \21559 , \21558 , \21121 );
and \U$21183 ( \21560 , \21099 , \21110 );
or \U$21184 ( \21561 , \21559 , \21560 );
not \U$21185 ( \21562 , \20963 );
not \U$21186 ( \21563 , \20939 );
and \U$21187 ( \21564 , \20953 , \21563 );
not \U$21188 ( \21565 , \20953 );
and \U$21189 ( \21566 , \21565 , \20939 );
nor \U$21190 ( \21567 , \21564 , \21566 );
not \U$21191 ( \21568 , \21567 );
or \U$21192 ( \21569 , \21562 , \21568 );
nand \U$21193 ( \21570 , \20953 , \21563 );
nand \U$21194 ( \21571 , \21569 , \21570 );
xor \U$21195 ( \21572 , \21561 , \21571 );
not \U$21196 ( \21573 , \20899 );
not \U$21197 ( \21574 , \20916 );
or \U$21198 ( \21575 , \21573 , \21574 );
not \U$21199 ( \21576 , \20902 );
nand \U$21200 ( \21577 , \21576 , \20912 );
nand \U$21201 ( \21578 , \21575 , \21577 );
xor \U$21202 ( \21579 , \21572 , \21578 );
not \U$21203 ( \21580 , \21579 );
not \U$21204 ( \21581 , \21122 );
nand \U$21205 ( \21582 , \21581 , \21131 );
not \U$21206 ( \21583 , \21582 );
not \U$21207 ( \21584 , \21141 );
or \U$21208 ( \21585 , \21583 , \21584 );
nand \U$21209 ( \21586 , \21130 , \21122 );
nand \U$21210 ( \21587 , \21585 , \21586 );
not \U$21211 ( \21588 , \21587 );
not \U$21212 ( \21589 , \21165 );
nand \U$21213 ( \21590 , \21589 , \15660 );
not \U$21214 ( \21591 , \21590 );
not \U$21215 ( \21592 , \21155 );
or \U$21216 ( \21593 , \21591 , \21592 );
not \U$21217 ( \21594 , \21589 );
nand \U$21218 ( \21595 , \21594 , \15657 );
nand \U$21219 ( \21596 , \21593 , \21595 );
not \U$21220 ( \21597 , \21596 );
not \U$21221 ( \21598 , \21597 );
or \U$21222 ( \21599 , \21588 , \21598 );
or \U$21223 ( \21600 , \21597 , \21587 );
nand \U$21224 ( \21601 , \21599 , \21600 );
not \U$21225 ( \21602 , \21601 );
not \U$21226 ( \21603 , \21602 );
or \U$21227 ( \21604 , \21580 , \21603 );
not \U$21228 ( \21605 , \21579 );
nand \U$21229 ( \21606 , \21605 , \21601 );
nand \U$21230 ( \21607 , \21604 , \21606 );
xor \U$21231 ( \21608 , \21557 , \21607 );
xor \U$21232 ( \21609 , \21539 , \21608 );
or \U$21233 ( \21610 , \20806 , \20815 );
nand \U$21234 ( \21611 , \21610 , \20820 );
nand \U$21235 ( \21612 , \20815 , \20806 );
nand \U$21236 ( \21613 , \21611 , \21612 );
xor \U$21237 ( \21614 , \21609 , \21613 );
not \U$21238 ( \21615 , \21283 );
not \U$21239 ( \21616 , \21091 );
or \U$21240 ( \21617 , \21615 , \21616 );
not \U$21241 ( \21618 , \21097 );
nand \U$21242 ( \21619 , \21618 , \21279 );
nand \U$21243 ( \21620 , \21617 , \21619 );
xor \U$21244 ( \21621 , \21614 , \21620 );
xor \U$21245 ( \21622 , \20821 , \21072 );
and \U$21246 ( \21623 , \21622 , \21080 );
and \U$21247 ( \21624 , \20821 , \21072 );
or \U$21248 ( \21625 , \21623 , \21624 );
xor \U$21249 ( \21626 , \21621 , \21625 );
not \U$21250 ( \21627 , \21626 );
xor \U$21251 ( \21628 , \20964 , \20968 );
and \U$21252 ( \21629 , \21628 , \20973 );
and \U$21253 ( \21630 , \20964 , \20968 );
or \U$21254 ( \21631 , \21629 , \21630 );
or \U$21255 ( \21632 , \20837 , \20842 );
nand \U$21256 ( \21633 , \21632 , \20847 );
nand \U$21257 ( \21634 , \20837 , \20842 );
nand \U$21258 ( \21635 , \21633 , \21634 );
and \U$21259 ( \21636 , \21631 , \21635 );
not \U$21260 ( \21637 , \21631 );
not \U$21261 ( \21638 , \21635 );
and \U$21262 ( \21639 , \21637 , \21638 );
nor \U$21263 ( \21640 , \21636 , \21639 );
not \U$21264 ( \21641 , \21640 );
not \U$21265 ( \21642 , \20930 );
not \U$21266 ( \21643 , \20925 );
or \U$21267 ( \21644 , \21642 , \21643 );
or \U$21268 ( \21645 , \20921 , \20888 );
nand \U$21269 ( \21646 , \21644 , \21645 );
not \U$21270 ( \21647 , \21646 );
and \U$21271 ( \21648 , \21641 , \21647 );
and \U$21272 ( \21649 , \21646 , \21640 );
nor \U$21273 ( \21650 , \21648 , \21649 );
buf \U$21274 ( \21651 , \20852 );
or \U$21275 ( \21652 , \20931 , \21651 );
nand \U$21276 ( \21653 , \21652 , \20856 );
nand \U$21277 ( \21654 , \20931 , \21651 );
nand \U$21278 ( \21655 , \21653 , \21654 );
xor \U$21279 ( \21656 , \21650 , \21655 );
xor \U$21280 ( \21657 , \20789 , \20798 );
and \U$21281 ( \21658 , \21657 , \20805 );
and \U$21282 ( \21659 , \20789 , \20798 );
or \U$21283 ( \21660 , \21658 , \21659 );
xnor \U$21284 ( \21661 , \21656 , \21660 );
not \U$21285 ( \21662 , \20831 );
not \U$21286 ( \21663 , \20932 );
or \U$21287 ( \21664 , \21662 , \21663 );
nand \U$21288 ( \21665 , \21664 , \21070 );
not \U$21289 ( \21666 , \20831 );
not \U$21290 ( \21667 , \20932 );
nand \U$21291 ( \21668 , \21666 , \21667 );
nand \U$21292 ( \21669 , \21665 , \21668 );
not \U$21293 ( \21670 , \21669 );
nand \U$21294 ( \21671 , \21661 , \21670 );
not \U$21295 ( \21672 , \21670 );
not \U$21296 ( \21673 , \21661 );
nand \U$21297 ( \21674 , \21672 , \21673 );
nand \U$21298 ( \21675 , \21671 , \21674 );
not \U$21299 ( \21676 , \21209 );
or \U$21300 ( \21677 , \21199 , \21189 );
not \U$21301 ( \21678 , \21677 );
or \U$21302 ( \21679 , \21676 , \21678 );
nand \U$21303 ( \21680 , \21199 , \21189 );
nand \U$21304 ( \21681 , \21679 , \21680 );
not \U$21305 ( \21682 , \20876 );
not \U$21306 ( \21683 , \20867 );
not \U$21307 ( \21684 , \21683 );
not \U$21308 ( \21685 , \20887 );
or \U$21309 ( \21686 , \21684 , \21685 );
or \U$21310 ( \21687 , \20887 , \21683 );
nand \U$21311 ( \21688 , \21686 , \21687 );
not \U$21312 ( \21689 , \21688 );
or \U$21313 ( \21690 , \21682 , \21689 );
nand \U$21314 ( \21691 , \20887 , \20867 );
nand \U$21315 ( \21692 , \21690 , \21691 );
xor \U$21316 ( \21693 , \21681 , \21692 );
xor \U$21317 ( \21694 , \21000 , \21009 );
and \U$21318 ( \21695 , \21694 , \21020 );
and \U$21319 ( \21696 , \21000 , \21009 );
or \U$21320 ( \21697 , \21695 , \21696 );
xor \U$21321 ( \21698 , \21693 , \21697 );
or \U$21322 ( \21699 , \10071 , \860 );
not \U$21323 ( \21700 , \1863 );
not \U$21324 ( \21701 , RIae793b8_143);
not \U$21325 ( \21702 , \4960 );
or \U$21326 ( \21703 , \21701 , \21702 );
nand \U$21327 ( \21704 , \17009 , \1884 );
nand \U$21328 ( \21705 , \21703 , \21704 );
not \U$21329 ( \21706 , \21705 );
or \U$21330 ( \21707 , \21700 , \21706 );
nand \U$21331 ( \21708 , \20863 , \1910 );
nand \U$21332 ( \21709 , \21707 , \21708 );
xor \U$21333 ( \21710 , \21699 , \21709 );
not \U$21334 ( \21711 , \2063 );
not \U$21335 ( \21712 , \20908 );
or \U$21336 ( \21713 , \21711 , \21712 );
and \U$21337 ( \21714 , \13999 , \2056 );
not \U$21338 ( \21715 , \13999 );
and \U$21339 ( \21716 , \21715 , RIae79610_148);
nor \U$21340 ( \21717 , \21714 , \21716 );
nand \U$21341 ( \21718 , \21717 , \2011 );
nand \U$21342 ( \21719 , \21713 , \21718 );
xnor \U$21343 ( \21720 , \21710 , \21719 );
not \U$21344 ( \21721 , \10451 );
not \U$21345 ( \21722 , RIae79160_138);
not \U$21346 ( \21723 , \12687 );
or \U$21347 ( \21724 , \21722 , \21723 );
or \U$21348 ( \21725 , \15217 , RIae79160_138);
nand \U$21349 ( \21726 , \21724 , \21725 );
not \U$21350 ( \21727 , \21726 );
or \U$21351 ( \21728 , \21721 , \21727 );
nand \U$21352 ( \21729 , \20885 , \1008 );
nand \U$21353 ( \21730 , \21728 , \21729 );
not \U$21354 ( \21731 , \1501 );
not \U$21355 ( \21732 , \13976 );
and \U$21356 ( \21733 , RIae79250_140, \21732 );
not \U$21357 ( \21734 , RIae79250_140);
and \U$21358 ( \21735 , \21734 , \15207 );
nor \U$21359 ( \21736 , \21733 , \21735 );
not \U$21360 ( \21737 , \21736 );
or \U$21361 ( \21738 , \21731 , \21737 );
nand \U$21362 ( \21739 , \20874 , \9403 );
nand \U$21363 ( \21740 , \21738 , \21739 );
xor \U$21364 ( \21741 , \21730 , \21740 );
not \U$21365 ( \21742 , \1049 );
not \U$21366 ( \21743 , \17387 );
not \U$21367 ( \21744 , \21743 );
and \U$21368 ( \21745 , RIae79070_136, \21744 );
not \U$21369 ( \21746 , RIae79070_136);
not \U$21370 ( \21747 , \12707 );
and \U$21371 ( \21748 , \21746 , \21747 );
or \U$21372 ( \21749 , \21745 , \21748 );
not \U$21373 ( \21750 , \21749 );
or \U$21374 ( \21751 , \21742 , \21750 );
nand \U$21375 ( \21752 , \20951 , \2276 );
nand \U$21376 ( \21753 , \21751 , \21752 );
xor \U$21377 ( \21754 , \21741 , \21753 );
xor \U$21378 ( \21755 , \21720 , \21754 );
not \U$21379 ( \21756 , \839 );
not \U$21380 ( \21757 , \3105 );
not \U$21381 ( \21758 , \14110 );
or \U$21382 ( \21759 , \21757 , \21758 );
nand \U$21383 ( \21760 , \20941 , RIae78f80_134);
nand \U$21384 ( \21761 , \21759 , \21760 );
not \U$21385 ( \21762 , \21761 );
or \U$21386 ( \21763 , \21756 , \21762 );
nand \U$21387 ( \21764 , \20961 , \796 );
nand \U$21388 ( \21765 , \21763 , \21764 );
not \U$21389 ( \21766 , \1320 );
not \U$21390 ( \21767 , \921 );
not \U$21391 ( \21768 , \12088 );
or \U$21392 ( \21769 , \21767 , \21768 );
not \U$21393 ( \21770 , \10936 );
nand \U$21394 ( \21771 , \21770 , RIae78e90_132);
nand \U$21395 ( \21772 , \21769 , \21771 );
not \U$21396 ( \21773 , \21772 );
or \U$21397 ( \21774 , \21766 , \21773 );
not \U$21398 ( \21775 , \20934 );
nand \U$21399 ( \21776 , \21775 , \1086 );
nand \U$21400 ( \21777 , \21774 , \21776 );
xor \U$21401 ( \21778 , \21765 , \21777 );
not \U$21402 ( \21779 , \16564 );
not \U$21403 ( \21780 , \21016 );
or \U$21404 ( \21781 , \21779 , \21780 );
nand \U$21405 ( \21782 , \11422 , RIae7a498_179);
nand \U$21406 ( \21783 , \21781 , \21782 );
xor \U$21407 ( \21784 , \21778 , \21783 );
xor \U$21408 ( \21785 , \21755 , \21784 );
xor \U$21409 ( \21786 , \21698 , \21785 );
xor \U$21410 ( \21787 , \21210 , \21240 );
and \U$21411 ( \21788 , \21787 , \21273 );
and \U$21412 ( \21789 , \21210 , \21240 );
or \U$21413 ( \21790 , \21788 , \21789 );
xor \U$21414 ( \21791 , \21786 , \21790 );
not \U$21415 ( \21792 , \20974 );
not \U$21416 ( \21793 , \21069 );
or \U$21417 ( \21794 , \21792 , \21793 );
not \U$21418 ( \21795 , \20978 );
nand \U$21419 ( \21796 , \21794 , \21795 );
or \U$21420 ( \21797 , \20974 , \21069 );
nand \U$21421 ( \21798 , \21796 , \21797 );
xor \U$21422 ( \21799 , \21791 , \21798 );
not \U$21423 ( \21800 , \21173 );
not \U$21424 ( \21801 , \21278 );
or \U$21425 ( \21802 , \21800 , \21801 );
not \U$21426 ( \21803 , \21274 );
nand \U$21427 ( \21804 , \21803 , \21179 );
nand \U$21428 ( \21805 , \21802 , \21804 );
xor \U$21429 ( \21806 , \21799 , \21805 );
buf \U$21430 ( \21807 , \21806 );
xor \U$21431 ( \21808 , \21675 , \21807 );
not \U$21432 ( \21809 , \21808 );
not \U$21433 ( \21810 , \20785 );
not \U$21434 ( \21811 , \21287 );
or \U$21435 ( \21812 , \21810 , \21811 );
or \U$21436 ( \21813 , \20785 , \21287 );
nand \U$21437 ( \21814 , \21813 , \21086 );
nand \U$21438 ( \21815 , \21812 , \21814 );
not \U$21439 ( \21816 , \21815 );
or \U$21440 ( \21817 , \21809 , \21816 );
or \U$21441 ( \21818 , \21808 , \21815 );
nand \U$21442 ( \21819 , \21817 , \21818 );
not \U$21443 ( \21820 , \21819 );
or \U$21444 ( \21821 , \21627 , \21820 );
not \U$21445 ( \21822 , \21808 );
nand \U$21446 ( \21823 , \21815 , \21822 );
nand \U$21447 ( \21824 , \21821 , \21823 );
xor \U$21448 ( \21825 , \21681 , \21692 );
and \U$21449 ( \21826 , \21825 , \21697 );
and \U$21450 ( \21827 , \21681 , \21692 );
or \U$21451 ( \21828 , \21826 , \21827 );
not \U$21452 ( \21829 , \21503 );
not \U$21453 ( \21830 , \21536 );
or \U$21454 ( \21831 , \21829 , \21830 );
not \U$21455 ( \21832 , \21472 );
nand \U$21456 ( \21833 , \21831 , \21832 );
not \U$21457 ( \21834 , \21503 );
nand \U$21458 ( \21835 , \21834 , \21537 );
nand \U$21459 ( \21836 , \21833 , \21835 );
xor \U$21460 ( \21837 , \21828 , \21836 );
xor \U$21461 ( \21838 , \21341 , \21382 );
and \U$21462 ( \21839 , \21838 , \21414 );
and \U$21463 ( \21840 , \21341 , \21382 );
or \U$21464 ( \21841 , \21839 , \21840 );
xor \U$21465 ( \21842 , \21837 , \21841 );
not \U$21466 ( \21843 , \21439 );
not \U$21467 ( \21844 , \21415 );
or \U$21468 ( \21845 , \21843 , \21844 );
or \U$21469 ( \21846 , \21415 , \21439 );
nand \U$21470 ( \21847 , \21846 , \21538 );
nand \U$21471 ( \21848 , \21845 , \21847 );
xnor \U$21472 ( \21849 , \21842 , \21848 );
not \U$21473 ( \21850 , \21849 );
not \U$21474 ( \21851 , \1501 );
not \U$21475 ( \21852 , \1503 );
not \U$21476 ( \21853 , \16311 );
or \U$21477 ( \21854 , \21852 , \21853 );
nand \U$21478 ( \21855 , \6257 , RIae79250_140);
nand \U$21479 ( \21856 , \21854 , \21855 );
not \U$21480 ( \21857 , \21856 );
or \U$21481 ( \21858 , \21851 , \21857 );
nand \U$21482 ( \21859 , \21736 , \9403 );
nand \U$21483 ( \21860 , \21858 , \21859 );
not \U$21484 ( \21861 , \2063 );
not \U$21485 ( \21862 , \21717 );
or \U$21486 ( \21863 , \21861 , \21862 );
and \U$21487 ( \21864 , \6674 , \2403 );
not \U$21488 ( \21865 , \6674 );
not \U$21489 ( \21866 , \2403 );
and \U$21490 ( \21867 , \21865 , \21866 );
nor \U$21491 ( \21868 , \21864 , \21867 );
nand \U$21492 ( \21869 , \21868 , \2011 );
nand \U$21493 ( \21870 , \21863 , \21869 );
xor \U$21494 ( \21871 , \21860 , \21870 );
not \U$21495 ( \21872 , \1864 );
buf \U$21496 ( \21873 , \6242 );
and \U$21497 ( \21874 , RIae793b8_143, \21873 );
not \U$21498 ( \21875 , RIae793b8_143);
and \U$21499 ( \21876 , \21875 , \4169 );
or \U$21500 ( \21877 , \21874 , \21876 );
not \U$21501 ( \21878 , \21877 );
or \U$21502 ( \21879 , \21872 , \21878 );
nand \U$21503 ( \21880 , \21705 , \1910 );
nand \U$21504 ( \21881 , \21879 , \21880 );
xor \U$21505 ( \21882 , \21871 , \21881 );
not \U$21506 ( \21883 , \21340 );
not \U$21507 ( \21884 , \21315 );
not \U$21508 ( \21885 , \21884 );
or \U$21509 ( \21886 , \21883 , \21885 );
nand \U$21510 ( \21887 , \21326 , \21335 );
nand \U$21511 ( \21888 , \21886 , \21887 );
xor \U$21512 ( \21889 , \21882 , \21888 );
not \U$21513 ( \21890 , \21365 );
not \U$21514 ( \21891 , \21362 );
or \U$21515 ( \21892 , \21890 , \21891 );
nand \U$21516 ( \21893 , \21892 , \21377 );
nand \U$21517 ( \21894 , \21361 , \21351 );
and \U$21518 ( \21895 , \21893 , \21894 );
not \U$21519 ( \21896 , \21895 );
xnor \U$21520 ( \21897 , \21889 , \21896 );
not \U$21521 ( \21898 , \2157 );
not \U$21522 ( \21899 , \21726 );
or \U$21523 ( \21900 , \21898 , \21899 );
and \U$21524 ( \21901 , RIae79160_138, \9291 );
not \U$21525 ( \21902 , RIae79160_138);
and \U$21526 ( \21903 , \21902 , \6345 );
or \U$21527 ( \21904 , \21901 , \21903 );
nand \U$21528 ( \21905 , \21904 , \10451 );
nand \U$21529 ( \21906 , \21900 , \21905 );
not \U$21530 ( \21907 , \839 );
not \U$21531 ( \21908 , \3105 );
not \U$21532 ( \21909 , \15088 );
or \U$21533 ( \21910 , \21908 , \21909 );
nand \U$21534 ( \21911 , \13287 , RIae78f80_134);
nand \U$21535 ( \21912 , \21910 , \21911 );
not \U$21536 ( \21913 , \21912 );
or \U$21537 ( \21914 , \21907 , \21913 );
nand \U$21538 ( \21915 , \21761 , \797 );
nand \U$21539 ( \21916 , \21914 , \21915 );
and \U$21540 ( \21917 , \21906 , \21916 );
not \U$21541 ( \21918 , \21906 );
not \U$21542 ( \21919 , \21916 );
and \U$21543 ( \21920 , \21918 , \21919 );
or \U$21544 ( \21921 , \21917 , \21920 );
not \U$21545 ( \21922 , \1062 );
not \U$21546 ( \21923 , \21749 );
or \U$21547 ( \21924 , \21922 , \21923 );
not \U$21548 ( \21925 , RIae79070_136);
not \U$21549 ( \21926 , \9316 );
or \U$21550 ( \21927 , \21925 , \21926 );
or \U$21551 ( \21928 , \9313 , RIae79070_136);
nand \U$21552 ( \21929 , \21927 , \21928 );
nand \U$21553 ( \21930 , \21929 , \1049 );
nand \U$21554 ( \21931 , \21924 , \21930 );
xor \U$21555 ( \21932 , \21921 , \21931 );
not \U$21556 ( \21933 , \21932 );
not \U$21557 ( \21934 , \951 );
not \U$21558 ( \21935 , \21446 );
or \U$21559 ( \21936 , \21934 , \21935 );
not \U$21560 ( \21937 , RIae78bc0_126);
not \U$21561 ( \21938 , \11804 );
or \U$21562 ( \21939 , \21937 , \21938 );
or \U$21563 ( \21940 , \9412 , RIae78bc0_126);
nand \U$21564 ( \21941 , \21939 , \21940 );
nand \U$21565 ( \21942 , \21941 , \1027 );
nand \U$21566 ( \21943 , \21936 , \21942 );
not \U$21567 ( \21944 , \21943 );
not \U$21568 ( \21945 , \5858 );
not \U$21569 ( \21946 , \21772 );
or \U$21570 ( \21947 , \21945 , \21946 );
not \U$21571 ( \21948 , \9455 );
and \U$21572 ( \21949 , RIae78e90_132, \21948 );
not \U$21573 ( \21950 , RIae78e90_132);
and \U$21574 ( \21951 , \21950 , \9459 );
or \U$21575 ( \21952 , \21949 , \21951 );
nand \U$21576 ( \21953 , \21952 , \1320 );
nand \U$21577 ( \21954 , \21947 , \21953 );
not \U$21578 ( \21955 , \21954 );
or \U$21579 ( \21956 , \21944 , \21955 );
or \U$21580 ( \21957 , \21954 , \21943 );
nand \U$21581 ( \21958 , \21956 , \21957 );
not \U$21582 ( \21959 , \14940 );
and \U$21583 ( \21960 , RIae79d90_164, \6147 );
not \U$21584 ( \21961 , RIae79d90_164);
and \U$21585 ( \21962 , \21961 , \2848 );
or \U$21586 ( \21963 , \21960 , \21962 );
not \U$21587 ( \21964 , \21963 );
or \U$21588 ( \21965 , \21959 , \21964 );
nand \U$21589 ( \21966 , \21458 , \6091 );
nand \U$21590 ( \21967 , \21965 , \21966 );
xor \U$21591 ( \21968 , \21958 , \21967 );
xnor \U$21592 ( \21969 , \21933 , \21968 );
not \U$21593 ( \21970 , \14580 );
not \U$21594 ( \21971 , \21321 );
or \U$21595 ( \21972 , \21970 , \21971 );
and \U$21596 ( \21973 , RIae798e0_154, \2835 );
not \U$21597 ( \21974 , RIae798e0_154);
and \U$21598 ( \21975 , \21974 , \3748 );
or \U$21599 ( \21976 , \21973 , \21975 );
nand \U$21600 ( \21977 , \21976 , \2322 );
nand \U$21601 ( \21978 , \21972 , \21977 );
not \U$21602 ( \21979 , \2007 );
and \U$21603 ( \21980 , RIae797f0_152, \2153 );
not \U$21604 ( \21981 , RIae797f0_152);
and \U$21605 ( \21982 , \21981 , \2955 );
or \U$21606 ( \21983 , \21980 , \21982 );
not \U$21607 ( \21984 , \21983 );
or \U$21608 ( \21985 , \21979 , \21984 );
nand \U$21609 ( \21986 , \21512 , \1989 );
nand \U$21610 ( \21987 , \21985 , \21986 );
xor \U$21611 ( \21988 , \21978 , \21987 );
not \U$21612 ( \21989 , \9499 );
not \U$21613 ( \21990 , \21311 );
or \U$21614 ( \21991 , \21989 , \21990 );
not \U$21615 ( \21992 , \11069 );
not \U$21616 ( \21993 , \883 );
or \U$21617 ( \21994 , \21992 , \21993 );
nand \U$21618 ( \21995 , \2175 , RIae79fe8_169);
nand \U$21619 ( \21996 , \21994 , \21995 );
nand \U$21620 ( \21997 , \21996 , \9518 );
nand \U$21621 ( \21998 , \21991 , \21997 );
xor \U$21622 ( \21999 , \21988 , \21998 );
not \U$21623 ( \22000 , \21999 );
and \U$21624 ( \22001 , \21969 , \22000 );
not \U$21625 ( \22002 , \21969 );
and \U$21626 ( \22003 , \22002 , \21999 );
nor \U$21627 ( \22004 , \22001 , \22003 );
not \U$21628 ( \22005 , \22004 );
and \U$21629 ( \22006 , \21897 , \22005 );
not \U$21630 ( \22007 , \21897 );
and \U$21631 ( \22008 , \22007 , \22004 );
nor \U$21632 ( \22009 , \22006 , \22008 );
xor \U$21633 ( \22010 , \21482 , \21492 );
and \U$21634 ( \22011 , \22010 , \21502 );
and \U$21635 ( \22012 , \21482 , \21492 );
or \U$21636 ( \22013 , \22011 , \22012 );
nor \U$21637 ( \22014 , \21535 , \21514 );
not \U$21638 ( \22015 , \21524 );
or \U$21639 ( \22016 , \22014 , \22015 );
nand \U$21640 ( \22017 , \21535 , \21514 );
nand \U$21641 ( \22018 , \22016 , \22017 );
xor \U$21642 ( \22019 , \22013 , \22018 );
not \U$21643 ( \22020 , \21393 );
not \U$21644 ( \22021 , \21413 );
or \U$21645 ( \22022 , \22020 , \22021 );
nand \U$21646 ( \22023 , \21412 , \21402 );
nand \U$21647 ( \22024 , \22022 , \22023 );
xnor \U$21648 ( \22025 , \22019 , \22024 );
and \U$21649 ( \22026 , \22009 , \22025 );
not \U$21650 ( \22027 , \22009 );
not \U$21651 ( \22028 , \22025 );
and \U$21652 ( \22029 , \22027 , \22028 );
nor \U$21653 ( \22030 , \22026 , \22029 );
not \U$21654 ( \22031 , \22030 );
and \U$21655 ( \22032 , \21850 , \22031 );
and \U$21656 ( \22033 , \21849 , \22030 );
nor \U$21657 ( \22034 , \22032 , \22033 );
not \U$21658 ( \22035 , \22034 );
not \U$21659 ( \22036 , \21798 );
not \U$21660 ( \22037 , \21805 );
not \U$21661 ( \22038 , \22037 );
or \U$21662 ( \22039 , \22036 , \22038 );
or \U$21663 ( \22040 , \22037 , \21798 );
nand \U$21664 ( \22041 , \22040 , \21791 );
nand \U$21665 ( \22042 , \22039 , \22041 );
not \U$21666 ( \22043 , \2189 );
not \U$21667 ( \22044 , \21347 );
or \U$21668 ( \22045 , \22043 , \22044 );
not \U$21669 ( \22046 , RIae79520_146);
not \U$21670 ( \22047 , \1788 );
or \U$21671 ( \22048 , \22046 , \22047 );
or \U$21672 ( \22049 , \1788 , RIae79520_146);
nand \U$21673 ( \22050 , \22048 , \22049 );
nand \U$21674 ( \22051 , \22050 , \2610 );
nand \U$21675 ( \22052 , \22045 , \22051 );
and \U$21676 ( \22053 , RIae7a150_172, RIae7a420_178);
nor \U$21677 ( \22054 , \22053 , \10625 );
nand \U$21678 ( \22055 , \10207 , RIae78b48_125);
xor \U$21679 ( \22056 , \22054 , \22055 );
not \U$21680 ( \22057 , \893 );
not \U$21681 ( \22058 , \21331 );
or \U$21682 ( \22059 , \22057 , \22058 );
and \U$21683 ( \22060 , \11186 , RIae78b48_125);
not \U$21684 ( \22061 , \11186 );
and \U$21685 ( \22062 , \22061 , \860 );
nor \U$21686 ( \22063 , \22060 , \22062 );
nand \U$21687 ( \22064 , \22063 , \867 );
nand \U$21688 ( \22065 , \22059 , \22064 );
xor \U$21689 ( \22066 , \22056 , \22065 );
nor \U$21690 ( \22067 , \22052 , \22066 );
not \U$21691 ( \22068 , \22067 );
nand \U$21692 ( \22069 , \22052 , \22066 );
nand \U$21693 ( \22070 , \22068 , \22069 );
not \U$21694 ( \22071 , \21709 );
xnor \U$21695 ( \22072 , \21699 , \21719 );
not \U$21696 ( \22073 , \22072 );
or \U$21697 ( \22074 , \22071 , \22073 );
not \U$21698 ( \22075 , \21699 );
nand \U$21699 ( \22076 , \22075 , \21719 );
nand \U$21700 ( \22077 , \22074 , \22076 );
xnor \U$21701 ( \22078 , \22070 , \22077 );
not \U$21702 ( \22079 , \21422 );
not \U$21703 ( \22080 , \21431 );
or \U$21704 ( \22081 , \22079 , \22080 );
not \U$21705 ( \22082 , \21422 );
nand \U$21706 ( \22083 , \22082 , \21428 , \21430 );
nand \U$21707 ( \22084 , \21438 , \22083 );
nand \U$21708 ( \22085 , \22081 , \22084 );
xor \U$21709 ( \22086 , \22078 , \22085 );
xor \U$21710 ( \22087 , \21720 , \21784 );
and \U$21711 ( \22088 , \22087 , \21754 );
and \U$21712 ( \22089 , \21720 , \21784 );
or \U$21713 ( \22090 , \22088 , \22089 );
xor \U$21714 ( \22091 , \22086 , \22090 );
not \U$21715 ( \22092 , \22091 );
not \U$21716 ( \22093 , \21579 );
not \U$21717 ( \22094 , \21601 );
or \U$21718 ( \22095 , \22093 , \22094 );
nand \U$21719 ( \22096 , \21596 , \21587 );
nand \U$21720 ( \22097 , \22095 , \22096 );
not \U$21721 ( \22098 , \22097 );
nand \U$21722 ( \22099 , \22092 , \22098 );
nand \U$21723 ( \22100 , \22091 , \22097 );
nand \U$21724 ( \22101 , \22099 , \22100 );
not \U$21725 ( \22102 , \21790 );
buf \U$21726 ( \22103 , \21785 );
or \U$21727 ( \22104 , \22102 , \22103 );
nand \U$21728 ( \22105 , \22104 , \21698 );
nand \U$21729 ( \22106 , \22102 , \22103 );
nand \U$21730 ( \22107 , \22105 , \22106 );
and \U$21731 ( \22108 , \22101 , \22107 );
not \U$21732 ( \22109 , \22101 );
not \U$21733 ( \22110 , \22107 );
and \U$21734 ( \22111 , \22109 , \22110 );
nor \U$21735 ( \22112 , \22108 , \22111 );
not \U$21736 ( \22113 , \22112 );
and \U$21737 ( \22114 , \22042 , \22113 );
not \U$21738 ( \22115 , \22042 );
and \U$21739 ( \22116 , \22115 , \22112 );
nor \U$21740 ( \22117 , \22114 , \22116 );
xnor \U$21741 ( \22118 , \22035 , \22117 );
not \U$21742 ( \22119 , \22118 );
not \U$21743 ( \22120 , \21539 );
not \U$21744 ( \22121 , \21608 );
or \U$21745 ( \22122 , \22120 , \22121 );
or \U$21746 ( \22123 , \21608 , \21539 );
nand \U$21747 ( \22124 , \22123 , \21613 );
nand \U$21748 ( \22125 , \22122 , \22124 );
not \U$21749 ( \22126 , \21607 );
not \U$21750 ( \22127 , \21557 );
or \U$21751 ( \22128 , \22126 , \22127 );
nand \U$21752 ( \22129 , \21545 , \21552 );
nand \U$21753 ( \22130 , \22128 , \22129 );
not \U$21754 ( \22131 , \4853 );
not \U$21755 ( \22132 , RIae79ca0_162);
not \U$21756 ( \22133 , \17067 );
or \U$21757 ( \22134 , \22132 , \22133 );
or \U$21758 ( \22135 , \3145 , RIae79ca0_162);
nand \U$21759 ( \22136 , \22134 , \22135 );
not \U$21760 ( \22137 , \22136 );
or \U$21761 ( \22138 , \22131 , \22137 );
nand \U$21762 ( \22139 , \21490 , \4154 );
nand \U$21763 ( \22140 , \22138 , \22139 );
not \U$21764 ( \22141 , \22140 );
not \U$21765 ( \22142 , \13720 );
not \U$21766 ( \22143 , \21398 );
or \U$21767 ( \22144 , \22142 , \22143 );
not \U$21768 ( \22145 , RIae7a240_174);
not \U$21769 ( \22146 , \11441 );
or \U$21770 ( \22147 , \22145 , \22146 );
or \U$21771 ( \22148 , \1158 , RIae7a240_174);
nand \U$21772 ( \22149 , \22147 , \22148 );
nand \U$21773 ( \22150 , \22149 , \9699 );
nand \U$21774 ( \22151 , \22144 , \22150 );
not \U$21775 ( \22152 , \22151 );
not \U$21776 ( \22153 , \22152 );
or \U$21777 ( \22154 , \22141 , \22153 );
or \U$21778 ( \22155 , \22152 , \22140 );
nand \U$21779 ( \22156 , \22154 , \22155 );
not \U$21780 ( \22157 , \2767 );
not \U$21781 ( \22158 , \21391 );
or \U$21782 ( \22159 , \22157 , \22158 );
not \U$21783 ( \22160 , \10584 );
not \U$21784 ( \22161 , \3294 );
or \U$21785 ( \22162 , \22160 , \22161 );
or \U$21786 ( \22163 , \1898 , \10584 );
nand \U$21787 ( \22164 , \22162 , \22163 );
nand \U$21788 ( \22165 , \22164 , \5324 );
nand \U$21789 ( \22166 , \22159 , \22165 );
xor \U$21790 ( \22167 , \22156 , \22166 );
not \U$21791 ( \22168 , \2545 );
not \U$21792 ( \22169 , \21531 );
or \U$21793 ( \22170 , \22168 , \22169 );
and \U$21794 ( \22171 , RIae79778_151, \18384 );
not \U$21795 ( \22172 , RIae79778_151);
and \U$21796 ( \22173 , \22172 , \2230 );
nor \U$21797 ( \22174 , \22171 , \22173 );
nand \U$21798 ( \22175 , \22174 , \11037 );
nand \U$21799 ( \22176 , \22170 , \22175 );
not \U$21800 ( \22177 , \9643 );
not \U$21801 ( \22178 , \21522 );
or \U$21802 ( \22179 , \22177 , \22178 );
xnor \U$21803 ( \22180 , RIae7a3a8_177, \779 );
nand \U$21804 ( \22181 , \22180 , \9622 );
nand \U$21805 ( \22182 , \22179 , \22181 );
nand \U$21806 ( \22183 , \21408 , \9792 );
not \U$21807 ( \22184 , \12184 );
not \U$21808 ( \22185 , \937 );
or \U$21809 ( \22186 , \22184 , \22185 );
not \U$21810 ( \22187 , \9810 );
nand \U$21811 ( \22188 , \22187 , \936 );
nand \U$21812 ( \22189 , \22186 , \22188 );
nand \U$21813 ( \22190 , \22189 , \16135 );
nand \U$21814 ( \22191 , \22183 , \22190 );
xor \U$21815 ( \22192 , \22182 , \22191 );
xor \U$21816 ( \22193 , \22176 , \22192 );
xor \U$21817 ( \22194 , \22167 , \22193 );
not \U$21818 ( \22195 , \1844 );
not \U$21819 ( \22196 , \21478 );
or \U$21820 ( \22197 , \22195 , \22196 );
and \U$21821 ( \22198 , \1969 , \2970 );
not \U$21822 ( \22199 , \1969 );
and \U$21823 ( \22200 , \22199 , RIae79688_149);
nor \U$21824 ( \22201 , \22198 , \22200 );
nand \U$21825 ( \22202 , \22201 , \1821 );
nand \U$21826 ( \22203 , \22197 , \22202 );
not \U$21827 ( \22204 , \2272 );
not \U$21828 ( \22205 , \21467 );
or \U$21829 ( \22206 , \22204 , \22205 );
and \U$21830 ( \22207 , RIae79ac0_158, \13008 );
not \U$21831 ( \22208 , RIae79ac0_158);
and \U$21832 ( \22209 , \22208 , \2089 );
or \U$21833 ( \22210 , \22207 , \22209 );
nand \U$21834 ( \22211 , \22210 , \2252 );
nand \U$21835 ( \22212 , \22206 , \22211 );
xor \U$21836 ( \22213 , \22203 , \22212 );
not \U$21837 ( \22214 , \12233 );
not \U$21838 ( \22215 , \10633 );
not \U$21839 ( \22216 , \991 );
or \U$21840 ( \22217 , \22215 , \22216 );
or \U$21841 ( \22218 , \991 , \14931 );
nand \U$21842 ( \22219 , \22217 , \22218 );
not \U$21843 ( \22220 , \22219 );
or \U$21844 ( \22221 , \22214 , \22220 );
nand \U$21845 ( \22222 , \21498 , \10638 );
nand \U$21846 ( \22223 , \22221 , \22222 );
not \U$21847 ( \22224 , \22223 );
xnor \U$21848 ( \22225 , \22213 , \22224 );
xor \U$21849 ( \22226 , \22194 , \22225 );
not \U$21850 ( \22227 , \21646 );
not \U$21851 ( \22228 , \21631 );
nand \U$21852 ( \22229 , \22228 , \21638 );
not \U$21853 ( \22230 , \22229 );
or \U$21854 ( \22231 , \22227 , \22230 );
buf \U$21855 ( \22232 , \21631 );
nand \U$21856 ( \22233 , \22232 , \21635 );
nand \U$21857 ( \22234 , \22231 , \22233 );
xor \U$21858 ( \22235 , \22226 , \22234 );
not \U$21859 ( \22236 , \1933 );
not \U$21860 ( \22237 , \21357 );
or \U$21861 ( \22238 , \22236 , \22237 );
not \U$21862 ( \22239 , RIae794a8_145);
not \U$21863 ( \22240 , \10608 );
or \U$21864 ( \22241 , \22239 , \22240 );
or \U$21865 ( \22242 , \10905 , RIae794a8_145);
nand \U$21866 ( \22243 , \22241 , \22242 );
nand \U$21867 ( \22244 , \22243 , \1919 );
nand \U$21868 ( \22245 , \22238 , \22244 );
xor \U$21869 ( \22246 , \21335 , \22245 );
not \U$21870 ( \22247 , \11409 );
not \U$21871 ( \22248 , \21373 );
or \U$21872 ( \22249 , \22247 , \22248 );
not \U$21873 ( \22250 , \6207 );
not \U$21874 ( \22251 , \11429 );
or \U$21875 ( \22252 , \22250 , \22251 );
or \U$21876 ( \22253 , \10645 , \6207 );
nand \U$21877 ( \22254 , \22252 , \22253 );
nand \U$21878 ( \22255 , \22254 , \6214 );
nand \U$21879 ( \22256 , \22249 , \22255 );
xor \U$21880 ( \22257 , \22246 , \22256 );
not \U$21881 ( \22258 , \21578 );
not \U$21882 ( \22259 , \21572 );
or \U$21883 ( \22260 , \22258 , \22259 );
nand \U$21884 ( \22261 , \21571 , \21561 );
nand \U$21885 ( \22262 , \22260 , \22261 );
not \U$21886 ( \22263 , \22262 );
xor \U$21887 ( \22264 , \22257 , \22263 );
xor \U$21888 ( \22265 , \21450 , \21460 );
and \U$21889 ( \22266 , \22265 , \21471 );
and \U$21890 ( \22267 , \21450 , \21460 );
or \U$21891 ( \22268 , \22266 , \22267 );
xor \U$21892 ( \22269 , \21765 , \21777 );
and \U$21893 ( \22270 , \22269 , \21783 );
and \U$21894 ( \22271 , \21765 , \21777 );
or \U$21895 ( \22272 , \22270 , \22271 );
xor \U$21896 ( \22273 , \22268 , \22272 );
xor \U$21897 ( \22274 , \21730 , \21740 );
and \U$21898 ( \22275 , \22274 , \21753 );
and \U$21899 ( \22276 , \21730 , \21740 );
or \U$21900 ( \22277 , \22275 , \22276 );
xor \U$21901 ( \22278 , \22273 , \22277 );
xnor \U$21902 ( \22279 , \22264 , \22278 );
xor \U$21903 ( \22280 , \22235 , \22279 );
xor \U$21904 ( \22281 , \22130 , \22280 );
or \U$21905 ( \22282 , \21660 , \21650 );
nand \U$21906 ( \22283 , \22282 , \21655 );
nand \U$21907 ( \22284 , \21660 , \21650 );
nand \U$21908 ( \22285 , \22283 , \22284 );
xor \U$21909 ( \22286 , \22281 , \22285 );
xor \U$21910 ( \22287 , \22125 , \22286 );
nand \U$21911 ( \22288 , \21806 , \21671 );
nand \U$21912 ( \22289 , \22288 , \21674 );
xnor \U$21913 ( \22290 , \22287 , \22289 );
not \U$21914 ( \22291 , \22290 );
or \U$21915 ( \22292 , \22119 , \22291 );
or \U$21916 ( \22293 , \22118 , \22290 );
nand \U$21917 ( \22294 , \22292 , \22293 );
not \U$21918 ( \22295 , \22294 );
and \U$21919 ( \22296 , \21620 , \21614 );
or \U$21920 ( \22297 , \22296 , \21625 );
or \U$21921 ( \22298 , \21614 , \21620 );
nand \U$21922 ( \22299 , \22297 , \22298 );
not \U$21923 ( \22300 , \22299 );
not \U$21924 ( \22301 , \22300 );
and \U$21925 ( \22302 , \22295 , \22301 );
and \U$21926 ( \22303 , \22294 , \22300 );
nor \U$21927 ( \22304 , \22302 , \22303 );
nor \U$21928 ( \22305 , \21824 , \22304 );
not \U$21929 ( \22306 , \22028 );
not \U$21930 ( \22307 , \22005 );
or \U$21931 ( \22308 , \22306 , \22307 );
not \U$21932 ( \22309 , \22004 );
not \U$21933 ( \22310 , \22025 );
or \U$21934 ( \22311 , \22309 , \22310 );
nand \U$21935 ( \22312 , \22311 , \21897 );
nand \U$21936 ( \22313 , \22308 , \22312 );
not \U$21937 ( \22314 , \21828 );
not \U$21938 ( \22315 , \22314 );
not \U$21939 ( \22316 , \21836 );
or \U$21940 ( \22317 , \22315 , \22316 );
nand \U$21941 ( \22318 , \22317 , \21841 );
nand \U$21942 ( \22319 , \21833 , \21835 , \21828 );
nand \U$21943 ( \22320 , \22318 , \22319 );
not \U$21944 ( \22321 , \22257 );
not \U$21945 ( \22322 , \22262 );
or \U$21946 ( \22323 , \22321 , \22322 );
not \U$21947 ( \22324 , \22278 );
nand \U$21948 ( \22325 , \22323 , \22324 );
not \U$21949 ( \22326 , \22257 );
nand \U$21950 ( \22327 , \22326 , \22263 );
nand \U$21951 ( \22328 , \22325 , \22327 );
and \U$21952 ( \22329 , \22320 , \22328 );
not \U$21953 ( \22330 , \22320 );
not \U$21954 ( \22331 , \22328 );
and \U$21955 ( \22332 , \22330 , \22331 );
nor \U$21956 ( \22333 , \22329 , \22332 );
xnor \U$21957 ( \22334 , \22313 , \22333 );
or \U$21958 ( \22335 , \21954 , \21943 );
not \U$21959 ( \22336 , \22335 );
not \U$21960 ( \22337 , \21967 );
or \U$21961 ( \22338 , \22336 , \22337 );
nand \U$21962 ( \22339 , \21954 , \21943 );
nand \U$21963 ( \22340 , \22338 , \22339 );
not \U$21964 ( \22341 , \1072 );
not \U$21965 ( \22342 , \9438 );
not \U$21966 ( \22343 , RIae78e90_132);
and \U$21967 ( \22344 , \22342 , \22343 );
and \U$21968 ( \22345 , \9438 , RIae78e90_132);
nor \U$21969 ( \22346 , \22344 , \22345 );
not \U$21970 ( \22347 , \22346 );
or \U$21971 ( \22348 , \22341 , \22347 );
nand \U$21972 ( \22349 , \21952 , \1086 );
nand \U$21973 ( \22350 , \22348 , \22349 );
not \U$21974 ( \22351 , \9947 );
not \U$21975 ( \22352 , RIae79070_136);
not \U$21976 ( \22353 , \6230 );
not \U$21977 ( \22354 , \22353 );
or \U$21978 ( \22355 , \22352 , \22354 );
not \U$21979 ( \22356 , \9298 );
or \U$21980 ( \22357 , \22356 , RIae79070_136);
nand \U$21981 ( \22358 , \22355 , \22357 );
not \U$21982 ( \22359 , \22358 );
or \U$21983 ( \22360 , \22351 , \22359 );
nand \U$21984 ( \22361 , \21929 , \1062 );
nand \U$21985 ( \22362 , \22360 , \22361 );
xor \U$21986 ( \22363 , \22350 , \22362 );
not \U$21987 ( \22364 , \5124 );
and \U$21988 ( \22365 , RIae78f80_134, \12707 );
not \U$21989 ( \22366 , RIae78f80_134);
and \U$21990 ( \22367 , \22366 , \21743 );
or \U$21991 ( \22368 , \22365 , \22367 );
not \U$21992 ( \22369 , \22368 );
or \U$21993 ( \22370 , \22364 , \22369 );
nand \U$21994 ( \22371 , \21912 , \796 );
nand \U$21995 ( \22372 , \22370 , \22371 );
xor \U$21996 ( \22373 , \22363 , \22372 );
xor \U$21997 ( \22374 , \22340 , \22373 );
not \U$21998 ( \22375 , \1919 );
not \U$21999 ( \22376 , RIae794a8_145);
not \U$22000 ( \22377 , \3098 );
or \U$22001 ( \22378 , \22376 , \22377 );
not \U$22002 ( \22379 , RIae794a8_145);
nand \U$22003 ( \22380 , \22379 , \1740 );
nand \U$22004 ( \22381 , \22378 , \22380 );
not \U$22005 ( \22382 , \22381 );
or \U$22006 ( \22383 , \22375 , \22382 );
nand \U$22007 ( \22384 , \22243 , \2457 );
nand \U$22008 ( \22385 , \22383 , \22384 );
not \U$22009 ( \22386 , \22385 );
not \U$22010 ( \22387 , \22386 );
not \U$22011 ( \22388 , \6214 );
not \U$22012 ( \22389 , RIae79ef8_167);
not \U$22013 ( \22390 , \22389 );
not \U$22014 ( \22391 , \1118 );
or \U$22015 ( \22392 , \22390 , \22391 );
or \U$22016 ( \22393 , \12801 , \22389 );
nand \U$22017 ( \22394 , \22392 , \22393 );
not \U$22018 ( \22395 , \22394 );
or \U$22019 ( \22396 , \22388 , \22395 );
nand \U$22020 ( \22397 , \15989 , \22254 );
nand \U$22021 ( \22398 , \22396 , \22397 );
not \U$22022 ( \22399 , \22398 );
or \U$22023 ( \22400 , \22387 , \22399 );
or \U$22024 ( \22401 , \22398 , \22386 );
nand \U$22025 ( \22402 , \22400 , \22401 );
not \U$22026 ( \22403 , \5049 );
not \U$22027 ( \22404 , RIae79d90_164);
not \U$22028 ( \22405 , \1186 );
or \U$22029 ( \22406 , \22404 , \22405 );
or \U$22030 ( \22407 , \3539 , RIae79d90_164);
nand \U$22031 ( \22408 , \22406 , \22407 );
not \U$22032 ( \22409 , \22408 );
or \U$22033 ( \22410 , \22403 , \22409 );
nand \U$22034 ( \22411 , \21963 , \5040 );
nand \U$22035 ( \22412 , \22410 , \22411 );
xor \U$22036 ( \22413 , \22402 , \22412 );
xor \U$22037 ( \22414 , \22374 , \22413 );
not \U$22038 ( \22415 , \22414 );
not \U$22039 ( \22416 , \22415 );
not \U$22040 ( \22417 , \21999 );
nand \U$22041 ( \22418 , \21932 , \21968 );
not \U$22042 ( \22419 , \22418 );
or \U$22043 ( \22420 , \22417 , \22419 );
not \U$22044 ( \22421 , \21968 );
nand \U$22045 ( \22422 , \22421 , \21933 );
nand \U$22046 ( \22423 , \22420 , \22422 );
xor \U$22047 ( \22424 , \21450 , \21460 );
and \U$22048 ( \22425 , \22424 , \21471 );
and \U$22049 ( \22426 , \21450 , \21460 );
or \U$22050 ( \22427 , \22425 , \22426 );
not \U$22051 ( \22428 , \22427 );
not \U$22052 ( \22429 , \22272 );
or \U$22053 ( \22430 , \22428 , \22429 );
not \U$22054 ( \22431 , \22277 );
nand \U$22055 ( \22432 , \22430 , \22431 );
not \U$22056 ( \22433 , \22272 );
not \U$22057 ( \22434 , \22427 );
nand \U$22058 ( \22435 , \22433 , \22434 );
nand \U$22059 ( \22436 , \22432 , \22435 );
xnor \U$22060 ( \22437 , \22423 , \22436 );
not \U$22061 ( \22438 , \22437 );
not \U$22062 ( \22439 , \22438 );
or \U$22063 ( \22440 , \22416 , \22439 );
nand \U$22064 ( \22441 , \22437 , \22414 );
nand \U$22065 ( \22442 , \22440 , \22441 );
not \U$22066 ( \22443 , \21895 );
not \U$22067 ( \22444 , \21888 );
or \U$22068 ( \22445 , \22443 , \22444 );
nand \U$22069 ( \22446 , \22445 , \21882 );
not \U$22070 ( \22447 , \21888 );
nand \U$22071 ( \22448 , \22447 , \21896 );
nand \U$22072 ( \22449 , \22446 , \22448 );
not \U$22073 ( \22450 , \22013 );
not \U$22074 ( \22451 , \22450 );
not \U$22075 ( \22452 , \22451 );
not \U$22076 ( \22453 , \22018 );
or \U$22077 ( \22454 , \22452 , \22453 );
not \U$22078 ( \22455 , \22450 );
not \U$22079 ( \22456 , \22018 );
not \U$22080 ( \22457 , \22456 );
or \U$22081 ( \22458 , \22455 , \22457 );
nand \U$22082 ( \22459 , \22458 , \22024 );
nand \U$22083 ( \22460 , \22454 , \22459 );
xor \U$22084 ( \22461 , \22449 , \22460 );
not \U$22085 ( \22462 , \21931 );
not \U$22086 ( \22463 , \21906 );
nand \U$22087 ( \22464 , \22463 , \21919 );
not \U$22088 ( \22465 , \22464 );
or \U$22089 ( \22466 , \22462 , \22465 );
nand \U$22090 ( \22467 , \21916 , \21906 );
nand \U$22091 ( \22468 , \22466 , \22467 );
xor \U$22092 ( \22469 , \21860 , \21870 );
and \U$22093 ( \22470 , \22469 , \21881 );
and \U$22094 ( \22471 , \21860 , \21870 );
or \U$22095 ( \22472 , \22470 , \22471 );
xor \U$22096 ( \22473 , \22468 , \22472 );
not \U$22097 ( \22474 , \22212 );
not \U$22098 ( \22475 , \22203 );
not \U$22099 ( \22476 , \22475 );
not \U$22100 ( \22477 , \22223 );
or \U$22101 ( \22478 , \22476 , \22477 );
or \U$22102 ( \22479 , \22223 , \22475 );
nand \U$22103 ( \22480 , \22478 , \22479 );
not \U$22104 ( \22481 , \22480 );
or \U$22105 ( \22482 , \22474 , \22481 );
not \U$22106 ( \22483 , \22224 );
nand \U$22107 ( \22484 , \22483 , \22203 );
nand \U$22108 ( \22485 , \22482 , \22484 );
xor \U$22109 ( \22486 , \22473 , \22485 );
xor \U$22110 ( \22487 , \22461 , \22486 );
xor \U$22111 ( \22488 , \22442 , \22487 );
xor \U$22112 ( \22489 , \22167 , \22193 );
and \U$22113 ( \22490 , \22489 , \22225 );
and \U$22114 ( \22491 , \22167 , \22193 );
or \U$22115 ( \22492 , \22490 , \22491 );
not \U$22116 ( \22493 , \22166 );
not \U$22117 ( \22494 , \22156 );
or \U$22118 ( \22495 , \22493 , \22494 );
nand \U$22119 ( \22496 , \22151 , \22140 );
nand \U$22120 ( \22497 , \22495 , \22496 );
not \U$22121 ( \22498 , \22497 );
nand \U$22122 ( \22499 , \22192 , \22176 );
not \U$22123 ( \22500 , \22190 );
not \U$22124 ( \22501 , \22183 );
or \U$22125 ( \22502 , \22500 , \22501 );
nand \U$22126 ( \22503 , \22502 , \22182 );
and \U$22127 ( \22504 , \22499 , \22503 );
not \U$22128 ( \22505 , \22504 );
or \U$22129 ( \22506 , \22498 , \22505 );
or \U$22130 ( \22507 , \22504 , \22497 );
nand \U$22131 ( \22508 , \22506 , \22507 );
not \U$22132 ( \22509 , \22508 );
xor \U$22133 ( \22510 , \21978 , \21987 );
and \U$22134 ( \22511 , \22510 , \21998 );
and \U$22135 ( \22512 , \21978 , \21987 );
or \U$22136 ( \22513 , \22511 , \22512 );
not \U$22137 ( \22514 , \22513 );
not \U$22138 ( \22515 , \22514 );
and \U$22139 ( \22516 , \22509 , \22515 );
and \U$22140 ( \22517 , \22508 , \22514 );
nor \U$22141 ( \22518 , \22516 , \22517 );
not \U$22142 ( \22519 , \22518 );
xor \U$22143 ( \22520 , \22492 , \22519 );
xor \U$22144 ( \22521 , \21335 , \22245 );
and \U$22145 ( \22522 , \22521 , \22256 );
and \U$22146 ( \22523 , \21335 , \22245 );
or \U$22147 ( \22524 , \22522 , \22523 );
not \U$22148 ( \22525 , \997 );
not \U$22149 ( \22526 , \5722 );
or \U$22150 ( \22527 , \22525 , \22526 );
nand \U$22151 ( \22528 , \12700 , RIae79160_138);
nand \U$22152 ( \22529 , \22527 , \22528 );
and \U$22153 ( \22530 , \10451 , \22529 );
and \U$22154 ( \22531 , \21904 , \1008 );
nor \U$22155 ( \22532 , \22530 , \22531 );
not \U$22156 ( \22533 , \1501 );
not \U$22157 ( \22534 , RIae79250_140);
not \U$22158 ( \22535 , \4960 );
or \U$22159 ( \22536 , \22534 , \22535 );
nand \U$22160 ( \22537 , \17009 , \1503 );
nand \U$22161 ( \22538 , \22536 , \22537 );
not \U$22162 ( \22539 , \22538 );
or \U$22163 ( \22540 , \22533 , \22539 );
nand \U$22164 ( \22541 , \21856 , \1499 );
nand \U$22165 ( \22542 , \22540 , \22541 );
xor \U$22166 ( \22543 , \22532 , \22542 );
not \U$22167 ( \22544 , \1910 );
not \U$22168 ( \22545 , \21877 );
or \U$22169 ( \22546 , \22544 , \22545 );
and \U$22170 ( \22547 , RIae793b8_143, \3207 );
not \U$22171 ( \22548 , RIae793b8_143);
and \U$22172 ( \22549 , \22548 , \9830 );
nor \U$22173 ( \22550 , \22547 , \22549 );
nand \U$22174 ( \22551 , \22550 , \1864 );
nand \U$22175 ( \22552 , \22546 , \22551 );
xnor \U$22176 ( \22553 , \22543 , \22552 );
xor \U$22177 ( \22554 , \22524 , \22553 );
not \U$22178 ( \22555 , \929 );
not \U$22179 ( \22556 , \1286 );
not \U$22180 ( \22557 , \15488 );
not \U$22181 ( \22558 , \22557 );
or \U$22182 ( \22559 , \22556 , \22558 );
buf \U$22183 ( \22560 , \10937 );
nand \U$22184 ( \22561 , \22560 , RIae78bc0_126);
nand \U$22185 ( \22562 , \22559 , \22561 );
not \U$22186 ( \22563 , \22562 );
or \U$22187 ( \22564 , \22555 , \22563 );
nand \U$22188 ( \22565 , \21941 , \952 );
nand \U$22189 ( \22566 , \22564 , \22565 );
not \U$22190 ( \22567 , \2096 );
xor \U$22191 ( \22568 , RIae78b48_125, \9607 );
not \U$22192 ( \22569 , \22568 );
or \U$22193 ( \22570 , \22567 , \22569 );
nand \U$22194 ( \22571 , \22063 , \893 );
nand \U$22195 ( \22572 , \22570 , \22571 );
not \U$22196 ( \22573 , \22572 );
xor \U$22197 ( \22574 , \22566 , \22573 );
not \U$22198 ( \22575 , \11400 );
not \U$22199 ( \22576 , \22219 );
or \U$22200 ( \22577 , \22575 , \22576 );
nand \U$22201 ( \22578 , \16358 , RIae7a510_180);
nand \U$22202 ( \22579 , \22577 , \22578 );
xnor \U$22203 ( \22580 , \22574 , \22579 );
xor \U$22204 ( \22581 , \22554 , \22580 );
xnor \U$22205 ( \22582 , \22520 , \22581 );
xor \U$22206 ( \22583 , \22488 , \22582 );
xor \U$22207 ( \22584 , \22334 , \22583 );
not \U$22208 ( \22585 , \22030 );
not \U$22209 ( \22586 , \22585 );
not \U$22210 ( \22587 , \21849 );
or \U$22211 ( \22588 , \22586 , \22587 );
not \U$22212 ( \22589 , \21842 );
nand \U$22213 ( \22590 , \22589 , \21848 );
nand \U$22214 ( \22591 , \22588 , \22590 );
xor \U$22215 ( \22592 , \22584 , \22591 );
buf \U$22216 ( \22593 , \22125 );
not \U$22217 ( \22594 , \22593 );
buf \U$22218 ( \22595 , \22286 );
not \U$22219 ( \22596 , \22595 );
or \U$22220 ( \22597 , \22594 , \22596 );
or \U$22221 ( \22598 , \22595 , \22593 );
nand \U$22222 ( \22599 , \22598 , \22289 );
nand \U$22223 ( \22600 , \22597 , \22599 );
xor \U$22224 ( \22601 , \22592 , \22600 );
xor \U$22225 ( \22602 , \22130 , \22280 );
and \U$22226 ( \22603 , \22602 , \22285 );
and \U$22227 ( \22604 , \22130 , \22280 );
or \U$22228 ( \22605 , \22603 , \22604 );
xor \U$22229 ( \22606 , \22226 , \22234 );
and \U$22230 ( \22607 , \22606 , \22279 );
and \U$22231 ( \22608 , \22226 , \22234 );
or \U$22232 ( \22609 , \22607 , \22608 );
not \U$22233 ( \22610 , \2252 );
xor \U$22234 ( \22611 , \11512 , RIae79ac0_158);
not \U$22235 ( \22612 , \22611 );
or \U$22236 ( \22613 , \22610 , \22612 );
nand \U$22237 ( \22614 , \22210 , \2272 );
nand \U$22238 ( \22615 , \22613 , \22614 );
nand \U$22239 ( \22616 , \22050 , \12680 );
not \U$22240 ( \22617 , \2183 );
not \U$22241 ( \22618 , \1808 );
or \U$22242 ( \22619 , \22617 , \22618 );
or \U$22243 ( \22620 , \1808 , \2183 );
nand \U$22244 ( \22621 , \22619 , \22620 );
nand \U$22245 ( \22622 , \22621 , \10223 );
and \U$22246 ( \22623 , \22616 , \22622 );
not \U$22247 ( \22624 , \22054 );
xnor \U$22248 ( \22625 , \22624 , \22055 );
not \U$22249 ( \22626 , \22625 );
not \U$22250 ( \22627 , \22065 );
or \U$22251 ( \22628 , \22626 , \22627 );
nand \U$22252 ( \22629 , \21106 , \22624 , RIae78b48_125);
nand \U$22253 ( \22630 , \22628 , \22629 );
xnor \U$22254 ( \22631 , \22623 , \22630 );
xor \U$22255 ( \22632 , \22615 , \22631 );
not \U$22256 ( \22633 , \1822 );
not \U$22257 ( \22634 , RIae79688_149);
not \U$22258 ( \22635 , \4112 );
or \U$22259 ( \22636 , \22634 , \22635 );
nand \U$22260 ( \22637 , \5115 , \3147 );
nand \U$22261 ( \22638 , \22636 , \22637 );
not \U$22262 ( \22639 , \22638 );
or \U$22263 ( \22640 , \22633 , \22639 );
nand \U$22264 ( \22641 , \22201 , \1844 );
nand \U$22265 ( \22642 , \22640 , \22641 );
not \U$22266 ( \22643 , \2011 );
and \U$22267 ( \22644 , RIae79610_148, \17596 );
not \U$22268 ( \22645 , RIae79610_148);
and \U$22269 ( \22646 , \22645 , \4100 );
nor \U$22270 ( \22647 , \22644 , \22646 );
not \U$22271 ( \22648 , \22647 );
or \U$22272 ( \22649 , \22643 , \22648 );
nand \U$22273 ( \22650 , \21868 , \2063 );
nand \U$22274 ( \22651 , \22649 , \22650 );
not \U$22275 ( \22652 , \22651 );
not \U$22276 ( \22653 , \6276 );
not \U$22277 ( \22654 , \22136 );
or \U$22278 ( \22655 , \22653 , \22654 );
and \U$22279 ( \22656 , RIae79ca0_162, \2025 );
not \U$22280 ( \22657 , RIae79ca0_162);
and \U$22281 ( \22658 , \22657 , \2030 );
nor \U$22282 ( \22659 , \22656 , \22658 );
nand \U$22283 ( \22660 , \4853 , \22659 );
nand \U$22284 ( \22661 , \22655 , \22660 );
not \U$22285 ( \22662 , \22661 );
not \U$22286 ( \22663 , \22662 );
or \U$22287 ( \22664 , \22652 , \22663 );
or \U$22288 ( \22665 , \22662 , \22651 );
nand \U$22289 ( \22666 , \22664 , \22665 );
xor \U$22290 ( \22667 , \22642 , \22666 );
xor \U$22291 ( \22668 , \22632 , \22667 );
not \U$22292 ( \22669 , \22067 );
not \U$22293 ( \22670 , \22669 );
not \U$22294 ( \22671 , \22077 );
or \U$22295 ( \22672 , \22670 , \22671 );
nand \U$22296 ( \22673 , \22672 , \22069 );
xor \U$22297 ( \22674 , \22668 , \22673 );
not \U$22298 ( \22675 , \13657 );
nand \U$22299 ( \22676 , \22675 , RIae78b48_125);
not \U$22300 ( \22677 , \9518 );
xor \U$22301 ( \22678 , RIae79fe8_169, \854 );
not \U$22302 ( \22679 , \22678 );
or \U$22303 ( \22680 , \22677 , \22679 );
nand \U$22304 ( \22681 , \21996 , \9499 );
nand \U$22305 ( \22682 , \22680 , \22681 );
xor \U$22306 ( \22683 , \22676 , \22682 );
not \U$22307 ( \22684 , \2450 );
and \U$22308 ( \22685 , RIae79778_151, \2207 );
not \U$22309 ( \22686 , RIae79778_151);
and \U$22310 ( \22687 , \22686 , \3051 );
nor \U$22311 ( \22688 , \22685 , \22687 );
not \U$22312 ( \22689 , \22688 );
or \U$22313 ( \22690 , \22684 , \22689 );
nand \U$22314 ( \22691 , \22174 , \2433 );
nand \U$22315 ( \22692 , \22690 , \22691 );
xnor \U$22316 ( \22693 , \22683 , \22692 );
not \U$22317 ( \22694 , \22693 );
not \U$22318 ( \22695 , \22694 );
not \U$22319 ( \22696 , \9699 );
not \U$22320 ( \22697 , RIae7a240_174);
not \U$22321 ( \22698 , \3999 );
or \U$22322 ( \22699 , \22697 , \22698 );
or \U$22323 ( \22700 , \1142 , RIae7a240_174);
nand \U$22324 ( \22701 , \22699 , \22700 );
not \U$22325 ( \22702 , \22701 );
or \U$22326 ( \22703 , \22696 , \22702 );
nand \U$22327 ( \22704 , \22149 , \13130 );
nand \U$22328 ( \22705 , \22703 , \22704 );
not \U$22329 ( \22706 , \2519 );
not \U$22330 ( \22707 , \2521 );
not \U$22331 ( \22708 , \10567 );
or \U$22332 ( \22709 , \22707 , \22708 );
nand \U$22333 ( \22710 , \10570 , RIae797f0_152);
nand \U$22334 ( \22711 , \22709 , \22710 );
not \U$22335 ( \22712 , \22711 );
or \U$22336 ( \22713 , \22706 , \22712 );
nand \U$22337 ( \22714 , \21983 , \1988 );
nand \U$22338 ( \22715 , \22713 , \22714 );
not \U$22339 ( \22716 , \10807 );
not \U$22340 ( \22717 , \21976 );
or \U$22341 ( \22718 , \22716 , \22717 );
and \U$22342 ( \22719 , RIae798e0_154, \2305 );
not \U$22343 ( \22720 , RIae798e0_154);
and \U$22344 ( \22721 , \22720 , \2309 );
or \U$22345 ( \22722 , \22719 , \22721 );
nand \U$22346 ( \22723 , \22722 , \2322 );
nand \U$22347 ( \22724 , \22718 , \22723 );
and \U$22348 ( \22725 , \22715 , \22724 );
not \U$22349 ( \22726 , \22715 );
not \U$22350 ( \22727 , \22724 );
and \U$22351 ( \22728 , \22726 , \22727 );
nor \U$22352 ( \22729 , \22725 , \22728 );
xor \U$22353 ( \22730 , \22705 , \22729 );
not \U$22354 ( \22731 , \22730 );
not \U$22355 ( \22732 , \22731 );
or \U$22356 ( \22733 , \22695 , \22732 );
nand \U$22357 ( \22734 , \22693 , \22730 );
nand \U$22358 ( \22735 , \22733 , \22734 );
not \U$22359 ( \22736 , \2776 );
and \U$22360 ( \22737 , RIae79c28_161, \4458 );
not \U$22361 ( \22738 , RIae79c28_161);
and \U$22362 ( \22739 , \22738 , \5162 );
or \U$22363 ( \22740 , \22737 , \22739 );
not \U$22364 ( \22741 , \22740 );
or \U$22365 ( \22742 , \22736 , \22741 );
nand \U$22366 ( \22743 , \22164 , \2767 );
nand \U$22367 ( \22744 , \22742 , \22743 );
not \U$22368 ( \22745 , \9622 );
not \U$22369 ( \22746 , RIae7a3a8_177);
not \U$22370 ( \22747 , \827 );
or \U$22371 ( \22748 , \22746 , \22747 );
or \U$22372 ( \22749 , \4413 , RIae7a3a8_177);
nand \U$22373 ( \22750 , \22748 , \22749 );
not \U$22374 ( \22751 , \22750 );
or \U$22375 ( \22752 , \22745 , \22751 );
nand \U$22376 ( \22753 , \22180 , \11014 );
nand \U$22377 ( \22754 , \22752 , \22753 );
xor \U$22378 ( \22755 , \22744 , \22754 );
and \U$22379 ( \22756 , RIae7a2b8_175, \15675 );
not \U$22380 ( \22757 , RIae7a2b8_175);
and \U$22381 ( \22758 , \22757 , \16589 );
nor \U$22382 ( \22759 , \22756 , \22758 );
not \U$22383 ( \22760 , \22759 );
not \U$22384 ( \22761 , \9814 );
or \U$22385 ( \22762 , \22760 , \22761 );
nand \U$22386 ( \22763 , \22189 , \9792 );
nand \U$22387 ( \22764 , \22762 , \22763 );
xor \U$22388 ( \22765 , \22755 , \22764 );
not \U$22389 ( \22766 , \22765 );
and \U$22390 ( \22767 , \22735 , \22766 );
not \U$22391 ( \22768 , \22735 );
and \U$22392 ( \22769 , \22768 , \22765 );
nor \U$22393 ( \22770 , \22767 , \22769 );
xor \U$22394 ( \22771 , \22674 , \22770 );
xor \U$22395 ( \22772 , \22078 , \22085 );
and \U$22396 ( \22773 , \22772 , \22090 );
and \U$22397 ( \22774 , \22078 , \22085 );
or \U$22398 ( \22775 , \22773 , \22774 );
xnor \U$22399 ( \22776 , \22771 , \22775 );
xor \U$22400 ( \22777 , \22609 , \22776 );
not \U$22401 ( \22778 , \22107 );
not \U$22402 ( \22779 , \22099 );
or \U$22403 ( \22780 , \22778 , \22779 );
nand \U$22404 ( \22781 , \22780 , \22100 );
xor \U$22405 ( \22782 , \22777 , \22781 );
xor \U$22406 ( \22783 , \22605 , \22782 );
not \U$22407 ( \22784 , \22113 );
not \U$22408 ( \22785 , \22035 );
or \U$22409 ( \22786 , \22784 , \22785 );
not \U$22410 ( \22787 , \22034 );
not \U$22411 ( \22788 , \22112 );
or \U$22412 ( \22789 , \22787 , \22788 );
not \U$22413 ( \22790 , \22042 );
nand \U$22414 ( \22791 , \22789 , \22790 );
nand \U$22415 ( \22792 , \22786 , \22791 );
xor \U$22416 ( \22793 , \22783 , \22792 );
xnor \U$22417 ( \22794 , \22601 , \22793 );
not \U$22418 ( \22795 , \22299 );
not \U$22419 ( \22796 , \22294 );
or \U$22420 ( \22797 , \22795 , \22796 );
not \U$22421 ( \22798 , \22118 );
nand \U$22422 ( \22799 , \22798 , \22290 );
nand \U$22423 ( \22800 , \22797 , \22799 );
nand \U$22424 ( \22801 , \22794 , \22800 );
not \U$22425 ( \22802 , \22801 );
nor \U$22426 ( \22803 , \22305 , \22802 );
not \U$22427 ( \22804 , \21303 );
buf \U$22428 ( \22805 , \20785 );
xor \U$22429 ( \22806 , \21293 , \22805 );
nand \U$22430 ( \22807 , \22806 , \21081 );
not \U$22431 ( \22808 , \22807 );
or \U$22432 ( \22809 , \22804 , \22808 );
or \U$22433 ( \22810 , \22806 , \21081 );
nand \U$22434 ( \22811 , \22809 , \22810 );
xnor \U$22435 ( \22812 , \21819 , \21626 );
nand \U$22436 ( \22813 , \22811 , \22812 );
and \U$22437 ( \22814 , \21306 , \22803 , \22813 );
not \U$22438 ( \22815 , \22814 );
not \U$22439 ( \22816 , \22815 );
nand \U$22440 ( \22817 , \15931 , \20772 , \22816 );
not \U$22441 ( \22818 , \22817 );
not \U$22442 ( \22819 , \2602 );
not \U$22443 ( \22820 , \5971 );
not \U$22444 ( \22821 , RIae79520_146);
and \U$22445 ( \22822 , \22820 , \22821 );
and \U$22446 ( \22823 , \3055 , RIae79520_146);
nor \U$22447 ( \22824 , \22822 , \22823 );
not \U$22448 ( \22825 , \22824 );
or \U$22449 ( \22826 , \22819 , \22825 );
nand \U$22450 ( \22827 , \6076 , \2610 );
nand \U$22451 ( \22828 , \22826 , \22827 );
not \U$22452 ( \22829 , \2767 );
not \U$22453 ( \22830 , RIae79c28_161);
not \U$22454 ( \22831 , \2169 );
or \U$22455 ( \22832 , \22830 , \22831 );
nand \U$22456 ( \22833 , \5191 , \10584 );
nand \U$22457 ( \22834 , \22832 , \22833 );
not \U$22458 ( \22835 , \22834 );
or \U$22459 ( \22836 , \22829 , \22835 );
nand \U$22460 ( \22837 , \6114 , \5324 );
nand \U$22461 ( \22838 , \22836 , \22837 );
nor \U$22462 ( \22839 , \22828 , \22838 );
buf \U$22463 ( \22840 , \22839 );
not \U$22464 ( \22841 , \2272 );
not \U$22465 ( \22842 , RIae79ac0_158);
not \U$22466 ( \22843 , \3071 );
or \U$22467 ( \22844 , \22842 , \22843 );
nand \U$22468 ( \22845 , \9501 , \2268 );
nand \U$22469 ( \22846 , \22844 , \22845 );
not \U$22470 ( \22847 , \22846 );
or \U$22471 ( \22848 , \22841 , \22847 );
nand \U$22472 ( \22849 , \6123 , \3015 );
nand \U$22473 ( \22850 , \22848 , \22849 );
not \U$22474 ( \22851 , \22850 );
or \U$22475 ( \22852 , \22840 , \22851 );
nand \U$22476 ( \22853 , \22828 , \22838 );
nand \U$22477 ( \22854 , \22852 , \22853 );
not \U$22478 ( \22855 , \1919 );
xor \U$22479 ( \22856 , \3146 , RIae794a8_145);
not \U$22480 ( \22857 , \22856 );
or \U$22481 ( \22858 , \22855 , \22857 );
and \U$22482 ( \22859 , RIae794a8_145, \4458 );
not \U$22483 ( \22860 , RIae794a8_145);
and \U$22484 ( \22861 , \22860 , \4198 );
or \U$22485 ( \22862 , \22859 , \22861 );
nand \U$22486 ( \22863 , \22862 , \9828 );
nand \U$22487 ( \22864 , \22858 , \22863 );
not \U$22488 ( \22865 , \22864 );
not \U$22489 ( \22866 , \6214 );
not \U$22490 ( \22867 , \6209 );
or \U$22491 ( \22868 , \22866 , \22867 );
not \U$22492 ( \22869 , RIae79ef8_167);
not \U$22493 ( \22870 , \16395 );
or \U$22494 ( \22871 , \22869 , \22870 );
or \U$22495 ( \22872 , \834 , RIae79ef8_167);
nand \U$22496 ( \22873 , \22871 , \22872 );
nand \U$22497 ( \22874 , \22873 , \6201 );
nand \U$22498 ( \22875 , \22868 , \22874 );
not \U$22499 ( \22876 , \22875 );
or \U$22500 ( \22877 , \22865 , \22876 );
not \U$22501 ( \22878 , \4842 );
not \U$22502 ( \22879 , RIae79ca0_162);
not \U$22503 ( \22880 , \3443 );
or \U$22504 ( \22881 , \22879 , \22880 );
not \U$22505 ( \22882 , \5958 );
nand \U$22506 ( \22883 , \22882 , \10892 );
nand \U$22507 ( \22884 , \22881 , \22883 );
not \U$22508 ( \22885 , \22884 );
or \U$22509 ( \22886 , \22878 , \22885 );
nand \U$22510 ( \22887 , \6275 , \4853 );
nand \U$22511 ( \22888 , \22886 , \22887 );
not \U$22512 ( \22889 , \22888 );
nand \U$22513 ( \22890 , \22877 , \22889 );
not \U$22514 ( \22891 , \22864 );
not \U$22515 ( \22892 , \22875 );
nand \U$22516 ( \22893 , \22891 , \22892 );
nand \U$22517 ( \22894 , \22890 , \22893 );
and \U$22518 ( \22895 , RIae79070_136, \1970 );
not \U$22519 ( \22896 , RIae79070_136);
and \U$22520 ( \22897 , \22896 , \1973 );
nor \U$22521 ( \22898 , \22895 , \22897 );
not \U$22522 ( \22899 , \22898 );
not \U$22523 ( \22900 , \1203 );
and \U$22524 ( \22901 , \22899 , \22900 );
and \U$22525 ( \22902 , RIae79070_136, \1860 );
not \U$22526 ( \22903 , RIae79070_136);
and \U$22527 ( \22904 , \22903 , \2385 );
or \U$22528 ( \22905 , \22902 , \22904 );
and \U$22529 ( \22906 , \22905 , \1062 );
nor \U$22530 ( \22907 , \22901 , \22906 );
not \U$22531 ( \22908 , \2157 );
and \U$22532 ( \22909 , RIae79160_138, \2358 );
not \U$22533 ( \22910 , RIae79160_138);
and \U$22534 ( \22911 , \22910 , \5115 );
or \U$22535 ( \22912 , \22909 , \22911 );
not \U$22536 ( \22913 , \22912 );
or \U$22537 ( \22914 , \22908 , \22913 );
and \U$22538 ( \22915 , RIae79160_138, \2786 );
not \U$22539 ( \22916 , RIae79160_138);
not \U$22540 ( \22917 , \14439 );
and \U$22541 ( \22918 , \22916 , \22917 );
or \U$22542 ( \22919 , \22915 , \22918 );
nand \U$22543 ( \22920 , \22919 , \1013 );
nand \U$22544 ( \22921 , \22914 , \22920 );
not \U$22545 ( \22922 , \22921 );
xor \U$22546 ( \22923 , \22907 , \22922 );
and \U$22547 ( \22924 , \6152 , \2322 );
not \U$22548 ( \22925 , \10807 );
and \U$22549 ( \22926 , RIae798e0_154, \2026 );
not \U$22550 ( \22927 , RIae798e0_154);
and \U$22551 ( \22928 , \22927 , \6359 );
nor \U$22552 ( \22929 , \22926 , \22928 );
nor \U$22553 ( \22930 , \22925 , \22929 );
nor \U$22554 ( \22931 , \22924 , \22930 );
and \U$22555 ( \22932 , \22923 , \22931 );
and \U$22556 ( \22933 , \22907 , \22922 );
or \U$22557 ( \22934 , \22932 , \22933 );
nor \U$22558 ( \22935 , \22894 , \22934 );
or \U$22559 ( \22936 , \22854 , \22935 );
nand \U$22560 ( \22937 , \22894 , \22934 );
nand \U$22561 ( \22938 , \22936 , \22937 );
xor \U$22562 ( \22939 , \6216 , \6265 );
xor \U$22563 ( \22940 , \22939 , \6306 );
xor \U$22564 ( \22941 , \22938 , \22940 );
xor \U$22565 ( \22942 , \6233 , \6263 );
xor \U$22566 ( \22943 , \22942 , \6249 );
not \U$22567 ( \22944 , \22943 );
not \U$22568 ( \22945 , \22944 );
nand \U$22569 ( \22946 , RIae7a2b8_175, RIae7a678_183);
and \U$22570 ( \22947 , \22946 , RIae79fe8_169);
not \U$22571 ( \22948 , \6246 );
not \U$22572 ( \22949 , \1320 );
not \U$22573 ( \22950 , \22949 );
and \U$22574 ( \22951 , \22948 , \22950 );
not \U$22575 ( \22952 , \10227 );
and \U$22576 ( \22953 , RIae78e90_132, \22952 );
not \U$22577 ( \22954 , RIae78e90_132);
and \U$22578 ( \22955 , \22954 , \4972 );
or \U$22579 ( \22956 , \22953 , \22955 );
and \U$22580 ( \22957 , \22956 , \5858 );
nor \U$22581 ( \22958 , \22951 , \22957 );
xor \U$22582 ( \22959 , \22947 , \22958 );
not \U$22583 ( \22960 , \797 );
not \U$22584 ( \22961 , \3208 );
and \U$22585 ( \22962 , \22961 , \3105 );
not \U$22586 ( \22963 , \22961 );
and \U$22587 ( \22964 , \22963 , RIae78f80_134);
nor \U$22588 ( \22965 , \22962 , \22964 );
not \U$22589 ( \22966 , \22965 );
or \U$22590 ( \22967 , \22960 , \22966 );
nand \U$22591 ( \22968 , \6066 , \839 );
nand \U$22592 ( \22969 , \22967 , \22968 );
not \U$22593 ( \22970 , \22969 );
and \U$22594 ( \22971 , \22959 , \22970 );
and \U$22595 ( \22972 , \22947 , \22958 );
nor \U$22596 ( \22973 , \22971 , \22972 );
not \U$22597 ( \22974 , \22973 );
xor \U$22598 ( \22975 , \6347 , RIae78b48_125);
not \U$22599 ( \22976 , \22975 );
nor \U$22600 ( \22977 , \22976 , \1959 );
xor \U$22601 ( \22978 , RIae78b48_125, \6232 );
not \U$22602 ( \22979 , \22978 );
nor \U$22603 ( \22980 , \22979 , \1128 );
nor \U$22604 ( \22981 , \22977 , \22980 );
not \U$22605 ( \22982 , \22981 );
nand \U$22606 ( \22983 , \15102 , RIae78b48_125);
not \U$22607 ( \22984 , \22983 );
nand \U$22608 ( \22985 , \6261 , \1027 );
not \U$22609 ( \22986 , \12838 );
not \U$22610 ( \22987 , \5722 );
or \U$22611 ( \22988 , \22986 , \22987 );
or \U$22612 ( \22989 , \21732 , \12843 );
nand \U$22613 ( \22990 , \22988 , \22989 );
nand \U$22614 ( \22991 , \22990 , \952 );
nand \U$22615 ( \22992 , \22985 , \22991 );
not \U$22616 ( \22993 , \22992 );
or \U$22617 ( \22994 , \22984 , \22993 );
or \U$22618 ( \22995 , \22992 , \22983 );
nand \U$22619 ( \22996 , \22994 , \22995 );
not \U$22620 ( \22997 , \22996 );
or \U$22621 ( \22998 , \22982 , \22997 );
nand \U$22622 ( \22999 , \22985 , \22991 , \22983 );
nand \U$22623 ( \23000 , \22998 , \22999 );
not \U$22624 ( \23001 , \23000 );
or \U$22625 ( \23002 , \22974 , \23001 );
or \U$22626 ( \23003 , \22973 , \23000 );
nand \U$22627 ( \23004 , \23002 , \23003 );
not \U$22628 ( \23005 , \23004 );
or \U$22629 ( \23006 , \22945 , \23005 );
not \U$22630 ( \23007 , \22973 );
nand \U$22631 ( \23008 , \23007 , \23000 );
nand \U$22632 ( \23009 , \23006 , \23008 );
xnor \U$22633 ( \23010 , \22941 , \23009 );
xor \U$22634 ( \23011 , \6373 , \6378 );
xor \U$22635 ( \23012 , \23011 , \6384 );
not \U$22636 ( \23013 , \6216 );
not \U$22637 ( \23014 , \1209 );
not \U$22638 ( \23015 , \6416 );
or \U$22639 ( \23016 , \23014 , \23015 );
nand \U$22640 ( \23017 , \22919 , \2157 );
nand \U$22641 ( \23018 , \23016 , \23017 );
not \U$22642 ( \23019 , \23018 );
not \U$22643 ( \23020 , \23019 );
or \U$22644 ( \23021 , \23013 , \23020 );
or \U$22645 ( \23022 , \6216 , \23019 );
not \U$22646 ( \23023 , \1501 );
not \U$22647 ( \23024 , \6402 );
or \U$22648 ( \23025 , \23023 , \23024 );
and \U$22649 ( \23026 , \10891 , RIae79250_140);
not \U$22650 ( \23027 , \10891 );
and \U$22651 ( \23028 , \23027 , \1503 );
nor \U$22652 ( \23029 , \23026 , \23028 );
nand \U$22653 ( \23030 , \23029 , \1499 );
nand \U$22654 ( \23031 , \23025 , \23030 );
not \U$22655 ( \23032 , \23031 );
nand \U$22656 ( \23033 , \23022 , \23032 );
nand \U$22657 ( \23034 , \23021 , \23033 );
xnor \U$22658 ( \23035 , \23012 , \23034 );
xor \U$22659 ( \23036 , \5927 , \5918 );
xnor \U$22660 ( \23037 , \23036 , \5935 );
xnor \U$22661 ( \23038 , \23035 , \23037 );
not \U$22662 ( \23039 , \1501 );
not \U$22663 ( \23040 , \23029 );
or \U$22664 ( \23041 , \23039 , \23040 );
and \U$22665 ( \23042 , RIae79250_140, \2676 );
not \U$22666 ( \23043 , RIae79250_140);
and \U$22667 ( \23044 , \23043 , \4837 );
or \U$22668 ( \23045 , \23042 , \23044 );
nand \U$22669 ( \23046 , \23045 , \2650 );
nand \U$22670 ( \23047 , \23041 , \23046 );
not \U$22671 ( \23048 , \11914 );
not \U$22672 ( \23049 , \11918 );
not \U$22673 ( \23050 , \992 );
or \U$22674 ( \23051 , \23049 , \23050 );
not \U$22675 ( \23052 , RIae79fe8_169);
or \U$22676 ( \23053 , \992 , \23052 );
nand \U$22677 ( \23054 , \23051 , \23053 );
not \U$22678 ( \23055 , \23054 );
or \U$22679 ( \23056 , \23048 , \23055 );
nand \U$22680 ( \23057 , \9518 , RIae79fe8_169);
nand \U$22681 ( \23058 , \23056 , \23057 );
and \U$22682 ( \23059 , \23047 , \23058 );
not \U$22683 ( \23060 , \868 );
not \U$22684 ( \23061 , \22978 );
or \U$22685 ( \23062 , \23060 , \23061 );
and \U$22686 ( \23063 , \860 , \14644 );
not \U$22687 ( \23064 , \860 );
and \U$22688 ( \23065 , \23064 , \9313 );
nor \U$22689 ( \23066 , \23063 , \23065 );
or \U$22690 ( \23067 , \23066 , \1976 );
nand \U$22691 ( \23068 , \23062 , \23067 );
not \U$22692 ( \23069 , \23068 );
not \U$22693 ( \23070 , \1320 );
not \U$22694 ( \23071 , \22956 );
or \U$22695 ( \23072 , \23070 , \23071 );
not \U$22696 ( \23073 , RIae78e90_132);
not \U$22697 ( \23074 , \13248 );
or \U$22698 ( \23075 , \23073 , \23074 );
or \U$22699 ( \23076 , \16310 , RIae78e90_132);
nand \U$22700 ( \23077 , \23075 , \23076 );
nand \U$22701 ( \23078 , \23077 , \1087 );
nand \U$22702 ( \23079 , \23072 , \23078 );
not \U$22703 ( \23080 , \23079 );
or \U$22704 ( \23081 , \23069 , \23080 );
or \U$22705 ( \23082 , \23079 , \23068 );
not \U$22706 ( \23083 , \5124 );
not \U$22707 ( \23084 , \22965 );
or \U$22708 ( \23085 , \23083 , \23084 );
and \U$22709 ( \23086 , RIae78f80_134, \6238 );
not \U$22710 ( \23087 , RIae78f80_134);
and \U$22711 ( \23088 , \23087 , \4169 );
or \U$22712 ( \23089 , \23086 , \23088 );
nand \U$22713 ( \23090 , \23089 , \797 );
nand \U$22714 ( \23091 , \23085 , \23090 );
nand \U$22715 ( \23092 , \23082 , \23091 );
nand \U$22716 ( \23093 , \23081 , \23092 );
or \U$22717 ( \23094 , \23059 , \23093 );
not \U$22718 ( \23095 , \23058 );
not \U$22719 ( \23096 , \23047 );
nand \U$22720 ( \23097 , \23095 , \23096 );
nand \U$22721 ( \23098 , \23094 , \23097 );
not \U$22722 ( \23099 , \23098 );
xor \U$22723 ( \23100 , \6068 , \6078 );
xor \U$22724 ( \23101 , \23100 , \6093 );
nand \U$22725 ( \23102 , \23099 , \23101 );
xor \U$22726 ( \23103 , \6167 , \6180 );
xor \U$22727 ( \23104 , \23103 , \6154 );
and \U$22728 ( \23105 , \23102 , \23104 );
nor \U$22729 ( \23106 , \23099 , \23101 );
nor \U$22730 ( \23107 , \23105 , \23106 );
xor \U$22731 ( \23108 , \6116 , \6127 );
xor \U$22732 ( \23109 , \23108 , \6109 );
xor \U$22733 ( \23110 , \6278 , \6287 );
xor \U$22734 ( \23111 , \23110 , \6303 );
nand \U$22735 ( \23112 , \23109 , \23111 );
not \U$22736 ( \23113 , \1049 );
not \U$22737 ( \23114 , \5914 );
or \U$22738 ( \23115 , \23113 , \23114 );
not \U$22739 ( \23116 , \22898 );
nand \U$22740 ( \23117 , \23116 , \1062 );
nand \U$22741 ( \23118 , \23115 , \23117 );
not \U$22742 ( \23119 , \1933 );
not \U$22743 ( \23120 , \22856 );
or \U$22744 ( \23121 , \23119 , \23120 );
nand \U$22745 ( \23122 , \6361 , \1919 );
nand \U$22746 ( \23123 , \23121 , \23122 );
not \U$22747 ( \23124 , \893 );
not \U$22748 ( \23125 , \22975 );
or \U$22749 ( \23126 , \23124 , \23125 );
nand \U$22750 ( \23127 , \6350 , \2096 );
nand \U$22751 ( \23128 , \23126 , \23127 );
and \U$22752 ( \23129 , \23123 , \23128 );
not \U$22753 ( \23130 , \23123 );
not \U$22754 ( \23131 , \23128 );
and \U$22755 ( \23132 , \23130 , \23131 );
nor \U$22756 ( \23133 , \23129 , \23132 );
xnor \U$22757 ( \23134 , \23118 , \23133 );
and \U$22758 ( \23135 , \23112 , \23134 );
nor \U$22759 ( \23136 , \23109 , \23111 );
nor \U$22760 ( \23137 , \23135 , \23136 );
not \U$22761 ( \23138 , \23137 );
and \U$22762 ( \23139 , \23107 , \23138 );
not \U$22763 ( \23140 , \23107 );
and \U$22764 ( \23141 , \23140 , \23137 );
nor \U$22765 ( \23142 , \23139 , \23141 );
xor \U$22766 ( \23143 , \23038 , \23142 );
xor \U$22767 ( \23144 , \23010 , \23143 );
xor \U$22768 ( \23145 , \6406 , \6418 );
xor \U$22769 ( \23146 , \23145 , \6424 );
xor \U$22770 ( \23147 , \5952 , \5964 );
xor \U$22771 ( \23148 , \23147 , \5976 );
xor \U$22772 ( \23149 , \23146 , \23148 );
not \U$22773 ( \23150 , \6001 );
nand \U$22774 ( \23151 , \23150 , \6011 );
xor \U$22775 ( \23152 , \23151 , \6009 );
xor \U$22776 ( \23153 , \23149 , \23152 );
not \U$22777 ( \23154 , \22969 );
buf \U$22778 ( \23155 , \22959 );
not \U$22779 ( \23156 , \23155 );
or \U$22780 ( \23157 , \23154 , \23156 );
or \U$22781 ( \23158 , \23155 , \22969 );
nand \U$22782 ( \23159 , \23157 , \23158 );
xnor \U$22783 ( \23160 , \22996 , \22981 );
not \U$22784 ( \23161 , \2341 );
not \U$22785 ( \23162 , RIae798e0_154);
not \U$22786 ( \23163 , \2593 );
or \U$22787 ( \23164 , \23162 , \23163 );
or \U$22788 ( \23165 , \3141 , RIae798e0_154);
nand \U$22789 ( \23166 , \23164 , \23165 );
not \U$22790 ( \23167 , \23166 );
or \U$22791 ( \23168 , \23161 , \23167 );
not \U$22792 ( \23169 , \22929 );
nand \U$22793 ( \23170 , \23169 , \2322 );
nand \U$22794 ( \23171 , \23168 , \23170 );
not \U$22795 ( \23172 , \23171 );
not \U$22796 ( \23173 , \952 );
not \U$22797 ( \23174 , \6346 );
xor \U$22798 ( \23175 , RIae78bc0_126, \23174 );
not \U$22799 ( \23176 , \23175 );
or \U$22800 ( \23177 , \23173 , \23176 );
nand \U$22801 ( \23178 , \22990 , \1027 );
nand \U$22802 ( \23179 , \23177 , \23178 );
not \U$22803 ( \23180 , \16977 );
nand \U$22804 ( \23181 , \23180 , RIae78b48_125);
and \U$22805 ( \23182 , \23179 , \23181 );
not \U$22806 ( \23183 , \23179 );
and \U$22807 ( \23184 , \15519 , RIae78b48_125);
and \U$22808 ( \23185 , \23183 , \23184 );
or \U$22809 ( \23186 , \23182 , \23185 );
not \U$22810 ( \23187 , \23186 );
or \U$22811 ( \23188 , \23172 , \23187 );
nand \U$22812 ( \23189 , \23179 , \23184 );
nand \U$22813 ( \23190 , \23188 , \23189 );
nand \U$22814 ( \23191 , \23160 , \23190 );
and \U$22815 ( \23192 , \23159 , \23191 );
nor \U$22816 ( \23193 , \23160 , \23190 );
nor \U$22817 ( \23194 , \23192 , \23193 );
not \U$22818 ( \23195 , \23194 );
not \U$22819 ( \23196 , \23004 );
not \U$22820 ( \23197 , \22943 );
and \U$22821 ( \23198 , \23196 , \23197 );
and \U$22822 ( \23199 , \23004 , \22943 );
nor \U$22823 ( \23200 , \23198 , \23199 );
not \U$22824 ( \23201 , \23200 );
or \U$22825 ( \23202 , \23195 , \23201 );
not \U$22826 ( \23203 , \14940 );
and \U$22827 ( \23204 , RIae79d90_164, \1141 );
not \U$22828 ( \23205 , RIae79d90_164);
and \U$22829 ( \23206 , \23205 , \1142 );
nor \U$22830 ( \23207 , \23204 , \23206 );
not \U$22831 ( \23208 , \23207 );
or \U$22832 ( \23209 , \23203 , \23208 );
not \U$22833 ( \23210 , RIae79d90_164);
not \U$22834 ( \23211 , \1158 );
or \U$22835 ( \23212 , \23210 , \23211 );
not \U$22836 ( \23213 , \3326 );
nand \U$22837 ( \23214 , \23213 , \4968 );
nand \U$22838 ( \23215 , \23212 , \23214 );
nand \U$22839 ( \23216 , \23215 , \5040 );
nand \U$22840 ( \23217 , \23209 , \23216 );
not \U$22841 ( \23218 , \3014 );
not \U$22842 ( \23219 , \22846 );
or \U$22843 ( \23220 , \23218 , \23219 );
not \U$22844 ( \23221 , \2268 );
not \U$22845 ( \23222 , \11071 );
or \U$22846 ( \23223 , \23221 , \23222 );
nand \U$22847 ( \23224 , \2153 , RIae79ac0_158);
nand \U$22848 ( \23225 , \23223 , \23224 );
nand \U$22849 ( \23226 , \23225 , \2272 );
nand \U$22850 ( \23227 , \23220 , \23226 );
or \U$22851 ( \23228 , \23217 , \23227 );
not \U$22852 ( \23229 , \11364 );
not \U$22853 ( \23230 , \22834 );
or \U$22854 ( \23231 , \23229 , \23230 );
not \U$22855 ( \23232 , \10688 );
not \U$22856 ( \23233 , RIae79c28_161);
and \U$22857 ( \23234 , \23232 , \23233 );
and \U$22858 ( \23235 , \3256 , RIae79c28_161);
nor \U$22859 ( \23236 , \23234 , \23235 );
nand \U$22860 ( \23237 , \23236 , \2767 );
nand \U$22861 ( \23238 , \23231 , \23237 );
nand \U$22862 ( \23239 , \23228 , \23238 );
buf \U$22863 ( \23240 , \23239 );
not \U$22864 ( \23241 , \1049 );
not \U$22865 ( \23242 , \22905 );
or \U$22866 ( \23243 , \23241 , \23242 );
and \U$22867 ( \23244 , RIae79070_136, \2402 );
not \U$22868 ( \23245 , RIae79070_136);
and \U$22869 ( \23246 , \23245 , \5673 );
or \U$22870 ( \23247 , \23244 , \23246 );
nand \U$22871 ( \23248 , \23247 , \1062 );
nand \U$22872 ( \23249 , \23243 , \23248 );
not \U$22873 ( \23250 , \1013 );
not \U$22874 ( \23251 , \22912 );
or \U$22875 ( \23252 , \23250 , \23251 );
and \U$22876 ( \23253 , RIae79160_138, \1973 );
not \U$22877 ( \23254 , RIae79160_138);
not \U$22878 ( \23255 , \14422 );
and \U$22879 ( \23256 , \23254 , \23255 );
nor \U$22880 ( \23257 , \23253 , \23256 );
nand \U$22881 ( \23258 , \23257 , \2157 );
nand \U$22882 ( \23259 , \23252 , \23258 );
xor \U$22883 ( \23260 , \23249 , \23259 );
not \U$22884 ( \23261 , \11409 );
not \U$22885 ( \23262 , \3283 );
not \U$22886 ( \23263 , RIae79ef8_167);
and \U$22887 ( \23264 , \23262 , \23263 );
and \U$22888 ( \23265 , \1994 , RIae79ef8_167);
nor \U$22889 ( \23266 , \23264 , \23265 );
not \U$22890 ( \23267 , \23266 );
or \U$22891 ( \23268 , \23261 , \23267 );
nand \U$22892 ( \23269 , \22873 , \6214 );
nand \U$22893 ( \23270 , \23268 , \23269 );
and \U$22894 ( \23271 , \23260 , \23270 );
and \U$22895 ( \23272 , \23249 , \23259 );
or \U$22896 ( \23273 , \23271 , \23272 );
not \U$22897 ( \23274 , \23273 );
nand \U$22898 ( \23275 , \23227 , \23217 );
buf \U$22899 ( \23276 , \23275 );
nand \U$22900 ( \23277 , \23240 , \23274 , \23276 );
and \U$22901 ( \23278 , \22824 , \2924 );
not \U$22902 ( \23279 , \2183 );
not \U$22903 ( \23280 , \2231 );
or \U$22904 ( \23281 , \23279 , \23280 );
nand \U$22905 ( \23282 , \3244 , RIae79520_146);
nand \U$22906 ( \23283 , \23281 , \23282 );
not \U$22907 ( \23284 , \23283 );
nor \U$22908 ( \23285 , \23284 , \6635 );
nor \U$22909 ( \23286 , \23278 , \23285 );
not \U$22910 ( \23287 , \23286 );
not \U$22911 ( \23288 , \4853 );
not \U$22912 ( \23289 , \22884 );
or \U$22913 ( \23290 , \23288 , \23289 );
and \U$22914 ( \23291 , RIae79ca0_162, \940 );
not \U$22915 ( \23292 , RIae79ca0_162);
and \U$22916 ( \23293 , \23292 , \3236 );
or \U$22917 ( \23294 , \23291 , \23293 );
nand \U$22918 ( \23295 , \23294 , \4842 );
nand \U$22919 ( \23296 , \23290 , \23295 );
not \U$22920 ( \23297 , \1919 );
not \U$22921 ( \23298 , \22862 );
or \U$22922 ( \23299 , \23297 , \23298 );
not \U$22923 ( \23300 , \3810 );
not \U$22924 ( \23301 , \3294 );
or \U$22925 ( \23302 , \23300 , \23301 );
or \U$22926 ( \23303 , \1899 , \3810 );
nand \U$22927 ( \23304 , \23302 , \23303 );
nand \U$22928 ( \23305 , \23304 , \1933 );
nand \U$22929 ( \23306 , \23299 , \23305 );
not \U$22930 ( \23307 , \23306 );
and \U$22931 ( \23308 , \23296 , \23307 );
not \U$22932 ( \23309 , \23296 );
and \U$22933 ( \23310 , \23309 , \23306 );
or \U$22934 ( \23311 , \23308 , \23310 );
not \U$22935 ( \23312 , \23311 );
or \U$22936 ( \23313 , \23287 , \23312 );
not \U$22937 ( \23314 , \23296 );
nand \U$22938 ( \23315 , \23314 , \23307 );
nand \U$22939 ( \23316 , \23313 , \23315 );
not \U$22940 ( \23317 , \23316 );
and \U$22941 ( \23318 , \23277 , \23317 );
and \U$22942 ( \23319 , \23240 , \23276 );
nor \U$22943 ( \23320 , \23319 , \23274 );
nor \U$22944 ( \23321 , \23318 , \23320 );
nand \U$22945 ( \23322 , \23202 , \23321 );
not \U$22946 ( \23323 , \23200 );
not \U$22947 ( \23324 , \23194 );
nand \U$22948 ( \23325 , \23323 , \23324 );
nand \U$22949 ( \23326 , \23322 , \23325 );
not \U$22950 ( \23327 , \23326 );
xor \U$22951 ( \23328 , \23153 , \23327 );
xor \U$22952 ( \23329 , \23144 , \23328 );
not \U$22953 ( \23330 , \23329 );
xor \U$22954 ( \23331 , \23324 , \23200 );
xor \U$22955 ( \23332 , \23331 , \23321 );
not \U$22956 ( \23333 , \23332 );
not \U$22957 ( \23334 , \23333 );
xor \U$22958 ( \23335 , \23134 , \23111 );
xnor \U$22959 ( \23336 , \23335 , \23109 );
not \U$22960 ( \23337 , \23336 );
not \U$22961 ( \23338 , \2450 );
and \U$22962 ( \23339 , RIae79778_151, \2917 );
not \U$22963 ( \23340 , RIae79778_151);
and \U$22964 ( \23341 , \23340 , \1119 );
nor \U$22965 ( \23342 , \23339 , \23341 );
not \U$22966 ( \23343 , \23342 );
or \U$22967 ( \23344 , \23338 , \23343 );
xor \U$22968 ( \23345 , RIae79778_151, \2262 );
nand \U$22969 ( \23346 , \23345 , \2433 );
nand \U$22970 ( \23347 , \23344 , \23346 );
not \U$22971 ( \23348 , \2011 );
and \U$22972 ( \23349 , RIae79610_148, \2857 );
not \U$22973 ( \23350 , RIae79610_148);
and \U$22974 ( \23351 , \23350 , \4023 );
or \U$22975 ( \23352 , \23349 , \23351 );
not \U$22976 ( \23353 , \23352 );
or \U$22977 ( \23354 , \23348 , \23353 );
not \U$22978 ( \23355 , \2056 );
not \U$22979 ( \23356 , \10908 );
or \U$22980 ( \23357 , \23355 , \23356 );
not \U$22981 ( \23358 , \10605 );
nand \U$22982 ( \23359 , \23358 , RIae79610_148);
nand \U$22983 ( \23360 , \23357 , \23359 );
nand \U$22984 ( \23361 , \23360 , \2063 );
nand \U$22985 ( \23362 , \23354 , \23361 );
not \U$22986 ( \23363 , \23362 );
not \U$22987 ( \23364 , \1844 );
and \U$22988 ( \23365 , RIae79688_149, \2287 );
not \U$22989 ( \23366 , RIae79688_149);
and \U$22990 ( \23367 , \23366 , \3748 );
or \U$22991 ( \23368 , \23365 , \23367 );
not \U$22992 ( \23369 , \23368 );
or \U$22993 ( \23370 , \23364 , \23369 );
not \U$22994 ( \23371 , \2970 );
not \U$22995 ( \23372 , \2310 );
or \U$22996 ( \23373 , \23371 , \23372 );
nand \U$22997 ( \23374 , \2305 , RIae79688_149);
nand \U$22998 ( \23375 , \23373 , \23374 );
nand \U$22999 ( \23376 , \23375 , \1821 );
nand \U$23000 ( \23377 , \23370 , \23376 );
and \U$23001 ( \23378 , \23363 , \23377 );
not \U$23002 ( \23379 , \23363 );
not \U$23003 ( \23380 , \23377 );
and \U$23004 ( \23381 , \23379 , \23380 );
or \U$23005 ( \23382 , \23378 , \23381 );
xnor \U$23006 ( \23383 , \23347 , \23382 );
xor \U$23007 ( \23384 , \23286 , \23311 );
xor \U$23008 ( \23385 , \23383 , \23384 );
not \U$23009 ( \23386 , \1049 );
not \U$23010 ( \23387 , RIae79070_136);
not \U$23011 ( \23388 , \10809 );
or \U$23012 ( \23389 , \23387 , \23388 );
not \U$23013 ( \23390 , \3207 );
not \U$23014 ( \23391 , \23390 );
nand \U$23015 ( \23392 , \23391 , \1039 );
nand \U$23016 ( \23393 , \23389 , \23392 );
not \U$23017 ( \23394 , \23393 );
or \U$23018 ( \23395 , \23386 , \23394 );
and \U$23019 ( \23396 , RIae79070_136, \6238 );
not \U$23020 ( \23397 , RIae79070_136);
and \U$23021 ( \23398 , \23397 , \4169 );
or \U$23022 ( \23399 , \23396 , \23398 );
nand \U$23023 ( \23400 , \23399 , \2276 );
nand \U$23024 ( \23401 , \23395 , \23400 );
not \U$23025 ( \23402 , \23401 );
not \U$23026 ( \23403 , \23402 );
not \U$23027 ( \23404 , \2063 );
and \U$23028 ( \23405 , RIae79610_148, \6398 );
not \U$23029 ( \23406 , RIae79610_148);
and \U$23030 ( \23407 , \23406 , \2697 );
nor \U$23031 ( \23408 , \23405 , \23407 );
not \U$23032 ( \23409 , \23408 );
or \U$23033 ( \23410 , \23404 , \23409 );
nand \U$23034 ( \23411 , \23360 , \2011 );
nand \U$23035 ( \23412 , \23410 , \23411 );
not \U$23036 ( \23413 , \23412 );
not \U$23037 ( \23414 , \23413 );
and \U$23038 ( \23415 , \23403 , \23414 );
and \U$23039 ( \23416 , \23412 , \23402 );
not \U$23040 ( \23417 , \23412 );
and \U$23041 ( \23418 , \23417 , \23401 );
nor \U$23042 ( \23419 , \23416 , \23418 );
not \U$23043 ( \23420 , \23419 );
not \U$23044 ( \23421 , \1910 );
not \U$23045 ( \23422 , \19456 );
and \U$23046 ( \23423 , RIae793b8_143, \23422 );
not \U$23047 ( \23424 , RIae793b8_143);
and \U$23048 ( \23425 , \23424 , \2564 );
nor \U$23049 ( \23426 , \23423 , \23425 );
not \U$23050 ( \23427 , \23426 );
or \U$23051 ( \23428 , \23421 , \23427 );
and \U$23052 ( \23429 , RIae793b8_143, \1789 );
not \U$23053 ( \23430 , RIae793b8_143);
and \U$23054 ( \23431 , \23430 , \13398 );
nor \U$23055 ( \23432 , \23429 , \23431 );
not \U$23056 ( \23433 , \23432 );
nand \U$23057 ( \23434 , \23433 , \1864 );
nand \U$23058 ( \23435 , \23428 , \23434 );
and \U$23059 ( \23436 , \23420 , \23435 );
nor \U$23060 ( \23437 , \23415 , \23436 );
and \U$23061 ( \23438 , \23385 , \23437 );
and \U$23062 ( \23439 , \23383 , \23384 );
or \U$23063 ( \23440 , \23438 , \23439 );
not \U$23064 ( \23441 , \23440 );
not \U$23065 ( \23442 , \23171 );
and \U$23066 ( \23443 , \23186 , \23442 );
not \U$23067 ( \23444 , \23186 );
and \U$23068 ( \23445 , \23444 , \23171 );
nor \U$23069 ( \23446 , \23443 , \23445 );
xor \U$23070 ( \23447 , \23091 , \23068 );
xnor \U$23071 ( \23448 , \23447 , \23079 );
xor \U$23072 ( \23449 , \23446 , \23448 );
and \U$23073 ( \23450 , RIae78b48_125, \14691 );
not \U$23074 ( \23451 , \2007 );
not \U$23075 ( \23452 , \2521 );
not \U$23076 ( \23453 , \1835 );
or \U$23077 ( \23454 , \23452 , \23453 );
nand \U$23078 ( \23455 , \1834 , RIae797f0_152);
nand \U$23079 ( \23456 , \23454 , \23455 );
not \U$23080 ( \23457 , \23456 );
or \U$23081 ( \23458 , \23451 , \23457 );
and \U$23082 ( \23459 , RIae797f0_152, \5134 );
not \U$23083 ( \23460 , RIae797f0_152);
and \U$23084 ( \23461 , \23460 , \14071 );
or \U$23085 ( \23462 , \23459 , \23461 );
nand \U$23086 ( \23463 , \23462 , \1989 );
nand \U$23087 ( \23464 , \23458 , \23463 );
xor \U$23088 ( \23465 , \23450 , \23464 );
not \U$23089 ( \23466 , \2650 );
and \U$23090 ( \23467 , RIae79250_140, \4113 );
not \U$23091 ( \23468 , RIae79250_140);
and \U$23092 ( \23469 , \23468 , \5115 );
or \U$23093 ( \23470 , \23467 , \23469 );
not \U$23094 ( \23471 , \23470 );
or \U$23095 ( \23472 , \23466 , \23471 );
and \U$23096 ( \23473 , RIae79250_140, \14439 );
not \U$23097 ( \23474 , RIae79250_140);
and \U$23098 ( \23475 , \23474 , \5891 );
or \U$23099 ( \23476 , \23473 , \23475 );
nand \U$23100 ( \23477 , \23476 , \1501 );
nand \U$23101 ( \23478 , \23472 , \23477 );
and \U$23102 ( \23479 , \23465 , \23478 );
and \U$23103 ( \23480 , \23450 , \23464 );
nor \U$23104 ( \23481 , \23479 , \23480 );
and \U$23105 ( \23482 , \23449 , \23481 );
and \U$23106 ( \23483 , \23446 , \23448 );
or \U$23107 ( \23484 , \23482 , \23483 );
not \U$23108 ( \23485 , \23484 );
not \U$23109 ( \23486 , \23485 );
not \U$23110 ( \23487 , \1209 );
not \U$23111 ( \23488 , \23257 );
or \U$23112 ( \23489 , \23487 , \23488 );
not \U$23113 ( \23490 , \997 );
not \U$23114 ( \23491 , \17596 );
or \U$23115 ( \23492 , \23490 , \23491 );
nand \U$23116 ( \23493 , \1860 , RIae79160_138);
nand \U$23117 ( \23494 , \23492 , \23493 );
nand \U$23118 ( \23495 , \23494 , \2157 );
nand \U$23119 ( \23496 , \23489 , \23495 );
not \U$23120 ( \23497 , \23496 );
not \U$23121 ( \23498 , \23497 );
not \U$23122 ( \23499 , \9518 );
not \U$23123 ( \23500 , \23054 );
or \U$23124 ( \23501 , \23499 , \23500 );
not \U$23125 ( \23502 , \834 );
and \U$23126 ( \23503 , RIae79fe8_169, \23502 );
not \U$23127 ( \23504 , RIae79fe8_169);
and \U$23128 ( \23505 , \23504 , \16395 );
nor \U$23129 ( \23506 , \23503 , \23505 );
nand \U$23130 ( \23507 , \23506 , \11914 );
nand \U$23131 ( \23508 , \23501 , \23507 );
not \U$23132 ( \23509 , \23508 );
not \U$23133 ( \23510 , \23509 );
or \U$23134 ( \23511 , \23498 , \23510 );
not \U$23135 ( \23512 , \23496 );
not \U$23136 ( \23513 , \23508 );
or \U$23137 ( \23514 , \23512 , \23513 );
and \U$23138 ( \23515 , \2322 , \23166 );
not \U$23139 ( \23516 , RIae798e0_154);
not \U$23140 ( \23517 , \1880 );
or \U$23141 ( \23518 , \23516 , \23517 );
or \U$23142 ( \23519 , \4458 , RIae798e0_154);
nand \U$23143 ( \23520 , \23518 , \23519 );
and \U$23144 ( \23521 , \23520 , \10807 );
nor \U$23145 ( \23522 , \23515 , \23521 );
nand \U$23146 ( \23523 , \23514 , \23522 );
nand \U$23147 ( \23524 , \23511 , \23523 );
not \U$23148 ( \23525 , \6091 );
and \U$23149 ( \23526 , \1439 , \13059 );
not \U$23150 ( \23527 , \1439 );
and \U$23151 ( \23528 , \23527 , RIae79d90_164);
nor \U$23152 ( \23529 , \23526 , \23528 );
not \U$23153 ( \23530 , \23529 );
or \U$23154 ( \23531 , \23525 , \23530 );
nand \U$23155 ( \23532 , \23215 , \6080 );
nand \U$23156 ( \23533 , \23531 , \23532 );
not \U$23157 ( \23534 , \4842 );
and \U$23158 ( \23535 , RIae79ca0_162, \854 );
not \U$23159 ( \23536 , RIae79ca0_162);
and \U$23160 ( \23537 , \23536 , \855 );
nor \U$23161 ( \23538 , \23535 , \23537 );
not \U$23162 ( \23539 , \23538 );
or \U$23163 ( \23540 , \23534 , \23539 );
nand \U$23164 ( \23541 , \23294 , \4853 );
nand \U$23165 ( \23542 , \23540 , \23541 );
xor \U$23166 ( \23543 , \23533 , \23542 );
not \U$23167 ( \23544 , \2458 );
not \U$23168 ( \23545 , RIae794a8_145);
not \U$23169 ( \23546 , \2212 );
or \U$23170 ( \23547 , \23545 , \23546 );
not \U$23171 ( \23548 , RIae794a8_145);
nand \U$23172 ( \23549 , \23548 , \4065 );
nand \U$23173 ( \23550 , \23547 , \23549 );
not \U$23174 ( \23551 , \23550 );
or \U$23175 ( \23552 , \23544 , \23551 );
nand \U$23176 ( \23553 , \23304 , \1919 );
nand \U$23177 ( \23554 , \23552 , \23553 );
and \U$23178 ( \23555 , \23543 , \23554 );
and \U$23179 ( \23556 , \23533 , \23542 );
nor \U$23180 ( \23557 , \23555 , \23556 );
xor \U$23181 ( \23558 , \23524 , \23557 );
not \U$23182 ( \23559 , \2767 );
xor \U$23183 ( \23560 , RIae79c28_161, \2917 );
not \U$23184 ( \23561 , \23560 );
or \U$23185 ( \23562 , \23559 , \23561 );
nand \U$23186 ( \23563 , \23236 , \5324 );
nand \U$23187 ( \23564 , \23562 , \23563 );
not \U$23188 ( \23565 , \23564 );
not \U$23189 ( \23566 , \23565 );
not \U$23190 ( \23567 , \6214 );
not \U$23191 ( \23568 , \23266 );
or \U$23192 ( \23569 , \23567 , \23568 );
and \U$23193 ( \23570 , \13733 , \1142 );
not \U$23194 ( \23571 , \13733 );
and \U$23195 ( \23572 , \23571 , \2640 );
nor \U$23196 ( \23573 , \23570 , \23572 );
nand \U$23197 ( \23574 , \23573 , \6201 );
nand \U$23198 ( \23575 , \23569 , \23574 );
not \U$23199 ( \23576 , \23575 );
not \U$23200 ( \23577 , RIae79520_146);
not \U$23201 ( \23578 , \2141 );
or \U$23202 ( \23579 , \23577 , \23578 );
or \U$23203 ( \23580 , \2137 , RIae79520_146);
nand \U$23204 ( \23581 , \23579 , \23580 );
nand \U$23205 ( \23582 , \23581 , \2189 );
nand \U$23206 ( \23583 , \23283 , \2610 );
nand \U$23207 ( \23584 , \23582 , \23583 );
not \U$23208 ( \23585 , \23584 );
not \U$23209 ( \23586 , \23585 );
or \U$23210 ( \23587 , \23576 , \23586 );
not \U$23211 ( \23588 , \23583 );
not \U$23212 ( \23589 , \23582 );
or \U$23213 ( \23590 , \23588 , \23589 );
not \U$23214 ( \23591 , \23575 );
nand \U$23215 ( \23592 , \23590 , \23591 );
nand \U$23216 ( \23593 , \23587 , \23592 );
not \U$23217 ( \23594 , \23593 );
or \U$23218 ( \23595 , \23566 , \23594 );
not \U$23219 ( \23596 , \23584 );
nand \U$23220 ( \23597 , \23596 , \23591 );
nand \U$23221 ( \23598 , \23595 , \23597 );
and \U$23222 ( \23599 , \23558 , \23598 );
and \U$23223 ( \23600 , \23524 , \23557 );
or \U$23224 ( \23601 , \23599 , \23600 );
not \U$23225 ( \23602 , \23601 );
or \U$23226 ( \23603 , \23486 , \23602 );
or \U$23227 ( \23604 , \23601 , \23485 );
nand \U$23228 ( \23605 , \23603 , \23604 );
not \U$23229 ( \23606 , \23605 );
or \U$23230 ( \23607 , \23441 , \23606 );
not \U$23231 ( \23608 , \23601 );
not \U$23232 ( \23609 , \23608 );
nand \U$23233 ( \23610 , \23609 , \23484 );
nand \U$23234 ( \23611 , \23607 , \23610 );
not \U$23235 ( \23612 , \23611 );
or \U$23236 ( \23613 , \23337 , \23612 );
or \U$23237 ( \23614 , \23336 , \23611 );
nand \U$23238 ( \23615 , \23613 , \23614 );
not \U$23239 ( \23616 , \23615 );
or \U$23240 ( \23617 , \23334 , \23616 );
not \U$23241 ( \23618 , \23336 );
nand \U$23242 ( \23619 , \23618 , \23611 );
nand \U$23243 ( \23620 , \23617 , \23619 );
not \U$23244 ( \23621 , \23620 );
or \U$23245 ( \23622 , \23330 , \23621 );
xor \U$23246 ( \23623 , \23328 , \23010 );
nand \U$23247 ( \23624 , \23623 , \23143 );
nand \U$23248 ( \23625 , \23622 , \23624 );
not \U$23249 ( \23626 , \23625 );
xor \U$23250 ( \23627 , \6437 , \6439 );
xor \U$23251 ( \23628 , \23627 , \6443 );
not \U$23252 ( \23629 , \23628 );
and \U$23253 ( \23630 , \6387 , \6367 );
not \U$23254 ( \23631 , \6387 );
and \U$23255 ( \23632 , \23631 , \6394 );
nor \U$23256 ( \23633 , \23630 , \23632 );
xor \U$23257 ( \23634 , \6391 , \23633 );
not \U$23258 ( \23635 , \23634 );
xor \U$23259 ( \23636 , \5939 , \5979 );
xor \U$23260 ( \23637 , \23636 , \6012 );
not \U$23261 ( \23638 , \23637 );
or \U$23262 ( \23639 , \23635 , \23638 );
or \U$23263 ( \23640 , \23637 , \23634 );
nand \U$23264 ( \23641 , \23639 , \23640 );
not \U$23265 ( \23642 , \23641 );
or \U$23266 ( \23643 , \23629 , \23642 );
or \U$23267 ( \23644 , \23641 , \23628 );
nand \U$23268 ( \23645 , \23643 , \23644 );
not \U$23269 ( \23646 , \23645 );
or \U$23270 ( \23647 , \23142 , \23038 );
not \U$23271 ( \23648 , \23138 );
buf \U$23272 ( \23649 , \23107 );
or \U$23273 ( \23650 , \23648 , \23649 );
nand \U$23274 ( \23651 , \23647 , \23650 );
xor \U$23275 ( \23652 , \6096 , \6183 );
buf \U$23276 ( \23653 , \6135 );
xnor \U$23277 ( \23654 , \23652 , \23653 );
not \U$23278 ( \23655 , \23654 );
not \U$23279 ( \23656 , \2063 );
not \U$23280 ( \23657 , \23352 );
or \U$23281 ( \23658 , \23656 , \23657 );
nand \U$23282 ( \23659 , \6159 , \2011 );
nand \U$23283 ( \23660 , \23658 , \23659 );
not \U$23284 ( \23661 , \1910 );
and \U$23285 ( \23662 , RIae793b8_143, \10883 );
not \U$23286 ( \23663 , RIae793b8_143);
and \U$23287 ( \23664 , \23663 , \3530 );
or \U$23288 ( \23665 , \23662 , \23664 );
not \U$23289 ( \23666 , \23665 );
or \U$23290 ( \23667 , \23661 , \23666 );
nand \U$23291 ( \23668 , \6178 , \1864 );
nand \U$23292 ( \23669 , \23667 , \23668 );
xor \U$23293 ( \23670 , \23660 , \23669 );
not \U$23294 ( \23671 , \2529 );
not \U$23295 ( \23672 , RIae797f0_152);
not \U$23296 ( \23673 , \1186 );
or \U$23297 ( \23674 , \23672 , \23673 );
or \U$23298 ( \23675 , \1186 , RIae797f0_152);
nand \U$23299 ( \23676 , \23674 , \23675 );
not \U$23300 ( \23677 , \23676 );
or \U$23301 ( \23678 , \23671 , \23677 );
nand \U$23302 ( \23679 , \6301 , \2007 );
nand \U$23303 ( \23680 , \23678 , \23679 );
and \U$23304 ( \23681 , \23670 , \23680 );
and \U$23305 ( \23682 , \23660 , \23669 );
or \U$23306 ( \23683 , \23681 , \23682 );
not \U$23307 ( \23684 , \23683 );
xor \U$23308 ( \23685 , \23018 , \23031 );
xnor \U$23309 ( \23686 , \23685 , \6216 );
not \U$23310 ( \23687 , \23686 );
or \U$23311 ( \23688 , \23684 , \23687 );
not \U$23312 ( \23689 , \1822 );
not \U$23313 ( \23690 , \6285 );
or \U$23314 ( \23691 , \23689 , \23690 );
nand \U$23315 ( \23692 , \23375 , \2966 );
nand \U$23316 ( \23693 , \23691 , \23692 );
not \U$23317 ( \23694 , \23693 );
and \U$23318 ( \23695 , \23342 , \2433 );
not \U$23319 ( \23696 , \2450 );
nor \U$23320 ( \23697 , \23696 , \6106 );
nor \U$23321 ( \23698 , \23695 , \23697 );
not \U$23322 ( \23699 , \5040 );
not \U$23323 ( \23700 , \23207 );
or \U$23324 ( \23701 , \23699 , \23700 );
nand \U$23325 ( \23702 , \6090 , \6080 );
nand \U$23326 ( \23703 , \23701 , \23702 );
xnor \U$23327 ( \23704 , \23698 , \23703 );
not \U$23328 ( \23705 , \23704 );
or \U$23329 ( \23706 , \23694 , \23705 );
and \U$23330 ( \23707 , \23342 , \2433 );
or \U$23331 ( \23708 , \23707 , \23697 );
nand \U$23332 ( \23709 , \23708 , \23703 );
nand \U$23333 ( \23710 , \23706 , \23709 );
not \U$23334 ( \23711 , \23710 );
nand \U$23335 ( \23712 , \23688 , \23711 );
not \U$23336 ( \23713 , \23683 );
not \U$23337 ( \23714 , \23686 );
nand \U$23338 ( \23715 , \23713 , \23714 );
nand \U$23339 ( \23716 , \23712 , \23715 );
not \U$23340 ( \23717 , \23123 );
not \U$23341 ( \23718 , \23118 );
or \U$23342 ( \23719 , \23717 , \23718 );
nand \U$23343 ( \23720 , \23719 , \23131 );
or \U$23344 ( \23721 , \23118 , \23123 );
nand \U$23345 ( \23722 , \23720 , \23721 );
xor \U$23346 ( \23723 , \6363 , \6353 );
xor \U$23347 ( \23724 , \23722 , \23723 );
xor \U$23348 ( \23725 , \5870 , \5880 );
xnor \U$23349 ( \23726 , \23725 , \5866 );
xnor \U$23350 ( \23727 , \23724 , \23726 );
xor \U$23351 ( \23728 , \23716 , \23727 );
not \U$23352 ( \23729 , \23728 );
or \U$23353 ( \23730 , \23655 , \23729 );
nand \U$23354 ( \23731 , \23727 , \23716 );
nand \U$23355 ( \23732 , \23730 , \23731 );
not \U$23356 ( \23733 , \23732 );
and \U$23357 ( \23734 , \23651 , \23733 );
not \U$23358 ( \23735 , \23651 );
and \U$23359 ( \23736 , \23735 , \23732 );
nor \U$23360 ( \23737 , \23734 , \23736 );
not \U$23361 ( \23738 , \23737 );
or \U$23362 ( \23739 , \23646 , \23738 );
or \U$23363 ( \23740 , \23645 , \23737 );
nand \U$23364 ( \23741 , \23739 , \23740 );
not \U$23365 ( \23742 , \23741 );
not \U$23366 ( \23743 , \22935 );
nand \U$23367 ( \23744 , \23743 , \22937 );
xor \U$23368 ( \23745 , \23744 , \22854 );
not \U$23369 ( \23746 , \23745 );
xor \U$23370 ( \23747 , \23660 , \23669 );
xor \U$23371 ( \23748 , \23747 , \23680 );
not \U$23372 ( \23749 , \23096 );
not \U$23373 ( \23750 , \23058 );
or \U$23374 ( \23751 , \23749 , \23750 );
not \U$23375 ( \23752 , \23095 );
or \U$23376 ( \23753 , \23752 , \23096 );
nand \U$23377 ( \23754 , \23751 , \23753 );
buf \U$23378 ( \23755 , \23093 );
xor \U$23379 ( \23756 , \23754 , \23755 );
xor \U$23380 ( \23757 , \23748 , \23756 );
not \U$23381 ( \23758 , \23066 );
not \U$23382 ( \23759 , \1959 );
and \U$23383 ( \23760 , \23758 , \23759 );
not \U$23384 ( \23761 , \860 );
not \U$23385 ( \23762 , \21743 );
or \U$23386 ( \23763 , \23761 , \23762 );
not \U$23387 ( \23764 , \23180 );
nand \U$23388 ( \23765 , \23764 , RIae78b48_125);
nand \U$23389 ( \23766 , \23763 , \23765 );
and \U$23390 ( \23767 , \23766 , \1129 );
nor \U$23391 ( \23768 , \23760 , \23767 );
not \U$23392 ( \23769 , \23768 );
not \U$23393 ( \23770 , \23769 );
not \U$23394 ( \23771 , \1074 );
not \U$23395 ( \23772 , \23077 );
or \U$23396 ( \23773 , \23771 , \23772 );
not \U$23397 ( \23774 , \1066 );
not \U$23398 ( \23775 , \9280 );
or \U$23399 ( \23776 , \23774 , \23775 );
nand \U$23400 ( \23777 , \10793 , RIae78e90_132);
nand \U$23401 ( \23778 , \23776 , \23777 );
nand \U$23402 ( \23779 , \23778 , \1087 );
nand \U$23403 ( \23780 , \23773 , \23779 );
and \U$23404 ( \23781 , \23175 , \1027 );
not \U$23405 ( \23782 , RIae78bc0_126);
not \U$23406 ( \23783 , \6231 );
or \U$23407 ( \23784 , \23782 , \23783 );
or \U$23408 ( \23785 , \22356 , RIae78bc0_126);
nand \U$23409 ( \23786 , \23784 , \23785 );
and \U$23410 ( \23787 , \23786 , \1036 );
nor \U$23411 ( \23788 , \23781 , \23787 );
and \U$23412 ( \23789 , \23780 , \23788 );
not \U$23413 ( \23790 , \23780 );
not \U$23414 ( \23791 , \23788 );
and \U$23415 ( \23792 , \23790 , \23791 );
or \U$23416 ( \23793 , \23789 , \23792 );
not \U$23417 ( \23794 , \23793 );
or \U$23418 ( \23795 , \23770 , \23794 );
nand \U$23419 ( \23796 , \23780 , \23791 );
nand \U$23420 ( \23797 , \23795 , \23796 );
not \U$23421 ( \23798 , \23797 );
not \U$23422 ( \23799 , \23752 );
not \U$23423 ( \23800 , \2276 );
not \U$23424 ( \23801 , \23393 );
or \U$23425 ( \23802 , \23800 , \23801 );
nand \U$23426 ( \23803 , \23247 , \1049 );
nand \U$23427 ( \23804 , \23802 , \23803 );
not \U$23428 ( \23805 , \23804 );
not \U$23429 ( \23806 , RIae7a240_174);
not \U$23430 ( \23807 , RIae7a1c8_173);
or \U$23431 ( \23808 , \23806 , \23807 );
nand \U$23432 ( \23809 , \23808 , RIae7a2b8_175);
not \U$23433 ( \23810 , \797 );
and \U$23434 ( \23811 , RIae78f80_134, \17010 );
not \U$23435 ( \23812 , RIae78f80_134);
and \U$23436 ( \23813 , \23812 , \10227 );
or \U$23437 ( \23814 , \23811 , \23813 );
not \U$23438 ( \23815 , \23814 );
or \U$23439 ( \23816 , \23810 , \23815 );
nand \U$23440 ( \23817 , \23089 , \839 );
nand \U$23441 ( \23818 , \23816 , \23817 );
and \U$23442 ( \23819 , \23809 , \23818 );
not \U$23443 ( \23820 , \23809 );
not \U$23444 ( \23821 , \23818 );
and \U$23445 ( \23822 , \23820 , \23821 );
nor \U$23446 ( \23823 , \23819 , \23822 );
not \U$23447 ( \23824 , \23823 );
or \U$23448 ( \23825 , \23805 , \23824 );
not \U$23449 ( \23826 , \23821 );
nand \U$23450 ( \23827 , \23826 , \23809 );
nand \U$23451 ( \23828 , \23825 , \23827 );
not \U$23452 ( \23829 , \23828 );
or \U$23453 ( \23830 , \23799 , \23829 );
or \U$23454 ( \23831 , \23828 , \23752 );
nand \U$23455 ( \23832 , \23830 , \23831 );
not \U$23456 ( \23833 , \23832 );
or \U$23457 ( \23834 , \23798 , \23833 );
nand \U$23458 ( \23835 , \23828 , \23095 );
nand \U$23459 ( \23836 , \23834 , \23835 );
and \U$23460 ( \23837 , \23757 , \23836 );
and \U$23461 ( \23838 , \23748 , \23756 );
or \U$23462 ( \23839 , \23837 , \23838 );
and \U$23463 ( \23840 , \23101 , \23098 );
not \U$23464 ( \23841 , \23101 );
and \U$23465 ( \23842 , \23841 , \23099 );
nor \U$23466 ( \23843 , \23840 , \23842 );
xor \U$23467 ( \23844 , \23843 , \23104 );
nand \U$23468 ( \23845 , \23839 , \23844 );
not \U$23469 ( \23846 , \23845 );
or \U$23470 ( \23847 , \23746 , \23846 );
or \U$23471 ( \23848 , \23839 , \23844 );
nand \U$23472 ( \23849 , \23847 , \23848 );
xor \U$23473 ( \23850 , \22864 , \22888 );
xnor \U$23474 ( \23851 , \23850 , \22892 );
xor \U$23475 ( \23852 , \23693 , \23704 );
xor \U$23476 ( \23853 , \23851 , \23852 );
not \U$23477 ( \23854 , \22839 );
nand \U$23478 ( \23855 , \23854 , \22853 );
not \U$23479 ( \23856 , \23855 );
xor \U$23480 ( \23857 , \22850 , \23856 );
and \U$23481 ( \23858 , \23853 , \23857 );
and \U$23482 ( \23859 , \23851 , \23852 );
or \U$23483 ( \23860 , \23858 , \23859 );
not \U$23484 ( \23861 , \23860 );
not \U$23485 ( \23862 , \23363 );
not \U$23486 ( \23863 , \23380 );
or \U$23487 ( \23864 , \23862 , \23863 );
nand \U$23488 ( \23865 , \23864 , \23347 );
nand \U$23489 ( \23866 , \23377 , \23362 );
and \U$23490 ( \23867 , \23865 , \23866 );
not \U$23491 ( \23868 , \1501 );
not \U$23492 ( \23869 , \23045 );
or \U$23493 ( \23870 , \23868 , \23869 );
nand \U$23494 ( \23871 , \23476 , \2650 );
nand \U$23495 ( \23872 , \23870 , \23871 );
not \U$23496 ( \23873 , \23872 );
not \U$23497 ( \23874 , \23432 );
not \U$23498 ( \23875 , \6846 );
and \U$23499 ( \23876 , \23874 , \23875 );
and \U$23500 ( \23877 , \23665 , \1864 );
nor \U$23501 ( \23878 , \23876 , \23877 );
not \U$23502 ( \23879 , \23878 );
not \U$23503 ( \23880 , \23879 );
or \U$23504 ( \23881 , \23873 , \23880 );
not \U$23505 ( \23882 , \2519 );
not \U$23506 ( \23883 , \23676 );
or \U$23507 ( \23884 , \23882 , \23883 );
nand \U$23508 ( \23885 , \23456 , \1989 );
nand \U$23509 ( \23886 , \23884 , \23885 );
not \U$23510 ( \23887 , \23872 );
nand \U$23511 ( \23888 , \23878 , \23887 );
nand \U$23512 ( \23889 , \23886 , \23888 );
nand \U$23513 ( \23890 , \23881 , \23889 );
not \U$23514 ( \23891 , \23890 );
xor \U$23515 ( \23892 , \23867 , \23891 );
xor \U$23516 ( \23893 , \22907 , \22922 );
xor \U$23517 ( \23894 , \23893 , \22931 );
and \U$23518 ( \23895 , \23892 , \23894 );
and \U$23519 ( \23896 , \23867 , \23891 );
or \U$23520 ( \23897 , \23895 , \23896 );
not \U$23521 ( \23898 , \23897 );
xor \U$23522 ( \23899 , \23683 , \23710 );
xnor \U$23523 ( \23900 , \23899 , \23714 );
nand \U$23524 ( \23901 , \23898 , \23900 );
nand \U$23525 ( \23902 , \23861 , \23901 );
not \U$23526 ( \23903 , \23900 );
nand \U$23527 ( \23904 , \23903 , \23897 );
nand \U$23528 ( \23905 , \23902 , \23904 );
not \U$23529 ( \23906 , \23654 );
not \U$23530 ( \23907 , \23728 );
not \U$23531 ( \23908 , \23907 );
or \U$23532 ( \23909 , \23906 , \23908 );
not \U$23533 ( \23910 , \23654 );
nand \U$23534 ( \23911 , \23910 , \23728 );
nand \U$23535 ( \23912 , \23909 , \23911 );
xor \U$23536 ( \23913 , \23905 , \23912 );
and \U$23537 ( \23914 , \23849 , \23913 );
and \U$23538 ( \23915 , \23912 , \23905 );
nor \U$23539 ( \23916 , \23914 , \23915 );
not \U$23540 ( \23917 , \23916 );
and \U$23541 ( \23918 , \23742 , \23917 );
and \U$23542 ( \23919 , \23916 , \23741 );
nor \U$23543 ( \23920 , \23918 , \23919 );
not \U$23544 ( \23921 , \23920 );
not \U$23545 ( \23922 , \23921 );
or \U$23546 ( \23923 , \23626 , \23922 );
not \U$23547 ( \23924 , \23916 );
nand \U$23548 ( \23925 , \23924 , \23741 );
nand \U$23549 ( \23926 , \23923 , \23925 );
not \U$23550 ( \23927 , \23926 );
not \U$23551 ( \23928 , \23927 );
not \U$23552 ( \23929 , \23009 );
nand \U$23553 ( \23930 , \23929 , \22940 );
not \U$23554 ( \23931 , \23930 );
not \U$23555 ( \23932 , \22938 );
or \U$23556 ( \23933 , \23931 , \23932 );
not \U$23557 ( \23934 , \22940 );
nand \U$23558 ( \23935 , \23934 , \23009 );
nand \U$23559 ( \23936 , \23933 , \23935 );
not \U$23560 ( \23937 , \23936 );
xor \U$23561 ( \23938 , \6427 , \6429 );
xor \U$23562 ( \23939 , \23938 , \6432 );
not \U$23563 ( \23940 , \23939 );
not \U$23564 ( \23941 , \6185 );
xnor \U$23565 ( \23942 , \5883 , \6060 );
not \U$23566 ( \23943 , \23942 );
not \U$23567 ( \23944 , \6309 );
or \U$23568 ( \23945 , \23943 , \23944 );
or \U$23569 ( \23946 , \6309 , \23942 );
nand \U$23570 ( \23947 , \23945 , \23946 );
not \U$23571 ( \23948 , \23947 );
or \U$23572 ( \23949 , \23941 , \23948 );
or \U$23573 ( \23950 , \23947 , \6185 );
nand \U$23574 ( \23951 , \23949 , \23950 );
not \U$23575 ( \23952 , \23951 );
or \U$23576 ( \23953 , \23940 , \23952 );
or \U$23577 ( \23954 , \23951 , \23939 );
nand \U$23578 ( \23955 , \23953 , \23954 );
not \U$23579 ( \23956 , \23955 );
or \U$23580 ( \23957 , \23937 , \23956 );
not \U$23581 ( \23958 , \23939 );
nand \U$23582 ( \23959 , \23958 , \23951 );
nand \U$23583 ( \23960 , \23957 , \23959 );
not \U$23584 ( \23961 , \23960 );
not \U$23585 ( \23962 , \6326 );
and \U$23586 ( \23963 , \6329 , \23962 );
not \U$23587 ( \23964 , \6329 );
and \U$23588 ( \23965 , \23964 , \6326 );
nor \U$23589 ( \23966 , \23963 , \23965 );
xor \U$23590 ( \23967 , \6322 , \23966 );
not \U$23591 ( \23968 , \23967 );
xor \U$23592 ( \23969 , \6056 , \6058 );
xor \U$23593 ( \23970 , \23969 , \6311 );
not \U$23594 ( \23971 , \23970 );
or \U$23595 ( \23972 , \23968 , \23971 );
or \U$23596 ( \23973 , \23970 , \23967 );
nand \U$23597 ( \23974 , \23972 , \23973 );
not \U$23598 ( \23975 , \23974 );
not \U$23599 ( \23976 , \23975 );
or \U$23600 ( \23977 , \23961 , \23976 );
not \U$23601 ( \23978 , \23960 );
nand \U$23602 ( \23979 , \23978 , \23974 );
nand \U$23603 ( \23980 , \23977 , \23979 );
xor \U$23604 ( \23981 , \23955 , \23936 );
not \U$23605 ( \23982 , \23981 );
not \U$23606 ( \23983 , \23010 );
not \U$23607 ( \23984 , \23328 );
or \U$23608 ( \23985 , \23983 , \23984 );
not \U$23609 ( \23986 , \23153 );
nand \U$23610 ( \23987 , \23986 , \23326 );
nand \U$23611 ( \23988 , \23985 , \23987 );
not \U$23612 ( \23989 , \23037 );
not \U$23613 ( \23990 , \23035 );
or \U$23614 ( \23991 , \23989 , \23990 );
not \U$23615 ( \23992 , \23012 );
nand \U$23616 ( \23993 , \23992 , \23034 );
nand \U$23617 ( \23994 , \23991 , \23993 );
not \U$23618 ( \23995 , \23994 );
xor \U$23619 ( \23996 , \23726 , \23722 );
not \U$23620 ( \23997 , \23723 );
and \U$23621 ( \23998 , \23996 , \23997 );
and \U$23622 ( \23999 , \23726 , \23722 );
or \U$23623 ( \24000 , \23998 , \23999 );
not \U$23624 ( \24001 , \24000 );
not \U$23625 ( \24002 , \24001 );
or \U$23626 ( \24003 , \23995 , \24002 );
or \U$23627 ( \24004 , \23994 , \24001 );
nand \U$23628 ( \24005 , \24003 , \24004 );
xor \U$23629 ( \24006 , \23146 , \23148 );
and \U$23630 ( \24007 , \24006 , \23152 );
and \U$23631 ( \24008 , \23146 , \23148 );
nor \U$23632 ( \24009 , \24007 , \24008 );
xor \U$23633 ( \24010 , \24005 , \24009 );
and \U$23634 ( \24011 , \23988 , \24010 );
not \U$23635 ( \24012 , \23988 );
not \U$23636 ( \24013 , \24010 );
and \U$23637 ( \24014 , \24012 , \24013 );
nor \U$23638 ( \24015 , \24011 , \24014 );
not \U$23639 ( \24016 , \24015 );
or \U$23640 ( \24017 , \23982 , \24016 );
buf \U$23641 ( \24018 , \23988 );
nand \U$23642 ( \24019 , \24018 , \24010 );
nand \U$23643 ( \24020 , \24017 , \24019 );
not \U$23644 ( \24021 , \24020 );
xor \U$23645 ( \24022 , \23980 , \24021 );
xor \U$23646 ( \24023 , \6396 , \6435 );
xor \U$23647 ( \24024 , \24023 , \6446 );
not \U$23648 ( \24025 , \24024 );
not \U$23649 ( \24026 , \24005 );
not \U$23650 ( \24027 , \24009 );
or \U$23651 ( \24028 , \24026 , \24027 );
nand \U$23652 ( \24029 , \23994 , \24000 );
nand \U$23653 ( \24030 , \24028 , \24029 );
not \U$23654 ( \24031 , \24030 );
or \U$23655 ( \24032 , \24025 , \24031 );
or \U$23656 ( \24033 , \24030 , \24024 );
nand \U$23657 ( \24034 , \24032 , \24033 );
not \U$23658 ( \24035 , \23628 );
not \U$23659 ( \24036 , \24035 );
not \U$23660 ( \24037 , \23641 );
or \U$23661 ( \24038 , \24036 , \24037 );
not \U$23662 ( \24039 , \23637 );
nand \U$23663 ( \24040 , \24039 , \23634 );
nand \U$23664 ( \24041 , \24038 , \24040 );
xnor \U$23665 ( \24042 , \24034 , \24041 );
not \U$23666 ( \24043 , \24042 );
not \U$23667 ( \24044 , \24043 );
not \U$23668 ( \24045 , \23737 );
not \U$23669 ( \24046 , \24045 );
not \U$23670 ( \24047 , \23645 );
or \U$23671 ( \24048 , \24046 , \24047 );
nand \U$23672 ( \24049 , \23732 , \23651 );
nand \U$23673 ( \24050 , \24048 , \24049 );
not \U$23674 ( \24051 , \24050 );
not \U$23675 ( \24052 , \24051 );
or \U$23676 ( \24053 , \24044 , \24052 );
nand \U$23677 ( \24054 , \24050 , \24042 );
nand \U$23678 ( \24055 , \24053 , \24054 );
xnor \U$23679 ( \24056 , \24022 , \24055 );
not \U$23680 ( \24057 , \24056 );
or \U$23681 ( \24058 , \23928 , \24057 );
or \U$23682 ( \24059 , \23927 , \24056 );
nand \U$23683 ( \24060 , \24058 , \24059 );
buf \U$23684 ( \24061 , \24060 );
xor \U$23685 ( \24062 , \23745 , \23844 );
xor \U$23686 ( \24063 , \24062 , \23839 );
not \U$23687 ( \24064 , \24063 );
xor \U$23688 ( \24065 , \23867 , \23891 );
xor \U$23689 ( \24066 , \24065 , \23894 );
not \U$23690 ( \24067 , \24066 );
nand \U$23691 ( \24068 , \23239 , \23275 );
and \U$23692 ( \24069 , \24068 , \23274 );
not \U$23693 ( \24070 , \24068 );
and \U$23694 ( \24071 , \24070 , \23273 );
nor \U$23695 ( \24072 , \24069 , \24071 );
xnor \U$23696 ( \24073 , \24072 , \23317 );
nand \U$23697 ( \24074 , \24067 , \24073 );
not \U$23698 ( \24075 , \24074 );
xor \U$23699 ( \24076 , \23249 , \23259 );
xor \U$23700 ( \24077 , \24076 , \23270 );
not \U$23701 ( \24078 , \24077 );
not \U$23702 ( \24079 , \2966 );
and \U$23703 ( \24080 , \1740 , RIae79688_149);
not \U$23704 ( \24081 , \1740 );
and \U$23705 ( \24082 , \24081 , \2970 );
nor \U$23706 ( \24083 , \24080 , \24082 );
not \U$23707 ( \24084 , \24083 );
or \U$23708 ( \24085 , \24079 , \24084 );
nand \U$23709 ( \24086 , \23368 , \3827 );
nand \U$23710 ( \24087 , \24085 , \24086 );
not \U$23711 ( \24088 , \2252 );
not \U$23712 ( \24089 , \23225 );
or \U$23713 ( \24090 , \24088 , \24089 );
and \U$23714 ( \24091 , \2309 , RIae79ac0_158);
not \U$23715 ( \24092 , \2309 );
and \U$23716 ( \24093 , \24092 , \2268 );
nor \U$23717 ( \24094 , \24091 , \24093 );
nand \U$23718 ( \24095 , \24094 , \2272 );
nand \U$23719 ( \24096 , \24090 , \24095 );
xor \U$23720 ( \24097 , \24087 , \24096 );
not \U$23721 ( \24098 , \2433 );
and \U$23722 ( \24099 , RIae79778_151, \3539 );
not \U$23723 ( \24100 , RIae79778_151);
and \U$23724 ( \24101 , \24100 , \10916 );
or \U$23725 ( \24102 , \24099 , \24101 );
not \U$23726 ( \24103 , \24102 );
or \U$23727 ( \24104 , \24098 , \24103 );
nand \U$23728 ( \24105 , \23345 , \2450 );
nand \U$23729 ( \24106 , \24104 , \24105 );
and \U$23730 ( \24107 , \24097 , \24106 );
and \U$23731 ( \24108 , \24087 , \24096 );
or \U$23732 ( \24109 , \24107 , \24108 );
not \U$23733 ( \24110 , \24109 );
not \U$23734 ( \24111 , \23238 );
xor \U$23735 ( \24112 , \23217 , \24111 );
xnor \U$23736 ( \24113 , \24112 , \23227 );
not \U$23737 ( \24114 , \24113 );
and \U$23738 ( \24115 , \24110 , \24114 );
not \U$23739 ( \24116 , \24110 );
and \U$23740 ( \24117 , \24116 , \24113 );
nor \U$23741 ( \24118 , \24115 , \24117 );
not \U$23742 ( \24119 , \24118 );
or \U$23743 ( \24120 , \24078 , \24119 );
nand \U$23744 ( \24121 , \24109 , \24113 );
nand \U$23745 ( \24122 , \24120 , \24121 );
not \U$23746 ( \24123 , \24122 );
not \U$23747 ( \24124 , \24123 );
or \U$23748 ( \24125 , \24075 , \24124 );
not \U$23749 ( \24126 , \24073 );
nand \U$23750 ( \24127 , \24126 , \24066 );
nand \U$23751 ( \24128 , \24125 , \24127 );
not \U$23752 ( \24129 , \24128 );
xor \U$23753 ( \24130 , \23897 , \23860 );
xnor \U$23754 ( \24131 , \24130 , \23900 );
not \U$23755 ( \24132 , \24131 );
or \U$23756 ( \24133 , \24129 , \24132 );
or \U$23757 ( \24134 , \24128 , \24131 );
nand \U$23758 ( \24135 , \24133 , \24134 );
not \U$23759 ( \24136 , \24135 );
or \U$23760 ( \24137 , \24064 , \24136 );
not \U$23761 ( \24138 , \24131 );
nand \U$23762 ( \24139 , \24138 , \24128 );
nand \U$23763 ( \24140 , \24137 , \24139 );
not \U$23764 ( \24141 , \24140 );
xnor \U$23765 ( \24142 , \23913 , \23849 );
not \U$23766 ( \24143 , \24142 );
or \U$23767 ( \24144 , \24141 , \24143 );
or \U$23768 ( \24145 , \24140 , \24142 );
nand \U$23769 ( \24146 , \24144 , \24145 );
not \U$23770 ( \24147 , \24146 );
xnor \U$23771 ( \24148 , \23329 , \23620 );
not \U$23772 ( \24149 , \24148 );
not \U$23773 ( \24150 , \24149 );
or \U$23774 ( \24151 , \24147 , \24150 );
not \U$23775 ( \24152 , \24142 );
nand \U$23776 ( \24153 , \24152 , \24140 );
nand \U$23777 ( \24154 , \24151 , \24153 );
not \U$23778 ( \24155 , \24154 );
xor \U$23779 ( \24156 , \24013 , \23981 );
xnor \U$23780 ( \24157 , \24156 , \24018 );
not \U$23781 ( \24158 , \24157 );
not \U$23782 ( \24159 , \24158 );
not \U$23783 ( \24160 , \23625 );
not \U$23784 ( \24161 , \24160 );
not \U$23785 ( \24162 , \23921 );
or \U$23786 ( \24163 , \24161 , \24162 );
nand \U$23787 ( \24164 , \23920 , \23625 );
nand \U$23788 ( \24165 , \24163 , \24164 );
not \U$23789 ( \24166 , \24165 );
or \U$23790 ( \24167 , \24159 , \24166 );
or \U$23791 ( \24168 , \24165 , \24158 );
nand \U$23792 ( \24169 , \24167 , \24168 );
not \U$23793 ( \24170 , \24169 );
or \U$23794 ( \24171 , \24155 , \24170 );
nand \U$23795 ( \24172 , \24165 , \24157 );
nand \U$23796 ( \24173 , \24171 , \24172 );
buf \U$23797 ( \24174 , \24173 );
nand \U$23798 ( \24175 , \24061 , \24174 );
nand \U$23799 ( \24176 , \24055 , \24021 );
not \U$23800 ( \24177 , \24176 );
not \U$23801 ( \24178 , \24055 );
nand \U$23802 ( \24179 , \24178 , \24020 );
not \U$23803 ( \24180 , \24179 );
or \U$23804 ( \24181 , \24177 , \24180 );
nand \U$23805 ( \24182 , \24181 , \23980 );
not \U$23806 ( \24183 , \24182 );
nand \U$23807 ( \24184 , \24056 , \23926 );
not \U$23808 ( \24185 , \24184 );
or \U$23809 ( \24186 , \24183 , \24185 );
not \U$23810 ( \24187 , \24020 );
not \U$23811 ( \24188 , \24055 );
or \U$23812 ( \24189 , \24187 , \24188 );
nand \U$23813 ( \24190 , \24050 , \24043 );
nand \U$23814 ( \24191 , \24189 , \24190 );
not \U$23815 ( \24192 , \24191 );
xor \U$23816 ( \24193 , \6055 , \6314 );
xor \U$23817 ( \24194 , \24193 , \6317 );
not \U$23818 ( \24195 , \23960 );
not \U$23819 ( \24196 , \23974 );
or \U$23820 ( \24197 , \24195 , \24196 );
not \U$23821 ( \24198 , \23970 );
nand \U$23822 ( \24199 , \24198 , \23967 );
nand \U$23823 ( \24200 , \24197 , \24199 );
not \U$23824 ( \24201 , \24200 );
xor \U$23825 ( \24202 , \24194 , \24201 );
not \U$23826 ( \24203 , \24041 );
not \U$23827 ( \24204 , \24034 );
or \U$23828 ( \24205 , \24203 , \24204 );
not \U$23829 ( \24206 , \24024 );
nand \U$23830 ( \24207 , \24206 , \24030 );
nand \U$23831 ( \24208 , \24205 , \24207 );
xor \U$23832 ( \24209 , \6332 , \6449 );
xor \U$23833 ( \24210 , \24209 , \6455 );
xnor \U$23834 ( \24211 , \24208 , \24210 );
xnor \U$23835 ( \24212 , \24202 , \24211 );
not \U$23836 ( \24213 , \24212 );
or \U$23837 ( \24214 , \24192 , \24213 );
or \U$23838 ( \24215 , \24191 , \24212 );
nand \U$23839 ( \24216 , \24214 , \24215 );
nand \U$23840 ( \24217 , \24186 , \24216 );
buf \U$23841 ( \24218 , \24217 );
xor \U$23842 ( \24219 , \6034 , \6025 );
xnor \U$23843 ( \24220 , \24219 , \5848 );
not \U$23844 ( \24221 , \6458 );
and \U$23845 ( \24222 , \6461 , \24221 );
not \U$23846 ( \24223 , \6461 );
and \U$23847 ( \24224 , \24223 , \6458 );
nor \U$23848 ( \24225 , \24222 , \24224 );
xor \U$23849 ( \24226 , \6320 , \24225 );
xor \U$23850 ( \24227 , \24220 , \24226 );
not \U$23851 ( \24228 , \24194 );
not \U$23852 ( \24229 , \24228 );
not \U$23853 ( \24230 , \24211 );
or \U$23854 ( \24231 , \24229 , \24230 );
not \U$23855 ( \24232 , \24210 );
nand \U$23856 ( \24233 , \24232 , \24208 );
nand \U$23857 ( \24234 , \24231 , \24233 );
xnor \U$23858 ( \24235 , \24227 , \24234 );
not \U$23859 ( \24236 , \24191 );
not \U$23860 ( \24237 , \24212 );
not \U$23861 ( \24238 , \24237 );
or \U$23862 ( \24239 , \24236 , \24238 );
and \U$23863 ( \24240 , \24211 , \24194 );
not \U$23864 ( \24241 , \24211 );
and \U$23865 ( \24242 , \24241 , \24228 );
or \U$23866 ( \24243 , \24240 , \24242 );
nand \U$23867 ( \24244 , \24243 , \24200 );
nand \U$23868 ( \24245 , \24239 , \24244 );
nand \U$23869 ( \24246 , \24235 , \24245 );
not \U$23870 ( \24247 , \24220 );
nand \U$23871 ( \24248 , \24247 , \24234 );
not \U$23872 ( \24249 , \24248 );
nand \U$23873 ( \24250 , \24234 , \24220 );
not \U$23874 ( \24251 , \24250 );
or \U$23875 ( \24252 , \24220 , \24234 );
not \U$23876 ( \24253 , \24252 );
or \U$23877 ( \24254 , \24251 , \24253 );
nand \U$23878 ( \24255 , \24254 , \24226 );
not \U$23879 ( \24256 , \24255 );
or \U$23880 ( \24257 , \24249 , \24256 );
xor \U$23881 ( \24258 , \6050 , \6464 );
xnor \U$23882 ( \24259 , \24258 , \6037 );
nand \U$23883 ( \24260 , \24257 , \24259 );
and \U$23884 ( \24261 , \24175 , \24218 , \24246 , \24260 );
xor \U$23885 ( \24262 , \22609 , \22776 );
and \U$23886 ( \24263 , \24262 , \22781 );
and \U$23887 ( \24264 , \22609 , \22776 );
or \U$23888 ( \24265 , \24263 , \24264 );
not \U$23889 ( \24266 , \22674 );
not \U$23890 ( \24267 , \24266 );
not \U$23891 ( \24268 , \22770 );
or \U$23892 ( \24269 , \24267 , \24268 );
nand \U$23893 ( \24270 , \24269 , \22775 );
or \U$23894 ( \24271 , \22770 , \24266 );
nand \U$23895 ( \24272 , \24270 , \24271 );
not \U$23896 ( \24273 , \22313 );
not \U$23897 ( \24274 , \22320 );
or \U$23898 ( \24275 , \24273 , \24274 );
or \U$23899 ( \24276 , \22313 , \22320 );
nand \U$23900 ( \24277 , \24276 , \22331 );
nand \U$23901 ( \24278 , \24275 , \24277 );
xor \U$23902 ( \24279 , \24272 , \24278 );
not \U$23903 ( \24280 , \1919 );
not \U$23904 ( \24281 , RIae794a8_145);
not \U$23905 ( \24282 , \2835 );
or \U$23906 ( \24283 , \24281 , \24282 );
or \U$23907 ( \24284 , \2835 , RIae794a8_145);
nand \U$23908 ( \24285 , \24283 , \24284 );
not \U$23909 ( \24286 , \24285 );
or \U$23910 ( \24287 , \24280 , \24286 );
nand \U$23911 ( \24288 , \22381 , \9828 );
nand \U$23912 ( \24289 , \24287 , \24288 );
not \U$23913 ( \24290 , \24289 );
not \U$23914 ( \24291 , \22676 );
and \U$23915 ( \24292 , \24290 , \24291 );
and \U$23916 ( \24293 , \24289 , \22676 );
nor \U$23917 ( \24294 , \24292 , \24293 );
and \U$23918 ( \24295 , \15989 , \22394 );
not \U$23919 ( \24296 , RIae79ef8_167);
not \U$23920 ( \24297 , \877 );
or \U$23921 ( \24298 , \24296 , \24297 );
or \U$23922 ( \24299 , \877 , RIae79ef8_167);
nand \U$23923 ( \24300 , \24298 , \24299 );
and \U$23924 ( \24301 , \24300 , \6214 );
nor \U$23925 ( \24302 , \24295 , \24301 );
xor \U$23926 ( \24303 , \24294 , \24302 );
not \U$23927 ( \24304 , \2776 );
not \U$23928 ( \24305 , RIae79c28_161);
not \U$23929 ( \24306 , \13033 );
or \U$23930 ( \24307 , \24305 , \24306 );
or \U$23931 ( \24308 , \2049 , RIae79c28_161);
nand \U$23932 ( \24309 , \24307 , \24308 );
not \U$23933 ( \24310 , \24309 );
or \U$23934 ( \24311 , \24304 , \24310 );
nand \U$23935 ( \24312 , \22740 , \2767 );
nand \U$23936 ( \24313 , \24311 , \24312 );
not \U$23937 ( \24314 , \9622 );
xor \U$23938 ( \24315 , RIae7a3a8_177, \991 );
not \U$23939 ( \24316 , \24315 );
or \U$23940 ( \24317 , \24314 , \24316 );
nand \U$23941 ( \24318 , \22750 , \11014 );
nand \U$23942 ( \24319 , \24317 , \24318 );
xor \U$23943 ( \24320 , \24313 , \24319 );
not \U$23944 ( \24321 , \2063 );
not \U$23945 ( \24322 , \22647 );
or \U$23946 ( \24323 , \24321 , \24322 );
and \U$23947 ( \24324 , RIae79610_148, \14422 );
not \U$23948 ( \24325 , RIae79610_148);
and \U$23949 ( \24326 , \24325 , \1970 );
nor \U$23950 ( \24327 , \24324 , \24326 );
nand \U$23951 ( \24328 , \24327 , \2011 );
nand \U$23952 ( \24329 , \24323 , \24328 );
xor \U$23953 ( \24330 , \24320 , \24329 );
xor \U$23954 ( \24331 , \24303 , \24330 );
not \U$23955 ( \24332 , \2322 );
and \U$23956 ( \24333 , RIae798e0_154, \2954 );
not \U$23957 ( \24334 , RIae798e0_154);
and \U$23958 ( \24335 , \24334 , \15033 );
or \U$23959 ( \24336 , \24333 , \24335 );
not \U$23960 ( \24337 , \24336 );
or \U$23961 ( \24338 , \24332 , \24337 );
nand \U$23962 ( \24339 , \22722 , \2340 );
nand \U$23963 ( \24340 , \24338 , \24339 );
not \U$23964 ( \24341 , \13121 );
not \U$23965 ( \24342 , \9532 );
not \U$23966 ( \24343 , RIae7a240_174);
and \U$23967 ( \24344 , \24342 , \24343 );
and \U$23968 ( \24345 , \781 , RIae7a240_174);
nor \U$23969 ( \24346 , \24344 , \24345 );
not \U$23970 ( \24347 , \24346 );
or \U$23971 ( \24348 , \24341 , \24347 );
nand \U$23972 ( \24349 , \22701 , \13720 );
nand \U$23973 ( \24350 , \24348 , \24349 );
xor \U$23974 ( \24351 , \24340 , \24350 );
not \U$23975 ( \24352 , \2519 );
not \U$23976 ( \24353 , \2521 );
not \U$23977 ( \24354 , \2230 );
not \U$23978 ( \24355 , \24354 );
or \U$23979 ( \24356 , \24353 , \24355 );
or \U$23980 ( \24357 , \2231 , \19713 );
nand \U$23981 ( \24358 , \24356 , \24357 );
not \U$23982 ( \24359 , \24358 );
or \U$23983 ( \24360 , \24352 , \24359 );
nand \U$23984 ( \24361 , \22711 , \1989 );
nand \U$23985 ( \24362 , \24360 , \24361 );
xor \U$23986 ( \24363 , \24351 , \24362 );
not \U$23987 ( \24364 , \24363 );
and \U$23988 ( \24365 , \24331 , \24364 );
not \U$23989 ( \24366 , \24331 );
and \U$23990 ( \24367 , \24366 , \24363 );
nor \U$23991 ( \24368 , \24365 , \24367 );
xor \U$23992 ( \24369 , \22632 , \22667 );
and \U$23993 ( \24370 , \24369 , \22673 );
and \U$23994 ( \24371 , \22632 , \22667 );
or \U$23995 ( \24372 , \24370 , \24371 );
not \U$23996 ( \24373 , \24372 );
and \U$23997 ( \24374 , RIae78b48_125, \9417 );
not \U$23998 ( \24375 , RIae78b48_125);
and \U$23999 ( \24376 , \24375 , \11198 );
nor \U$24000 ( \24377 , \24374 , \24376 );
not \U$24001 ( \24378 , \24377 );
not \U$24002 ( \24379 , \3267 );
and \U$24003 ( \24380 , \24378 , \24379 );
and \U$24004 ( \24381 , \22568 , \1129 );
nor \U$24005 ( \24382 , \24380 , \24381 );
not \U$24006 ( \24383 , \4853 );
not \U$24007 ( \24384 , RIae79ca0_162);
not \U$24008 ( \24385 , \2847 );
or \U$24009 ( \24386 , \24384 , \24385 );
or \U$24010 ( \24387 , \1833 , RIae79ca0_162);
nand \U$24011 ( \24388 , \24386 , \24387 );
not \U$24012 ( \24389 , \24388 );
or \U$24013 ( \24390 , \24383 , \24389 );
nand \U$24014 ( \24391 , \22659 , \11762 );
nand \U$24015 ( \24392 , \24390 , \24391 );
not \U$24016 ( \24393 , \24392 );
xor \U$24017 ( \24394 , \24382 , \24393 );
not \U$24018 ( \24395 , \1843 );
not \U$24019 ( \24396 , \22638 );
or \U$24020 ( \24397 , \24395 , \24396 );
not \U$24021 ( \24398 , RIae79688_149);
not \U$24022 ( \24399 , \13008 );
or \U$24023 ( \24400 , \24398 , \24399 );
nand \U$24024 ( \24401 , \14907 , \13986 );
nand \U$24025 ( \24402 , \24400 , \24401 );
nand \U$24026 ( \24403 , \1821 , \24402 );
nand \U$24027 ( \24404 , \24397 , \24403 );
not \U$24028 ( \24405 , \24404 );
xnor \U$24029 ( \24406 , \24394 , \24405 );
not \U$24030 ( \24407 , \9792 );
not \U$24031 ( \24408 , \22759 );
or \U$24032 ( \24409 , \24407 , \24408 );
not \U$24033 ( \24410 , RIae7a2b8_175);
not \U$24034 ( \24411 , \11441 );
or \U$24035 ( \24412 , \24410 , \24411 );
or \U$24036 ( \24413 , \1288 , RIae7a2b8_175);
nand \U$24037 ( \24414 , \24412 , \24413 );
nand \U$24038 ( \24415 , \24414 , \9814 );
nand \U$24039 ( \24416 , \24409 , \24415 );
not \U$24040 ( \24417 , \11914 );
not \U$24041 ( \24418 , \22678 );
or \U$24042 ( \24419 , \24417 , \24418 );
and \U$24043 ( \24420 , RIae79fe8_169, \9770 );
not \U$24044 ( \24421 , RIae79fe8_169);
and \U$24045 ( \24422 , \24421 , \18413 );
nor \U$24046 ( \24423 , \24420 , \24422 );
nand \U$24047 ( \24424 , \24423 , \9518 );
nand \U$24048 ( \24425 , \24419 , \24424 );
xor \U$24049 ( \24426 , \24416 , \24425 );
not \U$24050 ( \24427 , \2545 );
not \U$24051 ( \24428 , \22688 );
or \U$24052 ( \24429 , \24427 , \24428 );
not \U$24053 ( \24430 , \2447 );
not \U$24054 ( \24431 , \3294 );
or \U$24055 ( \24432 , \24430 , \24431 );
or \U$24056 ( \24433 , \13087 , \2504 );
nand \U$24057 ( \24434 , \24432 , \24433 );
nand \U$24058 ( \24435 , \24434 , \2450 );
nand \U$24059 ( \24436 , \24429 , \24435 );
xor \U$24060 ( \24437 , \24426 , \24436 );
xor \U$24061 ( \24438 , \24406 , \24437 );
buf \U$24062 ( \24439 , \24438 );
not \U$24063 ( \24440 , \2189 );
not \U$24064 ( \24441 , \22621 );
or \U$24065 ( \24442 , \24440 , \24441 );
and \U$24066 ( \24443 , RIae79520_146, \1760 );
not \U$24067 ( \24444 , RIae79520_146);
not \U$24068 ( \24445 , \4583 );
and \U$24069 ( \24446 , \24444 , \24445 );
or \U$24070 ( \24447 , \24443 , \24446 );
nand \U$24071 ( \24448 , \24447 , \3440 );
nand \U$24072 ( \24449 , \24442 , \24448 );
not \U$24073 ( \24450 , \2272 );
not \U$24074 ( \24451 , \22611 );
or \U$24075 ( \24452 , \24450 , \24451 );
not \U$24076 ( \24453 , RIae79ac0_158);
not \U$24077 ( \24454 , \1789 );
or \U$24078 ( \24455 , \24453 , \24454 );
nand \U$24079 ( \24456 , \13398 , \2268 );
nand \U$24080 ( \24457 , \24455 , \24456 );
nand \U$24081 ( \24458 , \24457 , \2252 );
nand \U$24082 ( \24459 , \24452 , \24458 );
xor \U$24083 ( \24460 , \24449 , \24459 );
not \U$24084 ( \24461 , \5040 );
not \U$24085 ( \24462 , \22408 );
or \U$24086 ( \24463 , \24461 , \24462 );
not \U$24087 ( \24464 , RIae79d90_164);
not \U$24088 ( \24465 , \975 );
or \U$24089 ( \24466 , \24464 , \24465 );
or \U$24090 ( \24467 , \16510 , RIae79d90_164);
nand \U$24091 ( \24468 , \24466 , \24467 );
nand \U$24092 ( \24469 , \24468 , \14940 );
nand \U$24093 ( \24470 , \24463 , \24469 );
xor \U$24094 ( \24471 , \24460 , \24470 );
buf \U$24095 ( \24472 , \24471 );
not \U$24096 ( \24473 , \24472 );
and \U$24097 ( \24474 , \24439 , \24473 );
not \U$24098 ( \24475 , \24439 );
and \U$24099 ( \24476 , \24475 , \24472 );
nor \U$24100 ( \24477 , \24474 , \24476 );
not \U$24101 ( \24478 , \24477 );
or \U$24102 ( \24479 , \24373 , \24478 );
or \U$24103 ( \24480 , \24372 , \24477 );
nand \U$24104 ( \24481 , \24479 , \24480 );
xnor \U$24105 ( \24482 , \24368 , \24481 );
buf \U$24106 ( \24483 , \24482 );
xor \U$24107 ( \24484 , \24279 , \24483 );
xor \U$24108 ( \24485 , \24265 , \24484 );
not \U$24109 ( \24486 , \22582 );
not \U$24110 ( \24487 , \22442 );
nand \U$24111 ( \24488 , \24487 , \22487 );
not \U$24112 ( \24489 , \24488 );
or \U$24113 ( \24490 , \24486 , \24489 );
not \U$24114 ( \24491 , \22487 );
nand \U$24115 ( \24492 , \24491 , \22442 );
nand \U$24116 ( \24493 , \24490 , \24492 );
not \U$24117 ( \24494 , \24493 );
not \U$24118 ( \24495 , \22460 );
not \U$24119 ( \24496 , \22486 );
or \U$24120 ( \24497 , \24495 , \24496 );
or \U$24121 ( \24498 , \22486 , \22460 );
nand \U$24122 ( \24499 , \24498 , \22449 );
nand \U$24123 ( \24500 , \24497 , \24499 );
not \U$24124 ( \24501 , \22492 );
not \U$24125 ( \24502 , \24501 );
not \U$24126 ( \24503 , \22518 );
or \U$24127 ( \24504 , \24502 , \24503 );
nand \U$24128 ( \24505 , \24504 , \22581 );
not \U$24129 ( \24506 , \24501 );
nand \U$24130 ( \24507 , \24506 , \22519 );
nand \U$24131 ( \24508 , \24505 , \24507 );
xor \U$24132 ( \24509 , \24500 , \24508 );
xor \U$24133 ( \24510 , \22350 , \22362 );
and \U$24134 ( \24511 , \24510 , \22372 );
and \U$24135 ( \24512 , \22350 , \22362 );
or \U$24136 ( \24513 , \24511 , \24512 );
not \U$24137 ( \24514 , \1910 );
not \U$24138 ( \24515 , \22550 );
or \U$24139 ( \24516 , \24514 , \24515 );
not \U$24140 ( \24517 , RIae793b8_143);
not \U$24141 ( \24518 , \2402 );
or \U$24142 ( \24519 , \24517 , \24518 );
or \U$24143 ( \24520 , \3270 , RIae793b8_143);
nand \U$24144 ( \24521 , \24519 , \24520 );
nand \U$24145 ( \24522 , \24521 , \1863 );
nand \U$24146 ( \24523 , \24516 , \24522 );
not \U$24147 ( \24524 , \24523 );
nand \U$24148 ( \24525 , \15504 , RIae78b48_125);
and \U$24149 ( \24526 , RIae7a498_179, RIae7a588_181);
nor \U$24150 ( \24527 , \24526 , \10633 );
or \U$24151 ( \24528 , \24525 , \24527 );
nand \U$24152 ( \24529 , \24525 , \24527 );
nand \U$24153 ( \24530 , \24528 , \24529 );
not \U$24154 ( \24531 , \24530 );
and \U$24155 ( \24532 , \24524 , \24531 );
and \U$24156 ( \24533 , \24523 , \24530 );
nor \U$24157 ( \24534 , \24532 , \24533 );
not \U$24158 ( \24535 , \24534 );
and \U$24159 ( \24536 , \24513 , \24535 );
not \U$24160 ( \24537 , \24513 );
and \U$24161 ( \24538 , \24537 , \24534 );
nor \U$24162 ( \24539 , \24536 , \24538 );
not \U$24163 ( \24540 , \22552 );
not \U$24164 ( \24541 , \22532 );
not \U$24165 ( \24542 , \22542 );
or \U$24166 ( \24543 , \24541 , \24542 );
or \U$24167 ( \24544 , \22542 , \22532 );
nand \U$24168 ( \24545 , \24543 , \24544 );
not \U$24169 ( \24546 , \24545 );
or \U$24170 ( \24547 , \24540 , \24546 );
not \U$24171 ( \24548 , \22532 );
nand \U$24172 ( \24549 , \24548 , \22542 );
nand \U$24173 ( \24550 , \24547 , \24549 );
and \U$24174 ( \24551 , \24539 , \24550 );
not \U$24175 ( \24552 , \24539 );
not \U$24176 ( \24553 , \24550 );
and \U$24177 ( \24554 , \24552 , \24553 );
nor \U$24178 ( \24555 , \24551 , \24554 );
not \U$24179 ( \24556 , \22513 );
not \U$24180 ( \24557 , \22508 );
or \U$24181 ( \24558 , \24556 , \24557 );
not \U$24182 ( \24559 , \22503 );
not \U$24183 ( \24560 , \22499 );
or \U$24184 ( \24561 , \24559 , \24560 );
nand \U$24185 ( \24562 , \24561 , \22497 );
nand \U$24186 ( \24563 , \24558 , \24562 );
xor \U$24187 ( \24564 , \24555 , \24563 );
xor \U$24188 ( \24565 , \22524 , \22553 );
and \U$24189 ( \24566 , \24565 , \22580 );
and \U$24190 ( \24567 , \22524 , \22553 );
or \U$24191 ( \24568 , \24566 , \24567 );
xnor \U$24192 ( \24569 , \24564 , \24568 );
xnor \U$24193 ( \24570 , \24509 , \24569 );
nand \U$24194 ( \24571 , \24494 , \24570 );
not \U$24195 ( \24572 , \24570 );
nand \U$24196 ( \24573 , \24572 , \24493 );
nand \U$24197 ( \24574 , \24571 , \24573 );
not \U$24198 ( \24575 , \22415 );
not \U$24199 ( \24576 , \22437 );
or \U$24200 ( \24577 , \24575 , \24576 );
not \U$24201 ( \24578 , \22423 );
nand \U$24202 ( \24579 , \24578 , \22436 );
nand \U$24203 ( \24580 , \24577 , \24579 );
xor \U$24204 ( \24581 , \22468 , \22472 );
and \U$24205 ( \24582 , \24581 , \22485 );
and \U$24206 ( \24583 , \22468 , \22472 );
or \U$24207 ( \24584 , \24582 , \24583 );
not \U$24208 ( \24585 , \22615 );
not \U$24209 ( \24586 , \22631 );
or \U$24210 ( \24587 , \24585 , \24586 );
not \U$24211 ( \24588 , \22622 );
not \U$24212 ( \24589 , \22616 );
or \U$24213 ( \24590 , \24588 , \24589 );
nand \U$24214 ( \24591 , \24590 , \22630 );
nand \U$24215 ( \24592 , \24587 , \24591 );
not \U$24216 ( \24593 , \22642 );
not \U$24217 ( \24594 , \22666 );
or \U$24218 ( \24595 , \24593 , \24594 );
nand \U$24219 ( \24596 , \22661 , \22651 );
nand \U$24220 ( \24597 , \24595 , \24596 );
xor \U$24221 ( \24598 , \24592 , \24597 );
not \U$24222 ( \24599 , \22412 );
not \U$24223 ( \24600 , \22402 );
or \U$24224 ( \24601 , \24599 , \24600 );
nand \U$24225 ( \24602 , \22398 , \22385 );
nand \U$24226 ( \24603 , \24601 , \24602 );
buf \U$24227 ( \24604 , \24603 );
xor \U$24228 ( \24605 , \24598 , \24604 );
xor \U$24229 ( \24606 , \24584 , \24605 );
not \U$24230 ( \24607 , \5858 );
not \U$24231 ( \24608 , \22346 );
or \U$24232 ( \24609 , \24607 , \24608 );
and \U$24233 ( \24610 , RIae78e90_132, \13287 );
not \U$24234 ( \24611 , RIae78e90_132);
and \U$24235 ( \24612 , \24611 , \14691 );
or \U$24236 ( \24613 , \24610 , \24612 );
nand \U$24237 ( \24614 , \24613 , \1072 );
nand \U$24238 ( \24615 , \24609 , \24614 );
not \U$24239 ( \24616 , \951 );
not \U$24240 ( \24617 , \22562 );
or \U$24241 ( \24618 , \24616 , \24617 );
and \U$24242 ( \24619 , RIae78bc0_126, \13301 );
not \U$24243 ( \24620 , RIae78bc0_126);
and \U$24244 ( \24621 , \24620 , \16786 );
or \U$24245 ( \24622 , \24619 , \24621 );
nand \U$24246 ( \24623 , \24622 , \927 );
nand \U$24247 ( \24624 , \24618 , \24623 );
xor \U$24248 ( \24625 , \24615 , \24624 );
not \U$24249 ( \24626 , \796 );
not \U$24250 ( \24627 , \22368 );
or \U$24251 ( \24628 , \24626 , \24627 );
and \U$24252 ( \24629 , RIae78f80_134, \9313 );
not \U$24253 ( \24630 , RIae78f80_134);
and \U$24254 ( \24631 , \24630 , \14644 );
or \U$24255 ( \24632 , \24629 , \24631 );
nand \U$24256 ( \24633 , \24632 , \5124 );
nand \U$24257 ( \24634 , \24628 , \24633 );
xor \U$24258 ( \24635 , \24625 , \24634 );
not \U$24259 ( \24636 , \22566 );
and \U$24260 ( \24637 , \22579 , \22572 );
not \U$24261 ( \24638 , \22579 );
and \U$24262 ( \24639 , \24638 , \22573 );
nor \U$24263 ( \24640 , \24637 , \24639 );
not \U$24264 ( \24641 , \24640 );
or \U$24265 ( \24642 , \24636 , \24641 );
nand \U$24266 ( \24643 , \22579 , \22572 );
nand \U$24267 ( \24644 , \24642 , \24643 );
and \U$24268 ( \24645 , \24635 , \24644 );
not \U$24269 ( \24646 , \24635 );
not \U$24270 ( \24647 , \24644 );
and \U$24271 ( \24648 , \24646 , \24647 );
nor \U$24272 ( \24649 , \24645 , \24648 );
not \U$24273 ( \24650 , \22729 );
not \U$24274 ( \24651 , \22705 );
or \U$24275 ( \24652 , \24650 , \24651 );
nand \U$24276 ( \24653 , \22715 , \22724 );
nand \U$24277 ( \24654 , \24652 , \24653 );
and \U$24278 ( \24655 , \24649 , \24654 );
not \U$24279 ( \24656 , \24649 );
not \U$24280 ( \24657 , \24654 );
and \U$24281 ( \24658 , \24656 , \24657 );
nor \U$24282 ( \24659 , \24655 , \24658 );
xor \U$24283 ( \24660 , \24606 , \24659 );
xor \U$24284 ( \24661 , \24580 , \24660 );
xor \U$24285 ( \24662 , \22340 , \22373 );
and \U$24286 ( \24663 , \24662 , \22413 );
and \U$24287 ( \24664 , \22340 , \22373 );
or \U$24288 ( \24665 , \24663 , \24664 );
not \U$24289 ( \24666 , \1062 );
not \U$24290 ( \24667 , \22358 );
or \U$24291 ( \24668 , \24666 , \24667 );
not \U$24292 ( \24669 , RIae79070_136);
not \U$24293 ( \24670 , \15117 );
or \U$24294 ( \24671 , \24669 , \24670 );
not \U$24295 ( \24672 , \9291 );
nand \U$24296 ( \24673 , \24672 , \1039 );
nand \U$24297 ( \24674 , \24671 , \24673 );
nand \U$24298 ( \24675 , \24674 , \1049 );
nand \U$24299 ( \24676 , \24668 , \24675 );
not \U$24300 ( \24677 , \1013 );
not \U$24301 ( \24678 , \997 );
not \U$24302 ( \24679 , \6257 );
not \U$24303 ( \24680 , \24679 );
or \U$24304 ( \24681 , \24678 , \24680 );
nand \U$24305 ( \24682 , \16310 , RIae79160_138);
nand \U$24306 ( \24683 , \24681 , \24682 );
not \U$24307 ( \24684 , \24683 );
or \U$24308 ( \24685 , \24677 , \24684 );
nand \U$24309 ( \24686 , \22529 , \2157 );
nand \U$24310 ( \24687 , \24685 , \24686 );
xor \U$24311 ( \24688 , \24676 , \24687 );
not \U$24312 ( \24689 , \1501 );
not \U$24313 ( \24690 , RIae79250_140);
not \U$24314 ( \24691 , \6238 );
or \U$24315 ( \24692 , \24690 , \24691 );
or \U$24316 ( \24693 , \6244 , RIae79250_140);
nand \U$24317 ( \24694 , \24692 , \24693 );
not \U$24318 ( \24695 , \24694 );
or \U$24319 ( \24696 , \24689 , \24695 );
nand \U$24320 ( \24697 , \22538 , \2650 );
nand \U$24321 ( \24698 , \24696 , \24697 );
xor \U$24322 ( \24699 , \24688 , \24698 );
xor \U$24323 ( \24700 , \22744 , \22754 );
and \U$24324 ( \24701 , \24700 , \22764 );
and \U$24325 ( \24702 , \22744 , \22754 );
or \U$24326 ( \24703 , \24701 , \24702 );
xor \U$24327 ( \24704 , \24699 , \24703 );
xor \U$24328 ( \24705 , \22682 , \22676 );
and \U$24329 ( \24706 , \24705 , \22692 );
and \U$24330 ( \24707 , \22682 , \22676 );
or \U$24331 ( \24708 , \24706 , \24707 );
xor \U$24332 ( \24709 , \24704 , \24708 );
xor \U$24333 ( \24710 , \24665 , \24709 );
not \U$24334 ( \24711 , \22765 );
not \U$24335 ( \24712 , \22735 );
or \U$24336 ( \24713 , \24711 , \24712 );
nand \U$24337 ( \24714 , \22730 , \22694 );
nand \U$24338 ( \24715 , \24713 , \24714 );
not \U$24339 ( \24716 , \24715 );
xor \U$24340 ( \24717 , \24710 , \24716 );
xnor \U$24341 ( \24718 , \24661 , \24717 );
and \U$24342 ( \24719 , \24574 , \24718 );
not \U$24343 ( \24720 , \24574 );
not \U$24344 ( \24721 , \24718 );
and \U$24345 ( \24722 , \24720 , \24721 );
nor \U$24346 ( \24723 , \24719 , \24722 );
and \U$24347 ( \24724 , \24485 , \24723 );
and \U$24348 ( \24725 , \24265 , \24484 );
or \U$24349 ( \24726 , \24724 , \24725 );
not \U$24350 ( \24727 , \24726 );
not \U$24351 ( \24728 , \24727 );
not \U$24352 ( \24729 , \24654 );
not \U$24353 ( \24730 , \24649 );
or \U$24354 ( \24731 , \24729 , \24730 );
nand \U$24355 ( \24732 , \24644 , \24635 );
nand \U$24356 ( \24733 , \24731 , \24732 );
not \U$24357 ( \24734 , \24529 );
not \U$24358 ( \24735 , \24523 );
or \U$24359 ( \24736 , \24734 , \24735 );
nand \U$24360 ( \24737 , \24736 , \24528 );
not \U$24361 ( \24738 , \24737 );
not \U$24362 ( \24739 , \1501 );
and \U$24363 ( \24740 , RIae79250_140, \22961 );
not \U$24364 ( \24741 , RIae79250_140);
not \U$24365 ( \24742 , \13999 );
and \U$24366 ( \24743 , \24741 , \24742 );
or \U$24367 ( \24744 , \24740 , \24743 );
not \U$24368 ( \24745 , \24744 );
or \U$24369 ( \24746 , \24739 , \24745 );
nand \U$24370 ( \24747 , \24694 , \2650 );
nand \U$24371 ( \24748 , \24746 , \24747 );
not \U$24372 ( \24749 , \24748 );
or \U$24373 ( \24750 , \24738 , \24749 );
or \U$24374 ( \24751 , \24737 , \24748 );
nand \U$24375 ( \24752 , \24750 , \24751 );
not \U$24376 ( \24753 , \24752 );
xor \U$24377 ( \24754 , \24676 , \24687 );
and \U$24378 ( \24755 , \24754 , \24698 );
and \U$24379 ( \24756 , \24676 , \24687 );
or \U$24380 ( \24757 , \24755 , \24756 );
not \U$24381 ( \24758 , \24757 );
not \U$24382 ( \24759 , \24758 );
and \U$24383 ( \24760 , \24753 , \24759 );
and \U$24384 ( \24761 , \24752 , \24758 );
nor \U$24385 ( \24762 , \24760 , \24761 );
not \U$24386 ( \24763 , \24550 );
not \U$24387 ( \24764 , \24539 );
or \U$24388 ( \24765 , \24763 , \24764 );
nand \U$24389 ( \24766 , \24513 , \24535 );
nand \U$24390 ( \24767 , \24765 , \24766 );
xnor \U$24391 ( \24768 , \24762 , \24767 );
xnor \U$24392 ( \24769 , \24733 , \24768 );
not \U$24393 ( \24770 , \24555 );
not \U$24394 ( \24771 , \24563 );
or \U$24395 ( \24772 , \24770 , \24771 );
or \U$24396 ( \24773 , \24563 , \24555 );
nand \U$24397 ( \24774 , \24773 , \24568 );
nand \U$24398 ( \24775 , \24772 , \24774 );
xor \U$24399 ( \24776 , \24769 , \24775 );
xor \U$24400 ( \24777 , \24584 , \24605 );
and \U$24401 ( \24778 , \24777 , \24659 );
and \U$24402 ( \24779 , \24584 , \24605 );
or \U$24403 ( \24780 , \24778 , \24779 );
xnor \U$24404 ( \24781 , \24776 , \24780 );
not \U$24405 ( \24782 , \24781 );
not \U$24406 ( \24783 , \24368 );
not \U$24407 ( \24784 , \24783 );
not \U$24408 ( \24785 , \24481 );
or \U$24409 ( \24786 , \24784 , \24785 );
not \U$24410 ( \24787 , \24477 );
nand \U$24411 ( \24788 , \24787 , \24372 );
nand \U$24412 ( \24789 , \24786 , \24788 );
not \U$24413 ( \24790 , \24789 );
not \U$24414 ( \24791 , \24665 );
not \U$24415 ( \24792 , \24791 );
not \U$24416 ( \24793 , \24716 );
or \U$24417 ( \24794 , \24792 , \24793 );
nand \U$24418 ( \24795 , \24794 , \24709 );
nand \U$24419 ( \24796 , \24715 , \24665 );
nand \U$24420 ( \24797 , \24795 , \24796 );
not \U$24421 ( \24798 , \24797 );
not \U$24422 ( \24799 , \24382 );
xor \U$24423 ( \24800 , \24799 , \24392 );
not \U$24424 ( \24801 , \24405 );
and \U$24425 ( \24802 , \24800 , \24801 );
and \U$24426 ( \24803 , \24799 , \24392 );
nor \U$24427 ( \24804 , \24802 , \24803 );
not \U$24428 ( \24805 , \927 );
and \U$24429 ( \24806 , \14110 , RIae78bc0_126);
not \U$24430 ( \24807 , \14110 );
and \U$24431 ( \24808 , \24807 , \1286 );
nor \U$24432 ( \24809 , \24806 , \24808 );
not \U$24433 ( \24810 , \24809 );
or \U$24434 ( \24811 , \24805 , \24810 );
nand \U$24435 ( \24812 , \24622 , \951 );
nand \U$24436 ( \24813 , \24811 , \24812 );
not \U$24437 ( \24814 , \1320 );
not \U$24438 ( \24815 , \9347 );
not \U$24439 ( \24816 , \24815 );
and \U$24440 ( \24817 , RIae78e90_132, \24816 );
not \U$24441 ( \24818 , RIae78e90_132);
and \U$24442 ( \24819 , \24818 , \21747 );
or \U$24443 ( \24820 , \24817 , \24819 );
not \U$24444 ( \24821 , \24820 );
or \U$24445 ( \24822 , \24814 , \24821 );
nand \U$24446 ( \24823 , \24613 , \5858 );
nand \U$24447 ( \24824 , \24822 , \24823 );
xor \U$24448 ( \24825 , \24813 , \24824 );
not \U$24449 ( \24826 , \12515 );
not \U$24450 ( \24827 , \24315 );
or \U$24451 ( \24828 , \24826 , \24827 );
nand \U$24452 ( \24829 , \9622 , RIae7a3a8_177);
nand \U$24453 ( \24830 , \24828 , \24829 );
xnor \U$24454 ( \24831 , \24825 , \24830 );
not \U$24455 ( \24832 , \24831 );
xor \U$24456 ( \24833 , \24804 , \24832 );
xor \U$24457 ( \24834 , \24449 , \24459 );
and \U$24458 ( \24835 , \24834 , \24470 );
and \U$24459 ( \24836 , \24449 , \24459 );
or \U$24460 ( \24837 , \24835 , \24836 );
not \U$24461 ( \24838 , \24837 );
xnor \U$24462 ( \24839 , \24833 , \24838 );
not \U$24463 ( \24840 , \24839 );
not \U$24464 ( \24841 , \24597 );
not \U$24465 ( \24842 , \24603 );
not \U$24466 ( \24843 , \24592 );
not \U$24467 ( \24844 , \24843 );
or \U$24468 ( \24845 , \24842 , \24844 );
or \U$24469 ( \24846 , \24603 , \24843 );
nand \U$24470 ( \24847 , \24845 , \24846 );
not \U$24471 ( \24848 , \24847 );
or \U$24472 ( \24849 , \24841 , \24848 );
not \U$24473 ( \24850 , \24843 );
nand \U$24474 ( \24851 , \24850 , \24604 );
nand \U$24475 ( \24852 , \24849 , \24851 );
not \U$24476 ( \24853 , \24852 );
and \U$24477 ( \24854 , \24438 , \24471 );
and \U$24478 ( \24855 , \24406 , \24437 );
nor \U$24479 ( \24856 , \24854 , \24855 );
not \U$24480 ( \24857 , \24856 );
or \U$24481 ( \24858 , \24853 , \24857 );
not \U$24482 ( \24859 , \24855 );
not \U$24483 ( \24860 , \24859 );
not \U$24484 ( \24861 , \24854 );
not \U$24485 ( \24862 , \24861 );
or \U$24486 ( \24863 , \24860 , \24862 );
not \U$24487 ( \24864 , \24852 );
nand \U$24488 ( \24865 , \24863 , \24864 );
nand \U$24489 ( \24866 , \24858 , \24865 );
not \U$24490 ( \24867 , \24866 );
or \U$24491 ( \24868 , \24840 , \24867 );
or \U$24492 ( \24869 , \24839 , \24866 );
nand \U$24493 ( \24870 , \24868 , \24869 );
not \U$24494 ( \24871 , \24870 );
not \U$24495 ( \24872 , \24871 );
or \U$24496 ( \24873 , \24798 , \24872 );
not \U$24497 ( \24874 , \24797 );
nand \U$24498 ( \24875 , \24874 , \24870 );
nand \U$24499 ( \24876 , \24873 , \24875 );
not \U$24500 ( \24877 , \24876 );
or \U$24501 ( \24878 , \24790 , \24877 );
or \U$24502 ( \24879 , \24876 , \24789 );
nand \U$24503 ( \24880 , \24878 , \24879 );
not \U$24504 ( \24881 , \24880 );
or \U$24505 ( \24882 , \24782 , \24881 );
or \U$24506 ( \24883 , \24781 , \24880 );
nand \U$24507 ( \24884 , \24882 , \24883 );
not \U$24508 ( \24885 , \24717 );
xnor \U$24509 ( \24886 , \24580 , \24660 );
not \U$24510 ( \24887 , \24886 );
or \U$24511 ( \24888 , \24885 , \24887 );
not \U$24512 ( \24889 , \24660 );
nand \U$24513 ( \24890 , \24889 , \24580 );
nand \U$24514 ( \24891 , \24888 , \24890 );
xor \U$24515 ( \24892 , \24884 , \24891 );
not \U$24516 ( \24893 , \24892 );
not \U$24517 ( \24894 , \24718 );
not \U$24518 ( \24895 , \24571 );
or \U$24519 ( \24896 , \24894 , \24895 );
nand \U$24520 ( \24897 , \24896 , \24573 );
not \U$24521 ( \24898 , \24897 );
not \U$24522 ( \24899 , \24898 );
or \U$24523 ( \24900 , \24294 , \24302 );
not \U$24524 ( \24901 , \24289 );
or \U$24525 ( \24902 , \24901 , \22676 );
nand \U$24526 ( \24903 , \24900 , \24902 );
not \U$24527 ( \24904 , \24903 );
xor \U$24528 ( \24905 , \24615 , \24634 );
and \U$24529 ( \24906 , \24905 , \24624 );
and \U$24530 ( \24907 , \24615 , \24634 );
nor \U$24531 ( \24908 , \24906 , \24907 );
not \U$24532 ( \24909 , \24908 );
or \U$24533 ( \24910 , \24904 , \24909 );
or \U$24534 ( \24911 , \24908 , \24903 );
nand \U$24535 ( \24912 , \24910 , \24911 );
not \U$24536 ( \24913 , \24912 );
not \U$24537 ( \24914 , \24436 );
not \U$24538 ( \24915 , \11914 );
not \U$24539 ( \24916 , \22678 );
or \U$24540 ( \24917 , \24915 , \24916 );
nand \U$24541 ( \24918 , \24917 , \24424 );
and \U$24542 ( \24919 , \24918 , \24416 );
not \U$24543 ( \24920 , \24918 );
not \U$24544 ( \24921 , \24416 );
and \U$24545 ( \24922 , \24920 , \24921 );
nor \U$24546 ( \24923 , \24919 , \24922 );
not \U$24547 ( \24924 , \24923 );
or \U$24548 ( \24925 , \24914 , \24924 );
nand \U$24549 ( \24926 , \24918 , \24416 );
nand \U$24550 ( \24927 , \24925 , \24926 );
not \U$24551 ( \24928 , \24927 );
not \U$24552 ( \24929 , \24928 );
and \U$24553 ( \24930 , \24913 , \24929 );
and \U$24554 ( \24931 , \24912 , \24928 );
nor \U$24555 ( \24932 , \24930 , \24931 );
xor \U$24556 ( \24933 , \24699 , \24703 );
and \U$24557 ( \24934 , \24933 , \24708 );
and \U$24558 ( \24935 , \24699 , \24703 );
or \U$24559 ( \24936 , \24934 , \24935 );
not \U$24560 ( \24937 , \24936 );
xor \U$24561 ( \24938 , \24932 , \24937 );
and \U$24562 ( \24939 , \24331 , \24363 );
and \U$24563 ( \24940 , \24303 , \24330 );
nor \U$24564 ( \24941 , \24939 , \24940 );
xor \U$24565 ( \24942 , \24938 , \24941 );
xor \U$24566 ( \24943 , \24340 , \24350 );
and \U$24567 ( \24944 , \24943 , \24362 );
and \U$24568 ( \24945 , \24340 , \24350 );
or \U$24569 ( \24946 , \24944 , \24945 );
and \U$24570 ( \24947 , RIae78b48_125, \9607 );
not \U$24571 ( \24948 , \2096 );
and \U$24572 ( \24949 , \22560 , \860 );
not \U$24573 ( \24950 , \22560 );
and \U$24574 ( \24951 , \24950 , RIae78b48_125);
nor \U$24575 ( \24952 , \24949 , \24951 );
not \U$24576 ( \24953 , \24952 );
or \U$24577 ( \24954 , \24948 , \24953 );
not \U$24578 ( \24955 , \24377 );
nand \U$24579 ( \24956 , \24955 , \893 );
nand \U$24580 ( \24957 , \24954 , \24956 );
xor \U$24581 ( \24958 , \24947 , \24957 );
not \U$24582 ( \24959 , \2776 );
not \U$24583 ( \24960 , RIae79c28_161);
not \U$24584 ( \24961 , \2026 );
or \U$24585 ( \24962 , \24960 , \24961 );
or \U$24586 ( \24963 , \16086 , RIae79c28_161);
nand \U$24587 ( \24964 , \24962 , \24963 );
not \U$24588 ( \24965 , \24964 );
or \U$24589 ( \24966 , \24959 , \24965 );
nand \U$24590 ( \24967 , \24309 , \2767 );
nand \U$24591 ( \24968 , \24966 , \24967 );
xor \U$24592 ( \24969 , \24958 , \24968 );
not \U$24593 ( \24970 , \24969 );
not \U$24594 ( \24971 , \5124 );
not \U$24595 ( \24972 , RIae78f80_134);
not \U$24596 ( \24973 , \14120 );
or \U$24597 ( \24974 , \24972 , \24973 );
nand \U$24598 ( \24975 , \6230 , \3105 );
nand \U$24599 ( \24976 , \24974 , \24975 );
not \U$24600 ( \24977 , \24976 );
or \U$24601 ( \24978 , \24971 , \24977 );
nand \U$24602 ( \24979 , \24632 , \796 );
nand \U$24603 ( \24980 , \24978 , \24979 );
not \U$24604 ( \24981 , \1062 );
not \U$24605 ( \24982 , \24674 );
or \U$24606 ( \24983 , \24981 , \24982 );
and \U$24607 ( \24984 , RIae79070_136, \13976 );
not \U$24608 ( \24985 , RIae79070_136);
and \U$24609 ( \24986 , \24985 , \5722 );
or \U$24610 ( \24987 , \24984 , \24986 );
nand \U$24611 ( \24988 , \24987 , \1049 );
nand \U$24612 ( \24989 , \24983 , \24988 );
xor \U$24613 ( \24990 , \24980 , \24989 );
xnor \U$24614 ( \24991 , RIae79160_138, \10226 );
not \U$24615 ( \24992 , \24991 );
not \U$24616 ( \24993 , \1013 );
or \U$24617 ( \24994 , \24992 , \24993 );
nand \U$24618 ( \24995 , \24683 , \2157 );
nand \U$24619 ( \24996 , \24994 , \24995 );
xor \U$24620 ( \24997 , \24990 , \24996 );
not \U$24621 ( \24998 , \24997 );
or \U$24622 ( \24999 , \24970 , \24998 );
or \U$24623 ( \25000 , \24997 , \24969 );
nand \U$24624 ( \25001 , \24999 , \25000 );
xor \U$24625 ( \25002 , \24946 , \25001 );
and \U$24626 ( \25003 , RIae79ef8_167, \9760 );
not \U$24627 ( \25004 , RIae79ef8_167);
and \U$24628 ( \25005 , \25004 , \854 );
or \U$24629 ( \25006 , \25003 , \25005 );
not \U$24630 ( \25007 , \25006 );
not \U$24631 ( \25008 , \10573 );
or \U$24632 ( \25009 , \25007 , \25008 );
nand \U$24633 ( \25010 , \24300 , \14768 );
nand \U$24634 ( \25011 , \25009 , \25010 );
not \U$24635 ( \25012 , \9814 );
not \U$24636 ( \25013 , \11054 );
not \U$24637 ( \25014 , \10551 );
or \U$24638 ( \25015 , \25013 , \25014 );
or \U$24639 ( \25016 , \10551 , \9804 );
nand \U$24640 ( \25017 , \25015 , \25016 );
not \U$24641 ( \25018 , \25017 );
or \U$24642 ( \25019 , \25012 , \25018 );
nand \U$24643 ( \25020 , \24414 , \9792 );
nand \U$24644 ( \25021 , \25019 , \25020 );
xor \U$24645 ( \25022 , \25011 , \25021 );
not \U$24646 ( \25023 , \2322 );
not \U$24647 ( \25024 , RIae798e0_154);
not \U$24648 ( \25025 , \12564 );
or \U$24649 ( \25026 , \25024 , \25025 );
or \U$24650 ( \25027 , \3071 , RIae798e0_154);
nand \U$24651 ( \25028 , \25026 , \25027 );
not \U$24652 ( \25029 , \25028 );
or \U$24653 ( \25030 , \25023 , \25029 );
nand \U$24654 ( \25031 , \24336 , \2341 );
nand \U$24655 ( \25032 , \25030 , \25031 );
or \U$24656 ( \25033 , \25022 , \25032 );
nand \U$24657 ( \25034 , \25022 , \25032 );
nand \U$24658 ( \25035 , \25033 , \25034 );
xor \U$24659 ( \25036 , \24313 , \24319 );
and \U$24660 ( \25037 , \25036 , \24329 );
and \U$24661 ( \25038 , \24313 , \24319 );
nor \U$24662 ( \25039 , \25037 , \25038 );
xor \U$24663 ( \25040 , \25035 , \25039 );
not \U$24664 ( \25041 , \9828 );
not \U$24665 ( \25042 , \24285 );
or \U$24666 ( \25043 , \25041 , \25042 );
not \U$24667 ( \25044 , \3039 );
not \U$24668 ( \25045 , \2309 );
or \U$24669 ( \25046 , \25044 , \25045 );
nand \U$24670 ( \25047 , \2305 , RIae794a8_145);
nand \U$24671 ( \25048 , \25046 , \25047 );
nand \U$24672 ( \25049 , \25048 , \1919 );
nand \U$24673 ( \25050 , \25043 , \25049 );
not \U$24674 ( \25051 , \2610 );
and \U$24675 ( \25052 , RIae79520_146, \1741 );
not \U$24676 ( \25053 , RIae79520_146);
and \U$24677 ( \25054 , \25053 , \4023 );
or \U$24678 ( \25055 , \25052 , \25054 );
not \U$24679 ( \25056 , \25055 );
or \U$24680 ( \25057 , \25051 , \25056 );
nand \U$24681 ( \25058 , \24447 , \2602 );
nand \U$24682 ( \25059 , \25057 , \25058 );
xor \U$24683 ( \25060 , \25050 , \25059 );
not \U$24684 ( \25061 , \14940 );
and \U$24685 ( \25062 , RIae79d90_164, \1118 );
not \U$24686 ( \25063 , RIae79d90_164);
and \U$24687 ( \25064 , \25063 , \2918 );
nor \U$24688 ( \25065 , \25062 , \25064 );
not \U$24689 ( \25066 , \25065 );
or \U$24690 ( \25067 , \25061 , \25066 );
nand \U$24691 ( \25068 , \24468 , \6091 );
nand \U$24692 ( \25069 , \25067 , \25068 );
not \U$24693 ( \25070 , \25069 );
xor \U$24694 ( \25071 , \25060 , \25070 );
xor \U$24695 ( \25072 , \25040 , \25071 );
xor \U$24696 ( \25073 , \25002 , \25072 );
not \U$24697 ( \25074 , \1864 );
and \U$24698 ( \25075 , RIae793b8_143, \1860 );
not \U$24699 ( \25076 , RIae793b8_143);
and \U$24700 ( \25077 , \25076 , \2385 );
or \U$24701 ( \25078 , \25075 , \25077 );
not \U$24702 ( \25079 , \25078 );
or \U$24703 ( \25080 , \25074 , \25079 );
nand \U$24704 ( \25081 , \24521 , \1910 );
nand \U$24705 ( \25082 , \25080 , \25081 );
not \U$24706 ( \25083 , \2011 );
not \U$24707 ( \25084 , \4113 );
not \U$24708 ( \25085 , RIae79610_148);
and \U$24709 ( \25086 , \25084 , \25085 );
and \U$24710 ( \25087 , \4113 , RIae79610_148);
nor \U$24711 ( \25088 , \25086 , \25087 );
not \U$24712 ( \25089 , \25088 );
not \U$24713 ( \25090 , \25089 );
or \U$24714 ( \25091 , \25083 , \25090 );
nand \U$24715 ( \25092 , \24327 , \2063 );
nand \U$24716 ( \25093 , \25091 , \25092 );
xor \U$24717 ( \25094 , \25082 , \25093 );
not \U$24718 ( \25095 , \13121 );
and \U$24719 ( \25096 , RIae7a240_174, \12522 );
not \U$24720 ( \25097 , RIae7a240_174);
and \U$24721 ( \25098 , \25097 , \827 );
nor \U$24722 ( \25099 , \25096 , \25098 );
not \U$24723 ( \25100 , \25099 );
or \U$24724 ( \25101 , \25095 , \25100 );
nand \U$24725 ( \25102 , \24346 , \9687 );
nand \U$24726 ( \25103 , \25101 , \25102 );
xor \U$24727 ( \25104 , \25094 , \25103 );
not \U$24728 ( \25105 , \3827 );
and \U$24729 ( \25106 , \3417 , RIae79688_149);
not \U$24730 ( \25107 , \3417 );
and \U$24731 ( \25108 , \25107 , \3147 );
or \U$24732 ( \25109 , \25106 , \25108 );
not \U$24733 ( \25110 , \25109 );
or \U$24734 ( \25111 , \25105 , \25110 );
nand \U$24735 ( \25112 , \24402 , \1844 );
nand \U$24736 ( \25113 , \25111 , \25112 );
and \U$24737 ( \25114 , \24457 , \2272 );
and \U$24738 ( \25115 , RIae79ac0_158, \2697 );
not \U$24739 ( \25116 , RIae79ac0_158);
and \U$24740 ( \25117 , \25116 , \3529 );
or \U$24741 ( \25118 , \25115 , \25117 );
and \U$24742 ( \25119 , \25118 , \3014 );
nor \U$24743 ( \25120 , \25114 , \25119 );
not \U$24744 ( \25121 , \25120 );
xor \U$24745 ( \25122 , \25113 , \25121 );
not \U$24746 ( \25123 , \4853 );
not \U$24747 ( \25124 , RIae79ca0_162);
not \U$24748 ( \25125 , \1186 );
or \U$24749 ( \25126 , \25124 , \25125 );
or \U$24750 ( \25127 , \1186 , RIae79ca0_162);
nand \U$24751 ( \25128 , \25126 , \25127 );
not \U$24752 ( \25129 , \25128 );
or \U$24753 ( \25130 , \25123 , \25129 );
nand \U$24754 ( \25131 , \24388 , \6276 );
nand \U$24755 ( \25132 , \25130 , \25131 );
xor \U$24756 ( \25133 , \25122 , \25132 );
xor \U$24757 ( \25134 , \25104 , \25133 );
not \U$24758 ( \25135 , \2450 );
and \U$24759 ( \25136 , \5944 , RIae79778_151);
not \U$24760 ( \25137 , \5944 );
and \U$24761 ( \25138 , \25137 , \2447 );
nor \U$24762 ( \25139 , \25136 , \25138 );
not \U$24763 ( \25140 , \25139 );
or \U$24764 ( \25141 , \25135 , \25140 );
nand \U$24765 ( \25142 , \9576 , \24434 );
nand \U$24766 ( \25143 , \25141 , \25142 );
not \U$24767 ( \25144 , \9518 );
and \U$24768 ( \25145 , \2471 , RIae79fe8_169);
not \U$24769 ( \25146 , \2471 );
and \U$24770 ( \25147 , \25146 , \11069 );
nor \U$24771 ( \25148 , \25145 , \25147 );
not \U$24772 ( \25149 , \25148 );
or \U$24773 ( \25150 , \25144 , \25149 );
nand \U$24774 ( \25151 , \24423 , \10709 );
nand \U$24775 ( \25152 , \25150 , \25151 );
xor \U$24776 ( \25153 , \25143 , \25152 );
not \U$24777 ( \25154 , \1989 );
not \U$24778 ( \25155 , \24358 );
or \U$24779 ( \25156 , \25154 , \25155 );
not \U$24780 ( \25157 , \2212 );
not \U$24781 ( \25158 , \1991 );
and \U$24782 ( \25159 , \25157 , \25158 );
and \U$24783 ( \25160 , \2629 , \1997 );
nor \U$24784 ( \25161 , \25159 , \25160 );
nand \U$24785 ( \25162 , \25161 , \2519 );
nand \U$24786 ( \25163 , \25156 , \25162 );
xor \U$24787 ( \25164 , \25153 , \25163 );
xor \U$24788 ( \25165 , \25134 , \25164 );
xnor \U$24789 ( \25166 , \25073 , \25165 );
xor \U$24790 ( \25167 , \24942 , \25166 );
not \U$24791 ( \25168 , \24500 );
nand \U$24792 ( \25169 , \25168 , \24505 , \24507 );
not \U$24793 ( \25170 , \24500 );
not \U$24794 ( \25171 , \24508 );
or \U$24795 ( \25172 , \25170 , \25171 );
nand \U$24796 ( \25173 , \25172 , \24569 );
nand \U$24797 ( \25174 , \25169 , \25173 );
xor \U$24798 ( \25175 , \25167 , \25174 );
not \U$24799 ( \25176 , \24278 );
not \U$24800 ( \25177 , \24270 );
not \U$24801 ( \25178 , \24271 );
or \U$24802 ( \25179 , \25177 , \25178 );
nand \U$24803 ( \25180 , \25179 , \24482 );
nand \U$24804 ( \25181 , \25176 , \25180 );
not \U$24805 ( \25182 , \24272 );
not \U$24806 ( \25183 , \24482 );
nand \U$24807 ( \25184 , \25182 , \25183 );
nand \U$24808 ( \25185 , \25181 , \25184 );
and \U$24809 ( \25186 , \25175 , \25185 );
not \U$24810 ( \25187 , \25175 );
not \U$24811 ( \25188 , \25185 );
and \U$24812 ( \25189 , \25187 , \25188 );
nor \U$24813 ( \25190 , \25186 , \25189 );
not \U$24814 ( \25191 , \25190 );
and \U$24815 ( \25192 , \24899 , \25191 );
and \U$24816 ( \25193 , \25190 , \24898 );
nor \U$24817 ( \25194 , \25192 , \25193 );
not \U$24818 ( \25195 , \25194 );
or \U$24819 ( \25196 , \24893 , \25195 );
or \U$24820 ( \25197 , \25194 , \24892 );
nand \U$24821 ( \25198 , \25196 , \25197 );
not \U$24822 ( \25199 , \25198 );
or \U$24823 ( \25200 , \24728 , \25199 );
not \U$24824 ( \25201 , \25194 );
nand \U$24825 ( \25202 , \25201 , \24892 );
nand \U$24826 ( \25203 , \25200 , \25202 );
not \U$24827 ( \25204 , \24897 );
not \U$24828 ( \25205 , \25190 );
or \U$24829 ( \25206 , \25204 , \25205 );
nand \U$24830 ( \25207 , \25175 , \25185 );
nand \U$24831 ( \25208 , \25206 , \25207 );
not \U$24832 ( \25209 , \24891 );
not \U$24833 ( \25210 , \24884 );
or \U$24834 ( \25211 , \25209 , \25210 );
not \U$24835 ( \25212 , \24781 );
nand \U$24836 ( \25213 , \24880 , \25212 );
nand \U$24837 ( \25214 , \25211 , \25213 );
and \U$24838 ( \25215 , \25208 , \25214 );
not \U$24839 ( \25216 , \25208 );
not \U$24840 ( \25217 , \25214 );
and \U$24841 ( \25218 , \25216 , \25217 );
nor \U$24842 ( \25219 , \25215 , \25218 );
xor \U$24843 ( \25220 , \24942 , \25166 );
and \U$24844 ( \25221 , \25220 , \25174 );
and \U$24845 ( \25222 , \24942 , \25166 );
or \U$24846 ( \25223 , \25221 , \25222 );
not \U$24847 ( \25224 , \1910 );
not \U$24848 ( \25225 , \25078 );
or \U$24849 ( \25226 , \25224 , \25225 );
not \U$24850 ( \25227 , RIae793b8_143);
not \U$24851 ( \25228 , \1970 );
or \U$24852 ( \25229 , \25227 , \25228 );
or \U$24853 ( \25230 , \1970 , RIae793b8_143);
nand \U$24854 ( \25231 , \25229 , \25230 );
nand \U$24855 ( \25232 , \25231 , \1863 );
nand \U$24856 ( \25233 , \25226 , \25232 );
not \U$24857 ( \25234 , RIae79610_148);
not \U$24858 ( \25235 , \5890 );
or \U$24859 ( \25236 , \25234 , \25235 );
or \U$24860 ( \25237 , \2785 , RIae79610_148);
nand \U$24861 ( \25238 , \25236 , \25237 );
not \U$24862 ( \25239 , \25238 );
not \U$24863 ( \25240 , \2011 );
or \U$24864 ( \25241 , \25239 , \25240 );
or \U$24865 ( \25242 , \25088 , \8320 );
nand \U$24866 ( \25243 , \25241 , \25242 );
xor \U$24867 ( \25244 , \25233 , \25243 );
not \U$24868 ( \25245 , \2767 );
not \U$24869 ( \25246 , \24964 );
or \U$24870 ( \25247 , \25245 , \25246 );
not \U$24871 ( \25248 , \10584 );
not \U$24872 ( \25249 , \3689 );
or \U$24873 ( \25250 , \25248 , \25249 );
nand \U$24874 ( \25251 , \6147 , RIae79c28_161);
nand \U$24875 ( \25252 , \25250 , \25251 );
not \U$24876 ( \25253 , \25252 );
or \U$24877 ( \25254 , \25253 , \2410 );
nand \U$24878 ( \25255 , \25247 , \25254 );
xor \U$24879 ( \25256 , \25244 , \25255 );
not \U$24880 ( \25257 , \2450 );
and \U$24881 ( \25258 , RIae79778_151, \2593 );
not \U$24882 ( \25259 , RIae79778_151);
and \U$24883 ( \25260 , \25259 , \2048 );
or \U$24884 ( \25261 , \25258 , \25260 );
not \U$24885 ( \25262 , \25261 );
or \U$24886 ( \25263 , \25257 , \25262 );
nand \U$24887 ( \25264 , \25139 , \9576 );
nand \U$24888 ( \25265 , \25263 , \25264 );
not \U$24889 ( \25266 , \9499 );
not \U$24890 ( \25267 , \25148 );
or \U$24891 ( \25268 , \25266 , \25267 );
not \U$24892 ( \25269 , RIae79fe8_169);
not \U$24893 ( \25270 , \2510 );
or \U$24894 ( \25271 , \25269 , \25270 );
or \U$24895 ( \25272 , \2331 , RIae79fe8_169);
nand \U$24896 ( \25273 , \25271 , \25272 );
nand \U$24897 ( \25274 , \25273 , \9517 );
nand \U$24898 ( \25275 , \25268 , \25274 );
xor \U$24899 ( \25276 , \25265 , \25275 );
not \U$24900 ( \25277 , \13130 );
not \U$24901 ( \25278 , \25099 );
or \U$24902 ( \25279 , \25277 , \25278 );
xor \U$24903 ( \25280 , RIae7a240_174, \991 );
nand \U$24904 ( \25281 , \25280 , \13121 );
nand \U$24905 ( \25282 , \25279 , \25281 );
xor \U$24906 ( \25283 , \25276 , \25282 );
xor \U$24907 ( \25284 , \25256 , \25283 );
not \U$24908 ( \25285 , \2322 );
not \U$24909 ( \25286 , \2334 );
not \U$24910 ( \25287 , \18384 );
or \U$24911 ( \25288 , \25286 , \25287 );
nand \U$24912 ( \25289 , \2993 , RIae798e0_154);
nand \U$24913 ( \25290 , \25288 , \25289 );
not \U$24914 ( \25291 , \25290 );
or \U$24915 ( \25292 , \25285 , \25291 );
nand \U$24916 ( \25293 , \25028 , \2341 );
nand \U$24917 ( \25294 , \25292 , \25293 );
not \U$24918 ( \25295 , \2529 );
not \U$24919 ( \25296 , \25161 );
or \U$24920 ( \25297 , \25295 , \25296 );
not \U$24921 ( \25298 , \2521 );
not \U$24922 ( \25299 , \1897 );
or \U$24923 ( \25300 , \25298 , \25299 );
or \U$24924 ( \25301 , \1898 , \2521 );
nand \U$24925 ( \25302 , \25300 , \25301 );
nand \U$24926 ( \25303 , \25302 , \2519 );
nand \U$24927 ( \25304 , \25297 , \25303 );
not \U$24928 ( \25305 , \11409 );
not \U$24929 ( \25306 , \25006 );
or \U$24930 ( \25307 , \25305 , \25306 );
and \U$24931 ( \25308 , RIae79ef8_167, \938 );
not \U$24932 ( \25309 , RIae79ef8_167);
and \U$24933 ( \25310 , \25309 , \18414 );
or \U$24934 ( \25311 , \25308 , \25310 );
nand \U$24935 ( \25312 , \25311 , \6214 );
nand \U$24936 ( \25313 , \25307 , \25312 );
and \U$24937 ( \25314 , \25304 , \25313 );
not \U$24938 ( \25315 , \25304 );
not \U$24939 ( \25316 , \25313 );
and \U$24940 ( \25317 , \25315 , \25316 );
nor \U$24941 ( \25318 , \25314 , \25317 );
xor \U$24942 ( \25319 , \25294 , \25318 );
xnor \U$24943 ( \25320 , \25284 , \25319 );
nor \U$24944 ( \25321 , \11195 , \860 );
not \U$24945 ( \25322 , \1129 );
not \U$24946 ( \25323 , \24952 );
or \U$24947 ( \25324 , \25322 , \25323 );
or \U$24948 ( \25325 , \16786 , RIae78b48_125);
nand \U$24949 ( \25326 , \19736 , RIae78b48_125);
nand \U$24950 ( \25327 , \25325 , \25326 , \2096 );
nand \U$24951 ( \25328 , \25324 , \25327 );
xor \U$24952 ( \25329 , \25321 , \25328 );
not \U$24953 ( \25330 , \951 );
not \U$24954 ( \25331 , \24809 );
or \U$24955 ( \25332 , \25330 , \25331 );
not \U$24956 ( \25333 , \15088 );
and \U$24957 ( \25334 , RIae78bc0_126, \25333 );
not \U$24958 ( \25335 , RIae78bc0_126);
and \U$24959 ( \25336 , \25335 , \15088 );
or \U$24960 ( \25337 , \25334 , \25336 );
nand \U$24961 ( \25338 , \25337 , \927 );
nand \U$24962 ( \25339 , \25332 , \25338 );
xor \U$24963 ( \25340 , \25329 , \25339 );
not \U$24964 ( \25341 , RIae7a600_182);
not \U$24965 ( \25342 , RIae7a510_180);
or \U$24966 ( \25343 , \25341 , \25342 );
nand \U$24967 ( \25344 , \25343 , RIae7a3a8_177);
not \U$24968 ( \25345 , \1499 );
not \U$24969 ( \25346 , \24744 );
or \U$24970 ( \25347 , \25345 , \25346 );
and \U$24971 ( \25348 , \2402 , \1503 );
not \U$24972 ( \25349 , \2402 );
and \U$24973 ( \25350 , \25349 , RIae79250_140);
nor \U$24974 ( \25351 , \25348 , \25350 );
nand \U$24975 ( \25352 , \25351 , \1501 );
nand \U$24976 ( \25353 , \25347 , \25352 );
xor \U$24977 ( \25354 , \25344 , \25353 );
not \U$24978 ( \25355 , \1009 );
and \U$24979 ( \25356 , RIae79160_138, \4960 );
not \U$24980 ( \25357 , RIae79160_138);
and \U$24981 ( \25358 , \25357 , \4972 );
or \U$24982 ( \25359 , \25356 , \25358 );
not \U$24983 ( \25360 , \25359 );
or \U$24984 ( \25361 , \25355 , \25360 );
not \U$24985 ( \25362 , RIae79160_138);
not \U$24986 ( \25363 , \4928 );
or \U$24987 ( \25364 , \25362 , \25363 );
or \U$24988 ( \25365 , \6238 , RIae79160_138);
nand \U$24989 ( \25366 , \25364 , \25365 );
nand \U$24990 ( \25367 , \25366 , \1209 );
nand \U$24991 ( \25368 , \25361 , \25367 );
xor \U$24992 ( \25369 , \25354 , \25368 );
xor \U$24993 ( \25370 , \25340 , \25369 );
not \U$24994 ( \25371 , \25121 );
not \U$24995 ( \25372 , \25132 );
or \U$24996 ( \25373 , \25371 , \25372 );
not \U$24997 ( \25374 , \25120 );
not \U$24998 ( \25375 , \25132 );
or \U$24999 ( \25376 , \25374 , \25375 );
or \U$25000 ( \25377 , \25120 , \25132 );
nand \U$25001 ( \25378 , \25376 , \25377 );
nand \U$25002 ( \25379 , \25378 , \25113 );
nand \U$25003 ( \25380 , \25373 , \25379 );
xnor \U$25004 ( \25381 , \25370 , \25380 );
not \U$25005 ( \25382 , \5950 );
not \U$25006 ( \25383 , \25055 );
or \U$25007 ( \25384 , \25382 , \25383 );
not \U$25008 ( \25385 , \2183 );
not \U$25009 ( \25386 , \3748 );
or \U$25010 ( \25387 , \25385 , \25386 );
nand \U$25011 ( \25388 , \2287 , RIae79520_146);
nand \U$25012 ( \25389 , \25387 , \25388 );
nand \U$25013 ( \25390 , \25389 , \10223 );
nand \U$25014 ( \25391 , \25384 , \25390 );
not \U$25015 ( \25392 , \2272 );
not \U$25016 ( \25393 , \25118 );
or \U$25017 ( \25394 , \25392 , \25393 );
and \U$25018 ( \25395 , RIae79ac0_158, \10605 );
not \U$25019 ( \25396 , RIae79ac0_158);
and \U$25020 ( \25397 , \25396 , \23358 );
nor \U$25021 ( \25398 , \25395 , \25397 );
nand \U$25022 ( \25399 , \25398 , \2252 );
nand \U$25023 ( \25400 , \25394 , \25399 );
xor \U$25024 ( \25401 , \25391 , \25400 );
not \U$25025 ( \25402 , \11761 );
not \U$25026 ( \25403 , \25128 );
or \U$25027 ( \25404 , \25402 , \25403 );
not \U$25028 ( \25405 , RIae79ca0_162);
not \U$25029 ( \25406 , \975 );
or \U$25030 ( \25407 , \25405 , \25406 );
or \U$25031 ( \25408 , \16510 , RIae79ca0_162);
nand \U$25032 ( \25409 , \25407 , \25408 );
nand \U$25033 ( \25410 , \25409 , \4853 );
nand \U$25034 ( \25411 , \25404 , \25410 );
xor \U$25035 ( \25412 , \25401 , \25411 );
xor \U$25036 ( \25413 , \25143 , \25152 );
and \U$25037 ( \25414 , \25413 , \25163 );
and \U$25038 ( \25415 , \25143 , \25152 );
or \U$25039 ( \25416 , \25414 , \25415 );
xor \U$25040 ( \25417 , \25412 , \25416 );
not \U$25041 ( \25418 , \6080 );
and \U$25042 ( \25419 , RIae79d90_164, \2175 );
not \U$25043 ( \25420 , RIae79d90_164);
and \U$25044 ( \25421 , \25420 , \883 );
or \U$25045 ( \25422 , \25419 , \25421 );
not \U$25046 ( \25423 , \25422 );
or \U$25047 ( \25424 , \25418 , \25423 );
nand \U$25048 ( \25425 , \25065 , \6091 );
nand \U$25049 ( \25426 , \25424 , \25425 );
xnor \U$25050 ( \25427 , RIae7a2b8_175, \1993 );
not \U$25051 ( \25428 , \25427 );
not \U$25052 ( \25429 , \9815 );
or \U$25053 ( \25430 , \25428 , \25429 );
nand \U$25054 ( \25431 , \25017 , \9792 );
nand \U$25055 ( \25432 , \25430 , \25431 );
xor \U$25056 ( \25433 , \25426 , \25432 );
not \U$25057 ( \25434 , \1919 );
not \U$25058 ( \25435 , \3039 );
not \U$25059 ( \25436 , \2955 );
or \U$25060 ( \25437 , \25435 , \25436 );
nand \U$25061 ( \25438 , \14712 , RIae794a8_145);
nand \U$25062 ( \25439 , \25437 , \25438 );
not \U$25063 ( \25440 , \25439 );
or \U$25064 ( \25441 , \25434 , \25440 );
nand \U$25065 ( \25442 , \25048 , \2458 );
nand \U$25066 ( \25443 , \25441 , \25442 );
xor \U$25067 ( \25444 , \25433 , \25443 );
xor \U$25068 ( \25445 , \25417 , \25444 );
xor \U$25069 ( \25446 , \25381 , \25445 );
xor \U$25070 ( \25447 , \25320 , \25446 );
not \U$25071 ( \25448 , \25165 );
not \U$25072 ( \25449 , \25002 );
not \U$25073 ( \25450 , \25072 );
xor \U$25074 ( \25451 , \25449 , \25450 );
not \U$25075 ( \25452 , \25451 );
or \U$25076 ( \25453 , \25448 , \25452 );
not \U$25077 ( \25454 , \25072 );
and \U$25078 ( \25455 , \25449 , \25454 );
not \U$25079 ( \25456 , \25455 );
nand \U$25080 ( \25457 , \25453 , \25456 );
xor \U$25081 ( \25458 , \25447 , \25457 );
not \U$25082 ( \25459 , \24839 );
not \U$25083 ( \25460 , \25459 );
not \U$25084 ( \25461 , \24866 );
or \U$25085 ( \25462 , \25460 , \25461 );
not \U$25086 ( \25463 , \24859 );
not \U$25087 ( \25464 , \24861 );
or \U$25088 ( \25465 , \25463 , \25464 );
nand \U$25089 ( \25466 , \25465 , \24852 );
nand \U$25090 ( \25467 , \25462 , \25466 );
not \U$25091 ( \25468 , \1822 );
and \U$25092 ( \25469 , \2758 , \21474 );
not \U$25093 ( \25470 , \2758 );
and \U$25094 ( \25471 , \25470 , RIae79688_149);
nor \U$25095 ( \25472 , \25469 , \25471 );
not \U$25096 ( \25473 , \25472 );
or \U$25097 ( \25474 , \25468 , \25473 );
nand \U$25098 ( \25475 , \25109 , \2966 );
nand \U$25099 ( \25476 , \25474 , \25475 );
xor \U$25100 ( \25477 , \24748 , \25476 );
xor \U$25101 ( \25478 , \24980 , \24989 );
and \U$25102 ( \25479 , \25478 , \24996 );
and \U$25103 ( \25480 , \24980 , \24989 );
or \U$25104 ( \25481 , \25479 , \25480 );
xor \U$25105 ( \25482 , \25477 , \25481 );
not \U$25106 ( \25483 , \24752 );
not \U$25107 ( \25484 , \24757 );
or \U$25108 ( \25485 , \25483 , \25484 );
not \U$25109 ( \25486 , \24748 );
nand \U$25110 ( \25487 , \25486 , \24737 );
nand \U$25111 ( \25488 , \25485 , \25487 );
xor \U$25112 ( \25489 , \25482 , \25488 );
not \U$25113 ( \25490 , \24927 );
not \U$25114 ( \25491 , \24912 );
or \U$25115 ( \25492 , \25490 , \25491 );
not \U$25116 ( \25493 , \24908 );
nand \U$25117 ( \25494 , \25493 , \24903 );
nand \U$25118 ( \25495 , \25492 , \25494 );
xor \U$25119 ( \25496 , \25489 , \25495 );
nand \U$25120 ( \25497 , \24733 , \24768 );
not \U$25121 ( \25498 , \24762 );
nand \U$25122 ( \25499 , \25498 , \24767 );
nand \U$25123 ( \25500 , \25497 , \25499 );
xor \U$25124 ( \25501 , \25496 , \25500 );
xor \U$25125 ( \25502 , \25467 , \25501 );
not \U$25126 ( \25503 , \25502 );
and \U$25127 ( \25504 , \25458 , \25503 );
not \U$25128 ( \25505 , \25458 );
and \U$25129 ( \25506 , \25505 , \25502 );
nor \U$25130 ( \25507 , \25504 , \25506 );
xor \U$25131 ( \25508 , \25223 , \25507 );
not \U$25132 ( \25509 , \24769 );
or \U$25133 ( \25510 , \24780 , \25509 );
nand \U$25134 ( \25511 , \25510 , \24775 );
nand \U$25135 ( \25512 , \24780 , \25509 );
and \U$25136 ( \25513 , \25511 , \25512 );
not \U$25137 ( \25514 , \25513 );
buf \U$25138 ( \25515 , \24797 );
not \U$25139 ( \25516 , \25515 );
buf \U$25140 ( \25517 , \24870 );
not \U$25141 ( \25518 , \25517 );
or \U$25142 ( \25519 , \25516 , \25518 );
or \U$25143 ( \25520 , \25517 , \25515 );
nand \U$25144 ( \25521 , \25520 , \24789 );
nand \U$25145 ( \25522 , \25519 , \25521 );
not \U$25146 ( \25523 , \25522 );
or \U$25147 ( \25524 , \25514 , \25523 );
or \U$25148 ( \25525 , \25522 , \25513 );
nand \U$25149 ( \25526 , \25524 , \25525 );
not \U$25150 ( \25527 , \25021 );
not \U$25151 ( \25528 , \25011 );
or \U$25152 ( \25529 , \25527 , \25528 );
nand \U$25153 ( \25530 , \25529 , \25034 );
not \U$25154 ( \25531 , \25530 );
not \U$25155 ( \25532 , \25531 );
not \U$25156 ( \25533 , \24824 );
xor \U$25157 ( \25534 , \24813 , \24830 );
not \U$25158 ( \25535 , \25534 );
or \U$25159 ( \25536 , \25533 , \25535 );
nand \U$25160 ( \25537 , \24813 , \24830 );
nand \U$25161 ( \25538 , \25536 , \25537 );
not \U$25162 ( \25539 , \25059 );
xor \U$25163 ( \25540 , \25069 , \25050 );
not \U$25164 ( \25541 , \25540 );
or \U$25165 ( \25542 , \25539 , \25541 );
not \U$25166 ( \25543 , \25070 );
nand \U$25167 ( \25544 , \25543 , \25050 );
nand \U$25168 ( \25545 , \25542 , \25544 );
and \U$25169 ( \25546 , \25538 , \25545 );
not \U$25170 ( \25547 , \25538 );
not \U$25171 ( \25548 , \25545 );
and \U$25172 ( \25549 , \25547 , \25548 );
nor \U$25173 ( \25550 , \25546 , \25549 );
not \U$25174 ( \25551 , \25550 );
or \U$25175 ( \25552 , \25532 , \25551 );
or \U$25176 ( \25553 , \25550 , \25531 );
nand \U$25177 ( \25554 , \25552 , \25553 );
or \U$25178 ( \25555 , \24969 , \24946 );
nand \U$25179 ( \25556 , \25555 , \24997 );
nand \U$25180 ( \25557 , \24946 , \24969 );
nand \U$25181 ( \25558 , \25556 , \25557 );
not \U$25182 ( \25559 , \25558 );
not \U$25183 ( \25560 , \24800 );
nor \U$25184 ( \25561 , \25560 , \24405 );
not \U$25185 ( \25562 , \25561 );
not \U$25186 ( \25563 , \24803 );
and \U$25187 ( \25564 , \25562 , \25563 );
nor \U$25188 ( \25565 , \25564 , \24831 );
not \U$25189 ( \25566 , \25565 );
not \U$25190 ( \25567 , \24804 );
not \U$25191 ( \25568 , \24831 );
or \U$25192 ( \25569 , \25567 , \25568 );
nand \U$25193 ( \25570 , \25569 , \24837 );
nand \U$25194 ( \25571 , \25566 , \25570 );
not \U$25195 ( \25572 , \25571 );
not \U$25196 ( \25573 , \25572 );
or \U$25197 ( \25574 , \25559 , \25573 );
not \U$25198 ( \25575 , \25558 );
nand \U$25199 ( \25576 , \25575 , \25571 );
nand \U$25200 ( \25577 , \25574 , \25576 );
xor \U$25201 ( \25578 , \25554 , \25577 );
not \U$25202 ( \25579 , \25578 );
xor \U$25203 ( \25580 , \24932 , \24937 );
and \U$25204 ( \25581 , \25580 , \24941 );
and \U$25205 ( \25582 , \24932 , \24937 );
or \U$25206 ( \25583 , \25581 , \25582 );
not \U$25207 ( \25584 , \25583 );
or \U$25208 ( \25585 , \25579 , \25584 );
or \U$25209 ( \25586 , \25583 , \25578 );
nand \U$25210 ( \25587 , \25585 , \25586 );
buf \U$25211 ( \25588 , \25587 );
xor \U$25212 ( \25589 , \25082 , \25093 );
and \U$25213 ( \25590 , \25589 , \25103 );
and \U$25214 ( \25591 , \25082 , \25093 );
or \U$25215 ( \25592 , \25590 , \25591 );
not \U$25216 ( \25593 , \797 );
not \U$25217 ( \25594 , \24976 );
or \U$25218 ( \25595 , \25593 , \25594 );
and \U$25219 ( \25596 , RIae78f80_134, \6346 );
not \U$25220 ( \25597 , RIae78f80_134);
and \U$25221 ( \25598 , \25597 , \9290 );
or \U$25222 ( \25599 , \25596 , \25598 );
nand \U$25223 ( \25600 , \25599 , \838 );
nand \U$25224 ( \25601 , \25595 , \25600 );
not \U$25225 ( \25602 , \5858 );
not \U$25226 ( \25603 , \24820 );
or \U$25227 ( \25604 , \25602 , \25603 );
and \U$25228 ( \25605 , RIae78e90_132, \9316 );
not \U$25229 ( \25606 , RIae78e90_132);
and \U$25230 ( \25607 , \25606 , \10386 );
or \U$25231 ( \25608 , \25605 , \25607 );
nand \U$25232 ( \25609 , \25608 , \1072 );
nand \U$25233 ( \25610 , \25604 , \25609 );
xor \U$25234 ( \25611 , \25601 , \25610 );
not \U$25235 ( \25612 , \1049 );
not \U$25236 ( \25613 , \1039 );
not \U$25237 ( \25614 , \24679 );
or \U$25238 ( \25615 , \25613 , \25614 );
nand \U$25239 ( \25616 , \15128 , RIae79070_136);
nand \U$25240 ( \25617 , \25615 , \25616 );
not \U$25241 ( \25618 , \25617 );
or \U$25242 ( \25619 , \25612 , \25618 );
nand \U$25243 ( \25620 , \24987 , \1062 );
nand \U$25244 ( \25621 , \25619 , \25620 );
xor \U$25245 ( \25622 , \25611 , \25621 );
xor \U$25246 ( \25623 , \24947 , \24957 );
and \U$25247 ( \25624 , \25623 , \24968 );
and \U$25248 ( \25625 , \24947 , \24957 );
or \U$25249 ( \25626 , \25624 , \25625 );
xor \U$25250 ( \25627 , \25622 , \25626 );
xor \U$25251 ( \25628 , \25592 , \25627 );
xor \U$25252 ( \25629 , \25035 , \25039 );
and \U$25253 ( \25630 , \25629 , \25071 );
and \U$25254 ( \25631 , \25035 , \25039 );
or \U$25255 ( \25632 , \25630 , \25631 );
not \U$25256 ( \25633 , \25632 );
xor \U$25257 ( \25634 , \25628 , \25633 );
xor \U$25258 ( \25635 , \25104 , \25133 );
and \U$25259 ( \25636 , \25635 , \25164 );
and \U$25260 ( \25637 , \25104 , \25133 );
or \U$25261 ( \25638 , \25636 , \25637 );
xor \U$25262 ( \25639 , \25634 , \25638 );
not \U$25263 ( \25640 , \25639 );
and \U$25264 ( \25641 , \25588 , \25640 );
not \U$25265 ( \25642 , \25588 );
and \U$25266 ( \25643 , \25642 , \25639 );
nor \U$25267 ( \25644 , \25641 , \25643 );
xor \U$25268 ( \25645 , \25526 , \25644 );
xor \U$25269 ( \25646 , \25508 , \25645 );
xor \U$25270 ( \25647 , \25219 , \25646 );
nand \U$25271 ( \25648 , \25203 , \25647 );
nor \U$25272 ( \25649 , \25198 , \24726 );
not \U$25273 ( \25650 , \25649 );
nand \U$25274 ( \25651 , \25198 , \24726 );
nand \U$25275 ( \25652 , \25650 , \25651 );
xor \U$25276 ( \25653 , \22605 , \22782 );
and \U$25277 ( \25654 , \25653 , \22792 );
and \U$25278 ( \25655 , \22605 , \22782 );
or \U$25279 ( \25656 , \25654 , \25655 );
xor \U$25280 ( \25657 , \22334 , \22583 );
and \U$25281 ( \25658 , \25657 , \22591 );
and \U$25282 ( \25659 , \22334 , \22583 );
or \U$25283 ( \25660 , \25658 , \25659 );
nand \U$25284 ( \25661 , \25656 , \25660 );
not \U$25285 ( \25662 , \25661 );
xor \U$25286 ( \25663 , \24265 , \24484 );
xor \U$25287 ( \25664 , \25663 , \24723 );
not \U$25288 ( \25665 , \25664 );
not \U$25289 ( \25666 , \25665 );
or \U$25290 ( \25667 , \25662 , \25666 );
nor \U$25291 ( \25668 , \25656 , \25660 );
not \U$25292 ( \25669 , \25668 );
nand \U$25293 ( \25670 , \25667 , \25669 );
nand \U$25294 ( \25671 , \25652 , \25670 );
not \U$25295 ( \25672 , \25646 );
not \U$25296 ( \25673 , \25219 );
or \U$25297 ( \25674 , \25672 , \25673 );
not \U$25298 ( \25675 , \25217 );
nand \U$25299 ( \25676 , \25675 , \25208 );
nand \U$25300 ( \25677 , \25674 , \25676 );
xor \U$25301 ( \25678 , \24748 , \25476 );
and \U$25302 ( \25679 , \25678 , \25481 );
and \U$25303 ( \25680 , \24748 , \25476 );
or \U$25304 ( \25681 , \25679 , \25680 );
not \U$25305 ( \25682 , \4853 );
not \U$25306 ( \25683 , RIae79ca0_162);
not \U$25307 ( \25684 , \1472 );
or \U$25308 ( \25685 , \25683 , \25684 );
or \U$25309 ( \25686 , \1119 , RIae79ca0_162);
nand \U$25310 ( \25687 , \25685 , \25686 );
not \U$25311 ( \25688 , \25687 );
or \U$25312 ( \25689 , \25682 , \25688 );
nand \U$25313 ( \25690 , \25409 , \6276 );
nand \U$25314 ( \25691 , \25689 , \25690 );
not \U$25315 ( \25692 , \2776 );
not \U$25316 ( \25693 , \10584 );
not \U$25317 ( \25694 , \3538 );
or \U$25318 ( \25695 , \25693 , \25694 );
nand \U$25319 ( \25696 , \1186 , RIae79c28_161);
nand \U$25320 ( \25697 , \25695 , \25696 );
not \U$25321 ( \25698 , \25697 );
or \U$25322 ( \25699 , \25692 , \25698 );
nand \U$25323 ( \25700 , \25252 , \2767 );
nand \U$25324 ( \25701 , \25699 , \25700 );
xor \U$25325 ( \25702 , \25691 , \25701 );
not \U$25326 ( \25703 , \2252 );
and \U$25327 ( \25704 , RIae79ac0_158, \4431 );
not \U$25328 ( \25705 , RIae79ac0_158);
and \U$25329 ( \25706 , \25705 , \1741 );
nor \U$25330 ( \25707 , \25704 , \25706 );
not \U$25331 ( \25708 , \25707 );
or \U$25332 ( \25709 , \25703 , \25708 );
nand \U$25333 ( \25710 , \25398 , \2272 );
nand \U$25334 ( \25711 , \25709 , \25710 );
xor \U$25335 ( \25712 , \25702 , \25711 );
xor \U$25336 ( \25713 , \25681 , \25712 );
or \U$25337 ( \25714 , \25610 , \25601 );
nand \U$25338 ( \25715 , \25714 , \25621 );
nand \U$25339 ( \25716 , \25610 , \25601 );
nand \U$25340 ( \25717 , \25715 , \25716 );
xor \U$25341 ( \25718 , \25321 , \25328 );
and \U$25342 ( \25719 , \25718 , \25339 );
and \U$25343 ( \25720 , \25321 , \25328 );
or \U$25344 ( \25721 , \25719 , \25720 );
xor \U$25345 ( \25722 , \25717 , \25721 );
xor \U$25346 ( \25723 , \25344 , \25353 );
and \U$25347 ( \25724 , \25723 , \25368 );
and \U$25348 ( \25725 , \25344 , \25353 );
or \U$25349 ( \25726 , \25724 , \25725 );
and \U$25350 ( \25727 , \25722 , \25726 );
not \U$25351 ( \25728 , \25722 );
not \U$25352 ( \25729 , \25726 );
and \U$25353 ( \25730 , \25728 , \25729 );
nor \U$25354 ( \25731 , \25727 , \25730 );
xor \U$25355 ( \25732 , \25713 , \25731 );
xor \U$25356 ( \25733 , \25482 , \25488 );
and \U$25357 ( \25734 , \25733 , \25495 );
and \U$25358 ( \25735 , \25482 , \25488 );
or \U$25359 ( \25736 , \25734 , \25735 );
not \U$25360 ( \25737 , \25736 );
xor \U$25361 ( \25738 , \25732 , \25737 );
not \U$25362 ( \25739 , \25554 );
not \U$25363 ( \25740 , \25577 );
or \U$25364 ( \25741 , \25739 , \25740 );
nand \U$25365 ( \25742 , \25571 , \25558 );
nand \U$25366 ( \25743 , \25741 , \25742 );
buf \U$25367 ( \25744 , \25743 );
xnor \U$25368 ( \25745 , \25738 , \25744 );
not \U$25369 ( \25746 , \25639 );
not \U$25370 ( \25747 , \25587 );
or \U$25371 ( \25748 , \25746 , \25747 );
not \U$25372 ( \25749 , \25583 );
nand \U$25373 ( \25750 , \25749 , \25578 );
nand \U$25374 ( \25751 , \25748 , \25750 );
xor \U$25375 ( \25752 , \25745 , \25751 );
xor \U$25376 ( \25753 , \25628 , \25633 );
and \U$25377 ( \25754 , \25753 , \25638 );
and \U$25378 ( \25755 , \25628 , \25633 );
or \U$25379 ( \25756 , \25754 , \25755 );
not \U$25380 ( \25757 , \25530 );
not \U$25381 ( \25758 , \25550 );
or \U$25382 ( \25759 , \25757 , \25758 );
not \U$25383 ( \25760 , \25548 );
nand \U$25384 ( \25761 , \25760 , \25538 );
nand \U$25385 ( \25762 , \25759 , \25761 );
not \U$25386 ( \25763 , \25762 );
not \U$25387 ( \25764 , \25592 );
not \U$25388 ( \25765 , \25627 );
or \U$25389 ( \25766 , \25764 , \25765 );
nand \U$25390 ( \25767 , \25622 , \25626 );
nand \U$25391 ( \25768 , \25766 , \25767 );
not \U$25392 ( \25769 , \25380 );
not \U$25393 ( \25770 , \25340 );
or \U$25394 ( \25771 , \25769 , \25770 );
or \U$25395 ( \25772 , \25380 , \25340 );
nand \U$25396 ( \25773 , \25772 , \25369 );
nand \U$25397 ( \25774 , \25771 , \25773 );
xnor \U$25398 ( \25775 , \25768 , \25774 );
not \U$25399 ( \25776 , \25775 );
or \U$25400 ( \25777 , \25763 , \25776 );
not \U$25401 ( \25778 , \25762 );
xor \U$25402 ( \25779 , \25768 , \25774 );
nand \U$25403 ( \25780 , \25778 , \25779 );
nand \U$25404 ( \25781 , \25777 , \25780 );
xor \U$25405 ( \25782 , \25756 , \25781 );
xor \U$25406 ( \25783 , \25412 , \25416 );
and \U$25407 ( \25784 , \25783 , \25444 );
and \U$25408 ( \25785 , \25412 , \25416 );
or \U$25409 ( \25786 , \25784 , \25785 );
not \U$25410 ( \25787 , \25294 );
not \U$25411 ( \25788 , \25318 );
or \U$25412 ( \25789 , \25787 , \25788 );
nand \U$25413 ( \25790 , \25304 , \25313 );
nand \U$25414 ( \25791 , \25789 , \25790 );
not \U$25415 ( \25792 , \2096 );
xor \U$25416 ( \25793 , RIae78b48_125, \12614 );
not \U$25417 ( \25794 , \25793 );
or \U$25418 ( \25795 , \25792 , \25794 );
not \U$25419 ( \25796 , RIae78b48_125);
nand \U$25420 ( \25797 , \25796 , \9456 );
nand \U$25421 ( \25798 , \25797 , \25326 , \893 );
nand \U$25422 ( \25799 , \25795 , \25798 );
not \U$25423 ( \25800 , \927 );
and \U$25424 ( \25801 , \21743 , RIae78bc0_126);
not \U$25425 ( \25802 , \21743 );
and \U$25426 ( \25803 , \25802 , \1286 );
nor \U$25427 ( \25804 , \25801 , \25803 );
not \U$25428 ( \25805 , \25804 );
or \U$25429 ( \25806 , \25800 , \25805 );
nand \U$25430 ( \25807 , \25337 , \952 );
nand \U$25431 ( \25808 , \25806 , \25807 );
not \U$25432 ( \25809 , \25808 );
xor \U$25433 ( \25810 , \25799 , \25809 );
not \U$25434 ( \25811 , \13130 );
not \U$25435 ( \25812 , \25280 );
or \U$25436 ( \25813 , \25811 , \25812 );
nand \U$25437 ( \25814 , \9699 , RIae7a240_174);
nand \U$25438 ( \25815 , \25813 , \25814 );
xor \U$25439 ( \25816 , \25810 , \25815 );
not \U$25440 ( \25817 , \25816 );
xor \U$25441 ( \25818 , \25233 , \25243 );
and \U$25442 ( \25819 , \25818 , \25255 );
and \U$25443 ( \25820 , \25233 , \25243 );
or \U$25444 ( \25821 , \25819 , \25820 );
not \U$25445 ( \25822 , \25821 );
or \U$25446 ( \25823 , \25817 , \25822 );
or \U$25447 ( \25824 , \25816 , \25821 );
nand \U$25448 ( \25825 , \25823 , \25824 );
xor \U$25449 ( \25826 , \25791 , \25825 );
xor \U$25450 ( \25827 , \25786 , \25826 );
or \U$25451 ( \25828 , \25319 , \25283 );
nand \U$25452 ( \25829 , \25828 , \25256 );
nand \U$25453 ( \25830 , \25319 , \25283 );
nand \U$25454 ( \25831 , \25829 , \25830 );
xnor \U$25455 ( \25832 , \25827 , \25831 );
not \U$25456 ( \25833 , \25832 );
xnor \U$25457 ( \25834 , \25782 , \25833 );
xor \U$25458 ( \25835 , \25752 , \25834 );
xor \U$25459 ( \25836 , \25223 , \25507 );
and \U$25460 ( \25837 , \25836 , \25645 );
and \U$25461 ( \25838 , \25223 , \25507 );
or \U$25462 ( \25839 , \25837 , \25838 );
xor \U$25463 ( \25840 , \25835 , \25839 );
xor \U$25464 ( \25841 , \25588 , \25639 );
not \U$25465 ( \25842 , \25841 );
not \U$25466 ( \25843 , \25526 );
or \U$25467 ( \25844 , \25842 , \25843 );
not \U$25468 ( \25845 , \25513 );
nand \U$25469 ( \25846 , \25845 , \25522 );
nand \U$25470 ( \25847 , \25844 , \25846 );
not \U$25471 ( \25848 , \25502 );
not \U$25472 ( \25849 , \25458 );
or \U$25473 ( \25850 , \25848 , \25849 );
nand \U$25474 ( \25851 , \25457 , \25447 );
nand \U$25475 ( \25852 , \25850 , \25851 );
not \U$25476 ( \25853 , \25852 );
not \U$25477 ( \25854 , \25501 );
not \U$25478 ( \25855 , \25467 );
or \U$25479 ( \25856 , \25854 , \25855 );
not \U$25480 ( \25857 , \25499 );
not \U$25481 ( \25858 , \25497 );
or \U$25482 ( \25859 , \25857 , \25858 );
nand \U$25483 ( \25860 , \25859 , \25496 );
nand \U$25484 ( \25861 , \25856 , \25860 );
not \U$25485 ( \25862 , \1320 );
and \U$25486 ( \25863 , RIae78e90_132, \6232 );
not \U$25487 ( \25864 , RIae78e90_132);
and \U$25488 ( \25865 , \25864 , \9299 );
nor \U$25489 ( \25866 , \25863 , \25865 );
not \U$25490 ( \25867 , \25866 );
or \U$25491 ( \25868 , \25862 , \25867 );
nand \U$25492 ( \25869 , \25608 , \5858 );
nand \U$25493 ( \25870 , \25868 , \25869 );
not \U$25494 ( \25871 , \839 );
and \U$25495 ( \25872 , RIae78f80_134, \12334 );
not \U$25496 ( \25873 , RIae78f80_134);
and \U$25497 ( \25874 , \25873 , \5722 );
or \U$25498 ( \25875 , \25872 , \25874 );
not \U$25499 ( \25876 , \25875 );
or \U$25500 ( \25877 , \25871 , \25876 );
nand \U$25501 ( \25878 , \25599 , \797 );
nand \U$25502 ( \25879 , \25877 , \25878 );
xor \U$25503 ( \25880 , \25870 , \25879 );
not \U$25504 ( \25881 , \1049 );
xnor \U$25505 ( \25882 , \4960 , RIae79070_136);
not \U$25506 ( \25883 , \25882 );
or \U$25507 ( \25884 , \25881 , \25883 );
nand \U$25508 ( \25885 , \25617 , \1062 );
nand \U$25509 ( \25886 , \25884 , \25885 );
xor \U$25510 ( \25887 , \25880 , \25886 );
xor \U$25511 ( \25888 , \25391 , \25400 );
and \U$25512 ( \25889 , \25888 , \25411 );
and \U$25513 ( \25890 , \25391 , \25400 );
or \U$25514 ( \25891 , \25889 , \25890 );
xor \U$25515 ( \25892 , \25887 , \25891 );
xor \U$25516 ( \25893 , \25426 , \25432 );
and \U$25517 ( \25894 , \25893 , \25443 );
and \U$25518 ( \25895 , \25426 , \25432 );
or \U$25519 ( \25896 , \25894 , \25895 );
xor \U$25520 ( \25897 , \25892 , \25896 );
not \U$25521 ( \25898 , \25265 );
not \U$25522 ( \25899 , \25282 );
or \U$25523 ( \25900 , \25898 , \25899 );
or \U$25524 ( \25901 , \25282 , \25265 );
nand \U$25525 ( \25902 , \25901 , \25275 );
nand \U$25526 ( \25903 , \25900 , \25902 );
not \U$25527 ( \25904 , \2011 );
not \U$25528 ( \25905 , \2056 );
not \U$25529 ( \25906 , \11512 );
or \U$25530 ( \25907 , \25905 , \25906 );
nand \U$25531 ( \25908 , \2676 , RIae79610_148);
nand \U$25532 ( \25909 , \25907 , \25908 );
not \U$25533 ( \25910 , \25909 );
or \U$25534 ( \25911 , \25904 , \25910 );
nand \U$25535 ( \25912 , \25238 , \2063 );
nand \U$25536 ( \25913 , \25911 , \25912 );
not \U$25537 ( \25914 , \25913 );
not \U$25538 ( \25915 , \25914 );
not \U$25539 ( \25916 , \2157 );
not \U$25540 ( \25917 , \25366 );
or \U$25541 ( \25918 , \25916 , \25917 );
and \U$25542 ( \25919 , RIae79160_138, \3207 );
not \U$25543 ( \25920 , RIae79160_138);
and \U$25544 ( \25921 , \25920 , \19325 );
nor \U$25545 ( \25922 , \25919 , \25921 );
nand \U$25546 ( \25923 , \25922 , \10451 );
nand \U$25547 ( \25924 , \25918 , \25923 );
not \U$25548 ( \25925 , \25924 );
not \U$25549 ( \25926 , \25925 );
or \U$25550 ( \25927 , \25915 , \25926 );
nand \U$25551 ( \25928 , \25924 , \25913 );
nand \U$25552 ( \25929 , \25927 , \25928 );
not \U$25553 ( \25930 , \1844 );
not \U$25554 ( \25931 , \25472 );
or \U$25555 ( \25932 , \25930 , \25931 );
not \U$25556 ( \25933 , \3147 );
not \U$25557 ( \25934 , \10884 );
or \U$25558 ( \25935 , \25933 , \25934 );
nand \U$25559 ( \25936 , \2697 , RIae79688_149);
nand \U$25560 ( \25937 , \25935 , \25936 );
nand \U$25561 ( \25938 , \25937 , \1822 );
nand \U$25562 ( \25939 , \25932 , \25938 );
xnor \U$25563 ( \25940 , \25929 , \25939 );
xor \U$25564 ( \25941 , \25903 , \25940 );
not \U$25565 ( \25942 , \10573 );
not \U$25566 ( \25943 , RIae79ef8_167);
not \U$25567 ( \25944 , \5958 );
or \U$25568 ( \25945 , \25943 , \25944 );
nand \U$25569 ( \25946 , \918 , \6207 );
nand \U$25570 ( \25947 , \25945 , \25946 );
not \U$25571 ( \25948 , \25947 );
or \U$25572 ( \25949 , \25942 , \25948 );
nand \U$25573 ( \25950 , \25311 , \6201 );
nand \U$25574 ( \25951 , \25949 , \25950 );
not \U$25575 ( \25952 , \5049 );
xor \U$25576 ( \25953 , \854 , RIae79d90_164);
not \U$25577 ( \25954 , \25953 );
or \U$25578 ( \25955 , \25952 , \25954 );
nand \U$25579 ( \25956 , \25422 , \6091 );
nand \U$25580 ( \25957 , \25955 , \25956 );
xor \U$25581 ( \25958 , \25951 , \25957 );
not \U$25582 ( \25959 , \10807 );
not \U$25583 ( \25960 , \25290 );
or \U$25584 ( \25961 , \25959 , \25960 );
not \U$25585 ( \25962 , RIae798e0_154);
not \U$25586 ( \25963 , \19373 );
or \U$25587 ( \25964 , \25962 , \25963 );
nand \U$25588 ( \25965 , \2207 , \2334 );
nand \U$25589 ( \25966 , \25964 , \25965 );
nand \U$25590 ( \25967 , \25966 , \2322 );
nand \U$25591 ( \25968 , \25961 , \25967 );
xnor \U$25592 ( \25969 , \25958 , \25968 );
xor \U$25593 ( \25970 , \25941 , \25969 );
xor \U$25594 ( \25971 , \25897 , \25970 );
not \U$25595 ( \25972 , \1501 );
and \U$25596 ( \25973 , RIae79250_140, \1859 );
not \U$25597 ( \25974 , RIae79250_140);
and \U$25598 ( \25975 , \25974 , \12502 );
or \U$25599 ( \25976 , \25973 , \25975 );
not \U$25600 ( \25977 , \25976 );
or \U$25601 ( \25978 , \25972 , \25977 );
nand \U$25602 ( \25979 , \25351 , \9403 );
nand \U$25603 ( \25980 , \25978 , \25979 );
not \U$25604 ( \25981 , \2007 );
and \U$25605 ( \25982 , RIae797f0_152, \1878 );
not \U$25606 ( \25983 , RIae797f0_152);
and \U$25607 ( \25984 , \25983 , \5944 );
or \U$25608 ( \25985 , \25982 , \25984 );
not \U$25609 ( \25986 , \25985 );
or \U$25610 ( \25987 , \25981 , \25986 );
nand \U$25611 ( \25988 , \25302 , \1988 );
nand \U$25612 ( \25989 , \25987 , \25988 );
xor \U$25613 ( \25990 , \25980 , \25989 );
not \U$25614 ( \25991 , \9814 );
not \U$25615 ( \25992 , RIae7a2b8_175);
not \U$25616 ( \25993 , \827 );
or \U$25617 ( \25994 , \25992 , \25993 );
or \U$25618 ( \25995 , \834 , RIae7a2b8_175);
nand \U$25619 ( \25996 , \25994 , \25995 );
not \U$25620 ( \25997 , \25996 );
or \U$25621 ( \25998 , \25991 , \25997 );
not \U$25622 ( \25999 , RIae7a2b8_175);
not \U$25623 ( \26000 , \1993 );
or \U$25624 ( \26001 , \25999 , \26000 );
or \U$25625 ( \26002 , \1993 , RIae7a2b8_175);
nand \U$25626 ( \26003 , \26001 , \26002 );
nand \U$25627 ( \26004 , \26003 , \9792 );
nand \U$25628 ( \26005 , \25998 , \26004 );
xor \U$25629 ( \26006 , \25990 , \26005 );
not \U$25630 ( \26007 , \1864 );
not \U$25631 ( \26008 , \1884 );
not \U$25632 ( \26009 , \5912 );
or \U$25633 ( \26010 , \26008 , \26009 );
nand \U$25634 ( \26011 , \4113 , RIae793b8_143);
nand \U$25635 ( \26012 , \26010 , \26011 );
not \U$25636 ( \26013 , \26012 );
or \U$25637 ( \26014 , \26007 , \26013 );
nand \U$25638 ( \26015 , \25231 , \1910 );
nand \U$25639 ( \26016 , \26014 , \26015 );
not \U$25640 ( \26017 , \19422 );
nand \U$25641 ( \26018 , \26017 , RIae78b48_125);
not \U$25642 ( \26019 , \26018 );
not \U$25643 ( \26020 , \2545 );
not \U$25644 ( \26021 , \25261 );
or \U$25645 ( \26022 , \26020 , \26021 );
and \U$25646 ( \26023 , RIae79778_151, \2026 );
not \U$25647 ( \26024 , RIae79778_151);
and \U$25648 ( \26025 , \26024 , \14071 );
or \U$25649 ( \26026 , \26023 , \26025 );
nand \U$25650 ( \26027 , \26026 , \11037 );
nand \U$25651 ( \26028 , \26022 , \26027 );
not \U$25652 ( \26029 , \26028 );
or \U$25653 ( \26030 , \26019 , \26029 );
or \U$25654 ( \26031 , \26028 , \26018 );
nand \U$25655 ( \26032 , \26030 , \26031 );
xor \U$25656 ( \26033 , \26016 , \26032 );
xor \U$25657 ( \26034 , \26006 , \26033 );
not \U$25658 ( \26035 , \1919 );
not \U$25659 ( \26036 , \3039 );
not \U$25660 ( \26037 , \2142 );
or \U$25661 ( \26038 , \26036 , \26037 );
not \U$25662 ( \26039 , \4081 );
nand \U$25663 ( \26040 , \26039 , RIae794a8_145);
nand \U$25664 ( \26041 , \26038 , \26040 );
not \U$25665 ( \26042 , \26041 );
or \U$25666 ( \26043 , \26035 , \26042 );
nand \U$25667 ( \26044 , \25439 , \2458 );
nand \U$25668 ( \26045 , \26043 , \26044 );
not \U$25669 ( \26046 , \2189 );
not \U$25670 ( \26047 , \25389 );
or \U$25671 ( \26048 , \26046 , \26047 );
and \U$25672 ( \26049 , RIae79520_146, \2305 );
not \U$25673 ( \26050 , RIae79520_146);
and \U$25674 ( \26051 , \26050 , \2309 );
or \U$25675 ( \26052 , \26049 , \26051 );
nand \U$25676 ( \26053 , \26052 , \2163 );
nand \U$25677 ( \26054 , \26048 , \26053 );
not \U$25678 ( \26055 , \10700 );
and \U$25679 ( \26056 , RIae79fe8_169, \3999 );
not \U$25680 ( \26057 , RIae79fe8_169);
and \U$25681 ( \26058 , \26057 , \1141 );
or \U$25682 ( \26059 , \26056 , \26058 );
not \U$25683 ( \26060 , \26059 );
or \U$25684 ( \26061 , \26055 , \26060 );
nand \U$25685 ( \26062 , \25273 , \11914 );
nand \U$25686 ( \26063 , \26061 , \26062 );
xor \U$25687 ( \26064 , \26054 , \26063 );
xor \U$25688 ( \26065 , \26045 , \26064 );
xor \U$25689 ( \26066 , \26034 , \26065 );
xor \U$25690 ( \26067 , \25971 , \26066 );
not \U$25691 ( \26068 , \26067 );
not \U$25692 ( \26069 , \25445 );
not \U$25693 ( \26070 , \26069 );
not \U$25694 ( \26071 , \25381 );
or \U$25695 ( \26072 , \26070 , \26071 );
or \U$25696 ( \26073 , \25381 , \26069 );
nand \U$25697 ( \26074 , \26073 , \25320 );
nand \U$25698 ( \26075 , \26072 , \26074 );
not \U$25699 ( \26076 , \26075 );
or \U$25700 ( \26077 , \26068 , \26076 );
or \U$25701 ( \26078 , \26075 , \26067 );
nand \U$25702 ( \26079 , \26077 , \26078 );
xnor \U$25703 ( \26080 , \25861 , \26079 );
not \U$25704 ( \26081 , \26080 );
and \U$25705 ( \26082 , \25853 , \26081 );
and \U$25706 ( \26083 , \25852 , \26080 );
nor \U$25707 ( \26084 , \26082 , \26083 );
xor \U$25708 ( \26085 , \25847 , \26084 );
xor \U$25709 ( \26086 , \25840 , \26085 );
nand \U$25710 ( \26087 , \25677 , \26086 );
or \U$25711 ( \26088 , \22592 , \22793 );
nand \U$25712 ( \26089 , \26088 , \22600 );
nand \U$25713 ( \26090 , \22793 , \22592 );
nand \U$25714 ( \26091 , \26089 , \26090 );
not \U$25715 ( \26092 , \26091 );
not \U$25716 ( \26093 , \25668 );
nand \U$25717 ( \26094 , \26093 , \25661 );
and \U$25718 ( \26095 , \26094 , \25665 );
not \U$25719 ( \26096 , \26094 );
and \U$25720 ( \26097 , \26096 , \25664 );
nor \U$25721 ( \26098 , \26095 , \26097 );
not \U$25722 ( \26099 , \26098 );
nand \U$25723 ( \26100 , \26092 , \26099 );
and \U$25724 ( \26101 , \25648 , \25671 , \26087 , \26100 );
not \U$25725 ( \26102 , \25762 );
not \U$25726 ( \26103 , \25779 );
or \U$25727 ( \26104 , \26102 , \26103 );
nand \U$25728 ( \26105 , \25774 , \25768 );
nand \U$25729 ( \26106 , \26104 , \26105 );
not \U$25730 ( \26107 , \1501 );
and \U$25731 ( \26108 , RIae79250_140, \3217 );
not \U$25732 ( \26109 , RIae79250_140);
and \U$25733 ( \26110 , \26109 , \1969 );
nor \U$25734 ( \26111 , \26108 , \26110 );
not \U$25735 ( \26112 , \26111 );
or \U$25736 ( \26113 , \26107 , \26112 );
nand \U$25737 ( \26114 , \25976 , \1499 );
nand \U$25738 ( \26115 , \26113 , \26114 );
not \U$25739 ( \26116 , \1910 );
not \U$25740 ( \26117 , \26012 );
or \U$25741 ( \26118 , \26116 , \26117 );
not \U$25742 ( \26119 , \2786 );
and \U$25743 ( \26120 , RIae793b8_143, \26119 );
not \U$25744 ( \26121 , RIae793b8_143);
and \U$25745 ( \26122 , \26121 , \2090 );
nor \U$25746 ( \26123 , \26120 , \26122 );
nand \U$25747 ( \26124 , \26123 , \1864 );
nand \U$25748 ( \26125 , \26118 , \26124 );
xor \U$25749 ( \26126 , \26115 , \26125 );
not \U$25750 ( \26127 , \9792 );
not \U$25751 ( \26128 , \25996 );
or \U$25752 ( \26129 , \26127 , \26128 );
not \U$25753 ( \26130 , \9804 );
not \U$25754 ( \26131 , \992 );
or \U$25755 ( \26132 , \26130 , \26131 );
or \U$25756 ( \26133 , \992 , \9810 );
nand \U$25757 ( \26134 , \26132 , \26133 );
nand \U$25758 ( \26135 , \26134 , \9814 );
nand \U$25759 ( \26136 , \26129 , \26135 );
xor \U$25760 ( \26137 , \26126 , \26136 );
not \U$25761 ( \26138 , \11914 );
not \U$25762 ( \26139 , \26059 );
or \U$25763 ( \26140 , \26138 , \26139 );
and \U$25764 ( \26141 , RIae79fe8_169, \780 );
not \U$25765 ( \26142 , RIae79fe8_169);
and \U$25766 ( \26143 , \26142 , \1994 );
or \U$25767 ( \26144 , \26141 , \26143 );
nand \U$25768 ( \26145 , \26144 , \9517 );
nand \U$25769 ( \26146 , \26140 , \26145 );
not \U$25770 ( \26147 , \6091 );
not \U$25771 ( \26148 , \25953 );
or \U$25772 ( \26149 , \26147 , \26148 );
and \U$25773 ( \26150 , \3236 , RIae79d90_164);
not \U$25774 ( \26151 , \3236 );
and \U$25775 ( \26152 , \26151 , \10900 );
nor \U$25776 ( \26153 , \26150 , \26152 );
nand \U$25777 ( \26154 , \26153 , \5049 );
nand \U$25778 ( \26155 , \26149 , \26154 );
xor \U$25779 ( \26156 , \26146 , \26155 );
not \U$25780 ( \26157 , \2458 );
not \U$25781 ( \26158 , \26041 );
or \U$25782 ( \26159 , \26157 , \26158 );
not \U$25783 ( \26160 , \3039 );
not \U$25784 ( \26161 , \11056 );
or \U$25785 ( \26162 , \26160 , \26161 );
not \U$25786 ( \26163 , \2994 );
nand \U$25787 ( \26164 , \26163 , RIae794a8_145);
nand \U$25788 ( \26165 , \26162 , \26164 );
nand \U$25789 ( \26166 , \26165 , \1919 );
nand \U$25790 ( \26167 , \26159 , \26166 );
xor \U$25791 ( \26168 , \26156 , \26167 );
xor \U$25792 ( \26169 , \26137 , \26168 );
not \U$25793 ( \26170 , \25726 );
not \U$25794 ( \26171 , \25722 );
or \U$25795 ( \26172 , \26170 , \26171 );
not \U$25796 ( \26173 , \25716 );
not \U$25797 ( \26174 , \25715 );
or \U$25798 ( \26175 , \26173 , \26174 );
nand \U$25799 ( \26176 , \26175 , \25721 );
nand \U$25800 ( \26177 , \26172 , \26176 );
xor \U$25801 ( \26178 , \26169 , \26177 );
xor \U$25802 ( \26179 , \25681 , \25712 );
and \U$25803 ( \26180 , \26179 , \25731 );
and \U$25804 ( \26181 , \25681 , \25712 );
or \U$25805 ( \26182 , \26180 , \26181 );
xor \U$25806 ( \26183 , \26178 , \26182 );
and \U$25807 ( \26184 , \26106 , \26183 );
and \U$25808 ( \26185 , \26178 , \26182 );
nor \U$25809 ( \26186 , \26184 , \26185 );
xor \U$25810 ( \26187 , \25980 , \25989 );
and \U$25811 ( \26188 , \26187 , \26005 );
and \U$25812 ( \26189 , \25980 , \25989 );
or \U$25813 ( \26190 , \26188 , \26189 );
or \U$25814 ( \26191 , \25968 , \25951 );
nand \U$25815 ( \26192 , \26191 , \25957 );
nand \U$25816 ( \26193 , \25968 , \25951 );
nand \U$25817 ( \26194 , \26192 , \26193 );
xor \U$25818 ( \26195 , \26190 , \26194 );
not \U$25819 ( \26196 , \25939 );
not \U$25820 ( \26197 , \25929 );
or \U$25821 ( \26198 , \26196 , \26197 );
buf \U$25822 ( \26199 , \25925 );
nand \U$25823 ( \26200 , \26199 , \25913 );
nand \U$25824 ( \26201 , \26198 , \26200 );
xor \U$25825 ( \26202 , \26195 , \26201 );
not \U$25826 ( \26203 , \26202 );
not \U$25827 ( \26204 , \26203 );
not \U$25828 ( \26205 , \2450 );
and \U$25829 ( \26206 , RIae79778_151, \1834 );
not \U$25830 ( \26207 , RIae79778_151);
and \U$25831 ( \26208 , \26207 , \2848 );
or \U$25832 ( \26209 , \26206 , \26208 );
not \U$25833 ( \26210 , \26209 );
or \U$25834 ( \26211 , \26205 , \26210 );
nand \U$25835 ( \26212 , \26026 , \2433 );
nand \U$25836 ( \26213 , \26211 , \26212 );
not \U$25837 ( \26214 , \25326 );
not \U$25838 ( \26215 , \26214 );
nand \U$25839 ( \26216 , \25793 , \1129 );
xor \U$25840 ( \26217 , RIae78b48_125, \14691 );
nand \U$25841 ( \26218 , \26217 , \2096 );
nand \U$25842 ( \26219 , \26216 , \26218 );
not \U$25843 ( \26220 , \26219 );
not \U$25844 ( \26221 , \26220 );
or \U$25845 ( \26222 , \26215 , \26221 );
not \U$25846 ( \26223 , \26218 );
not \U$25847 ( \26224 , \26216 );
or \U$25848 ( \26225 , \26223 , \26224 );
nand \U$25849 ( \26226 , \26225 , \25326 );
nand \U$25850 ( \26227 , \26222 , \26226 );
not \U$25851 ( \26228 , \26227 );
and \U$25852 ( \26229 , \26213 , \26228 );
not \U$25853 ( \26230 , \26213 );
and \U$25854 ( \26231 , \26230 , \26227 );
nor \U$25855 ( \26232 , \26229 , \26231 );
not \U$25856 ( \26233 , \26232 );
not \U$25857 ( \26234 , \952 );
not \U$25858 ( \26235 , \25804 );
or \U$25859 ( \26236 , \26234 , \26235 );
and \U$25860 ( \26237 , RIae78bc0_126, \9316 );
not \U$25861 ( \26238 , RIae78bc0_126);
and \U$25862 ( \26239 , \26238 , \10386 );
or \U$25863 ( \26240 , \26237 , \26239 );
nand \U$25864 ( \26241 , \26240 , \927 );
nand \U$25865 ( \26242 , \26236 , \26241 );
not \U$25866 ( \26243 , \1086 );
not \U$25867 ( \26244 , \25866 );
or \U$25868 ( \26245 , \26243 , \26244 );
not \U$25869 ( \26246 , RIae78e90_132);
not \U$25870 ( \26247 , \9286 );
or \U$25871 ( \26248 , \26246 , \26247 );
or \U$25872 ( \26249 , \14630 , RIae78e90_132);
nand \U$25873 ( \26250 , \26248 , \26249 );
nand \U$25874 ( \26251 , \1320 , \26250 );
nand \U$25875 ( \26252 , \26245 , \26251 );
not \U$25876 ( \26253 , \838 );
not \U$25877 ( \26254 , \3105 );
not \U$25878 ( \26255 , \6256 );
or \U$25879 ( \26256 , \26254 , \26255 );
nand \U$25880 ( \26257 , \5108 , RIae78f80_134);
nand \U$25881 ( \26258 , \26256 , \26257 );
not \U$25882 ( \26259 , \26258 );
or \U$25883 ( \26260 , \26253 , \26259 );
nand \U$25884 ( \26261 , \25875 , \796 );
nand \U$25885 ( \26262 , \26260 , \26261 );
xor \U$25886 ( \26263 , \26252 , \26262 );
xor \U$25887 ( \26264 , \26242 , \26263 );
not \U$25888 ( \26265 , \26264 );
and \U$25889 ( \26266 , \26233 , \26265 );
and \U$25890 ( \26267 , \26264 , \26232 );
nor \U$25891 ( \26268 , \26266 , \26267 );
not \U$25892 ( \26269 , \25711 );
not \U$25893 ( \26270 , \25702 );
or \U$25894 ( \26271 , \26269 , \26270 );
nand \U$25895 ( \26272 , \25701 , \25691 );
nand \U$25896 ( \26273 , \26271 , \26272 );
xor \U$25897 ( \26274 , \26268 , \26273 );
not \U$25898 ( \26275 , \26274 );
or \U$25899 ( \26276 , \26204 , \26275 );
not \U$25900 ( \26277 , \1843 );
not \U$25901 ( \26278 , \25937 );
or \U$25902 ( \26279 , \26277 , \26278 );
xor \U$25903 ( \26280 , \10605 , RIae79688_149);
nand \U$25904 ( \26281 , \26280 , \1821 );
nand \U$25905 ( \26282 , \26279 , \26281 );
not \U$25906 ( \26283 , \2011 );
not \U$25907 ( \26284 , RIae79610_148);
not \U$25908 ( \26285 , \2577 );
or \U$25909 ( \26286 , \26284 , \26285 );
nand \U$25910 ( \26287 , \10891 , \2056 );
nand \U$25911 ( \26288 , \26286 , \26287 );
not \U$25912 ( \26289 , \26288 );
or \U$25913 ( \26290 , \26283 , \26289 );
nand \U$25914 ( \26291 , \25909 , \2063 );
nand \U$25915 ( \26292 , \26290 , \26291 );
xor \U$25916 ( \26293 , \26282 , \26292 );
not \U$25917 ( \26294 , \2767 );
not \U$25918 ( \26295 , \25697 );
or \U$25919 ( \26296 , \26294 , \26295 );
and \U$25920 ( \26297 , \16510 , \10584 );
not \U$25921 ( \26298 , \16510 );
and \U$25922 ( \26299 , \26298 , RIae79c28_161);
nor \U$25923 ( \26300 , \26297 , \26299 );
nand \U$25924 ( \26301 , \26300 , \11364 );
nand \U$25925 ( \26302 , \26296 , \26301 );
xor \U$25926 ( \26303 , \26293 , \26302 );
not \U$25927 ( \26304 , \26303 );
not \U$25928 ( \26305 , \26304 );
not \U$25929 ( \26306 , \4842 );
not \U$25930 ( \26307 , \25687 );
or \U$25931 ( \26308 , \26306 , \26307 );
not \U$25932 ( \26309 , \2406 );
not \U$25933 ( \26310 , \10688 );
or \U$25934 ( \26311 , \26309 , \26310 );
not \U$25935 ( \26312 , RIae79ca0_162);
or \U$25936 ( \26313 , \3256 , \26312 );
nand \U$25937 ( \26314 , \26311 , \26313 );
nand \U$25938 ( \26315 , \26314 , \4853 );
nand \U$25939 ( \26316 , \26308 , \26315 );
not \U$25940 ( \26317 , \26316 );
not \U$25941 ( \26318 , \2272 );
not \U$25942 ( \26319 , \25707 );
or \U$25943 ( \26320 , \26318 , \26319 );
not \U$25944 ( \26321 , RIae79ac0_158);
not \U$25945 ( \26322 , \2836 );
or \U$25946 ( \26323 , \26321 , \26322 );
or \U$25947 ( \26324 , \10534 , RIae79ac0_158);
nand \U$25948 ( \26325 , \26323 , \26324 );
nand \U$25949 ( \26326 , \26325 , \10414 );
nand \U$25950 ( \26327 , \26320 , \26326 );
not \U$25951 ( \26328 , \10223 );
not \U$25952 ( \26329 , \2153 );
not \U$25953 ( \26330 , \26329 );
and \U$25954 ( \26331 , RIae79520_146, \26330 );
not \U$25955 ( \26332 , RIae79520_146);
and \U$25956 ( \26333 , \26332 , \2955 );
or \U$25957 ( \26334 , \26331 , \26333 );
not \U$25958 ( \26335 , \26334 );
or \U$25959 ( \26336 , \26328 , \26335 );
nand \U$25960 ( \26337 , \26052 , \5950 );
nand \U$25961 ( \26338 , \26336 , \26337 );
xor \U$25962 ( \26339 , \26327 , \26338 );
not \U$25963 ( \26340 , \26339 );
not \U$25964 ( \26341 , \26340 );
or \U$25965 ( \26342 , \26317 , \26341 );
not \U$25966 ( \26343 , \26316 );
nand \U$25967 ( \26344 , \26343 , \26339 );
nand \U$25968 ( \26345 , \26342 , \26344 );
not \U$25969 ( \26346 , \26345 );
not \U$25970 ( \26347 , \26346 );
or \U$25971 ( \26348 , \26305 , \26347 );
nand \U$25972 ( \26349 , \26345 , \26303 );
nand \U$25973 ( \26350 , \26348 , \26349 );
not \U$25974 ( \26351 , \2519 );
and \U$25975 ( \26352 , RIae797f0_152, \13033 );
not \U$25976 ( \26353 , RIae797f0_152);
and \U$25977 ( \26354 , \26353 , \3146 );
or \U$25978 ( \26355 , \26352 , \26354 );
not \U$25979 ( \26356 , \26355 );
or \U$25980 ( \26357 , \26351 , \26356 );
nand \U$25981 ( \26358 , \25985 , \1989 );
nand \U$25982 ( \26359 , \26357 , \26358 );
not \U$25983 ( \26360 , \11409 );
not \U$25984 ( \26361 , \25947 );
or \U$25985 ( \26362 , \26360 , \26361 );
and \U$25986 ( \26363 , RIae79ef8_167, \2510 );
not \U$25987 ( \26364 , RIae79ef8_167);
and \U$25988 ( \26365 , \26364 , \1159 );
nor \U$25989 ( \26366 , \26363 , \26365 );
not \U$25990 ( \26367 , \26366 );
nand \U$25991 ( \26368 , \26367 , \6214 );
nand \U$25992 ( \26369 , \26362 , \26368 );
xor \U$25993 ( \26370 , \26359 , \26369 );
not \U$25994 ( \26371 , \2341 );
not \U$25995 ( \26372 , \25966 );
or \U$25996 ( \26373 , \26371 , \26372 );
xor \U$25997 ( \26374 , RIae798e0_154, \3294 );
nand \U$25998 ( \26375 , \26374 , \2322 );
nand \U$25999 ( \26376 , \26373 , \26375 );
xnor \U$26000 ( \26377 , \26370 , \26376 );
xor \U$26001 ( \26378 , \26350 , \26377 );
nand \U$26002 ( \26379 , \26276 , \26378 );
or \U$26003 ( \26380 , \26274 , \26203 );
nand \U$26004 ( \26381 , \26379 , \26380 );
and \U$26005 ( \26382 , \26064 , \26045 );
and \U$26006 ( \26383 , \26054 , \26063 );
nor \U$26007 ( \26384 , \26382 , \26383 );
not \U$26008 ( \26385 , \26384 );
not \U$26009 ( \26386 , \26385 );
not \U$26010 ( \26387 , \26016 );
not \U$26011 ( \26388 , \26032 );
or \U$26012 ( \26389 , \26387 , \26388 );
not \U$26013 ( \26390 , \26018 );
nand \U$26014 ( \26391 , \26390 , \26028 );
nand \U$26015 ( \26392 , \26389 , \26391 );
or \U$26016 ( \26393 , \19466 , \9699 );
nand \U$26017 ( \26394 , \26393 , RIae7a240_174);
not \U$26018 ( \26395 , \2276 );
not \U$26019 ( \26396 , \25882 );
or \U$26020 ( \26397 , \26395 , \26396 );
nand \U$26021 ( \26398 , \23399 , \1049 );
nand \U$26022 ( \26399 , \26397 , \26398 );
xor \U$26023 ( \26400 , \26394 , \26399 );
not \U$26024 ( \26401 , \26400 );
not \U$26025 ( \26402 , \1009 );
not \U$26026 ( \26403 , \25922 );
or \U$26027 ( \26404 , \26402 , \26403 );
and \U$26028 ( \26405 , \2403 , \997 );
not \U$26029 ( \26406 , \2403 );
and \U$26030 ( \26407 , \26406 , RIae79160_138);
nor \U$26031 ( \26408 , \26405 , \26407 );
nand \U$26032 ( \26409 , \26408 , \1013 );
nand \U$26033 ( \26410 , \26404 , \26409 );
not \U$26034 ( \26411 , \26410 );
not \U$26035 ( \26412 , \26411 );
and \U$26036 ( \26413 , \26401 , \26412 );
and \U$26037 ( \26414 , \26400 , \26411 );
nor \U$26038 ( \26415 , \26413 , \26414 );
xnor \U$26039 ( \26416 , \26392 , \26415 );
not \U$26040 ( \26417 , \26416 );
or \U$26041 ( \26418 , \26386 , \26417 );
not \U$26042 ( \26419 , \26415 );
nand \U$26043 ( \26420 , \26419 , \26392 );
nand \U$26044 ( \26421 , \26418 , \26420 );
not \U$26045 ( \26422 , \26410 );
not \U$26046 ( \26423 , \26400 );
or \U$26047 ( \26424 , \26422 , \26423 );
nand \U$26048 ( \26425 , \26399 , \26394 );
nand \U$26049 ( \26426 , \26424 , \26425 );
not \U$26050 ( \26427 , \1864 );
not \U$26051 ( \26428 , \23426 );
or \U$26052 ( \26429 , \26427 , \26428 );
nand \U$26053 ( \26430 , \26123 , \1910 );
nand \U$26054 ( \26431 , \26429 , \26430 );
xor \U$26055 ( \26432 , \26431 , \23402 );
xor \U$26056 ( \26433 , \26426 , \26432 );
not \U$26057 ( \26434 , \26268 );
not \U$26058 ( \26435 , \26434 );
not \U$26059 ( \26436 , \26273 );
or \U$26060 ( \26437 , \26435 , \26436 );
not \U$26061 ( \26438 , \26232 );
nand \U$26062 ( \26439 , \26438 , \26264 );
nand \U$26063 ( \26440 , \26437 , \26439 );
xor \U$26064 ( \26441 , \26433 , \26440 );
xor \U$26065 ( \26442 , \26421 , \26441 );
xor \U$26066 ( \26443 , \26381 , \26442 );
not \U$26067 ( \26444 , \26033 );
or \U$26068 ( \26445 , \26065 , \26006 );
not \U$26069 ( \26446 , \26445 );
or \U$26070 ( \26447 , \26444 , \26446 );
nand \U$26071 ( \26448 , \26065 , \26006 );
nand \U$26072 ( \26449 , \26447 , \26448 );
not \U$26073 ( \26450 , \26449 );
not \U$26074 ( \26451 , \25940 );
nor \U$26075 ( \26452 , \26451 , \25903 );
or \U$26076 ( \26453 , \26452 , \25969 );
not \U$26077 ( \26454 , \25940 );
nand \U$26078 ( \26455 , \26454 , \25903 );
nand \U$26079 ( \26456 , \26453 , \26455 );
not \U$26080 ( \26457 , \26456 );
not \U$26081 ( \26458 , \26416 );
not \U$26082 ( \26459 , \26384 );
and \U$26083 ( \26460 , \26458 , \26459 );
and \U$26084 ( \26461 , \26416 , \26384 );
nor \U$26085 ( \26462 , \26460 , \26461 );
not \U$26086 ( \26463 , \26462 );
or \U$26087 ( \26464 , \26457 , \26463 );
or \U$26088 ( \26465 , \26462 , \26456 );
nand \U$26089 ( \26466 , \26464 , \26465 );
not \U$26090 ( \26467 , \26466 );
or \U$26091 ( \26468 , \26450 , \26467 );
not \U$26092 ( \26469 , \26462 );
nand \U$26093 ( \26470 , \26469 , \26456 );
nand \U$26094 ( \26471 , \26468 , \26470 );
xor \U$26095 ( \26472 , \26443 , \26471 );
xor \U$26096 ( \26473 , \26186 , \26472 );
xor \U$26097 ( \26474 , \25887 , \25891 );
and \U$26098 ( \26475 , \26474 , \25896 );
and \U$26099 ( \26476 , \25887 , \25891 );
or \U$26100 ( \26477 , \26475 , \26476 );
not \U$26101 ( \26478 , \25791 );
not \U$26102 ( \26479 , \25825 );
or \U$26103 ( \26480 , \26478 , \26479 );
not \U$26104 ( \26481 , \25816 );
nand \U$26105 ( \26482 , \26481 , \25821 );
nand \U$26106 ( \26483 , \26480 , \26482 );
xor \U$26107 ( \26484 , \26477 , \26483 );
xor \U$26108 ( \26485 , \25870 , \25879 );
and \U$26109 ( \26486 , \26485 , \25886 );
and \U$26110 ( \26487 , \25870 , \25879 );
or \U$26111 ( \26488 , \26486 , \26487 );
xor \U$26112 ( \26489 , \26199 , \26488 );
not \U$26113 ( \26490 , \25799 );
xnor \U$26114 ( \26491 , \25809 , \25815 );
not \U$26115 ( \26492 , \26491 );
or \U$26116 ( \26493 , \26490 , \26492 );
nand \U$26117 ( \26494 , \25815 , \25808 );
nand \U$26118 ( \26495 , \26493 , \26494 );
xor \U$26119 ( \26496 , \26489 , \26495 );
xnor \U$26120 ( \26497 , \26484 , \26496 );
not \U$26121 ( \26498 , \25786 );
not \U$26122 ( \26499 , \25826 );
or \U$26123 ( \26500 , \26498 , \26499 );
or \U$26124 ( \26501 , \25826 , \25786 );
nand \U$26125 ( \26502 , \26501 , \25831 );
nand \U$26126 ( \26503 , \26500 , \26502 );
or \U$26127 ( \26504 , \26497 , \26503 );
not \U$26128 ( \26505 , \26449 );
not \U$26129 ( \26506 , \26466 );
not \U$26130 ( \26507 , \26506 );
or \U$26131 ( \26508 , \26505 , \26507 );
not \U$26132 ( \26509 , \26449 );
nand \U$26133 ( \26510 , \26509 , \26466 );
nand \U$26134 ( \26511 , \26508 , \26510 );
nand \U$26135 ( \26512 , \26504 , \26511 );
nand \U$26136 ( \26513 , \26503 , \26497 );
nand \U$26137 ( \26514 , \26512 , \26513 );
not \U$26138 ( \26515 , \26514 );
xnor \U$26139 ( \26516 , \26473 , \26515 );
xor \U$26140 ( \26517 , \25897 , \25970 );
and \U$26141 ( \26518 , \26517 , \26066 );
and \U$26142 ( \26519 , \25897 , \25970 );
or \U$26143 ( \26520 , \26518 , \26519 );
not \U$26144 ( \26521 , \26520 );
not \U$26145 ( \26522 , \26378 );
not \U$26146 ( \26523 , \26202 );
not \U$26147 ( \26524 , \26274 );
or \U$26148 ( \26525 , \26523 , \26524 );
or \U$26149 ( \26526 , \26274 , \26202 );
nand \U$26150 ( \26527 , \26525 , \26526 );
not \U$26151 ( \26528 , \26527 );
or \U$26152 ( \26529 , \26522 , \26528 );
or \U$26153 ( \26530 , \26527 , \26378 );
nand \U$26154 ( \26531 , \26529 , \26530 );
buf \U$26155 ( \26532 , \26531 );
nand \U$26156 ( \26533 , \26521 , \26532 );
not \U$26157 ( \26534 , \25743 );
nand \U$26158 ( \26535 , \26534 , \25737 );
nand \U$26159 ( \26536 , \26533 , \26535 , \25732 );
nand \U$26160 ( \26537 , \26533 , \25744 , \25736 );
not \U$26161 ( \26538 , \26532 );
nand \U$26162 ( \26539 , \26538 , \26520 );
nand \U$26163 ( \26540 , \26536 , \26537 , \26539 );
not \U$26164 ( \26541 , \26540 );
not \U$26165 ( \26542 , \26541 );
not \U$26166 ( \26543 , \2322 );
not \U$26167 ( \26544 , \23520 );
or \U$26168 ( \26545 , \26543 , \26544 );
nand \U$26169 ( \26546 , \26374 , \14580 );
nand \U$26170 ( \26547 , \26545 , \26546 );
not \U$26171 ( \26548 , \26547 );
not \U$26172 ( \26549 , \14940 );
not \U$26173 ( \26550 , \23529 );
or \U$26174 ( \26551 , \26549 , \26550 );
nand \U$26175 ( \26552 , \26153 , \6091 );
nand \U$26176 ( \26553 , \26551 , \26552 );
xor \U$26177 ( \26554 , \26548 , \26553 );
not \U$26178 ( \26555 , \9518 );
not \U$26179 ( \26556 , \23506 );
or \U$26180 ( \26557 , \26555 , \26556 );
nand \U$26181 ( \26558 , \26144 , \10709 );
nand \U$26182 ( \26559 , \26557 , \26558 );
not \U$26183 ( \26560 , \26559 );
not \U$26184 ( \26561 , \26560 );
xor \U$26185 ( \26562 , \26554 , \26561 );
not \U$26186 ( \26563 , \26562 );
not \U$26187 ( \26564 , \26563 );
and \U$26188 ( \26565 , \23573 , \6214 );
not \U$26189 ( \26566 , \6201 );
nor \U$26190 ( \26567 , \26566 , \26366 );
nor \U$26191 ( \26568 , \26565 , \26567 );
not \U$26192 ( \26569 , \2776 );
not \U$26193 ( \26570 , \23560 );
or \U$26194 ( \26571 , \26569 , \26570 );
nand \U$26195 ( \26572 , \26300 , \2767 );
nand \U$26196 ( \26573 , \26571 , \26572 );
xnor \U$26197 ( \26574 , \26568 , \26573 );
not \U$26198 ( \26575 , \3015 );
not \U$26199 ( \26576 , \24094 );
or \U$26200 ( \26577 , \26575 , \26576 );
nand \U$26201 ( \26578 , \26325 , \2272 );
nand \U$26202 ( \26579 , \26577 , \26578 );
xor \U$26203 ( \26580 , \26574 , \26579 );
not \U$26204 ( \26581 , \26580 );
not \U$26205 ( \26582 , \26581 );
or \U$26206 ( \26583 , \26564 , \26582 );
nand \U$26207 ( \26584 , \26580 , \26562 );
nand \U$26208 ( \26585 , \26583 , \26584 );
not \U$26209 ( \26586 , \3827 );
not \U$26210 ( \26587 , \24083 );
or \U$26211 ( \26588 , \26586 , \26587 );
nand \U$26212 ( \26589 , \26280 , \1844 );
nand \U$26213 ( \26590 , \26588 , \26589 );
not \U$26214 ( \26591 , \2011 );
not \U$26215 ( \26592 , \23408 );
or \U$26216 ( \26593 , \26591 , \26592 );
nand \U$26217 ( \26594 , \26288 , \2063 );
nand \U$26218 ( \26595 , \26593 , \26594 );
xor \U$26219 ( \26596 , \26590 , \26595 );
not \U$26220 ( \26597 , \2450 );
not \U$26221 ( \26598 , \24102 );
or \U$26222 ( \26599 , \26597 , \26598 );
nand \U$26223 ( \26600 , \26209 , \2545 );
nand \U$26224 ( \26601 , \26599 , \26600 );
xor \U$26225 ( \26602 , \26596 , \26601 );
and \U$26226 ( \26603 , \26585 , \26602 );
not \U$26227 ( \26604 , \26585 );
not \U$26228 ( \26605 , \26602 );
and \U$26229 ( \26606 , \26604 , \26605 );
nor \U$26230 ( \26607 , \26603 , \26606 );
not \U$26231 ( \26608 , \26304 );
not \U$26232 ( \26609 , \26346 );
or \U$26233 ( \26610 , \26608 , \26609 );
not \U$26234 ( \26611 , \26377 );
nand \U$26235 ( \26612 , \26610 , \26611 );
nand \U$26236 ( \26613 , \26612 , \26349 );
not \U$26237 ( \26614 , \26613 );
not \U$26238 ( \26615 , \26213 );
not \U$26239 ( \26616 , \26227 );
or \U$26240 ( \26617 , \26615 , \26616 );
nand \U$26241 ( \26618 , \26219 , \26214 );
nand \U$26242 ( \26619 , \26617 , \26618 );
not \U$26243 ( \26620 , \26619 );
not \U$26244 ( \26621 , \26620 );
not \U$26245 ( \26622 , \927 );
not \U$26246 ( \26623 , \23786 );
or \U$26247 ( \26624 , \26622 , \26623 );
nand \U$26248 ( \26625 , \26240 , \951 );
nand \U$26249 ( \26626 , \26624 , \26625 );
not \U$26250 ( \26627 , \5858 );
not \U$26251 ( \26628 , \26250 );
or \U$26252 ( \26629 , \26627 , \26628 );
nand \U$26253 ( \26630 , \23778 , \1072 );
nand \U$26254 ( \26631 , \26629 , \26630 );
xor \U$26255 ( \26632 , \26626 , \26631 );
not \U$26256 ( \26633 , \26632 );
not \U$26257 ( \26634 , \5124 );
not \U$26258 ( \26635 , \23814 );
or \U$26259 ( \26636 , \26634 , \26635 );
nand \U$26260 ( \26637 , \26258 , \797 );
nand \U$26261 ( \26638 , \26636 , \26637 );
not \U$26262 ( \26639 , \26638 );
not \U$26263 ( \26640 , \26639 );
and \U$26264 ( \26641 , \26633 , \26640 );
and \U$26265 ( \26642 , \26632 , \26639 );
nor \U$26266 ( \26643 , \26641 , \26642 );
not \U$26267 ( \26644 , \26643 );
not \U$26268 ( \26645 , \26644 );
or \U$26269 ( \26646 , \26621 , \26645 );
nand \U$26270 ( \26647 , \26643 , \26619 );
nand \U$26271 ( \26648 , \26646 , \26647 );
not \U$26272 ( \26649 , \26316 );
not \U$26273 ( \26650 , \26339 );
or \U$26274 ( \26651 , \26649 , \26650 );
nand \U$26275 ( \26652 , \26338 , \26327 );
nand \U$26276 ( \26653 , \26651 , \26652 );
not \U$26277 ( \26654 , \26653 );
and \U$26278 ( \26655 , \26648 , \26654 );
not \U$26279 ( \26656 , \26648 );
and \U$26280 ( \26657 , \26656 , \26653 );
nor \U$26281 ( \26658 , \26655 , \26657 );
not \U$26282 ( \26659 , \26658 );
and \U$26283 ( \26660 , \26614 , \26659 );
and \U$26284 ( \26661 , \26613 , \26658 );
nor \U$26285 ( \26662 , \26660 , \26661 );
xnor \U$26286 ( \26663 , \26607 , \26662 );
xor \U$26287 ( \26664 , \26190 , \26194 );
and \U$26288 ( \26665 , \26664 , \26201 );
and \U$26289 ( \26666 , \26190 , \26194 );
or \U$26290 ( \26667 , \26665 , \26666 );
xor \U$26291 ( \26668 , \26115 , \26125 );
and \U$26292 ( \26669 , \26668 , \26136 );
and \U$26293 ( \26670 , \26115 , \26125 );
or \U$26294 ( \26671 , \26669 , \26670 );
not \U$26295 ( \26672 , \26359 );
not \U$26296 ( \26673 , \26376 );
or \U$26297 ( \26674 , \26672 , \26673 );
or \U$26298 ( \26675 , \26359 , \26376 );
nand \U$26299 ( \26676 , \26675 , \26369 );
nand \U$26300 ( \26677 , \26674 , \26676 );
xor \U$26301 ( \26678 , \26671 , \26677 );
xor \U$26302 ( \26679 , \26146 , \26155 );
and \U$26303 ( \26680 , \26679 , \26167 );
and \U$26304 ( \26681 , \26146 , \26155 );
or \U$26305 ( \26682 , \26680 , \26681 );
xor \U$26306 ( \26683 , \26678 , \26682 );
xor \U$26307 ( \26684 , \26667 , \26683 );
not \U$26308 ( \26685 , \26242 );
not \U$26309 ( \26686 , \26263 );
or \U$26310 ( \26687 , \26685 , \26686 );
nand \U$26311 ( \26688 , \26262 , \26252 );
nand \U$26312 ( \26689 , \26687 , \26688 );
and \U$26313 ( \26690 , RIae78b48_125, \12614 );
not \U$26314 ( \26691 , \868 );
not \U$26315 ( \26692 , \23766 );
or \U$26316 ( \26693 , \26691 , \26692 );
nand \U$26317 ( \26694 , \26217 , \1129 );
nand \U$26318 ( \26695 , \26693 , \26694 );
xor \U$26319 ( \26696 , \26690 , \26695 );
not \U$26320 ( \26697 , \9792 );
not \U$26321 ( \26698 , \26134 );
or \U$26322 ( \26699 , \26697 , \26698 );
nand \U$26323 ( \26700 , \9814 , RIae7a2b8_175);
nand \U$26324 ( \26701 , \26699 , \26700 );
xor \U$26325 ( \26702 , \26696 , \26701 );
xor \U$26326 ( \26703 , \26689 , \26702 );
not \U$26327 ( \26704 , \1843 );
not \U$26328 ( \26705 , \25937 );
or \U$26329 ( \26706 , \26704 , \26705 );
nand \U$26330 ( \26707 , \26706 , \26281 );
and \U$26331 ( \26708 , \26707 , \26292 );
nor \U$26332 ( \26709 , \26708 , \26302 );
nor \U$26333 ( \26710 , \26707 , \26292 );
nor \U$26334 ( \26711 , \26709 , \26710 );
xor \U$26335 ( \26712 , \26703 , \26711 );
xor \U$26336 ( \26713 , \26684 , \26712 );
and \U$26337 ( \26714 , \26663 , \26713 );
not \U$26338 ( \26715 , \26663 );
not \U$26339 ( \26716 , \26713 );
and \U$26340 ( \26717 , \26715 , \26716 );
nor \U$26341 ( \26718 , \26714 , \26717 );
not \U$26342 ( \26719 , \26718 );
not \U$26343 ( \26720 , \26719 );
and \U$26344 ( \26721 , \26137 , \26168 );
or \U$26345 ( \26722 , \26177 , \26721 );
or \U$26346 ( \26723 , \26168 , \26137 );
nand \U$26347 ( \26724 , \26722 , \26723 );
not \U$26348 ( \26725 , \26724 );
not \U$26349 ( \26726 , \2924 );
not \U$26350 ( \26727 , \23581 );
or \U$26351 ( \26728 , \26726 , \26727 );
nand \U$26352 ( \26729 , \26334 , \2189 );
nand \U$26353 ( \26730 , \26728 , \26729 );
not \U$26354 ( \26731 , \10451 );
not \U$26355 ( \26732 , \23494 );
or \U$26356 ( \26733 , \26731 , \26732 );
nand \U$26357 ( \26734 , \26408 , \1008 );
nand \U$26358 ( \26735 , \26733 , \26734 );
not \U$26359 ( \26736 , \1989 );
not \U$26360 ( \26737 , \26355 );
or \U$26361 ( \26738 , \26736 , \26737 );
nand \U$26362 ( \26739 , \23462 , \2519 );
nand \U$26363 ( \26740 , \26738 , \26739 );
xor \U$26364 ( \26741 , \26735 , \26740 );
not \U$26365 ( \26742 , \1501 );
not \U$26366 ( \26743 , \23470 );
or \U$26367 ( \26744 , \26742 , \26743 );
nand \U$26368 ( \26745 , \26111 , \2650 );
nand \U$26369 ( \26746 , \26744 , \26745 );
xor \U$26370 ( \26747 , \26741 , \26746 );
xor \U$26371 ( \26748 , \26730 , \26747 );
not \U$26372 ( \26749 , \4853 );
not \U$26373 ( \26750 , \23538 );
or \U$26374 ( \26751 , \26749 , \26750 );
nand \U$26375 ( \26752 , \26314 , \11761 );
nand \U$26376 ( \26753 , \26751 , \26752 );
not \U$26377 ( \26754 , \5285 );
not \U$26378 ( \26755 , \23550 );
or \U$26379 ( \26756 , \26754 , \26755 );
nand \U$26380 ( \26757 , \26165 , \2458 );
nand \U$26381 ( \26758 , \26756 , \26757 );
xor \U$26382 ( \26759 , \26753 , \26758 );
xnor \U$26383 ( \26760 , \26748 , \26759 );
not \U$26384 ( \26761 , \26760 );
not \U$26385 ( \26762 , \26761 );
not \U$26386 ( \26763 , \26488 );
not \U$26387 ( \26764 , \26199 );
not \U$26388 ( \26765 , \26495 );
or \U$26389 ( \26766 , \26764 , \26765 );
or \U$26390 ( \26767 , \26495 , \26199 );
nand \U$26391 ( \26768 , \26766 , \26767 );
not \U$26392 ( \26769 , \26768 );
or \U$26393 ( \26770 , \26763 , \26769 );
not \U$26394 ( \26771 , \26199 );
nand \U$26395 ( \26772 , \26771 , \26495 );
nand \U$26396 ( \26773 , \26770 , \26772 );
not \U$26397 ( \26774 , \26773 );
not \U$26398 ( \26775 , \26774 );
or \U$26399 ( \26776 , \26762 , \26775 );
nand \U$26400 ( \26777 , \26773 , \26760 );
nand \U$26401 ( \26778 , \26776 , \26777 );
xor \U$26402 ( \26779 , \26725 , \26778 );
not \U$26403 ( \26780 , \26483 );
xnor \U$26404 ( \26781 , \26477 , \26496 );
not \U$26405 ( \26782 , \26781 );
or \U$26406 ( \26783 , \26780 , \26782 );
not \U$26407 ( \26784 , \26496 );
nand \U$26408 ( \26785 , \26784 , \26477 );
nand \U$26409 ( \26786 , \26783 , \26785 );
xnor \U$26410 ( \26787 , \26779 , \26786 );
not \U$26411 ( \26788 , \26787 );
or \U$26412 ( \26789 , \26720 , \26788 );
not \U$26413 ( \26790 , \26787 );
nand \U$26414 ( \26791 , \26790 , \26718 );
nand \U$26415 ( \26792 , \26789 , \26791 );
not \U$26416 ( \26793 , \26792 );
not \U$26417 ( \26794 , \26793 );
or \U$26418 ( \26795 , \26542 , \26794 );
nand \U$26419 ( \26796 , \26792 , \26540 );
nand \U$26420 ( \26797 , \26795 , \26796 );
not \U$26421 ( \26798 , \26797 );
not \U$26422 ( \26799 , \25832 );
not \U$26423 ( \26800 , \25781 );
not \U$26424 ( \26801 , \26800 );
or \U$26425 ( \26802 , \26799 , \26801 );
nand \U$26426 ( \26803 , \26802 , \25756 );
not \U$26427 ( \26804 , \26183 );
xor \U$26428 ( \26805 , \26106 , \26804 );
nand \U$26429 ( \26806 , \25781 , \25833 );
and \U$26430 ( \26807 , \26803 , \26805 , \26806 );
xor \U$26431 ( \26808 , \26497 , \26503 );
not \U$26432 ( \26809 , \26511 );
and \U$26433 ( \26810 , \26808 , \26809 );
not \U$26434 ( \26811 , \26808 );
not \U$26435 ( \26812 , \26809 );
and \U$26436 ( \26813 , \26811 , \26812 );
nor \U$26437 ( \26814 , \26810 , \26813 );
or \U$26438 ( \26815 , \26807 , \26814 );
xor \U$26439 ( \26816 , \26106 , \26183 );
nand \U$26440 ( \26817 , \26803 , \26806 );
nand \U$26441 ( \26818 , \26816 , \26817 );
nand \U$26442 ( \26819 , \26815 , \26818 );
not \U$26443 ( \26820 , \26819 );
not \U$26444 ( \26821 , \26820 );
and \U$26445 ( \26822 , \26798 , \26821 );
and \U$26446 ( \26823 , \26797 , \26820 );
nor \U$26447 ( \26824 , \26822 , \26823 );
xor \U$26448 ( \26825 , \26516 , \26824 );
not \U$26449 ( \26826 , \26067 );
nand \U$26450 ( \26827 , \26826 , \26075 );
not \U$26451 ( \26828 , \26827 );
not \U$26452 ( \26829 , \25861 );
or \U$26453 ( \26830 , \26828 , \26829 );
not \U$26454 ( \26831 , \26075 );
nand \U$26455 ( \26832 , \26831 , \26067 );
nand \U$26456 ( \26833 , \26830 , \26832 );
not \U$26457 ( \26834 , \26833 );
not \U$26458 ( \26835 , \26531 );
not \U$26459 ( \26836 , \26520 );
and \U$26460 ( \26837 , \26835 , \26836 );
and \U$26461 ( \26838 , \26520 , \26531 );
nor \U$26462 ( \26839 , \26837 , \26838 );
not \U$26463 ( \26840 , \26839 );
not \U$26464 ( \26841 , \25736 );
not \U$26465 ( \26842 , \25743 );
or \U$26466 ( \26843 , \26841 , \26842 );
not \U$26467 ( \26844 , \25732 );
nand \U$26468 ( \26845 , \26843 , \26844 );
nand \U$26469 ( \26846 , \26535 , \26845 );
not \U$26470 ( \26847 , \26846 );
and \U$26471 ( \26848 , \26840 , \26847 );
and \U$26472 ( \26849 , \26846 , \26839 );
nor \U$26473 ( \26850 , \26848 , \26849 );
not \U$26474 ( \26851 , \26850 );
nand \U$26475 ( \26852 , \26834 , \26851 );
not \U$26476 ( \26853 , \26852 );
nor \U$26477 ( \26854 , \25751 , \25745 );
or \U$26478 ( \26855 , \25834 , \26854 );
nand \U$26479 ( \26856 , \25751 , \25745 );
nand \U$26480 ( \26857 , \26855 , \26856 );
not \U$26481 ( \26858 , \26857 );
or \U$26482 ( \26859 , \26853 , \26858 );
not \U$26483 ( \26860 , \26851 );
nand \U$26484 ( \26861 , \26860 , \26833 );
nand \U$26485 ( \26862 , \26859 , \26861 );
not \U$26486 ( \26863 , \26862 );
xor \U$26487 ( \26864 , \26825 , \26863 );
not \U$26488 ( \26865 , \26864 );
xnor \U$26489 ( \26866 , \26833 , \26850 );
xnor \U$26490 ( \26867 , \26866 , \26857 );
not \U$26491 ( \26868 , \26867 );
not \U$26492 ( \26869 , \26807 );
nand \U$26493 ( \26870 , \26869 , \26818 );
not \U$26494 ( \26871 , \26814 );
and \U$26495 ( \26872 , \26870 , \26871 );
not \U$26496 ( \26873 , \26870 );
and \U$26497 ( \26874 , \26873 , \26814 );
nor \U$26498 ( \26875 , \26872 , \26874 );
not \U$26499 ( \26876 , \26875 );
and \U$26500 ( \26877 , \26868 , \26876 );
and \U$26501 ( \26878 , \26867 , \26875 );
nor \U$26502 ( \26879 , \26877 , \26878 );
not \U$26503 ( \26880 , \26879 );
not \U$26504 ( \26881 , \25847 );
not \U$26505 ( \26882 , \26084 );
not \U$26506 ( \26883 , \26882 );
or \U$26507 ( \26884 , \26881 , \26883 );
not \U$26508 ( \26885 , \26080 );
nand \U$26509 ( \26886 , \26885 , \25852 );
nand \U$26510 ( \26887 , \26884 , \26886 );
not \U$26511 ( \26888 , \26887 );
not \U$26512 ( \26889 , \26888 );
and \U$26513 ( \26890 , \26880 , \26889 );
not \U$26514 ( \26891 , \26867 );
nor \U$26515 ( \26892 , \26891 , \26875 );
nor \U$26516 ( \26893 , \26890 , \26892 );
not \U$26517 ( \26894 , \26893 );
or \U$26518 ( \26895 , \26865 , \26894 );
not \U$26519 ( \26896 , \26879 );
not \U$26520 ( \26897 , \26887 );
and \U$26521 ( \26898 , \26896 , \26897 );
and \U$26522 ( \26899 , \26879 , \26887 );
nor \U$26523 ( \26900 , \26898 , \26899 );
xor \U$26524 ( \26901 , \25835 , \25839 );
and \U$26525 ( \26902 , \26901 , \26085 );
and \U$26526 ( \26903 , \25835 , \25839 );
or \U$26527 ( \26904 , \26902 , \26903 );
nand \U$26528 ( \26905 , \26900 , \26904 );
nand \U$26529 ( \26906 , \26895 , \26905 );
not \U$26530 ( \26907 , \26906 );
not \U$26531 ( \26908 , \26820 );
nand \U$26532 ( \26909 , \26793 , \26540 );
not \U$26533 ( \26910 , \26909 );
or \U$26534 ( \26911 , \26908 , \26910 );
not \U$26535 ( \26912 , \26540 );
nand \U$26536 ( \26913 , \26912 , \26792 );
nand \U$26537 ( \26914 , \26911 , \26913 );
not \U$26538 ( \26915 , \26914 );
not \U$26539 ( \26916 , \26725 );
not \U$26540 ( \26917 , \26778 );
nand \U$26541 ( \26918 , \26916 , \26917 );
not \U$26542 ( \26919 , \26918 );
not \U$26543 ( \26920 , \26786 );
or \U$26544 ( \26921 , \26919 , \26920 );
not \U$26545 ( \26922 , \26917 );
nand \U$26546 ( \26923 , \26922 , \26725 );
nand \U$26547 ( \26924 , \26921 , \26923 );
xor \U$26548 ( \26925 , \26667 , \26683 );
and \U$26549 ( \26926 , \26925 , \26712 );
and \U$26550 ( \26927 , \26667 , \26683 );
or \U$26551 ( \26928 , \26926 , \26927 );
not \U$26552 ( \26929 , \26432 );
not \U$26553 ( \26930 , \26426 );
or \U$26554 ( \26931 , \26929 , \26930 );
nand \U$26555 ( \26932 , \23402 , \26431 );
nand \U$26556 ( \26933 , \26931 , \26932 );
not \U$26557 ( \26934 , \26653 );
not \U$26558 ( \26935 , \26648 );
or \U$26559 ( \26936 , \26934 , \26935 );
nand \U$26560 ( \26937 , \26644 , \26619 );
nand \U$26561 ( \26938 , \26936 , \26937 );
xor \U$26562 ( \26939 , \26933 , \26938 );
xor \U$26563 ( \26940 , \26689 , \26702 );
and \U$26564 ( \26941 , \26940 , \26711 );
and \U$26565 ( \26942 , \26689 , \26702 );
or \U$26566 ( \26943 , \26941 , \26942 );
and \U$26567 ( \26944 , \26939 , \26943 );
not \U$26568 ( \26945 , \26939 );
not \U$26569 ( \26946 , \26943 );
and \U$26570 ( \26947 , \26945 , \26946 );
nor \U$26571 ( \26948 , \26944 , \26947 );
xor \U$26572 ( \26949 , \26928 , \26948 );
xor \U$26573 ( \26950 , \26671 , \26677 );
and \U$26574 ( \26951 , \26950 , \26682 );
and \U$26575 ( \26952 , \26671 , \26677 );
or \U$26576 ( \26953 , \26951 , \26952 );
not \U$26577 ( \26954 , \26638 );
not \U$26578 ( \26955 , \26632 );
or \U$26579 ( \26956 , \26954 , \26955 );
nand \U$26580 ( \26957 , \26631 , \26626 );
nand \U$26581 ( \26958 , \26956 , \26957 );
xor \U$26582 ( \26959 , \26690 , \26695 );
and \U$26583 ( \26960 , \26959 , \26701 );
and \U$26584 ( \26961 , \26690 , \26695 );
or \U$26585 ( \26962 , \26960 , \26961 );
xor \U$26586 ( \26963 , \26958 , \26962 );
not \U$26587 ( \26964 , \23793 );
xor \U$26588 ( \26965 , \23768 , \26964 );
xor \U$26589 ( \26966 , \26963 , \26965 );
xor \U$26590 ( \26967 , \26953 , \26966 );
not \U$26591 ( \26968 , \26602 );
not \U$26592 ( \26969 , \26585 );
or \U$26593 ( \26970 , \26968 , \26969 );
nand \U$26594 ( \26971 , \26580 , \26563 );
nand \U$26595 ( \26972 , \26970 , \26971 );
xor \U$26596 ( \26973 , \26967 , \26972 );
xor \U$26597 ( \26974 , \26949 , \26973 );
xor \U$26598 ( \26975 , \26924 , \26974 );
xor \U$26599 ( \26976 , \26381 , \26442 );
and \U$26600 ( \26977 , \26976 , \26471 );
and \U$26601 ( \26978 , \26381 , \26442 );
or \U$26602 ( \26979 , \26977 , \26978 );
xor \U$26603 ( \26980 , \26975 , \26979 );
not \U$26604 ( \26981 , \26980 );
not \U$26605 ( \26982 , \26716 );
not \U$26606 ( \26983 , \26787 );
or \U$26607 ( \26984 , \26982 , \26983 );
nand \U$26608 ( \26985 , \26984 , \26663 );
nand \U$26609 ( \26986 , \26790 , \26713 );
nand \U$26610 ( \26987 , \26985 , \26986 );
not \U$26611 ( \26988 , \26987 );
not \U$26612 ( \26989 , \26662 );
and \U$26613 ( \26990 , \26989 , \26607 );
and \U$26614 ( \26991 , \26612 , \26349 );
nor \U$26615 ( \26992 , \26991 , \26658 );
nor \U$26616 ( \26993 , \26990 , \26992 );
not \U$26617 ( \26994 , \26590 );
xor \U$26618 ( \26995 , \26601 , \26595 );
not \U$26619 ( \26996 , \26995 );
or \U$26620 ( \26997 , \26994 , \26996 );
nand \U$26621 ( \26998 , \26601 , \26595 );
nand \U$26622 ( \26999 , \26997 , \26998 );
not \U$26623 ( \27000 , \26999 );
not \U$26624 ( \27001 , \27000 );
xor \U$26625 ( \27002 , \26735 , \26740 );
and \U$26626 ( \27003 , \27002 , \26746 );
and \U$26627 ( \27004 , \26735 , \26740 );
nor \U$26628 ( \27005 , \27003 , \27004 );
not \U$26629 ( \27006 , \27005 );
xor \U$26630 ( \27007 , \23823 , \23804 );
not \U$26631 ( \27008 , \27007 );
or \U$26632 ( \27009 , \27006 , \27008 );
or \U$26633 ( \27010 , \27007 , \27005 );
nand \U$26634 ( \27011 , \27009 , \27010 );
not \U$26635 ( \27012 , \27011 );
and \U$26636 ( \27013 , \27001 , \27012 );
and \U$26637 ( \27014 , \27011 , \27000 );
nor \U$26638 ( \27015 , \27013 , \27014 );
not \U$26639 ( \27016 , \27015 );
not \U$26640 ( \27017 , \26548 );
not \U$26641 ( \27018 , \26560 );
or \U$26642 ( \27019 , \27017 , \27018 );
not \U$26643 ( \27020 , \26547 );
not \U$26644 ( \27021 , \26559 );
or \U$26645 ( \27022 , \27020 , \27021 );
not \U$26646 ( \27023 , \26553 );
nand \U$26647 ( \27024 , \27022 , \27023 );
nand \U$26648 ( \27025 , \27019 , \27024 );
not \U$26649 ( \27026 , \27025 );
not \U$26650 ( \27027 , \26579 );
not \U$26651 ( \27028 , \26574 );
or \U$26652 ( \27029 , \27027 , \27028 );
not \U$26653 ( \27030 , \26568 );
nand \U$26654 ( \27031 , \27030 , \26573 );
nand \U$26655 ( \27032 , \27029 , \27031 );
xor \U$26656 ( \27033 , \27026 , \27032 );
not \U$26657 ( \27034 , \26730 );
not \U$26658 ( \27035 , \26759 );
or \U$26659 ( \27036 , \27034 , \27035 );
nand \U$26660 ( \27037 , \26758 , \26753 );
nand \U$26661 ( \27038 , \27036 , \27037 );
not \U$26662 ( \27039 , \27038 );
xnor \U$26663 ( \27040 , \27033 , \27039 );
not \U$26664 ( \27041 , \27040 );
or \U$26665 ( \27042 , \27016 , \27041 );
or \U$26666 ( \27043 , \27040 , \27015 );
nand \U$26667 ( \27044 , \27042 , \27043 );
not \U$26668 ( \27045 , \27044 );
not \U$26669 ( \27046 , \26761 );
not \U$26670 ( \27047 , \26773 );
or \U$26671 ( \27048 , \27046 , \27047 );
not \U$26672 ( \27049 , \26730 );
nand \U$26673 ( \27050 , \27049 , \26759 );
not \U$26674 ( \27051 , \27050 );
not \U$26675 ( \27052 , \26759 );
nand \U$26676 ( \27053 , \27052 , \26730 );
not \U$26677 ( \27054 , \27053 );
or \U$26678 ( \27055 , \27051 , \27054 );
nand \U$26679 ( \27056 , \27055 , \26747 );
nand \U$26680 ( \27057 , \27048 , \27056 );
not \U$26681 ( \27058 , \27057 );
not \U$26682 ( \27059 , \27058 );
and \U$26683 ( \27060 , \27045 , \27059 );
and \U$26684 ( \27061 , \27058 , \27044 );
nor \U$26685 ( \27062 , \27060 , \27061 );
xor \U$26686 ( \27063 , \26993 , \27062 );
and \U$26687 ( \27064 , \26441 , \26421 );
and \U$26688 ( \27065 , \26433 , \26440 );
nor \U$26689 ( \27066 , \27064 , \27065 );
not \U$26690 ( \27067 , \23435 );
not \U$26691 ( \27068 , \23419 );
or \U$26692 ( \27069 , \27067 , \27068 );
or \U$26693 ( \27070 , \23435 , \23419 );
nand \U$26694 ( \27071 , \27069 , \27070 );
not \U$26695 ( \27072 , \27071 );
xor \U$26696 ( \27073 , \23450 , \23478 );
xnor \U$26697 ( \27074 , \27073 , \23464 );
not \U$26698 ( \27075 , \27074 );
and \U$26699 ( \27076 , \27072 , \27075 );
and \U$26700 ( \27077 , \27074 , \27071 );
nor \U$26701 ( \27078 , \27076 , \27077 );
xor \U$26702 ( \27079 , \23533 , \23542 );
xor \U$26703 ( \27080 , \27079 , \23554 );
xor \U$26704 ( \27081 , \27078 , \27080 );
not \U$26705 ( \27082 , \27081 );
not \U$26706 ( \27083 , \23509 );
not \U$26707 ( \27084 , \23496 );
not \U$26708 ( \27085 , \23522 );
or \U$26709 ( \27086 , \27084 , \27085 );
or \U$26710 ( \27087 , \23522 , \23496 );
nand \U$26711 ( \27088 , \27086 , \27087 );
not \U$26712 ( \27089 , \27088 );
or \U$26713 ( \27090 , \27083 , \27089 );
or \U$26714 ( \27091 , \27088 , \23509 );
nand \U$26715 ( \27092 , \27090 , \27091 );
xor \U$26716 ( \27093 , \23593 , \23564 );
xor \U$26717 ( \27094 , \27092 , \27093 );
xor \U$26718 ( \27095 , \24087 , \24096 );
xor \U$26719 ( \27096 , \27095 , \24106 );
xor \U$26720 ( \27097 , \27094 , \27096 );
not \U$26721 ( \27098 , \27097 );
or \U$26722 ( \27099 , \27082 , \27098 );
or \U$26723 ( \27100 , \27097 , \27081 );
nand \U$26724 ( \27101 , \27099 , \27100 );
xor \U$26725 ( \27102 , \27066 , \27101 );
xor \U$26726 ( \27103 , \27063 , \27102 );
not \U$26727 ( \27104 , \27103 );
and \U$26728 ( \27105 , \26988 , \27104 );
and \U$26729 ( \27106 , \26987 , \27103 );
nor \U$26730 ( \27107 , \27105 , \27106 );
not \U$26731 ( \27108 , \26186 );
not \U$26732 ( \27109 , \26515 );
or \U$26733 ( \27110 , \27108 , \27109 );
nand \U$26734 ( \27111 , \27110 , \26472 );
not \U$26735 ( \27112 , \26186 );
nand \U$26736 ( \27113 , \27112 , \26514 );
nand \U$26737 ( \27114 , \27111 , \27113 );
and \U$26738 ( \27115 , \27107 , \27114 );
not \U$26739 ( \27116 , \27107 );
not \U$26740 ( \27117 , \27114 );
and \U$26741 ( \27118 , \27116 , \27117 );
nor \U$26742 ( \27119 , \27115 , \27118 );
not \U$26743 ( \27120 , \27119 );
or \U$26744 ( \27121 , \26981 , \27120 );
or \U$26745 ( \27122 , \27119 , \26980 );
nand \U$26746 ( \27123 , \27121 , \27122 );
not \U$26747 ( \27124 , \27123 );
or \U$26748 ( \27125 , \26915 , \27124 );
not \U$26749 ( \27126 , \27119 );
or \U$26750 ( \27127 , \27126 , \26980 );
nand \U$26751 ( \27128 , \27125 , \27127 );
not \U$26752 ( \27129 , \27040 );
not \U$26753 ( \27130 , \27057 );
or \U$26754 ( \27131 , \27129 , \27130 );
nand \U$26755 ( \27132 , \27131 , \27015 );
not \U$26756 ( \27133 , \27040 );
nand \U$26757 ( \27134 , \27133 , \27058 );
and \U$26758 ( \27135 , \27132 , \27134 );
xor \U$26759 ( \27136 , \23446 , \23448 );
xor \U$26760 ( \27137 , \27136 , \23481 );
xor \U$26761 ( \27138 , \27092 , \27093 );
and \U$26762 ( \27139 , \27138 , \27096 );
and \U$26763 ( \27140 , \27092 , \27093 );
or \U$26764 ( \27141 , \27139 , \27140 );
not \U$26765 ( \27142 , \27141 );
xor \U$26766 ( \27143 , \27137 , \27142 );
not \U$26767 ( \27144 , \27071 );
not \U$26768 ( \27145 , \27144 );
not \U$26769 ( \27146 , \27074 );
and \U$26770 ( \27147 , \27145 , \27146 );
not \U$26771 ( \27148 , \27078 );
and \U$26772 ( \27149 , \27148 , \27080 );
nor \U$26773 ( \27150 , \27147 , \27149 );
xor \U$26774 ( \27151 , \27143 , \27150 );
not \U$26775 ( \27152 , \27151 );
nand \U$26776 ( \27153 , \27135 , \27152 );
not \U$26777 ( \27154 , \27134 );
not \U$26778 ( \27155 , \27132 );
or \U$26779 ( \27156 , \27154 , \27155 );
nand \U$26780 ( \27157 , \27156 , \27151 );
nand \U$26781 ( \27158 , \27153 , \27157 );
not \U$26782 ( \27159 , \27066 );
not \U$26783 ( \27160 , \27159 );
not \U$26784 ( \27161 , \27101 );
or \U$26785 ( \27162 , \27160 , \27161 );
not \U$26786 ( \27163 , \27081 );
nand \U$26787 ( \27164 , \27163 , \27097 );
nand \U$26788 ( \27165 , \27162 , \27164 );
and \U$26789 ( \27166 , \27158 , \27165 );
not \U$26790 ( \27167 , \27158 );
not \U$26791 ( \27168 , \27165 );
and \U$26792 ( \27169 , \27167 , \27168 );
nor \U$26793 ( \27170 , \27166 , \27169 );
not \U$26794 ( \27171 , \27170 );
not \U$26795 ( \27172 , \27171 );
xor \U$26796 ( \27173 , \26993 , \27062 );
and \U$26797 ( \27174 , \27173 , \27102 );
and \U$26798 ( \27175 , \26993 , \27062 );
or \U$26799 ( \27176 , \27174 , \27175 );
not \U$26800 ( \27177 , \27176 );
or \U$26801 ( \27178 , \27172 , \27177 );
not \U$26802 ( \27179 , \27176 );
nand \U$26803 ( \27180 , \27179 , \27170 );
nand \U$26804 ( \27181 , \27178 , \27180 );
xor \U$26805 ( \27182 , \26924 , \26974 );
and \U$26806 ( \27183 , \27182 , \26979 );
and \U$26807 ( \27184 , \26924 , \26974 );
or \U$26808 ( \27185 , \27183 , \27184 );
xor \U$26809 ( \27186 , \27181 , \27185 );
not \U$26810 ( \27187 , \27186 );
xor \U$26811 ( \27188 , \26928 , \26948 );
and \U$26812 ( \27189 , \27188 , \26973 );
and \U$26813 ( \27190 , \26928 , \26948 );
or \U$26814 ( \27191 , \27189 , \27190 );
xor \U$26815 ( \27192 , \23383 , \23384 );
xor \U$26816 ( \27193 , \27192 , \23437 );
not \U$26817 ( \27194 , \24077 );
and \U$26818 ( \27195 , \24118 , \27194 );
not \U$26819 ( \27196 , \24118 );
and \U$26820 ( \27197 , \27196 , \24077 );
nor \U$26821 ( \27198 , \27195 , \27197 );
xor \U$26822 ( \27199 , \27193 , \27198 );
or \U$26823 ( \27200 , \26933 , \26938 );
and \U$26824 ( \27201 , \27200 , \26943 );
and \U$26825 ( \27202 , \26933 , \26938 );
nor \U$26826 ( \27203 , \27201 , \27202 );
xor \U$26827 ( \27204 , \27199 , \27203 );
not \U$26828 ( \27205 , \27204 );
and \U$26829 ( \27206 , \27191 , \27205 );
not \U$26830 ( \27207 , \27191 );
and \U$26831 ( \27208 , \27207 , \27204 );
nor \U$26832 ( \27209 , \27206 , \27208 );
and \U$26833 ( \27210 , \23879 , \23872 );
not \U$26834 ( \27211 , \23879 );
and \U$26835 ( \27212 , \27211 , \23887 );
nor \U$26836 ( \27213 , \27210 , \27212 );
xnor \U$26837 ( \27214 , \23886 , \27213 );
not \U$26838 ( \27215 , \26999 );
not \U$26839 ( \27216 , \27011 );
or \U$26840 ( \27217 , \27215 , \27216 );
not \U$26841 ( \27218 , \27005 );
nand \U$26842 ( \27219 , \27218 , \27007 );
nand \U$26843 ( \27220 , \27217 , \27219 );
not \U$26844 ( \27221 , \27220 );
xor \U$26845 ( \27222 , \27214 , \27221 );
xor \U$26846 ( \27223 , \23095 , \23797 );
xnor \U$26847 ( \27224 , \27223 , \23828 );
xor \U$26848 ( \27225 , \27222 , \27224 );
xor \U$26849 ( \27226 , \26953 , \26966 );
and \U$26850 ( \27227 , \27226 , \26972 );
and \U$26851 ( \27228 , \26953 , \26966 );
or \U$26852 ( \27229 , \27227 , \27228 );
not \U$26853 ( \27230 , \27229 );
and \U$26854 ( \27231 , \27225 , \27230 );
not \U$26855 ( \27232 , \27225 );
and \U$26856 ( \27233 , \27232 , \27229 );
nor \U$26857 ( \27234 , \27231 , \27233 );
and \U$26858 ( \27235 , \26963 , \26965 );
and \U$26859 ( \27236 , \26958 , \26962 );
nor \U$26860 ( \27237 , \27235 , \27236 );
not \U$26861 ( \27238 , \27026 );
not \U$26862 ( \27239 , \27032 );
or \U$26863 ( \27240 , \27238 , \27239 );
nand \U$26864 ( \27241 , \27240 , \27039 );
not \U$26865 ( \27242 , \27032 );
nand \U$26866 ( \27243 , \27242 , \27025 );
nand \U$26867 ( \27244 , \27241 , \27243 );
xor \U$26868 ( \27245 , \27237 , \27244 );
xor \U$26869 ( \27246 , \23524 , \23557 );
xor \U$26870 ( \27247 , \27246 , \23598 );
xnor \U$26871 ( \27248 , \27245 , \27247 );
not \U$26872 ( \27249 , \27248 );
not \U$26873 ( \27250 , \27249 );
and \U$26874 ( \27251 , \27234 , \27250 );
not \U$26875 ( \27252 , \27234 );
and \U$26876 ( \27253 , \27252 , \27249 );
nor \U$26877 ( \27254 , \27251 , \27253 );
and \U$26878 ( \27255 , \27209 , \27254 );
not \U$26879 ( \27256 , \27209 );
not \U$26880 ( \27257 , \27254 );
and \U$26881 ( \27258 , \27256 , \27257 );
or \U$26882 ( \27259 , \27255 , \27258 );
not \U$26883 ( \27260 , \27259 );
not \U$26884 ( \27261 , \27113 );
not \U$26885 ( \27262 , \27111 );
or \U$26886 ( \27263 , \27261 , \27262 );
nand \U$26887 ( \27264 , \26985 , \27103 , \26986 );
nand \U$26888 ( \27265 , \27263 , \27264 );
not \U$26889 ( \27266 , \27103 );
nand \U$26890 ( \27267 , \27266 , \26987 );
nand \U$26891 ( \27268 , \27265 , \27267 );
not \U$26892 ( \27269 , \27268 );
or \U$26893 ( \27270 , \27260 , \27269 );
or \U$26894 ( \27271 , \27268 , \27259 );
nand \U$26895 ( \27272 , \27270 , \27271 );
not \U$26896 ( \27273 , \27272 );
or \U$26897 ( \27274 , \27187 , \27273 );
or \U$26898 ( \27275 , \27186 , \27272 );
nand \U$26899 ( \27276 , \27274 , \27275 );
nand \U$26900 ( \27277 , \27128 , \27276 );
xor \U$26901 ( \27278 , \26516 , \26824 );
and \U$26902 ( \27279 , \27278 , \26863 );
and \U$26903 ( \27280 , \26516 , \26824 );
or \U$26904 ( \27281 , \27279 , \27280 );
not \U$26905 ( \27282 , \26914 );
xor \U$26906 ( \27283 , \26980 , \27282 );
xnor \U$26907 ( \27284 , \27283 , \27126 );
nand \U$26908 ( \27285 , \27281 , \27284 );
nand \U$26909 ( \27286 , \27277 , \27285 );
not \U$26910 ( \27287 , \27286 );
and \U$26911 ( \27288 , \26101 , \26907 , \27287 );
not \U$26912 ( \27289 , \27230 );
not \U$26913 ( \27290 , \27249 );
or \U$26914 ( \27291 , \27289 , \27290 );
not \U$26915 ( \27292 , \27229 );
not \U$26916 ( \27293 , \27248 );
or \U$26917 ( \27294 , \27292 , \27293 );
nand \U$26918 ( \27295 , \27294 , \27225 );
nand \U$26919 ( \27296 , \27291 , \27295 );
xor \U$26920 ( \27297 , \27193 , \27198 );
and \U$26921 ( \27298 , \27297 , \27203 );
and \U$26922 ( \27299 , \27193 , \27198 );
or \U$26923 ( \27300 , \27298 , \27299 );
not \U$26924 ( \27301 , \27300 );
and \U$26925 ( \27302 , \27296 , \27301 );
not \U$26926 ( \27303 , \27296 );
and \U$26927 ( \27304 , \27303 , \27300 );
nor \U$26928 ( \27305 , \27302 , \27304 );
not \U$26929 ( \27306 , \27305 );
not \U$26930 ( \27307 , \27306 );
xor \U$26931 ( \27308 , \23748 , \23756 );
xor \U$26932 ( \27309 , \27308 , \23836 );
not \U$26933 ( \27310 , \27247 );
buf \U$26934 ( \27311 , \27237 );
or \U$26935 ( \27312 , \27244 , \27311 );
not \U$26936 ( \27313 , \27312 );
or \U$26937 ( \27314 , \27310 , \27313 );
nand \U$26938 ( \27315 , \27244 , \27311 );
nand \U$26939 ( \27316 , \27314 , \27315 );
xor \U$26940 ( \27317 , \27309 , \27316 );
xor \U$26941 ( \27318 , \23484 , \23440 );
xnor \U$26942 ( \27319 , \27318 , \23608 );
xnor \U$26943 ( \27320 , \27317 , \27319 );
not \U$26944 ( \27321 , \27320 );
or \U$26945 ( \27322 , \27307 , \27321 );
not \U$26946 ( \27323 , \27301 );
nand \U$26947 ( \27324 , \27323 , \27296 );
nand \U$26948 ( \27325 , \27322 , \27324 );
xor \U$26949 ( \27326 , \23160 , \23190 );
xor \U$26950 ( \27327 , \27326 , \23159 );
not \U$26951 ( \27328 , \27327 );
xor \U$26952 ( \27329 , \23851 , \23852 );
xor \U$26953 ( \27330 , \27329 , \23857 );
not \U$26954 ( \27331 , \27330 );
or \U$26955 ( \27332 , \27328 , \27331 );
or \U$26956 ( \27333 , \27330 , \27327 );
nand \U$26957 ( \27334 , \27332 , \27333 );
not \U$26958 ( \27335 , \27334 );
xor \U$26959 ( \27336 , \27214 , \27221 );
and \U$26960 ( \27337 , \27336 , \27224 );
and \U$26961 ( \27338 , \27214 , \27221 );
or \U$26962 ( \27339 , \27337 , \27338 );
not \U$26963 ( \27340 , \27339 );
not \U$26964 ( \27341 , \27340 );
or \U$26965 ( \27342 , \27335 , \27341 );
or \U$26966 ( \27343 , \27340 , \27334 );
nand \U$26967 ( \27344 , \27342 , \27343 );
not \U$26968 ( \27345 , \27344 );
not \U$26969 ( \27346 , \24122 );
not \U$26970 ( \27347 , \24066 );
not \U$26971 ( \27348 , \24073 );
or \U$26972 ( \27349 , \27347 , \27348 );
or \U$26973 ( \27350 , \24066 , \24073 );
nand \U$26974 ( \27351 , \27349 , \27350 );
not \U$26975 ( \27352 , \27351 );
or \U$26976 ( \27353 , \27346 , \27352 );
or \U$26977 ( \27354 , \27351 , \24122 );
nand \U$26978 ( \27355 , \27353 , \27354 );
not \U$26979 ( \27356 , \27355 );
xor \U$26980 ( \27357 , \27137 , \27142 );
and \U$26981 ( \27358 , \27357 , \27150 );
and \U$26982 ( \27359 , \27137 , \27142 );
or \U$26983 ( \27360 , \27358 , \27359 );
not \U$26984 ( \27361 , \27360 );
not \U$26985 ( \27362 , \27361 );
and \U$26986 ( \27363 , \27356 , \27362 );
and \U$26987 ( \27364 , \27355 , \27361 );
nor \U$26988 ( \27365 , \27363 , \27364 );
not \U$26989 ( \27366 , \27365 );
not \U$26990 ( \27367 , \27366 );
or \U$26991 ( \27368 , \27345 , \27367 );
not \U$26992 ( \27369 , \27361 );
nand \U$26993 ( \27370 , \27369 , \27355 );
nand \U$26994 ( \27371 , \27368 , \27370 );
not \U$26995 ( \27372 , \27371 );
xnor \U$26996 ( \27373 , \24135 , \24063 );
not \U$26997 ( \27374 , \27373 );
and \U$26998 ( \27375 , \27372 , \27374 );
and \U$26999 ( \27376 , \27371 , \27373 );
nor \U$27000 ( \27377 , \27375 , \27376 );
xor \U$27001 ( \27378 , \27325 , \27377 );
not \U$27002 ( \27379 , \27378 );
not \U$27003 ( \27380 , \27168 );
not \U$27004 ( \27381 , \27153 );
or \U$27005 ( \27382 , \27380 , \27381 );
nand \U$27006 ( \27383 , \27382 , \27157 );
not \U$27007 ( \27384 , \27383 );
not \U$27008 ( \27385 , \27365 );
not \U$27009 ( \27386 , \27344 );
and \U$27010 ( \27387 , \27385 , \27386 );
and \U$27011 ( \27388 , \27365 , \27344 );
nor \U$27012 ( \27389 , \27387 , \27388 );
not \U$27013 ( \27390 , \27389 );
or \U$27014 ( \27391 , \27384 , \27390 );
or \U$27015 ( \27392 , \27383 , \27389 );
nand \U$27016 ( \27393 , \27391 , \27392 );
not \U$27017 ( \27394 , \27393 );
not \U$27018 ( \27395 , \27320 );
not \U$27019 ( \27396 , \27305 );
or \U$27020 ( \27397 , \27395 , \27396 );
or \U$27021 ( \27398 , \27320 , \27305 );
nand \U$27022 ( \27399 , \27397 , \27398 );
not \U$27023 ( \27400 , \27399 );
or \U$27024 ( \27401 , \27394 , \27400 );
not \U$27025 ( \27402 , \27389 );
nand \U$27026 ( \27403 , \27402 , \27383 );
nand \U$27027 ( \27404 , \27401 , \27403 );
not \U$27028 ( \27405 , \27334 );
not \U$27029 ( \27406 , \27339 );
or \U$27030 ( \27407 , \27405 , \27406 );
not \U$27031 ( \27408 , \27330 );
nand \U$27032 ( \27409 , \27408 , \27327 );
nand \U$27033 ( \27410 , \27407 , \27409 );
xor \U$27034 ( \27411 , \23332 , \27410 );
not \U$27035 ( \27412 , \23615 );
xor \U$27036 ( \27413 , \27411 , \27412 );
not \U$27037 ( \27414 , \27413 );
xor \U$27038 ( \27415 , \27309 , \23440 );
xnor \U$27039 ( \27416 , \27415 , \23605 );
not \U$27040 ( \27417 , \27416 );
not \U$27041 ( \27418 , \27316 );
or \U$27042 ( \27419 , \27417 , \27418 );
not \U$27043 ( \27420 , \27309 );
nand \U$27044 ( \27421 , \27420 , \27319 );
nand \U$27045 ( \27422 , \27419 , \27421 );
not \U$27046 ( \27423 , \27422 );
not \U$27047 ( \27424 , \27423 );
and \U$27048 ( \27425 , \27414 , \27424 );
and \U$27049 ( \27426 , \27413 , \27423 );
nor \U$27050 ( \27427 , \27425 , \27426 );
xnor \U$27051 ( \27428 , \27404 , \27427 );
not \U$27052 ( \27429 , \27428 );
or \U$27053 ( \27430 , \27379 , \27429 );
or \U$27054 ( \27431 , \27378 , \27428 );
nand \U$27055 ( \27432 , \27430 , \27431 );
not \U$27056 ( \27433 , \27393 );
not \U$27057 ( \27434 , \27433 );
buf \U$27058 ( \27435 , \27399 );
not \U$27059 ( \27436 , \27435 );
or \U$27060 ( \27437 , \27434 , \27436 );
or \U$27061 ( \27438 , \27435 , \27433 );
nand \U$27062 ( \27439 , \27437 , \27438 );
not \U$27063 ( \27440 , \27439 );
not \U$27064 ( \27441 , \27176 );
not \U$27065 ( \27442 , \27170 );
or \U$27066 ( \27443 , \27441 , \27442 );
nand \U$27067 ( \27444 , \27443 , \27185 );
nand \U$27068 ( \27445 , \27171 , \27179 );
nand \U$27069 ( \27446 , \27444 , \27445 );
not \U$27070 ( \27447 , \27209 );
not \U$27071 ( \27448 , \27257 );
or \U$27072 ( \27449 , \27447 , \27448 );
not \U$27073 ( \27450 , \27191 );
nand \U$27074 ( \27451 , \27450 , \27204 );
nand \U$27075 ( \27452 , \27449 , \27451 );
xor \U$27076 ( \27453 , \27446 , \27452 );
not \U$27077 ( \27454 , \27453 );
not \U$27078 ( \27455 , \27454 );
or \U$27079 ( \27456 , \27440 , \27455 );
nand \U$27080 ( \27457 , \27444 , \27445 , \27452 );
nand \U$27081 ( \27458 , \27456 , \27457 );
nand \U$27082 ( \27459 , \27432 , \27458 );
not \U$27083 ( \27460 , \27272 );
not \U$27084 ( \27461 , \27186 );
not \U$27085 ( \27462 , \27461 );
or \U$27086 ( \27463 , \27460 , \27462 );
nand \U$27087 ( \27464 , \27265 , \27267 , \27259 );
nand \U$27088 ( \27465 , \27463 , \27464 );
xnor \U$27089 ( \27466 , \27439 , \27453 );
nand \U$27090 ( \27467 , \27465 , \27466 );
nand \U$27091 ( \27468 , \27459 , \27467 );
not \U$27092 ( \27469 , \27377 );
not \U$27093 ( \27470 , \27469 );
not \U$27094 ( \27471 , \27325 );
or \U$27095 ( \27472 , \27470 , \27471 );
not \U$27096 ( \27473 , \27373 );
nand \U$27097 ( \27474 , \27473 , \27371 );
nand \U$27098 ( \27475 , \27472 , \27474 );
not \U$27099 ( \27476 , \27475 );
not \U$27100 ( \27477 , \27422 );
not \U$27101 ( \27478 , \27413 );
or \U$27102 ( \27479 , \27477 , \27478 );
nand \U$27103 ( \27480 , \27412 , \23333 );
not \U$27104 ( \27481 , \27480 );
not \U$27105 ( \27482 , \27412 );
nand \U$27106 ( \27483 , \27482 , \23332 );
not \U$27107 ( \27484 , \27483 );
or \U$27108 ( \27485 , \27481 , \27484 );
nand \U$27109 ( \27486 , \27485 , \27410 );
nand \U$27110 ( \27487 , \27479 , \27486 );
not \U$27111 ( \27488 , \27487 );
not \U$27112 ( \27489 , \24148 );
not \U$27113 ( \27490 , \24146 );
and \U$27114 ( \27491 , \27489 , \27490 );
and \U$27115 ( \27492 , \24148 , \24146 );
nor \U$27116 ( \27493 , \27491 , \27492 );
not \U$27117 ( \27494 , \27493 );
or \U$27118 ( \27495 , \27488 , \27494 );
or \U$27119 ( \27496 , \27487 , \27493 );
nand \U$27120 ( \27497 , \27495 , \27496 );
not \U$27121 ( \27498 , \27497 );
or \U$27122 ( \27499 , \27476 , \27498 );
not \U$27123 ( \27500 , \27493 );
nand \U$27124 ( \27501 , \27500 , \27487 );
nand \U$27125 ( \27502 , \27499 , \27501 );
not \U$27126 ( \27503 , \27502 );
xor \U$27127 ( \27504 , \24157 , \24154 );
not \U$27128 ( \27505 , \24165 );
xnor \U$27129 ( \27506 , \27504 , \27505 );
not \U$27130 ( \27507 , \27506 );
or \U$27131 ( \27508 , \27503 , \27507 );
not \U$27132 ( \27509 , \27475 );
not \U$27133 ( \27510 , \27509 );
not \U$27134 ( \27511 , \27497 );
or \U$27135 ( \27512 , \27510 , \27511 );
or \U$27136 ( \27513 , \27497 , \27509 );
nand \U$27137 ( \27514 , \27512 , \27513 );
not \U$27138 ( \27515 , \27378 );
not \U$27139 ( \27516 , \27515 );
not \U$27140 ( \27517 , \27428 );
or \U$27141 ( \27518 , \27516 , \27517 );
not \U$27142 ( \27519 , \27427 );
nand \U$27143 ( \27520 , \27519 , \27404 );
nand \U$27144 ( \27521 , \27518 , \27520 );
nand \U$27145 ( \27522 , \27514 , \27521 );
nand \U$27146 ( \27523 , \27508 , \27522 );
nor \U$27147 ( \27524 , \27468 , \27523 );
and \U$27148 ( \27525 , \24261 , \27288 , \27524 );
not \U$27149 ( \27526 , \9644 );
not \U$27150 ( \27527 , RIae7a3a8_177);
not \U$27151 ( \27528 , \9657 );
or \U$27152 ( \27529 , \27527 , \27528 );
or \U$27153 ( \27530 , \1859 , RIae7a3a8_177);
nand \U$27154 ( \27531 , \27529 , \27530 );
not \U$27155 ( \27532 , \27531 );
or \U$27156 ( \27533 , \27526 , \27532 );
and \U$27157 ( \27534 , RIae7a3a8_177, \9672 );
not \U$27158 ( \27535 , RIae7a3a8_177);
and \U$27159 ( \27536 , \27535 , \17052 );
or \U$27160 ( \27537 , \27534 , \27536 );
nand \U$27161 ( \27538 , \27537 , \9622 );
nand \U$27162 ( \27539 , \27533 , \27538 );
not \U$27163 ( \27540 , \10667 );
and \U$27164 ( \27541 , RIae7a150_172, \1809 );
not \U$27165 ( \27542 , RIae7a150_172);
and \U$27166 ( \27543 , \27542 , \4036 );
or \U$27167 ( \27544 , \27541 , \27543 );
not \U$27168 ( \27545 , \27544 );
or \U$27169 ( \27546 , \27540 , \27545 );
and \U$27170 ( \27547 , \10658 , \4583 );
not \U$27171 ( \27548 , \10658 );
and \U$27172 ( \27549 , \27548 , \4582 );
nor \U$27173 ( \27550 , \27547 , \27549 );
nand \U$27174 ( \27551 , \27550 , \9776 );
nand \U$27175 ( \27552 , \27546 , \27551 );
xor \U$27176 ( \27553 , \27539 , \27552 );
not \U$27177 ( \27554 , \10519 );
and \U$27178 ( \27555 , RIae7a7e0_186, \2155 );
not \U$27179 ( \27556 , RIae7a7e0_186);
and \U$27180 ( \27557 , \27556 , \26329 );
or \U$27181 ( \27558 , \27555 , \27557 );
not \U$27182 ( \27559 , \27558 );
or \U$27183 ( \27560 , \27554 , \27559 );
not \U$27184 ( \27561 , \9529 );
not \U$27185 ( \27562 , \2309 );
or \U$27186 ( \27563 , \27561 , \27562 );
or \U$27187 ( \27564 , \2309 , \17112 );
nand \U$27188 ( \27565 , \27563 , \27564 );
nand \U$27189 ( \27566 , \27565 , \11851 );
nand \U$27190 ( \27567 , \27560 , \27566 );
xnor \U$27191 ( \27568 , \27553 , \27567 );
not \U$27192 ( \27569 , \27568 );
not \U$27193 ( \27570 , \27569 );
or \U$27194 ( \27571 , RIae79610_148, RIae799d0_156);
nand \U$27195 ( \27572 , \27571 , \12857 );
nand \U$27196 ( \27573 , \27572 , \8933 );
not \U$27197 ( \27574 , \27573 );
not \U$27198 ( \27575 , \1863 );
and \U$27199 ( \27576 , \16006 , \1902 );
not \U$27200 ( \27577 , \16006 );
and \U$27201 ( \27578 , \27577 , RIae793b8_143);
nor \U$27202 ( \27579 , \27576 , \27578 );
not \U$27203 ( \27580 , \27579 );
or \U$27204 ( \27581 , \27575 , \27580 );
and \U$27205 ( \27582 , RIae793b8_143, \12857 );
not \U$27206 ( \27583 , RIae793b8_143);
and \U$27207 ( \27584 , \27583 , \14601 );
nor \U$27208 ( \27585 , \27582 , \27584 );
nand \U$27209 ( \27586 , \27585 , \1909 );
nand \U$27210 ( \27587 , \27581 , \27586 );
nand \U$27211 ( \27588 , \27574 , \27587 );
not \U$27212 ( \27589 , \27588 );
not \U$27213 ( \27590 , \1820 );
and \U$27214 ( \27591 , RIae79688_149, \16909 );
not \U$27215 ( \27592 , RIae79688_149);
and \U$27216 ( \27593 , \27592 , \10042 );
or \U$27217 ( \27594 , \27591 , \27593 );
not \U$27218 ( \27595 , \27594 );
or \U$27219 ( \27596 , \27590 , \27595 );
not \U$27220 ( \27597 , \2970 );
not \U$27221 ( \27598 , \16035 );
or \U$27222 ( \27599 , \27597 , \27598 );
nand \U$27223 ( \27600 , \16036 , RIae79688_149);
nand \U$27224 ( \27601 , \27599 , \27600 );
nand \U$27225 ( \27602 , \27601 , \1842 );
nand \U$27226 ( \27603 , \27596 , \27602 );
not \U$27227 ( \27604 , \27603 );
or \U$27228 ( \27605 , \27589 , \27604 );
or \U$27229 ( \27606 , \27603 , \27588 );
nand \U$27230 ( \27607 , \27605 , \27606 );
buf \U$27231 ( \27608 , \27607 );
not \U$27232 ( \27609 , \2272 );
xor \U$27233 ( \27610 , RIae79ac0_158, \10031 );
not \U$27234 ( \27611 , \27610 );
or \U$27235 ( \27612 , \27609 , \27611 );
and \U$27236 ( \27613 , RIae79ac0_158, \10142 );
not \U$27237 ( \27614 , RIae79ac0_158);
and \U$27238 ( \27615 , \27614 , \10149 );
nor \U$27239 ( \27616 , \27613 , \27615 );
nand \U$27240 ( \27617 , \27616 , \2249 );
nand \U$27241 ( \27618 , \27612 , \27617 );
not \U$27242 ( \27619 , \27618 );
and \U$27243 ( \27620 , \27608 , \27619 );
not \U$27244 ( \27621 , \27608 );
and \U$27245 ( \27622 , \27621 , \27618 );
nor \U$27246 ( \27623 , \27620 , \27622 );
not \U$27247 ( \27624 , \27623 );
not \U$27248 ( \27625 , \11434 );
and \U$27249 ( \27626 , \2675 , RIae7a498_179);
not \U$27250 ( \27627 , \2675 );
not \U$27251 ( \27628 , RIae7a498_179);
and \U$27252 ( \27629 , \27627 , \27628 );
nor \U$27253 ( \27630 , \27626 , \27629 );
not \U$27254 ( \27631 , \27630 );
or \U$27255 ( \27632 , \27625 , \27631 );
and \U$27256 ( \27633 , RIae7a498_179, \18029 );
not \U$27257 ( \27634 , RIae7a498_179);
and \U$27258 ( \27635 , \27634 , \11681 );
nor \U$27259 ( \27636 , \27633 , \27635 );
nand \U$27260 ( \27637 , \27636 , \10675 );
nand \U$27261 ( \27638 , \27632 , \27637 );
not \U$27262 ( \27639 , \27638 );
or \U$27263 ( \27640 , \27624 , \27639 );
or \U$27264 ( \27641 , \27638 , \27623 );
nand \U$27265 ( \27642 , \27640 , \27641 );
not \U$27266 ( \27643 , \9478 );
not \U$27267 ( \27644 , RIae7a6f0_184);
not \U$27268 ( \27645 , \27644 );
not \U$27269 ( \27646 , \2994 );
or \U$27270 ( \27647 , \27645 , \27646 );
not \U$27271 ( \27648 , \11056 );
nand \U$27272 ( \27649 , \27648 , RIae7a6f0_184);
nand \U$27273 ( \27650 , \27647 , \27649 );
not \U$27274 ( \27651 , \27650 );
or \U$27275 ( \27652 , \27643 , \27651 );
not \U$27276 ( \27653 , RIae7a6f0_184);
not \U$27277 ( \27654 , \2140 );
or \U$27278 ( \27655 , \27653 , \27654 );
or \U$27279 ( \27656 , \19403 , RIae7a6f0_184);
nand \U$27280 ( \27657 , \27655 , \27656 );
nand \U$27281 ( \27658 , \27657 , \9473 );
nand \U$27282 ( \27659 , \27652 , \27658 );
and \U$27283 ( \27660 , \27642 , \27659 );
not \U$27284 ( \27661 , \27642 );
not \U$27285 ( \27662 , \27659 );
and \U$27286 ( \27663 , \27661 , \27662 );
nor \U$27287 ( \27664 , \27660 , \27663 );
not \U$27288 ( \27665 , \27664 );
not \U$27289 ( \27666 , \27665 );
or \U$27290 ( \27667 , \27570 , \27666 );
nand \U$27291 ( \27668 , \27664 , \27568 );
nand \U$27292 ( \27669 , \27667 , \27668 );
not \U$27293 ( \27670 , \10223 );
not \U$27294 ( \27671 , \16193 );
not \U$27295 ( \27672 , \27671 );
and \U$27296 ( \27673 , RIae79520_146, \27672 );
not \U$27297 ( \27674 , RIae79520_146);
not \U$27298 ( \27675 , \19035 );
and \U$27299 ( \27676 , \27674 , \27675 );
or \U$27300 ( \27677 , \27673 , \27676 );
not \U$27301 ( \27678 , \27677 );
or \U$27302 ( \27679 , \27670 , \27678 );
not \U$27303 ( \27680 , RIae79520_146);
not \U$27304 ( \27681 , \10149 );
or \U$27305 ( \27682 , \27680 , \27681 );
or \U$27306 ( \27683 , \10149 , RIae79520_146);
nand \U$27307 ( \27684 , \27682 , \27683 );
nand \U$27308 ( \27685 , \27684 , \12680 );
nand \U$27309 ( \27686 , \27679 , \27685 );
not \U$27310 ( \27687 , \2322 );
xnor \U$27311 ( \27688 , \11562 , RIae798e0_154);
not \U$27312 ( \27689 , \27688 );
or \U$27313 ( \27690 , \27687 , \27689 );
not \U$27314 ( \27691 , RIae798e0_154);
not \U$27315 ( \27692 , \9897 );
or \U$27316 ( \27693 , \27691 , \27692 );
or \U$27317 ( \27694 , \9897 , RIae798e0_154);
nand \U$27318 ( \27695 , \27693 , \27694 );
nand \U$27319 ( \27696 , \27695 , \2339 );
nand \U$27320 ( \27697 , \27690 , \27696 );
xor \U$27321 ( \27698 , \27686 , \27697 );
not \U$27322 ( \27699 , \2467 );
and \U$27323 ( \27700 , RIae794a8_145, \10750 );
not \U$27324 ( \27701 , RIae794a8_145);
and \U$27325 ( \27702 , \27701 , \9868 );
or \U$27326 ( \27703 , \27700 , \27702 );
not \U$27327 ( \27704 , \27703 );
or \U$27328 ( \27705 , \27699 , \27704 );
not \U$27329 ( \27706 , RIae794a8_145);
not \U$27330 ( \27707 , \9999 );
or \U$27331 ( \27708 , \27706 , \27707 );
or \U$27332 ( \27709 , \10000 , RIae794a8_145);
nand \U$27333 ( \27710 , \27708 , \27709 );
nand \U$27334 ( \27711 , \27710 , \1933 );
nand \U$27335 ( \27712 , \27705 , \27711 );
xor \U$27336 ( \27713 , \27698 , \27712 );
not \U$27337 ( \27714 , \27713 );
not \U$27338 ( \27715 , \10709 );
and \U$27339 ( \27716 , \6230 , RIae79fe8_169);
not \U$27340 ( \27717 , \6230 );
and \U$27341 ( \27718 , \27717 , \9504 );
nor \U$27342 ( \27719 , \27716 , \27718 );
not \U$27343 ( \27720 , \27719 );
or \U$27344 ( \27721 , \27715 , \27720 );
not \U$27345 ( \27722 , RIae79fe8_169);
not \U$27346 ( \27723 , \9286 );
or \U$27347 ( \27724 , \27722 , \27723 );
nand \U$27348 ( \27725 , \6345 , \18027 );
nand \U$27349 ( \27726 , \27724 , \27725 );
nand \U$27350 ( \27727 , \27726 , \9518 );
nand \U$27351 ( \27728 , \27721 , \27727 );
not \U$27352 ( \27729 , \27728 );
not \U$27353 ( \27730 , \14768 );
and \U$27354 ( \27731 , RIae79ef8_167, \15519 );
not \U$27355 ( \27732 , RIae79ef8_167);
and \U$27356 ( \27733 , \27732 , \17387 );
nor \U$27357 ( \27734 , \27731 , \27733 );
not \U$27358 ( \27735 , \27734 );
or \U$27359 ( \27736 , \27730 , \27735 );
and \U$27360 ( \27737 , \22389 , \16271 );
not \U$27361 ( \27738 , \22389 );
and \U$27362 ( \27739 , \27738 , \16274 );
nor \U$27363 ( \27740 , \27737 , \27739 );
nand \U$27364 ( \27741 , \27740 , \6214 );
nand \U$27365 ( \27742 , \27736 , \27741 );
not \U$27366 ( \27743 , \1820 );
xnor \U$27367 ( \27744 , RIae79688_149, \17155 );
not \U$27368 ( \27745 , \27744 );
or \U$27369 ( \27746 , \27743 , \27745 );
not \U$27370 ( \27747 , RIae79688_149);
not \U$27371 ( \27748 , \10844 );
or \U$27372 ( \27749 , \27747 , \27748 );
or \U$27373 ( \27750 , \10844 , RIae79688_149);
nand \U$27374 ( \27751 , \27749 , \27750 );
nand \U$27375 ( \27752 , \27751 , \1842 );
nand \U$27376 ( \27753 , \27746 , \27752 );
not \U$27377 ( \27754 , \27753 );
not \U$27378 ( \27755 , \2011 );
not \U$27379 ( \27756 , RIae79610_148);
not \U$27380 ( \27757 , \12750 );
or \U$27381 ( \27758 , \27756 , \27757 );
or \U$27382 ( \27759 , \12750 , RIae79610_148);
nand \U$27383 ( \27760 , \27758 , \27759 );
not \U$27384 ( \27761 , \27760 );
or \U$27385 ( \27762 , \27755 , \27761 );
or \U$27386 ( \27763 , \12857 , \2056 );
or \U$27387 ( \27764 , \16890 , RIae79610_148);
nand \U$27388 ( \27765 , \27763 , \27764 );
nand \U$27389 ( \27766 , \27765 , \2062 );
nand \U$27390 ( \27767 , \27762 , \27766 );
not \U$27391 ( \27768 , \2057 );
not \U$27392 ( \27769 , \2970 );
or \U$27393 ( \27770 , \27768 , \27769 );
nand \U$27394 ( \27771 , \27770 , \12857 );
nand \U$27395 ( \27772 , \27771 , \8668 );
xor \U$27396 ( \27773 , \27767 , \27772 );
not \U$27397 ( \27774 , \27773 );
or \U$27398 ( \27775 , \27754 , \27774 );
or \U$27399 ( \27776 , \27753 , \27773 );
nand \U$27400 ( \27777 , \27775 , \27776 );
not \U$27401 ( \27778 , \27777 );
not \U$27402 ( \27779 , \2162 );
and \U$27403 ( \27780 , RIae79520_146, \10337 );
not \U$27404 ( \27781 , RIae79520_146);
and \U$27405 ( \27782 , \27781 , \10031 );
or \U$27406 ( \27783 , \27780 , \27782 );
not \U$27407 ( \27784 , \27783 );
or \U$27408 ( \27785 , \27779 , \27784 );
not \U$27409 ( \27786 , RIae79520_146);
not \U$27410 ( \27787 , \27786 );
not \U$27411 ( \27788 , \10047 );
or \U$27412 ( \27789 , \27787 , \27788 );
or \U$27413 ( \27790 , \16912 , \2183 );
nand \U$27414 ( \27791 , \27789 , \27790 );
nand \U$27415 ( \27792 , \27791 , \2188 );
nand \U$27416 ( \27793 , \27785 , \27792 );
not \U$27417 ( \27794 , \27793 );
or \U$27418 ( \27795 , \27778 , \27794 );
not \U$27419 ( \27796 , \27773 );
nand \U$27420 ( \27797 , \27796 , \27753 );
nand \U$27421 ( \27798 , \27795 , \27797 );
and \U$27422 ( \27799 , \27742 , \27798 );
not \U$27423 ( \27800 , \27742 );
not \U$27424 ( \27801 , \27798 );
and \U$27425 ( \27802 , \27800 , \27801 );
nor \U$27426 ( \27803 , \27799 , \27802 );
not \U$27427 ( \27804 , \27803 );
or \U$27428 ( \27805 , \27729 , \27804 );
not \U$27429 ( \27806 , \27742 );
not \U$27430 ( \27807 , \27806 );
nand \U$27431 ( \27808 , \27807 , \27798 );
nand \U$27432 ( \27809 , \27805 , \27808 );
not \U$27433 ( \27810 , \27809 );
or \U$27434 ( \27811 , \27714 , \27810 );
or \U$27435 ( \27812 , \27809 , \27713 );
not \U$27436 ( \27813 , \9643 );
xor \U$27437 ( \27814 , RIae7a3a8_177, \10328 );
not \U$27438 ( \27815 , \27814 );
or \U$27439 ( \27816 , \27813 , \27815 );
not \U$27440 ( \27817 , RIae7a3a8_177);
not \U$27441 ( \27818 , \3270 );
or \U$27442 ( \27819 , \27817 , \27818 );
or \U$27443 ( \27820 , \2402 , RIae7a3a8_177);
nand \U$27444 ( \27821 , \27819 , \27820 );
nand \U$27445 ( \27822 , \27821 , \9622 );
nand \U$27446 ( \27823 , \27816 , \27822 );
not \U$27447 ( \27824 , \27823 );
not \U$27448 ( \27825 , \9814 );
not \U$27449 ( \27826 , RIae7a2b8_175);
not \U$27450 ( \27827 , \6256 );
not \U$27451 ( \27828 , \27827 );
or \U$27452 ( \27829 , \27826 , \27828 );
or \U$27453 ( \27830 , \27827 , RIae7a2b8_175);
nand \U$27454 ( \27831 , \27829 , \27830 );
not \U$27455 ( \27832 , \27831 );
or \U$27456 ( \27833 , \27825 , \27832 );
and \U$27457 ( \27834 , RIae7a2b8_175, \12334 );
not \U$27458 ( \27835 , RIae7a2b8_175);
and \U$27459 ( \27836 , \27835 , \5722 );
or \U$27460 ( \27837 , \27834 , \27836 );
nand \U$27461 ( \27838 , \27837 , \9792 );
nand \U$27462 ( \27839 , \27833 , \27838 );
not \U$27463 ( \27840 , \27839 );
or \U$27464 ( \27841 , \27824 , \27840 );
and \U$27465 ( \27842 , RIae7a240_174, \6238 );
not \U$27466 ( \27843 , RIae7a240_174);
and \U$27467 ( \27844 , \27843 , \4169 );
or \U$27468 ( \27845 , \27842 , \27844 );
and \U$27469 ( \27846 , \9699 , \27845 );
xor \U$27470 ( \27847 , \10829 , RIae7a240_174);
not \U$27471 ( \27848 , \27847 );
and \U$27472 ( \27849 , \27848 , \19466 );
nor \U$27473 ( \27850 , \27846 , \27849 );
nand \U$27474 ( \27851 , \27841 , \27850 );
not \U$27475 ( \27852 , \27823 );
not \U$27476 ( \27853 , \27839 );
nand \U$27477 ( \27854 , \27852 , \27853 );
and \U$27478 ( \27855 , \27851 , \27854 );
nand \U$27479 ( \27856 , \27812 , \27855 );
nand \U$27480 ( \27857 , \27811 , \27856 );
nand \U$27481 ( \27858 , \27669 , \27857 );
not \U$27482 ( \27859 , RIae7aab0_192);
and \U$27483 ( \27860 , \13032 , RIae7aa38_191);
not \U$27484 ( \27861 , \13032 );
and \U$27485 ( \27862 , \27861 , \11326 );
nor \U$27486 ( \27863 , \27860 , \27862 );
not \U$27487 ( \27864 , \27863 );
or \U$27488 ( \27865 , \27859 , \27864 );
xnor \U$27489 ( \27866 , RIae7aa38_191, \1878 );
nand \U$27490 ( \27867 , \27866 , \14668 );
nand \U$27491 ( \27868 , \27865 , \27867 );
not \U$27492 ( \27869 , \9730 );
and \U$27493 ( \27870 , RIae7a060_170, \4024 );
not \U$27494 ( \27871 , RIae7a060_170);
and \U$27495 ( \27872 , \27871 , \4023 );
or \U$27496 ( \27873 , \27870 , \27872 );
not \U$27497 ( \27874 , \27873 );
or \U$27498 ( \27875 , \27869 , \27874 );
xor \U$27499 ( \27876 , RIae7a060_170, \3747 );
nand \U$27500 ( \27877 , \27876 , \9745 );
nand \U$27501 ( \27878 , \27875 , \27877 );
xor \U$27502 ( \27879 , \27868 , \27878 );
not \U$27503 ( \27880 , \17847 );
not \U$27504 ( \27881 , RIae7a8d0_188);
not \U$27505 ( \27882 , \9797 );
or \U$27506 ( \27883 , \27881 , \27882 );
or \U$27507 ( \27884 , \9797 , RIae7a8d0_188);
nand \U$27508 ( \27885 , \27883 , \27884 );
not \U$27509 ( \27886 , \27885 );
or \U$27510 ( \27887 , \27880 , \27886 );
and \U$27511 ( \27888 , RIae7a8d0_188, \1898 );
not \U$27512 ( \27889 , RIae7a8d0_188);
and \U$27513 ( \27890 , \27889 , \9806 );
nor \U$27514 ( \27891 , \27888 , \27890 );
nand \U$27515 ( \27892 , \27891 , \10275 );
nand \U$27516 ( \27893 , \27887 , \27892 );
xor \U$27517 ( \27894 , \27879 , \27893 );
not \U$27518 ( \27895 , \27894 );
not \U$27519 ( \27896 , \27895 );
not \U$27520 ( \27897 , \10631 );
and \U$27521 ( \27898 , RIae7a510_180, \4112 );
not \U$27522 ( \27899 , RIae7a510_180);
and \U$27523 ( \27900 , \27899 , \2356 );
or \U$27524 ( \27901 , \27898 , \27900 );
not \U$27525 ( \27902 , \27901 );
or \U$27526 ( \27903 , \27897 , \27902 );
not \U$27527 ( \27904 , RIae7a510_180);
not \U$27528 ( \27905 , \1969 );
or \U$27529 ( \27906 , \27904 , \27905 );
or \U$27530 ( \27907 , \1969 , RIae7a510_180);
nand \U$27531 ( \27908 , \27906 , \27907 );
nand \U$27532 ( \27909 , \27908 , \10638 );
nand \U$27533 ( \27910 , \27903 , \27909 );
not \U$27534 ( \27911 , \27910 );
not \U$27535 ( \27912 , \9527 );
not \U$27536 ( \27913 , \27565 );
or \U$27537 ( \27914 , \27912 , \27913 );
not \U$27538 ( \27915 , RIae7a7e0_186);
not \U$27539 ( \27916 , \10534 );
or \U$27540 ( \27917 , \27915 , \27916 );
or \U$27541 ( \27918 , \2835 , RIae7a7e0_186);
nand \U$27542 ( \27919 , \27917 , \27918 );
nand \U$27543 ( \27920 , \27919 , \10510 );
nand \U$27544 ( \27921 , \27914 , \27920 );
not \U$27545 ( \27922 , \4853 );
and \U$27546 ( \27923 , RIae79ca0_162, \9438 );
not \U$27547 ( \27924 , RIae79ca0_162);
and \U$27548 ( \27925 , \27924 , \20941 );
nor \U$27549 ( \27926 , \27923 , \27925 );
not \U$27550 ( \27927 , \27926 );
or \U$27551 ( \27928 , \27922 , \27927 );
not \U$27552 ( \27929 , RIae79ca0_162);
not \U$27553 ( \27930 , \21948 );
or \U$27554 ( \27931 , \27929 , \27930 );
nand \U$27555 ( \27932 , \9459 , \11755 );
nand \U$27556 ( \27933 , \27931 , \27932 );
nand \U$27557 ( \27934 , \27933 , \11762 );
nand \U$27558 ( \27935 , \27928 , \27934 );
and \U$27559 ( \27936 , \27921 , \27935 );
not \U$27560 ( \27937 , \27921 );
not \U$27561 ( \27938 , \27935 );
and \U$27562 ( \27939 , \27937 , \27938 );
nor \U$27563 ( \27940 , \27936 , \27939 );
not \U$27564 ( \27941 , \27940 );
or \U$27565 ( \27942 , \27911 , \27941 );
not \U$27566 ( \27943 , \27938 );
nand \U$27567 ( \27944 , \27943 , \27921 );
nand \U$27568 ( \27945 , \27942 , \27944 );
not \U$27569 ( \27946 , \27945 );
not \U$27570 ( \27947 , \27946 );
or \U$27571 ( \27948 , \27896 , \27947 );
not \U$27572 ( \27949 , \27894 );
not \U$27573 ( \27950 , \27945 );
or \U$27574 ( \27951 , \27949 , \27950 );
not \U$27575 ( \27952 , \10676 );
not \U$27576 ( \27953 , \27630 );
or \U$27577 ( \27954 , \27952 , \27953 );
not \U$27578 ( \27955 , RIae7a498_179);
not \U$27579 ( \27956 , \13008 );
or \U$27580 ( \27957 , \27955 , \27956 );
nand \U$27581 ( \27958 , \2093 , \27628 );
nand \U$27582 ( \27959 , \27957 , \27958 );
nand \U$27583 ( \27960 , \27959 , \16564 );
nand \U$27584 ( \27961 , \27954 , \27960 );
not \U$27585 ( \27962 , \27961 );
nand \U$27586 ( \27963 , \12857 , \1863 );
not \U$27587 ( \27964 , \27963 );
not \U$27588 ( \27965 , \2011 );
not \U$27589 ( \27966 , RIae79610_148);
not \U$27590 ( \27967 , \10844 );
or \U$27591 ( \27968 , \27966 , \27967 );
or \U$27592 ( \27969 , \16165 , RIae79610_148);
nand \U$27593 ( \27970 , \27968 , \27969 );
not \U$27594 ( \27971 , \27970 );
or \U$27595 ( \27972 , \27965 , \27971 );
nand \U$27596 ( \27973 , \27760 , \2062 );
nand \U$27597 ( \27974 , \27972 , \27973 );
not \U$27598 ( \27975 , \27974 );
or \U$27599 ( \27976 , \27964 , \27975 );
or \U$27600 ( \27977 , \27974 , \27963 );
nand \U$27601 ( \27978 , \27976 , \27977 );
not \U$27602 ( \27979 , \27744 );
not \U$27603 ( \27980 , \1842 );
or \U$27604 ( \27981 , \27979 , \27980 );
not \U$27605 ( \27982 , \11317 );
not \U$27606 ( \27983 , \2970 );
and \U$27607 ( \27984 , \27982 , \27983 );
and \U$27608 ( \27985 , \10272 , \2970 );
nor \U$27609 ( \27986 , \27984 , \27985 );
or \U$27610 ( \27987 , \27986 , \1819 );
nand \U$27611 ( \27988 , \27981 , \27987 );
xor \U$27612 ( \27989 , \27978 , \27988 );
not \U$27613 ( \27990 , \1932 );
not \U$27614 ( \27991 , RIae794a8_145);
not \U$27615 ( \27992 , \16193 );
or \U$27616 ( \27993 , \27991 , \27992 );
or \U$27617 ( \27994 , \9989 , RIae794a8_145);
nand \U$27618 ( \27995 , \27993 , \27994 );
not \U$27619 ( \27996 , \27995 );
or \U$27620 ( \27997 , \27990 , \27996 );
nand \U$27621 ( \27998 , \27710 , \1919 );
nand \U$27622 ( \27999 , \27997 , \27998 );
xor \U$27623 ( \28000 , \27989 , \27999 );
not \U$27624 ( \28001 , \2339 );
xnor \U$27625 ( \28002 , \10749 , RIae798e0_154);
not \U$27626 ( \28003 , \28002 );
or \U$27627 ( \28004 , \28001 , \28003 );
nand \U$27628 ( \28005 , \27695 , \2321 );
nand \U$27629 ( \28006 , \28004 , \28005 );
and \U$27630 ( \28007 , \28000 , \28006 );
and \U$27631 ( \28008 , \27989 , \27999 );
nor \U$27632 ( \28009 , \28007 , \28008 );
not \U$27633 ( \28010 , \28009 );
not \U$27634 ( \28011 , RIae797f0_152);
not \U$27635 ( \28012 , \16826 );
or \U$27636 ( \28013 , \28011 , \28012 );
not \U$27637 ( \28014 , \9917 );
not \U$27638 ( \28015 , \9919 );
and \U$27639 ( \28016 , \28014 , \28015 );
and \U$27640 ( \28017 , \9917 , \9919 );
nor \U$27641 ( \28018 , \28016 , \28017 );
not \U$27642 ( \28019 , \28018 );
nand \U$27643 ( \28020 , \28019 , \2521 );
nand \U$27644 ( \28021 , \28013 , \28020 );
and \U$27645 ( \28022 , \2007 , \28021 );
not \U$27646 ( \28023 , RIae797f0_152);
not \U$27647 ( \28024 , \10083 );
or \U$27648 ( \28025 , \28023 , \28024 );
nand \U$27649 ( \28026 , \10207 , \2521 );
nand \U$27650 ( \28027 , \28025 , \28026 );
and \U$27651 ( \28028 , \28027 , \1988 );
nor \U$27652 ( \28029 , \28022 , \28028 );
not \U$27653 ( \28030 , \28029 );
not \U$27654 ( \28031 , \27988 );
not \U$27655 ( \28032 , \27978 );
or \U$27656 ( \28033 , \28031 , \28032 );
not \U$27657 ( \28034 , \27963 );
nand \U$27658 ( \28035 , \28034 , \27974 );
nand \U$27659 ( \28036 , \28033 , \28035 );
not \U$27660 ( \28037 , \2249 );
not \U$27661 ( \28038 , \27610 );
or \U$27662 ( \28039 , \28037 , \28038 );
and \U$27663 ( \28040 , RIae79ac0_158, \10042 );
not \U$27664 ( \28041 , RIae79ac0_158);
not \U$27665 ( \28042 , \10042 );
and \U$27666 ( \28043 , \28041 , \28042 );
nor \U$27667 ( \28044 , \28040 , \28043 );
nand \U$27668 ( \28045 , \28044 , \2272 );
nand \U$27669 ( \28046 , \28039 , \28045 );
xor \U$27670 ( \28047 , \28036 , \28046 );
not \U$27671 ( \28048 , \28047 );
or \U$27672 ( \28049 , \28030 , \28048 );
or \U$27673 ( \28050 , \28029 , \28047 );
nand \U$27674 ( \28051 , \28049 , \28050 );
not \U$27675 ( \28052 , \28051 );
or \U$27676 ( \28053 , \28010 , \28052 );
or \U$27677 ( \28054 , \28051 , \28009 );
nand \U$27678 ( \28055 , \28053 , \28054 );
not \U$27679 ( \28056 , \28055 );
or \U$27680 ( \28057 , \27962 , \28056 );
not \U$27681 ( \28058 , \28009 );
nand \U$27682 ( \28059 , \28058 , \28051 );
nand \U$27683 ( \28060 , \28057 , \28059 );
not \U$27684 ( \28061 , \28060 );
nand \U$27685 ( \28062 , \27951 , \28061 );
nand \U$27686 ( \28063 , \27948 , \28062 );
nand \U$27687 ( \28064 , \27664 , \27569 );
and \U$27688 ( \28065 , \27858 , \28063 , \28064 );
not \U$27689 ( \28066 , \28065 );
not \U$27690 ( \28067 , \28064 );
not \U$27691 ( \28068 , \27858 );
or \U$27692 ( \28069 , \28067 , \28068 );
not \U$27693 ( \28070 , \28063 );
nand \U$27694 ( \28071 , \28069 , \28070 );
not \U$27695 ( \28072 , \13121 );
not \U$27696 ( \28073 , RIae7a240_174);
not \U$27697 ( \28074 , \9657 );
or \U$27698 ( \28075 , \28073 , \28074 );
or \U$27699 ( \28076 , \9657 , RIae7a240_174);
nand \U$27700 ( \28077 , \28075 , \28076 );
not \U$27701 ( \28078 , \28077 );
or \U$27702 ( \28079 , \28072 , \28078 );
xnor \U$27703 ( \28080 , \2402 , RIae7a240_174);
nand \U$27704 ( \28081 , \28080 , \9688 );
nand \U$27705 ( \28082 , \28079 , \28081 );
not \U$27706 ( \28083 , \9622 );
xor \U$27707 ( \28084 , RIae7a3a8_177, \2356 );
not \U$27708 ( \28085 , \28084 );
or \U$27709 ( \28086 , \28083 , \28085 );
nand \U$27710 ( \28087 , \27537 , \9644 );
nand \U$27711 ( \28088 , \28086 , \28087 );
xor \U$27712 ( \28089 , \28082 , \28088 );
not \U$27713 ( \28090 , \10519 );
not \U$27714 ( \28091 , RIae7a7e0_186);
not \U$27715 ( \28092 , \10570 );
or \U$27716 ( \28093 , \28091 , \28092 );
or \U$27717 ( \28094 , \19400 , RIae7a7e0_186);
nand \U$27718 ( \28095 , \28093 , \28094 );
not \U$27719 ( \28096 , \28095 );
or \U$27720 ( \28097 , \28090 , \28096 );
nand \U$27721 ( \28098 , \27558 , \11851 );
nand \U$27722 ( \28099 , \28097 , \28098 );
xor \U$27723 ( \28100 , \28089 , \28099 );
not \U$27724 ( \28101 , \4853 );
not \U$27725 ( \28102 , \9347 );
xor \U$27726 ( \28103 , RIae79ca0_162, \28102 );
not \U$27727 ( \28104 , \28103 );
or \U$27728 ( \28105 , \28101 , \28104 );
xnor \U$27729 ( \28106 , \16254 , RIae79ca0_162);
nand \U$27730 ( \28107 , \28106 , \16804 );
nand \U$27731 ( \28108 , \28105 , \28107 );
not \U$27732 ( \28109 , \16358 );
not \U$27733 ( \28110 , RIae7a510_180);
not \U$27734 ( \28111 , \3417 );
or \U$27735 ( \28112 , \28110 , \28111 );
or \U$27736 ( \28113 , \13942 , RIae7a510_180);
nand \U$27737 ( \28114 , \28112 , \28113 );
not \U$27738 ( \28115 , \28114 );
or \U$27739 ( \28116 , \28109 , \28115 );
not \U$27740 ( \28117 , RIae7a510_180);
not \U$27741 ( \28118 , \14439 );
or \U$27742 ( \28119 , \28117 , \28118 );
or \U$27743 ( \28120 , \14439 , RIae7a510_180);
nand \U$27744 ( \28121 , \28119 , \28120 );
nand \U$27745 ( \28122 , \10637 , \28121 );
nand \U$27746 ( \28123 , \28116 , \28122 );
and \U$27747 ( \28124 , \28108 , \28123 );
not \U$27748 ( \28125 , \28108 );
not \U$27749 ( \28126 , \28123 );
and \U$27750 ( \28127 , \28125 , \28126 );
nor \U$27751 ( \28128 , \28124 , \28127 );
not \U$27752 ( \28129 , \14667 );
not \U$27753 ( \28130 , \27863 );
or \U$27754 ( \28131 , \28129 , \28130 );
not \U$27755 ( \28132 , RIae7aa38_191);
not \U$27756 ( \28133 , \10444 );
or \U$27757 ( \28134 , \28132 , \28133 );
or \U$27758 ( \28135 , \2030 , RIae7aa38_191);
nand \U$27759 ( \28136 , \28134 , \28135 );
nand \U$27760 ( \28137 , \28136 , RIae7aab0_192);
nand \U$27761 ( \28138 , \28131 , \28137 );
not \U$27762 ( \28139 , \28138 );
and \U$27763 ( \28140 , \28128 , \28139 );
not \U$27764 ( \28141 , \28128 );
and \U$27765 ( \28142 , \28141 , \28138 );
nor \U$27766 ( \28143 , \28140 , \28142 );
not \U$27767 ( \28144 , \28143 );
not \U$27768 ( \28145 , \10275 );
not \U$27769 ( \28146 , RIae7a8d0_188);
not \U$27770 ( \28147 , \4197 );
or \U$27771 ( \28148 , \28146 , \28147 );
or \U$27772 ( \28149 , \4197 , RIae7a8d0_188);
nand \U$27773 ( \28150 , \28148 , \28149 );
not \U$27774 ( \28151 , \28150 );
or \U$27775 ( \28152 , \28145 , \28151 );
nand \U$27776 ( \28153 , \27891 , \14510 );
nand \U$27777 ( \28154 , \28152 , \28153 );
not \U$27778 ( \28155 , \9729 );
not \U$27779 ( \28156 , \27876 );
or \U$27780 ( \28157 , \28155 , \28156 );
not \U$27781 ( \28158 , \9749 );
not \U$27782 ( \28159 , \2309 );
or \U$27783 ( \28160 , \28158 , \28159 );
nand \U$27784 ( \28161 , \2305 , RIae7a060_170);
nand \U$27785 ( \28162 , \28160 , \28161 );
nand \U$27786 ( \28163 , \28162 , \9745 );
nand \U$27787 ( \28164 , \28157 , \28163 );
xor \U$27788 ( \28165 , \28154 , \28164 );
not \U$27789 ( \28166 , \9776 );
not \U$27790 ( \28167 , \10658 );
not \U$27791 ( \28168 , \4023 );
or \U$27792 ( \28169 , \28167 , \28168 );
or \U$27793 ( \28170 , \4023 , \10658 );
nand \U$27794 ( \28171 , \28169 , \28170 );
not \U$27795 ( \28172 , \28171 );
or \U$27796 ( \28173 , \28166 , \28172 );
nand \U$27797 ( \28174 , \27550 , \9758 );
nand \U$27798 ( \28175 , \28173 , \28174 );
xnor \U$27799 ( \28176 , \28165 , \28175 );
not \U$27800 ( \28177 , \28176 );
and \U$27801 ( \28178 , \28144 , \28177 );
not \U$27802 ( \28179 , \28144 );
and \U$27803 ( \28180 , \28179 , \28176 );
nor \U$27804 ( \28181 , \28178 , \28180 );
not \U$27805 ( \28182 , \28181 );
xor \U$27806 ( \28183 , \28100 , \28182 );
nand \U$27807 ( \28184 , \28071 , \28183 );
nand \U$27808 ( \28185 , \28066 , \28184 );
not \U$27809 ( \28186 , \28185 );
not \U$27810 ( \28187 , \9792 );
not \U$27811 ( \28188 , RIae7a2b8_175);
not \U$27812 ( \28189 , \10226 );
or \U$27813 ( \28190 , \28188 , \28189 );
or \U$27814 ( \28191 , \4960 , RIae7a2b8_175);
nand \U$27815 ( \28192 , \28190 , \28191 );
not \U$27816 ( \28193 , \28192 );
or \U$27817 ( \28194 , \28187 , \28193 );
not \U$27818 ( \28195 , RIae7a2b8_175);
not \U$27819 ( \28196 , \6238 );
or \U$27820 ( \28197 , \28195 , \28196 );
not \U$27821 ( \28198 , RIae7a2b8_175);
nand \U$27822 ( \28199 , \4169 , \28198 );
nand \U$27823 ( \28200 , \28197 , \28199 );
nand \U$27824 ( \28201 , \28200 , \16135 );
nand \U$27825 ( \28202 , \28194 , \28201 );
not \U$27826 ( \28203 , \28202 );
not \U$27827 ( \28204 , \2432 );
and \U$27828 ( \28205 , \9607 , RIae79778_151);
not \U$27829 ( \28206 , \9607 );
and \U$27830 ( \28207 , \28206 , \2447 );
nor \U$27831 ( \28208 , \28205 , \28207 );
not \U$27832 ( \28209 , \28208 );
or \U$27833 ( \28210 , \28204 , \28209 );
not \U$27834 ( \28211 , \2447 );
not \U$27835 ( \28212 , \15947 );
or \U$27836 ( \28213 , \28211 , \28212 );
or \U$27837 ( \28214 , \11803 , \2447 );
nand \U$27838 ( \28215 , \28213 , \28214 );
nand \U$27839 ( \28216 , \28215 , \15337 );
nand \U$27840 ( \28217 , \28210 , \28216 );
not \U$27841 ( \28218 , \2417 );
not \U$27842 ( \28219 , RIae79c28_161);
not \U$27843 ( \28220 , \15488 );
or \U$27844 ( \28221 , \28219 , \28220 );
or \U$27845 ( \28222 , \15488 , RIae79c28_161);
nand \U$27846 ( \28223 , \28221 , \28222 );
not \U$27847 ( \28224 , \28223 );
or \U$27848 ( \28225 , \28218 , \28224 );
not \U$27849 ( \28226 , RIae79c28_161);
not \U$27850 ( \28227 , \9456 );
or \U$27851 ( \28228 , \28226 , \28227 );
nand \U$27852 ( \28229 , \9455 , \10584 );
nand \U$27853 ( \28230 , \28228 , \28229 );
nand \U$27854 ( \28231 , \28230 , \2418 );
nand \U$27855 ( \28232 , \28225 , \28231 );
and \U$27856 ( \28233 , \28217 , \28232 );
not \U$27857 ( \28234 , \28233 );
and \U$27858 ( \28235 , \28203 , \28234 );
nor \U$27859 ( \28236 , \28232 , \28217 );
nor \U$27860 ( \28237 , \28235 , \28236 );
not \U$27861 ( \28238 , \28237 );
not \U$27862 ( \28239 , \1863 );
not \U$27863 ( \28240 , RIae793b8_143);
not \U$27864 ( \28241 , \16651 );
or \U$27865 ( \28242 , \28240 , \28241 );
not \U$27866 ( \28243 , \16164 );
or \U$27867 ( \28244 , \28243 , RIae793b8_143);
nand \U$27868 ( \28245 , \28242 , \28244 );
not \U$27869 ( \28246 , \28245 );
or \U$27870 ( \28247 , \28239 , \28246 );
nand \U$27871 ( \28248 , \27579 , \1909 );
nand \U$27872 ( \28249 , \28247 , \28248 );
and \U$27873 ( \28250 , \12857 , \1501 );
nor \U$27874 ( \28251 , \28249 , \28250 );
not \U$27875 ( \28252 , \28251 );
nand \U$27876 ( \28253 , \28249 , \28250 );
nand \U$27877 ( \28254 , \28252 , \28253 );
not \U$27878 ( \28255 , \10272 );
not \U$27879 ( \28256 , \2056 );
and \U$27880 ( \28257 , \28255 , \28256 );
not \U$27881 ( \28258 , \11317 );
not \U$27882 ( \28259 , \28258 );
and \U$27883 ( \28260 , \28259 , \10957 );
nor \U$27884 ( \28261 , \28257 , \28260 );
not \U$27885 ( \28262 , \28261 );
not \U$27886 ( \28263 , \7887 );
and \U$27887 ( \28264 , \28262 , \28263 );
and \U$27888 ( \28265 , RIae79610_148, \10259 );
not \U$27889 ( \28266 , RIae79610_148);
not \U$27890 ( \28267 , \10259 );
and \U$27891 ( \28268 , \28266 , \28267 );
nor \U$27892 ( \28269 , \28265 , \28268 );
nor \U$27893 ( \28270 , \28269 , \8320 );
nor \U$27894 ( \28271 , \28264 , \28270 );
xor \U$27895 ( \28272 , \28254 , \28271 );
not \U$27896 ( \28273 , \2188 );
not \U$27897 ( \28274 , \27677 );
or \U$27898 ( \28275 , \28273 , \28274 );
not \U$27899 ( \28276 , RIae79520_146);
not \U$27900 ( \28277 , \16719 );
or \U$27901 ( \28278 , \28276 , \28277 );
or \U$27902 ( \28279 , \10000 , RIae79520_146);
nand \U$27903 ( \28280 , \28278 , \28279 );
nand \U$27904 ( \28281 , \28280 , \2163 );
nand \U$27905 ( \28282 , \28275 , \28281 );
nand \U$27906 ( \28283 , \28272 , \28282 );
not \U$27907 ( \28284 , \28283 );
and \U$27908 ( \28285 , \28021 , \1989 );
and \U$27909 ( \28286 , \10464 , \2521 );
not \U$27910 ( \28287 , \10464 );
and \U$27911 ( \28288 , \28287 , RIae797f0_152);
nor \U$27912 ( \28289 , \28286 , \28288 );
and \U$27913 ( \28290 , \28289 , \2007 );
nor \U$27914 ( \28291 , \28285 , \28290 );
not \U$27915 ( \28292 , \28291 );
or \U$27916 ( \28293 , \28284 , \28292 );
or \U$27917 ( \28294 , \28282 , \28272 );
nand \U$27918 ( \28295 , \28293 , \28294 );
not \U$27919 ( \28296 , \14768 );
and \U$27920 ( \28297 , \16260 , \12209 );
not \U$27921 ( \28298 , \16260 );
and \U$27922 ( \28299 , \28298 , RIae79ef8_167);
nor \U$27923 ( \28300 , \28297 , \28299 );
not \U$27924 ( \28301 , \28300 );
or \U$27925 ( \28302 , \28296 , \28301 );
not \U$27926 ( \28303 , RIae79ef8_167);
not \U$27927 ( \28304 , \28303 );
not \U$27928 ( \28305 , \10406 );
not \U$27929 ( \28306 , \28305 );
or \U$27930 ( \28307 , \28304 , \28306 );
nand \U$27931 ( \28308 , \6346 , RIae79ef8_167);
nand \U$27932 ( \28309 , \28307 , \28308 );
nand \U$27933 ( \28310 , \28309 , \10573 );
nand \U$27934 ( \28311 , \28302 , \28310 );
not \U$27935 ( \28312 , \6091 );
not \U$27936 ( \28313 , RIae79d90_164);
not \U$27937 ( \28314 , \12707 );
or \U$27938 ( \28315 , \28313 , \28314 );
or \U$27939 ( \28316 , \24816 , RIae79d90_164);
nand \U$27940 ( \28317 , \28315 , \28316 );
not \U$27941 ( \28318 , \28317 );
or \U$27942 ( \28319 , \28312 , \28318 );
and \U$27943 ( \28320 , RIae79d90_164, \9316 );
not \U$27944 ( \28321 , RIae79d90_164);
and \U$27945 ( \28322 , \28321 , \14644 );
or \U$27946 ( \28323 , \28320 , \28322 );
nand \U$27947 ( \28324 , \5048 , \28323 );
nand \U$27948 ( \28325 , \28319 , \28324 );
xor \U$27949 ( \28326 , \28311 , \28325 );
not \U$27950 ( \28327 , \9517 );
not \U$27951 ( \28328 , \18027 );
not \U$27952 ( \28329 , \24679 );
or \U$27953 ( \28330 , \28328 , \28329 );
nand \U$27954 ( \28331 , \15128 , RIae79fe8_169);
nand \U$27955 ( \28332 , \28330 , \28331 );
not \U$27956 ( \28333 , \28332 );
or \U$27957 ( \28334 , \28327 , \28333 );
not \U$27958 ( \28335 , \9504 );
not \U$27959 ( \28336 , \21732 );
or \U$27960 ( \28337 , \28335 , \28336 );
not \U$27961 ( \28338 , \9280 );
nand \U$27962 ( \28339 , \28338 , RIae79fe8_169);
nand \U$27963 ( \28340 , \28337 , \28339 );
nand \U$27964 ( \28341 , \28340 , \11913 );
nand \U$27965 ( \28342 , \28334 , \28341 );
and \U$27966 ( \28343 , \28326 , \28342 );
and \U$27967 ( \28344 , \28311 , \28325 );
or \U$27968 ( \28345 , \28343 , \28344 );
not \U$27969 ( \28346 , \28345 );
xor \U$27970 ( \28347 , \28295 , \28346 );
not \U$27971 ( \28348 , \28347 );
or \U$27972 ( \28349 , \28238 , \28348 );
or \U$27973 ( \28350 , \28347 , \28237 );
nand \U$27974 ( \28351 , \28349 , \28350 );
not \U$27975 ( \28352 , \27618 );
not \U$27976 ( \28353 , \27607 );
or \U$27977 ( \28354 , \28352 , \28353 );
not \U$27978 ( \28355 , \27588 );
nand \U$27979 ( \28356 , \28355 , \27603 );
nand \U$27980 ( \28357 , \28354 , \28356 );
not \U$27981 ( \28358 , \28357 );
not \U$27982 ( \28359 , \1820 );
not \U$27983 ( \28360 , \2970 );
not \U$27984 ( \28361 , \10338 );
or \U$27985 ( \28362 , \28360 , \28361 );
or \U$27986 ( \28363 , \10856 , \21474 );
nand \U$27987 ( \28364 , \28362 , \28363 );
not \U$27988 ( \28365 , \28364 );
or \U$27989 ( \28366 , \28359 , \28365 );
nand \U$27990 ( \28367 , \27594 , \1843 );
nand \U$27991 ( \28368 , \28366 , \28367 );
not \U$27992 ( \28369 , \28368 );
not \U$27993 ( \28370 , \1863 );
not \U$27994 ( \28371 , RIae793b8_143);
not \U$27995 ( \28372 , \10259 );
or \U$27996 ( \28373 , \28371 , \28372 );
or \U$27997 ( \28374 , \10259 , RIae793b8_143);
nand \U$27998 ( \28375 , \28373 , \28374 );
not \U$27999 ( \28376 , \28375 );
or \U$28000 ( \28377 , \28370 , \28376 );
nand \U$28001 ( \28378 , \28245 , \1909 );
nand \U$28002 ( \28379 , \28377 , \28378 );
not \U$28003 ( \28380 , \28379 );
not \U$28004 ( \28381 , RIae79250_140);
not \U$28005 ( \28382 , \16006 );
or \U$28006 ( \28383 , \28381 , \28382 );
or \U$28007 ( \28384 , \16006 , RIae79250_140);
nand \U$28008 ( \28385 , \28383 , \28384 );
not \U$28009 ( \28386 , \28385 );
or \U$28010 ( \28387 , \28386 , \1502 );
and \U$28011 ( \28388 , RIae79250_140, \17971 );
not \U$28012 ( \28389 , RIae79250_140);
and \U$28013 ( \28390 , \28389 , \12857 );
nor \U$28014 ( \28391 , \28388 , \28390 );
or \U$28015 ( \28392 , \28391 , \1496 );
nand \U$28016 ( \28393 , \28387 , \28392 );
not \U$28017 ( \28394 , \28393 );
or \U$28018 ( \28395 , RIae79340_142, RIae793b8_143);
nand \U$28019 ( \28396 , \28395 , \12857 );
nand \U$28020 ( \28397 , \28396 , \1435 );
not \U$28021 ( \28398 , \28397 );
and \U$28022 ( \28399 , \28394 , \28398 );
and \U$28023 ( \28400 , \28393 , \28397 );
nor \U$28024 ( \28401 , \28399 , \28400 );
not \U$28025 ( \28402 , \28401 );
and \U$28026 ( \28403 , \28380 , \28402 );
and \U$28027 ( \28404 , \28379 , \28401 );
nor \U$28028 ( \28405 , \28403 , \28404 );
not \U$28029 ( \28406 , \28405 );
and \U$28030 ( \28407 , \28369 , \28406 );
and \U$28031 ( \28408 , \28368 , \28405 );
nor \U$28032 ( \28409 , \28407 , \28408 );
not \U$28033 ( \28410 , \28409 );
or \U$28034 ( \28411 , \28358 , \28410 );
or \U$28035 ( \28412 , \28357 , \28409 );
nand \U$28036 ( \28413 , \28411 , \28412 );
not \U$28037 ( \28414 , \5048 );
not \U$28038 ( \28415 , RIae79d90_164);
not \U$28039 ( \28416 , \9299 );
or \U$28040 ( \28417 , \28415 , \28416 );
or \U$28041 ( \28418 , \17245 , RIae79d90_164);
nand \U$28042 ( \28419 , \28417 , \28418 );
not \U$28043 ( \28420 , \28419 );
or \U$28044 ( \28421 , \28414 , \28420 );
nand \U$28045 ( \28422 , \28323 , \5039 );
nand \U$28046 ( \28423 , \28421 , \28422 );
not \U$28047 ( \28424 , \28423 );
and \U$28048 ( \28425 , \28413 , \28424 );
not \U$28049 ( \28426 , \28413 );
and \U$28050 ( \28427 , \28426 , \28423 );
nor \U$28051 ( \28428 , \28425 , \28427 );
or \U$28052 ( \28429 , \27868 , \27878 );
nand \U$28053 ( \28430 , \28429 , \27893 );
nand \U$28054 ( \28431 , \27878 , \27868 );
nand \U$28055 ( \28432 , \28430 , \28431 );
xor \U$28056 ( \28433 , \28428 , \28432 );
not \U$28057 ( \28434 , \27623 );
nand \U$28058 ( \28435 , \28434 , \27638 );
not \U$28059 ( \28436 , \28435 );
not \U$28060 ( \28437 , \27662 );
or \U$28061 ( \28438 , \28436 , \28437 );
not \U$28062 ( \28439 , \27638 );
nand \U$28063 ( \28440 , \28439 , \27623 );
nand \U$28064 ( \28441 , \28438 , \28440 );
xnor \U$28065 ( \28442 , \28433 , \28441 );
xor \U$28066 ( \28443 , \28351 , \28442 );
not \U$28067 ( \28444 , \2007 );
not \U$28068 ( \28445 , \2521 );
not \U$28069 ( \28446 , \12482 );
or \U$28070 ( \28447 , \28445 , \28446 );
or \U$28071 ( \28448 , \9607 , \2521 );
nand \U$28072 ( \28449 , \28447 , \28448 );
not \U$28073 ( \28450 , \28449 );
or \U$28074 ( \28451 , \28444 , \28450 );
nand \U$28075 ( \28452 , \28289 , \1988 );
nand \U$28076 ( \28453 , \28451 , \28452 );
not \U$28077 ( \28454 , \2450 );
not \U$28078 ( \28455 , \2442 );
not \U$28079 ( \28456 , \12600 );
or \U$28080 ( \28457 , \28455 , \28456 );
or \U$28081 ( \28458 , \9395 , \2447 );
nand \U$28082 ( \28459 , \28457 , \28458 );
not \U$28083 ( \28460 , \28459 );
or \U$28084 ( \28461 , \28454 , \28460 );
nand \U$28085 ( \28462 , \28215 , \2431 );
nand \U$28086 ( \28463 , \28461 , \28462 );
xor \U$28087 ( \28464 , \28453 , \28463 );
not \U$28088 ( \28465 , \28464 );
not \U$28089 ( \28466 , \2776 );
and \U$28090 ( \28467 , RIae79c28_161, \12615 );
not \U$28091 ( \28468 , RIae79c28_161);
and \U$28092 ( \28469 , \28468 , \12614 );
or \U$28093 ( \28470 , \28467 , \28469 );
not \U$28094 ( \28471 , \28470 );
or \U$28095 ( \28472 , \28466 , \28471 );
nand \U$28096 ( \28473 , \28230 , \2767 );
nand \U$28097 ( \28474 , \28472 , \28473 );
not \U$28098 ( \28475 , \28474 );
not \U$28099 ( \28476 , \28475 );
and \U$28100 ( \28477 , \28465 , \28476 );
and \U$28101 ( \28478 , \28464 , \28475 );
nor \U$28102 ( \28479 , \28477 , \28478 );
or \U$28103 ( \28480 , \27567 , \27539 );
nand \U$28104 ( \28481 , \28480 , \27552 );
nand \U$28105 ( \28482 , \27567 , \27539 );
nand \U$28106 ( \28483 , \28481 , \28482 );
xor \U$28107 ( \28484 , \28479 , \28483 );
not \U$28108 ( \28485 , \10573 );
and \U$28109 ( \28486 , RIae79ef8_167, \13976 );
not \U$28110 ( \28487 , RIae79ef8_167);
and \U$28111 ( \28488 , \28487 , \5722 );
or \U$28112 ( \28489 , \28486 , \28488 );
not \U$28113 ( \28490 , \28489 );
or \U$28114 ( \28491 , \28485 , \28490 );
nand \U$28115 ( \28492 , \28309 , \19362 );
nand \U$28116 ( \28493 , \28491 , \28492 );
not \U$28117 ( \28494 , \9814 );
not \U$28118 ( \28495 , \11054 );
not \U$28119 ( \28496 , \4982 );
or \U$28120 ( \28497 , \28495 , \28496 );
or \U$28121 ( \28498 , \17338 , \9799 );
nand \U$28122 ( \28499 , \28497 , \28498 );
not \U$28123 ( \28500 , \28499 );
or \U$28124 ( \28501 , \28494 , \28500 );
nand \U$28125 ( \28502 , \28200 , \9792 );
nand \U$28126 ( \28503 , \28501 , \28502 );
xor \U$28127 ( \28504 , \28493 , \28503 );
not \U$28128 ( \28505 , \10700 );
not \U$28129 ( \28506 , RIae79fe8_169);
not \U$28130 ( \28507 , \4960 );
or \U$28131 ( \28508 , \28506 , \28507 );
or \U$28132 ( \28509 , \10829 , RIae79fe8_169);
nand \U$28133 ( \28510 , \28508 , \28509 );
not \U$28134 ( \28511 , \28510 );
or \U$28135 ( \28512 , \28505 , \28511 );
nand \U$28136 ( \28513 , \28332 , \11914 );
nand \U$28137 ( \28514 , \28512 , \28513 );
xor \U$28138 ( \28515 , \28504 , \28514 );
xor \U$28139 ( \28516 , \28484 , \28515 );
and \U$28140 ( \28517 , \28443 , \28516 );
and \U$28141 ( \28518 , \28351 , \28442 );
or \U$28142 ( \28519 , \28517 , \28518 );
not \U$28143 ( \28520 , \28519 );
not \U$28144 ( \28521 , \28520 );
not \U$28145 ( \28522 , \2007 );
xor \U$28146 ( \28523 , \15947 , RIae797f0_152);
not \U$28147 ( \28524 , \28523 );
or \U$28148 ( \28525 , \28522 , \28524 );
nand \U$28149 ( \28526 , \28449 , \1988 );
nand \U$28150 ( \28527 , \28525 , \28526 );
not \U$28151 ( \28528 , \28527 );
not \U$28152 ( \28529 , \2431 );
not \U$28153 ( \28530 , \28459 );
or \U$28154 ( \28531 , \28529 , \28530 );
xor \U$28155 ( \28532 , \9455 , RIae79778_151);
nand \U$28156 ( \28533 , \28532 , \2450 );
nand \U$28157 ( \28534 , \28531 , \28533 );
not \U$28158 ( \28535 , \28534 );
not \U$28159 ( \28536 , \28535 );
or \U$28160 ( \28537 , \28528 , \28536 );
not \U$28161 ( \28538 , \28527 );
nand \U$28162 ( \28539 , \28538 , \28534 );
nand \U$28163 ( \28540 , \28537 , \28539 );
not \U$28164 ( \28541 , \28540 );
not \U$28165 ( \28542 , \9792 );
not \U$28166 ( \28543 , \28499 );
or \U$28167 ( \28544 , \28542 , \28543 );
not \U$28168 ( \28545 , \11054 );
not \U$28169 ( \28546 , \5673 );
or \U$28170 ( \28547 , \28545 , \28546 );
nand \U$28171 ( \28548 , \3270 , RIae7a2b8_175);
nand \U$28172 ( \28549 , \28547 , \28548 );
nand \U$28173 ( \28550 , \28549 , \9814 );
nand \U$28174 ( \28551 , \28544 , \28550 );
not \U$28175 ( \28552 , \28551 );
not \U$28176 ( \28553 , \28552 );
and \U$28177 ( \28554 , \28541 , \28553 );
and \U$28178 ( \28555 , \28552 , \28540 );
nor \U$28179 ( \28556 , \28554 , \28555 );
not \U$28180 ( \28557 , \6091 );
not \U$28181 ( \28558 , \28419 );
or \U$28182 ( \28559 , \28557 , \28558 );
not \U$28183 ( \28560 , RIae79d90_164);
not \U$28184 ( \28561 , \15117 );
or \U$28185 ( \28562 , \28560 , \28561 );
or \U$28186 ( \28563 , \10406 , RIae79d90_164);
nand \U$28187 ( \28564 , \28562 , \28563 );
nand \U$28188 ( \28565 , \28564 , \5048 );
nand \U$28189 ( \28566 , \28559 , \28565 );
not \U$28190 ( \28567 , \10573 );
not \U$28191 ( \28568 , RIae79ef8_167);
not \U$28192 ( \28569 , \6257 );
or \U$28193 ( \28570 , \28568 , \28569 );
or \U$28194 ( \28571 , \15128 , RIae79ef8_167);
nand \U$28195 ( \28572 , \28570 , \28571 );
not \U$28196 ( \28573 , \28572 );
or \U$28197 ( \28574 , \28567 , \28573 );
nand \U$28198 ( \28575 , \28489 , \19362 );
nand \U$28199 ( \28576 , \28574 , \28575 );
xor \U$28200 ( \28577 , \28566 , \28576 );
not \U$28201 ( \28578 , \9517 );
and \U$28202 ( \28579 , RIae79fe8_169, \6238 );
not \U$28203 ( \28580 , RIae79fe8_169);
and \U$28204 ( \28581 , \28580 , \4169 );
or \U$28205 ( \28582 , \28579 , \28581 );
not \U$28206 ( \28583 , \28582 );
or \U$28207 ( \28584 , \28578 , \28583 );
nand \U$28208 ( \28585 , \28510 , \11913 );
nand \U$28209 ( \28586 , \28584 , \28585 );
xor \U$28210 ( \28587 , \28577 , \28586 );
xor \U$28211 ( \28588 , \28556 , \28587 );
not \U$28212 ( \28589 , \9473 );
not \U$28213 ( \28590 , \27650 );
or \U$28214 ( \28591 , \28589 , \28590 );
not \U$28215 ( \28592 , RIae7a6f0_184);
not \U$28216 ( \28593 , \9797 );
or \U$28217 ( \28594 , \28592 , \28593 );
or \U$28218 ( \28595 , \3051 , RIae7a6f0_184);
nand \U$28219 ( \28596 , \28594 , \28595 );
nand \U$28220 ( \28597 , \28596 , \9705 );
nand \U$28221 ( \28598 , \28591 , \28597 );
not \U$28222 ( \28599 , \28598 );
or \U$28223 ( \28600 , \28271 , \28251 );
nand \U$28224 ( \28601 , \28600 , \28253 );
not \U$28225 ( \28602 , \28601 );
not \U$28226 ( \28603 , \2011 );
and \U$28227 ( \28604 , RIae79610_148, \16036 );
not \U$28228 ( \28605 , RIae79610_148);
and \U$28229 ( \28606 , \28605 , \11576 );
or \U$28230 ( \28607 , \28604 , \28606 );
not \U$28231 ( \28608 , \28607 );
or \U$28232 ( \28609 , \28603 , \28608 );
not \U$28233 ( \28610 , \28261 );
nand \U$28234 ( \28611 , \28610 , \2063 );
nand \U$28235 ( \28612 , \28609 , \28611 );
not \U$28236 ( \28613 , \28612 );
not \U$28237 ( \28614 , \28613 );
and \U$28238 ( \28615 , \28602 , \28614 );
and \U$28239 ( \28616 , \28601 , \28613 );
nor \U$28240 ( \28617 , \28615 , \28616 );
not \U$28241 ( \28618 , \2321 );
not \U$28242 ( \28619 , RIae798e0_154);
not \U$28243 ( \28620 , \10724 );
or \U$28244 ( \28621 , \28619 , \28620 );
or \U$28245 ( \28622 , \19015 , RIae798e0_154);
nand \U$28246 ( \28623 , \28621 , \28622 );
not \U$28247 ( \28624 , \28623 );
or \U$28248 ( \28625 , \28618 , \28624 );
not \U$28249 ( \28626 , RIae798e0_154);
not \U$28250 ( \28627 , \11387 );
or \U$28251 ( \28628 , \28626 , \28627 );
or \U$28252 ( \28629 , \10084 , RIae798e0_154);
nand \U$28253 ( \28630 , \28628 , \28629 );
nand \U$28254 ( \28631 , \28630 , \2339 );
nand \U$28255 ( \28632 , \28625 , \28631 );
xnor \U$28256 ( \28633 , \28617 , \28632 );
not \U$28257 ( \28634 , \28633 );
not \U$28258 ( \28635 , \10696 );
not \U$28259 ( \28636 , \27636 );
or \U$28260 ( \28637 , \28635 , \28636 );
and \U$28261 ( \28638 , RIae7a498_179, \3529 );
not \U$28262 ( \28639 , RIae7a498_179);
and \U$28263 ( \28640 , \28639 , \3524 );
nor \U$28264 ( \28641 , \28638 , \28640 );
nand \U$28265 ( \28642 , \28641 , \10676 );
nand \U$28266 ( \28643 , \28637 , \28642 );
not \U$28267 ( \28644 , \28643 );
not \U$28268 ( \28645 , \28644 );
or \U$28269 ( \28646 , \28634 , \28645 );
or \U$28270 ( \28647 , \28644 , \28633 );
nand \U$28271 ( \28648 , \28646 , \28647 );
not \U$28272 ( \28649 , \28648 );
or \U$28273 ( \28650 , \28599 , \28649 );
not \U$28274 ( \28651 , \28644 );
nand \U$28275 ( \28652 , \28651 , \28633 );
nand \U$28276 ( \28653 , \28650 , \28652 );
not \U$28277 ( \28654 , \28653 );
xnor \U$28278 ( \28655 , \28588 , \28654 );
not \U$28279 ( \28656 , \28144 );
not \U$28280 ( \28657 , \28177 );
or \U$28281 ( \28658 , \28656 , \28657 );
not \U$28282 ( \28659 , \28143 );
not \U$28283 ( \28660 , \28176 );
or \U$28284 ( \28661 , \28659 , \28660 );
nand \U$28285 ( \28662 , \28661 , \28100 );
nand \U$28286 ( \28663 , \28658 , \28662 );
xor \U$28287 ( \28664 , \28655 , \28663 );
not \U$28288 ( \28665 , \28483 );
not \U$28289 ( \28666 , \28479 );
not \U$28290 ( \28667 , \28515 );
or \U$28291 ( \28668 , \28666 , \28667 );
or \U$28292 ( \28669 , \28515 , \28479 );
nand \U$28293 ( \28670 , \28668 , \28669 );
not \U$28294 ( \28671 , \28670 );
or \U$28295 ( \28672 , \28665 , \28671 );
not \U$28296 ( \28673 , \28479 );
nand \U$28297 ( \28674 , \28673 , \28515 );
nand \U$28298 ( \28675 , \28672 , \28674 );
xor \U$28299 ( \28676 , \28664 , \28675 );
not \U$28300 ( \28677 , \28676 );
or \U$28301 ( \28678 , \28521 , \28677 );
or \U$28302 ( \28679 , \28676 , \28520 );
nand \U$28303 ( \28680 , \28678 , \28679 );
not \U$28304 ( \28681 , \28680 );
or \U$28305 ( \28682 , \28186 , \28681 );
nand \U$28306 ( \28683 , \28519 , \28676 );
nand \U$28307 ( \28684 , \28682 , \28683 );
not \U$28308 ( \28685 , \28684 );
not \U$28309 ( \28686 , \28685 );
not \U$28310 ( \28687 , \28655 );
not \U$28311 ( \28688 , \28663 );
not \U$28312 ( \28689 , \28688 );
or \U$28313 ( \28690 , \28687 , \28689 );
nand \U$28314 ( \28691 , \28690 , \28675 );
not \U$28315 ( \28692 , \28655 );
nand \U$28316 ( \28693 , \28692 , \28663 );
nand \U$28317 ( \28694 , \28691 , \28693 );
nand \U$28318 ( \28695 , \28150 , \14510 );
not \U$28319 ( \28696 , \17067 );
xor \U$28320 ( \28697 , RIae7a8d0_188, \28696 );
nand \U$28321 ( \28698 , \28697 , \10275 );
nand \U$28322 ( \28699 , \28695 , \28698 );
not \U$28323 ( \28700 , \19466 );
not \U$28324 ( \28701 , \28077 );
or \U$28325 ( \28702 , \28700 , \28701 );
and \U$28326 ( \28703 , RIae7a240_174, \17052 );
not \U$28327 ( \28704 , RIae7a240_174);
and \U$28328 ( \28705 , \28704 , \9671 );
nor \U$28329 ( \28706 , \28703 , \28705 );
nand \U$28330 ( \28707 , \28706 , \9699 );
nand \U$28331 ( \28708 , \28702 , \28707 );
and \U$28332 ( \28709 , \28699 , \28708 );
not \U$28333 ( \28710 , \28699 );
not \U$28334 ( \28711 , \28708 );
and \U$28335 ( \28712 , \28710 , \28711 );
nor \U$28336 ( \28713 , \28709 , \28712 );
not \U$28337 ( \28714 , \9745 );
not \U$28338 ( \28715 , RIae7a060_170);
not \U$28339 ( \28716 , \2153 );
or \U$28340 ( \28717 , \28715 , \28716 );
or \U$28341 ( \28718 , \14712 , RIae7a060_170);
nand \U$28342 ( \28719 , \28717 , \28718 );
not \U$28343 ( \28720 , \28719 );
or \U$28344 ( \28721 , \28714 , \28720 );
nand \U$28345 ( \28722 , \28162 , \9730 );
nand \U$28346 ( \28723 , \28721 , \28722 );
xor \U$28347 ( \28724 , \28713 , \28723 );
not \U$28348 ( \28725 , \9473 );
not \U$28349 ( \28726 , \28596 );
or \U$28350 ( \28727 , \28725 , \28726 );
not \U$28351 ( \28728 , \16101 );
not \U$28352 ( \28729 , \1897 );
or \U$28353 ( \28730 , \28728 , \28729 );
not \U$28354 ( \28731 , RIae7a6f0_184);
or \U$28355 ( \28732 , \1898 , \28731 );
nand \U$28356 ( \28733 , \28730 , \28732 );
nand \U$28357 ( \28734 , \28733 , \9478 );
nand \U$28358 ( \28735 , \28727 , \28734 );
not \U$28359 ( \28736 , \28735 );
not \U$28360 ( \28737 , \2011 );
and \U$28361 ( \28738 , RIae79610_148, \16909 );
not \U$28362 ( \28739 , RIae79610_148);
and \U$28363 ( \28740 , \28739 , \10042 );
or \U$28364 ( \28741 , \28738 , \28740 );
not \U$28365 ( \28742 , \28741 );
or \U$28366 ( \28743 , \28737 , \28742 );
nand \U$28367 ( \28744 , \28607 , \2063 );
nand \U$28368 ( \28745 , \28743 , \28744 );
not \U$28369 ( \28746 , \28397 );
nand \U$28370 ( \28747 , \28746 , \28393 );
xor \U$28371 ( \28748 , \28745 , \28747 );
not \U$28372 ( \28749 , \1843 );
not \U$28373 ( \28750 , \28364 );
or \U$28374 ( \28751 , \28749 , \28750 );
and \U$28375 ( \28752 , RIae79688_149, \10149 );
not \U$28376 ( \28753 , RIae79688_149);
and \U$28377 ( \28754 , \28753 , \10142 );
or \U$28378 ( \28755 , \28752 , \28754 );
nand \U$28379 ( \28756 , \28755 , \1820 );
nand \U$28380 ( \28757 , \28751 , \28756 );
xor \U$28381 ( \28758 , \28748 , \28757 );
not \U$28382 ( \28759 , \28758 );
not \U$28383 ( \28760 , \10667 );
not \U$28384 ( \28761 , \28171 );
or \U$28385 ( \28762 , \28760 , \28761 );
not \U$28386 ( \28763 , RIae7a150_172);
not \U$28387 ( \28764 , \2285 );
or \U$28388 ( \28765 , \28763 , \28764 );
nand \U$28389 ( \28766 , \3747 , \10672 );
nand \U$28390 ( \28767 , \28765 , \28766 );
nand \U$28391 ( \28768 , \28767 , \9776 );
nand \U$28392 ( \28769 , \28762 , \28768 );
not \U$28393 ( \28770 , \28769 );
or \U$28394 ( \28771 , \28759 , \28770 );
or \U$28395 ( \28772 , \28769 , \28758 );
nand \U$28396 ( \28773 , \28771 , \28772 );
not \U$28397 ( \28774 , \28773 );
not \U$28398 ( \28775 , \28774 );
and \U$28399 ( \28776 , \28736 , \28775 );
and \U$28400 ( \28777 , \28735 , \28774 );
nor \U$28401 ( \28778 , \28776 , \28777 );
xor \U$28402 ( \28779 , \28724 , \28778 );
not \U$28403 ( \28780 , \9644 );
not \U$28404 ( \28781 , \28084 );
or \U$28405 ( \28782 , \28780 , \28781 );
xor \U$28406 ( \28783 , RIae7a3a8_177, \2093 );
nand \U$28407 ( \28784 , \28783 , \9622 );
nand \U$28408 ( \28785 , \28782 , \28784 );
not \U$28409 ( \28786 , \10631 );
not \U$28410 ( \28787 , RIae7a510_180);
not \U$28411 ( \28788 , \11681 );
or \U$28412 ( \28789 , \28787 , \28788 );
not \U$28413 ( \28790 , \10583 );
or \U$28414 ( \28791 , \28790 , RIae7a510_180);
nand \U$28415 ( \28792 , \28789 , \28791 );
not \U$28416 ( \28793 , \28792 );
or \U$28417 ( \28794 , \28786 , \28793 );
nand \U$28418 ( \28795 , \28114 , \10637 );
nand \U$28419 ( \28796 , \28794 , \28795 );
xor \U$28420 ( \28797 , \28785 , \28796 );
not \U$28421 ( \28798 , \9527 );
not \U$28422 ( \28799 , \9529 );
not \U$28423 ( \28800 , \11885 );
or \U$28424 ( \28801 , \28799 , \28800 );
or \U$28425 ( \28802 , \11888 , \17112 );
nand \U$28426 ( \28803 , \28801 , \28802 );
not \U$28427 ( \28804 , \28803 );
or \U$28428 ( \28805 , \28798 , \28804 );
nand \U$28429 ( \28806 , \28095 , \11851 );
nand \U$28430 ( \28807 , \28805 , \28806 );
xor \U$28431 ( \28808 , \28797 , \28807 );
xor \U$28432 ( \28809 , \28779 , \28808 );
not \U$28433 ( \28810 , \28809 );
not \U$28434 ( \28811 , \28810 );
and \U$28435 ( \28812 , \2101 , RIae7aa38_191);
nor \U$28436 ( \28813 , \2849 , RIae7aa38_191);
nor \U$28437 ( \28814 , \28812 , \28813 );
or \U$28438 ( \28815 , \28814 , \14666 );
nand \U$28439 ( \28816 , \28136 , \16383 );
nand \U$28440 ( \28817 , \28815 , \28816 );
not \U$28441 ( \28818 , \28817 );
nand \U$28442 ( \28819 , \28103 , \11761 );
not \U$28443 ( \28820 , RIae79ca0_162);
not \U$28444 ( \28821 , \9316 );
or \U$28445 ( \28822 , \28820 , \28821 );
nand \U$28446 ( \28823 , \16274 , \4844 );
nand \U$28447 ( \28824 , \28822 , \28823 );
nand \U$28448 ( \28825 , \28824 , \4853 );
and \U$28449 ( \28826 , \28819 , \28825 );
not \U$28450 ( \28827 , \28405 );
not \U$28451 ( \28828 , \28827 );
not \U$28452 ( \28829 , \28368 );
or \U$28453 ( \28830 , \28828 , \28829 );
not \U$28454 ( \28831 , \28401 );
nand \U$28455 ( \28832 , \28831 , \28379 );
nand \U$28456 ( \28833 , \28830 , \28832 );
xnor \U$28457 ( \28834 , \28826 , \28833 );
xor \U$28458 ( \28835 , \28818 , \28834 );
not \U$28459 ( \28836 , \28164 );
not \U$28460 ( \28837 , \28175 );
or \U$28461 ( \28838 , \28836 , \28837 );
or \U$28462 ( \28839 , \28175 , \28164 );
nand \U$28463 ( \28840 , \28839 , \28154 );
nand \U$28464 ( \28841 , \28838 , \28840 );
xnor \U$28465 ( \28842 , \28835 , \28841 );
not \U$28466 ( \28843 , \28088 );
not \U$28467 ( \28844 , \28082 );
not \U$28468 ( \28845 , \28844 );
not \U$28469 ( \28846 , \28099 );
or \U$28470 ( \28847 , \28845 , \28846 );
or \U$28471 ( \28848 , \28099 , \28844 );
nand \U$28472 ( \28849 , \28847 , \28848 );
not \U$28473 ( \28850 , \28849 );
or \U$28474 ( \28851 , \28843 , \28850 );
nand \U$28475 ( \28852 , \28099 , \28082 );
nand \U$28476 ( \28853 , \28851 , \28852 );
xnor \U$28477 ( \28854 , \28842 , \28853 );
not \U$28478 ( \28855 , \28854 );
not \U$28479 ( \28856 , \28855 );
or \U$28480 ( \28857 , \28811 , \28856 );
not \U$28481 ( \28858 , \28809 );
not \U$28482 ( \28859 , \28854 );
or \U$28483 ( \28860 , \28858 , \28859 );
xor \U$28484 ( \28861 , \28648 , \28598 );
not \U$28485 ( \28862 , \28047 );
not \U$28486 ( \28863 , \28029 );
not \U$28487 ( \28864 , \28863 );
or \U$28488 ( \28865 , \28862 , \28864 );
nand \U$28489 ( \28866 , \28046 , \28036 );
nand \U$28490 ( \28867 , \28865 , \28866 );
xor \U$28491 ( \28868 , \27686 , \27697 );
and \U$28492 ( \28869 , \28868 , \27712 );
and \U$28493 ( \28870 , \27686 , \27697 );
or \U$28494 ( \28871 , \28869 , \28870 );
nor \U$28495 ( \28872 , \28867 , \28871 );
not \U$28496 ( \28873 , \28872 );
not \U$28497 ( \28874 , \28873 );
not \U$28498 ( \28875 , \9517 );
not \U$28499 ( \28876 , \28340 );
or \U$28500 ( \28877 , \28875 , \28876 );
nand \U$28501 ( \28878 , \27726 , \11913 );
nand \U$28502 ( \28879 , \28877 , \28878 );
not \U$28503 ( \28880 , \28879 );
not \U$28504 ( \28881 , \27573 );
not \U$28505 ( \28882 , \27587 );
or \U$28506 ( \28883 , \28881 , \28882 );
or \U$28507 ( \28884 , \27587 , \27573 );
nand \U$28508 ( \28885 , \28883 , \28884 );
not \U$28509 ( \28886 , \2011 );
not \U$28510 ( \28887 , \28269 );
not \U$28511 ( \28888 , \28887 );
or \U$28512 ( \28889 , \28886 , \28888 );
nand \U$28513 ( \28890 , \27970 , \2063 );
nand \U$28514 ( \28891 , \28889 , \28890 );
xor \U$28515 ( \28892 , \28885 , \28891 );
not \U$28516 ( \28893 , \1843 );
not \U$28517 ( \28894 , \27986 );
not \U$28518 ( \28895 , \28894 );
or \U$28519 ( \28896 , \28893 , \28895 );
nand \U$28520 ( \28897 , \27601 , \1820 );
nand \U$28521 ( \28898 , \28896 , \28897 );
xor \U$28522 ( \28899 , \28892 , \28898 );
not \U$28523 ( \28900 , \28899 );
not \U$28524 ( \28901 , \2418 );
not \U$28525 ( \28902 , \28223 );
or \U$28526 ( \28903 , \28901 , \28902 );
not \U$28527 ( \28904 , RIae79c28_161);
not \U$28528 ( \28905 , \15944 );
or \U$28529 ( \28906 , \28904 , \28905 );
or \U$28530 ( \28907 , \15944 , RIae79c28_161);
nand \U$28531 ( \28908 , \28906 , \28907 );
nand \U$28532 ( \28909 , \28908 , \2417 );
nand \U$28533 ( \28910 , \28903 , \28909 );
not \U$28534 ( \28911 , \28910 );
not \U$28535 ( \28912 , \28911 );
or \U$28536 ( \28913 , \28900 , \28912 );
not \U$28537 ( \28914 , \28899 );
nand \U$28538 ( \28915 , \28914 , \28910 );
nand \U$28539 ( \28916 , \28913 , \28915 );
not \U$28540 ( \28917 , \28916 );
or \U$28541 ( \28918 , \28880 , \28917 );
nand \U$28542 ( \28919 , \28910 , \28899 );
nand \U$28543 ( \28920 , \28918 , \28919 );
not \U$28544 ( \28921 , \28920 );
or \U$28545 ( \28922 , \28874 , \28921 );
nand \U$28546 ( \28923 , \28867 , \28871 );
nand \U$28547 ( \28924 , \28922 , \28923 );
nor \U$28548 ( \28925 , \28861 , \28924 );
not \U$28549 ( \28926 , \28925 );
not \U$28550 ( \28927 , \28926 );
nand \U$28551 ( \28928 , \28294 , \28283 );
xor \U$28552 ( \28929 , \28928 , \28291 );
not \U$28553 ( \28930 , \2339 );
not \U$28554 ( \28931 , \27688 );
or \U$28555 ( \28932 , \28930 , \28931 );
nand \U$28556 ( \28933 , \28630 , \2322 );
nand \U$28557 ( \28934 , \28932 , \28933 );
not \U$28558 ( \28935 , \9828 );
not \U$28559 ( \28936 , \27703 );
or \U$28560 ( \28937 , \28935 , \28936 );
xor \U$28561 ( \28938 , \17185 , RIae794a8_145);
nand \U$28562 ( \28939 , \28938 , \1919 );
nand \U$28563 ( \28940 , \28937 , \28939 );
xor \U$28564 ( \28941 , \28934 , \28940 );
not \U$28565 ( \28942 , \13720 );
not \U$28566 ( \28943 , RIae7a240_174);
not \U$28567 ( \28944 , \22961 );
or \U$28568 ( \28945 , \28943 , \28944 );
nand \U$28569 ( \28946 , \3208 , \11114 );
nand \U$28570 ( \28947 , \28945 , \28946 );
not \U$28571 ( \28948 , \28947 );
or \U$28572 ( \28949 , \28942 , \28948 );
nand \U$28573 ( \28950 , \28080 , \13121 );
nand \U$28574 ( \28951 , \28949 , \28950 );
xor \U$28575 ( \28952 , \28941 , \28951 );
xor \U$28576 ( \28953 , \28929 , \28952 );
not \U$28577 ( \28954 , \10573 );
not \U$28578 ( \28955 , \28300 );
or \U$28579 ( \28956 , \28954 , \28955 );
nand \U$28580 ( \28957 , \27740 , \15989 );
nand \U$28581 ( \28958 , \28956 , \28957 );
not \U$28582 ( \28959 , \28958 );
not \U$28583 ( \28960 , \14940 );
not \U$28584 ( \28961 , \28317 );
or \U$28585 ( \28962 , \28960 , \28961 );
not \U$28586 ( \28963 , \4968 );
not \U$28587 ( \28964 , \14691 );
or \U$28588 ( \28965 , \28963 , \28964 );
or \U$28589 ( \28966 , \14691 , \4968 );
nand \U$28590 ( \28967 , \28965 , \28966 );
nand \U$28591 ( \28968 , \28967 , \6091 );
nand \U$28592 ( \28969 , \28962 , \28968 );
not \U$28593 ( \28970 , \27772 );
nand \U$28594 ( \28971 , \28970 , \27767 );
not \U$28595 ( \28972 , \28971 );
not \U$28596 ( \28973 , \2249 );
not \U$28597 ( \28974 , \28044 );
or \U$28598 ( \28975 , \28973 , \28974 );
not \U$28599 ( \28976 , \10419 );
not \U$28600 ( \28977 , \10193 );
or \U$28601 ( \28978 , \28976 , \28977 );
nand \U$28602 ( \28979 , \19689 , RIae79ac0_158);
nand \U$28603 ( \28980 , \28978 , \28979 );
nand \U$28604 ( \28981 , \28980 , \2272 );
nand \U$28605 ( \28982 , \28975 , \28981 );
not \U$28606 ( \28983 , \28982 );
or \U$28607 ( \28984 , \28972 , \28983 );
or \U$28608 ( \28985 , \28982 , \28971 );
nand \U$28609 ( \28986 , \28984 , \28985 );
not \U$28610 ( \28987 , \28986 );
not \U$28611 ( \28988 , \2188 );
not \U$28612 ( \28989 , \27783 );
or \U$28613 ( \28990 , \28988 , \28989 );
nand \U$28614 ( \28991 , \27684 , \2162 );
nand \U$28615 ( \28992 , \28990 , \28991 );
not \U$28616 ( \28993 , \28992 );
or \U$28617 ( \28994 , \28987 , \28993 );
not \U$28618 ( \28995 , \28971 );
nand \U$28619 ( \28996 , \28995 , \28982 );
nand \U$28620 ( \28997 , \28994 , \28996 );
xor \U$28621 ( \28998 , \28969 , \28997 );
not \U$28622 ( \28999 , \28998 );
or \U$28623 ( \29000 , \28959 , \28999 );
nand \U$28624 ( \29001 , \28969 , \28997 );
nand \U$28625 ( \29002 , \29000 , \29001 );
and \U$28626 ( \29003 , \28953 , \29002 );
and \U$28627 ( \29004 , \28929 , \28952 );
or \U$28628 ( \29005 , \29003 , \29004 );
not \U$28629 ( \29006 , \29005 );
or \U$28630 ( \29007 , \28927 , \29006 );
nand \U$28631 ( \29008 , \28861 , \28924 );
nand \U$28632 ( \29009 , \29007 , \29008 );
nand \U$28633 ( \29010 , \28860 , \29009 );
nand \U$28634 ( \29011 , \28857 , \29010 );
xor \U$28635 ( \29012 , \28694 , \29011 );
not \U$28636 ( \29013 , \28808 );
nand \U$28637 ( \29014 , \29013 , \28778 );
not \U$28638 ( \29015 , \29014 );
not \U$28639 ( \29016 , \28724 );
or \U$28640 ( \29017 , \29015 , \29016 );
not \U$28641 ( \29018 , \28778 );
nand \U$28642 ( \29019 , \29018 , \28808 );
nand \U$28643 ( \29020 , \29017 , \29019 );
not \U$28644 ( \29021 , \29020 );
not \U$28645 ( \29022 , \29021 );
buf \U$28646 ( \29023 , \28556 );
not \U$28647 ( \29024 , \29023 );
not \U$28648 ( \29025 , \28654 );
or \U$28649 ( \29026 , \29024 , \29025 );
nand \U$28650 ( \29027 , \29026 , \28587 );
not \U$28651 ( \29028 , \29023 );
nand \U$28652 ( \29029 , \29028 , \28653 );
nand \U$28653 ( \29030 , \29027 , \29029 );
not \U$28654 ( \29031 , RIae79ef8_167);
not \U$28655 ( \29032 , \10829 );
or \U$28656 ( \29033 , \29031 , \29032 );
or \U$28657 ( \29034 , \10829 , RIae79ef8_167);
nand \U$28658 ( \29035 , \29033 , \29034 );
and \U$28659 ( \29036 , \6214 , \29035 );
and \U$28660 ( \29037 , \28572 , \11409 );
nor \U$28661 ( \29038 , \29036 , \29037 );
not \U$28662 ( \29039 , \29038 );
not \U$28663 ( \29040 , \2776 );
and \U$28664 ( \29041 , \23180 , \10584 );
not \U$28665 ( \29042 , \23180 );
and \U$28666 ( \29043 , \29042 , RIae79c28_161);
or \U$28667 ( \29044 , \29041 , \29043 );
not \U$28668 ( \29045 , \29044 );
or \U$28669 ( \29046 , \29040 , \29045 );
not \U$28670 ( \29047 , \10584 );
not \U$28671 ( \29048 , \14691 );
or \U$28672 ( \29049 , \29047 , \29048 );
not \U$28673 ( \29050 , \14691 );
nand \U$28674 ( \29051 , \29050 , RIae79c28_161);
nand \U$28675 ( \29052 , \29049 , \29051 );
nand \U$28676 ( \29053 , \29052 , \2767 );
nand \U$28677 ( \29054 , \29046 , \29053 );
not \U$28678 ( \29055 , \29054 );
not \U$28679 ( \29056 , \29055 );
not \U$28680 ( \29057 , \11913 );
not \U$28681 ( \29058 , \28582 );
or \U$28682 ( \29059 , \29057 , \29058 );
not \U$28683 ( \29060 , RIae79fe8_169);
not \U$28684 ( \29061 , \3207 );
not \U$28685 ( \29062 , \29061 );
or \U$28686 ( \29063 , \29060 , \29062 );
or \U$28687 ( \29064 , \23390 , RIae79fe8_169);
nand \U$28688 ( \29065 , \29063 , \29064 );
nand \U$28689 ( \29066 , \29065 , \9517 );
nand \U$28690 ( \29067 , \29059 , \29066 );
not \U$28691 ( \29068 , \29067 );
or \U$28692 ( \29069 , \29056 , \29068 );
or \U$28693 ( \29070 , \29067 , \29055 );
nand \U$28694 ( \29071 , \29069 , \29070 );
not \U$28695 ( \29072 , \29071 );
or \U$28696 ( \29073 , \29039 , \29072 );
or \U$28697 ( \29074 , \29071 , \29038 );
nand \U$28698 ( \29075 , \29073 , \29074 );
not \U$28699 ( \29076 , \29075 );
not \U$28700 ( \29077 , \5048 );
xor \U$28701 ( \29078 , RIae79d90_164, \5722 );
not \U$28702 ( \29079 , \29078 );
or \U$28703 ( \29080 , \29077 , \29079 );
nand \U$28704 ( \29081 , \28564 , \6091 );
nand \U$28705 ( \29082 , \29080 , \29081 );
not \U$28706 ( \29083 , \1007 );
and \U$28707 ( \29084 , RIae79160_138, \12858 );
not \U$28708 ( \29085 , RIae79160_138);
and \U$28709 ( \29086 , \29085 , \17971 );
nor \U$28710 ( \29087 , \29084 , \29086 );
not \U$28711 ( \29088 , \29087 );
or \U$28712 ( \29089 , \29083 , \29088 );
not \U$28713 ( \29090 , RIae79160_138);
not \U$28714 ( \29091 , \16005 );
or \U$28715 ( \29092 , \29090 , \29091 );
or \U$28716 ( \29093 , \12750 , RIae79160_138);
nand \U$28717 ( \29094 , \29092 , \29093 );
nand \U$28718 ( \29095 , \29094 , \1012 );
nand \U$28719 ( \29096 , \29089 , \29095 );
not \U$28720 ( \29097 , \29096 );
or \U$28721 ( \29098 , \2217 , \1004 );
or \U$28722 ( \29099 , RIae791d8_139, RIae79250_140);
nand \U$28723 ( \29100 , \29099 , \12857 );
nand \U$28724 ( \29101 , \29098 , \29100 , RIae79160_138);
not \U$28725 ( \29102 , \29101 );
and \U$28726 ( \29103 , \29097 , \29102 );
and \U$28727 ( \29104 , \29096 , \29101 );
nor \U$28728 ( \29105 , \29103 , \29104 );
not \U$28729 ( \29106 , \29105 );
not \U$28730 ( \29107 , \1501 );
xnor \U$28731 ( \29108 , \17155 , RIae79250_140);
not \U$28732 ( \29109 , \29108 );
or \U$28733 ( \29110 , \29107 , \29109 );
not \U$28734 ( \29111 , \1503 );
not \U$28735 ( \29112 , \10845 );
or \U$28736 ( \29113 , \29111 , \29112 );
nand \U$28737 ( \29114 , \28243 , RIae79250_140);
nand \U$28738 ( \29115 , \29113 , \29114 );
nand \U$28739 ( \29116 , \29115 , \1497 );
nand \U$28740 ( \29117 , \29110 , \29116 );
not \U$28741 ( \29118 , \29117 );
or \U$28742 ( \29119 , \29106 , \29118 );
or \U$28743 ( \29120 , \29117 , \29105 );
nand \U$28744 ( \29121 , \29119 , \29120 );
not \U$28745 ( \29122 , \2011 );
and \U$28746 ( \29123 , \10031 , RIae79610_148);
not \U$28747 ( \29124 , \10031 );
and \U$28748 ( \29125 , \29124 , \2053 );
nor \U$28749 ( \29126 , \29123 , \29125 );
not \U$28750 ( \29127 , \29126 );
or \U$28751 ( \29128 , \29122 , \29127 );
nand \U$28752 ( \29129 , \28741 , \2063 );
nand \U$28753 ( \29130 , \29128 , \29129 );
and \U$28754 ( \29131 , \29121 , \29130 );
not \U$28755 ( \29132 , \29121 );
not \U$28756 ( \29133 , \29130 );
and \U$28757 ( \29134 , \29132 , \29133 );
nor \U$28758 ( \29135 , \29131 , \29134 );
xor \U$28759 ( \29136 , \29082 , \29135 );
not \U$28760 ( \29137 , \29136 );
not \U$28761 ( \29138 , \4853 );
not \U$28762 ( \29139 , RIae79ca0_162);
not \U$28763 ( \29140 , \9298 );
not \U$28764 ( \29141 , \29140 );
or \U$28765 ( \29142 , \29139 , \29141 );
or \U$28766 ( \29143 , \22353 , RIae79ca0_162);
nand \U$28767 ( \29144 , \29142 , \29143 );
not \U$28768 ( \29145 , \29144 );
or \U$28769 ( \29146 , \29138 , \29145 );
nand \U$28770 ( \29147 , \28824 , \11761 );
nand \U$28771 ( \29148 , \29146 , \29147 );
not \U$28772 ( \29149 , \29148 );
not \U$28773 ( \29150 , \29149 );
and \U$28774 ( \29151 , \29137 , \29150 );
and \U$28775 ( \29152 , \29136 , \29149 );
nor \U$28776 ( \29153 , \29151 , \29152 );
not \U$28777 ( \29154 , \29153 );
not \U$28778 ( \29155 , \2322 );
and \U$28779 ( \29156 , \9607 , \2981 );
not \U$28780 ( \29157 , \9607 );
and \U$28781 ( \29158 , \29157 , RIae798e0_154);
or \U$28782 ( \29159 , \29156 , \29158 );
not \U$28783 ( \29160 , \29159 );
or \U$28784 ( \29161 , \29155 , \29160 );
not \U$28785 ( \29162 , RIae798e0_154);
not \U$28786 ( \29163 , \10461 );
or \U$28787 ( \29164 , \29162 , \29163 );
nand \U$28788 ( \29165 , \9944 , \2334 );
nand \U$28789 ( \29166 , \29164 , \29165 );
nand \U$28790 ( \29167 , \29166 , \2339 );
nand \U$28791 ( \29168 , \29161 , \29167 );
not \U$28792 ( \29169 , \15337 );
and \U$28793 ( \29170 , \9441 , RIae79778_151);
not \U$28794 ( \29171 , \9441 );
and \U$28795 ( \29172 , \29171 , \2447 );
nor \U$28796 ( \29173 , \29170 , \29172 );
not \U$28797 ( \29174 , \29173 );
or \U$28798 ( \29175 , \29169 , \29174 );
nand \U$28799 ( \29176 , \28532 , \2432 );
nand \U$28800 ( \29177 , \29175 , \29176 );
xor \U$28801 ( \29178 , \29168 , \29177 );
not \U$28802 ( \29179 , \2519 );
not \U$28803 ( \29180 , \2521 );
not \U$28804 ( \29181 , \14156 );
not \U$28805 ( \29182 , \29181 );
or \U$28806 ( \29183 , \29180 , \29182 );
nand \U$28807 ( \29184 , \9398 , RIae797f0_152);
nand \U$28808 ( \29185 , \29183 , \29184 );
not \U$28809 ( \29186 , \29185 );
or \U$28810 ( \29187 , \29179 , \29186 );
nand \U$28811 ( \29188 , \28523 , \1988 );
nand \U$28812 ( \29189 , \29187 , \29188 );
not \U$28813 ( \29190 , \29189 );
not \U$28814 ( \29191 , \29190 );
xor \U$28815 ( \29192 , \29178 , \29191 );
not \U$28816 ( \29193 , \29192 );
and \U$28817 ( \29194 , \29154 , \29193 );
and \U$28818 ( \29195 , \29153 , \29192 );
nor \U$28819 ( \29196 , \29194 , \29195 );
not \U$28820 ( \29197 , \29196 );
or \U$28821 ( \29198 , \29076 , \29197 );
or \U$28822 ( \29199 , \29196 , \29075 );
nand \U$28823 ( \29200 , \29198 , \29199 );
xor \U$28824 ( \29201 , \29030 , \29200 );
not \U$28825 ( \29202 , \29201 );
or \U$28826 ( \29203 , \29022 , \29202 );
or \U$28827 ( \29204 , \29021 , \29201 );
nand \U$28828 ( \29205 , \29203 , \29204 );
xnor \U$28829 ( \29206 , \29012 , \29205 );
not \U$28830 ( \29207 , \29206 );
or \U$28831 ( \29208 , \28686 , \29207 );
not \U$28832 ( \29209 , \28684 );
or \U$28833 ( \29210 , \29206 , \29209 );
nand \U$28834 ( \29211 , \29208 , \29210 );
not \U$28835 ( \29212 , \29211 );
xor \U$28836 ( \29213 , \28992 , \28986 );
not \U$28837 ( \29214 , \9777 );
not \U$28838 ( \29215 , RIae7a150_172);
not \U$28839 ( \29216 , \1789 );
or \U$28840 ( \29217 , \29215 , \29216 );
or \U$28841 ( \29218 , \1789 , RIae7a150_172);
nand \U$28842 ( \29219 , \29217 , \29218 );
not \U$28843 ( \29220 , \29219 );
or \U$28844 ( \29221 , \29214 , \29220 );
not \U$28845 ( \29222 , \2564 );
xor \U$28846 ( \29223 , RIae7a150_172, \29222 );
nand \U$28847 ( \29224 , \29223 , \13158 );
nand \U$28848 ( \29225 , \29221 , \29224 );
xor \U$28849 ( \29226 , \29213 , \29225 );
not \U$28850 ( \29227 , \16383 );
not \U$28851 ( \29228 , RIae7aa38_191);
not \U$28852 ( \29229 , \3051 );
or \U$28853 ( \29230 , \29228 , \29229 );
or \U$28854 ( \29231 , \2208 , RIae7aa38_191);
nand \U$28855 ( \29232 , \29230 , \29231 );
not \U$28856 ( \29233 , \29232 );
or \U$28857 ( \29234 , \29227 , \29233 );
xor \U$28858 ( \29235 , RIae7aa38_191, \1897 );
nand \U$28859 ( \29236 , \29235 , RIae7aab0_192);
nand \U$28860 ( \29237 , \29234 , \29236 );
and \U$28861 ( \29238 , \29226 , \29237 );
and \U$28862 ( \29239 , \29213 , \29225 );
or \U$28863 ( \29240 , \29238 , \29239 );
not \U$28864 ( \29241 , \2418 );
not \U$28865 ( \29242 , \28908 );
or \U$28866 ( \29243 , \29241 , \29242 );
not \U$28867 ( \29244 , RIae79c28_161);
not \U$28868 ( \29245 , \12483 );
or \U$28869 ( \29246 , \29244 , \29245 );
not \U$28870 ( \29247 , \12482 );
or \U$28871 ( \29248 , \29247 , RIae79c28_161);
nand \U$28872 ( \29249 , \29246 , \29248 );
nand \U$28873 ( \29250 , \29249 , \2417 );
nand \U$28874 ( \29251 , \29243 , \29250 );
not \U$28875 ( \29252 , \29251 );
not \U$28876 ( \29253 , \2431 );
and \U$28877 ( \29254 , RIae79778_151, \12644 );
not \U$28878 ( \29255 , RIae79778_151);
and \U$28879 ( \29256 , \29255 , \19015 );
nor \U$28880 ( \29257 , \29254 , \29256 );
not \U$28881 ( \29258 , \29257 );
or \U$28882 ( \29259 , \29253 , \29258 );
and \U$28883 ( \29260 , \10464 , \2447 );
not \U$28884 ( \29261 , \10464 );
and \U$28885 ( \29262 , \29261 , RIae79778_151);
nor \U$28886 ( \29263 , \29260 , \29262 );
nand \U$28887 ( \29264 , \29263 , \2450 );
nand \U$28888 ( \29265 , \29259 , \29264 );
not \U$28889 ( \29266 , \1988 );
xor \U$28890 ( \29267 , \10066 , RIae797f0_152);
not \U$28891 ( \29268 , \29267 );
or \U$28892 ( \29269 , \29266 , \29268 );
nand \U$28893 ( \29270 , \28027 , \2007 );
nand \U$28894 ( \29271 , \29269 , \29270 );
and \U$28895 ( \29272 , \29265 , \29271 );
not \U$28896 ( \29273 , \29265 );
not \U$28897 ( \29274 , \29271 );
and \U$28898 ( \29275 , \29273 , \29274 );
nor \U$28899 ( \29276 , \29272 , \29275 );
not \U$28900 ( \29277 , \29276 );
or \U$28901 ( \29278 , \29252 , \29277 );
nand \U$28902 ( \29279 , \29265 , \29271 );
nand \U$28903 ( \29280 , \29278 , \29279 );
nor \U$28904 ( \29281 , \29240 , \29280 );
not \U$28905 ( \29282 , \4154 );
not \U$28906 ( \29283 , RIae79ca0_162);
not \U$28907 ( \29284 , \14156 );
or \U$28908 ( \29285 , \29283 , \29284 );
not \U$28909 ( \29286 , \10936 );
or \U$28910 ( \29287 , \29286 , RIae79ca0_162);
nand \U$28911 ( \29288 , \29285 , \29287 );
not \U$28912 ( \29289 , \29288 );
or \U$28913 ( \29290 , \29282 , \29289 );
nand \U$28914 ( \29291 , \27933 , \4853 );
nand \U$28915 ( \29292 , \29290 , \29291 );
not \U$28916 ( \29293 , \5048 );
not \U$28917 ( \29294 , \28967 );
or \U$28918 ( \29295 , \29293 , \29294 );
not \U$28919 ( \29296 , \4968 );
not \U$28920 ( \29297 , \9438 );
or \U$28921 ( \29298 , \29296 , \29297 );
nand \U$28922 ( \29299 , \9442 , RIae79d90_164);
nand \U$28923 ( \29300 , \29298 , \29299 );
nand \U$28924 ( \29301 , \29300 , \6091 );
nand \U$28925 ( \29302 , \29295 , \29301 );
xor \U$28926 ( \29303 , \29292 , \29302 );
not \U$28927 ( \29304 , \10631 );
not \U$28928 ( \29305 , \27908 );
or \U$28929 ( \29306 , \29304 , \29305 );
not \U$28930 ( \29307 , \17324 );
not \U$28931 ( \29308 , \12502 );
or \U$28932 ( \29309 , \29307 , \29308 );
or \U$28933 ( \29310 , \17596 , \14931 );
nand \U$28934 ( \29311 , \29309 , \29310 );
nand \U$28935 ( \29312 , \29311 , \10927 );
nand \U$28936 ( \29313 , \29306 , \29312 );
and \U$28937 ( \29314 , \29303 , \29313 );
and \U$28938 ( \29315 , \29292 , \29302 );
or \U$28939 ( \29316 , \29314 , \29315 );
not \U$28940 ( \29317 , \29316 );
or \U$28941 ( \29318 , \29281 , \29317 );
nand \U$28942 ( \29319 , \29240 , \29280 );
nand \U$28943 ( \29320 , \29318 , \29319 );
xor \U$28944 ( \29321 , \28311 , \28325 );
xor \U$28945 ( \29322 , \29321 , \28342 );
not \U$28946 ( \29323 , \29322 );
not \U$28947 ( \29324 , \9621 );
not \U$28948 ( \29325 , \27531 );
or \U$28949 ( \29326 , \29324 , \29325 );
nand \U$28950 ( \29327 , \27821 , \11013 );
nand \U$28951 ( \29328 , \29326 , \29327 );
not \U$28952 ( \29329 , RIae7aab0_192);
not \U$28953 ( \29330 , \27866 );
or \U$28954 ( \29331 , \29329 , \29330 );
nand \U$28955 ( \29332 , \29235 , \14667 );
nand \U$28956 ( \29333 , \29331 , \29332 );
xor \U$28957 ( \29334 , \29328 , \29333 );
not \U$28958 ( \29335 , \9744 );
not \U$28959 ( \29336 , \27873 );
or \U$28960 ( \29337 , \29335 , \29336 );
not \U$28961 ( \29338 , \9749 );
not \U$28962 ( \29339 , \24445 );
or \U$28963 ( \29340 , \29338 , \29339 );
nand \U$28964 ( \29341 , \10905 , RIae7a060_170);
nand \U$28965 ( \29342 , \29340 , \29341 );
nand \U$28966 ( \29343 , \29342 , \9730 );
nand \U$28967 ( \29344 , \29337 , \29343 );
and \U$28968 ( \29345 , \29334 , \29344 );
and \U$28969 ( \29346 , \29328 , \29333 );
or \U$28970 ( \29347 , \29345 , \29346 );
not \U$28971 ( \29348 , \28202 );
xor \U$28972 ( \29349 , \28217 , \28232 );
not \U$28973 ( \29350 , \29349 );
or \U$28974 ( \29351 , \29348 , \29350 );
or \U$28975 ( \29352 , \28202 , \29349 );
nand \U$28976 ( \29353 , \29351 , \29352 );
xor \U$28977 ( \29354 , \29347 , \29353 );
not \U$28978 ( \29355 , \29354 );
or \U$28979 ( \29356 , \29323 , \29355 );
or \U$28980 ( \29357 , \29322 , \29354 );
nand \U$28981 ( \29358 , \29356 , \29357 );
xor \U$28982 ( \29359 , \29320 , \29358 );
not \U$28983 ( \29360 , \15382 );
and \U$28984 ( \29361 , \1956 , RIae7a498_179);
not \U$28985 ( \29362 , \1956 );
and \U$28986 ( \29363 , \29362 , \11427 );
nor \U$28987 ( \29364 , \29361 , \29363 );
not \U$28988 ( \29365 , \29364 );
or \U$28989 ( \29366 , \29360 , \29365 );
nand \U$28990 ( \29367 , \27959 , \10675 );
nand \U$28991 ( \29368 , \29366 , \29367 );
not \U$28992 ( \29369 , \29368 );
not \U$28993 ( \29370 , \2322 );
not \U$28994 ( \29371 , \28002 );
or \U$28995 ( \29372 , \29370 , \29371 );
and \U$28996 ( \29373 , \10000 , \21036 );
not \U$28997 ( \29374 , \10000 );
and \U$28998 ( \29375 , \29374 , RIae798e0_154);
nor \U$28999 ( \29376 , \29373 , \29375 );
nand \U$29000 ( \29377 , \29376 , \2339 );
nand \U$29001 ( \29378 , \29372 , \29377 );
not \U$29002 ( \29379 , \29378 );
not \U$29003 ( \29380 , \2249 );
not \U$29004 ( \29381 , \28980 );
or \U$29005 ( \29382 , \29380 , \29381 );
not \U$29006 ( \29383 , \2268 );
not \U$29007 ( \29384 , \10272 );
or \U$29008 ( \29385 , \29383 , \29384 );
or \U$29009 ( \29386 , \10272 , \2268 );
nand \U$29010 ( \29387 , \29385 , \29386 );
nand \U$29011 ( \29388 , \29387 , \2272 );
nand \U$29012 ( \29389 , \29382 , \29388 );
not \U$29013 ( \29390 , \2249 );
not \U$29014 ( \29391 , \29387 );
or \U$29015 ( \29392 , \29390 , \29391 );
not \U$29016 ( \29393 , \17155 );
xor \U$29017 ( \29394 , RIae79ac0_158, \29393 );
nand \U$29018 ( \29395 , \29394 , \2272 );
nand \U$29019 ( \29396 , \29392 , \29395 );
not \U$29020 ( \29397 , \29396 );
not \U$29021 ( \29398 , \1818 );
not \U$29022 ( \29399 , \27751 );
or \U$29023 ( \29400 , \29398 , \29399 );
and \U$29024 ( \29401 , \3147 , \12750 );
not \U$29025 ( \29402 , \3147 );
and \U$29026 ( \29403 , \29402 , \18985 );
nor \U$29027 ( \29404 , \29401 , \29403 );
nand \U$29028 ( \29405 , \29404 , \1842 );
nand \U$29029 ( \29406 , \29400 , \29405 );
not \U$29030 ( \29407 , \29406 );
and \U$29031 ( \29408 , \12857 , \2011 );
not \U$29032 ( \29409 , \29408 );
and \U$29033 ( \29410 , \29407 , \29409 );
not \U$29034 ( \29411 , \29407 );
and \U$29035 ( \29412 , \29411 , \29408 );
nor \U$29036 ( \29413 , \29410 , \29412 );
not \U$29037 ( \29414 , \29413 );
or \U$29038 ( \29415 , \29397 , \29414 );
nand \U$29039 ( \29416 , \29406 , \29408 );
nand \U$29040 ( \29417 , \29415 , \29416 );
xor \U$29041 ( \29418 , \29389 , \29417 );
not \U$29042 ( \29419 , \29418 );
or \U$29043 ( \29420 , \29379 , \29419 );
nand \U$29044 ( \29421 , \29417 , \29389 );
nand \U$29045 ( \29422 , \29420 , \29421 );
not \U$29046 ( \29423 , \9478 );
and \U$29047 ( \29424 , RIae7a6f0_184, \2955 );
not \U$29048 ( \29425 , RIae7a6f0_184);
and \U$29049 ( \29426 , \29425 , \2954 );
nor \U$29050 ( \29427 , \29424 , \29426 );
not \U$29051 ( \29428 , \29427 );
or \U$29052 ( \29429 , \29423 , \29428 );
and \U$29053 ( \29430 , \16101 , \2309 );
not \U$29054 ( \29431 , \16101 );
and \U$29055 ( \29432 , \29431 , \2305 );
or \U$29056 ( \29433 , \29430 , \29432 );
nand \U$29057 ( \29434 , \29433 , \9473 );
nand \U$29058 ( \29435 , \29429 , \29434 );
and \U$29059 ( \29436 , \29422 , \29435 );
not \U$29060 ( \29437 , \29422 );
not \U$29061 ( \29438 , \29435 );
and \U$29062 ( \29439 , \29437 , \29438 );
nor \U$29063 ( \29440 , \29436 , \29439 );
not \U$29064 ( \29441 , \29440 );
or \U$29065 ( \29442 , \29369 , \29441 );
nand \U$29066 ( \29443 , \29435 , \29422 );
nand \U$29067 ( \29444 , \29442 , \29443 );
not \U$29068 ( \29445 , \2450 );
not \U$29069 ( \29446 , \28208 );
or \U$29070 ( \29447 , \29445 , \29446 );
nand \U$29071 ( \29448 , \29263 , \2431 );
nand \U$29072 ( \29449 , \29447 , \29448 );
not \U$29073 ( \29450 , \9814 );
not \U$29074 ( \29451 , \28192 );
or \U$29075 ( \29452 , \29450 , \29451 );
nand \U$29076 ( \29453 , \27831 , \9792 );
nand \U$29077 ( \29454 , \29452 , \29453 );
xor \U$29078 ( \29455 , \29449 , \29454 );
not \U$29079 ( \29456 , \13130 );
not \U$29080 ( \29457 , \27845 );
or \U$29081 ( \29458 , \29456 , \29457 );
nand \U$29082 ( \29459 , \28947 , \13121 );
nand \U$29083 ( \29460 , \29458 , \29459 );
xor \U$29084 ( \29461 , \29455 , \29460 );
xor \U$29085 ( \29462 , \29444 , \29461 );
not \U$29086 ( \29463 , \9776 );
not \U$29087 ( \29464 , \27544 );
or \U$29088 ( \29465 , \29463 , \29464 );
nand \U$29089 ( \29466 , \29219 , \10667 );
nand \U$29090 ( \29467 , \29465 , \29466 );
not \U$29091 ( \29468 , \10275 );
not \U$29092 ( \29469 , \27885 );
or \U$29093 ( \29470 , \29468 , \29469 );
not \U$29094 ( \29471 , \18088 );
not \U$29095 ( \29472 , \3765 );
or \U$29096 ( \29473 , \29471 , \29472 );
nand \U$29097 ( \29474 , \2993 , RIae7a8d0_188);
nand \U$29098 ( \29475 , \29473 , \29474 );
nand \U$29099 ( \29476 , \29475 , \14510 );
nand \U$29100 ( \29477 , \29470 , \29476 );
xor \U$29101 ( \29478 , \29467 , \29477 );
not \U$29102 ( \29479 , \9705 );
not \U$29103 ( \29480 , \27657 );
or \U$29104 ( \29481 , \29479 , \29480 );
nand \U$29105 ( \29482 , \29427 , \9473 );
nand \U$29106 ( \29483 , \29481 , \29482 );
xor \U$29107 ( \29484 , \29478 , \29483 );
and \U$29108 ( \29485 , \29462 , \29484 );
and \U$29109 ( \29486 , \29444 , \29461 );
or \U$29110 ( \29487 , \29485 , \29486 );
and \U$29111 ( \29488 , \29359 , \29487 );
and \U$29112 ( \29489 , \29320 , \29358 );
or \U$29113 ( \29490 , \29488 , \29489 );
not \U$29114 ( \29491 , \29005 );
not \U$29115 ( \29492 , \29491 );
not \U$29116 ( \29493 , \28925 );
nand \U$29117 ( \29494 , \29493 , \29008 );
not \U$29118 ( \29495 , \29494 );
and \U$29119 ( \29496 , \29492 , \29495 );
and \U$29120 ( \29497 , \29494 , \29491 );
nor \U$29121 ( \29498 , \29496 , \29497 );
nor \U$29122 ( \29499 , \29490 , \29498 );
not \U$29123 ( \29500 , \17847 );
not \U$29124 ( \29501 , \9501 );
not \U$29125 ( \29502 , RIae7a8d0_188);
and \U$29126 ( \29503 , \29501 , \29502 );
and \U$29127 ( \29504 , \3070 , RIae7a8d0_188);
nor \U$29128 ( \29505 , \29503 , \29504 );
not \U$29129 ( \29506 , \29505 );
or \U$29130 ( \29507 , \29500 , \29506 );
nand \U$29131 ( \29508 , \29475 , \10275 );
nand \U$29132 ( \29509 , \29507 , \29508 );
not \U$29133 ( \29510 , \9549 );
not \U$29134 ( \29511 , \9529 );
not \U$29135 ( \29512 , \3094 );
or \U$29136 ( \29513 , \29511 , \29512 );
or \U$29137 ( \29514 , \13671 , \9541 );
nand \U$29138 ( \29515 , \29513 , \29514 );
not \U$29139 ( \29516 , \29515 );
or \U$29140 ( \29517 , \29510 , \29516 );
not \U$29141 ( \29518 , \9526 );
buf \U$29142 ( \29519 , \29518 );
nand \U$29143 ( \29520 , \27919 , \29519 );
nand \U$29144 ( \29521 , \29517 , \29520 );
or \U$29145 ( \29522 , \29509 , \29521 );
not \U$29146 ( \29523 , \9730 );
and \U$29147 ( \29524 , RIae7a060_170, \3524 );
not \U$29148 ( \29525 , RIae7a060_170);
and \U$29149 ( \29526 , \29525 , \10884 );
or \U$29150 ( \29527 , \29524 , \29526 );
not \U$29151 ( \29528 , \29527 );
or \U$29152 ( \29529 , \29523 , \29528 );
nand \U$29153 ( \29530 , \29342 , \9744 );
nand \U$29154 ( \29531 , \29529 , \29530 );
nand \U$29155 ( \29532 , \29522 , \29531 );
nand \U$29156 ( \29533 , \29509 , \29521 );
nand \U$29157 ( \29534 , \29532 , \29533 );
not \U$29158 ( \29535 , \29534 );
xnor \U$29159 ( \29536 , \28916 , \28879 );
not \U$29160 ( \29537 , \29536 );
xor \U$29161 ( \29538 , \28997 , \28958 );
xor \U$29162 ( \29539 , \29538 , \28969 );
not \U$29163 ( \29540 , \29539 );
or \U$29164 ( \29541 , \29537 , \29540 );
or \U$29165 ( \29542 , \29539 , \29536 );
nand \U$29166 ( \29543 , \29541 , \29542 );
not \U$29167 ( \29544 , \29543 );
or \U$29168 ( \29545 , \29535 , \29544 );
not \U$29169 ( \29546 , \29536 );
nand \U$29170 ( \29547 , \29546 , \29539 );
nand \U$29171 ( \29548 , \29545 , \29547 );
not \U$29172 ( \29549 , \29548 );
not \U$29173 ( \29550 , \28872 );
nand \U$29174 ( \29551 , \29550 , \28923 );
xor \U$29175 ( \29552 , \28920 , \29551 );
not \U$29176 ( \29553 , \29552 );
xor \U$29177 ( \29554 , \28929 , \28952 );
xor \U$29178 ( \29555 , \29554 , \29002 );
not \U$29179 ( \29556 , \29555 );
or \U$29180 ( \29557 , \29553 , \29556 );
or \U$29181 ( \29558 , \29555 , \29552 );
nand \U$29182 ( \29559 , \29557 , \29558 );
not \U$29183 ( \29560 , \29559 );
or \U$29184 ( \29561 , \29549 , \29560 );
not \U$29185 ( \29562 , \29552 );
nand \U$29186 ( \29563 , \29562 , \29555 );
nand \U$29187 ( \29564 , \29561 , \29563 );
not \U$29188 ( \29565 , \29564 );
or \U$29189 ( \29566 , \29499 , \29565 );
nand \U$29190 ( \29567 , \29490 , \29498 );
nand \U$29191 ( \29568 , \29566 , \29567 );
and \U$29192 ( \29569 , \29009 , \28854 );
not \U$29193 ( \29570 , \29009 );
and \U$29194 ( \29571 , \29570 , \28855 );
or \U$29195 ( \29572 , \29569 , \29571 );
and \U$29196 ( \29573 , \29572 , \28810 );
not \U$29197 ( \29574 , \29572 );
and \U$29198 ( \29575 , \29574 , \28809 );
nor \U$29199 ( \29576 , \29573 , \29575 );
nand \U$29200 ( \29577 , \29568 , \29576 );
not \U$29201 ( \29578 , \28617 );
not \U$29202 ( \29579 , \29578 );
not \U$29203 ( \29580 , \28632 );
or \U$29204 ( \29581 , \29579 , \29580 );
nand \U$29205 ( \29582 , \28601 , \28612 );
nand \U$29206 ( \29583 , \29581 , \29582 );
not \U$29207 ( \29584 , \2249 );
not \U$29208 ( \29585 , \10419 );
not \U$29209 ( \29586 , \10743 );
or \U$29210 ( \29587 , \29585 , \29586 );
nand \U$29211 ( \29588 , \16193 , RIae79ac0_158);
nand \U$29212 ( \29589 , \29587 , \29588 );
not \U$29213 ( \29590 , \29589 );
or \U$29214 ( \29591 , \29584 , \29590 );
nand \U$29215 ( \29592 , \27616 , \2272 );
nand \U$29216 ( \29593 , \29591 , \29592 );
not \U$29217 ( \29594 , \2162 );
not \U$29218 ( \29595 , RIae79520_146);
not \U$29219 ( \29596 , \9875 );
or \U$29220 ( \29597 , \29595 , \29596 );
or \U$29221 ( \29598 , \9875 , RIae79520_146);
nand \U$29222 ( \29599 , \29597 , \29598 );
not \U$29223 ( \29600 , \29599 );
or \U$29224 ( \29601 , \29594 , \29600 );
nand \U$29225 ( \29602 , \28280 , \2188 );
nand \U$29226 ( \29603 , \29601 , \29602 );
xor \U$29227 ( \29604 , \29593 , \29603 );
not \U$29228 ( \29605 , \1919 );
not \U$29229 ( \29606 , RIae794a8_145);
not \U$29230 ( \29607 , \11230 );
or \U$29231 ( \29608 , \29606 , \29607 );
or \U$29232 ( \29609 , \11562 , RIae794a8_145);
nand \U$29233 ( \29610 , \29608 , \29609 );
not \U$29234 ( \29611 , \29610 );
or \U$29235 ( \29612 , \29605 , \29611 );
nand \U$29236 ( \29613 , \28938 , \1932 );
nand \U$29237 ( \29614 , \29612 , \29613 );
and \U$29238 ( \29615 , \29604 , \29614 );
and \U$29239 ( \29616 , \29593 , \29603 );
nor \U$29240 ( \29617 , \29615 , \29616 );
and \U$29241 ( \29618 , \29583 , \29617 );
not \U$29242 ( \29619 , \29583 );
not \U$29243 ( \29620 , \29617 );
and \U$29244 ( \29621 , \29619 , \29620 );
or \U$29245 ( \29622 , \29618 , \29621 );
not \U$29246 ( \29623 , \10696 );
not \U$29247 ( \29624 , \28641 );
or \U$29248 ( \29625 , \29623 , \29624 );
not \U$29249 ( \29626 , \10625 );
not \U$29250 ( \29627 , \1759 );
or \U$29251 ( \29628 , \29626 , \29627 );
nand \U$29252 ( \29629 , \10608 , RIae7a498_179);
nand \U$29253 ( \29630 , \29628 , \29629 );
nand \U$29254 ( \29631 , \29630 , \10675 );
nand \U$29255 ( \29632 , \29625 , \29631 );
xor \U$29256 ( \29633 , \29622 , \29632 );
not \U$29257 ( \29634 , \28428 );
not \U$29258 ( \29635 , \29634 );
not \U$29259 ( \29636 , \28432 );
or \U$29260 ( \29637 , \29635 , \29636 );
nand \U$29261 ( \29638 , \29637 , \28441 );
nand \U$29262 ( \29639 , \28430 , \28431 , \28428 );
and \U$29263 ( \29640 , \29638 , \29639 );
xor \U$29264 ( \29641 , \29633 , \29640 );
not \U$29265 ( \29642 , \28237 );
and \U$29266 ( \29643 , \28347 , \29642 );
and \U$29267 ( \29644 , \28295 , \28346 );
nor \U$29268 ( \29645 , \29643 , \29644 );
xor \U$29269 ( \29646 , \29641 , \29645 );
xor \U$29270 ( \29647 , \29593 , \29614 );
xnor \U$29271 ( \29648 , \29647 , \29603 );
not \U$29272 ( \29649 , \29648 );
not \U$29273 ( \29650 , \10638 );
not \U$29274 ( \29651 , \27901 );
or \U$29275 ( \29652 , \29650 , \29651 );
nand \U$29276 ( \29653 , \28121 , \16358 );
nand \U$29277 ( \29654 , \29652 , \29653 );
not \U$29278 ( \29655 , \29654 );
xor \U$29279 ( \29656 , \28885 , \28891 );
and \U$29280 ( \29657 , \29656 , \28898 );
and \U$29281 ( \29658 , \28885 , \28891 );
nor \U$29282 ( \29659 , \29657 , \29658 );
not \U$29283 ( \29660 , \29659 );
not \U$29284 ( \29661 , \11761 );
not \U$29285 ( \29662 , \27926 );
or \U$29286 ( \29663 , \29661 , \29662 );
nand \U$29287 ( \29664 , \28106 , \4853 );
nand \U$29288 ( \29665 , \29663 , \29664 );
not \U$29289 ( \29666 , \29665 );
or \U$29290 ( \29667 , \29660 , \29666 );
or \U$29291 ( \29668 , \29665 , \29659 );
nand \U$29292 ( \29669 , \29667 , \29668 );
not \U$29293 ( \29670 , \29669 );
or \U$29294 ( \29671 , \29655 , \29670 );
not \U$29295 ( \29672 , \29659 );
nand \U$29296 ( \29673 , \29672 , \29665 );
nand \U$29297 ( \29674 , \29671 , \29673 );
nor \U$29298 ( \29675 , \29649 , \29674 );
nand \U$29299 ( \29676 , \28951 , \28941 );
nand \U$29300 ( \29677 , \28940 , \28934 );
and \U$29301 ( \29678 , \29676 , \29677 );
or \U$29302 ( \29679 , \29675 , \29678 );
not \U$29303 ( \29680 , \29648 );
nand \U$29304 ( \29681 , \29680 , \29674 );
nand \U$29305 ( \29682 , \29679 , \29681 );
not \U$29306 ( \29683 , \1932 );
not \U$29307 ( \29684 , \29610 );
or \U$29308 ( \29685 , \29683 , \29684 );
not \U$29309 ( \29686 , RIae794a8_145);
not \U$29310 ( \29687 , \10084 );
or \U$29311 ( \29688 , \29686 , \29687 );
or \U$29312 ( \29689 , \10084 , RIae794a8_145);
nand \U$29313 ( \29690 , \29688 , \29689 );
nand \U$29314 ( \29691 , \29690 , \1919 );
nand \U$29315 ( \29692 , \29685 , \29691 );
and \U$29316 ( \29693 , \12857 , \1012 );
not \U$29317 ( \29694 , \1501 );
not \U$29318 ( \29695 , \29115 );
or \U$29319 ( \29696 , \29694 , \29695 );
nand \U$29320 ( \29697 , \28385 , \1497 );
nand \U$29321 ( \29698 , \29696 , \29697 );
xor \U$29322 ( \29699 , \29693 , \29698 );
not \U$29323 ( \29700 , \1863 );
not \U$29324 ( \29701 , \12842 );
not \U$29325 ( \29702 , RIae793b8_143);
and \U$29326 ( \29703 , \29701 , \29702 );
and \U$29327 ( \29704 , \11318 , RIae793b8_143);
nor \U$29328 ( \29705 , \29703 , \29704 );
not \U$29329 ( \29706 , \29705 );
or \U$29330 ( \29707 , \29700 , \29706 );
nand \U$29331 ( \29708 , \28375 , \1909 );
nand \U$29332 ( \29709 , \29707 , \29708 );
xor \U$29333 ( \29710 , \29699 , \29709 );
and \U$29334 ( \29711 , \29692 , \29710 );
not \U$29335 ( \29712 , \29692 );
not \U$29336 ( \29713 , \29710 );
and \U$29337 ( \29714 , \29712 , \29713 );
nor \U$29338 ( \29715 , \29711 , \29714 );
buf \U$29339 ( \29716 , \29715 );
not \U$29340 ( \29717 , \2339 );
not \U$29341 ( \29718 , \28623 );
or \U$29342 ( \29719 , \29717 , \29718 );
nand \U$29343 ( \29720 , \29166 , \2322 );
nand \U$29344 ( \29721 , \29719 , \29720 );
and \U$29345 ( \29722 , \29716 , \29721 );
not \U$29346 ( \29723 , \29716 );
not \U$29347 ( \29724 , \29721 );
and \U$29348 ( \29725 , \29723 , \29724 );
nor \U$29349 ( \29726 , \29722 , \29725 );
not \U$29350 ( \29727 , \2776 );
not \U$29351 ( \29728 , \29052 );
or \U$29352 ( \29729 , \29727 , \29728 );
nand \U$29353 ( \29730 , \28470 , \2767 );
nand \U$29354 ( \29731 , \29729 , \29730 );
not \U$29355 ( \29732 , \29589 );
not \U$29356 ( \29733 , \29732 );
not \U$29357 ( \29734 , \3510 );
and \U$29358 ( \29735 , \29733 , \29734 );
not \U$29359 ( \29736 , RIae79ac0_158);
not \U$29360 ( \29737 , \16719 );
or \U$29361 ( \29738 , \29736 , \29737 );
or \U$29362 ( \29739 , \10000 , RIae79ac0_158);
nand \U$29363 ( \29740 , \29738 , \29739 );
and \U$29364 ( \29741 , \29740 , \10414 );
nor \U$29365 ( \29742 , \29735 , \29741 );
not \U$29366 ( \29743 , \29742 );
not \U$29367 ( \29744 , \2602 );
not \U$29368 ( \29745 , \29599 );
or \U$29369 ( \29746 , \29744 , \29745 );
not \U$29370 ( \29747 , RIae79520_146);
not \U$29371 ( \29748 , \10168 );
or \U$29372 ( \29749 , \29747 , \29748 );
nand \U$29373 ( \29750 , \14546 , \4653 );
nand \U$29374 ( \29751 , \29749 , \29750 );
nand \U$29375 ( \29752 , \29751 , \2163 );
nand \U$29376 ( \29753 , \29746 , \29752 );
not \U$29377 ( \29754 , \29753 );
or \U$29378 ( \29755 , \29743 , \29754 );
or \U$29379 ( \29756 , \29753 , \29742 );
nand \U$29380 ( \29757 , \29755 , \29756 );
and \U$29381 ( \29758 , \29731 , \29757 );
not \U$29382 ( \29759 , \29731 );
not \U$29383 ( \29760 , \29757 );
and \U$29384 ( \29761 , \29759 , \29760 );
nor \U$29385 ( \29762 , \29758 , \29761 );
xor \U$29386 ( \29763 , \29726 , \29762 );
not \U$29387 ( \29764 , \29763 );
not \U$29388 ( \29765 , \28139 );
not \U$29389 ( \29766 , \28126 );
or \U$29390 ( \29767 , \29765 , \29766 );
nand \U$29391 ( \29768 , \29767 , \28108 );
nand \U$29392 ( \29769 , \28123 , \28138 );
nand \U$29393 ( \29770 , \29768 , \29769 );
not \U$29394 ( \29771 , \29770 );
not \U$29395 ( \29772 , \29771 );
or \U$29396 ( \29773 , \29764 , \29772 );
not \U$29397 ( \29774 , \29763 );
nand \U$29398 ( \29775 , \29774 , \29770 );
nand \U$29399 ( \29776 , \29773 , \29775 );
xor \U$29400 ( \29777 , \29682 , \29776 );
not \U$29401 ( \29778 , \28423 );
not \U$29402 ( \29779 , \28413 );
or \U$29403 ( \29780 , \29778 , \29779 );
not \U$29404 ( \29781 , \28409 );
nand \U$29405 ( \29782 , \29781 , \28357 );
nand \U$29406 ( \29783 , \29780 , \29782 );
not \U$29407 ( \29784 , \29783 );
and \U$29408 ( \29785 , \28464 , \28474 );
and \U$29409 ( \29786 , \28453 , \28463 );
nor \U$29410 ( \29787 , \29785 , \29786 );
not \U$29411 ( \29788 , \29787 );
or \U$29412 ( \29789 , \29784 , \29788 );
or \U$29413 ( \29790 , \29787 , \29783 );
nand \U$29414 ( \29791 , \29789 , \29790 );
not \U$29415 ( \29792 , \28514 );
not \U$29416 ( \29793 , \28493 );
not \U$29417 ( \29794 , \29793 );
not \U$29418 ( \29795 , \28503 );
or \U$29419 ( \29796 , \29794 , \29795 );
or \U$29420 ( \29797 , \28503 , \29793 );
nand \U$29421 ( \29798 , \29796 , \29797 );
not \U$29422 ( \29799 , \29798 );
or \U$29423 ( \29800 , \29792 , \29799 );
nand \U$29424 ( \29801 , \28503 , \28493 );
nand \U$29425 ( \29802 , \29800 , \29801 );
not \U$29426 ( \29803 , \29802 );
and \U$29427 ( \29804 , \29791 , \29803 );
not \U$29428 ( \29805 , \29791 );
and \U$29429 ( \29806 , \29805 , \29802 );
or \U$29430 ( \29807 , \29804 , \29806 );
xor \U$29431 ( \29808 , \29777 , \29807 );
xor \U$29432 ( \29809 , \29646 , \29808 );
nor \U$29433 ( \29810 , \29347 , \29322 );
or \U$29434 ( \29811 , \29810 , \29353 );
nand \U$29435 ( \29812 , \29322 , \29347 );
nand \U$29436 ( \29813 , \29811 , \29812 );
not \U$29437 ( \29814 , \29813 );
xor \U$29438 ( \29815 , \29648 , \29674 );
xnor \U$29439 ( \29816 , \29815 , \29678 );
nand \U$29440 ( \29817 , \29814 , \29816 );
not \U$29441 ( \29818 , \29817 );
xor \U$29442 ( \29819 , \29669 , \29654 );
not \U$29443 ( \29820 , \29819 );
xor \U$29444 ( \29821 , \29449 , \29454 );
and \U$29445 ( \29822 , \29821 , \29460 );
and \U$29446 ( \29823 , \29449 , \29454 );
nor \U$29447 ( \29824 , \29822 , \29823 );
not \U$29448 ( \29825 , \29824 );
xor \U$29449 ( \29826 , \29467 , \29477 );
and \U$29450 ( \29827 , \29826 , \29483 );
and \U$29451 ( \29828 , \29467 , \29477 );
or \U$29452 ( \29829 , \29827 , \29828 );
not \U$29453 ( \29830 , \29829 );
or \U$29454 ( \29831 , \29825 , \29830 );
or \U$29455 ( \29832 , \29824 , \29829 );
nand \U$29456 ( \29833 , \29831 , \29832 );
not \U$29457 ( \29834 , \29833 );
or \U$29458 ( \29835 , \29820 , \29834 );
not \U$29459 ( \29836 , \29824 );
nand \U$29460 ( \29837 , \29836 , \29829 );
nand \U$29461 ( \29838 , \29835 , \29837 );
not \U$29462 ( \29839 , \29838 );
or \U$29463 ( \29840 , \29818 , \29839 );
not \U$29464 ( \29841 , \29816 );
nand \U$29465 ( \29842 , \29841 , \29813 );
nand \U$29466 ( \29843 , \29840 , \29842 );
not \U$29467 ( \29844 , \29843 );
and \U$29468 ( \29845 , \29809 , \29844 );
not \U$29469 ( \29846 , \29809 );
and \U$29470 ( \29847 , \29846 , \29843 );
nor \U$29471 ( \29848 , \29845 , \29847 );
and \U$29472 ( \29849 , \29577 , \29848 );
nor \U$29473 ( \29850 , \29568 , \29576 );
nor \U$29474 ( \29851 , \29849 , \29850 );
buf \U$29475 ( \29852 , \29851 );
not \U$29476 ( \29853 , \29852 );
and \U$29477 ( \29854 , \29212 , \29853 );
and \U$29478 ( \29855 , \29852 , \29211 );
nor \U$29479 ( \29856 , \29854 , \29855 );
not \U$29480 ( \29857 , \29856 );
not \U$29481 ( \29858 , \29646 );
not \U$29482 ( \29859 , \29808 );
or \U$29483 ( \29860 , \29858 , \29859 );
or \U$29484 ( \29861 , \29808 , \29646 );
nand \U$29485 ( \29862 , \29861 , \29843 );
nand \U$29486 ( \29863 , \29860 , \29862 );
not \U$29487 ( \29864 , \10631 );
not \U$29488 ( \29865 , \17324 );
not \U$29489 ( \29866 , \4036 );
or \U$29490 ( \29867 , \29865 , \29866 );
nand \U$29491 ( \29868 , \3524 , RIae7a510_180);
nand \U$29492 ( \29869 , \29867 , \29868 );
not \U$29493 ( \29870 , \29869 );
or \U$29494 ( \29871 , \29864 , \29870 );
nand \U$29495 ( \29872 , \28792 , \10927 );
nand \U$29496 ( \29873 , \29871 , \29872 );
not \U$29497 ( \29874 , \28757 );
not \U$29498 ( \29875 , \28748 );
not \U$29499 ( \29876 , \29875 );
or \U$29500 ( \29877 , \29874 , \29876 );
not \U$29501 ( \29878 , \28747 );
nand \U$29502 ( \29879 , \29878 , \28745 );
nand \U$29503 ( \29880 , \29877 , \29879 );
not \U$29504 ( \29881 , \29880 );
not \U$29505 ( \29882 , \16594 );
not \U$29506 ( \29883 , \28697 );
or \U$29507 ( \29884 , \29882 , \29883 );
not \U$29508 ( \29885 , \18088 );
not \U$29509 ( \29886 , \2025 );
or \U$29510 ( \29887 , \29885 , \29886 );
or \U$29511 ( \29888 , \2025 , \11207 );
nand \U$29512 ( \29889 , \29887 , \29888 );
nand \U$29513 ( \29890 , \29889 , \10275 );
nand \U$29514 ( \29891 , \29884 , \29890 );
not \U$29515 ( \29892 , \29891 );
not \U$29516 ( \29893 , \29892 );
or \U$29517 ( \29894 , \29881 , \29893 );
or \U$29518 ( \29895 , \29892 , \29880 );
nand \U$29519 ( \29896 , \29894 , \29895 );
xor \U$29520 ( \29897 , \29873 , \29896 );
not \U$29521 ( \29898 , \29897 );
not \U$29522 ( \29899 , \28817 );
not \U$29523 ( \29900 , \28834 );
or \U$29524 ( \29901 , \29899 , \29900 );
not \U$29525 ( \29902 , \28825 );
not \U$29526 ( \29903 , \28819 );
or \U$29527 ( \29904 , \29902 , \29903 );
nand \U$29528 ( \29905 , \29904 , \28833 );
nand \U$29529 ( \29906 , \29901 , \29905 );
not \U$29530 ( \29907 , \29906 );
not \U$29531 ( \29908 , \29907 );
or \U$29532 ( \29909 , \29898 , \29908 );
or \U$29533 ( \29910 , \29907 , \29897 );
nand \U$29534 ( \29911 , \29909 , \29910 );
not \U$29535 ( \29912 , \9622 );
and \U$29536 ( \29913 , RIae7a3a8_177, \2676 );
not \U$29537 ( \29914 , RIae7a3a8_177);
and \U$29538 ( \29915 , \29914 , \4837 );
or \U$29539 ( \29916 , \29913 , \29915 );
not \U$29540 ( \29917 , \29916 );
or \U$29541 ( \29918 , \29912 , \29917 );
nand \U$29542 ( \29919 , \28783 , \9644 );
nand \U$29543 ( \29920 , \29918 , \29919 );
not \U$29544 ( \29921 , \13121 );
and \U$29545 ( \29922 , RIae7a240_174, \1956 );
not \U$29546 ( \29923 , RIae7a240_174);
and \U$29547 ( \29924 , \29923 , \4113 );
nor \U$29548 ( \29925 , \29922 , \29924 );
not \U$29549 ( \29926 , \29925 );
or \U$29550 ( \29927 , \29921 , \29926 );
nand \U$29551 ( \29928 , \28706 , \19466 );
nand \U$29552 ( \29929 , \29927 , \29928 );
nor \U$29553 ( \29930 , \29920 , \29929 );
not \U$29554 ( \29931 , \29930 );
nand \U$29555 ( \29932 , \29920 , \29929 );
nand \U$29556 ( \29933 , \29931 , \29932 );
not \U$29557 ( \29934 , \10519 );
not \U$29558 ( \29935 , RIae7a7e0_186);
not \U$29559 ( \29936 , \9797 );
or \U$29560 ( \29937 , \29935 , \29936 );
nand \U$29561 ( \29938 , \2628 , \9537 );
nand \U$29562 ( \29939 , \29937 , \29938 );
not \U$29563 ( \29940 , \29939 );
or \U$29564 ( \29941 , \29934 , \29940 );
nand \U$29565 ( \29942 , \28803 , \10510 );
nand \U$29566 ( \29943 , \29941 , \29942 );
not \U$29567 ( \29944 , \29943 );
and \U$29568 ( \29945 , \29933 , \29944 );
not \U$29569 ( \29946 , \29933 );
and \U$29570 ( \29947 , \29946 , \29943 );
nor \U$29571 ( \29948 , \29945 , \29947 );
xnor \U$29572 ( \29949 , \29911 , \29948 );
not \U$29573 ( \29950 , \29949 );
not \U$29574 ( \29951 , \29950 );
not \U$29575 ( \29952 , \29632 );
not \U$29576 ( \29953 , \29952 );
not \U$29577 ( \29954 , \29617 );
or \U$29578 ( \29955 , \29953 , \29954 );
nand \U$29579 ( \29956 , \29955 , \29583 );
nand \U$29580 ( \29957 , \29620 , \29632 );
and \U$29581 ( \29958 , \29956 , \29957 );
not \U$29582 ( \29959 , \11422 );
and \U$29583 ( \29960 , RIae7a498_179, \21317 );
not \U$29584 ( \29961 , RIae7a498_179);
and \U$29585 ( \29962 , \29961 , \13671 );
or \U$29586 ( \29963 , \29960 , \29962 );
not \U$29587 ( \29964 , \29963 );
or \U$29588 ( \29965 , \29959 , \29964 );
nand \U$29589 ( \29966 , \29630 , \10696 );
nand \U$29590 ( \29967 , \29965 , \29966 );
not \U$29591 ( \29968 , \29967 );
not \U$29592 ( \29969 , \9478 );
not \U$29593 ( \29970 , \1878 );
xor \U$29594 ( \29971 , RIae7a6f0_184, \29970 );
not \U$29595 ( \29972 , \29971 );
or \U$29596 ( \29973 , \29969 , \29972 );
nand \U$29597 ( \29974 , \28733 , \9473 );
nand \U$29598 ( \29975 , \29973 , \29974 );
not \U$29599 ( \29976 , \29975 );
not \U$29600 ( \29977 , \29976 );
and \U$29601 ( \29978 , \29968 , \29977 );
and \U$29602 ( \29979 , \29967 , \29976 );
nor \U$29603 ( \29980 , \29978 , \29979 );
not \U$29604 ( \29981 , RIae7aab0_192);
not \U$29605 ( \29982 , RIae7aa38_191);
not \U$29606 ( \29983 , \1185 );
or \U$29607 ( \29984 , \29982 , \29983 );
or \U$29608 ( \29985 , \1186 , RIae7aa38_191);
nand \U$29609 ( \29986 , \29984 , \29985 );
not \U$29610 ( \29987 , \29986 );
or \U$29611 ( \29988 , \29981 , \29987 );
not \U$29612 ( \29989 , \28814 );
nand \U$29613 ( \29990 , \29989 , \14669 );
nand \U$29614 ( \29991 , \29988 , \29990 );
xnor \U$29615 ( \29992 , \29980 , \29991 );
xor \U$29616 ( \29993 , \29958 , \29992 );
not \U$29617 ( \29994 , \16135 );
not \U$29618 ( \29995 , RIae7a2b8_175);
and \U$29619 ( \29996 , \1859 , \29995 );
not \U$29620 ( \29997 , \1859 );
and \U$29621 ( \29998 , \29997 , RIae7a2b8_175);
nor \U$29622 ( \29999 , \29996 , \29998 );
not \U$29623 ( \30000 , \29999 );
or \U$29624 ( \30001 , \29994 , \30000 );
nand \U$29625 ( \30002 , \28549 , \9792 );
nand \U$29626 ( \30003 , \30001 , \30002 );
not \U$29627 ( \30004 , \9776 );
not \U$29628 ( \30005 , \10658 );
not \U$29629 ( \30006 , \2309 );
or \U$29630 ( \30007 , \30005 , \30006 );
nand \U$29631 ( \30008 , \2305 , RIae7a150_172);
nand \U$29632 ( \30009 , \30007 , \30008 );
not \U$29633 ( \30010 , \30009 );
or \U$29634 ( \30011 , \30004 , \30010 );
nand \U$29635 ( \30012 , \28767 , \9758 );
nand \U$29636 ( \30013 , \30011 , \30012 );
not \U$29637 ( \30014 , \30013 );
xor \U$29638 ( \30015 , \30003 , \30014 );
not \U$29639 ( \30016 , \11098 );
not \U$29640 ( \30017 , RIae7a060_170);
not \U$29641 ( \30018 , \19400 );
or \U$29642 ( \30019 , \30017 , \30018 );
or \U$29643 ( \30020 , \2136 , RIae7a060_170);
nand \U$29644 ( \30021 , \30019 , \30020 );
not \U$29645 ( \30022 , \30021 );
or \U$29646 ( \30023 , \30016 , \30022 );
nand \U$29647 ( \30024 , \28719 , \17797 );
nand \U$29648 ( \30025 , \30023 , \30024 );
xnor \U$29649 ( \30026 , \30015 , \30025 );
xnor \U$29650 ( \30027 , \29993 , \30026 );
not \U$29651 ( \30028 , \30027 );
not \U$29652 ( \30029 , \30028 );
or \U$29653 ( \30030 , \29951 , \30029 );
nand \U$29654 ( \30031 , \30027 , \29949 );
nand \U$29655 ( \30032 , \30030 , \30031 );
not \U$29656 ( \30033 , \29776 );
and \U$29657 ( \30034 , \29807 , \29682 );
not \U$29658 ( \30035 , \29807 );
not \U$29659 ( \30036 , \29682 );
and \U$29660 ( \30037 , \30035 , \30036 );
nor \U$29661 ( \30038 , \30034 , \30037 );
not \U$29662 ( \30039 , \30038 );
or \U$29663 ( \30040 , \30033 , \30039 );
nand \U$29664 ( \30041 , \29807 , \29682 );
nand \U$29665 ( \30042 , \30040 , \30041 );
not \U$29666 ( \30043 , \30042 );
xor \U$29667 ( \30044 , \30032 , \30043 );
not \U$29668 ( \30045 , \30044 );
xor \U$29669 ( \30046 , \29863 , \30045 );
xor \U$29670 ( \30047 , \29633 , \29640 );
and \U$29671 ( \30048 , \30047 , \29645 );
and \U$29672 ( \30049 , \29633 , \29640 );
or \U$29673 ( \30050 , \30048 , \30049 );
not \U$29674 ( \30051 , \30050 );
not \U$29675 ( \30052 , \30051 );
not \U$29676 ( \30053 , \29791 );
not \U$29677 ( \30054 , \29802 );
or \U$29678 ( \30055 , \30053 , \30054 );
not \U$29679 ( \30056 , \29787 );
nand \U$29680 ( \30057 , \30056 , \29783 );
nand \U$29681 ( \30058 , \30055 , \30057 );
not \U$29682 ( \30059 , \30058 );
not \U$29683 ( \30060 , \29721 );
not \U$29684 ( \30061 , \29715 );
or \U$29685 ( \30062 , \30060 , \30061 );
nand \U$29686 ( \30063 , \29692 , \29710 );
nand \U$29687 ( \30064 , \30062 , \30063 );
not \U$29688 ( \30065 , \10223 );
xnor \U$29689 ( \30066 , \10065 , RIae79520_146);
not \U$29690 ( \30067 , \30066 );
not \U$29691 ( \30068 , \30067 );
or \U$29692 ( \30069 , \30065 , \30068 );
nand \U$29693 ( \30070 , \29751 , \2602 );
nand \U$29694 ( \30071 , \30069 , \30070 );
not \U$29695 ( \30072 , \30071 );
not \U$29696 ( \30073 , \30072 );
not \U$29697 ( \30074 , \29709 );
not \U$29698 ( \30075 , \29699 );
or \U$29699 ( \30076 , \30074 , \30075 );
nand \U$29700 ( \30077 , \29698 , \29693 );
nand \U$29701 ( \30078 , \30076 , \30077 );
not \U$29702 ( \30079 , \1863 );
not \U$29703 ( \30080 , \1884 );
not \U$29704 ( \30081 , \19689 );
not \U$29705 ( \30082 , \30081 );
or \U$29706 ( \30083 , \30080 , \30082 );
nand \U$29707 ( \30084 , \11577 , RIae793b8_143);
nand \U$29708 ( \30085 , \30083 , \30084 );
not \U$29709 ( \30086 , \30085 );
or \U$29710 ( \30087 , \30079 , \30086 );
nand \U$29711 ( \30088 , \29705 , \1910 );
nand \U$29712 ( \30089 , \30087 , \30088 );
xor \U$29713 ( \30090 , \30078 , \30089 );
not \U$29714 ( \30091 , \30090 );
or \U$29715 ( \30092 , \30073 , \30091 );
or \U$29716 ( \30093 , \30090 , \30072 );
nand \U$29717 ( \30094 , \30092 , \30093 );
xor \U$29718 ( \30095 , \30064 , \30094 );
buf \U$29719 ( \30096 , \30095 );
not \U$29720 ( \30097 , \29757 );
not \U$29721 ( \30098 , \29731 );
or \U$29722 ( \30099 , \30097 , \30098 );
not \U$29723 ( \30100 , \29742 );
nand \U$29724 ( \30101 , \30100 , \29753 );
nand \U$29725 ( \30102 , \30099 , \30101 );
not \U$29726 ( \30103 , \30102 );
and \U$29727 ( \30104 , \30096 , \30103 );
not \U$29728 ( \30105 , \30096 );
and \U$29729 ( \30106 , \30105 , \30102 );
nor \U$29730 ( \30107 , \30104 , \30106 );
not \U$29731 ( \30108 , \30107 );
and \U$29732 ( \30109 , \30059 , \30108 );
and \U$29733 ( \30110 , \30107 , \30058 );
nor \U$29734 ( \30111 , \30109 , \30110 );
not \U$29735 ( \30112 , \1820 );
and \U$29736 ( \30113 , RIae79688_149, \16194 );
not \U$29737 ( \30114 , RIae79688_149);
and \U$29738 ( \30115 , \30114 , \10740 );
nor \U$29739 ( \30116 , \30113 , \30115 );
not \U$29740 ( \30117 , \30116 );
or \U$29741 ( \30118 , \30112 , \30117 );
nand \U$29742 ( \30119 , \28755 , \1843 );
nand \U$29743 ( \30120 , \30118 , \30119 );
not \U$29744 ( \30121 , \2249 );
not \U$29745 ( \30122 , RIae79ac0_158);
not \U$29746 ( \30123 , \10749 );
or \U$29747 ( \30124 , \30122 , \30123 );
or \U$29748 ( \30125 , \9875 , RIae79ac0_158);
nand \U$29749 ( \30126 , \30124 , \30125 );
not \U$29750 ( \30127 , \30126 );
or \U$29751 ( \30128 , \30121 , \30127 );
nand \U$29752 ( \30129 , \29740 , \2272 );
nand \U$29753 ( \30130 , \30128 , \30129 );
xor \U$29754 ( \30131 , \30120 , \30130 );
not \U$29755 ( \30132 , \1919 );
not \U$29756 ( \30133 , \3810 );
not \U$29757 ( \30134 , \28019 );
or \U$29758 ( \30135 , \30133 , \30134 );
or \U$29759 ( \30136 , \28019 , \3039 );
nand \U$29760 ( \30137 , \30135 , \30136 );
not \U$29761 ( \30138 , \30137 );
or \U$29762 ( \30139 , \30132 , \30138 );
nand \U$29763 ( \30140 , \29690 , \1932 );
nand \U$29764 ( \30141 , \30139 , \30140 );
not \U$29765 ( \30142 , \30141 );
xor \U$29766 ( \30143 , \30131 , \30142 );
not \U$29767 ( \30144 , \30143 );
not \U$29768 ( \30145 , \28540 );
not \U$29769 ( \30146 , \28551 );
or \U$29770 ( \30147 , \30145 , \30146 );
nand \U$29771 ( \30148 , \28534 , \28527 );
nand \U$29772 ( \30149 , \30147 , \30148 );
xor \U$29773 ( \30150 , \30144 , \30149 );
xor \U$29774 ( \30151 , \28566 , \28576 );
and \U$29775 ( \30152 , \30151 , \28586 );
and \U$29776 ( \30153 , \28566 , \28576 );
or \U$29777 ( \30154 , \30152 , \30153 );
buf \U$29778 ( \30155 , \30154 );
xnor \U$29779 ( \30156 , \30150 , \30155 );
and \U$29780 ( \30157 , \30111 , \30156 );
not \U$29781 ( \30158 , \30111 );
not \U$29782 ( \30159 , \30156 );
and \U$29783 ( \30160 , \30158 , \30159 );
nor \U$29784 ( \30161 , \30157 , \30160 );
not \U$29785 ( \30162 , \30161 );
or \U$29786 ( \30163 , \30052 , \30162 );
or \U$29787 ( \30164 , \30161 , \30051 );
nand \U$29788 ( \30165 , \30163 , \30164 );
not \U$29789 ( \30166 , \30165 );
and \U$29790 ( \30167 , \29770 , \29763 );
and \U$29791 ( \30168 , \29726 , \29762 );
nor \U$29792 ( \30169 , \30167 , \30168 );
not \U$29793 ( \30170 , \28773 );
not \U$29794 ( \30171 , \28735 );
or \U$29795 ( \30172 , \30170 , \30171 );
not \U$29796 ( \30173 , \28758 );
nand \U$29797 ( \30174 , \30173 , \28769 );
nand \U$29798 ( \30175 , \30172 , \30174 );
not \U$29799 ( \30176 , \28723 );
not \U$29800 ( \30177 , \30176 );
not \U$29801 ( \30178 , \28713 );
or \U$29802 ( \30179 , \30177 , \30178 );
nand \U$29803 ( \30180 , \28711 , \28695 , \28698 );
nand \U$29804 ( \30181 , \30179 , \30180 );
xor \U$29805 ( \30182 , \30175 , \30181 );
xor \U$29806 ( \30183 , \28785 , \28796 );
and \U$29807 ( \30184 , \30183 , \28807 );
and \U$29808 ( \30185 , \28785 , \28796 );
or \U$29809 ( \30186 , \30184 , \30185 );
xnor \U$29810 ( \30187 , \30182 , \30186 );
xor \U$29811 ( \30188 , \30169 , \30187 );
not \U$29812 ( \30189 , \28853 );
not \U$29813 ( \30190 , \28842 );
or \U$29814 ( \30191 , \30189 , \30190 );
not \U$29815 ( \30192 , \28834 );
nand \U$29816 ( \30193 , \30192 , \28817 );
not \U$29817 ( \30194 , \30193 );
nand \U$29818 ( \30195 , \28834 , \28818 );
not \U$29819 ( \30196 , \30195 );
or \U$29820 ( \30197 , \30194 , \30196 );
nand \U$29821 ( \30198 , \30197 , \28841 );
nand \U$29822 ( \30199 , \30191 , \30198 );
not \U$29823 ( \30200 , \30199 );
xnor \U$29824 ( \30201 , \30188 , \30200 );
not \U$29825 ( \30202 , \30201 );
not \U$29826 ( \30203 , \30202 );
not \U$29827 ( \30204 , \30203 );
or \U$29828 ( \30205 , \30166 , \30204 );
or \U$29829 ( \30206 , \30203 , \30165 );
nand \U$29830 ( \30207 , \30205 , \30206 );
xnor \U$29831 ( \30208 , \30046 , \30207 );
not \U$29832 ( \30209 , \30208 );
not \U$29833 ( \30210 , \30209 );
not \U$29834 ( \30211 , \28185 );
not \U$29835 ( \30212 , \28680 );
not \U$29836 ( \30213 , \30212 );
or \U$29837 ( \30214 , \30211 , \30213 );
not \U$29838 ( \30215 , \28185 );
nand \U$29839 ( \30216 , \30215 , \28680 );
nand \U$29840 ( \30217 , \30214 , \30216 );
not \U$29841 ( \30218 , \30217 );
and \U$29842 ( \30219 , \27669 , \27857 );
not \U$29843 ( \30220 , \27669 );
not \U$29844 ( \30221 , \27857 );
and \U$29845 ( \30222 , \30220 , \30221 );
nor \U$29846 ( \30223 , \30219 , \30222 );
not \U$29847 ( \30224 , \30223 );
not \U$29848 ( \30225 , \27961 );
not \U$29849 ( \30226 , \30225 );
not \U$29850 ( \30227 , \28055 );
or \U$29851 ( \30228 , \30226 , \30227 );
or \U$29852 ( \30229 , \28055 , \30225 );
nand \U$29853 ( \30230 , \30228 , \30229 );
xor \U$29854 ( \30231 , \29328 , \29333 );
xor \U$29855 ( \30232 , \30231 , \29344 );
nor \U$29856 ( \30233 , \30230 , \30232 );
xnor \U$29857 ( \30234 , \27940 , \27910 );
or \U$29858 ( \30235 , \30233 , \30234 );
nand \U$29859 ( \30236 , \30230 , \30232 );
nand \U$29860 ( \30237 , \30235 , \30236 );
buf \U$29861 ( \30238 , \30237 );
xor \U$29862 ( \30239 , \29819 , \29829 );
xor \U$29863 ( \30240 , \30239 , \29824 );
not \U$29864 ( \30241 , \30240 );
xor \U$29865 ( \30242 , \30238 , \30241 );
not \U$29866 ( \30243 , \30242 );
or \U$29867 ( \30244 , \30224 , \30243 );
not \U$29868 ( \30245 , \30240 );
and \U$29869 ( \30246 , \30238 , \30245 );
not \U$29870 ( \30247 , \30246 );
nand \U$29871 ( \30248 , \30244 , \30247 );
not \U$29872 ( \30249 , \30248 );
and \U$29873 ( \30250 , \29814 , \29841 );
not \U$29874 ( \30251 , \29814 );
and \U$29875 ( \30252 , \30251 , \29816 );
nor \U$29876 ( \30253 , \30250 , \30252 );
xor \U$29877 ( \30254 , \29838 , \30253 );
not \U$29878 ( \30255 , \30254 );
xor \U$29879 ( \30256 , \28351 , \28442 );
xor \U$29880 ( \30257 , \30256 , \28516 );
not \U$29881 ( \30258 , \30257 );
not \U$29882 ( \30259 , \30258 );
or \U$29883 ( \30260 , \30255 , \30259 );
not \U$29884 ( \30261 , \30254 );
nand \U$29885 ( \30262 , \30261 , \30257 );
nand \U$29886 ( \30263 , \30260 , \30262 );
not \U$29887 ( \30264 , \30263 );
or \U$29888 ( \30265 , \30249 , \30264 );
not \U$29889 ( \30266 , \30254 );
nand \U$29890 ( \30267 , \30266 , \30258 );
nand \U$29891 ( \30268 , \30265 , \30267 );
not \U$29892 ( \30269 , \30268 );
not \U$29893 ( \30270 , \30269 );
or \U$29894 ( \30271 , \30218 , \30270 );
xor \U$29895 ( \30272 , \29271 , \29251 );
xor \U$29896 ( \30273 , \30272 , \29265 );
not \U$29897 ( \30274 , \1919 );
not \U$29898 ( \30275 , \27995 );
or \U$29899 ( \30276 , \30274 , \30275 );
not \U$29900 ( \30277 , RIae794a8_145);
not \U$29901 ( \30278 , \10149 );
or \U$29902 ( \30279 , \30277 , \30278 );
or \U$29903 ( \30280 , \10149 , RIae794a8_145);
nand \U$29904 ( \30281 , \30279 , \30280 );
nand \U$29905 ( \30282 , \30281 , \2457 );
nand \U$29906 ( \30283 , \30276 , \30282 );
not \U$29907 ( \30284 , \2007 );
not \U$29908 ( \30285 , \29267 );
or \U$29909 ( \30286 , \30284 , \30285 );
not \U$29910 ( \30287 , \9896 );
xor \U$29911 ( \30288 , RIae797f0_152, \30287 );
nand \U$29912 ( \30289 , \30288 , \1988 );
nand \U$29913 ( \30290 , \30286 , \30289 );
xor \U$29914 ( \30291 , \30283 , \30290 );
not \U$29915 ( \30292 , \15337 );
not \U$29916 ( \30293 , \29257 );
or \U$29917 ( \30294 , \30292 , \30293 );
not \U$29918 ( \30295 , \2447 );
not \U$29919 ( \30296 , \11386 );
or \U$29920 ( \30297 , \30295 , \30296 );
or \U$29921 ( \30298 , \15650 , \2447 );
nand \U$29922 ( \30299 , \30297 , \30298 );
nand \U$29923 ( \30300 , \30299 , \2431 );
nand \U$29924 ( \30301 , \30294 , \30300 );
and \U$29925 ( \30302 , \30291 , \30301 );
and \U$29926 ( \30303 , \30283 , \30290 );
or \U$29927 ( \30304 , \30302 , \30303 );
or \U$29928 ( \30305 , \30273 , \30304 );
not \U$29929 ( \30306 , \10573 );
not \U$29930 ( \30307 , \27734 );
or \U$29931 ( \30308 , \30306 , \30307 );
not \U$29932 ( \30309 , \6203 );
not \U$29933 ( \30310 , \9367 );
or \U$29934 ( \30311 , \30309 , \30310 );
or \U$29935 ( \30312 , \9367 , \9560 );
nand \U$29936 ( \30313 , \30311 , \30312 );
nand \U$29937 ( \30314 , \30313 , \11409 );
nand \U$29938 ( \30315 , \30308 , \30314 );
not \U$29939 ( \30316 , \30315 );
not \U$29940 ( \30317 , \5049 );
not \U$29941 ( \30318 , \29300 );
or \U$29942 ( \30319 , \30317 , \30318 );
xnor \U$29943 ( \30320 , \10361 , RIae79d90_164);
nand \U$29944 ( \30321 , \30320 , \6091 );
nand \U$29945 ( \30322 , \30319 , \30321 );
not \U$29946 ( \30323 , \30322 );
not \U$29947 ( \30324 , \29404 );
or \U$29948 ( \30325 , \30324 , \1819 );
and \U$29949 ( \30326 , RIae79688_149, \14601 );
not \U$29950 ( \30327 , RIae79688_149);
and \U$29951 ( \30328 , \30327 , \12857 );
nor \U$29952 ( \30329 , \30326 , \30328 );
not \U$29953 ( \30330 , \1842 );
or \U$29954 ( \30331 , \30329 , \30330 );
nand \U$29955 ( \30332 , \30325 , \30331 );
not \U$29956 ( \30333 , \30332 );
or \U$29957 ( \30334 , \10419 , \1816 );
not \U$29958 ( \30335 , \1816 );
not \U$29959 ( \30336 , \2268 );
or \U$29960 ( \30337 , \30335 , \30336 );
nand \U$29961 ( \30338 , \30337 , \12857 );
nand \U$29962 ( \30339 , \30334 , \30338 , RIae79688_149);
nor \U$29963 ( \30340 , \30333 , \30339 );
not \U$29964 ( \30341 , \1932 );
and \U$29965 ( \30342 , RIae794a8_145, \10031 );
not \U$29966 ( \30343 , RIae794a8_145);
and \U$29967 ( \30344 , \30343 , \10337 );
nor \U$29968 ( \30345 , \30342 , \30344 );
not \U$29969 ( \30346 , \30345 );
or \U$29970 ( \30347 , \30341 , \30346 );
nand \U$29971 ( \30348 , \30281 , \1919 );
nand \U$29972 ( \30349 , \30347 , \30348 );
xor \U$29973 ( \30350 , \30340 , \30349 );
not \U$29974 ( \30351 , \2162 );
not \U$29975 ( \30352 , \27791 );
or \U$29976 ( \30353 , \30351 , \30352 );
and \U$29977 ( \30354 , RIae79520_146, \10193 );
not \U$29978 ( \30355 , RIae79520_146);
and \U$29979 ( \30356 , \30355 , \10194 );
nor \U$29980 ( \30357 , \30354 , \30356 );
nand \U$29981 ( \30358 , \30357 , \2188 );
nand \U$29982 ( \30359 , \30353 , \30358 );
and \U$29983 ( \30360 , \30350 , \30359 );
and \U$29984 ( \30361 , \30340 , \30349 );
or \U$29985 ( \30362 , \30360 , \30361 );
not \U$29986 ( \30363 , \30362 );
not \U$29987 ( \30364 , \30363 );
or \U$29988 ( \30365 , \30323 , \30364 );
or \U$29989 ( \30366 , \30322 , \30363 );
nand \U$29990 ( \30367 , \30365 , \30366 );
not \U$29991 ( \30368 , \30367 );
or \U$29992 ( \30369 , \30316 , \30368 );
not \U$29993 ( \30370 , \30363 );
nand \U$29994 ( \30371 , \30370 , \30322 );
nand \U$29995 ( \30372 , \30369 , \30371 );
nand \U$29996 ( \30373 , \30305 , \30372 );
nand \U$29997 ( \30374 , \30273 , \30304 );
nand \U$29998 ( \30375 , \30373 , \30374 );
not \U$29999 ( \30376 , \30375 );
not \U$30000 ( \30377 , \30376 );
not \U$30001 ( \30378 , \16358 );
not \U$30002 ( \30379 , \29311 );
or \U$30003 ( \30380 , \30378 , \30379 );
and \U$30004 ( \30381 , RIae7a510_180, \2402 );
not \U$30005 ( \30382 , RIae7a510_180);
and \U$30006 ( \30383 , \30382 , \3269 );
or \U$30007 ( \30384 , \30381 , \30383 );
nand \U$30008 ( \30385 , \30384 , \11400 );
nand \U$30009 ( \30386 , \30380 , \30385 );
not \U$30010 ( \30387 , \4853 );
not \U$30011 ( \30388 , \29288 );
or \U$30012 ( \30389 , \30387 , \30388 );
and \U$30013 ( \30390 , RIae79ca0_162, \9416 );
not \U$30014 ( \30391 , RIae79ca0_162);
and \U$30015 ( \30392 , \30391 , \9412 );
or \U$30016 ( \30393 , \30390 , \30392 );
not \U$30017 ( \30394 , \30393 );
nand \U$30018 ( \30395 , \30394 , \4154 );
nand \U$30019 ( \30396 , \30389 , \30395 );
xor \U$30020 ( \30397 , \30386 , \30396 );
not \U$30021 ( \30398 , \30397 );
not \U$30022 ( \30399 , \10275 );
not \U$30023 ( \30400 , \29505 );
or \U$30024 ( \30401 , \30399 , \30400 );
and \U$30025 ( \30402 , RIae7a8d0_188, \2154 );
not \U$30026 ( \30403 , RIae7a8d0_188);
and \U$30027 ( \30404 , \30403 , \13142 );
nor \U$30028 ( \30405 , \30402 , \30404 );
nand \U$30029 ( \30406 , \30405 , \11205 );
nand \U$30030 ( \30407 , \30401 , \30406 );
not \U$30031 ( \30408 , \30407 );
or \U$30032 ( \30409 , \30398 , \30408 );
nand \U$30033 ( \30410 , \30396 , \30386 );
nand \U$30034 ( \30411 , \30409 , \30410 );
not \U$30035 ( \30412 , \30411 );
not \U$30036 ( \30413 , \9527 );
not \U$30037 ( \30414 , \29515 );
or \U$30038 ( \30415 , \30413 , \30414 );
not \U$30039 ( \30416 , \10608 );
and \U$30040 ( \30417 , RIae7a7e0_186, \30416 );
not \U$30041 ( \30418 , RIae7a7e0_186);
and \U$30042 ( \30419 , \30418 , \10905 );
nor \U$30043 ( \30420 , \30417 , \30419 );
nand \U$30044 ( \30421 , \30420 , \9549 );
nand \U$30045 ( \30422 , \30415 , \30421 );
not \U$30046 ( \30423 , \9744 );
not \U$30047 ( \30424 , \29527 );
or \U$30048 ( \30425 , \30423 , \30424 );
not \U$30049 ( \30426 , RIae7a060_170);
not \U$30050 ( \30427 , \1789 );
or \U$30051 ( \30428 , \30426 , \30427 );
or \U$30052 ( \30429 , \28790 , RIae7a060_170);
nand \U$30053 ( \30430 , \30428 , \30429 );
nand \U$30054 ( \30431 , \30430 , \9730 );
nand \U$30055 ( \30432 , \30425 , \30431 );
xor \U$30056 ( \30433 , \30422 , \30432 );
not \U$30057 ( \30434 , RIae7aab0_192);
not \U$30058 ( \30435 , \29232 );
or \U$30059 ( \30436 , \30434 , \30435 );
not \U$30060 ( \30437 , \11326 );
not \U$30061 ( \30438 , \18384 );
or \U$30062 ( \30439 , \30437 , \30438 );
nand \U$30063 ( \30440 , \2230 , RIae7aa38_191);
nand \U$30064 ( \30441 , \30439 , \30440 );
nand \U$30065 ( \30442 , \30441 , \14667 );
nand \U$30066 ( \30443 , \30436 , \30442 );
and \U$30067 ( \30444 , \30433 , \30443 );
and \U$30068 ( \30445 , \30422 , \30432 );
or \U$30069 ( \30446 , \30444 , \30445 );
not \U$30070 ( \30447 , \30446 );
nand \U$30071 ( \30448 , \30412 , \30447 );
not \U$30072 ( \30449 , \9776 );
not \U$30073 ( \30450 , \29223 );
or \U$30074 ( \30451 , \30449 , \30450 );
not \U$30075 ( \30452 , \14907 );
not \U$30076 ( \30453 , RIae7a150_172);
and \U$30077 ( \30454 , \30452 , \30453 );
and \U$30078 ( \30455 , \2093 , RIae7a150_172);
nor \U$30079 ( \30456 , \30454 , \30455 );
nand \U$30080 ( \30457 , \30456 , \11087 );
nand \U$30081 ( \30458 , \30451 , \30457 );
not \U$30082 ( \30459 , \9473 );
and \U$30083 ( \30460 , \3748 , RIae7a6f0_184);
not \U$30084 ( \30461 , \3748 );
and \U$30085 ( \30462 , \30461 , \16101 );
nor \U$30086 ( \30463 , \30460 , \30462 );
not \U$30087 ( \30464 , \30463 );
or \U$30088 ( \30465 , \30459 , \30464 );
nand \U$30089 ( \30466 , \29433 , \9478 );
nand \U$30090 ( \30467 , \30465 , \30466 );
nor \U$30091 ( \30468 , \30458 , \30467 );
and \U$30092 ( \30469 , \12371 , \29364 );
and \U$30093 ( \30470 , \1970 , \10625 );
not \U$30094 ( \30471 , \1970 );
and \U$30095 ( \30472 , \30471 , RIae7a498_179);
nor \U$30096 ( \30473 , \30470 , \30472 );
and \U$30097 ( \30474 , \30473 , \11434 );
nor \U$30098 ( \30475 , \30469 , \30474 );
or \U$30099 ( \30476 , \30468 , \30475 );
nand \U$30100 ( \30477 , \30458 , \30467 );
nand \U$30101 ( \30478 , \30476 , \30477 );
and \U$30102 ( \30479 , \30448 , \30478 );
nand \U$30103 ( \30480 , \30411 , \30446 );
not \U$30104 ( \30481 , \30480 );
nor \U$30105 ( \30482 , \30479 , \30481 );
not \U$30106 ( \30483 , \30482 );
not \U$30107 ( \30484 , \30483 );
not \U$30108 ( \30485 , \30484 );
or \U$30109 ( \30486 , \30377 , \30485 );
not \U$30110 ( \30487 , \30375 );
not \U$30111 ( \30488 , \30483 );
or \U$30112 ( \30489 , \30487 , \30488 );
xor \U$30113 ( \30490 , \27793 , \27777 );
not \U$30114 ( \30491 , \16135 );
not \U$30115 ( \30492 , \27837 );
or \U$30116 ( \30493 , \30491 , \30492 );
xor \U$30117 ( \30494 , RIae7a2b8_175, \9289 );
nand \U$30118 ( \30495 , \30494 , \9792 );
nand \U$30119 ( \30496 , \30493 , \30495 );
xor \U$30120 ( \30497 , \30490 , \30496 );
not \U$30121 ( \30498 , \10700 );
not \U$30122 ( \30499 , \27719 );
or \U$30123 ( \30500 , \30498 , \30499 );
and \U$30124 ( \30501 , RIae79fe8_169, \9316 );
not \U$30125 ( \30502 , RIae79fe8_169);
and \U$30126 ( \30503 , \30502 , \14644 );
or \U$30127 ( \30504 , \30501 , \30503 );
nand \U$30128 ( \30505 , \30504 , \11914 );
nand \U$30129 ( \30506 , \30500 , \30505 );
and \U$30130 ( \30507 , \30497 , \30506 );
and \U$30131 ( \30508 , \30490 , \30496 );
nor \U$30132 ( \30509 , \30507 , \30508 );
not \U$30133 ( \30510 , \30509 );
not \U$30134 ( \30511 , \30510 );
not \U$30135 ( \30512 , \2776 );
not \U$30136 ( \30513 , \29249 );
or \U$30137 ( \30514 , \30512 , \30513 );
not \U$30138 ( \30515 , \16837 );
not \U$30139 ( \30516 , RIae79c28_161);
and \U$30140 ( \30517 , \30515 , \30516 );
and \U$30141 ( \30518 , \11186 , RIae79c28_161);
nor \U$30142 ( \30519 , \30517 , \30518 );
nand \U$30143 ( \30520 , \30519 , \2417 );
nand \U$30144 ( \30521 , \30514 , \30520 );
not \U$30145 ( \30522 , \9621 );
not \U$30146 ( \30523 , \27814 );
or \U$30147 ( \30524 , \30522 , \30523 );
nor \U$30148 ( \30525 , \4168 , \13165 );
not \U$30149 ( \30526 , \30525 );
nand \U$30150 ( \30527 , \4168 , \11690 );
nand \U$30151 ( \30528 , \30526 , \30527 );
nand \U$30152 ( \30529 , \30528 , \9644 );
nand \U$30153 ( \30530 , \30524 , \30529 );
xor \U$30154 ( \30531 , \30521 , \30530 );
not \U$30155 ( \30532 , \9699 );
or \U$30156 ( \30533 , \27847 , \30532 );
xor \U$30157 ( \30534 , RIae7a240_174, \5107 );
nand \U$30158 ( \30535 , \30534 , \19466 );
nand \U$30159 ( \30536 , \30533 , \30535 );
and \U$30160 ( \30537 , \30531 , \30536 );
and \U$30161 ( \30538 , \30521 , \30530 );
or \U$30162 ( \30539 , \30537 , \30538 );
not \U$30163 ( \30540 , \30539 );
xnor \U$30164 ( \30541 , \28000 , \28006 );
and \U$30165 ( \30542 , \30540 , \30541 );
not \U$30166 ( \30543 , \30540 );
not \U$30167 ( \30544 , \30541 );
and \U$30168 ( \30545 , \30543 , \30544 );
nor \U$30169 ( \30546 , \30542 , \30545 );
not \U$30170 ( \30547 , \30546 );
or \U$30171 ( \30548 , \30511 , \30547 );
nand \U$30172 ( \30549 , \30539 , \30544 );
nand \U$30173 ( \30550 , \30548 , \30549 );
not \U$30174 ( \30551 , \30550 );
nand \U$30175 ( \30552 , \30489 , \30551 );
nand \U$30176 ( \30553 , \30486 , \30552 );
xnor \U$30177 ( \30554 , \28060 , \27946 );
and \U$30178 ( \30555 , \30554 , \27895 );
not \U$30179 ( \30556 , \30554 );
and \U$30180 ( \30557 , \30556 , \27894 );
nor \U$30181 ( \30558 , \30555 , \30557 );
nand \U$30182 ( \30559 , \30553 , \30558 );
not \U$30183 ( \30560 , \30559 );
xor \U$30184 ( \30561 , \29559 , \29548 );
not \U$30185 ( \30562 , \30561 );
or \U$30186 ( \30563 , \30560 , \30562 );
or \U$30187 ( \30564 , \30553 , \30558 );
nand \U$30188 ( \30565 , \30563 , \30564 );
not \U$30189 ( \30566 , \30565 );
not \U$30190 ( \30567 , \28065 );
nand \U$30191 ( \30568 , \30567 , \28071 );
xor \U$30192 ( \30569 , \30568 , \28183 );
not \U$30193 ( \30570 , \30569 );
nand \U$30194 ( \30571 , \30566 , \30570 );
not \U$30195 ( \30572 , \30571 );
xor \U$30196 ( \30573 , \29498 , \29490 );
xnor \U$30197 ( \30574 , \30573 , \29565 );
not \U$30198 ( \30575 , \30574 );
or \U$30199 ( \30576 , \30572 , \30575 );
nand \U$30200 ( \30577 , \30565 , \30569 );
nand \U$30201 ( \30578 , \30576 , \30577 );
nand \U$30202 ( \30579 , \30271 , \30578 );
not \U$30203 ( \30580 , \30217 );
nand \U$30204 ( \30581 , \30580 , \30268 );
and \U$30205 ( \30582 , \30579 , \30581 );
not \U$30206 ( \30583 , \30582 );
or \U$30207 ( \30584 , \30210 , \30583 );
not \U$30208 ( \30585 , \30579 );
not \U$30209 ( \30586 , \30581 );
or \U$30210 ( \30587 , \30585 , \30586 );
nand \U$30211 ( \30588 , \30587 , \30208 );
nand \U$30212 ( \30589 , \30584 , \30588 );
not \U$30213 ( \30590 , \30589 );
or \U$30214 ( \30591 , \29857 , \30590 );
or \U$30215 ( \30592 , \30589 , \29856 );
nand \U$30216 ( \30593 , \30591 , \30592 );
xor \U$30217 ( \30594 , \30375 , \30550 );
xnor \U$30218 ( \30595 , \30594 , \30482 );
not \U$30219 ( \30596 , \30595 );
xor \U$30220 ( \30597 , \29444 , \29461 );
xor \U$30221 ( \30598 , \30597 , \29484 );
xor \U$30222 ( \30599 , \30283 , \30290 );
xor \U$30223 ( \30600 , \30599 , \30301 );
not \U$30224 ( \30601 , \30600 );
not \U$30225 ( \30602 , \29418 );
not \U$30226 ( \30603 , \29378 );
not \U$30227 ( \30604 , \30603 );
or \U$30228 ( \30605 , \30602 , \30604 );
or \U$30229 ( \30606 , \30603 , \29418 );
nand \U$30230 ( \30607 , \30605 , \30606 );
not \U$30231 ( \30608 , \2321 );
not \U$30232 ( \30609 , \29376 );
or \U$30233 ( \30610 , \30608 , \30609 );
not \U$30234 ( \30611 , \5344 );
not \U$30235 ( \30612 , \16194 );
or \U$30236 ( \30613 , \30611 , \30612 );
or \U$30237 ( \30614 , \27671 , \2334 );
nand \U$30238 ( \30615 , \30613 , \30614 );
nand \U$30239 ( \30616 , \30615 , \2339 );
nand \U$30240 ( \30617 , \30610 , \30616 );
not \U$30241 ( \30618 , \30617 );
not \U$30242 ( \30619 , \29396 );
not \U$30243 ( \30620 , \30619 );
not \U$30244 ( \30621 , \29413 );
and \U$30245 ( \30622 , \30620 , \30621 );
and \U$30246 ( \30623 , \29413 , \30619 );
nor \U$30247 ( \30624 , \30622 , \30623 );
not \U$30248 ( \30625 , \30624 );
not \U$30249 ( \30626 , \1988 );
xor \U$30250 ( \30627 , RIae797f0_152, \9867 );
not \U$30251 ( \30628 , \30627 );
or \U$30252 ( \30629 , \30626 , \30628 );
not \U$30253 ( \30630 , \2518 );
nand \U$30254 ( \30631 , \30630 , \30288 );
nand \U$30255 ( \30632 , \30629 , \30631 );
not \U$30256 ( \30633 , \30632 );
or \U$30257 ( \30634 , \30625 , \30633 );
or \U$30258 ( \30635 , \30632 , \30624 );
nand \U$30259 ( \30636 , \30634 , \30635 );
not \U$30260 ( \30637 , \30636 );
or \U$30261 ( \30638 , \30618 , \30637 );
not \U$30262 ( \30639 , \30624 );
nand \U$30263 ( \30640 , \30639 , \30632 );
nand \U$30264 ( \30641 , \30638 , \30640 );
xor \U$30265 ( \30642 , \30607 , \30641 );
not \U$30266 ( \30643 , \30642 );
or \U$30267 ( \30644 , \30601 , \30643 );
nand \U$30268 ( \30645 , \30641 , \30607 );
nand \U$30269 ( \30646 , \30644 , \30645 );
not \U$30270 ( \30647 , \30646 );
not \U$30271 ( \30648 , \30647 );
not \U$30272 ( \30649 , \6200 );
not \U$30273 ( \30650 , \6207 );
not \U$30274 ( \30651 , \9441 );
or \U$30275 ( \30652 , \30650 , \30651 );
or \U$30276 ( \30653 , \9441 , \13733 );
nand \U$30277 ( \30654 , \30652 , \30653 );
not \U$30278 ( \30655 , \30654 );
or \U$30279 ( \30656 , \30649 , \30655 );
nand \U$30280 ( \30657 , \30313 , \6212 );
nand \U$30281 ( \30658 , \30656 , \30657 );
not \U$30282 ( \30659 , \30658 );
not \U$30283 ( \30660 , \30332 );
not \U$30284 ( \30661 , \30339 );
and \U$30285 ( \30662 , \30660 , \30661 );
and \U$30286 ( \30663 , \30332 , \30339 );
nor \U$30287 ( \30664 , \30662 , \30663 );
not \U$30288 ( \30665 , \30664 );
not \U$30289 ( \30666 , \2249 );
not \U$30290 ( \30667 , \29394 );
or \U$30291 ( \30668 , \30666 , \30667 );
not \U$30292 ( \30669 , RIae79ac0_158);
not \U$30293 ( \30670 , \16165 );
or \U$30294 ( \30671 , \30669 , \30670 );
or \U$30295 ( \30672 , \17166 , RIae79ac0_158);
nand \U$30296 ( \30673 , \30671 , \30672 );
nand \U$30297 ( \30674 , \30673 , \2272 );
nand \U$30298 ( \30675 , \30668 , \30674 );
not \U$30299 ( \30676 , \30675 );
or \U$30300 ( \30677 , \30665 , \30676 );
or \U$30301 ( \30678 , \30675 , \30664 );
nand \U$30302 ( \30679 , \30677 , \30678 );
not \U$30303 ( \30680 , \30679 );
not \U$30304 ( \30681 , \1932 );
not \U$30305 ( \30682 , \3810 );
not \U$30306 ( \30683 , \11665 );
or \U$30307 ( \30684 , \30682 , \30683 );
or \U$30308 ( \30685 , \10047 , \3039 );
nand \U$30309 ( \30686 , \30684 , \30685 );
not \U$30310 ( \30687 , \30686 );
or \U$30311 ( \30688 , \30681 , \30687 );
nand \U$30312 ( \30689 , \30345 , \1919 );
nand \U$30313 ( \30690 , \30688 , \30689 );
not \U$30314 ( \30691 , \30690 );
or \U$30315 ( \30692 , \30680 , \30691 );
not \U$30316 ( \30693 , \30664 );
nand \U$30317 ( \30694 , \30693 , \30675 );
nand \U$30318 ( \30695 , \30692 , \30694 );
not \U$30319 ( \30696 , \30695 );
not \U$30320 ( \30697 , \30696 );
or \U$30321 ( \30698 , \30659 , \30697 );
or \U$30322 ( \30699 , \30658 , \30696 );
nand \U$30323 ( \30700 , \30698 , \30699 );
not \U$30324 ( \30701 , \30700 );
not \U$30325 ( \30702 , \11913 );
not \U$30326 ( \30703 , RIae79fe8_169);
not \U$30327 ( \30704 , \12707 );
or \U$30328 ( \30705 , \30703 , \30704 );
or \U$30329 ( \30706 , \24816 , RIae79fe8_169);
nand \U$30330 ( \30707 , \30705 , \30706 );
not \U$30331 ( \30708 , \30707 );
or \U$30332 ( \30709 , \30702 , \30708 );
nand \U$30333 ( \30710 , \30504 , \9517 );
nand \U$30334 ( \30711 , \30709 , \30710 );
not \U$30335 ( \30712 , \30711 );
or \U$30336 ( \30713 , \30701 , \30712 );
nand \U$30337 ( \30714 , \30658 , \30695 );
nand \U$30338 ( \30715 , \30713 , \30714 );
not \U$30339 ( \30716 , \2432 );
and \U$30340 ( \30717 , RIae79778_151, \10067 );
not \U$30341 ( \30718 , RIae79778_151);
and \U$30342 ( \30719 , \30718 , \10070 );
or \U$30343 ( \30720 , \30717 , \30719 );
not \U$30344 ( \30721 , \30720 );
or \U$30345 ( \30722 , \30716 , \30721 );
nand \U$30346 ( \30723 , \30299 , \15337 );
nand \U$30347 ( \30724 , \30722 , \30723 );
not \U$30348 ( \30725 , \30724 );
not \U$30349 ( \30726 , \2417 );
not \U$30350 ( \30727 , \10584 );
not \U$30351 ( \30728 , \28019 );
or \U$30352 ( \30729 , \30727 , \30728 );
or \U$30353 ( \30730 , \28019 , \10584 );
nand \U$30354 ( \30731 , \30729 , \30730 );
not \U$30355 ( \30732 , \30731 );
or \U$30356 ( \30733 , \30726 , \30732 );
nand \U$30357 ( \30734 , \30519 , \2418 );
nand \U$30358 ( \30735 , \30733 , \30734 );
not \U$30359 ( \30736 , \30735 );
not \U$30360 ( \30737 , \30736 );
or \U$30361 ( \30738 , \30725 , \30737 );
or \U$30362 ( \30739 , \30736 , \30724 );
nand \U$30363 ( \30740 , \30738 , \30739 );
not \U$30364 ( \30741 , \30740 );
not \U$30365 ( \30742 , \11014 );
and \U$30366 ( \30743 , RIae7a3a8_177, \13985 );
not \U$30367 ( \30744 , RIae7a3a8_177);
and \U$30368 ( \30745 , \30744 , \10829 );
nor \U$30369 ( \30746 , \30743 , \30745 );
not \U$30370 ( \30747 , \30746 );
or \U$30371 ( \30748 , \30742 , \30747 );
nand \U$30372 ( \30749 , \30528 , \9622 );
nand \U$30373 ( \30750 , \30748 , \30749 );
not \U$30374 ( \30751 , \30750 );
or \U$30375 ( \30752 , \30741 , \30751 );
nand \U$30376 ( \30753 , \30735 , \30724 );
nand \U$30377 ( \30754 , \30752 , \30753 );
or \U$30378 ( \30755 , \30715 , \30754 );
not \U$30379 ( \30756 , \9792 );
and \U$30380 ( \30757 , RIae7a2b8_175, \9298 );
not \U$30381 ( \30758 , RIae7a2b8_175);
and \U$30382 ( \30759 , \30758 , \17242 );
nor \U$30383 ( \30760 , \30757 , \30759 );
not \U$30384 ( \30761 , \30760 );
or \U$30385 ( \30762 , \30756 , \30761 );
nand \U$30386 ( \30763 , \30494 , \16135 );
nand \U$30387 ( \30764 , \30762 , \30763 );
not \U$30388 ( \30765 , \9699 );
not \U$30389 ( \30766 , \30534 );
or \U$30390 ( \30767 , \30765 , \30766 );
and \U$30391 ( \30768 , \12700 , \11114 );
not \U$30392 ( \30769 , \12700 );
and \U$30393 ( \30770 , \30769 , RIae7a240_174);
nor \U$30394 ( \30771 , \30768 , \30770 );
nand \U$30395 ( \30772 , \30771 , \9687 );
nand \U$30396 ( \30773 , \30767 , \30772 );
xor \U$30397 ( \30774 , \30764 , \30773 );
not \U$30398 ( \30775 , \10638 );
xor \U$30399 ( \30776 , RIae7a510_180, \4982 );
not \U$30400 ( \30777 , \30776 );
or \U$30401 ( \30778 , \30775 , \30777 );
nand \U$30402 ( \30779 , \30384 , \10631 );
nand \U$30403 ( \30780 , \30778 , \30779 );
and \U$30404 ( \30781 , \30774 , \30780 );
and \U$30405 ( \30782 , \30764 , \30773 );
or \U$30406 ( \30783 , \30781 , \30782 );
nand \U$30407 ( \30784 , \30755 , \30783 );
nand \U$30408 ( \30785 , \30715 , \30754 );
nand \U$30409 ( \30786 , \30784 , \30785 );
not \U$30410 ( \30787 , \30786 );
or \U$30411 ( \30788 , \30648 , \30787 );
or \U$30412 ( \30789 , \30786 , \30647 );
nand \U$30413 ( \30790 , \30788 , \30789 );
not \U$30414 ( \30791 , \30790 );
xnor \U$30415 ( \30792 , \30315 , \30367 );
not \U$30416 ( \30793 , \30792 );
xnor \U$30417 ( \30794 , \30506 , \30497 );
not \U$30418 ( \30795 , \30794 );
nand \U$30419 ( \30796 , \30793 , \30795 );
not \U$30420 ( \30797 , \30794 );
not \U$30421 ( \30798 , \30792 );
or \U$30422 ( \30799 , \30797 , \30798 );
xor \U$30423 ( \30800 , \30521 , \30530 );
xor \U$30424 ( \30801 , \30800 , \30536 );
nand \U$30425 ( \30802 , \30799 , \30801 );
nand \U$30426 ( \30803 , \30796 , \30802 );
not \U$30427 ( \30804 , \30803 );
or \U$30428 ( \30805 , \30791 , \30804 );
not \U$30429 ( \30806 , \30785 );
not \U$30430 ( \30807 , \30784 );
or \U$30431 ( \30808 , \30806 , \30807 );
nand \U$30432 ( \30809 , \30808 , \30646 );
nand \U$30433 ( \30810 , \30805 , \30809 );
xor \U$30434 ( \30811 , \30598 , \30810 );
not \U$30435 ( \30812 , \30811 );
or \U$30436 ( \30813 , \30596 , \30812 );
nand \U$30437 ( \30814 , \30598 , \30810 );
nand \U$30438 ( \30815 , \30813 , \30814 );
xor \U$30439 ( \30816 , \30237 , \30223 );
xnor \U$30440 ( \30817 , \30816 , \30240 );
xor \U$30441 ( \30818 , \30815 , \30817 );
not \U$30442 ( \30819 , \9478 );
not \U$30443 ( \30820 , \30463 );
or \U$30444 ( \30821 , \30819 , \30820 );
and \U$30445 ( \30822 , RIae7a6f0_184, \3098 );
not \U$30446 ( \30823 , RIae7a6f0_184);
and \U$30447 ( \30824 , \30823 , \6171 );
or \U$30448 ( \30825 , \30822 , \30824 );
nand \U$30449 ( \30826 , \30825 , \9473 );
nand \U$30450 ( \30827 , \30821 , \30826 );
xor \U$30451 ( \30828 , \30340 , \30349 );
xor \U$30452 ( \30829 , \30828 , \30359 );
nor \U$30453 ( \30830 , \30827 , \30829 );
not \U$30454 ( \30831 , \10667 );
xor \U$30455 ( \30832 , RIae7a150_172, \1956 );
not \U$30456 ( \30833 , \30832 );
or \U$30457 ( \30834 , \30831 , \30833 );
nand \U$30458 ( \30835 , \30456 , \9777 );
nand \U$30459 ( \30836 , \30834 , \30835 );
not \U$30460 ( \30837 , \30836 );
or \U$30461 ( \30838 , \30830 , \30837 );
nand \U$30462 ( \30839 , \30827 , \30829 );
nand \U$30463 ( \30840 , \30838 , \30839 );
not \U$30464 ( \30841 , \30840 );
not \U$30465 ( \30842 , \11439 );
xnor \U$30466 ( \30843 , RIae7a7e0_186, \3524 );
not \U$30467 ( \30844 , \30843 );
or \U$30468 ( \30845 , \30842 , \30844 );
nand \U$30469 ( \30846 , \30420 , \10519 );
nand \U$30470 ( \30847 , \30845 , \30846 );
not \U$30471 ( \30848 , \30847 );
not \U$30472 ( \30849 , \5039 );
and \U$30473 ( \30850 , RIae79d90_164, \10937 );
not \U$30474 ( \30851 , RIae79d90_164);
and \U$30475 ( \30852 , \30851 , \12600 );
or \U$30476 ( \30853 , \30850 , \30852 );
not \U$30477 ( \30854 , \30853 );
or \U$30478 ( \30855 , \30849 , \30854 );
nand \U$30479 ( \30856 , \30320 , \5049 );
nand \U$30480 ( \30857 , \30855 , \30856 );
not \U$30481 ( \30858 , \30857 );
not \U$30482 ( \30859 , \30393 );
not \U$30483 ( \30860 , \4852 );
and \U$30484 ( \30861 , \30859 , \30860 );
not \U$30485 ( \30862 , \12484 );
not \U$30486 ( \30863 , \10892 );
and \U$30487 ( \30864 , \30862 , \30863 );
and \U$30488 ( \30865 , \14148 , \6270 );
nor \U$30489 ( \30866 , \30864 , \30865 );
nor \U$30490 ( \30867 , \30866 , \11760 );
nor \U$30491 ( \30868 , \30861 , \30867 );
not \U$30492 ( \30869 , \30868 );
and \U$30493 ( \30870 , \30858 , \30869 );
and \U$30494 ( \30871 , \30857 , \30868 );
nor \U$30495 ( \30872 , \30870 , \30871 );
not \U$30496 ( \30873 , \30872 );
not \U$30497 ( \30874 , \30873 );
or \U$30498 ( \30875 , \30848 , \30874 );
not \U$30499 ( \30876 , \30868 );
nand \U$30500 ( \30877 , \30876 , \30857 );
nand \U$30501 ( \30878 , \30875 , \30877 );
not \U$30502 ( \30879 , \30878 );
not \U$30503 ( \30880 , \30879 );
not \U$30504 ( \30881 , \10275 );
not \U$30505 ( \30882 , \30405 );
or \U$30506 ( \30883 , \30881 , \30882 );
not \U$30507 ( \30884 , \11207 );
not \U$30508 ( \30885 , \2309 );
or \U$30509 ( \30886 , \30884 , \30885 );
or \U$30510 ( \30887 , \2309 , \18088 );
nand \U$30511 ( \30888 , \30886 , \30887 );
nand \U$30512 ( \30889 , \30888 , \17847 );
nand \U$30513 ( \30890 , \30883 , \30889 );
not \U$30514 ( \30891 , \9728 );
and \U$30515 ( \30892 , RIae7a060_170, \4837 );
not \U$30516 ( \30893 , RIae7a060_170);
and \U$30517 ( \30894 , \30893 , \2564 );
nor \U$30518 ( \30895 , \30892 , \30894 );
not \U$30519 ( \30896 , \30895 );
or \U$30520 ( \30897 , \30891 , \30896 );
nand \U$30521 ( \30898 , \30430 , \11098 );
nand \U$30522 ( \30899 , \30897 , \30898 );
xor \U$30523 ( \30900 , \30890 , \30899 );
not \U$30524 ( \30901 , \16383 );
not \U$30525 ( \30902 , \14671 );
not \U$30526 ( \30903 , \14023 );
or \U$30527 ( \30904 , \30902 , \30903 );
or \U$30528 ( \30905 , \3070 , \14671 );
nand \U$30529 ( \30906 , \30904 , \30905 );
not \U$30530 ( \30907 , \30906 );
or \U$30531 ( \30908 , \30901 , \30907 );
nand \U$30532 ( \30909 , \30441 , RIae7aab0_192);
nand \U$30533 ( \30910 , \30908 , \30909 );
and \U$30534 ( \30911 , \30900 , \30910 );
and \U$30535 ( \30912 , \30890 , \30899 );
or \U$30536 ( \30913 , \30911 , \30912 );
not \U$30537 ( \30914 , \30913 );
or \U$30538 ( \30915 , \30880 , \30914 );
or \U$30539 ( \30916 , \30913 , \30879 );
nand \U$30540 ( \30917 , \30915 , \30916 );
not \U$30541 ( \30918 , \30917 );
or \U$30542 ( \30919 , \30841 , \30918 );
not \U$30543 ( \30920 , \30879 );
nand \U$30544 ( \30921 , \30920 , \30913 );
nand \U$30545 ( \30922 , \30919 , \30921 );
not \U$30546 ( \30923 , \30922 );
xor \U$30547 ( \30924 , \30541 , \30540 );
xnor \U$30548 ( \30925 , \30924 , \30509 );
xor \U$30549 ( \30926 , \30304 , \30273 );
xor \U$30550 ( \30927 , \30926 , \30372 );
and \U$30551 ( \30928 , \30925 , \30927 );
not \U$30552 ( \30929 , \30925 );
not \U$30553 ( \30930 , \30927 );
and \U$30554 ( \30931 , \30929 , \30930 );
nor \U$30555 ( \30932 , \30928 , \30931 );
not \U$30556 ( \30933 , \30932 );
or \U$30557 ( \30934 , \30923 , \30933 );
nand \U$30558 ( \30935 , \30925 , \30927 );
nand \U$30559 ( \30936 , \30934 , \30935 );
not \U$30560 ( \30937 , \30936 );
xor \U$30561 ( \30938 , \29292 , \29302 );
xor \U$30562 ( \30939 , \30938 , \29313 );
not \U$30563 ( \30940 , \30939 );
xor \U$30564 ( \30941 , \27728 , \27801 );
xnor \U$30565 ( \30942 , \30941 , \27806 );
not \U$30566 ( \30943 , \30942 );
not \U$30567 ( \30944 , \30943 );
or \U$30568 ( \30945 , \30940 , \30944 );
not \U$30569 ( \30946 , \30939 );
not \U$30570 ( \30947 , \30946 );
not \U$30571 ( \30948 , \30942 );
or \U$30572 ( \30949 , \30947 , \30948 );
and \U$30573 ( \30950 , \27823 , \27853 );
not \U$30574 ( \30951 , \27823 );
and \U$30575 ( \30952 , \30951 , \27839 );
or \U$30576 ( \30953 , \30950 , \30952 );
xnor \U$30577 ( \30954 , \30953 , \27850 );
nand \U$30578 ( \30955 , \30949 , \30954 );
nand \U$30579 ( \30956 , \30945 , \30955 );
xor \U$30580 ( \30957 , \27713 , \27809 );
xnor \U$30581 ( \30958 , \30957 , \27855 );
xor \U$30582 ( \30959 , \30956 , \30958 );
xor \U$30583 ( \30960 , \29280 , \29317 );
xor \U$30584 ( \30961 , \30960 , \29240 );
xnor \U$30585 ( \30962 , \30959 , \30961 );
not \U$30586 ( \30963 , \30962 );
not \U$30587 ( \30964 , \30963 );
or \U$30588 ( \30965 , \30937 , \30964 );
or \U$30589 ( \30966 , \30963 , \30936 );
xor \U$30590 ( \30967 , \30939 , \30943 );
xor \U$30591 ( \30968 , \30967 , \30954 );
xor \U$30592 ( \30969 , \30478 , \30446 );
xor \U$30593 ( \30970 , \30969 , \30411 );
xor \U$30594 ( \30971 , \30968 , \30970 );
not \U$30595 ( \30972 , \30468 );
nand \U$30596 ( \30973 , \30972 , \30477 );
xor \U$30597 ( \30974 , \30973 , \30475 );
not \U$30598 ( \30975 , \30974 );
not \U$30599 ( \30976 , \30407 );
not \U$30600 ( \30977 , \30397 );
xor \U$30601 ( \30978 , \30976 , \30977 );
not \U$30602 ( \30979 , \2007 );
not \U$30603 ( \30980 , \30627 );
or \U$30604 ( \30981 , \30979 , \30980 );
xor \U$30605 ( \30982 , \10007 , RIae797f0_152);
nand \U$30606 ( \30983 , \30982 , \1988 );
nand \U$30607 ( \30984 , \30981 , \30983 );
not \U$30608 ( \30985 , \30984 );
not \U$30609 ( \30986 , \2162 );
not \U$30610 ( \30987 , \30357 );
or \U$30611 ( \30988 , \30986 , \30987 );
not \U$30612 ( \30989 , \27786 );
not \U$30613 ( \30990 , \11321 );
or \U$30614 ( \30991 , \30989 , \30990 );
not \U$30615 ( \30992 , RIae79520_146);
or \U$30616 ( \30993 , \10272 , \30992 );
nand \U$30617 ( \30994 , \30991 , \30993 );
nand \U$30618 ( \30995 , \30994 , \2188 );
nand \U$30619 ( \30996 , \30988 , \30995 );
not \U$30620 ( \30997 , \30996 );
and \U$30621 ( \30998 , \12857 , \1820 );
not \U$30622 ( \30999 , \2249 );
not \U$30623 ( \31000 , \30673 );
or \U$30624 ( \31001 , \30999 , \31000 );
not \U$30625 ( \31002 , RIae79ac0_158);
not \U$30626 ( \31003 , \16006 );
or \U$30627 ( \31004 , \31002 , \31003 );
or \U$30628 ( \31005 , \16006 , RIae79ac0_158);
nand \U$30629 ( \31006 , \31004 , \31005 );
nand \U$30630 ( \31007 , \31006 , \2271 );
nand \U$30631 ( \31008 , \31001 , \31007 );
xor \U$30632 ( \31009 , \30998 , \31008 );
not \U$30633 ( \31010 , \2162 );
not \U$30634 ( \31011 , \30994 );
or \U$30635 ( \31012 , \31010 , \31011 );
not \U$30636 ( \31013 , RIae79520_146);
not \U$30637 ( \31014 , \10259 );
or \U$30638 ( \31015 , \31013 , \31014 );
or \U$30639 ( \31016 , \10259 , RIae79520_146);
nand \U$30640 ( \31017 , \31015 , \31016 );
nand \U$30641 ( \31018 , \31017 , \2188 );
nand \U$30642 ( \31019 , \31012 , \31018 );
and \U$30643 ( \31020 , \31009 , \31019 );
and \U$30644 ( \31021 , \30998 , \31008 );
nor \U$30645 ( \31022 , \31020 , \31021 );
not \U$30646 ( \31023 , \31022 );
or \U$30647 ( \31024 , \30997 , \31023 );
or \U$30648 ( \31025 , \31022 , \30996 );
nand \U$30649 ( \31026 , \31024 , \31025 );
not \U$30650 ( \31027 , \31026 );
or \U$30651 ( \31028 , \30985 , \31027 );
not \U$30652 ( \31029 , \31022 );
nand \U$30653 ( \31030 , \31029 , \30996 );
nand \U$30654 ( \31031 , \31028 , \31030 );
not \U$30655 ( \31032 , \2322 );
not \U$30656 ( \31033 , \30615 );
or \U$30657 ( \31034 , \31032 , \31033 );
xor \U$30658 ( \31035 , \10142 , RIae798e0_154);
nand \U$30659 ( \31036 , \31035 , \2339 );
nand \U$30660 ( \31037 , \31034 , \31036 );
not \U$30661 ( \31038 , \2450 );
and \U$30662 ( \31039 , RIae79778_151, \10066 );
not \U$30663 ( \31040 , RIae79778_151);
and \U$30664 ( \31041 , \31040 , \11230 );
nor \U$30665 ( \31042 , \31039 , \31041 );
not \U$30666 ( \31043 , \31042 );
or \U$30667 ( \31044 , \31038 , \31043 );
and \U$30668 ( \31045 , RIae79778_151, \14546 );
not \U$30669 ( \31046 , RIae79778_151);
and \U$30670 ( \31047 , \31046 , \9897 );
nor \U$30671 ( \31048 , \31045 , \31047 );
nand \U$30672 ( \31049 , \31048 , \2431 );
nand \U$30673 ( \31050 , \31044 , \31049 );
xor \U$30674 ( \31051 , \31037 , \31050 );
not \U$30675 ( \31052 , \2776 );
not \U$30676 ( \31053 , \30731 );
or \U$30677 ( \31054 , \31052 , \31053 );
and \U$30678 ( \31055 , \10208 , RIae79c28_161);
not \U$30679 ( \31056 , \10208 );
and \U$30680 ( \31057 , \31056 , \10584 );
nor \U$30681 ( \31058 , \31055 , \31057 );
nand \U$30682 ( \31059 , \31058 , \2417 );
nand \U$30683 ( \31060 , \31054 , \31059 );
and \U$30684 ( \31061 , \31051 , \31060 );
and \U$30685 ( \31062 , \31037 , \31050 );
or \U$30686 ( \31063 , \31061 , \31062 );
xor \U$30687 ( \31064 , \31031 , \31063 );
not \U$30688 ( \31065 , \10696 );
and \U$30689 ( \31066 , RIae7a498_179, \1859 );
not \U$30690 ( \31067 , RIae7a498_179);
and \U$30691 ( \31068 , \31067 , \12502 );
or \U$30692 ( \31069 , \31066 , \31068 );
not \U$30693 ( \31070 , \31069 );
or \U$30694 ( \31071 , \31065 , \31070 );
nand \U$30695 ( \31072 , \30473 , \11422 );
nand \U$30696 ( \31073 , \31071 , \31072 );
and \U$30697 ( \31074 , \31064 , \31073 );
and \U$30698 ( \31075 , \31031 , \31063 );
nor \U$30699 ( \31076 , \31074 , \31075 );
xnor \U$30700 ( \31077 , \30978 , \31076 );
not \U$30701 ( \31078 , \31077 );
or \U$30702 ( \31079 , \30975 , \31078 );
not \U$30703 ( \31080 , \31076 );
xor \U$30704 ( \31081 , \30977 , \30976 );
nand \U$30705 ( \31082 , \31080 , \31081 );
nand \U$30706 ( \31083 , \31079 , \31082 );
and \U$30707 ( \31084 , \30971 , \31083 );
and \U$30708 ( \31085 , \30968 , \30970 );
or \U$30709 ( \31086 , \31084 , \31085 );
nand \U$30710 ( \31087 , \30966 , \31086 );
nand \U$30711 ( \31088 , \30965 , \31087 );
and \U$30712 ( \31089 , \30818 , \31088 );
and \U$30713 ( \31090 , \30815 , \30817 );
or \U$30714 ( \31091 , \31089 , \31090 );
not \U$30715 ( \31092 , \31091 );
not \U$30716 ( \31093 , \31092 );
xnor \U$30717 ( \31094 , \30263 , \30248 );
not \U$30718 ( \31095 , \31094 );
or \U$30719 ( \31096 , \31093 , \31095 );
not \U$30720 ( \31097 , \29534 );
and \U$30721 ( \31098 , \29543 , \31097 );
not \U$30722 ( \31099 , \29543 );
and \U$30723 ( \31100 , \31099 , \29534 );
nor \U$30724 ( \31101 , \31098 , \31100 );
not \U$30725 ( \31102 , \30234 );
not \U$30726 ( \31103 , \30233 );
nand \U$30727 ( \31104 , \31103 , \30236 );
not \U$30728 ( \31105 , \31104 );
or \U$30729 ( \31106 , \31102 , \31105 );
or \U$30730 ( \31107 , \31104 , \30234 );
nand \U$30731 ( \31108 , \31106 , \31107 );
xor \U$30732 ( \31109 , \31101 , \31108 );
xor \U$30733 ( \31110 , \29440 , \29368 );
not \U$30734 ( \31111 , \31110 );
not \U$30735 ( \31112 , \29531 );
not \U$30736 ( \31113 , \29521 );
not \U$30737 ( \31114 , \31113 );
and \U$30738 ( \31115 , \31112 , \31114 );
and \U$30739 ( \31116 , \29531 , \31113 );
nor \U$30740 ( \31117 , \31115 , \31116 );
xor \U$30741 ( \31118 , \29509 , \31117 );
not \U$30742 ( \31119 , \31118 );
xor \U$30743 ( \31120 , \29213 , \29225 );
xor \U$30744 ( \31121 , \31120 , \29237 );
not \U$30745 ( \31122 , \31121 );
or \U$30746 ( \31123 , \31119 , \31122 );
or \U$30747 ( \31124 , \31121 , \31118 );
nand \U$30748 ( \31125 , \31123 , \31124 );
not \U$30749 ( \31126 , \31125 );
or \U$30750 ( \31127 , \31111 , \31126 );
not \U$30751 ( \31128 , \31118 );
nand \U$30752 ( \31129 , \31128 , \31121 );
nand \U$30753 ( \31130 , \31127 , \31129 );
not \U$30754 ( \31131 , \31130 );
and \U$30755 ( \31132 , \31109 , \31131 );
and \U$30756 ( \31133 , \31101 , \31108 );
or \U$30757 ( \31134 , \31132 , \31133 );
not \U$30758 ( \31135 , \31134 );
not \U$30759 ( \31136 , \31135 );
not \U$30760 ( \31137 , \30958 );
not \U$30761 ( \31138 , \30961 );
or \U$30762 ( \31139 , \31137 , \31138 );
nand \U$30763 ( \31140 , \31139 , \30956 );
or \U$30764 ( \31141 , \30958 , \30961 );
nand \U$30765 ( \31142 , \31140 , \31141 );
not \U$30766 ( \31143 , \31142 );
not \U$30767 ( \31144 , \31143 );
xor \U$30768 ( \31145 , \29320 , \29358 );
xor \U$30769 ( \31146 , \31145 , \29487 );
not \U$30770 ( \31147 , \31146 );
or \U$30771 ( \31148 , \31144 , \31147 );
or \U$30772 ( \31149 , \31146 , \31143 );
nand \U$30773 ( \31150 , \31148 , \31149 );
not \U$30774 ( \31151 , \31150 );
or \U$30775 ( \31152 , \31136 , \31151 );
nand \U$30776 ( \31153 , \31146 , \31142 );
nand \U$30777 ( \31154 , \31152 , \31153 );
buf \U$30778 ( \31155 , \31154 );
nand \U$30779 ( \31156 , \31096 , \31155 );
not \U$30780 ( \31157 , \31094 );
nand \U$30781 ( \31158 , \31157 , \31091 );
nand \U$30782 ( \31159 , \31156 , \31158 );
not \U$30783 ( \31160 , \29850 );
nand \U$30784 ( \31161 , \31160 , \29577 );
not \U$30785 ( \31162 , \31161 );
not \U$30786 ( \31163 , \29848 );
and \U$30787 ( \31164 , \31162 , \31163 );
and \U$30788 ( \31165 , \31161 , \29848 );
nor \U$30789 ( \31166 , \31164 , \31165 );
nand \U$30790 ( \31167 , \31159 , \31166 );
not \U$30791 ( \31168 , \31167 );
xor \U$30792 ( \31169 , \30217 , \30269 );
xnor \U$30793 ( \31170 , \31169 , \30578 );
not \U$30794 ( \31171 , \31170 );
or \U$30795 ( \31172 , \31168 , \31171 );
not \U$30796 ( \31173 , \31166 );
not \U$30797 ( \31174 , \31159 );
nand \U$30798 ( \31175 , \31173 , \31174 );
nand \U$30799 ( \31176 , \31172 , \31175 );
nand \U$30800 ( \31177 , \30593 , \31176 );
xor \U$30801 ( \31178 , \31166 , \31174 );
xnor \U$30802 ( \31179 , \31178 , \31170 );
not \U$30803 ( \31180 , \30574 );
xnor \U$30804 ( \31181 , \30569 , \30565 );
not \U$30805 ( \31182 , \31181 );
or \U$30806 ( \31183 , \31180 , \31182 );
or \U$30807 ( \31184 , \31181 , \30574 );
nand \U$30808 ( \31185 , \31183 , \31184 );
not \U$30809 ( \31186 , \31185 );
xor \U$30810 ( \31187 , \31154 , \31091 );
xnor \U$30811 ( \31188 , \31187 , \31094 );
not \U$30812 ( \31189 , \31188 );
nand \U$30813 ( \31190 , \31186 , \31189 );
not \U$30814 ( \31191 , \31185 );
not \U$30815 ( \31192 , \31188 );
or \U$30816 ( \31193 , \31191 , \31192 );
xor \U$30817 ( \31194 , \30558 , \30553 );
xnor \U$30818 ( \31195 , \31194 , \30561 );
not \U$30819 ( \31196 , \31195 );
xor \U$30820 ( \31197 , \31142 , \31134 );
xnor \U$30821 ( \31198 , \31197 , \31146 );
buf \U$30822 ( \31199 , \31198 );
nand \U$30823 ( \31200 , \31196 , \31199 );
xor \U$30824 ( \31201 , \30815 , \30817 );
xor \U$30825 ( \31202 , \31201 , \31088 );
not \U$30826 ( \31203 , \31198 );
nand \U$30827 ( \31204 , \31203 , \31195 );
nand \U$30828 ( \31205 , \31202 , \31204 );
and \U$30829 ( \31206 , \31200 , \31205 );
nand \U$30830 ( \31207 , \31193 , \31206 );
nand \U$30831 ( \31208 , \31190 , \31207 );
nor \U$30832 ( \31209 , \31179 , \31208 );
nand \U$30833 ( \31210 , \31177 , \31209 );
not \U$30834 ( \31211 , \31210 );
not \U$30835 ( \31212 , \31176 );
not \U$30836 ( \31213 , \30593 );
nand \U$30837 ( \31214 , \31212 , \31213 );
not \U$30838 ( \31215 , \29856 );
not \U$30839 ( \31216 , \31215 );
not \U$30840 ( \31217 , \30589 );
or \U$30841 ( \31218 , \31216 , \31217 );
nand \U$30842 ( \31219 , \30579 , \30208 , \30581 );
nand \U$30843 ( \31220 , \31218 , \31219 );
not \U$30844 ( \31221 , \31220 );
not \U$30845 ( \31222 , \30071 );
not \U$30846 ( \31223 , \30090 );
or \U$30847 ( \31224 , \31222 , \31223 );
nand \U$30848 ( \31225 , \30078 , \30089 );
nand \U$30849 ( \31226 , \31224 , \31225 );
not \U$30850 ( \31227 , \31226 );
not \U$30851 ( \31228 , \29168 );
not \U$30852 ( \31229 , \29177 );
or \U$30853 ( \31230 , \31228 , \31229 );
nand \U$30854 ( \31231 , \31230 , \29190 );
or \U$30855 ( \31232 , \29177 , \29168 );
nand \U$30856 ( \31233 , \31231 , \31232 );
xnor \U$30857 ( \31234 , \31227 , \31233 );
not \U$30858 ( \31235 , \29054 );
not \U$30859 ( \31236 , \29067 );
or \U$30860 ( \31237 , \31235 , \31236 );
nand \U$30861 ( \31238 , \31237 , \29038 );
not \U$30862 ( \31239 , \29067 );
nand \U$30863 ( \31240 , \31239 , \29055 );
nand \U$30864 ( \31241 , \31238 , \31240 );
xor \U$30865 ( \31242 , \31234 , \31241 );
not \U$30866 ( \31243 , \30149 );
xnor \U$30867 ( \31244 , \30143 , \30154 );
not \U$30868 ( \31245 , \31244 );
or \U$30869 ( \31246 , \31243 , \31245 );
nand \U$30870 ( \31247 , \30155 , \30144 );
nand \U$30871 ( \31248 , \31246 , \31247 );
not \U$30872 ( \31249 , \31248 );
xor \U$30873 ( \31250 , \31242 , \31249 );
not \U$30874 ( \31251 , \29075 );
not \U$30875 ( \31252 , \29196 );
not \U$30876 ( \31253 , \31252 );
or \U$30877 ( \31254 , \31251 , \31253 );
not \U$30878 ( \31255 , \29153 );
nand \U$30879 ( \31256 , \31255 , \29192 );
nand \U$30880 ( \31257 , \31254 , \31256 );
xnor \U$30881 ( \31258 , \31250 , \31257 );
not \U$30882 ( \31259 , \29020 );
not \U$30883 ( \31260 , \29201 );
or \U$30884 ( \31261 , \31259 , \31260 );
nand \U$30885 ( \31262 , \29200 , \29030 );
nand \U$30886 ( \31263 , \31261 , \31262 );
not \U$30887 ( \31264 , \31263 );
xor \U$30888 ( \31265 , \31258 , \31264 );
not \U$30889 ( \31266 , \30187 );
not \U$30890 ( \31267 , \30169 );
not \U$30891 ( \31268 , \30199 );
or \U$30892 ( \31269 , \31267 , \31268 );
or \U$30893 ( \31270 , \30199 , \30169 );
nand \U$30894 ( \31271 , \31269 , \31270 );
not \U$30895 ( \31272 , \31271 );
or \U$30896 ( \31273 , \31266 , \31272 );
not \U$30897 ( \31274 , \30169 );
nand \U$30898 ( \31275 , \31274 , \30199 );
nand \U$30899 ( \31276 , \31273 , \31275 );
xor \U$30900 ( \31277 , \31265 , \31276 );
not \U$30901 ( \31278 , \29863 );
not \U$30902 ( \31279 , \30045 );
or \U$30903 ( \31280 , \31278 , \31279 );
not \U$30904 ( \31281 , \29863 );
not \U$30905 ( \31282 , \31281 );
not \U$30906 ( \31283 , \30044 );
or \U$30907 ( \31284 , \31282 , \31283 );
nand \U$30908 ( \31285 , \31284 , \30207 );
nand \U$30909 ( \31286 , \31280 , \31285 );
xor \U$30910 ( \31287 , \31277 , \31286 );
not \U$30911 ( \31288 , \29992 );
not \U$30912 ( \31289 , \29958 );
not \U$30913 ( \31290 , \30026 );
or \U$30914 ( \31291 , \31289 , \31290 );
or \U$30915 ( \31292 , \30026 , \29958 );
nand \U$30916 ( \31293 , \31291 , \31292 );
not \U$30917 ( \31294 , \31293 );
or \U$30918 ( \31295 , \31288 , \31294 );
not \U$30919 ( \31296 , \29958 );
nand \U$30920 ( \31297 , \31296 , \30026 );
nand \U$30921 ( \31298 , \31295 , \31297 );
not \U$30922 ( \31299 , \31298 );
not \U$30923 ( \31300 , \29148 );
not \U$30924 ( \31301 , \29136 );
or \U$30925 ( \31302 , \31300 , \31301 );
nand \U$30926 ( \31303 , \29082 , \29135 );
nand \U$30927 ( \31304 , \31302 , \31303 );
not \U$30928 ( \31305 , \2450 );
and \U$30929 ( \31306 , RIae79778_151, \13287 );
not \U$30930 ( \31307 , RIae79778_151);
and \U$30931 ( \31308 , \31307 , \14691 );
or \U$30932 ( \31309 , \31306 , \31308 );
not \U$30933 ( \31310 , \31309 );
or \U$30934 ( \31311 , \31305 , \31310 );
nand \U$30935 ( \31312 , \29173 , \2432 );
nand \U$30936 ( \31313 , \31311 , \31312 );
not \U$30937 ( \31314 , \1501 );
not \U$30938 ( \31315 , \1503 );
not \U$30939 ( \31316 , \11317 );
or \U$30940 ( \31317 , \31315 , \31316 );
or \U$30941 ( \31318 , \11317 , \8789 );
nand \U$30942 ( \31319 , \31317 , \31318 );
not \U$30943 ( \31320 , \31319 );
or \U$30944 ( \31321 , \31314 , \31320 );
nand \U$30945 ( \31322 , \29108 , \1497 );
nand \U$30946 ( \31323 , \31321 , \31322 );
not \U$30947 ( \31324 , \31323 );
not \U$30948 ( \31325 , \31324 );
not \U$30949 ( \31326 , \1012 );
not \U$30950 ( \31327 , RIae79160_138);
not \U$30951 ( \31328 , \10844 );
or \U$30952 ( \31329 , \31327 , \31328 );
or \U$30953 ( \31330 , \10844 , RIae79160_138);
nand \U$30954 ( \31331 , \31329 , \31330 );
not \U$30955 ( \31332 , \31331 );
or \U$30956 ( \31333 , \31326 , \31332 );
nand \U$30957 ( \31334 , \29094 , \1007 );
nand \U$30958 ( \31335 , \31333 , \31334 );
not \U$30959 ( \31336 , \31335 );
nand \U$30960 ( \31337 , \12857 , \1048 );
not \U$30961 ( \31338 , \31337 );
and \U$30962 ( \31339 , \31336 , \31338 );
and \U$30963 ( \31340 , \31335 , \31337 );
nor \U$30964 ( \31341 , \31339 , \31340 );
not \U$30965 ( \31342 , \31341 );
not \U$30966 ( \31343 , \31342 );
or \U$30967 ( \31344 , \31325 , \31343 );
nand \U$30968 ( \31345 , \31341 , \31323 );
nand \U$30969 ( \31346 , \31344 , \31345 );
not \U$30970 ( \31347 , \31346 );
and \U$30971 ( \31348 , \2183 , \10083 );
not \U$30972 ( \31349 , \2183 );
and \U$30973 ( \31350 , \31349 , \10207 );
nor \U$30974 ( \31351 , \31348 , \31350 );
nand \U$30975 ( \31352 , \31351 , \2162 );
not \U$30976 ( \31353 , \31352 );
not \U$30977 ( \31354 , \2188 );
nor \U$30978 ( \31355 , \31354 , \30066 );
nor \U$30979 ( \31356 , \31353 , \31355 );
not \U$30980 ( \31357 , \31356 );
or \U$30981 ( \31358 , \31347 , \31357 );
not \U$30982 ( \31359 , \31352 );
not \U$30983 ( \31360 , \31355 );
not \U$30984 ( \31361 , \31360 );
or \U$30985 ( \31362 , \31359 , \31361 );
not \U$30986 ( \31363 , \31346 );
nand \U$30987 ( \31364 , \31362 , \31363 );
nand \U$30988 ( \31365 , \31358 , \31364 );
not \U$30989 ( \31366 , \2272 );
not \U$30990 ( \31367 , \30126 );
or \U$30991 ( \31368 , \31366 , \31367 );
and \U$30992 ( \31369 , RIae79ac0_158, \9897 );
not \U$30993 ( \31370 , RIae79ac0_158);
and \U$30994 ( \31371 , \31370 , \17185 );
or \U$30995 ( \31372 , \31369 , \31371 );
nand \U$30996 ( \31373 , \31372 , \2249 );
nand \U$30997 ( \31374 , \31368 , \31373 );
xnor \U$30998 ( \31375 , \31365 , \31374 );
xor \U$30999 ( \31376 , \31313 , \31375 );
not \U$31000 ( \31377 , \1843 );
not \U$31001 ( \31378 , \30116 );
or \U$31002 ( \31379 , \31377 , \31378 );
not \U$31003 ( \31380 , RIae79688_149);
not \U$31004 ( \31381 , \10000 );
or \U$31005 ( \31382 , \31380 , \31381 );
or \U$31006 ( \31383 , \16719 , RIae79688_149);
nand \U$31007 ( \31384 , \31382 , \31383 );
nand \U$31008 ( \31385 , \31384 , \1820 );
nand \U$31009 ( \31386 , \31379 , \31385 );
not \U$31010 ( \31387 , \2457 );
not \U$31011 ( \31388 , \30137 );
or \U$31012 ( \31389 , \31387 , \31388 );
and \U$31013 ( \31390 , \3810 , \10464 );
not \U$31014 ( \31391 , \3810 );
and \U$31015 ( \31392 , \31391 , \16837 );
nor \U$31016 ( \31393 , \31390 , \31392 );
nand \U$31017 ( \31394 , \31393 , \1919 );
nand \U$31018 ( \31395 , \31389 , \31394 );
and \U$31019 ( \31396 , \31386 , \31395 );
not \U$31020 ( \31397 , \31386 );
not \U$31021 ( \31398 , \31395 );
and \U$31022 ( \31399 , \31397 , \31398 );
nor \U$31023 ( \31400 , \31396 , \31399 );
buf \U$31024 ( \31401 , \31400 );
xnor \U$31025 ( \31402 , \31376 , \31401 );
xnor \U$31026 ( \31403 , \31304 , \31402 );
not \U$31027 ( \31404 , \31403 );
not \U$31028 ( \31405 , \30175 );
not \U$31029 ( \31406 , \31405 );
not \U$31030 ( \31407 , \31406 );
not \U$31031 ( \31408 , \30186 );
or \U$31032 ( \31409 , \31407 , \31408 );
not \U$31033 ( \31410 , \30186 );
not \U$31034 ( \31411 , \31410 );
not \U$31035 ( \31412 , \31405 );
or \U$31036 ( \31413 , \31411 , \31412 );
not \U$31037 ( \31414 , \30181 );
nand \U$31038 ( \31415 , \31413 , \31414 );
nand \U$31039 ( \31416 , \31409 , \31415 );
not \U$31040 ( \31417 , \31416 );
or \U$31041 ( \31418 , \31404 , \31417 );
or \U$31042 ( \31419 , \31416 , \31403 );
nand \U$31043 ( \31420 , \31418 , \31419 );
not \U$31044 ( \31421 , \31420 );
not \U$31045 ( \31422 , \31421 );
and \U$31046 ( \31423 , \31299 , \31422 );
and \U$31047 ( \31424 , \31298 , \31421 );
nor \U$31048 ( \31425 , \31423 , \31424 );
not \U$31049 ( \31426 , \29948 );
not \U$31050 ( \31427 , \29911 );
or \U$31051 ( \31428 , \31426 , \31427 );
nand \U$31052 ( \31429 , \29906 , \29897 );
nand \U$31053 ( \31430 , \31428 , \31429 );
not \U$31054 ( \31431 , \29873 );
not \U$31055 ( \31432 , \29896 );
or \U$31056 ( \31433 , \31431 , \31432 );
nand \U$31057 ( \31434 , \29891 , \29880 );
nand \U$31058 ( \31435 , \31433 , \31434 );
not \U$31059 ( \31436 , \30003 );
not \U$31060 ( \31437 , \30025 );
or \U$31061 ( \31438 , \31436 , \31437 );
nand \U$31062 ( \31439 , \31438 , \30014 );
not \U$31063 ( \31440 , \30025 );
not \U$31064 ( \31441 , \30003 );
nand \U$31065 ( \31442 , \31440 , \31441 );
nand \U$31066 ( \31443 , \31439 , \31442 );
not \U$31067 ( \31444 , \31443 );
xor \U$31068 ( \31445 , \31435 , \31444 );
not \U$31069 ( \31446 , \29932 );
not \U$31070 ( \31447 , \29944 );
or \U$31071 ( \31448 , \31446 , \31447 );
not \U$31072 ( \31449 , \29930 );
nand \U$31073 ( \31450 , \31448 , \31449 );
xnor \U$31074 ( \31451 , \31445 , \31450 );
xor \U$31075 ( \31452 , \31430 , \31451 );
not \U$31076 ( \31453 , \10275 );
not \U$31077 ( \31454 , RIae7a8d0_188);
not \U$31078 ( \31455 , \1405 );
or \U$31079 ( \31456 , \31454 , \31455 );
or \U$31080 ( \31457 , \2101 , RIae7a8d0_188);
nand \U$31081 ( \31458 , \31456 , \31457 );
not \U$31082 ( \31459 , \31458 );
or \U$31083 ( \31460 , \31453 , \31459 );
nand \U$31084 ( \31461 , \29889 , \14510 );
nand \U$31085 ( \31462 , \31460 , \31461 );
not \U$31086 ( \31463 , \31462 );
not \U$31087 ( \31464 , \4842 );
not \U$31088 ( \31465 , \29144 );
or \U$31089 ( \31466 , \31464 , \31465 );
not \U$31090 ( \31467 , RIae79ca0_162);
not \U$31091 ( \31468 , \10409 );
or \U$31092 ( \31469 , \31467 , \31468 );
not \U$31093 ( \31470 , \9290 );
or \U$31094 ( \31471 , \31470 , RIae79ca0_162);
nand \U$31095 ( \31472 , \31469 , \31471 );
nand \U$31096 ( \31473 , \31472 , \4853 );
nand \U$31097 ( \31474 , \31466 , \31473 );
not \U$31098 ( \31475 , \31474 );
not \U$31099 ( \31476 , \29121 );
not \U$31100 ( \31477 , \29130 );
or \U$31101 ( \31478 , \31476 , \31477 );
not \U$31102 ( \31479 , \29105 );
nand \U$31103 ( \31480 , \31479 , \29117 );
nand \U$31104 ( \31481 , \31478 , \31480 );
not \U$31105 ( \31482 , \31481 );
not \U$31106 ( \31483 , \31482 );
and \U$31107 ( \31484 , \31475 , \31483 );
and \U$31108 ( \31485 , \31474 , \31482 );
nor \U$31109 ( \31486 , \31484 , \31485 );
not \U$31110 ( \31487 , \31486 );
or \U$31111 ( \31488 , \31463 , \31487 );
or \U$31112 ( \31489 , \31462 , \31486 );
nand \U$31113 ( \31490 , \31488 , \31489 );
not \U$31114 ( \31491 , \29967 );
nand \U$31115 ( \31492 , \31491 , \29976 );
not \U$31116 ( \31493 , \31492 );
not \U$31117 ( \31494 , \29991 );
or \U$31118 ( \31495 , \31493 , \31494 );
or \U$31119 ( \31496 , \31491 , \29976 );
nand \U$31120 ( \31497 , \31495 , \31496 );
xor \U$31121 ( \31498 , \31490 , \31497 );
not \U$31122 ( \31499 , \5049 );
not \U$31123 ( \31500 , RIae79d90_164);
not \U$31124 ( \31501 , \16310 );
or \U$31125 ( \31502 , \31500 , \31501 );
or \U$31126 ( \31503 , \27827 , RIae79d90_164);
nand \U$31127 ( \31504 , \31502 , \31503 );
not \U$31128 ( \31505 , \31504 );
or \U$31129 ( \31506 , \31499 , \31505 );
nand \U$31130 ( \31507 , \29078 , \6091 );
nand \U$31131 ( \31508 , \31506 , \31507 );
not \U$31132 ( \31509 , \31508 );
not \U$31133 ( \31510 , \19362 );
not \U$31134 ( \31511 , \29035 );
or \U$31135 ( \31512 , \31510 , \31511 );
not \U$31136 ( \31513 , RIae79ef8_167);
not \U$31137 ( \31514 , \4928 );
or \U$31138 ( \31515 , \31513 , \31514 );
nand \U$31139 ( \31516 , \4168 , \6203 );
nand \U$31140 ( \31517 , \31515 , \31516 );
nand \U$31141 ( \31518 , \31517 , \10573 );
nand \U$31142 ( \31519 , \31512 , \31518 );
not \U$31143 ( \31520 , \31519 );
xor \U$31144 ( \31521 , \31509 , \31520 );
not \U$31145 ( \31522 , \11914 );
not \U$31146 ( \31523 , \29065 );
or \U$31147 ( \31524 , \31522 , \31523 );
and \U$31148 ( \31525 , \10492 , \11069 );
not \U$31149 ( \31526 , \10492 );
and \U$31150 ( \31527 , \31526 , RIae79fe8_169);
nor \U$31151 ( \31528 , \31525 , \31527 );
nand \U$31152 ( \31529 , \31528 , \9517 );
nand \U$31153 ( \31530 , \31524 , \31529 );
xnor \U$31154 ( \31531 , \31521 , \31530 );
xor \U$31155 ( \31532 , \31498 , \31531 );
xnor \U$31156 ( \31533 , \31452 , \31532 );
xor \U$31157 ( \31534 , \31425 , \31533 );
not \U$31158 ( \31535 , \30042 );
not \U$31159 ( \31536 , \30032 );
or \U$31160 ( \31537 , \31535 , \31536 );
not \U$31161 ( \31538 , \30028 );
nand \U$31162 ( \31539 , \31538 , \29950 );
nand \U$31163 ( \31540 , \31537 , \31539 );
not \U$31164 ( \31541 , \31540 );
xnor \U$31165 ( \31542 , \31534 , \31541 );
xnor \U$31166 ( \31543 , \31287 , \31542 );
not \U$31167 ( \31544 , \31543 );
not \U$31168 ( \31545 , \28684 );
not \U$31169 ( \31546 , \29206 );
or \U$31170 ( \31547 , \31545 , \31546 );
nand \U$31171 ( \31548 , \31547 , \29851 );
not \U$31172 ( \31549 , \29206 );
nand \U$31173 ( \31550 , \31549 , \29209 );
nand \U$31174 ( \31551 , \31548 , \31550 );
not \U$31175 ( \31552 , \31551 );
not \U$31176 ( \31553 , \2322 );
and \U$31177 ( \31554 , RIae798e0_154, \9412 );
not \U$31178 ( \31555 , RIae798e0_154);
and \U$31179 ( \31556 , \31555 , \11803 );
or \U$31180 ( \31557 , \31554 , \31556 );
not \U$31181 ( \31558 , \31557 );
or \U$31182 ( \31559 , \31553 , \31558 );
nand \U$31183 ( \31560 , \29159 , \14580 );
nand \U$31184 ( \31561 , \31559 , \31560 );
nand \U$31185 ( \31562 , \29185 , \1988 );
and \U$31186 ( \31563 , RIae797f0_152, \9456 );
not \U$31187 ( \31564 , RIae797f0_152);
and \U$31188 ( \31565 , \31564 , \9455 );
or \U$31189 ( \31566 , \31563 , \31565 );
nand \U$31190 ( \31567 , \31566 , \2007 );
nand \U$31191 ( \31568 , \31562 , \31567 );
xor \U$31192 ( \31569 , \31561 , \31568 );
not \U$31193 ( \31570 , \2767 );
not \U$31194 ( \31571 , \29044 );
or \U$31195 ( \31572 , \31570 , \31571 );
and \U$31196 ( \31573 , RIae79c28_161, \9316 );
not \U$31197 ( \31574 , RIae79c28_161);
and \U$31198 ( \31575 , \31574 , \16274 );
or \U$31199 ( \31576 , \31573 , \31575 );
nand \U$31200 ( \31577 , \31576 , \2776 );
nand \U$31201 ( \31578 , \31572 , \31577 );
xnor \U$31202 ( \31579 , \31569 , \31578 );
not \U$31203 ( \31580 , \30120 );
not \U$31204 ( \31581 , \30130 );
or \U$31205 ( \31582 , \31580 , \31581 );
or \U$31206 ( \31583 , \30130 , \30120 );
nand \U$31207 ( \31584 , \31583 , \30141 );
nand \U$31208 ( \31585 , \31582 , \31584 );
not \U$31209 ( \31586 , \9478 );
and \U$31210 ( \31587 , RIae7a6f0_184, \9696 );
not \U$31211 ( \31588 , RIae7a6f0_184);
and \U$31212 ( \31589 , \31588 , \17068 );
or \U$31213 ( \31590 , \31587 , \31589 );
not \U$31214 ( \31591 , \31590 );
or \U$31215 ( \31592 , \31586 , \31591 );
nand \U$31216 ( \31593 , \29971 , \9473 );
nand \U$31217 ( \31594 , \31592 , \31593 );
not \U$31218 ( \31595 , \31594 );
xor \U$31219 ( \31596 , \31585 , \31595 );
not \U$31220 ( \31597 , \11434 );
not \U$31221 ( \31598 , \29963 );
or \U$31222 ( \31599 , \31597 , \31598 );
not \U$31223 ( \31600 , \10625 );
not \U$31224 ( \31601 , \3748 );
or \U$31225 ( \31602 , \31600 , \31601 );
nand \U$31226 ( \31603 , \2835 , RIae7a498_179);
nand \U$31227 ( \31604 , \31602 , \31603 );
nand \U$31228 ( \31605 , \31604 , \10677 );
nand \U$31229 ( \31606 , \31599 , \31605 );
xnor \U$31230 ( \31607 , \31596 , \31606 );
xor \U$31231 ( \31608 , \31579 , \31607 );
not \U$31232 ( \31609 , \10638 );
not \U$31233 ( \31610 , \29869 );
or \U$31234 ( \31611 , \31609 , \31610 );
and \U$31235 ( \31612 , RIae7a510_180, \10905 );
not \U$31236 ( \31613 , RIae7a510_180);
and \U$31237 ( \31614 , \31613 , \10605 );
or \U$31238 ( \31615 , \31612 , \31614 );
nand \U$31239 ( \31616 , \31615 , \16358 );
nand \U$31240 ( \31617 , \31611 , \31616 );
not \U$31241 ( \31618 , \9622 );
and \U$31242 ( \31619 , \2576 , RIae7a3a8_177);
not \U$31243 ( \31620 , \2576 );
and \U$31244 ( \31621 , \31620 , \11690 );
nor \U$31245 ( \31622 , \31619 , \31621 );
not \U$31246 ( \31623 , \31622 );
or \U$31247 ( \31624 , \31618 , \31623 );
nand \U$31248 ( \31625 , \29916 , \9644 );
nand \U$31249 ( \31626 , \31624 , \31625 );
xor \U$31250 ( \31627 , \31617 , \31626 );
not \U$31251 ( \31628 , \11851 );
not \U$31252 ( \31629 , \29939 );
or \U$31253 ( \31630 , \31628 , \31629 );
not \U$31254 ( \31631 , \9537 );
not \U$31255 ( \31632 , \9807 );
or \U$31256 ( \31633 , \31631 , \31632 );
or \U$31257 ( \31634 , \9807 , \9537 );
nand \U$31258 ( \31635 , \31633 , \31634 );
nand \U$31259 ( \31636 , \31635 , \9527 );
nand \U$31260 ( \31637 , \31630 , \31636 );
xor \U$31261 ( \31638 , \31627 , \31637 );
xnor \U$31262 ( \31639 , \31608 , \31638 );
not \U$31263 ( \31640 , \30102 );
not \U$31264 ( \31641 , \30095 );
or \U$31265 ( \31642 , \31640 , \31641 );
nand \U$31266 ( \31643 , \30064 , \30094 );
nand \U$31267 ( \31644 , \31642 , \31643 );
not \U$31268 ( \31645 , \9792 );
not \U$31269 ( \31646 , \29999 );
or \U$31270 ( \31647 , \31645 , \31646 );
not \U$31271 ( \31648 , RIae7a2b8_175);
not \U$31272 ( \31649 , \3216 );
or \U$31273 ( \31650 , \31648 , \31649 );
or \U$31274 ( \31651 , \3216 , RIae7a2b8_175);
nand \U$31275 ( \31652 , \31650 , \31651 );
nand \U$31276 ( \31653 , \31652 , \9814 );
nand \U$31277 ( \31654 , \31647 , \31653 );
not \U$31278 ( \31655 , \13720 );
not \U$31279 ( \31656 , \29925 );
or \U$31280 ( \31657 , \31655 , \31656 );
and \U$31281 ( \31658 , RIae7a240_174, \14439 );
not \U$31282 ( \31659 , RIae7a240_174);
and \U$31283 ( \31660 , \31659 , \22917 );
or \U$31284 ( \31661 , \31658 , \31660 );
nand \U$31285 ( \31662 , \31661 , \13121 );
nand \U$31286 ( \31663 , \31657 , \31662 );
xor \U$31287 ( \31664 , \31654 , \31663 );
not \U$31288 ( \31665 , \9745 );
not \U$31289 ( \31666 , \11102 );
not \U$31290 ( \31667 , \11885 );
or \U$31291 ( \31668 , \31666 , \31667 );
or \U$31292 ( \31669 , \19857 , \11102 );
nand \U$31293 ( \31670 , \31668 , \31669 );
not \U$31294 ( \31671 , \31670 );
or \U$31295 ( \31672 , \31665 , \31671 );
nand \U$31296 ( \31673 , \30021 , \9730 );
nand \U$31297 ( \31674 , \31672 , \31673 );
xor \U$31298 ( \31675 , \31664 , \31674 );
xor \U$31299 ( \31676 , \31644 , \31675 );
not \U$31300 ( \31677 , \29096 );
nor \U$31301 ( \31678 , \31677 , \29101 );
not \U$31302 ( \31679 , \1863 );
not \U$31303 ( \31680 , \1884 );
not \U$31304 ( \31681 , \10042 );
or \U$31305 ( \31682 , \31680 , \31681 );
or \U$31306 ( \31683 , \10042 , \1884 );
nand \U$31307 ( \31684 , \31682 , \31683 );
not \U$31308 ( \31685 , \31684 );
or \U$31309 ( \31686 , \31679 , \31685 );
nand \U$31310 ( \31687 , \30085 , \1910 );
nand \U$31311 ( \31688 , \31686 , \31687 );
xor \U$31312 ( \31689 , \31678 , \31688 );
not \U$31313 ( \31690 , \2063 );
not \U$31314 ( \31691 , \29126 );
or \U$31315 ( \31692 , \31690 , \31691 );
and \U$31316 ( \31693 , \10149 , \2056 );
not \U$31317 ( \31694 , \10149 );
and \U$31318 ( \31695 , \31694 , RIae79610_148);
nor \U$31319 ( \31696 , \31693 , \31695 );
nand \U$31320 ( \31697 , \31696 , \2011 );
nand \U$31321 ( \31698 , \31692 , \31697 );
not \U$31322 ( \31699 , \31698 );
xor \U$31323 ( \31700 , \31689 , \31699 );
not \U$31324 ( \31701 , \9776 );
not \U$31325 ( \31702 , RIae7a150_172);
not \U$31326 ( \31703 , \2954 );
or \U$31327 ( \31704 , \31702 , \31703 );
or \U$31328 ( \31705 , \2155 , RIae7a150_172);
nand \U$31329 ( \31706 , \31704 , \31705 );
not \U$31330 ( \31707 , \31706 );
or \U$31331 ( \31708 , \31701 , \31707 );
nand \U$31332 ( \31709 , \30009 , \10667 );
nand \U$31333 ( \31710 , \31708 , \31709 );
not \U$31334 ( \31711 , \31710 );
xor \U$31335 ( \31712 , \31700 , \31711 );
not \U$31336 ( \31713 , \16383 );
not \U$31337 ( \31714 , \29986 );
or \U$31338 ( \31715 , \31713 , \31714 );
xor \U$31339 ( \31716 , \1124 , RIae7aa38_191);
nand \U$31340 ( \31717 , \31716 , RIae7aab0_192);
nand \U$31341 ( \31718 , \31715 , \31717 );
xor \U$31342 ( \31719 , \31712 , \31718 );
xnor \U$31343 ( \31720 , \31676 , \31719 );
not \U$31344 ( \31721 , \31720 );
xor \U$31345 ( \31722 , \31639 , \31721 );
or \U$31346 ( \31723 , \30111 , \30156 );
not \U$31347 ( \31724 , \30107 );
nand \U$31348 ( \31725 , \31724 , \30058 );
nand \U$31349 ( \31726 , \31723 , \31725 );
not \U$31350 ( \31727 , \31726 );
xnor \U$31351 ( \31728 , \31722 , \31727 );
not \U$31352 ( \31729 , \30051 );
not \U$31353 ( \31730 , \30201 );
or \U$31354 ( \31731 , \31729 , \31730 );
nand \U$31355 ( \31732 , \31731 , \30161 );
nand \U$31356 ( \31733 , \30202 , \30050 );
and \U$31357 ( \31734 , \31732 , \31733 );
xor \U$31358 ( \31735 , \31728 , \31734 );
not \U$31359 ( \31736 , \29011 );
not \U$31360 ( \31737 , \28694 );
not \U$31361 ( \31738 , \31737 );
not \U$31362 ( \31739 , \29205 );
or \U$31363 ( \31740 , \31738 , \31739 );
or \U$31364 ( \31741 , \29205 , \31737 );
nand \U$31365 ( \31742 , \31740 , \31741 );
not \U$31366 ( \31743 , \31742 );
or \U$31367 ( \31744 , \31736 , \31743 );
nand \U$31368 ( \31745 , \29205 , \28694 );
nand \U$31369 ( \31746 , \31744 , \31745 );
xor \U$31370 ( \31747 , \31735 , \31746 );
not \U$31371 ( \31748 , \31747 );
or \U$31372 ( \31749 , \31552 , \31748 );
or \U$31373 ( \31750 , \31551 , \31747 );
nand \U$31374 ( \31751 , \31749 , \31750 );
not \U$31375 ( \31752 , \31751 );
not \U$31376 ( \31753 , \31752 );
or \U$31377 ( \31754 , \31544 , \31753 );
not \U$31378 ( \31755 , \31543 );
nand \U$31379 ( \31756 , \31751 , \31755 );
nand \U$31380 ( \31757 , \31754 , \31756 );
not \U$31381 ( \31758 , \31757 );
nand \U$31382 ( \31759 , \31221 , \31758 );
not \U$31383 ( \31760 , \31277 );
not \U$31384 ( \31761 , \31542 );
or \U$31385 ( \31762 , \31760 , \31761 );
nand \U$31386 ( \31763 , \31762 , \31286 );
or \U$31387 ( \31764 , \31542 , \31277 );
not \U$31388 ( \31765 , RIae7aab0_192);
and \U$31389 ( \31766 , RIae7aa38_191, \12801 );
not \U$31390 ( \31767 , RIae7aa38_191);
and \U$31391 ( \31768 , \31767 , \12800 );
nor \U$31392 ( \31769 , \31766 , \31768 );
not \U$31393 ( \31770 , \31769 );
or \U$31394 ( \31771 , \31765 , \31770 );
nand \U$31395 ( \31772 , \31716 , \14667 );
nand \U$31396 ( \31773 , \31771 , \31772 );
not \U$31397 ( \31774 , \31323 );
not \U$31398 ( \31775 , \31342 );
or \U$31399 ( \31776 , \31774 , \31775 );
not \U$31400 ( \31777 , \31337 );
nand \U$31401 ( \31778 , \31777 , \31335 );
nand \U$31402 ( \31779 , \31776 , \31778 );
not \U$31403 ( \31780 , \1863 );
not \U$31404 ( \31781 , \19667 );
or \U$31405 ( \31782 , \31780 , \31781 );
nand \U$31406 ( \31783 , \31684 , \1910 );
nand \U$31407 ( \31784 , \31782 , \31783 );
xor \U$31408 ( \31785 , \31779 , \31784 );
not \U$31409 ( \31786 , \31785 );
not \U$31410 ( \31787 , \2249 );
xor \U$31411 ( \31788 , RIae79ac0_158, \10070 );
not \U$31412 ( \31789 , \31788 );
or \U$31413 ( \31790 , \31787 , \31789 );
nand \U$31414 ( \31791 , \31372 , \2272 );
nand \U$31415 ( \31792 , \31790 , \31791 );
not \U$31416 ( \31793 , \31792 );
not \U$31417 ( \31794 , \31793 );
and \U$31418 ( \31795 , \31786 , \31794 );
and \U$31419 ( \31796 , \31785 , \31793 );
nor \U$31420 ( \31797 , \31795 , \31796 );
not \U$31421 ( \31798 , \31374 );
not \U$31422 ( \31799 , \31365 );
or \U$31423 ( \31800 , \31798 , \31799 );
not \U$31424 ( \31801 , \31352 );
not \U$31425 ( \31802 , \31360 );
or \U$31426 ( \31803 , \31801 , \31802 );
nand \U$31427 ( \31804 , \31803 , \31346 );
nand \U$31428 ( \31805 , \31800 , \31804 );
not \U$31429 ( \31806 , \31805 );
and \U$31430 ( \31807 , \31797 , \31806 );
not \U$31431 ( \31808 , \31797 );
and \U$31432 ( \31809 , \31808 , \31805 );
nor \U$31433 ( \31810 , \31807 , \31809 );
xor \U$31434 ( \31811 , \31773 , \31810 );
not \U$31435 ( \31812 , \10700 );
and \U$31436 ( \31813 , RIae79fe8_169, \1859 );
not \U$31437 ( \31814 , RIae79fe8_169);
and \U$31438 ( \31815 , \31814 , \12502 );
or \U$31439 ( \31816 , \31813 , \31815 );
not \U$31440 ( \31817 , \31816 );
or \U$31441 ( \31818 , \31812 , \31817 );
nand \U$31442 ( \31819 , \31528 , \11914 );
nand \U$31443 ( \31820 , \31818 , \31819 );
not \U$31444 ( \31821 , \9814 );
not \U$31445 ( \31822 , RIae7a2b8_175);
not \U$31446 ( \31823 , \4112 );
or \U$31447 ( \31824 , \31822 , \31823 );
or \U$31448 ( \31825 , \2357 , RIae7a2b8_175);
nand \U$31449 ( \31826 , \31824 , \31825 );
not \U$31450 ( \31827 , \31826 );
or \U$31451 ( \31828 , \31821 , \31827 );
nand \U$31452 ( \31829 , \31652 , \9792 );
nand \U$31453 ( \31830 , \31828 , \31829 );
xor \U$31454 ( \31831 , \31820 , \31830 );
not \U$31455 ( \31832 , \9745 );
and \U$31456 ( \31833 , RIae7a060_170, \2207 );
not \U$31457 ( \31834 , RIae7a060_170);
and \U$31458 ( \31835 , \31834 , \2629 );
nor \U$31459 ( \31836 , \31833 , \31835 );
not \U$31460 ( \31837 , \31836 );
or \U$31461 ( \31838 , \31832 , \31837 );
nand \U$31462 ( \31839 , \31670 , \17797 );
nand \U$31463 ( \31840 , \31838 , \31839 );
xor \U$31464 ( \31841 , \31831 , \31840 );
xor \U$31465 ( \31842 , \31811 , \31841 );
not \U$31466 ( \31843 , \31304 );
not \U$31467 ( \31844 , \31402 );
or \U$31468 ( \31845 , \31843 , \31844 );
not \U$31469 ( \31846 , \31375 );
xor \U$31470 ( \31847 , \31313 , \31401 );
nand \U$31471 ( \31848 , \31846 , \31847 );
nand \U$31472 ( \31849 , \31845 , \31848 );
xnor \U$31473 ( \31850 , \31842 , \31849 );
not \U$31474 ( \31851 , \31606 );
not \U$31475 ( \31852 , \31585 );
not \U$31476 ( \31853 , \31852 );
not \U$31477 ( \31854 , \31594 );
or \U$31478 ( \31855 , \31853 , \31854 );
or \U$31479 ( \31856 , \31594 , \31852 );
nand \U$31480 ( \31857 , \31855 , \31856 );
not \U$31481 ( \31858 , \31857 );
or \U$31482 ( \31859 , \31851 , \31858 );
nand \U$31483 ( \31860 , \31594 , \31585 );
nand \U$31484 ( \31861 , \31859 , \31860 );
not \U$31485 ( \31862 , \31861 );
not \U$31486 ( \31863 , \10696 );
not \U$31487 ( \31864 , \31604 );
or \U$31488 ( \31865 , \31863 , \31864 );
and \U$31489 ( \31866 , RIae7a498_179, \2305 );
not \U$31490 ( \31867 , RIae7a498_179);
and \U$31491 ( \31868 , \31867 , \2309 );
or \U$31492 ( \31869 , \31866 , \31868 );
nand \U$31493 ( \31870 , \31869 , \10675 );
nand \U$31494 ( \31871 , \31865 , \31870 );
not \U$31495 ( \31872 , \9478 );
not \U$31496 ( \31873 , \12183 );
xor \U$31497 ( \31874 , RIae7a6f0_184, \31873 );
not \U$31498 ( \31875 , \31874 );
or \U$31499 ( \31876 , \31872 , \31875 );
nand \U$31500 ( \31877 , \31590 , \9473 );
nand \U$31501 ( \31878 , \31876 , \31877 );
xor \U$31502 ( \31879 , \31871 , \31878 );
not \U$31503 ( \31880 , \9776 );
not \U$31504 ( \31881 , RIae7a150_172);
not \U$31505 ( \31882 , \2140 );
or \U$31506 ( \31883 , \31881 , \31882 );
or \U$31507 ( \31884 , \2136 , RIae7a150_172);
nand \U$31508 ( \31885 , \31883 , \31884 );
not \U$31509 ( \31886 , \31885 );
or \U$31510 ( \31887 , \31880 , \31886 );
nand \U$31511 ( \31888 , \31706 , \9758 );
nand \U$31512 ( \31889 , \31887 , \31888 );
xor \U$31513 ( \31890 , \31879 , \31889 );
xor \U$31514 ( \31891 , \31862 , \31890 );
and \U$31515 ( \31892 , \31689 , \31698 );
and \U$31516 ( \31893 , \31678 , \31688 );
nor \U$31517 ( \31894 , \31892 , \31893 );
not \U$31518 ( \31895 , \12233 );
not \U$31519 ( \31896 , \17324 );
not \U$31520 ( \31897 , \6171 );
or \U$31521 ( \31898 , \31896 , \31897 );
or \U$31522 ( \31899 , \4431 , \14931 );
nand \U$31523 ( \31900 , \31898 , \31899 );
not \U$31524 ( \31901 , \31900 );
or \U$31525 ( \31902 , \31895 , \31901 );
nand \U$31526 ( \31903 , \31615 , \10927 );
nand \U$31527 ( \31904 , \31902 , \31903 );
xor \U$31528 ( \31905 , \31894 , \31904 );
not \U$31529 ( \31906 , \10275 );
and \U$31530 ( \31907 , RIae7a8d0_188, \10916 );
not \U$31531 ( \31908 , RIae7a8d0_188);
and \U$31532 ( \31909 , \31908 , \1186 );
nor \U$31533 ( \31910 , \31907 , \31909 );
not \U$31534 ( \31911 , \31910 );
or \U$31535 ( \31912 , \31906 , \31911 );
nand \U$31536 ( \31913 , \31458 , \11205 );
nand \U$31537 ( \31914 , \31912 , \31913 );
xnor \U$31538 ( \31915 , \31905 , \31914 );
xnor \U$31539 ( \31916 , \31891 , \31915 );
xor \U$31540 ( \31917 , \31850 , \31916 );
not \U$31541 ( \31918 , \31257 );
xor \U$31542 ( \31919 , \31242 , \31248 );
not \U$31543 ( \31920 , \31919 );
or \U$31544 ( \31921 , \31918 , \31920 );
nand \U$31545 ( \31922 , \31248 , \31242 );
nand \U$31546 ( \31923 , \31921 , \31922 );
xnor \U$31547 ( \31924 , \31917 , \31923 );
not \U$31548 ( \31925 , \31264 );
not \U$31549 ( \31926 , \31276 );
not \U$31550 ( \31927 , \31926 );
or \U$31551 ( \31928 , \31925 , \31927 );
not \U$31552 ( \31929 , \31276 );
not \U$31553 ( \31930 , \31263 );
or \U$31554 ( \31931 , \31929 , \31930 );
not \U$31555 ( \31932 , \31258 );
nand \U$31556 ( \31933 , \31931 , \31932 );
nand \U$31557 ( \31934 , \31928 , \31933 );
xor \U$31558 ( \31935 , \31924 , \31934 );
not \U$31559 ( \31936 , \31451 );
xnor \U$31560 ( \31937 , \31430 , \31532 );
not \U$31561 ( \31938 , \31937 );
or \U$31562 ( \31939 , \31936 , \31938 );
not \U$31563 ( \31940 , \31532 );
nand \U$31564 ( \31941 , \31940 , \31430 );
nand \U$31565 ( \31942 , \31939 , \31941 );
not \U$31566 ( \31943 , \31298 );
not \U$31567 ( \31944 , \31420 );
or \U$31568 ( \31945 , \31943 , \31944 );
not \U$31569 ( \31946 , \31403 );
nand \U$31570 ( \31947 , \31946 , \31416 );
nand \U$31571 ( \31948 , \31945 , \31947 );
not \U$31572 ( \31949 , \31948 );
not \U$31573 ( \31950 , \2011 );
and \U$31574 ( \31951 , RIae79610_148, \10740 );
not \U$31575 ( \31952 , RIae79610_148);
and \U$31576 ( \31953 , \31952 , \10743 );
or \U$31577 ( \31954 , \31951 , \31953 );
not \U$31578 ( \31955 , \31954 );
or \U$31579 ( \31956 , \31950 , \31955 );
nand \U$31580 ( \31957 , \31696 , \2063 );
nand \U$31581 ( \31958 , \31956 , \31957 );
not \U$31582 ( \31959 , \1820 );
not \U$31583 ( \31960 , RIae79688_149);
not \U$31584 ( \31961 , \10749 );
or \U$31585 ( \31962 , \31960 , \31961 );
or \U$31586 ( \31963 , \10749 , RIae79688_149);
nand \U$31587 ( \31964 , \31962 , \31963 );
not \U$31588 ( \31965 , \31964 );
or \U$31589 ( \31966 , \31959 , \31965 );
nand \U$31590 ( \31967 , \31384 , \1843 );
nand \U$31591 ( \31968 , \31966 , \31967 );
not \U$31592 ( \31969 , \31968 );
xor \U$31593 ( \31970 , \31958 , \31969 );
not \U$31594 ( \31971 , \10223 );
not \U$31595 ( \31972 , \2183 );
not \U$31596 ( \31973 , \28019 );
or \U$31597 ( \31974 , \31972 , \31973 );
or \U$31598 ( \31975 , \28019 , \2183 );
nand \U$31599 ( \31976 , \31974 , \31975 );
not \U$31600 ( \31977 , \31976 );
or \U$31601 ( \31978 , \31971 , \31977 );
nand \U$31602 ( \31979 , \31351 , \2188 );
nand \U$31603 ( \31980 , \31978 , \31979 );
xnor \U$31604 ( \31981 , \31970 , \31980 );
not \U$31605 ( \31982 , \31981 );
not \U$31606 ( \31983 , \31313 );
not \U$31607 ( \31984 , \31400 );
or \U$31608 ( \31985 , \31983 , \31984 );
not \U$31609 ( \31986 , \31398 );
nand \U$31610 ( \31987 , \31986 , \31386 );
nand \U$31611 ( \31988 , \31985 , \31987 );
not \U$31612 ( \31989 , \31988 );
not \U$31613 ( \31990 , \31989 );
or \U$31614 ( \31991 , \31982 , \31990 );
or \U$31615 ( \31992 , \31989 , \31981 );
nand \U$31616 ( \31993 , \31991 , \31992 );
not \U$31617 ( \31994 , \31578 );
not \U$31618 ( \31995 , \31561 );
nand \U$31619 ( \31996 , \31995 , \31562 , \31567 );
not \U$31620 ( \31997 , \31996 );
or \U$31621 ( \31998 , \31994 , \31997 );
nand \U$31622 ( \31999 , \31568 , \31561 );
nand \U$31623 ( \32000 , \31998 , \31999 );
xnor \U$31624 ( \32001 , \31993 , \32000 );
not \U$31625 ( \32002 , \31233 );
nand \U$31626 ( \32003 , \32002 , \31226 );
not \U$31627 ( \32004 , \32003 );
not \U$31628 ( \32005 , \31241 );
or \U$31629 ( \32006 , \32004 , \32005 );
nand \U$31630 ( \32007 , \31233 , \31227 );
nand \U$31631 ( \32008 , \32006 , \32007 );
xor \U$31632 ( \32009 , \32001 , \32008 );
nor \U$31633 ( \32010 , \31444 , \31435 );
or \U$31634 ( \32011 , \31450 , \32010 );
nand \U$31635 ( \32012 , \31444 , \31435 );
nand \U$31636 ( \32013 , \32011 , \32012 );
not \U$31637 ( \32014 , \32013 );
and \U$31638 ( \32015 , \32009 , \32014 );
not \U$31639 ( \32016 , \32009 );
and \U$31640 ( \32017 , \32016 , \32013 );
nor \U$31641 ( \32018 , \32015 , \32017 );
and \U$31642 ( \32019 , \31949 , \32018 );
not \U$31643 ( \32020 , \31949 );
not \U$31644 ( \32021 , \32018 );
and \U$31645 ( \32022 , \32020 , \32021 );
nor \U$31646 ( \32023 , \32019 , \32022 );
xnor \U$31647 ( \32024 , \31942 , \32023 );
xnor \U$31648 ( \32025 , \31935 , \32024 );
and \U$31649 ( \32026 , \31763 , \31764 , \32025 );
not \U$31650 ( \32027 , \32026 );
not \U$31651 ( \32028 , \31764 );
not \U$31652 ( \32029 , \31763 );
or \U$31653 ( \32030 , \32028 , \32029 );
not \U$31654 ( \32031 , \32025 );
nand \U$31655 ( \32032 , \32030 , \32031 );
nand \U$31656 ( \32033 , \32027 , \32032 );
not \U$31657 ( \32034 , \31425 );
not \U$31658 ( \32035 , \31541 );
or \U$31659 ( \32036 , \32034 , \32035 );
not \U$31660 ( \32037 , \31425 );
not \U$31661 ( \32038 , \32037 );
not \U$31662 ( \32039 , \31540 );
or \U$31663 ( \32040 , \32038 , \32039 );
not \U$31664 ( \32041 , \31533 );
nand \U$31665 ( \32042 , \32040 , \32041 );
nand \U$31666 ( \32043 , \32036 , \32042 );
not \U$31667 ( \32044 , \31639 );
nand \U$31668 ( \32045 , \32044 , \31720 );
not \U$31669 ( \32046 , \32045 );
not \U$31670 ( \32047 , \31726 );
or \U$31671 ( \32048 , \32046 , \32047 );
nand \U$31672 ( \32049 , \31721 , \31639 );
nand \U$31673 ( \32050 , \32048 , \32049 );
not \U$31674 ( \32051 , \32050 );
not \U$31675 ( \32052 , \31579 );
not \U$31676 ( \32053 , \32052 );
not \U$31677 ( \32054 , \31638 );
or \U$31678 ( \32055 , \32053 , \32054 );
not \U$31679 ( \32056 , \31607 );
nand \U$31680 ( \32057 , \32055 , \32056 );
not \U$31681 ( \32058 , \31638 );
nand \U$31682 ( \32059 , \32058 , \31579 );
and \U$31683 ( \32060 , \32057 , \32059 );
not \U$31684 ( \32061 , \31486 );
not \U$31685 ( \32062 , \32061 );
not \U$31686 ( \32063 , \31462 );
or \U$31687 ( \32064 , \32062 , \32063 );
not \U$31688 ( \32065 , \31482 );
nand \U$31689 ( \32066 , \32065 , \31474 );
nand \U$31690 ( \32067 , \32064 , \32066 );
not \U$31691 ( \32068 , \31530 );
and \U$31692 ( \32069 , \31520 , \31509 );
not \U$31693 ( \32070 , \31520 );
and \U$31694 ( \32071 , \32070 , \31508 );
nor \U$31695 ( \32072 , \32069 , \32071 );
not \U$31696 ( \32073 , \32072 );
or \U$31697 ( \32074 , \32068 , \32073 );
nand \U$31698 ( \32075 , \31519 , \31508 );
nand \U$31699 ( \32076 , \32074 , \32075 );
not \U$31700 ( \32077 , \32076 );
xor \U$31701 ( \32078 , \32067 , \32077 );
xor \U$31702 ( \32079 , \31617 , \31626 );
and \U$31703 ( \32080 , \32079 , \31637 );
and \U$31704 ( \32081 , \31617 , \31626 );
or \U$31705 ( \32082 , \32080 , \32081 );
xnor \U$31706 ( \32083 , \32078 , \32082 );
xor \U$31707 ( \32084 , \32060 , \32083 );
or \U$31708 ( \32085 , \31719 , \31644 );
nand \U$31709 ( \32086 , \32085 , \31675 );
nand \U$31710 ( \32087 , \31719 , \31644 );
nand \U$31711 ( \32088 , \32086 , \32087 );
xnor \U$31712 ( \32089 , \32084 , \32088 );
not \U$31713 ( \32090 , \32089 );
or \U$31714 ( \32091 , \32051 , \32090 );
or \U$31715 ( \32092 , \32050 , \32089 );
nand \U$31716 ( \32093 , \32091 , \32092 );
not \U$31717 ( \32094 , \32093 );
not \U$31718 ( \32095 , \2007 );
and \U$31719 ( \32096 , RIae797f0_152, \9442 );
not \U$31720 ( \32097 , RIae797f0_152);
and \U$31721 ( \32098 , \32097 , \9438 );
or \U$31722 ( \32099 , \32096 , \32098 );
not \U$31723 ( \32100 , \32099 );
or \U$31724 ( \32101 , \32095 , \32100 );
nand \U$31725 ( \32102 , \31566 , \1988 );
nand \U$31726 ( \32103 , \32101 , \32102 );
not \U$31727 ( \32104 , \2322 );
not \U$31728 ( \32105 , RIae798e0_154);
not \U$31729 ( \32106 , \10937 );
or \U$31730 ( \32107 , \32105 , \32106 );
or \U$31731 ( \32108 , \16766 , RIae798e0_154);
nand \U$31732 ( \32109 , \32107 , \32108 );
not \U$31733 ( \32110 , \32109 );
or \U$31734 ( \32111 , \32104 , \32110 );
nand \U$31735 ( \32112 , \31557 , \10807 );
nand \U$31736 ( \32113 , \32111 , \32112 );
not \U$31737 ( \32114 , \32113 );
xor \U$31738 ( \32115 , \32103 , \32114 );
not \U$31739 ( \32116 , \2450 );
xor \U$31740 ( \32117 , RIae79778_151, \9350 );
not \U$31741 ( \32118 , \32117 );
or \U$31742 ( \32119 , \32116 , \32118 );
nand \U$31743 ( \32120 , \31309 , \9576 );
nand \U$31744 ( \32121 , \32119 , \32120 );
xnor \U$31745 ( \32122 , \32115 , \32121 );
not \U$31746 ( \32123 , \1919 );
not \U$31747 ( \32124 , \3810 );
not \U$31748 ( \32125 , \12482 );
or \U$31749 ( \32126 , \32124 , \32125 );
or \U$31750 ( \32127 , \9607 , \3039 );
nand \U$31751 ( \32128 , \32126 , \32127 );
not \U$31752 ( \32129 , \32128 );
or \U$31753 ( \32130 , \32123 , \32129 );
nand \U$31754 ( \32131 , \31393 , \1932 );
nand \U$31755 ( \32132 , \32130 , \32131 );
not \U$31756 ( \32133 , \2776 );
and \U$31757 ( \32134 , RIae79c28_161, \16260 );
not \U$31758 ( \32135 , RIae79c28_161);
and \U$31759 ( \32136 , \32135 , \9298 );
or \U$31760 ( \32137 , \32134 , \32136 );
not \U$31761 ( \32138 , \32137 );
or \U$31762 ( \32139 , \32133 , \32138 );
nand \U$31763 ( \32140 , \31576 , \2417 );
nand \U$31764 ( \32141 , \32139 , \32140 );
xor \U$31765 ( \32142 , \32132 , \32141 );
not \U$31766 ( \32143 , \10573 );
xor \U$31767 ( \32144 , RIae79ef8_167, \10328 );
not \U$31768 ( \32145 , \32144 );
or \U$31769 ( \32146 , \32143 , \32145 );
nand \U$31770 ( \32147 , \31517 , \19362 );
nand \U$31771 ( \32148 , \32146 , \32147 );
xor \U$31772 ( \32149 , \32142 , \32148 );
xor \U$31773 ( \32150 , \32122 , \32149 );
not \U$31774 ( \32151 , \9527 );
and \U$31775 ( \32152 , RIae7a7e0_186, \16561 );
not \U$31776 ( \32153 , RIae7a7e0_186);
and \U$31777 ( \32154 , \32153 , \5162 );
or \U$31778 ( \32155 , \32152 , \32154 );
not \U$31779 ( \32156 , \32155 );
or \U$31780 ( \32157 , \32151 , \32156 );
nand \U$31781 ( \32158 , \31635 , \11851 );
nand \U$31782 ( \32159 , \32157 , \32158 );
not \U$31783 ( \32160 , \13121 );
and \U$31784 ( \32161 , RIae7a240_174, \2676 );
not \U$31785 ( \32162 , RIae7a240_174);
and \U$31786 ( \32163 , \32162 , \4837 );
or \U$31787 ( \32164 , \32161 , \32163 );
not \U$31788 ( \32165 , \32164 );
or \U$31789 ( \32166 , \32160 , \32165 );
nand \U$31790 ( \32167 , \31661 , \13130 );
nand \U$31791 ( \32168 , \32166 , \32167 );
xor \U$31792 ( \32169 , \32159 , \32168 );
not \U$31793 ( \32170 , \11014 );
not \U$31794 ( \32171 , \31622 );
or \U$31795 ( \32172 , \32170 , \32171 );
xor \U$31796 ( \32173 , RIae7a3a8_177, \1808 );
nand \U$31797 ( \32174 , \32173 , \9621 );
nand \U$31798 ( \32175 , \32172 , \32174 );
xor \U$31799 ( \32176 , \32169 , \32175 );
xor \U$31800 ( \32177 , \32150 , \32176 );
not \U$31801 ( \32178 , \1501 );
not \U$31802 ( \32179 , \19693 );
or \U$31803 ( \32180 , \32178 , \32179 );
nand \U$31804 ( \32181 , \31319 , \1497 );
nand \U$31805 ( \32182 , \32180 , \32181 );
not \U$31806 ( \32183 , \19683 );
not \U$31807 ( \32184 , \19676 );
and \U$31808 ( \32185 , \32183 , \32184 );
and \U$31809 ( \32186 , \19683 , \19676 );
nor \U$31810 ( \32187 , \32185 , \32186 );
not \U$31811 ( \32188 , \32187 );
not \U$31812 ( \32189 , \1012 );
not \U$31813 ( \32190 , \18973 );
or \U$31814 ( \32191 , \32189 , \32190 );
nand \U$31815 ( \32192 , \31331 , \1007 );
nand \U$31816 ( \32193 , \32191 , \32192 );
not \U$31817 ( \32194 , \32193 );
or \U$31818 ( \32195 , \32188 , \32194 );
or \U$31819 ( \32196 , \32193 , \32187 );
nand \U$31820 ( \32197 , \32195 , \32196 );
xor \U$31821 ( \32198 , \32182 , \32197 );
not \U$31822 ( \32199 , \4853 );
and \U$31823 ( \32200 , RIae79ca0_162, \12700 );
not \U$31824 ( \32201 , RIae79ca0_162);
and \U$31825 ( \32202 , \32201 , \9280 );
or \U$31826 ( \32203 , \32200 , \32202 );
not \U$31827 ( \32204 , \32203 );
or \U$31828 ( \32205 , \32199 , \32204 );
nand \U$31829 ( \32206 , \31472 , \4842 );
nand \U$31830 ( \32207 , \32205 , \32206 );
xor \U$31831 ( \32208 , \32198 , \32207 );
not \U$31832 ( \32209 , \5048 );
and \U$31833 ( \32210 , RIae79d90_164, \4960 );
not \U$31834 ( \32211 , RIae79d90_164);
and \U$31835 ( \32212 , \32211 , \17009 );
or \U$31836 ( \32213 , \32210 , \32212 );
not \U$31837 ( \32214 , \32213 );
or \U$31838 ( \32215 , \32209 , \32214 );
nand \U$31839 ( \32216 , \31504 , \6091 );
nand \U$31840 ( \32217 , \32215 , \32216 );
xor \U$31841 ( \32218 , \32208 , \32217 );
nand \U$31842 ( \32219 , \31711 , \31700 );
not \U$31843 ( \32220 , \32219 );
not \U$31844 ( \32221 , \31718 );
or \U$31845 ( \32222 , \32220 , \32221 );
not \U$31846 ( \32223 , \31700 );
nand \U$31847 ( \32224 , \32223 , \31710 );
nand \U$31848 ( \32225 , \32222 , \32224 );
not \U$31849 ( \32226 , \32225 );
not \U$31850 ( \32227 , \32226 );
xor \U$31851 ( \32228 , \32218 , \32227 );
xor \U$31852 ( \32229 , \31654 , \31663 );
and \U$31853 ( \32230 , \32229 , \31674 );
and \U$31854 ( \32231 , \31654 , \31663 );
or \U$31855 ( \32232 , \32230 , \32231 );
xnor \U$31856 ( \32233 , \32228 , \32232 );
xor \U$31857 ( \32234 , \32177 , \32233 );
not \U$31858 ( \32235 , \31497 );
not \U$31859 ( \32236 , \31531 );
and \U$31860 ( \32237 , \31490 , \32236 );
not \U$31861 ( \32238 , \31490 );
and \U$31862 ( \32239 , \32238 , \31531 );
nor \U$31863 ( \32240 , \32237 , \32239 );
not \U$31864 ( \32241 , \32240 );
or \U$31865 ( \32242 , \32235 , \32241 );
nand \U$31866 ( \32243 , \32236 , \31490 );
nand \U$31867 ( \32244 , \32242 , \32243 );
xor \U$31868 ( \32245 , \32234 , \32244 );
not \U$31869 ( \32246 , \32245 );
and \U$31870 ( \32247 , \32094 , \32246 );
and \U$31871 ( \32248 , \32093 , \32245 );
nor \U$31872 ( \32249 , \32247 , \32248 );
not \U$31873 ( \32250 , \32249 );
xor \U$31874 ( \32251 , \32043 , \32250 );
not \U$31875 ( \32252 , \31728 );
nand \U$31876 ( \32253 , \32252 , \31734 );
not \U$31877 ( \32254 , \32253 );
not \U$31878 ( \32255 , \31746 );
or \U$31879 ( \32256 , \32254 , \32255 );
not \U$31880 ( \32257 , \31734 );
nand \U$31881 ( \32258 , \32257 , \31728 );
nand \U$31882 ( \32259 , \32256 , \32258 );
xor \U$31883 ( \32260 , \32251 , \32259 );
not \U$31884 ( \32261 , \32260 );
and \U$31885 ( \32262 , \32033 , \32261 );
not \U$31886 ( \32263 , \32033 );
and \U$31887 ( \32264 , \32263 , \32260 );
nor \U$31888 ( \32265 , \32262 , \32264 );
not \U$31889 ( \32266 , \32265 );
not \U$31890 ( \32267 , \31543 );
not \U$31891 ( \32268 , \31751 );
or \U$31892 ( \32269 , \32267 , \32268 );
nand \U$31893 ( \32270 , \31747 , \31548 , \31550 );
nand \U$31894 ( \32271 , \32269 , \32270 );
not \U$31895 ( \32272 , \32271 );
nand \U$31896 ( \32273 , \32266 , \32272 );
nand \U$31897 ( \32274 , \31214 , \31759 , \32273 );
not \U$31898 ( \32275 , \32274 );
not \U$31899 ( \32276 , \32275 );
or \U$31900 ( \32277 , \31211 , \32276 );
nand \U$31901 ( \32278 , \31757 , \31220 );
not \U$31902 ( \32279 , \32278 );
nand \U$31903 ( \32280 , \32265 , \32271 );
not \U$31904 ( \32281 , \32280 );
or \U$31905 ( \32282 , \32279 , \32281 );
buf \U$31906 ( \32283 , \32273 );
nand \U$31907 ( \32284 , \32282 , \32283 );
nand \U$31908 ( \32285 , \32277 , \32284 );
nand \U$31909 ( \32286 , \31179 , \31208 );
and \U$31910 ( \32287 , \32286 , \31177 );
xor \U$31911 ( \32288 , \30803 , \30790 );
xor \U$31912 ( \32289 , \30890 , \30899 );
xor \U$31913 ( \32290 , \32289 , \30910 );
not \U$31914 ( \32291 , \32290 );
not \U$31915 ( \32292 , \31026 );
not \U$31916 ( \32293 , \30984 );
not \U$31917 ( \32294 , \32293 );
or \U$31918 ( \32295 , \32292 , \32294 );
or \U$31919 ( \32296 , \32293 , \31026 );
nand \U$31920 ( \32297 , \32295 , \32296 );
not \U$31921 ( \32298 , \32297 );
not \U$31922 ( \32299 , \10676 );
not \U$31923 ( \32300 , \31069 );
or \U$31924 ( \32301 , \32299 , \32300 );
and \U$31925 ( \32302 , \10625 , \10492 );
not \U$31926 ( \32303 , \10625 );
and \U$31927 ( \32304 , \32303 , \3273 );
nor \U$31928 ( \32305 , \32302 , \32304 );
nand \U$31929 ( \32306 , \32305 , \11434 );
nand \U$31930 ( \32307 , \32301 , \32306 );
not \U$31931 ( \32308 , \32307 );
nand \U$31932 ( \32309 , \32298 , \32308 );
not \U$31933 ( \32310 , \32309 );
not \U$31934 ( \32311 , \9478 );
not \U$31935 ( \32312 , \30825 );
or \U$31936 ( \32313 , \32311 , \32312 );
not \U$31937 ( \32314 , \16101 );
not \U$31938 ( \32315 , \1759 );
or \U$31939 ( \32316 , \32314 , \32315 );
or \U$31940 ( \32317 , \4584 , \28731 );
nand \U$31941 ( \32318 , \32316 , \32317 );
nand \U$31942 ( \32319 , \32318 , \9473 );
nand \U$31943 ( \32320 , \32313 , \32319 );
not \U$31944 ( \32321 , \32320 );
or \U$31945 ( \32322 , \32310 , \32321 );
nand \U$31946 ( \32323 , \32297 , \32307 );
nand \U$31947 ( \32324 , \32322 , \32323 );
not \U$31948 ( \32325 , \30847 );
not \U$31949 ( \32326 , \30872 );
or \U$31950 ( \32327 , \32325 , \32326 );
or \U$31951 ( \32328 , \30847 , \30872 );
nand \U$31952 ( \32329 , \32327 , \32328 );
xor \U$31953 ( \32330 , \32324 , \32329 );
not \U$31954 ( \32331 , \32330 );
or \U$31955 ( \32332 , \32291 , \32331 );
nand \U$31956 ( \32333 , \32329 , \32324 );
nand \U$31957 ( \32334 , \32332 , \32333 );
not \U$31958 ( \32335 , \30792 );
not \U$31959 ( \32336 , \30801 );
or \U$31960 ( \32337 , \32335 , \32336 );
or \U$31961 ( \32338 , \30801 , \30792 );
nand \U$31962 ( \32339 , \32337 , \32338 );
and \U$31963 ( \32340 , \32339 , \30795 );
not \U$31964 ( \32341 , \32339 );
and \U$31965 ( \32342 , \32341 , \30794 );
nor \U$31966 ( \32343 , \32340 , \32342 );
xor \U$31967 ( \32344 , \32334 , \32343 );
xor \U$31968 ( \32345 , \30840 , \30917 );
and \U$31969 ( \32346 , \32344 , \32345 );
and \U$31970 ( \32347 , \32334 , \32343 );
or \U$31971 ( \32348 , \32346 , \32347 );
xor \U$31972 ( \32349 , \32288 , \32348 );
xor \U$31973 ( \32350 , \30922 , \30932 );
and \U$31974 ( \32351 , \32349 , \32350 );
and \U$31975 ( \32352 , \32288 , \32348 );
nor \U$31976 ( \32353 , \32351 , \32352 );
not \U$31977 ( \32354 , \32353 );
xor \U$31978 ( \32355 , \31101 , \31108 );
xor \U$31979 ( \32356 , \32355 , \31131 );
not \U$31980 ( \32357 , \32356 );
not \U$31981 ( \32358 , \11205 );
xor \U$31982 ( \32359 , \3748 , RIae7a8d0_188);
not \U$31983 ( \32360 , \32359 );
or \U$31984 ( \32361 , \32358 , \32360 );
nand \U$31985 ( \32362 , \30888 , \10275 );
nand \U$31986 ( \32363 , \32361 , \32362 );
not \U$31987 ( \32364 , \32363 );
not \U$31988 ( \32365 , \9776 );
not \U$31989 ( \32366 , \30832 );
or \U$31990 ( \32367 , \32365 , \32366 );
and \U$31991 ( \32368 , RIae7a150_172, \14422 );
not \U$31992 ( \32369 , RIae7a150_172);
and \U$31993 ( \32370 , \32369 , \1969 );
or \U$31994 ( \32371 , \32368 , \32370 );
not \U$31995 ( \32372 , \32371 );
nand \U$31996 ( \32373 , \32372 , \10667 );
nand \U$31997 ( \32374 , \32367 , \32373 );
not \U$31998 ( \32375 , \9745 );
not \U$31999 ( \32376 , \30895 );
or \U$32000 ( \32377 , \32375 , \32376 );
and \U$32001 ( \32378 , RIae7a060_170, \2093 );
not \U$32002 ( \32379 , RIae7a060_170);
and \U$32003 ( \32380 , \32379 , \13008 );
nor \U$32004 ( \32381 , \32378 , \32380 );
nand \U$32005 ( \32382 , \32381 , \9728 );
nand \U$32006 ( \32383 , \32377 , \32382 );
xor \U$32007 ( \32384 , \32374 , \32383 );
not \U$32008 ( \32385 , \32384 );
or \U$32009 ( \32386 , \32364 , \32385 );
nand \U$32010 ( \32387 , \32383 , \32374 );
nand \U$32011 ( \32388 , \32386 , \32387 );
not \U$32012 ( \32389 , \32388 );
buf \U$32013 ( \32390 , \30700 );
xor \U$32014 ( \32391 , \30711 , \32390 );
xor \U$32015 ( \32392 , \30764 , \30773 );
xor \U$32016 ( \32393 , \32392 , \30780 );
xor \U$32017 ( \32394 , \32391 , \32393 );
not \U$32018 ( \32395 , \32394 );
or \U$32019 ( \32396 , \32389 , \32395 );
nand \U$32020 ( \32397 , \32393 , \32391 );
nand \U$32021 ( \32398 , \32396 , \32397 );
not \U$32022 ( \32399 , \32398 );
xor \U$32023 ( \32400 , \30783 , \30715 );
buf \U$32024 ( \32401 , \30754 );
not \U$32025 ( \32402 , \32401 );
and \U$32026 ( \32403 , \32400 , \32402 );
not \U$32027 ( \32404 , \32400 );
and \U$32028 ( \32405 , \32404 , \32401 );
nor \U$32029 ( \32406 , \32403 , \32405 );
not \U$32030 ( \32407 , \32406 );
not \U$32031 ( \32408 , \9699 );
not \U$32032 ( \32409 , \30771 );
or \U$32033 ( \32410 , \32408 , \32409 );
and \U$32034 ( \32411 , RIae7a240_174, \15117 );
not \U$32035 ( \32412 , RIae7a240_174);
and \U$32036 ( \32413 , \32412 , \9290 );
or \U$32037 ( \32414 , \32411 , \32413 );
nand \U$32038 ( \32415 , \32414 , \13720 );
nand \U$32039 ( \32416 , \32410 , \32415 );
not \U$32040 ( \32417 , \9622 );
not \U$32041 ( \32418 , \30746 );
or \U$32042 ( \32419 , \32417 , \32418 );
and \U$32043 ( \32420 , RIae7a3a8_177, \13248 );
not \U$32044 ( \32421 , RIae7a3a8_177);
and \U$32045 ( \32422 , \32421 , \16311 );
or \U$32046 ( \32423 , \32420 , \32422 );
nand \U$32047 ( \32424 , \32423 , \9644 );
nand \U$32048 ( \32425 , \32419 , \32424 );
xor \U$32049 ( \32426 , \32416 , \32425 );
and \U$32050 ( \32427 , \4169 , RIae7a510_180);
not \U$32051 ( \32428 , \4169 );
and \U$32052 ( \32429 , \32428 , \17324 );
nor \U$32053 ( \32430 , \32427 , \32429 );
not \U$32054 ( \32431 , \32430 );
not \U$32055 ( \32432 , \10927 );
or \U$32056 ( \32433 , \32431 , \32432 );
nand \U$32057 ( \32434 , \30776 , \12233 );
nand \U$32058 ( \32435 , \32433 , \32434 );
and \U$32059 ( \32436 , \32426 , \32435 );
and \U$32060 ( \32437 , \32416 , \32425 );
or \U$32061 ( \32438 , \32436 , \32437 );
not \U$32062 ( \32439 , \32438 );
not \U$32063 ( \32440 , \32439 );
not \U$32064 ( \32441 , \4853 );
not \U$32065 ( \32442 , \30866 );
not \U$32066 ( \32443 , \32442 );
or \U$32067 ( \32444 , \32441 , \32443 );
and \U$32068 ( \32445 , \10464 , \4844 );
not \U$32069 ( \32446 , \10464 );
and \U$32070 ( \32447 , \32446 , RIae79ca0_162);
nor \U$32071 ( \32448 , \32445 , \32447 );
nand \U$32072 ( \32449 , \32448 , \11761 );
nand \U$32073 ( \32450 , \32444 , \32449 );
not \U$32074 ( \32451 , \10510 );
and \U$32075 ( \32452 , RIae7a7e0_186, \2576 );
not \U$32076 ( \32453 , RIae7a7e0_186);
and \U$32077 ( \32454 , \32453 , \1789 );
nor \U$32078 ( \32455 , \32452 , \32454 );
not \U$32079 ( \32456 , \32455 );
or \U$32080 ( \32457 , \32451 , \32456 );
nand \U$32081 ( \32458 , \30843 , \29519 );
nand \U$32082 ( \32459 , \32457 , \32458 );
xor \U$32083 ( \32460 , \32450 , \32459 );
not \U$32084 ( \32461 , RIae7aab0_192);
not \U$32085 ( \32462 , \30906 );
or \U$32086 ( \32463 , \32461 , \32462 );
not \U$32087 ( \32464 , RIae7aa38_191);
not \U$32088 ( \32465 , \26330 );
or \U$32089 ( \32466 , \32464 , \32465 );
or \U$32090 ( \32467 , \13142 , RIae7aa38_191);
nand \U$32091 ( \32468 , \32466 , \32467 );
nand \U$32092 ( \32469 , \32468 , \14667 );
nand \U$32093 ( \32470 , \32463 , \32469 );
and \U$32094 ( \32471 , \32460 , \32470 );
and \U$32095 ( \32472 , \32450 , \32459 );
or \U$32096 ( \32473 , \32471 , \32472 );
not \U$32097 ( \32474 , \32473 );
not \U$32098 ( \32475 , \10700 );
not \U$32099 ( \32476 , \30707 );
or \U$32100 ( \32477 , \32475 , \32476 );
not \U$32101 ( \32478 , \11918 );
not \U$32102 ( \32479 , \9363 );
or \U$32103 ( \32480 , \32478 , \32479 );
not \U$32104 ( \32481 , \16254 );
or \U$32105 ( \32482 , \32481 , \11069 );
nand \U$32106 ( \32483 , \32480 , \32482 );
nand \U$32107 ( \32484 , \32483 , \10709 );
nand \U$32108 ( \32485 , \32477 , \32484 );
not \U$32109 ( \32486 , \32485 );
not \U$32110 ( \32487 , \16135 );
not \U$32111 ( \32488 , \30760 );
or \U$32112 ( \32489 , \32487 , \32488 );
and \U$32113 ( \32490 , RIae7a2b8_175, \19661 );
not \U$32114 ( \32491 , RIae7a2b8_175);
and \U$32115 ( \32492 , \32491 , \16274 );
or \U$32116 ( \32493 , \32490 , \32492 );
nand \U$32117 ( \32494 , \32493 , \9792 );
nand \U$32118 ( \32495 , \32489 , \32494 );
not \U$32119 ( \32496 , \32495 );
xor \U$32120 ( \32497 , \30690 , \30679 );
not \U$32121 ( \32498 , \32497 );
and \U$32122 ( \32499 , \32496 , \32498 );
not \U$32123 ( \32500 , \32496 );
and \U$32124 ( \32501 , \32500 , \32497 );
nor \U$32125 ( \32502 , \32499 , \32501 );
not \U$32126 ( \32503 , \32502 );
or \U$32127 ( \32504 , \32486 , \32503 );
not \U$32128 ( \32505 , \32496 );
nand \U$32129 ( \32506 , \32505 , \32497 );
nand \U$32130 ( \32507 , \32504 , \32506 );
not \U$32131 ( \32508 , \32507 );
nand \U$32132 ( \32509 , \32474 , \32508 );
nand \U$32133 ( \32510 , \32440 , \32509 );
nand \U$32134 ( \32511 , \32473 , \32507 );
nand \U$32135 ( \32512 , \32510 , \32511 );
not \U$32136 ( \32513 , \32512 );
or \U$32137 ( \32514 , \32407 , \32513 );
or \U$32138 ( \32515 , \32512 , \32406 );
nand \U$32139 ( \32516 , \32514 , \32515 );
not \U$32140 ( \32517 , \32516 );
or \U$32141 ( \32518 , \32399 , \32517 );
not \U$32142 ( \32519 , \32406 );
nand \U$32143 ( \32520 , \32519 , \32512 );
nand \U$32144 ( \32521 , \32518 , \32520 );
not \U$32145 ( \32522 , \32521 );
not \U$32146 ( \32523 , \6214 );
not \U$32147 ( \32524 , \30654 );
or \U$32148 ( \32525 , \32523 , \32524 );
not \U$32149 ( \32526 , \9455 );
and \U$32150 ( \32527 , RIae79ef8_167, \32526 );
not \U$32151 ( \32528 , RIae79ef8_167);
and \U$32152 ( \32529 , \32528 , \9459 );
or \U$32153 ( \32530 , \32527 , \32529 );
nand \U$32154 ( \32531 , \32530 , \19362 );
nand \U$32155 ( \32532 , \32525 , \32531 );
not \U$32156 ( \32533 , \2339 );
not \U$32157 ( \32534 , \11589 );
and \U$32158 ( \32535 , RIae798e0_154, \32534 );
not \U$32159 ( \32536 , RIae798e0_154);
and \U$32160 ( \32537 , \32536 , \10337 );
nor \U$32161 ( \32538 , \32535 , \32537 );
not \U$32162 ( \32539 , \32538 );
or \U$32163 ( \32540 , \32533 , \32539 );
nand \U$32164 ( \32541 , \31035 , \2321 );
nand \U$32165 ( \32542 , \32540 , \32541 );
not \U$32166 ( \32543 , \32542 );
or \U$32167 ( \32544 , RIae79520_146, RIae79a48_157);
nand \U$32168 ( \32545 , \32544 , \12857 );
nand \U$32169 ( \32546 , \32545 , \7625 );
not \U$32170 ( \32547 , \32546 );
not \U$32171 ( \32548 , \2271 );
not \U$32172 ( \32549 , \2268 );
not \U$32173 ( \32550 , \12857 );
or \U$32174 ( \32551 , \32549 , \32550 );
or \U$32175 ( \32552 , \12857 , \10419 );
nand \U$32176 ( \32553 , \32551 , \32552 );
not \U$32177 ( \32554 , \32553 );
or \U$32178 ( \32555 , \32548 , \32554 );
nand \U$32179 ( \32556 , \31006 , \2249 );
nand \U$32180 ( \32557 , \32555 , \32556 );
nand \U$32181 ( \32558 , \32547 , \32557 );
not \U$32182 ( \32559 , \32558 );
not \U$32183 ( \32560 , \1919 );
not \U$32184 ( \32561 , \30686 );
or \U$32185 ( \32562 , \32560 , \32561 );
and \U$32186 ( \32563 , RIae794a8_145, \19689 );
not \U$32187 ( \32564 , RIae794a8_145);
not \U$32188 ( \32565 , \11581 );
and \U$32189 ( \32566 , \32564 , \32565 );
or \U$32190 ( \32567 , \32563 , \32566 );
nand \U$32191 ( \32568 , \32567 , \1932 );
nand \U$32192 ( \32569 , \32562 , \32568 );
not \U$32193 ( \32570 , \32569 );
or \U$32194 ( \32571 , \32559 , \32570 );
or \U$32195 ( \32572 , \32569 , \32558 );
nand \U$32196 ( \32573 , \32571 , \32572 );
not \U$32197 ( \32574 , \32573 );
or \U$32198 ( \32575 , \32543 , \32574 );
not \U$32199 ( \32576 , \32558 );
nand \U$32200 ( \32577 , \32576 , \32569 );
nand \U$32201 ( \32578 , \32575 , \32577 );
xor \U$32202 ( \32579 , \32532 , \32578 );
not \U$32203 ( \32580 , \30853 );
not \U$32204 ( \32581 , \5049 );
or \U$32205 ( \32582 , \32580 , \32581 );
not \U$32206 ( \32583 , RIae79d90_164);
not \U$32207 ( \32584 , \9412 );
or \U$32208 ( \32585 , \32583 , \32584 );
or \U$32209 ( \32586 , \9412 , RIae79d90_164);
nand \U$32210 ( \32587 , \32585 , \32586 );
not \U$32211 ( \32588 , \32587 );
or \U$32212 ( \32589 , \32588 , \19330 );
nand \U$32213 ( \32590 , \32582 , \32589 );
and \U$32214 ( \32591 , \32579 , \32590 );
and \U$32215 ( \32592 , \32532 , \32578 );
or \U$32216 ( \32593 , \32591 , \32592 );
not \U$32217 ( \32594 , \32593 );
xnor \U$32218 ( \32595 , \30636 , \30617 );
not \U$32219 ( \32596 , \32595 );
not \U$32220 ( \32597 , \32596 );
xor \U$32221 ( \32598 , \30750 , \30740 );
not \U$32222 ( \32599 , \32598 );
not \U$32223 ( \32600 , \32599 );
or \U$32224 ( \32601 , \32597 , \32600 );
nand \U$32225 ( \32602 , \32598 , \32595 );
nand \U$32226 ( \32603 , \32601 , \32602 );
not \U$32227 ( \32604 , \32603 );
or \U$32228 ( \32605 , \32594 , \32604 );
nand \U$32229 ( \32606 , \32598 , \32596 );
nand \U$32230 ( \32607 , \32605 , \32606 );
not \U$32231 ( \32608 , \32607 );
xor \U$32232 ( \32609 , \30607 , \30641 );
xnor \U$32233 ( \32610 , \32609 , \30600 );
not \U$32234 ( \32611 , \32610 );
xor \U$32235 ( \32612 , \30422 , \30432 );
xor \U$32236 ( \32613 , \32612 , \30443 );
not \U$32237 ( \32614 , \32613 );
or \U$32238 ( \32615 , \32611 , \32614 );
or \U$32239 ( \32616 , \32613 , \32610 );
nand \U$32240 ( \32617 , \32615 , \32616 );
not \U$32241 ( \32618 , \32617 );
or \U$32242 ( \32619 , \32608 , \32618 );
not \U$32243 ( \32620 , \32610 );
nand \U$32244 ( \32621 , \32620 , \32613 );
nand \U$32245 ( \32622 , \32619 , \32621 );
not \U$32246 ( \32623 , \32622 );
not \U$32247 ( \32624 , \32623 );
xor \U$32248 ( \32625 , \31110 , \31118 );
xnor \U$32249 ( \32626 , \32625 , \31121 );
not \U$32250 ( \32627 , \32626 );
or \U$32251 ( \32628 , \32624 , \32627 );
or \U$32252 ( \32629 , \32626 , \32623 );
nand \U$32253 ( \32630 , \32628 , \32629 );
not \U$32254 ( \32631 , \32630 );
or \U$32255 ( \32632 , \32522 , \32631 );
nand \U$32256 ( \32633 , \32626 , \32622 );
nand \U$32257 ( \32634 , \32632 , \32633 );
not \U$32258 ( \32635 , \32634 );
or \U$32259 ( \32636 , \32357 , \32635 );
or \U$32260 ( \32637 , \32634 , \32356 );
nand \U$32261 ( \32638 , \32636 , \32637 );
not \U$32262 ( \32639 , \32638 );
or \U$32263 ( \32640 , \32354 , \32639 );
or \U$32264 ( \32641 , \32638 , \32353 );
nand \U$32265 ( \32642 , \32640 , \32641 );
not \U$32266 ( \32643 , \32642 );
xnor \U$32267 ( \32644 , \32350 , \32349 );
not \U$32268 ( \32645 , \32644 );
not \U$32269 ( \32646 , \32645 );
xor \U$32270 ( \32647 , \32516 , \32398 );
not \U$32271 ( \32648 , \32647 );
xor \U$32272 ( \32649 , \32617 , \32607 );
xnor \U$32273 ( \32650 , \32603 , \32593 );
not \U$32274 ( \32651 , \32650 );
not \U$32275 ( \32652 , \32394 );
not \U$32276 ( \32653 , \32388 );
not \U$32277 ( \32654 , \32653 );
and \U$32278 ( \32655 , \32652 , \32654 );
and \U$32279 ( \32656 , \32394 , \32653 );
nor \U$32280 ( \32657 , \32655 , \32656 );
not \U$32281 ( \32658 , \32657 );
or \U$32282 ( \32659 , \32651 , \32658 );
xor \U$32283 ( \32660 , \32450 , \32459 );
xor \U$32284 ( \32661 , \32660 , \32470 );
not \U$32285 ( \32662 , \32661 );
xor \U$32286 ( \32663 , \32416 , \32425 );
xor \U$32287 ( \32664 , \32663 , \32435 );
not \U$32288 ( \32665 , \32664 );
xor \U$32289 ( \32666 , \32532 , \32578 );
xor \U$32290 ( \32667 , \32666 , \32590 );
not \U$32291 ( \32668 , \32667 );
nand \U$32292 ( \32669 , \32665 , \32668 );
not \U$32293 ( \32670 , \32669 );
or \U$32294 ( \32671 , \32662 , \32670 );
nand \U$32295 ( \32672 , \32664 , \32667 );
nand \U$32296 ( \32673 , \32671 , \32672 );
nand \U$32297 ( \32674 , \32659 , \32673 );
not \U$32298 ( \32675 , \32650 );
not \U$32299 ( \32676 , \32657 );
nand \U$32300 ( \32677 , \32675 , \32676 );
nand \U$32301 ( \32678 , \32674 , \32677 );
xor \U$32302 ( \32679 , \32649 , \32678 );
not \U$32303 ( \32680 , \32679 );
or \U$32304 ( \32681 , \32648 , \32680 );
not \U$32305 ( \32682 , \32677 );
not \U$32306 ( \32683 , \32674 );
or \U$32307 ( \32684 , \32682 , \32683 );
nand \U$32308 ( \32685 , \32684 , \32649 );
nand \U$32309 ( \32686 , \32681 , \32685 );
not \U$32310 ( \32687 , \32686 );
or \U$32311 ( \32688 , \32646 , \32687 );
not \U$32312 ( \32689 , \32686 );
not \U$32313 ( \32690 , \32689 );
not \U$32314 ( \32691 , \32644 );
or \U$32315 ( \32692 , \32690 , \32691 );
xor \U$32316 ( \32693 , \31031 , \31063 );
xnor \U$32317 ( \32694 , \32693 , \31073 );
not \U$32318 ( \32695 , \30830 );
nand \U$32319 ( \32696 , \32695 , \30839 );
xor \U$32320 ( \32697 , \32696 , \30836 );
xor \U$32321 ( \32698 , \32694 , \32697 );
not \U$32322 ( \32699 , \19466 );
not \U$32323 ( \32700 , RIae7a240_174);
not \U$32324 ( \32701 , \9299 );
or \U$32325 ( \32702 , \32700 , \32701 );
or \U$32326 ( \32703 , \6231 , RIae7a240_174);
nand \U$32327 ( \32704 , \32702 , \32703 );
not \U$32328 ( \32705 , \32704 );
or \U$32329 ( \32706 , \32699 , \32705 );
nand \U$32330 ( \32707 , \32414 , \9699 );
nand \U$32331 ( \32708 , \32706 , \32707 );
not \U$32332 ( \32709 , \32708 );
not \U$32333 ( \32710 , \9792 );
not \U$32334 ( \32711 , \9804 );
not \U$32335 ( \32712 , \24815 );
or \U$32336 ( \32713 , \32711 , \32712 );
or \U$32337 ( \32714 , \9350 , \9810 );
nand \U$32338 ( \32715 , \32713 , \32714 );
not \U$32339 ( \32716 , \32715 );
or \U$32340 ( \32717 , \32710 , \32716 );
nand \U$32341 ( \32718 , \32493 , \9814 );
nand \U$32342 ( \32719 , \32717 , \32718 );
not \U$32343 ( \32720 , \32719 );
nand \U$32344 ( \32721 , \32709 , \32720 );
not \U$32345 ( \32722 , \32721 );
not \U$32346 ( \32723 , \9622 );
not \U$32347 ( \32724 , \32423 );
or \U$32348 ( \32725 , \32723 , \32724 );
not \U$32349 ( \32726 , \13165 );
not \U$32350 ( \32727 , \5722 );
or \U$32351 ( \32728 , \32726 , \32727 );
nand \U$32352 ( \32729 , \15207 , RIae7a3a8_177);
nand \U$32353 ( \32730 , \32728 , \32729 );
nand \U$32354 ( \32731 , \32730 , \9644 );
nand \U$32355 ( \32732 , \32725 , \32731 );
not \U$32356 ( \32733 , \32732 );
or \U$32357 ( \32734 , \32722 , \32733 );
not \U$32358 ( \32735 , \32720 );
nand \U$32359 ( \32736 , \32735 , \32708 );
nand \U$32360 ( \32737 , \32734 , \32736 );
not \U$32361 ( \32738 , \32737 );
xor \U$32362 ( \32739 , \31037 , \31050 );
xor \U$32363 ( \32740 , \32739 , \31060 );
not \U$32364 ( \32741 , \32740 );
xnor \U$32365 ( \32742 , \31009 , \31019 );
not \U$32366 ( \32743 , \32742 );
not \U$32367 ( \32744 , \2431 );
not \U$32368 ( \32745 , RIae79778_151);
not \U$32369 ( \32746 , \9875 );
or \U$32370 ( \32747 , \32745 , \32746 );
or \U$32371 ( \32748 , \10749 , RIae79778_151);
nand \U$32372 ( \32749 , \32747 , \32748 );
not \U$32373 ( \32750 , \32749 );
or \U$32374 ( \32751 , \32744 , \32750 );
nand \U$32375 ( \32752 , \31048 , \2450 );
nand \U$32376 ( \32753 , \32751 , \32752 );
not \U$32377 ( \32754 , \32753 );
or \U$32378 ( \32755 , \32743 , \32754 );
or \U$32379 ( \32756 , \32753 , \32742 );
nand \U$32380 ( \32757 , \32755 , \32756 );
not \U$32381 ( \32758 , \2417 );
xor \U$32382 ( \32759 , \10070 , RIae79c28_161);
not \U$32383 ( \32760 , \32759 );
or \U$32384 ( \32761 , \32758 , \32760 );
nand \U$32385 ( \32762 , \31058 , \2418 );
nand \U$32386 ( \32763 , \32761 , \32762 );
nand \U$32387 ( \32764 , \32757 , \32763 );
not \U$32388 ( \32765 , \32742 );
nand \U$32389 ( \32766 , \32765 , \32753 );
and \U$32390 ( \32767 , \32764 , \32766 );
not \U$32391 ( \32768 , \32767 );
or \U$32392 ( \32769 , \32741 , \32768 );
not \U$32393 ( \32770 , \32766 );
not \U$32394 ( \32771 , \32764 );
or \U$32395 ( \32772 , \32770 , \32771 );
not \U$32396 ( \32773 , \32740 );
nand \U$32397 ( \32774 , \32772 , \32773 );
nand \U$32398 ( \32775 , \32769 , \32774 );
not \U$32399 ( \32776 , \32775 );
or \U$32400 ( \32777 , \32738 , \32776 );
not \U$32401 ( \32778 , \32767 );
nand \U$32402 ( \32779 , \32778 , \32740 );
nand \U$32403 ( \32780 , \32777 , \32779 );
not \U$32404 ( \32781 , \32780 );
xor \U$32405 ( \32782 , \32698 , \32781 );
not \U$32406 ( \32783 , \32782 );
not \U$32407 ( \32784 , \32783 );
not \U$32408 ( \32785 , \32308 );
not \U$32409 ( \32786 , \32297 );
or \U$32410 ( \32787 , \32785 , \32786 );
or \U$32411 ( \32788 , \32297 , \32308 );
nand \U$32412 ( \32789 , \32787 , \32788 );
not \U$32413 ( \32790 , \32789 );
not \U$32414 ( \32791 , \32320 );
and \U$32415 ( \32792 , \32790 , \32791 );
and \U$32416 ( \32793 , \32789 , \32320 );
nor \U$32417 ( \32794 , \32792 , \32793 );
not \U$32418 ( \32795 , \2776 );
not \U$32419 ( \32796 , \32759 );
or \U$32420 ( \32797 , \32795 , \32796 );
and \U$32421 ( \32798 , RIae79c28_161, \11272 );
not \U$32422 ( \32799 , RIae79c28_161);
and \U$32423 ( \32800 , \32799 , \10168 );
nor \U$32424 ( \32801 , \32798 , \32800 );
nand \U$32425 ( \32802 , \32801 , \2417 );
nand \U$32426 ( \32803 , \32797 , \32802 );
not \U$32427 ( \32804 , \32803 );
not \U$32428 ( \32805 , \1919 );
not \U$32429 ( \32806 , \32567 );
or \U$32430 ( \32807 , \32805 , \32806 );
not \U$32431 ( \32808 , \10272 );
and \U$32432 ( \32809 , \3039 , \32808 );
not \U$32433 ( \32810 , \3039 );
and \U$32434 ( \32811 , \32810 , \10272 );
nor \U$32435 ( \32812 , \32809 , \32811 );
nand \U$32436 ( \32813 , \32812 , \1932 );
nand \U$32437 ( \32814 , \32807 , \32813 );
not \U$32438 ( \32815 , \32814 );
not \U$32439 ( \32816 , \1919 );
not \U$32440 ( \32817 , \32812 );
or \U$32441 ( \32818 , \32816 , \32817 );
and \U$32442 ( \32819 , RIae794a8_145, \10259 );
not \U$32443 ( \32820 , RIae794a8_145);
and \U$32444 ( \32821 , \32820 , \18971 );
or \U$32445 ( \32822 , \32819 , \32821 );
nand \U$32446 ( \32823 , \32822 , \1932 );
nand \U$32447 ( \32824 , \32818 , \32823 );
not \U$32448 ( \32825 , \32824 );
and \U$32449 ( \32826 , \12857 , \2249 );
not \U$32450 ( \32827 , \32826 );
not \U$32451 ( \32828 , \2161 );
xor \U$32452 ( \32829 , \2183 , \16651 );
not \U$32453 ( \32830 , \32829 );
or \U$32454 ( \32831 , \32828 , \32830 );
not \U$32455 ( \32832 , RIae79520_146);
not \U$32456 ( \32833 , \12750 );
or \U$32457 ( \32834 , \32832 , \32833 );
or \U$32458 ( \32835 , \16006 , RIae79520_146);
nand \U$32459 ( \32836 , \32834 , \32835 );
nand \U$32460 ( \32837 , \32836 , \2188 );
nand \U$32461 ( \32838 , \32831 , \32837 );
not \U$32462 ( \32839 , \32838 );
not \U$32463 ( \32840 , \32839 );
or \U$32464 ( \32841 , \32827 , \32840 );
or \U$32465 ( \32842 , \32839 , \32826 );
nand \U$32466 ( \32843 , \32841 , \32842 );
not \U$32467 ( \32844 , \32843 );
or \U$32468 ( \32845 , \32825 , \32844 );
nand \U$32469 ( \32846 , \32838 , \32826 );
nand \U$32470 ( \32847 , \32845 , \32846 );
not \U$32471 ( \32848 , \32847 );
not \U$32472 ( \32849 , \32848 );
or \U$32473 ( \32850 , \32815 , \32849 );
not \U$32474 ( \32851 , \32814 );
nand \U$32475 ( \32852 , \32851 , \32847 );
nand \U$32476 ( \32853 , \32850 , \32852 );
not \U$32477 ( \32854 , \32853 );
or \U$32478 ( \32855 , \32804 , \32854 );
nand \U$32479 ( \32856 , \32847 , \32814 );
nand \U$32480 ( \32857 , \32855 , \32856 );
not \U$32481 ( \32858 , \4853 );
and \U$32482 ( \32859 , RIae79ca0_162, \12644 );
not \U$32483 ( \32860 , RIae79ca0_162);
and \U$32484 ( \32861 , \32860 , \16826 );
nor \U$32485 ( \32862 , \32859 , \32861 );
not \U$32486 ( \32863 , \32862 );
or \U$32487 ( \32864 , \32858 , \32863 );
and \U$32488 ( \32865 , \10208 , RIae79ca0_162);
not \U$32489 ( \32866 , \10208 );
and \U$32490 ( \32867 , \32866 , \11755 );
nor \U$32491 ( \32868 , \32865 , \32867 );
nand \U$32492 ( \32869 , \32868 , \4154 );
nand \U$32493 ( \32870 , \32864 , \32869 );
not \U$32494 ( \32871 , \32870 );
not \U$32495 ( \32872 , \2007 );
and \U$32496 ( \32873 , RIae797f0_152, \17423 );
not \U$32497 ( \32874 , RIae797f0_152);
and \U$32498 ( \32875 , \32874 , \16193 );
nor \U$32499 ( \32876 , \32873 , \32875 );
not \U$32500 ( \32877 , \32876 );
or \U$32501 ( \32878 , \32872 , \32877 );
and \U$32502 ( \32879 , \10149 , \2521 );
not \U$32503 ( \32880 , \10149 );
and \U$32504 ( \32881 , \32880 , RIae797f0_152);
nor \U$32505 ( \32882 , \32879 , \32881 );
nand \U$32506 ( \32883 , \32882 , \1988 );
nand \U$32507 ( \32884 , \32878 , \32883 );
not \U$32508 ( \32885 , \32884 );
not \U$32509 ( \32886 , \32885 );
not \U$32510 ( \32887 , \15337 );
not \U$32511 ( \32888 , \32749 );
or \U$32512 ( \32889 , \32887 , \32888 );
not \U$32513 ( \32890 , \2447 );
not \U$32514 ( \32891 , \10007 );
or \U$32515 ( \32892 , \32890 , \32891 );
or \U$32516 ( \32893 , \10007 , \2504 );
nand \U$32517 ( \32894 , \32892 , \32893 );
nand \U$32518 ( \32895 , \32894 , \2432 );
nand \U$32519 ( \32896 , \32889 , \32895 );
not \U$32520 ( \32897 , \32896 );
or \U$32521 ( \32898 , \32886 , \32897 );
or \U$32522 ( \32899 , \32896 , \32885 );
nand \U$32523 ( \32900 , \32898 , \32899 );
not \U$32524 ( \32901 , \32900 );
or \U$32525 ( \32902 , \32871 , \32901 );
nand \U$32526 ( \32903 , \32896 , \32884 );
nand \U$32527 ( \32904 , \32902 , \32903 );
xor \U$32528 ( \32905 , \32857 , \32904 );
not \U$32529 ( \32906 , \32905 );
not \U$32530 ( \32907 , \11434 );
and \U$32531 ( \32908 , \4169 , RIae7a498_179);
not \U$32532 ( \32909 , \4169 );
and \U$32533 ( \32910 , \32909 , \27628 );
nor \U$32534 ( \32911 , \32908 , \32910 );
not \U$32535 ( \32912 , \32911 );
or \U$32536 ( \32913 , \32907 , \32912 );
xor \U$32537 ( \32914 , RIae7a498_179, \3207 );
nand \U$32538 ( \32915 , \32914 , \12371 );
nand \U$32539 ( \32916 , \32913 , \32915 );
not \U$32540 ( \32917 , \32916 );
not \U$32541 ( \32918 , \2321 );
not \U$32542 ( \32919 , \32538 );
or \U$32543 ( \32920 , \32918 , \32919 );
not \U$32544 ( \32921 , \10043 );
not \U$32545 ( \32922 , \2334 );
or \U$32546 ( \32923 , \32921 , \32922 );
or \U$32547 ( \32924 , \16912 , \2334 );
nand \U$32548 ( \32925 , \32923 , \32924 );
nand \U$32549 ( \32926 , \32925 , \2339 );
nand \U$32550 ( \32927 , \32920 , \32926 );
not \U$32551 ( \32928 , \32557 );
not \U$32552 ( \32929 , \32546 );
and \U$32553 ( \32930 , \32928 , \32929 );
and \U$32554 ( \32931 , \32557 , \32546 );
nor \U$32555 ( \32932 , \32930 , \32931 );
not \U$32556 ( \32933 , \32932 );
not \U$32557 ( \32934 , \2162 );
not \U$32558 ( \32935 , \31017 );
or \U$32559 ( \32936 , \32934 , \32935 );
nand \U$32560 ( \32937 , \32829 , \2188 );
nand \U$32561 ( \32938 , \32936 , \32937 );
not \U$32562 ( \32939 , \32938 );
or \U$32563 ( \32940 , \32933 , \32939 );
or \U$32564 ( \32941 , \32938 , \32932 );
nand \U$32565 ( \32942 , \32940 , \32941 );
not \U$32566 ( \32943 , \32942 );
and \U$32567 ( \32944 , \32927 , \32943 );
not \U$32568 ( \32945 , \32927 );
and \U$32569 ( \32946 , \32945 , \32942 );
nor \U$32570 ( \32947 , \32944 , \32946 );
not \U$32571 ( \32948 , \32947 );
not \U$32572 ( \32949 , \9814 );
not \U$32573 ( \32950 , \32715 );
or \U$32574 ( \32951 , \32949 , \32950 );
xor \U$32575 ( \32952 , RIae7a2b8_175, \32481 );
nand \U$32576 ( \32953 , \32952 , \9792 );
nand \U$32577 ( \32954 , \32951 , \32953 );
not \U$32578 ( \32955 , \32954 );
or \U$32579 ( \32956 , \32948 , \32955 );
or \U$32580 ( \32957 , \32954 , \32947 );
nand \U$32581 ( \32958 , \32956 , \32957 );
not \U$32582 ( \32959 , \32958 );
or \U$32583 ( \32960 , \32917 , \32959 );
not \U$32584 ( \32961 , \32947 );
nand \U$32585 ( \32962 , \32961 , \32954 );
nand \U$32586 ( \32963 , \32960 , \32962 );
not \U$32587 ( \32964 , \32963 );
or \U$32588 ( \32965 , \32906 , \32964 );
nand \U$32589 ( \32966 , \32904 , \32857 );
nand \U$32590 ( \32967 , \32965 , \32966 );
xor \U$32591 ( \32968 , \32794 , \32967 );
xor \U$32592 ( \32969 , \32363 , \32384 );
and \U$32593 ( \32970 , \32968 , \32969 );
and \U$32594 ( \32971 , \32794 , \32967 );
or \U$32595 ( \32972 , \32970 , \32971 );
not \U$32596 ( \32973 , \32330 );
not \U$32597 ( \32974 , \32290 );
not \U$32598 ( \32975 , \32974 );
and \U$32599 ( \32976 , \32973 , \32975 );
and \U$32600 ( \32977 , \32330 , \32974 );
nor \U$32601 ( \32978 , \32976 , \32977 );
xnor \U$32602 ( \32979 , \32972 , \32978 );
not \U$32603 ( \32980 , \32979 );
or \U$32604 ( \32981 , \32784 , \32980 );
not \U$32605 ( \32982 , \32978 );
nand \U$32606 ( \32983 , \32982 , \32972 );
nand \U$32607 ( \32984 , \32981 , \32983 );
xor \U$32608 ( \32985 , \32334 , \32343 );
xor \U$32609 ( \32986 , \32985 , \32345 );
nor \U$32610 ( \32987 , \32984 , \32986 );
not \U$32611 ( \32988 , \30974 );
and \U$32612 ( \32989 , \31077 , \32988 );
not \U$32613 ( \32990 , \31077 );
and \U$32614 ( \32991 , \32990 , \30974 );
nor \U$32615 ( \32992 , \32989 , \32991 );
xor \U$32616 ( \32993 , \32694 , \32697 );
and \U$32617 ( \32994 , \32993 , \32781 );
and \U$32618 ( \32995 , \32694 , \32697 );
or \U$32619 ( \32996 , \32994 , \32995 );
nand \U$32620 ( \32997 , \32992 , \32996 );
not \U$32621 ( \32998 , \32992 );
not \U$32622 ( \32999 , \32996 );
nand \U$32623 ( \33000 , \32998 , \32999 );
nand \U$32624 ( \33001 , \32997 , \33000 );
not \U$32625 ( \33002 , \9473 );
not \U$32626 ( \33003 , RIae7a6f0_184);
not \U$32627 ( \33004 , \2697 );
or \U$32628 ( \33005 , \33003 , \33004 );
or \U$32629 ( \33006 , \2697 , RIae7a6f0_184);
nand \U$32630 ( \33007 , \33005 , \33006 );
not \U$32631 ( \33008 , \33007 );
or \U$32632 ( \33009 , \33002 , \33008 );
nand \U$32633 ( \33010 , \32318 , \9705 );
nand \U$32634 ( \33011 , \33009 , \33010 );
not \U$32635 ( \33012 , \33011 );
not \U$32636 ( \33013 , RIae7a150_172);
not \U$32637 ( \33014 , \1860 );
or \U$32638 ( \33015 , \33013 , \33014 );
or \U$32639 ( \33016 , \1859 , RIae7a150_172);
nand \U$32640 ( \33017 , \33015 , \33016 );
and \U$32641 ( \33018 , \33017 , \13158 );
not \U$32642 ( \33019 , \9776 );
nor \U$32643 ( \33020 , \33019 , \32371 );
nor \U$32644 ( \33021 , \33018 , \33020 );
not \U$32645 ( \33022 , \33021 );
not \U$32646 ( \33023 , RIae7aab0_192);
not \U$32647 ( \33024 , \32468 );
or \U$32648 ( \33025 , \33023 , \33024 );
and \U$32649 ( \33026 , \2309 , RIae7aa38_191);
not \U$32650 ( \33027 , \2309 );
and \U$32651 ( \33028 , \33027 , \11326 );
nor \U$32652 ( \33029 , \33026 , \33028 );
nand \U$32653 ( \33030 , \33029 , \16383 );
nand \U$32654 ( \33031 , \33025 , \33030 );
not \U$32655 ( \33032 , \33031 );
or \U$32656 ( \33033 , \33022 , \33032 );
or \U$32657 ( \33034 , \33031 , \33021 );
nand \U$32658 ( \33035 , \33033 , \33034 );
not \U$32659 ( \33036 , \33035 );
or \U$32660 ( \33037 , \33012 , \33036 );
not \U$32661 ( \33038 , \33021 );
nand \U$32662 ( \33039 , \33038 , \33031 );
nand \U$32663 ( \33040 , \33037 , \33039 );
not \U$32664 ( \33041 , \33040 );
not \U$32665 ( \33042 , \9518 );
not \U$32666 ( \33043 , \32483 );
or \U$32667 ( \33044 , \33042 , \33043 );
xor \U$32668 ( \33045 , RIae79fe8_169, \9438 );
nand \U$32669 ( \33046 , \33045 , \9499 );
nand \U$32670 ( \33047 , \33044 , \33046 );
not \U$32671 ( \33048 , \33047 );
not \U$32672 ( \33049 , \33048 );
not \U$32673 ( \33050 , \4968 );
not \U$32674 ( \33051 , \9609 );
or \U$32675 ( \33052 , \33050 , \33051 );
or \U$32676 ( \33053 , \9609 , \4968 );
nand \U$32677 ( \33054 , \33052 , \33053 );
not \U$32678 ( \33055 , \33054 );
not \U$32679 ( \33056 , \5039 );
or \U$32680 ( \33057 , \33055 , \33056 );
nand \U$32681 ( \33058 , \32587 , \5049 );
nand \U$32682 ( \33059 , \33057 , \33058 );
not \U$32683 ( \33060 , \33059 );
or \U$32684 ( \33061 , \33049 , \33060 );
or \U$32685 ( \33062 , \33048 , \33059 );
nand \U$32686 ( \33063 , \33061 , \33062 );
not \U$32687 ( \33064 , \33063 );
not \U$32688 ( \33065 , \10519 );
not \U$32689 ( \33066 , \32455 );
or \U$32690 ( \33067 , \33065 , \33066 );
not \U$32691 ( \33068 , RIae7a7e0_186);
not \U$32692 ( \33069 , \3417 );
or \U$32693 ( \33070 , \33068 , \33069 );
or \U$32694 ( \33071 , \13942 , RIae7a7e0_186);
nand \U$32695 ( \33072 , \33070 , \33071 );
nand \U$32696 ( \33073 , \33072 , \11851 );
nand \U$32697 ( \33074 , \33067 , \33073 );
not \U$32698 ( \33075 , \33074 );
or \U$32699 ( \33076 , \33064 , \33075 );
nand \U$32700 ( \33077 , \33047 , \33059 );
nand \U$32701 ( \33078 , \33076 , \33077 );
not \U$32702 ( \33079 , \32485 );
not \U$32703 ( \33080 , \33079 );
not \U$32704 ( \33081 , \32502 );
or \U$32705 ( \33082 , \33080 , \33081 );
or \U$32706 ( \33083 , \32502 , \33079 );
nand \U$32707 ( \33084 , \33082 , \33083 );
xor \U$32708 ( \33085 , \33078 , \33084 );
not \U$32709 ( \33086 , \33085 );
or \U$32710 ( \33087 , \33041 , \33086 );
nand \U$32711 ( \33088 , \33078 , \33084 );
nand \U$32712 ( \33089 , \33087 , \33088 );
not \U$32713 ( \33090 , \33089 );
and \U$32714 ( \33091 , \32507 , \32439 );
not \U$32715 ( \33092 , \32507 );
and \U$32716 ( \33093 , \33092 , \32438 );
nor \U$32717 ( \33094 , \33091 , \33093 );
xor \U$32718 ( \33095 , \33094 , \32473 );
nand \U$32719 ( \33096 , \33090 , \33095 );
not \U$32720 ( \33097 , \33096 );
not \U$32721 ( \33098 , \17847 );
and \U$32722 ( \33099 , \6642 , RIae7a8d0_188);
not \U$32723 ( \33100 , \6642 );
and \U$32724 ( \33101 , \33100 , \18088 );
nor \U$32725 ( \33102 , \33099 , \33101 );
not \U$32726 ( \33103 , \33102 );
or \U$32727 ( \33104 , \33098 , \33103 );
nand \U$32728 ( \33105 , \32359 , \10275 );
nand \U$32729 ( \33106 , \33104 , \33105 );
not \U$32730 ( \33107 , \33106 );
not \U$32731 ( \33108 , \32542 );
not \U$32732 ( \33109 , \33108 );
not \U$32733 ( \33110 , \32573 );
or \U$32734 ( \33111 , \33109 , \33110 );
or \U$32735 ( \33112 , \32573 , \33108 );
nand \U$32736 ( \33113 , \33111 , \33112 );
not \U$32737 ( \33114 , \33113 );
not \U$32738 ( \33115 , \9729 );
xor \U$32739 ( \33116 , RIae7a060_170, \5911 );
not \U$32740 ( \33117 , \33116 );
or \U$32741 ( \33118 , \33115 , \33117 );
nand \U$32742 ( \33119 , \32381 , \11098 );
nand \U$32743 ( \33120 , \33118 , \33119 );
not \U$32744 ( \33121 , \33120 );
not \U$32745 ( \33122 , \33121 );
or \U$32746 ( \33123 , \33114 , \33122 );
not \U$32747 ( \33124 , \33113 );
nand \U$32748 ( \33125 , \33124 , \33120 );
nand \U$32749 ( \33126 , \33123 , \33125 );
not \U$32750 ( \33127 , \33126 );
or \U$32751 ( \33128 , \33107 , \33127 );
nand \U$32752 ( \33129 , \33120 , \33113 );
nand \U$32753 ( \33130 , \33128 , \33129 );
not \U$32754 ( \33131 , \33130 );
not \U$32755 ( \33132 , \32942 );
not \U$32756 ( \33133 , \32927 );
or \U$32757 ( \33134 , \33132 , \33133 );
not \U$32758 ( \33135 , \32932 );
nand \U$32759 ( \33136 , \33135 , \32938 );
nand \U$32760 ( \33137 , \33134 , \33136 );
not \U$32761 ( \33138 , \33137 );
not \U$32762 ( \33139 , \33138 );
not \U$32763 ( \33140 , \19362 );
xor \U$32764 ( \33141 , RIae79ef8_167, \9395 );
not \U$32765 ( \33142 , \33141 );
or \U$32766 ( \33143 , \33140 , \33142 );
nand \U$32767 ( \33144 , \32530 , \6212 );
nand \U$32768 ( \33145 , \33143 , \33144 );
not \U$32769 ( \33146 , \33145 );
or \U$32770 ( \33147 , \33139 , \33146 );
or \U$32771 ( \33148 , \33145 , \33138 );
nand \U$32772 ( \33149 , \33147 , \33148 );
not \U$32773 ( \33150 , \33149 );
not \U$32774 ( \33151 , \16564 );
not \U$32775 ( \33152 , \32914 );
or \U$32776 ( \33153 , \33151 , \33152 );
nand \U$32777 ( \33154 , \32305 , \11422 );
nand \U$32778 ( \33155 , \33153 , \33154 );
not \U$32779 ( \33156 , \33155 );
or \U$32780 ( \33157 , \33150 , \33156 );
not \U$32781 ( \33158 , \33138 );
nand \U$32782 ( \33159 , \33158 , \33145 );
nand \U$32783 ( \33160 , \33157 , \33159 );
not \U$32784 ( \33161 , \33160 );
nand \U$32785 ( \33162 , \32430 , \10631 );
not \U$32786 ( \33163 , \33162 );
not \U$32787 ( \33164 , RIae7a510_180);
not \U$32788 ( \33165 , \10829 );
or \U$32789 ( \33166 , \33164 , \33165 );
or \U$32790 ( \33167 , \10226 , RIae7a510_180);
nand \U$32791 ( \33168 , \33166 , \33167 );
nand \U$32792 ( \33169 , \33168 , \10637 );
not \U$32793 ( \33170 , \33169 );
or \U$32794 ( \33171 , \33163 , \33170 );
not \U$32795 ( \33172 , \2007 );
not \U$32796 ( \33173 , \30982 );
or \U$32797 ( \33174 , \33172 , \33173 );
nand \U$32798 ( \33175 , \32876 , \1988 );
nand \U$32799 ( \33176 , \33174 , \33175 );
not \U$32800 ( \33177 , \33176 );
not \U$32801 ( \33178 , \4154 );
not \U$32802 ( \33179 , \32862 );
or \U$32803 ( \33180 , \33178 , \33179 );
nand \U$32804 ( \33181 , \32448 , \4853 );
nand \U$32805 ( \33182 , \33180 , \33181 );
not \U$32806 ( \33183 , \33182 );
not \U$32807 ( \33184 , \33183 );
or \U$32808 ( \33185 , \33177 , \33184 );
not \U$32809 ( \33186 , \33176 );
nand \U$32810 ( \33187 , \33186 , \33182 );
nand \U$32811 ( \33188 , \33185 , \33187 );
nand \U$32812 ( \33189 , \33171 , \33188 );
nand \U$32813 ( \33190 , \33182 , \33176 );
and \U$32814 ( \33191 , \33189 , \33190 );
not \U$32815 ( \33192 , \33191 );
or \U$32816 ( \33193 , \33161 , \33192 );
not \U$32817 ( \33194 , \33190 );
not \U$32818 ( \33195 , \33189 );
or \U$32819 ( \33196 , \33194 , \33195 );
not \U$32820 ( \33197 , \33160 );
nand \U$32821 ( \33198 , \33196 , \33197 );
nand \U$32822 ( \33199 , \33193 , \33198 );
not \U$32823 ( \33200 , \33199 );
or \U$32824 ( \33201 , \33131 , \33200 );
not \U$32825 ( \33202 , \33190 );
not \U$32826 ( \33203 , \33189 );
or \U$32827 ( \33204 , \33202 , \33203 );
nand \U$32828 ( \33205 , \33204 , \33160 );
nand \U$32829 ( \33206 , \33201 , \33205 );
not \U$32830 ( \33207 , \33206 );
or \U$32831 ( \33208 , \33097 , \33207 );
not \U$32832 ( \33209 , \33095 );
nand \U$32833 ( \33210 , \33209 , \33089 );
nand \U$32834 ( \33211 , \33208 , \33210 );
buf \U$32835 ( \33212 , \33211 );
xor \U$32836 ( \33213 , \33001 , \33212 );
or \U$32837 ( \33214 , \32987 , \33213 );
nand \U$32838 ( \33215 , \32984 , \32986 );
nand \U$32839 ( \33216 , \33214 , \33215 );
nand \U$32840 ( \33217 , \32692 , \33216 );
nand \U$32841 ( \33218 , \32688 , \33217 );
not \U$32842 ( \33219 , \33218 );
not \U$32843 ( \33220 , \33219 );
or \U$32844 ( \33221 , \32643 , \33220 );
or \U$32845 ( \33222 , \33219 , \32642 );
nand \U$32846 ( \33223 , \33221 , \33222 );
not \U$32847 ( \33224 , \33223 );
buf \U$32848 ( \33225 , \30595 );
xnor \U$32849 ( \33226 , \30811 , \33225 );
not \U$32850 ( \33227 , \33226 );
not \U$32851 ( \33228 , \30936 );
not \U$32852 ( \33229 , \30962 );
or \U$32853 ( \33230 , \33228 , \33229 );
or \U$32854 ( \33231 , \30962 , \30936 );
nand \U$32855 ( \33232 , \33230 , \33231 );
and \U$32856 ( \33233 , \33232 , \31086 );
not \U$32857 ( \33234 , \33232 );
not \U$32858 ( \33235 , \31086 );
and \U$32859 ( \33236 , \33234 , \33235 );
nor \U$32860 ( \33237 , \33233 , \33236 );
not \U$32861 ( \33238 , \33237 );
or \U$32862 ( \33239 , \33227 , \33238 );
or \U$32863 ( \33240 , \33237 , \33226 );
nand \U$32864 ( \33241 , \33239 , \33240 );
buf \U$32865 ( \33242 , \33241 );
xor \U$32866 ( \33243 , \32521 , \32630 );
not \U$32867 ( \33244 , \33243 );
xor \U$32868 ( \33245 , \30968 , \30970 );
xor \U$32869 ( \33246 , \33245 , \31083 );
not \U$32870 ( \33247 , \32997 );
not \U$32871 ( \33248 , \33211 );
or \U$32872 ( \33249 , \33247 , \33248 );
nand \U$32873 ( \33250 , \33249 , \33000 );
xor \U$32874 ( \33251 , \33246 , \33250 );
not \U$32875 ( \33252 , \33251 );
or \U$32876 ( \33253 , \33244 , \33252 );
nand \U$32877 ( \33254 , \33246 , \33250 );
nand \U$32878 ( \33255 , \33253 , \33254 );
not \U$32879 ( \33256 , \33255 );
and \U$32880 ( \33257 , \33242 , \33256 );
not \U$32881 ( \33258 , \33242 );
and \U$32882 ( \33259 , \33258 , \33255 );
nor \U$32883 ( \33260 , \33257 , \33259 );
not \U$32884 ( \33261 , \33260 );
and \U$32885 ( \33262 , \33224 , \33261 );
and \U$32886 ( \33263 , \33223 , \33260 );
nor \U$32887 ( \33264 , \33262 , \33263 );
xor \U$32888 ( \33265 , \33251 , \33243 );
and \U$32889 ( \33266 , \32979 , \32783 );
not \U$32890 ( \33267 , \32979 );
and \U$32891 ( \33268 , \33267 , \32782 );
nor \U$32892 ( \33269 , \33266 , \33268 );
not \U$32893 ( \33270 , \32673 );
not \U$32894 ( \33271 , \32650 );
and \U$32895 ( \33272 , \33270 , \33271 );
and \U$32896 ( \33273 , \32673 , \32650 );
nor \U$32897 ( \33274 , \33272 , \33273 );
not \U$32898 ( \33275 , \32676 );
and \U$32899 ( \33276 , \33274 , \33275 );
not \U$32900 ( \33277 , \33274 );
and \U$32901 ( \33278 , \33277 , \32676 );
nor \U$32902 ( \33279 , \33276 , \33278 );
or \U$32903 ( \33280 , \33269 , \33279 );
xor \U$32904 ( \33281 , \32794 , \32967 );
xor \U$32905 ( \33282 , \33281 , \32969 );
not \U$32906 ( \33283 , \33282 );
nand \U$32907 ( \33284 , \32669 , \32672 );
not \U$32908 ( \33285 , \32661 );
and \U$32909 ( \33286 , \33284 , \33285 );
not \U$32910 ( \33287 , \33284 );
and \U$32911 ( \33288 , \33287 , \32661 );
nor \U$32912 ( \33289 , \33286 , \33288 );
buf \U$32913 ( \33290 , \33085 );
and \U$32914 ( \33291 , \33290 , \33040 );
not \U$32915 ( \33292 , \33290 );
not \U$32916 ( \33293 , \33040 );
and \U$32917 ( \33294 , \33292 , \33293 );
nor \U$32918 ( \33295 , \33291 , \33294 );
xor \U$32919 ( \33296 , \33289 , \33295 );
not \U$32920 ( \33297 , \33296 );
or \U$32921 ( \33298 , \33283 , \33297 );
nand \U$32922 ( \33299 , \33289 , \33295 );
nand \U$32923 ( \33300 , \33298 , \33299 );
nand \U$32924 ( \33301 , \33280 , \33300 );
nand \U$32925 ( \33302 , \33269 , \33279 );
nand \U$32926 ( \33303 , \33301 , \33302 );
xor \U$32927 ( \33304 , \32647 , \32679 );
or \U$32928 ( \33305 , \33303 , \33304 );
xor \U$32929 ( \33306 , \33089 , \33206 );
xor \U$32930 ( \33307 , \33306 , \33209 );
not \U$32931 ( \33308 , \33307 );
not \U$32932 ( \33309 , \9699 );
not \U$32933 ( \33310 , \32704 );
or \U$32934 ( \33311 , \33309 , \33310 );
and \U$32935 ( \33312 , RIae7a240_174, \15102 );
not \U$32936 ( \33313 , RIae7a240_174);
and \U$32937 ( \33314 , \33313 , \9313 );
nor \U$32938 ( \33315 , \33312 , \33314 );
nand \U$32939 ( \33316 , \33315 , \9688 );
nand \U$32940 ( \33317 , \33311 , \33316 );
not \U$32941 ( \33318 , \11014 );
and \U$32942 ( \33319 , RIae7a3a8_177, \14630 );
not \U$32943 ( \33320 , RIae7a3a8_177);
and \U$32944 ( \33321 , \33320 , \9290 );
or \U$32945 ( \33322 , \33319 , \33321 );
not \U$32946 ( \33323 , \33322 );
or \U$32947 ( \33324 , \33318 , \33323 );
nand \U$32948 ( \33325 , \32730 , \9622 );
nand \U$32949 ( \33326 , \33324 , \33325 );
xor \U$32950 ( \33327 , \33317 , \33326 );
not \U$32951 ( \33328 , \33168 );
or \U$32952 ( \33329 , \33328 , \12232 );
not \U$32953 ( \33330 , RIae7a510_180);
not \U$32954 ( \33331 , \27827 );
or \U$32955 ( \33332 , \33330 , \33331 );
or \U$32956 ( \33333 , \6257 , RIae7a510_180);
nand \U$32957 ( \33334 , \33332 , \33333 );
not \U$32958 ( \33335 , \33334 );
not \U$32959 ( \33336 , \10638 );
or \U$32960 ( \33337 , \33335 , \33336 );
nand \U$32961 ( \33338 , \33329 , \33337 );
and \U$32962 ( \33339 , \33327 , \33338 );
and \U$32963 ( \33340 , \33317 , \33326 );
or \U$32964 ( \33341 , \33339 , \33340 );
not \U$32965 ( \33342 , \33341 );
xnor \U$32966 ( \33343 , \32757 , \32763 );
not \U$32967 ( \33344 , \33343 );
nand \U$32968 ( \33345 , \33169 , \33162 );
xor \U$32969 ( \33346 , \33188 , \33345 );
not \U$32970 ( \33347 , \33346 );
or \U$32971 ( \33348 , \33344 , \33347 );
or \U$32972 ( \33349 , \33346 , \33343 );
nand \U$32973 ( \33350 , \33348 , \33349 );
not \U$32974 ( \33351 , \33350 );
or \U$32975 ( \33352 , \33342 , \33351 );
not \U$32976 ( \33353 , \33343 );
buf \U$32977 ( \33354 , \33346 );
nand \U$32978 ( \33355 , \33353 , \33354 );
nand \U$32979 ( \33356 , \33352 , \33355 );
not \U$32980 ( \33357 , \33356 );
not \U$32981 ( \33358 , \33130 );
not \U$32982 ( \33359 , \33358 );
not \U$32983 ( \33360 , \33199 );
or \U$32984 ( \33361 , \33359 , \33360 );
or \U$32985 ( \33362 , \33199 , \33358 );
nand \U$32986 ( \33363 , \33361 , \33362 );
not \U$32987 ( \33364 , \33363 );
not \U$32988 ( \33365 , \33364 );
or \U$32989 ( \33366 , \33357 , \33365 );
not \U$32990 ( \33367 , \33356 );
nand \U$32991 ( \33368 , \33367 , \33363 );
nand \U$32992 ( \33369 , \33366 , \33368 );
not \U$32993 ( \33370 , \14668 );
xor \U$32994 ( \33371 , \3748 , RIae7aa38_191);
not \U$32995 ( \33372 , \33371 );
or \U$32996 ( \33373 , \33370 , \33372 );
nand \U$32997 ( \33374 , \33029 , RIae7aab0_192);
nand \U$32998 ( \33375 , \33373 , \33374 );
not \U$32999 ( \33376 , \33375 );
not \U$33000 ( \33377 , \9777 );
not \U$33001 ( \33378 , \33017 );
or \U$33002 ( \33379 , \33377 , \33378 );
not \U$33003 ( \33380 , RIae7a150_172);
not \U$33004 ( \33381 , \2402 );
or \U$33005 ( \33382 , \33380 , \33381 );
or \U$33006 ( \33383 , \5674 , RIae7a150_172);
nand \U$33007 ( \33384 , \33382 , \33383 );
nand \U$33008 ( \33385 , \33384 , \9758 );
nand \U$33009 ( \33386 , \33379 , \33385 );
not \U$33010 ( \33387 , \9745 );
not \U$33011 ( \33388 , \33116 );
or \U$33012 ( \33389 , \33387 , \33388 );
not \U$33013 ( \33390 , \9749 );
not \U$33014 ( \33391 , \1973 );
or \U$33015 ( \33392 , \33390 , \33391 );
nand \U$33016 ( \33393 , \1970 , RIae7a060_170);
nand \U$33017 ( \33394 , \33392 , \33393 );
nand \U$33018 ( \33395 , \33394 , \9730 );
nand \U$33019 ( \33396 , \33389 , \33395 );
xor \U$33020 ( \33397 , \33386 , \33396 );
not \U$33021 ( \33398 , \33397 );
or \U$33022 ( \33399 , \33376 , \33398 );
nand \U$33023 ( \33400 , \33396 , \33386 );
nand \U$33024 ( \33401 , \33399 , \33400 );
not \U$33025 ( \33402 , \33401 );
buf \U$33026 ( \33403 , \33149 );
not \U$33027 ( \33404 , \33403 );
and \U$33028 ( \33405 , \33155 , \33404 );
not \U$33029 ( \33406 , \33155 );
and \U$33030 ( \33407 , \33406 , \33403 );
nor \U$33031 ( \33408 , \33405 , \33407 );
not \U$33032 ( \33409 , \33408 );
not \U$33033 ( \33410 , \33409 );
not \U$33034 ( \33411 , \1988 );
and \U$33035 ( \33412 , RIae797f0_152, \16922 );
not \U$33036 ( \33413 , RIae797f0_152);
not \U$33037 ( \33414 , \10031 );
not \U$33038 ( \33415 , \33414 );
and \U$33039 ( \33416 , \33413 , \33415 );
or \U$33040 ( \33417 , \33412 , \33416 );
not \U$33041 ( \33418 , \33417 );
or \U$33042 ( \33419 , \33411 , \33418 );
not \U$33043 ( \33420 , \32882 );
or \U$33044 ( \33421 , \33420 , \2518 );
nand \U$33045 ( \33422 , \33419 , \33421 );
not \U$33046 ( \33423 , \33422 );
not \U$33047 ( \33424 , \2322 );
not \U$33048 ( \33425 , \32925 );
or \U$33049 ( \33426 , \33424 , \33425 );
and \U$33050 ( \33427 , RIae798e0_154, \10195 );
not \U$33051 ( \33428 , RIae798e0_154);
and \U$33052 ( \33429 , \33428 , \11240 );
nor \U$33053 ( \33430 , \33427 , \33429 );
nand \U$33054 ( \33431 , \33430 , \2339 );
nand \U$33055 ( \33432 , \33426 , \33431 );
not \U$33056 ( \33433 , \33432 );
or \U$33057 ( \33434 , \3039 , \2184 );
or \U$33058 ( \33435 , RIae79430_144, RIae794a8_145);
nand \U$33059 ( \33436 , \33435 , \12857 );
nand \U$33060 ( \33437 , \33434 , \33436 , RIae79520_146);
not \U$33061 ( \33438 , \33437 );
not \U$33062 ( \33439 , \2188 );
or \U$33063 ( \33440 , \12857 , \4653 );
or \U$33064 ( \33441 , \17971 , RIae79520_146);
nand \U$33065 ( \33442 , \33440 , \33441 );
not \U$33066 ( \33443 , \33442 );
or \U$33067 ( \33444 , \33439 , \33443 );
nand \U$33068 ( \33445 , \32836 , \2161 );
nand \U$33069 ( \33446 , \33444 , \33445 );
nand \U$33070 ( \33447 , \33438 , \33446 );
not \U$33071 ( \33448 , \33447 );
and \U$33072 ( \33449 , \33433 , \33448 );
and \U$33073 ( \33450 , \33432 , \33447 );
nor \U$33074 ( \33451 , \33449 , \33450 );
not \U$33075 ( \33452 , \33451 );
not \U$33076 ( \33453 , \33452 );
or \U$33077 ( \33454 , \33423 , \33453 );
not \U$33078 ( \33455 , \33447 );
nand \U$33079 ( \33456 , \33455 , \33432 );
nand \U$33080 ( \33457 , \33454 , \33456 );
not \U$33081 ( \33458 , \33457 );
not \U$33082 ( \33459 , \6214 );
not \U$33083 ( \33460 , \33141 );
or \U$33084 ( \33461 , \33459 , \33460 );
not \U$33085 ( \33462 , RIae79ef8_167);
not \U$33086 ( \33463 , \9412 );
or \U$33087 ( \33464 , \33462 , \33463 );
or \U$33088 ( \33465 , \9417 , RIae79ef8_167);
nand \U$33089 ( \33466 , \33464 , \33465 );
nand \U$33090 ( \33467 , \33466 , \14768 );
nand \U$33091 ( \33468 , \33461 , \33467 );
not \U$33092 ( \33469 , \9517 );
not \U$33093 ( \33470 , \33045 );
or \U$33094 ( \33471 , \33469 , \33470 );
not \U$33095 ( \33472 , \18027 );
not \U$33096 ( \33473 , \9455 );
or \U$33097 ( \33474 , \33472 , \33473 );
or \U$33098 ( \33475 , \9459 , \11918 );
nand \U$33099 ( \33476 , \33474 , \33475 );
nand \U$33100 ( \33477 , \33476 , \10709 );
nand \U$33101 ( \33478 , \33471 , \33477 );
xor \U$33102 ( \33479 , \33468 , \33478 );
not \U$33103 ( \33480 , \33479 );
or \U$33104 ( \33481 , \33458 , \33480 );
nand \U$33105 ( \33482 , \33478 , \33468 );
nand \U$33106 ( \33483 , \33481 , \33482 );
not \U$33107 ( \33484 , \33483 );
not \U$33108 ( \33485 , \33484 );
or \U$33109 ( \33486 , \33410 , \33485 );
nand \U$33110 ( \33487 , \33483 , \33408 );
nand \U$33111 ( \33488 , \33486 , \33487 );
not \U$33112 ( \33489 , \33488 );
or \U$33113 ( \33490 , \33402 , \33489 );
nand \U$33114 ( \33491 , \33409 , \33483 );
nand \U$33115 ( \33492 , \33490 , \33491 );
nand \U$33116 ( \33493 , \33369 , \33492 );
nand \U$33117 ( \33494 , \33363 , \33356 );
and \U$33118 ( \33495 , \33493 , \33494 );
xor \U$33119 ( \33496 , \32737 , \32775 );
not \U$33120 ( \33497 , \33496 );
xor \U$33121 ( \33498 , \32719 , \32708 );
not \U$33122 ( \33499 , \32732 );
and \U$33123 ( \33500 , \33498 , \33499 );
not \U$33124 ( \33501 , \33498 );
and \U$33125 ( \33502 , \33501 , \32732 );
nor \U$33126 ( \33503 , \33500 , \33502 );
not \U$33127 ( \33504 , \33503 );
not \U$33128 ( \33505 , \33063 );
not \U$33129 ( \33506 , \33505 );
not \U$33130 ( \33507 , \33074 );
and \U$33131 ( \33508 , \33506 , \33507 );
and \U$33132 ( \33509 , \33074 , \33505 );
nor \U$33133 ( \33510 , \33508 , \33509 );
not \U$33134 ( \33511 , \33510 );
or \U$33135 ( \33512 , \33504 , \33511 );
not \U$33136 ( \33513 , \5049 );
not \U$33137 ( \33514 , \33054 );
or \U$33138 ( \33515 , \33513 , \33514 );
and \U$33139 ( \33516 , \10461 , \10900 );
not \U$33140 ( \33517 , \10461 );
and \U$33141 ( \33518 , \33517 , RIae79d90_164);
nor \U$33142 ( \33519 , \33516 , \33518 );
not \U$33143 ( \33520 , \33519 );
or \U$33144 ( \33521 , \33520 , \19330 );
nand \U$33145 ( \33522 , \33515 , \33521 );
not \U$33146 ( \33523 , \33522 );
not \U$33147 ( \33524 , \10519 );
not \U$33148 ( \33525 , \33072 );
or \U$33149 ( \33526 , \33524 , \33525 );
and \U$33150 ( \33527 , RIae7a7e0_186, \2090 );
not \U$33151 ( \33528 , RIae7a7e0_186);
and \U$33152 ( \33529 , \33528 , \22917 );
or \U$33153 ( \33530 , \33527 , \33529 );
nand \U$33154 ( \33531 , \33530 , \9549 );
nand \U$33155 ( \33532 , \33526 , \33531 );
not \U$33156 ( \33533 , \33532 );
or \U$33157 ( \33534 , \33523 , \33533 );
or \U$33158 ( \33535 , \33532 , \33522 );
not \U$33159 ( \33536 , \10275 );
not \U$33160 ( \33537 , \33102 );
or \U$33161 ( \33538 , \33536 , \33537 );
and \U$33162 ( \33539 , \1754 , \11207 );
not \U$33163 ( \33540 , \1754 );
and \U$33164 ( \33541 , \33540 , RIae7a8d0_188);
nor \U$33165 ( \33542 , \33539 , \33541 );
nand \U$33166 ( \33543 , \33542 , \16594 );
nand \U$33167 ( \33544 , \33538 , \33543 );
nand \U$33168 ( \33545 , \33535 , \33544 );
nand \U$33169 ( \33546 , \33534 , \33545 );
nand \U$33170 ( \33547 , \33512 , \33546 );
not \U$33171 ( \33548 , \33503 );
not \U$33172 ( \33549 , \33510 );
nand \U$33173 ( \33550 , \33548 , \33549 );
nand \U$33174 ( \33551 , \33547 , \33550 );
not \U$33175 ( \33552 , \33551 );
or \U$33176 ( \33553 , \33497 , \33552 );
not \U$33177 ( \33554 , \9478 );
not \U$33178 ( \33555 , \33007 );
or \U$33179 ( \33556 , \33554 , \33555 );
and \U$33180 ( \33557 , RIae7a6f0_184, \2759 );
not \U$33181 ( \33558 , RIae7a6f0_184);
and \U$33182 ( \33559 , \33558 , \5020 );
nor \U$33183 ( \33560 , \33557 , \33559 );
nand \U$33184 ( \33561 , \33560 , \9473 );
nand \U$33185 ( \33562 , \33556 , \33561 );
not \U$33186 ( \33563 , \33562 );
not \U$33187 ( \33564 , \32853 );
not \U$33188 ( \33565 , \32803 );
not \U$33189 ( \33566 , \33565 );
or \U$33190 ( \33567 , \33564 , \33566 );
or \U$33191 ( \33568 , \33565 , \32853 );
nand \U$33192 ( \33569 , \33567 , \33568 );
not \U$33193 ( \33570 , \2417 );
xor \U$33194 ( \33571 , RIae79c28_161, \9868 );
not \U$33195 ( \33572 , \33571 );
or \U$33196 ( \33573 , \33570 , \33572 );
nand \U$33197 ( \33574 , \32801 , \2418 );
nand \U$33198 ( \33575 , \33573 , \33574 );
not \U$33199 ( \33576 , \32824 );
not \U$33200 ( \33577 , \33576 );
not \U$33201 ( \33578 , \32843 );
or \U$33202 ( \33579 , \33577 , \33578 );
not \U$33203 ( \33580 , \32843 );
nand \U$33204 ( \33581 , \33580 , \32824 );
nand \U$33205 ( \33582 , \33579 , \33581 );
and \U$33206 ( \33583 , \33575 , \33582 );
not \U$33207 ( \33584 , \33575 );
not \U$33208 ( \33585 , \33582 );
and \U$33209 ( \33586 , \33584 , \33585 );
nor \U$33210 ( \33587 , \33583 , \33586 );
not \U$33211 ( \33588 , \33587 );
not \U$33212 ( \33589 , \6091 );
and \U$33213 ( \33590 , RIae79d90_164, \12644 );
not \U$33214 ( \33591 , RIae79d90_164);
not \U$33215 ( \33592 , \10724 );
not \U$33216 ( \33593 , \33592 );
and \U$33217 ( \33594 , \33591 , \33593 );
nor \U$33218 ( \33595 , \33590 , \33594 );
not \U$33219 ( \33596 , \33595 );
or \U$33220 ( \33597 , \33589 , \33596 );
nand \U$33221 ( \33598 , \5048 , \33519 );
nand \U$33222 ( \33599 , \33597 , \33598 );
not \U$33223 ( \33600 , \33599 );
or \U$33224 ( \33601 , \33588 , \33600 );
nand \U$33225 ( \33602 , \33575 , \33582 );
nand \U$33226 ( \33603 , \33601 , \33602 );
xor \U$33227 ( \33604 , \33569 , \33603 );
not \U$33228 ( \33605 , \33604 );
or \U$33229 ( \33606 , \33563 , \33605 );
nand \U$33230 ( \33607 , \33603 , \33569 );
nand \U$33231 ( \33608 , \33606 , \33607 );
xor \U$33232 ( \33609 , \33106 , \33126 );
xor \U$33233 ( \33610 , \33608 , \33609 );
xor \U$33234 ( \33611 , \33035 , \33011 );
and \U$33235 ( \33612 , \33610 , \33611 );
and \U$33236 ( \33613 , \33608 , \33609 );
nor \U$33237 ( \33614 , \33612 , \33613 );
not \U$33238 ( \33615 , \33614 );
nand \U$33239 ( \33616 , \33547 , \33550 );
not \U$33240 ( \33617 , \33496 );
and \U$33241 ( \33618 , \33616 , \33617 );
not \U$33242 ( \33619 , \33616 );
and \U$33243 ( \33620 , \33619 , \33496 );
or \U$33244 ( \33621 , \33618 , \33620 );
nand \U$33245 ( \33622 , \33615 , \33621 );
nand \U$33246 ( \33623 , \33553 , \33622 );
not \U$33247 ( \33624 , \33623 );
and \U$33248 ( \33625 , \33495 , \33624 );
not \U$33249 ( \33626 , \33495 );
and \U$33250 ( \33627 , \33626 , \33623 );
nor \U$33251 ( \33628 , \33625 , \33627 );
not \U$33252 ( \33629 , \33628 );
or \U$33253 ( \33630 , \33308 , \33629 );
not \U$33254 ( \33631 , \33494 );
not \U$33255 ( \33632 , \33493 );
or \U$33256 ( \33633 , \33631 , \33632 );
nand \U$33257 ( \33634 , \33633 , \33623 );
nand \U$33258 ( \33635 , \33630 , \33634 );
nand \U$33259 ( \33636 , \33305 , \33635 );
nand \U$33260 ( \33637 , \33304 , \33303 );
nand \U$33261 ( \33638 , \33636 , \33637 );
xor \U$33262 ( \33639 , \33265 , \33638 );
not \U$33263 ( \33640 , \33216 );
xor \U$33264 ( \33641 , \32686 , \33640 );
xor \U$33265 ( \33642 , \33641 , \32645 );
not \U$33266 ( \33643 , \33642 );
and \U$33267 ( \33644 , \33639 , \33643 );
and \U$33268 ( \33645 , \33265 , \33638 );
nor \U$33269 ( \33646 , \33644 , \33645 );
nor \U$33270 ( \33647 , \33264 , \33646 );
not \U$33271 ( \33648 , \32987 );
nand \U$33272 ( \33649 , \33648 , \33215 );
and \U$33273 ( \33650 , \33649 , \33213 );
not \U$33274 ( \33651 , \33649 );
not \U$33275 ( \33652 , \33213 );
and \U$33276 ( \33653 , \33651 , \33652 );
or \U$33277 ( \33654 , \33650 , \33653 );
xnor \U$33278 ( \33655 , \33628 , \33307 );
not \U$33279 ( \33656 , \33655 );
not \U$33280 ( \33657 , \33614 );
not \U$33281 ( \33658 , \33621 );
or \U$33282 ( \33659 , \33657 , \33658 );
or \U$33283 ( \33660 , \33621 , \33614 );
nand \U$33284 ( \33661 , \33659 , \33660 );
not \U$33285 ( \33662 , \33661 );
not \U$33286 ( \33663 , \33369 );
not \U$33287 ( \33664 , \33492 );
not \U$33288 ( \33665 , \33664 );
and \U$33289 ( \33666 , \33663 , \33665 );
and \U$33290 ( \33667 , \33369 , \33664 );
nor \U$33291 ( \33668 , \33666 , \33667 );
xor \U$33292 ( \33669 , \32870 , \32900 );
not \U$33293 ( \33670 , \9499 );
and \U$33294 ( \33671 , RIae79fe8_169, \29181 );
not \U$33295 ( \33672 , RIae79fe8_169);
and \U$33296 ( \33673 , \33672 , \16766 );
nor \U$33297 ( \33674 , \33671 , \33673 );
not \U$33298 ( \33675 , \33674 );
or \U$33299 ( \33676 , \33670 , \33675 );
nand \U$33300 ( \33677 , \33476 , \9517 );
nand \U$33301 ( \33678 , \33676 , \33677 );
not \U$33302 ( \33679 , \33678 );
not \U$33303 ( \33680 , \2322 );
not \U$33304 ( \33681 , \33430 );
or \U$33305 ( \33682 , \33680 , \33681 );
not \U$33306 ( \33683 , \5344 );
not \U$33307 ( \33684 , \11318 );
or \U$33308 ( \33685 , \33683 , \33684 );
or \U$33309 ( \33686 , \11321 , \19255 );
nand \U$33310 ( \33687 , \33685 , \33686 );
nand \U$33311 ( \33688 , \33687 , \2339 );
nand \U$33312 ( \33689 , \33682 , \33688 );
not \U$33313 ( \33690 , \33689 );
xor \U$33314 ( \33691 , \33446 , \33437 );
not \U$33315 ( \33692 , \33691 );
not \U$33316 ( \33693 , \1919 );
not \U$33317 ( \33694 , \32822 );
or \U$33318 ( \33695 , \33693 , \33694 );
and \U$33319 ( \33696 , \16651 , \3039 );
not \U$33320 ( \33697 , \16651 );
and \U$33321 ( \33698 , \33697 , RIae794a8_145);
nor \U$33322 ( \33699 , \33696 , \33698 );
nand \U$33323 ( \33700 , \33699 , \1932 );
nand \U$33324 ( \33701 , \33695 , \33700 );
not \U$33325 ( \33702 , \33701 );
or \U$33326 ( \33703 , \33692 , \33702 );
or \U$33327 ( \33704 , \33701 , \33691 );
nand \U$33328 ( \33705 , \33703 , \33704 );
not \U$33329 ( \33706 , \33705 );
or \U$33330 ( \33707 , \33690 , \33706 );
not \U$33331 ( \33708 , \33691 );
nand \U$33332 ( \33709 , \33708 , \33701 );
nand \U$33333 ( \33710 , \33707 , \33709 );
not \U$33334 ( \33711 , \33710 );
not \U$33335 ( \33712 , \33711 );
not \U$33336 ( \33713 , \6201 );
not \U$33337 ( \33714 , RIae79ef8_167);
not \U$33338 ( \33715 , \10453 );
or \U$33339 ( \33716 , \33714 , \33715 );
or \U$33340 ( \33717 , \29247 , RIae79ef8_167);
nand \U$33341 ( \33718 , \33716 , \33717 );
not \U$33342 ( \33719 , \33718 );
or \U$33343 ( \33720 , \33713 , \33719 );
nand \U$33344 ( \33721 , \33466 , \6214 );
nand \U$33345 ( \33722 , \33720 , \33721 );
not \U$33346 ( \33723 , \33722 );
or \U$33347 ( \33724 , \33712 , \33723 );
or \U$33348 ( \33725 , \33722 , \33711 );
nand \U$33349 ( \33726 , \33724 , \33725 );
not \U$33350 ( \33727 , \33726 );
or \U$33351 ( \33728 , \33679 , \33727 );
nand \U$33352 ( \33729 , \33722 , \33710 );
nand \U$33353 ( \33730 , \33728 , \33729 );
xor \U$33354 ( \33731 , \33669 , \33730 );
not \U$33355 ( \33732 , \4844 );
not \U$33356 ( \33733 , \10070 );
or \U$33357 ( \33734 , \33732 , \33733 );
not \U$33358 ( \33735 , \10067 );
or \U$33359 ( \33736 , \33735 , \2406 );
nand \U$33360 ( \33737 , \33734 , \33736 );
not \U$33361 ( \33738 , \33737 );
not \U$33362 ( \33739 , \4154 );
or \U$33363 ( \33740 , \33738 , \33739 );
nand \U$33364 ( \33741 , \32868 , \4853 );
nand \U$33365 ( \33742 , \33740 , \33741 );
not \U$33366 ( \33743 , \33742 );
not \U$33367 ( \33744 , \2432 );
xnor \U$33368 ( \33745 , \10740 , RIae79778_151);
not \U$33369 ( \33746 , \33745 );
or \U$33370 ( \33747 , \33744 , \33746 );
nand \U$33371 ( \33748 , \32894 , \15337 );
nand \U$33372 ( \33749 , \33747 , \33748 );
not \U$33373 ( \33750 , \33749 );
and \U$33374 ( \33751 , \33743 , \33750 );
not \U$33375 ( \33752 , \10631 );
not \U$33376 ( \33753 , \33334 );
or \U$33377 ( \33754 , \33752 , \33753 );
not \U$33378 ( \33755 , RIae7a510_180);
not \U$33379 ( \33756 , \28338 );
or \U$33380 ( \33757 , \33755 , \33756 );
or \U$33381 ( \33758 , \28338 , RIae7a510_180);
nand \U$33382 ( \33759 , \33757 , \33758 );
nand \U$33383 ( \33760 , \33759 , \10638 );
nand \U$33384 ( \33761 , \33754 , \33760 );
not \U$33385 ( \33762 , \33761 );
nand \U$33386 ( \33763 , \33742 , \33749 );
and \U$33387 ( \33764 , \33762 , \33763 );
nor \U$33388 ( \33765 , \33751 , \33764 );
and \U$33389 ( \33766 , \33731 , \33765 );
and \U$33390 ( \33767 , \33669 , \33730 );
or \U$33391 ( \33768 , \33766 , \33767 );
not \U$33392 ( \33769 , \33768 );
not \U$33393 ( \33770 , \32905 );
and \U$33394 ( \33771 , \32963 , \33770 );
not \U$33395 ( \33772 , \32963 );
and \U$33396 ( \33773 , \33772 , \32905 );
nor \U$33397 ( \33774 , \33771 , \33773 );
not \U$33398 ( \33775 , \33774 );
or \U$33399 ( \33776 , \33769 , \33775 );
or \U$33400 ( \33777 , \33768 , \33774 );
nand \U$33401 ( \33778 , \33776 , \33777 );
not \U$33402 ( \33779 , \33778 );
xor \U$33403 ( \33780 , \33343 , \33341 );
xnor \U$33404 ( \33781 , \33780 , \33354 );
not \U$33405 ( \33782 , \33781 );
or \U$33406 ( \33783 , \33779 , \33782 );
not \U$33407 ( \33784 , \33774 );
nand \U$33408 ( \33785 , \33784 , \33768 );
nand \U$33409 ( \33786 , \33783 , \33785 );
not \U$33410 ( \33787 , \33786 );
and \U$33411 ( \33788 , \33668 , \33787 );
not \U$33412 ( \33789 , \33668 );
and \U$33413 ( \33790 , \33789 , \33786 );
nor \U$33414 ( \33791 , \33788 , \33790 );
not \U$33415 ( \33792 , \33791 );
or \U$33416 ( \33793 , \33662 , \33792 );
not \U$33417 ( \33794 , \33668 );
nand \U$33418 ( \33795 , \33794 , \33786 );
nand \U$33419 ( \33796 , \33793 , \33795 );
not \U$33420 ( \33797 , \33796 );
not \U$33421 ( \33798 , \33797 );
or \U$33422 ( \33799 , \33656 , \33798 );
xnor \U$33423 ( \33800 , \33397 , \33375 );
xor \U$33424 ( \33801 , \33522 , \33544 );
xnor \U$33425 ( \33802 , \33801 , \33532 );
xor \U$33426 ( \33803 , \33800 , \33802 );
not \U$33427 ( \33804 , \2321 );
not \U$33428 ( \33805 , \33687 );
or \U$33429 ( \33806 , \33804 , \33805 );
and \U$33430 ( \33807 , \10259 , \21036 );
not \U$33431 ( \33808 , \10259 );
and \U$33432 ( \33809 , \33808 , RIae798e0_154);
nor \U$33433 ( \33810 , \33807 , \33809 );
nand \U$33434 ( \33811 , \33810 , \2338 );
nand \U$33435 ( \33812 , \33806 , \33811 );
not \U$33436 ( \33813 , \33812 );
and \U$33437 ( \33814 , \12857 , \2161 );
not \U$33438 ( \33815 , \1918 );
not \U$33439 ( \33816 , \33699 );
or \U$33440 ( \33817 , \33815 , \33816 );
not \U$33441 ( \33818 , RIae794a8_145);
not \U$33442 ( \33819 , \12750 );
or \U$33443 ( \33820 , \33818 , \33819 );
or \U$33444 ( \33821 , \16006 , RIae794a8_145);
nand \U$33445 ( \33822 , \33820 , \33821 );
nand \U$33446 ( \33823 , \33822 , \1931 );
nand \U$33447 ( \33824 , \33817 , \33823 );
not \U$33448 ( \33825 , \33824 );
and \U$33449 ( \33826 , \33814 , \33825 );
not \U$33450 ( \33827 , \33814 );
and \U$33451 ( \33828 , \33827 , \33824 );
or \U$33452 ( \33829 , \33826 , \33828 );
not \U$33453 ( \33830 , \33829 );
or \U$33454 ( \33831 , \33813 , \33830 );
nand \U$33455 ( \33832 , \33824 , \33814 );
nand \U$33456 ( \33833 , \33831 , \33832 );
not \U$33457 ( \33834 , \2007 );
not \U$33458 ( \33835 , \33417 );
or \U$33459 ( \33836 , \33834 , \33835 );
not \U$33460 ( \33837 , \2521 );
not \U$33461 ( \33838 , \11665 );
or \U$33462 ( \33839 , \33837 , \33838 );
or \U$33463 ( \33840 , \10042 , \2521 );
nand \U$33464 ( \33841 , \33839 , \33840 );
nand \U$33465 ( \33842 , \33841 , \1988 );
nand \U$33466 ( \33843 , \33836 , \33842 );
xor \U$33467 ( \33844 , \33833 , \33843 );
not \U$33468 ( \33845 , \33844 );
not \U$33469 ( \33846 , \14940 );
not \U$33470 ( \33847 , \33595 );
or \U$33471 ( \33848 , \33846 , \33847 );
not \U$33472 ( \33849 , \6084 );
not \U$33473 ( \33850 , \10087 );
or \U$33474 ( \33851 , \33849 , \33850 );
or \U$33475 ( \33852 , \10208 , \4968 );
nand \U$33476 ( \33853 , \33851 , \33852 );
nand \U$33477 ( \33854 , \33853 , \5039 );
nand \U$33478 ( \33855 , \33848 , \33854 );
not \U$33479 ( \33856 , \33855 );
or \U$33480 ( \33857 , \33845 , \33856 );
nand \U$33481 ( \33858 , \33843 , \33833 );
nand \U$33482 ( \33859 , \33857 , \33858 );
not \U$33483 ( \33860 , RIae7aab0_192);
not \U$33484 ( \33861 , \33371 );
or \U$33485 ( \33862 , \33860 , \33861 );
not \U$33486 ( \33863 , \14671 );
not \U$33487 ( \33864 , \4023 );
or \U$33488 ( \33865 , \33863 , \33864 );
or \U$33489 ( \33866 , \3094 , \14671 );
nand \U$33490 ( \33867 , \33865 , \33866 );
nand \U$33491 ( \33868 , \33867 , \14668 );
nand \U$33492 ( \33869 , \33862 , \33868 );
xor \U$33493 ( \33870 , \33859 , \33869 );
not \U$33494 ( \33871 , \9473 );
not \U$33495 ( \33872 , \16101 );
not \U$33496 ( \33873 , \23422 );
or \U$33497 ( \33874 , \33872 , \33873 );
nand \U$33498 ( \33875 , \2564 , RIae7a6f0_184);
nand \U$33499 ( \33876 , \33874 , \33875 );
not \U$33500 ( \33877 , \33876 );
or \U$33501 ( \33878 , \33871 , \33877 );
nand \U$33502 ( \33879 , \33560 , \17507 );
nand \U$33503 ( \33880 , \33878 , \33879 );
and \U$33504 ( \33881 , \33870 , \33880 );
and \U$33505 ( \33882 , \33859 , \33869 );
nor \U$33506 ( \33883 , \33881 , \33882 );
and \U$33507 ( \33884 , \33803 , \33883 );
and \U$33508 ( \33885 , \33800 , \33802 );
or \U$33509 ( \33886 , \33884 , \33885 );
not \U$33510 ( \33887 , \33886 );
not \U$33511 ( \33888 , \33887 );
xor \U$33512 ( \33889 , \33317 , \33326 );
xor \U$33513 ( \33890 , \33889 , \33338 );
not \U$33514 ( \33891 , \33890 );
not \U$33515 ( \33892 , \9687 );
and \U$33516 ( \33893 , RIae7a240_174, \21744 );
not \U$33517 ( \33894 , RIae7a240_174);
and \U$33518 ( \33895 , \33894 , \15519 );
or \U$33519 ( \33896 , \33893 , \33895 );
not \U$33520 ( \33897 , \33896 );
or \U$33521 ( \33898 , \33892 , \33897 );
nand \U$33522 ( \33899 , \33315 , \13121 );
nand \U$33523 ( \33900 , \33898 , \33899 );
not \U$33524 ( \33901 , \33900 );
not \U$33525 ( \33902 , \9621 );
not \U$33526 ( \33903 , \33322 );
or \U$33527 ( \33904 , \33902 , \33903 );
not \U$33528 ( \33905 , RIae7a3a8_177);
not \U$33529 ( \33906 , \17242 );
or \U$33530 ( \33907 , \33905 , \33906 );
or \U$33531 ( \33908 , \12687 , RIae7a3a8_177);
nand \U$33532 ( \33909 , \33907 , \33908 );
nand \U$33533 ( \33910 , \33909 , \11014 );
nand \U$33534 ( \33911 , \33904 , \33910 );
not \U$33535 ( \33912 , \33911 );
not \U$33536 ( \33913 , \9792 );
and \U$33537 ( \33914 , \14110 , RIae7a2b8_175);
not \U$33538 ( \33915 , \14110 );
and \U$33539 ( \33916 , \33915 , \28198 );
nor \U$33540 ( \33917 , \33914 , \33916 );
not \U$33541 ( \33918 , \33917 );
or \U$33542 ( \33919 , \33913 , \33918 );
nand \U$33543 ( \33920 , \32952 , \16135 );
nand \U$33544 ( \33921 , \33919 , \33920 );
not \U$33545 ( \33922 , \33921 );
not \U$33546 ( \33923 , \33922 );
or \U$33547 ( \33924 , \33912 , \33923 );
or \U$33548 ( \33925 , \33911 , \33922 );
nand \U$33549 ( \33926 , \33924 , \33925 );
not \U$33550 ( \33927 , \33926 );
or \U$33551 ( \33928 , \33901 , \33927 );
nand \U$33552 ( \33929 , \33921 , \33911 );
nand \U$33553 ( \33930 , \33928 , \33929 );
not \U$33554 ( \33931 , \33930 );
or \U$33555 ( \33932 , \33891 , \33931 );
or \U$33556 ( \33933 , \33930 , \33890 );
buf \U$33557 ( \33934 , \32958 );
not \U$33558 ( \33935 , \32916 );
and \U$33559 ( \33936 , \33934 , \33935 );
not \U$33560 ( \33937 , \33934 );
and \U$33561 ( \33938 , \33937 , \32916 );
nor \U$33562 ( \33939 , \33936 , \33938 );
not \U$33563 ( \33940 , \33939 );
nand \U$33564 ( \33941 , \33933 , \33940 );
nand \U$33565 ( \33942 , \33932 , \33941 );
not \U$33566 ( \33943 , \33942 );
not \U$33567 ( \33944 , \33943 );
and \U$33568 ( \33945 , \33422 , \33451 );
not \U$33569 ( \33946 , \33422 );
and \U$33570 ( \33947 , \33946 , \33452 );
or \U$33571 ( \33948 , \33945 , \33947 );
not \U$33572 ( \33949 , \11205 );
and \U$33573 ( \33950 , RIae7a8d0_188, \3530 );
not \U$33574 ( \33951 , RIae7a8d0_188);
and \U$33575 ( \33952 , \33951 , \3525 );
nor \U$33576 ( \33953 , \33950 , \33952 );
not \U$33577 ( \33954 , \33953 );
or \U$33578 ( \33955 , \33949 , \33954 );
nand \U$33579 ( \33956 , \33542 , \10275 );
nand \U$33580 ( \33957 , \33955 , \33956 );
xor \U$33581 ( \33958 , \33948 , \33957 );
and \U$33582 ( \33959 , \33394 , \9745 );
and \U$33583 ( \33960 , RIae7a060_170, \17596 );
not \U$33584 ( \33961 , RIae7a060_170);
and \U$33585 ( \33962 , \33961 , \1860 );
nor \U$33586 ( \33963 , \33960 , \33962 );
and \U$33587 ( \33964 , \33963 , \17797 );
nor \U$33588 ( \33965 , \33959 , \33964 );
not \U$33589 ( \33966 , \33965 );
and \U$33590 ( \33967 , \33958 , \33966 );
and \U$33591 ( \33968 , \33948 , \33957 );
nor \U$33592 ( \33969 , \33967 , \33968 );
not \U$33593 ( \33970 , \33969 );
not \U$33594 ( \33971 , \33970 );
not \U$33595 ( \33972 , \9758 );
and \U$33596 ( \33973 , RIae7a150_172, \19325 );
not \U$33597 ( \33974 , RIae7a150_172);
and \U$33598 ( \33975 , \33974 , \10812 );
or \U$33599 ( \33976 , \33973 , \33975 );
not \U$33600 ( \33977 , \33976 );
or \U$33601 ( \33978 , \33972 , \33977 );
nand \U$33602 ( \33979 , \33384 , \9776 );
nand \U$33603 ( \33980 , \33978 , \33979 );
not \U$33604 ( \33981 , \10677 );
not \U$33605 ( \33982 , \32911 );
or \U$33606 ( \33983 , \33981 , \33982 );
and \U$33607 ( \33984 , RIae7a498_179, \22952 );
not \U$33608 ( \33985 , RIae7a498_179);
and \U$33609 ( \33986 , \33985 , \12724 );
or \U$33610 ( \33987 , \33984 , \33986 );
nand \U$33611 ( \33988 , \33987 , \11434 );
nand \U$33612 ( \33989 , \33983 , \33988 );
xor \U$33613 ( \33990 , \33980 , \33989 );
not \U$33614 ( \33991 , \10510 );
not \U$33615 ( \33992 , \9529 );
not \U$33616 ( \33993 , \1956 );
or \U$33617 ( \33994 , \33992 , \33993 );
or \U$33618 ( \33995 , \5912 , \9529 );
nand \U$33619 ( \33996 , \33994 , \33995 );
not \U$33620 ( \33997 , \33996 );
or \U$33621 ( \33998 , \33991 , \33997 );
nand \U$33622 ( \33999 , \33530 , \10519 );
nand \U$33623 ( \34000 , \33998 , \33999 );
nand \U$33624 ( \34001 , \33990 , \34000 );
nand \U$33625 ( \34002 , \33989 , \33980 );
and \U$33626 ( \34003 , \34001 , \34002 );
and \U$33627 ( \34004 , \33479 , \33457 );
not \U$33628 ( \34005 , \33479 );
not \U$33629 ( \34006 , \33457 );
and \U$33630 ( \34007 , \34005 , \34006 );
nor \U$33631 ( \34008 , \34004 , \34007 );
not \U$33632 ( \34009 , \34008 );
and \U$33633 ( \34010 , \34003 , \34009 );
not \U$33634 ( \34011 , \34003 );
and \U$33635 ( \34012 , \34011 , \34008 );
nor \U$33636 ( \34013 , \34010 , \34012 );
not \U$33637 ( \34014 , \34013 );
or \U$33638 ( \34015 , \33971 , \34014 );
not \U$33639 ( \34016 , \34002 );
not \U$33640 ( \34017 , \34001 );
or \U$33641 ( \34018 , \34016 , \34017 );
nand \U$33642 ( \34019 , \34018 , \34008 );
nand \U$33643 ( \34020 , \34015 , \34019 );
not \U$33644 ( \34021 , \34020 );
or \U$33645 ( \34022 , \33944 , \34021 );
or \U$33646 ( \34023 , \34020 , \33943 );
nand \U$33647 ( \34024 , \34022 , \34023 );
not \U$33648 ( \34025 , \34024 );
or \U$33649 ( \34026 , \33888 , \34025 );
nand \U$33650 ( \34027 , \34020 , \33942 );
nand \U$33651 ( \34028 , \34026 , \34027 );
not \U$33652 ( \34029 , \33401 );
and \U$33653 ( \34030 , \33488 , \34029 );
not \U$33654 ( \34031 , \33488 );
and \U$33655 ( \34032 , \34031 , \33401 );
nor \U$33656 ( \34033 , \34030 , \34032 );
not \U$33657 ( \34034 , \34033 );
not \U$33658 ( \34035 , \33546 );
not \U$33659 ( \34036 , \33503 );
or \U$33660 ( \34037 , \34035 , \34036 );
or \U$33661 ( \34038 , \33546 , \33503 );
nand \U$33662 ( \34039 , \34037 , \34038 );
and \U$33663 ( \34040 , \34039 , \33549 );
not \U$33664 ( \34041 , \34039 );
and \U$33665 ( \34042 , \34041 , \33510 );
nor \U$33666 ( \34043 , \34040 , \34042 );
not \U$33667 ( \34044 , \34043 );
or \U$33668 ( \34045 , \34034 , \34044 );
or \U$33669 ( \34046 , \34043 , \34033 );
nand \U$33670 ( \34047 , \34045 , \34046 );
not \U$33671 ( \34048 , \34047 );
not \U$33672 ( \34049 , \10573 );
not \U$33673 ( \34050 , \33718 );
or \U$33674 ( \34051 , \34049 , \34050 );
and \U$33675 ( \34052 , RIae79ef8_167, \11186 );
not \U$33676 ( \34053 , RIae79ef8_167);
and \U$33677 ( \34054 , \34053 , \11187 );
nor \U$33678 ( \34055 , \34052 , \34054 );
nand \U$33679 ( \34056 , \34055 , \15989 );
nand \U$33680 ( \34057 , \34051 , \34056 );
not \U$33681 ( \34058 , \34057 );
not \U$33682 ( \34059 , \34058 );
not \U$33683 ( \34060 , \2431 );
and \U$33684 ( \34061 , RIae79778_151, \33414 );
not \U$33685 ( \34062 , RIae79778_151);
and \U$33686 ( \34063 , \34062 , \10031 );
or \U$33687 ( \34064 , \34061 , \34063 );
not \U$33688 ( \34065 , \34064 );
or \U$33689 ( \34066 , \34060 , \34065 );
xor \U$33690 ( \34067 , \10142 , RIae79778_151);
nand \U$33691 ( \34068 , \34067 , \15337 );
nand \U$33692 ( \34069 , \34066 , \34068 );
not \U$33693 ( \34070 , \34069 );
or \U$33694 ( \34071 , \16890 , \1916 );
nand \U$33695 ( \34072 , \34071 , \6997 );
not \U$33696 ( \34073 , \34072 );
not \U$33697 ( \34074 , \1918 );
not \U$33698 ( \34075 , \33822 );
or \U$33699 ( \34076 , \34074 , \34075 );
and \U$33700 ( \34077 , RIae794a8_145, \12857 );
not \U$33701 ( \34078 , RIae794a8_145);
and \U$33702 ( \34079 , \34078 , \17971 );
nor \U$33703 ( \34080 , \34077 , \34079 );
nand \U$33704 ( \34081 , \34080 , \1931 );
nand \U$33705 ( \34082 , \34076 , \34081 );
nand \U$33706 ( \34083 , \34073 , \34082 );
not \U$33707 ( \34084 , \34083 );
not \U$33708 ( \34085 , \2007 );
not \U$33709 ( \34086 , \33841 );
or \U$33710 ( \34087 , \34085 , \34086 );
and \U$33711 ( \34088 , RIae797f0_152, \11240 );
not \U$33712 ( \34089 , RIae797f0_152);
and \U$33713 ( \34090 , \34089 , \32565 );
or \U$33714 ( \34091 , \34088 , \34090 );
nand \U$33715 ( \34092 , \34091 , \1988 );
nand \U$33716 ( \34093 , \34087 , \34092 );
not \U$33717 ( \34094 , \34093 );
or \U$33718 ( \34095 , \34084 , \34094 );
or \U$33719 ( \34096 , \34093 , \34083 );
nand \U$33720 ( \34097 , \34095 , \34096 );
not \U$33721 ( \34098 , \34097 );
or \U$33722 ( \34099 , \34070 , \34098 );
not \U$33723 ( \34100 , \34083 );
nand \U$33724 ( \34101 , \34100 , \34093 );
nand \U$33725 ( \34102 , \34099 , \34101 );
not \U$33726 ( \34103 , \34102 );
or \U$33727 ( \34104 , \34059 , \34103 );
or \U$33728 ( \34105 , \34102 , \34058 );
nand \U$33729 ( \34106 , \34104 , \34105 );
not \U$33730 ( \34107 , \34106 );
not \U$33731 ( \34108 , \9758 );
not \U$33732 ( \34109 , RIae7a150_172);
not \U$33733 ( \34110 , \21873 );
or \U$33734 ( \34111 , \34109 , \34110 );
nand \U$33735 ( \34112 , \4169 , \10672 );
nand \U$33736 ( \34113 , \34111 , \34112 );
not \U$33737 ( \34114 , \34113 );
or \U$33738 ( \34115 , \34108 , \34114 );
nand \U$33739 ( \34116 , \33976 , \9777 );
nand \U$33740 ( \34117 , \34115 , \34116 );
not \U$33741 ( \34118 , \34117 );
or \U$33742 ( \34119 , \34107 , \34118 );
nand \U$33743 ( \34120 , \34102 , \34057 );
nand \U$33744 ( \34121 , \34119 , \34120 );
not \U$33745 ( \34122 , \34121 );
buf \U$33746 ( \34123 , \33587 );
xor \U$33747 ( \34124 , \33599 , \34123 );
not \U$33748 ( \34125 , \34124 );
and \U$33749 ( \34126 , \33674 , \9517 );
not \U$33750 ( \34127 , \10709 );
not \U$33751 ( \34128 , \9417 );
not \U$33752 ( \34129 , RIae79fe8_169);
and \U$33753 ( \34130 , \34128 , \34129 );
and \U$33754 ( \34131 , \9412 , RIae79fe8_169);
nor \U$33755 ( \34132 , \34130 , \34131 );
nor \U$33756 ( \34133 , \34127 , \34132 );
nor \U$33757 ( \34134 , \34126 , \34133 );
not \U$33758 ( \34135 , \34134 );
not \U$33759 ( \34136 , \16135 );
not \U$33760 ( \34137 , \33917 );
or \U$33761 ( \34138 , \34136 , \34137 );
not \U$33762 ( \34139 , RIae7a2b8_175);
not \U$33763 ( \34140 , \13302 );
or \U$33764 ( \34141 , \34139 , \34140 );
nand \U$33765 ( \34142 , \9455 , \28198 );
nand \U$33766 ( \34143 , \34141 , \34142 );
nand \U$33767 ( \34144 , \34143 , \9792 );
nand \U$33768 ( \34145 , \34138 , \34144 );
not \U$33769 ( \34146 , \34145 );
not \U$33770 ( \34147 , \34146 );
or \U$33771 ( \34148 , \34135 , \34147 );
not \U$33772 ( \34149 , \13121 );
not \U$33773 ( \34150 , \33896 );
or \U$33774 ( \34151 , \34149 , \34150 );
not \U$33775 ( \34152 , \11114 );
not \U$33776 ( \34153 , \15088 );
or \U$33777 ( \34154 , \34152 , \34153 );
not \U$33778 ( \34155 , \13290 );
nand \U$33779 ( \34156 , \34155 , RIae7a240_174);
nand \U$33780 ( \34157 , \34154 , \34156 );
nand \U$33781 ( \34158 , \34157 , \19466 );
nand \U$33782 ( \34159 , \34151 , \34158 );
nand \U$33783 ( \34160 , \34148 , \34159 );
not \U$33784 ( \34161 , \34134 );
nand \U$33785 ( \34162 , \34145 , \34161 );
nand \U$33786 ( \34163 , \34160 , \34162 );
not \U$33787 ( \34164 , \34163 );
not \U$33788 ( \34165 , \34164 );
or \U$33789 ( \34166 , \34125 , \34165 );
not \U$33790 ( \34167 , \34162 );
not \U$33791 ( \34168 , \34160 );
or \U$33792 ( \34169 , \34167 , \34168 );
not \U$33793 ( \34170 , \34124 );
nand \U$33794 ( \34171 , \34169 , \34170 );
nand \U$33795 ( \34172 , \34166 , \34171 );
not \U$33796 ( \34173 , \34172 );
or \U$33797 ( \34174 , \34122 , \34173 );
nand \U$33798 ( \34175 , \34163 , \34124 );
nand \U$33799 ( \34176 , \34174 , \34175 );
not \U$33800 ( \34177 , \34176 );
nand \U$33801 ( \34178 , \33909 , \9621 );
not \U$33802 ( \34179 , \11690 );
not \U$33803 ( \34180 , \9317 );
or \U$33804 ( \34181 , \34179 , \34180 );
or \U$33805 ( \34182 , \9317 , \11690 );
nand \U$33806 ( \34183 , \34181 , \34182 );
nand \U$33807 ( \34184 , \34183 , \9644 );
nand \U$33808 ( \34185 , \34178 , \34184 );
not \U$33809 ( \34186 , \33689 );
xor \U$33810 ( \34187 , \33705 , \34186 );
or \U$33811 ( \34188 , \34185 , \34187 );
not \U$33812 ( \34189 , \34184 );
not \U$33813 ( \34190 , \34178 );
or \U$33814 ( \34191 , \34189 , \34190 );
nand \U$33815 ( \34192 , \34191 , \34187 );
nand \U$33816 ( \34193 , \34188 , \34192 );
not \U$33817 ( \34194 , \34193 );
not \U$33818 ( \34195 , \10631 );
not \U$33819 ( \34196 , \33759 );
or \U$33820 ( \34197 , \34195 , \34196 );
and \U$33821 ( \34198 , RIae7a510_180, \6346 );
not \U$33822 ( \34199 , RIae7a510_180);
and \U$33823 ( \34200 , \34199 , \28305 );
or \U$33824 ( \34201 , \34198 , \34200 );
nand \U$33825 ( \34202 , \34201 , \11400 );
nand \U$33826 ( \34203 , \34197 , \34202 );
not \U$33827 ( \34204 , \34203 );
or \U$33828 ( \34205 , \34194 , \34204 );
not \U$33829 ( \34206 , \34184 );
not \U$33830 ( \34207 , \34178 );
or \U$33831 ( \34208 , \34206 , \34207 );
not \U$33832 ( \34209 , \34187 );
nand \U$33833 ( \34210 , \34208 , \34209 );
nand \U$33834 ( \34211 , \34205 , \34210 );
not \U$33835 ( \34212 , \34211 );
not \U$33836 ( \34213 , \2450 );
not \U$33837 ( \34214 , \33745 );
or \U$33838 ( \34215 , \34213 , \34214 );
nand \U$33839 ( \34216 , \34067 , \2432 );
nand \U$33840 ( \34217 , \34215 , \34216 );
not \U$33841 ( \34218 , \2776 );
not \U$33842 ( \34219 , \33571 );
or \U$33843 ( \34220 , \34218 , \34219 );
and \U$33844 ( \34221 , \10000 , \10584 );
not \U$33845 ( \34222 , \10000 );
and \U$33846 ( \34223 , \34222 , RIae79c28_161);
nor \U$33847 ( \34224 , \34221 , \34223 );
nand \U$33848 ( \34225 , \34224 , \2417 );
nand \U$33849 ( \34226 , \34220 , \34225 );
xor \U$33850 ( \34227 , \34217 , \34226 );
not \U$33851 ( \34228 , \4853 );
not \U$33852 ( \34229 , \33737 );
or \U$33853 ( \34230 , \34228 , \34229 );
not \U$33854 ( \34231 , \2406 );
not \U$33855 ( \34232 , \14546 );
or \U$33856 ( \34233 , \34231 , \34232 );
not \U$33857 ( \34234 , \4844 );
nand \U$33858 ( \34235 , \34234 , \10168 );
nand \U$33859 ( \34236 , \34233 , \34235 );
nand \U$33860 ( \34237 , \34236 , \4154 );
nand \U$33861 ( \34238 , \34230 , \34237 );
and \U$33862 ( \34239 , \34227 , \34238 );
and \U$33863 ( \34240 , \34217 , \34226 );
or \U$33864 ( \34241 , \34239 , \34240 );
not \U$33865 ( \34242 , \34241 );
not \U$33866 ( \34243 , \34242 );
xor \U$33867 ( \34244 , \33749 , \33742 );
and \U$33868 ( \34245 , \34244 , \33762 );
not \U$33869 ( \34246 , \34244 );
and \U$33870 ( \34247 , \34246 , \33761 );
or \U$33871 ( \34248 , \34245 , \34247 );
not \U$33872 ( \34249 , \34248 );
or \U$33873 ( \34250 , \34243 , \34249 );
or \U$33874 ( \34251 , \34248 , \34242 );
nand \U$33875 ( \34252 , \34250 , \34251 );
not \U$33876 ( \34253 , \34252 );
or \U$33877 ( \34254 , \34212 , \34253 );
nand \U$33878 ( \34255 , \34248 , \34241 );
nand \U$33879 ( \34256 , \34254 , \34255 );
not \U$33880 ( \34257 , \34256 );
not \U$33881 ( \34258 , \33562 );
and \U$33882 ( \34259 , \33604 , \34258 );
not \U$33883 ( \34260 , \33604 );
and \U$33884 ( \34261 , \34260 , \33562 );
nor \U$33885 ( \34262 , \34259 , \34261 );
not \U$33886 ( \34263 , \34262 );
and \U$33887 ( \34264 , \34257 , \34263 );
and \U$33888 ( \34265 , \34256 , \34262 );
nor \U$33889 ( \34266 , \34264 , \34265 );
not \U$33890 ( \34267 , \34266 );
not \U$33891 ( \34268 , \34267 );
or \U$33892 ( \34269 , \34177 , \34268 );
not \U$33893 ( \34270 , \34262 );
nand \U$33894 ( \34271 , \34270 , \34256 );
nand \U$33895 ( \34272 , \34269 , \34271 );
not \U$33896 ( \34273 , \34272 );
or \U$33897 ( \34274 , \34048 , \34273 );
not \U$33898 ( \34275 , \34033 );
nand \U$33899 ( \34276 , \34275 , \34043 );
nand \U$33900 ( \34277 , \34274 , \34276 );
or \U$33901 ( \34278 , \34028 , \34277 );
and \U$33902 ( \34279 , \33296 , \33282 );
not \U$33903 ( \34280 , \33296 );
not \U$33904 ( \34281 , \33282 );
and \U$33905 ( \34282 , \34280 , \34281 );
nor \U$33906 ( \34283 , \34279 , \34282 );
nand \U$33907 ( \34284 , \34278 , \34283 );
nand \U$33908 ( \34285 , \34028 , \34277 );
nand \U$33909 ( \34286 , \34284 , \34285 );
nand \U$33910 ( \34287 , \33799 , \34286 );
not \U$33911 ( \34288 , \33655 );
nand \U$33912 ( \34289 , \34288 , \33796 );
and \U$33913 ( \34290 , \34287 , \34289 );
xor \U$33914 ( \34291 , \33654 , \34290 );
xor \U$33915 ( \34292 , \33304 , \33635 );
not \U$33916 ( \34293 , \34292 );
not \U$33917 ( \34294 , \33303 );
not \U$33918 ( \34295 , \34294 );
and \U$33919 ( \34296 , \34293 , \34295 );
and \U$33920 ( \34297 , \34292 , \34294 );
nor \U$33921 ( \34298 , \34296 , \34297 );
and \U$33922 ( \34299 , \34291 , \34298 );
and \U$33923 ( \34300 , \33654 , \34290 );
or \U$33924 ( \34301 , \34299 , \34300 );
xor \U$33925 ( \34302 , \33639 , \33642 );
nor \U$33926 ( \34303 , \34301 , \34302 );
or \U$33927 ( \34304 , \33647 , \34303 );
nand \U$33928 ( \34305 , \33264 , \33646 );
nand \U$33929 ( \34306 , \34304 , \34305 );
not \U$33930 ( \34307 , \33260 );
not \U$33931 ( \34308 , \34307 );
not \U$33932 ( \34309 , \33223 );
or \U$33933 ( \34310 , \34308 , \34309 );
nand \U$33934 ( \34311 , \33218 , \32642 );
nand \U$33935 ( \34312 , \34310 , \34311 );
not \U$33936 ( \34313 , \32353 );
not \U$33937 ( \34314 , \34313 );
not \U$33938 ( \34315 , \32638 );
or \U$33939 ( \34316 , \34314 , \34315 );
not \U$33940 ( \34317 , \32356 );
nand \U$33941 ( \34318 , \34317 , \32634 );
nand \U$33942 ( \34319 , \34316 , \34318 );
not \U$33943 ( \34320 , \34319 );
nand \U$33944 ( \34321 , \33241 , \33255 );
not \U$33945 ( \34322 , \33226 );
nand \U$33946 ( \34323 , \34322 , \33237 );
and \U$33947 ( \34324 , \34321 , \34323 );
not \U$33948 ( \34325 , \34324 );
or \U$33949 ( \34326 , \34320 , \34325 );
not \U$33950 ( \34327 , \34323 );
not \U$33951 ( \34328 , \34321 );
or \U$33952 ( \34329 , \34327 , \34328 );
not \U$33953 ( \34330 , \34319 );
nand \U$33954 ( \34331 , \34329 , \34330 );
nand \U$33955 ( \34332 , \34326 , \34331 );
nand \U$33956 ( \34333 , \31200 , \31204 );
buf \U$33957 ( \34334 , \31202 );
not \U$33958 ( \34335 , \34334 );
and \U$33959 ( \34336 , \34333 , \34335 );
not \U$33960 ( \34337 , \34333 );
and \U$33961 ( \34338 , \34337 , \34334 );
nor \U$33962 ( \34339 , \34336 , \34338 );
xor \U$33963 ( \34340 , \34332 , \34339 );
nor \U$33964 ( \34341 , \34312 , \34340 );
or \U$33965 ( \34342 , \34306 , \34341 );
not \U$33966 ( \34343 , \31206 );
not \U$33967 ( \34344 , \31185 );
and \U$33968 ( \34345 , \34343 , \34344 );
and \U$33969 ( \34346 , \31206 , \31185 );
nor \U$33970 ( \34347 , \34345 , \34346 );
and \U$33971 ( \34348 , \34347 , \31189 );
not \U$33972 ( \34349 , \34347 );
and \U$33973 ( \34350 , \34349 , \31188 );
nor \U$33974 ( \34351 , \34348 , \34350 );
not \U$33975 ( \34352 , \34332 );
not \U$33976 ( \34353 , \34339 );
or \U$33977 ( \34354 , \34352 , \34353 );
not \U$33978 ( \34355 , \34323 );
not \U$33979 ( \34356 , \34321 );
or \U$33980 ( \34357 , \34355 , \34356 );
nand \U$33981 ( \34358 , \34357 , \34319 );
nand \U$33982 ( \34359 , \34354 , \34358 );
nand \U$33983 ( \34360 , \34351 , \34359 );
nand \U$33984 ( \34361 , \34340 , \34312 );
and \U$33985 ( \34362 , \34360 , \34361 );
nand \U$33986 ( \34363 , \34342 , \34362 );
not \U$33987 ( \34364 , \34351 );
not \U$33988 ( \34365 , \34359 );
nand \U$33989 ( \34366 , \34364 , \34365 );
and \U$33990 ( \34367 , \32280 , \32278 , \34366 );
nand \U$33991 ( \34368 , \32287 , \34363 , \34367 );
nand \U$33992 ( \34369 , \32285 , \34368 );
not \U$33993 ( \34370 , \32043 );
not \U$33994 ( \34371 , \32249 );
or \U$33995 ( \34372 , \34370 , \34371 );
nand \U$33996 ( \34373 , \34372 , \32259 );
or \U$33997 ( \34374 , \32249 , \32043 );
nand \U$33998 ( \34375 , \34373 , \34374 );
not \U$33999 ( \34376 , \34375 );
buf \U$34000 ( \34377 , \31924 );
not \U$34001 ( \34378 , \34377 );
not \U$34002 ( \34379 , \34378 );
not \U$34003 ( \34380 , \32024 );
or \U$34004 ( \34381 , \34379 , \34380 );
not \U$34005 ( \34382 , \31934 );
nand \U$34006 ( \34383 , \34381 , \34382 );
not \U$34007 ( \34384 , \32024 );
nand \U$34008 ( \34385 , \34384 , \34377 );
nand \U$34009 ( \34386 , \34383 , \34385 );
not \U$34010 ( \34387 , \34386 );
or \U$34011 ( \34388 , \34376 , \34387 );
not \U$34012 ( \34389 , \34386 );
not \U$34013 ( \34390 , \34389 );
not \U$34014 ( \34391 , \34375 );
and \U$34015 ( \34392 , \34390 , \34391 );
and \U$34016 ( \34393 , \34375 , \34389 );
nor \U$34017 ( \34394 , \34392 , \34393 );
not \U$34018 ( \34395 , \32245 );
not \U$34019 ( \34396 , \34395 );
not \U$34020 ( \34397 , \32093 );
or \U$34021 ( \34398 , \34396 , \34397 );
not \U$34022 ( \34399 , \32089 );
nand \U$34023 ( \34400 , \34399 , \32050 );
nand \U$34024 ( \34401 , \34398 , \34400 );
not \U$34025 ( \34402 , \34401 );
not \U$34026 ( \34403 , \32060 );
not \U$34027 ( \34404 , \32083 );
or \U$34028 ( \34405 , \34403 , \34404 );
or \U$34029 ( \34406 , \32060 , \32083 );
nand \U$34030 ( \34407 , \34406 , \32088 );
nand \U$34031 ( \34408 , \34405 , \34407 );
not \U$34032 ( \34409 , \31923 );
not \U$34033 ( \34410 , \31850 );
not \U$34034 ( \34411 , \31916 );
or \U$34035 ( \34412 , \34410 , \34411 );
or \U$34036 ( \34413 , \31850 , \31916 );
nand \U$34037 ( \34414 , \34412 , \34413 );
not \U$34038 ( \34415 , \34414 );
or \U$34039 ( \34416 , \34409 , \34415 );
not \U$34040 ( \34417 , \31850 );
nand \U$34041 ( \34418 , \34417 , \31916 );
nand \U$34042 ( \34419 , \34416 , \34418 );
xor \U$34043 ( \34420 , \34408 , \34419 );
not \U$34044 ( \34421 , \31841 );
or \U$34045 ( \34422 , \31849 , \31811 );
not \U$34046 ( \34423 , \34422 );
or \U$34047 ( \34424 , \34421 , \34423 );
nand \U$34048 ( \34425 , \31849 , \31811 );
nand \U$34049 ( \34426 , \34424 , \34425 );
not \U$34050 ( \34427 , \2767 );
not \U$34051 ( \34428 , \32137 );
or \U$34052 ( \34429 , \34427 , \34428 );
nand \U$34053 ( \34430 , \19773 , \2418 );
nand \U$34054 ( \34431 , \34429 , \34430 );
not \U$34055 ( \34432 , \14768 );
not \U$34056 ( \34433 , \32144 );
or \U$34057 ( \34434 , \34432 , \34433 );
nand \U$34058 ( \34435 , \19866 , \6214 );
nand \U$34059 ( \34436 , \34434 , \34435 );
xor \U$34060 ( \34437 , \34431 , \34436 );
xor \U$34061 ( \34438 , \4169 , RIae79d90_164);
not \U$34062 ( \34439 , \34438 );
not \U$34063 ( \34440 , \5048 );
or \U$34064 ( \34441 , \34439 , \34440 );
nand \U$34065 ( \34442 , \32213 , \5040 );
nand \U$34066 ( \34443 , \34441 , \34442 );
xor \U$34067 ( \34444 , \34437 , \34443 );
xor \U$34068 ( \34445 , \31871 , \31878 );
and \U$34069 ( \34446 , \34445 , \31889 );
and \U$34070 ( \34447 , \31871 , \31878 );
or \U$34071 ( \34448 , \34446 , \34447 );
xor \U$34072 ( \34449 , \34444 , \34448 );
not \U$34073 ( \34450 , \11205 );
not \U$34074 ( \34451 , \31910 );
or \U$34075 ( \34452 , \34450 , \34451 );
nand \U$34076 ( \34453 , \19932 , \10275 );
nand \U$34077 ( \34454 , \34452 , \34453 );
not \U$34078 ( \34455 , \32182 );
not \U$34079 ( \34456 , \32197 );
or \U$34080 ( \34457 , \34455 , \34456 );
not \U$34081 ( \34458 , \32187 );
nand \U$34082 ( \34459 , \34458 , \32193 );
nand \U$34083 ( \34460 , \34457 , \34459 );
not \U$34084 ( \34461 , \4853 );
not \U$34085 ( \34462 , \19784 );
or \U$34086 ( \34463 , \34461 , \34462 );
nand \U$34087 ( \34464 , \32203 , \16804 );
nand \U$34088 ( \34465 , \34463 , \34464 );
xor \U$34089 ( \34466 , \34460 , \34465 );
xor \U$34090 ( \34467 , \34454 , \34466 );
xnor \U$34091 ( \34468 , \34449 , \34467 );
xor \U$34092 ( \34469 , \34426 , \34468 );
not \U$34093 ( \34470 , \9320 );
not \U$34094 ( \34471 , \31964 );
or \U$34095 ( \34472 , \34470 , \34471 );
nand \U$34096 ( \34473 , \18957 , \1820 );
nand \U$34097 ( \34474 , \34472 , \34473 );
xor \U$34098 ( \34475 , \18994 , \18975 );
xor \U$34099 ( \34476 , \34474 , \34475 );
not \U$34100 ( \34477 , \2272 );
not \U$34101 ( \34478 , \31788 );
or \U$34102 ( \34479 , \34477 , \34478 );
nand \U$34103 ( \34480 , \19027 , \2251 );
nand \U$34104 ( \34481 , \34479 , \34480 );
xor \U$34105 ( \34482 , \34476 , \34481 );
xor \U$34106 ( \34483 , \32159 , \32168 );
and \U$34107 ( \34484 , \34483 , \32175 );
and \U$34108 ( \34485 , \32159 , \32168 );
or \U$34109 ( \34486 , \34484 , \34485 );
xor \U$34110 ( \34487 , \34482 , \34486 );
xor \U$34111 ( \34488 , \31904 , \31914 );
not \U$34112 ( \34489 , \31894 );
and \U$34113 ( \34490 , \34488 , \34489 );
and \U$34114 ( \34491 , \31904 , \31914 );
or \U$34115 ( \34492 , \34490 , \34491 );
xor \U$34116 ( \34493 , \34487 , \34492 );
xnor \U$34117 ( \34494 , \34469 , \34493 );
xor \U$34118 ( \34495 , \34420 , \34494 );
not \U$34119 ( \34496 , \34495 );
or \U$34120 ( \34497 , \34402 , \34496 );
or \U$34121 ( \34498 , \34495 , \34401 );
nand \U$34122 ( \34499 , \34497 , \34498 );
nand \U$34123 ( \34500 , \31949 , \32018 );
nand \U$34124 ( \34501 , \31942 , \34500 );
nand \U$34125 ( \34502 , \32021 , \31948 );
nand \U$34126 ( \34503 , \34501 , \34502 );
not \U$34127 ( \34504 , \10638 );
not \U$34128 ( \34505 , \31900 );
or \U$34129 ( \34506 , \34504 , \34505 );
nand \U$34130 ( \34507 , \19908 , \16358 );
nand \U$34131 ( \34508 , \34506 , \34507 );
not \U$34132 ( \34509 , \34508 );
not \U$34133 ( \34510 , \9643 );
not \U$34134 ( \34511 , \32173 );
or \U$34135 ( \34512 , \34510 , \34511 );
nand \U$34136 ( \34513 , \19616 , \9622 );
nand \U$34137 ( \34514 , \34512 , \34513 );
not \U$34138 ( \34515 , \34514 );
not \U$34139 ( \34516 , \34515 );
or \U$34140 ( \34517 , \34509 , \34516 );
not \U$34141 ( \34518 , \34508 );
nand \U$34142 ( \34519 , \34514 , \34518 );
nand \U$34143 ( \34520 , \34517 , \34519 );
not \U$34144 ( \34521 , \9527 );
not \U$34145 ( \34522 , \19604 );
or \U$34146 ( \34523 , \34521 , \34522 );
nand \U$34147 ( \34524 , \32155 , \11439 );
nand \U$34148 ( \34525 , \34523 , \34524 );
not \U$34149 ( \34526 , \34525 );
and \U$34150 ( \34527 , \34520 , \34526 );
not \U$34151 ( \34528 , \34520 );
and \U$34152 ( \34529 , \34528 , \34525 );
nor \U$34153 ( \34530 , \34527 , \34529 );
not \U$34154 ( \34531 , \34530 );
not \U$34155 ( \34532 , \31810 );
not \U$34156 ( \34533 , \31773 );
or \U$34157 ( \34534 , \34532 , \34533 );
not \U$34158 ( \34535 , \31797 );
nand \U$34159 ( \34536 , \34535 , \31805 );
nand \U$34160 ( \34537 , \34534 , \34536 );
not \U$34161 ( \34538 , \34537 );
or \U$34162 ( \34539 , \34531 , \34538 );
or \U$34163 ( \34540 , \34537 , \34530 );
nand \U$34164 ( \34541 , \34539 , \34540 );
not \U$34165 ( \34542 , \9792 );
not \U$34166 ( \34543 , \31826 );
or \U$34167 ( \34544 , \34542 , \34543 );
nand \U$34168 ( \34545 , \19819 , \9814 );
nand \U$34169 ( \34546 , \34544 , \34545 );
not \U$34170 ( \34547 , \13121 );
not \U$34171 ( \34548 , \19625 );
or \U$34172 ( \34549 , \34547 , \34548 );
nand \U$34173 ( \34550 , \32164 , \9688 );
nand \U$34174 ( \34551 , \34549 , \34550 );
not \U$34175 ( \34552 , \34551 );
xor \U$34176 ( \34553 , \34546 , \34552 );
not \U$34177 ( \34554 , \17797 );
not \U$34178 ( \34555 , \31836 );
or \U$34179 ( \34556 , \34554 , \34555 );
nand \U$34180 ( \34557 , \19830 , \11098 );
nand \U$34181 ( \34558 , \34556 , \34557 );
xnor \U$34182 ( \34559 , \34553 , \34558 );
and \U$34183 ( \34560 , \34541 , \34559 );
not \U$34184 ( \34561 , \34541 );
not \U$34185 ( \34562 , \34559 );
and \U$34186 ( \34563 , \34561 , \34562 );
nor \U$34187 ( \34564 , \34560 , \34563 );
nor \U$34188 ( \34565 , \32001 , \32008 );
or \U$34189 ( \34566 , \32013 , \34565 );
nand \U$34190 ( \34567 , \32001 , \32008 );
nand \U$34191 ( \34568 , \34566 , \34567 );
not \U$34192 ( \34569 , \34568 );
xor \U$34193 ( \34570 , \34564 , \34569 );
not \U$34194 ( \34571 , \32000 );
not \U$34195 ( \34572 , \31993 );
or \U$34196 ( \34573 , \34571 , \34572 );
not \U$34197 ( \34574 , \31989 );
nand \U$34198 ( \34575 , \34574 , \31981 );
nand \U$34199 ( \34576 , \34573 , \34575 );
not \U$34200 ( \34577 , \11913 );
not \U$34201 ( \34578 , \31816 );
or \U$34202 ( \34579 , \34577 , \34578 );
nand \U$34203 ( \34580 , \19841 , \9518 );
nand \U$34204 ( \34581 , \34579 , \34580 );
not \U$34205 ( \34582 , \17507 );
and \U$34206 ( \34583 , RIae7a6f0_184, \6147 );
not \U$34207 ( \34584 , RIae7a6f0_184);
and \U$34208 ( \34585 , \34584 , \3689 );
or \U$34209 ( \34586 , \34583 , \34585 );
not \U$34210 ( \34587 , \34586 );
or \U$34211 ( \34588 , \34582 , \34587 );
nand \U$34212 ( \34589 , \9473 , \31874 );
nand \U$34213 ( \34590 , \34588 , \34589 );
xor \U$34214 ( \34591 , \34581 , \34590 );
not \U$34215 ( \34592 , \11087 );
not \U$34216 ( \34593 , \31885 );
or \U$34217 ( \34594 , \34592 , \34593 );
nand \U$34218 ( \34595 , \19859 , \9776 );
nand \U$34219 ( \34596 , \34594 , \34595 );
xor \U$34220 ( \34597 , \34591 , \34596 );
xor \U$34221 ( \34598 , \34576 , \34597 );
not \U$34222 ( \34599 , \31958 );
and \U$34223 ( \34600 , \31980 , \31968 );
not \U$34224 ( \34601 , \31980 );
and \U$34225 ( \34602 , \34601 , \31969 );
nor \U$34226 ( \34603 , \34600 , \34602 );
not \U$34227 ( \34604 , \34603 );
or \U$34228 ( \34605 , \34599 , \34604 );
nand \U$34229 ( \34606 , \31980 , \31968 );
nand \U$34230 ( \34607 , \34605 , \34606 );
not \U$34231 ( \34608 , \34607 );
and \U$34232 ( \34609 , \31792 , \31785 );
and \U$34233 ( \34610 , \31784 , \31779 );
nor \U$34234 ( \34611 , \34609 , \34610 );
not \U$34235 ( \34612 , \34611 );
and \U$34236 ( \34613 , \34608 , \34612 );
and \U$34237 ( \34614 , \34607 , \34611 );
nor \U$34238 ( \34615 , \34613 , \34614 );
not \U$34239 ( \34616 , \32103 );
not \U$34240 ( \34617 , \32113 );
or \U$34241 ( \34618 , \34616 , \34617 );
not \U$34242 ( \34619 , \32103 );
nand \U$34243 ( \34620 , \34619 , \32114 );
nand \U$34244 ( \34621 , \32121 , \34620 );
nand \U$34245 ( \34622 , \34618 , \34621 );
not \U$34246 ( \34623 , \34622 );
and \U$34247 ( \34624 , \34615 , \34623 );
not \U$34248 ( \34625 , \34615 );
and \U$34249 ( \34626 , \34625 , \34622 );
nor \U$34250 ( \34627 , \34624 , \34626 );
xnor \U$34251 ( \34628 , \34598 , \34627 );
not \U$34252 ( \34629 , \34628 );
xnor \U$34253 ( \34630 , \34570 , \34629 );
or \U$34254 ( \34631 , \34503 , \34630 );
not \U$34255 ( \34632 , \34502 );
not \U$34256 ( \34633 , \34501 );
or \U$34257 ( \34634 , \34632 , \34633 );
nand \U$34258 ( \34635 , \34634 , \34630 );
nand \U$34259 ( \34636 , \34631 , \34635 );
xor \U$34260 ( \34637 , \32082 , \32067 );
not \U$34261 ( \34638 , \32077 );
and \U$34262 ( \34639 , \34637 , \34638 );
and \U$34263 ( \34640 , \32082 , \32067 );
or \U$34264 ( \34641 , \34639 , \34640 );
not \U$34265 ( \34642 , \34641 );
not \U$34266 ( \34643 , \34642 );
xor \U$34267 ( \34644 , \32132 , \32141 );
and \U$34268 ( \34645 , \34644 , \32148 );
and \U$34269 ( \34646 , \32132 , \32141 );
or \U$34270 ( \34647 , \34645 , \34646 );
not \U$34271 ( \34648 , \9576 );
not \U$34272 ( \34649 , \32117 );
or \U$34273 ( \34650 , \34648 , \34649 );
nand \U$34274 ( \34651 , \19663 , \2450 );
nand \U$34275 ( \34652 , \34650 , \34651 );
not \U$34276 ( \34653 , \34652 );
not \U$34277 ( \34654 , \2011 );
not \U$34278 ( \34655 , \19055 );
or \U$34279 ( \34656 , \34654 , \34655 );
nand \U$34280 ( \34657 , \31954 , \2063 );
nand \U$34281 ( \34658 , \34656 , \34657 );
not \U$34282 ( \34659 , \2188 );
not \U$34283 ( \34660 , \31976 );
or \U$34284 ( \34661 , \34659 , \34660 );
nand \U$34285 ( \34662 , \19729 , \2162 );
nand \U$34286 ( \34663 , \34661 , \34662 );
not \U$34287 ( \34664 , \34663 );
and \U$34288 ( \34665 , \34658 , \34664 );
not \U$34289 ( \34666 , \34658 );
and \U$34290 ( \34667 , \34666 , \34663 );
nor \U$34291 ( \34668 , \34665 , \34667 );
not \U$34292 ( \34669 , \34668 );
and \U$34293 ( \34670 , \34653 , \34669 );
and \U$34294 ( \34671 , \34652 , \34668 );
nor \U$34295 ( \34672 , \34670 , \34671 );
not \U$34296 ( \34673 , \34672 );
and \U$34297 ( \34674 , \34647 , \34673 );
not \U$34298 ( \34675 , \34647 );
and \U$34299 ( \34676 , \34675 , \34672 );
nor \U$34300 ( \34677 , \34674 , \34676 );
not \U$34301 ( \34678 , \32217 );
not \U$34302 ( \34679 , \32208 );
or \U$34303 ( \34680 , \34678 , \34679 );
nand \U$34304 ( \34681 , \32207 , \32198 );
nand \U$34305 ( \34682 , \34680 , \34681 );
not \U$34306 ( \34683 , \34682 );
and \U$34307 ( \34684 , \34677 , \34683 );
not \U$34308 ( \34685 , \34677 );
and \U$34309 ( \34686 , \34685 , \34682 );
nor \U$34310 ( \34687 , \34684 , \34686 );
not \U$34311 ( \34688 , \34687 );
not \U$34312 ( \34689 , \32232 );
or \U$34313 ( \34690 , \32225 , \32218 );
not \U$34314 ( \34691 , \34690 );
or \U$34315 ( \34692 , \34689 , \34691 );
nand \U$34316 ( \34693 , \32218 , \32225 );
nand \U$34317 ( \34694 , \34692 , \34693 );
not \U$34318 ( \34695 , \34694 );
or \U$34319 ( \34696 , \34688 , \34695 );
or \U$34320 ( \34697 , \34694 , \34687 );
nand \U$34321 ( \34698 , \34696 , \34697 );
not \U$34322 ( \34699 , \34698 );
or \U$34323 ( \34700 , \34643 , \34699 );
or \U$34324 ( \34701 , \34698 , \34642 );
nand \U$34325 ( \34702 , \34700 , \34701 );
not \U$34326 ( \34703 , \34702 );
not \U$34327 ( \34704 , \34703 );
nor \U$34328 ( \34705 , \32244 , \32177 );
or \U$34329 ( \34706 , \34705 , \32233 );
nand \U$34330 ( \34707 , \32244 , \32177 );
nand \U$34331 ( \34708 , \34706 , \34707 );
not \U$34332 ( \34709 , \34708 );
or \U$34333 ( \34710 , \34704 , \34709 );
not \U$34334 ( \34711 , \34708 );
nand \U$34335 ( \34712 , \34711 , \34702 );
nand \U$34336 ( \34713 , \34710 , \34712 );
not \U$34337 ( \34714 , \34713 );
xor \U$34338 ( \34715 , \32122 , \32149 );
and \U$34339 ( \34716 , \34715 , \32176 );
and \U$34340 ( \34717 , \32122 , \32149 );
or \U$34341 ( \34718 , \34716 , \34717 );
not \U$34342 ( \34719 , \31890 );
nor \U$34343 ( \34720 , \34719 , \31862 );
or \U$34344 ( \34721 , \34720 , \31915 );
nand \U$34345 ( \34722 , \34719 , \31862 );
nand \U$34346 ( \34723 , \34721 , \34722 );
xor \U$34347 ( \34724 , \34718 , \34723 );
not \U$34348 ( \34725 , \10677 );
not \U$34349 ( \34726 , \19879 );
or \U$34350 ( \34727 , \34725 , \34726 );
nand \U$34351 ( \34728 , \31869 , \10696 );
nand \U$34352 ( \34729 , \34727 , \34728 );
buf \U$34353 ( \34730 , \19699 );
buf \U$34354 ( \34731 , \19671 );
not \U$34355 ( \34732 , \34731 );
and \U$34356 ( \34733 , \34730 , \34732 );
not \U$34357 ( \34734 , \34730 );
and \U$34358 ( \34735 , \34734 , \34731 );
nor \U$34359 ( \34736 , \34733 , \34735 );
not \U$34360 ( \34737 , \16383 );
not \U$34361 ( \34738 , \31769 );
or \U$34362 ( \34739 , \34737 , \34738 );
not \U$34363 ( \34740 , RIae7aa38_191);
not \U$34364 ( \34741 , \2175 );
or \U$34365 ( \34742 , \34740 , \34741 );
or \U$34366 ( \34743 , \2175 , RIae7aa38_191);
nand \U$34367 ( \34744 , \34742 , \34743 );
nand \U$34368 ( \34745 , \34744 , RIae7aab0_192);
nand \U$34369 ( \34746 , \34739 , \34745 );
xnor \U$34370 ( \34747 , \34736 , \34746 );
xor \U$34371 ( \34748 , \34729 , \34747 );
not \U$34372 ( \34749 , \2467 );
not \U$34373 ( \34750 , \19764 );
or \U$34374 ( \34751 , \34749 , \34750 );
nand \U$34375 ( \34752 , \32128 , \9828 );
nand \U$34376 ( \34753 , \34751 , \34752 );
not \U$34377 ( \34754 , \2339 );
not \U$34378 ( \34755 , \32109 );
or \U$34379 ( \34756 , \34754 , \34755 );
nand \U$34380 ( \34757 , \19738 , \2322 );
nand \U$34381 ( \34758 , \34756 , \34757 );
not \U$34382 ( \34759 , \34758 );
xor \U$34383 ( \34760 , \34753 , \34759 );
not \U$34384 ( \34761 , \1988 );
not \U$34385 ( \34762 , \32099 );
or \U$34386 ( \34763 , \34761 , \34762 );
nand \U$34387 ( \34764 , \19715 , \2007 );
nand \U$34388 ( \34765 , \34763 , \34764 );
xor \U$34389 ( \34766 , \34760 , \34765 );
not \U$34390 ( \34767 , \34766 );
xor \U$34391 ( \34768 , \31820 , \31830 );
and \U$34392 ( \34769 , \34768 , \31840 );
and \U$34393 ( \34770 , \31820 , \31830 );
or \U$34394 ( \34771 , \34769 , \34770 );
not \U$34395 ( \34772 , \34771 );
or \U$34396 ( \34773 , \34767 , \34772 );
or \U$34397 ( \34774 , \34771 , \34766 );
nand \U$34398 ( \34775 , \34773 , \34774 );
xnor \U$34399 ( \34776 , \34748 , \34775 );
not \U$34400 ( \34777 , \34776 );
xor \U$34401 ( \34778 , \34724 , \34777 );
not \U$34402 ( \34779 , \34778 );
and \U$34403 ( \34780 , \34714 , \34779 );
and \U$34404 ( \34781 , \34713 , \34778 );
nor \U$34405 ( \34782 , \34780 , \34781 );
not \U$34406 ( \34783 , \34782 );
and \U$34407 ( \34784 , \34636 , \34783 );
not \U$34408 ( \34785 , \34636 );
and \U$34409 ( \34786 , \34785 , \34782 );
nor \U$34410 ( \34787 , \34784 , \34786 );
not \U$34411 ( \34788 , \34787 );
and \U$34412 ( \34789 , \34499 , \34788 );
not \U$34413 ( \34790 , \34499 );
and \U$34414 ( \34791 , \34790 , \34787 );
nor \U$34415 ( \34792 , \34789 , \34791 );
not \U$34416 ( \34793 , \34792 );
or \U$34417 ( \34794 , \34394 , \34793 );
nand \U$34418 ( \34795 , \34388 , \34794 );
not \U$34419 ( \34796 , \34795 );
not \U$34420 ( \34797 , \34466 );
not \U$34421 ( \34798 , \34454 );
or \U$34422 ( \34799 , \34797 , \34798 );
nand \U$34423 ( \34800 , \34465 , \34460 );
nand \U$34424 ( \34801 , \34799 , \34800 );
xor \U$34425 ( \34802 , \19608 , \19618 );
xor \U$34426 ( \34803 , \34802 , \19629 );
xor \U$34427 ( \34804 , \34801 , \34803 );
not \U$34428 ( \34805 , \9705 );
not \U$34429 ( \34806 , \19066 );
or \U$34430 ( \34807 , \34805 , \34806 );
nand \U$34431 ( \34808 , \34586 , \9473 );
nand \U$34432 ( \34809 , \34807 , \34808 );
not \U$34433 ( \34810 , RIae7aab0_192);
not \U$34434 ( \34811 , \19392 );
or \U$34435 ( \34812 , \34810 , \34811 );
nand \U$34436 ( \34813 , \34744 , \14669 );
nand \U$34437 ( \34814 , \34812 , \34813 );
or \U$34438 ( \34815 , \34474 , \34475 );
nand \U$34439 ( \34816 , \34815 , \34481 );
nand \U$34440 ( \34817 , \34474 , \34475 );
nand \U$34441 ( \34818 , \34816 , \34817 );
xor \U$34442 ( \34819 , \34814 , \34818 );
buf \U$34443 ( \34820 , \34819 );
xor \U$34444 ( \34821 , \34809 , \34820 );
xor \U$34445 ( \34822 , \34804 , \34821 );
or \U$34446 ( \34823 , \34623 , \34615 );
not \U$34447 ( \34824 , \34607 );
or \U$34448 ( \34825 , \34824 , \34611 );
nand \U$34449 ( \34826 , \34823 , \34825 );
not \U$34450 ( \34827 , \34682 );
not \U$34451 ( \34828 , \34677 );
or \U$34452 ( \34829 , \34827 , \34828 );
nand \U$34453 ( \34830 , \34647 , \34673 );
nand \U$34454 ( \34831 , \34829 , \34830 );
xor \U$34455 ( \34832 , \34826 , \34831 );
xor \U$34456 ( \34833 , \34482 , \34486 );
and \U$34457 ( \34834 , \34833 , \34492 );
and \U$34458 ( \34835 , \34482 , \34486 );
or \U$34459 ( \34836 , \34834 , \34835 );
and \U$34460 ( \34837 , \34832 , \34836 );
not \U$34461 ( \34838 , \34832 );
not \U$34462 ( \34839 , \34836 );
and \U$34463 ( \34840 , \34838 , \34839 );
nor \U$34464 ( \34841 , \34837 , \34840 );
xor \U$34465 ( \34842 , \34822 , \34841 );
not \U$34466 ( \34843 , \34641 );
not \U$34467 ( \34844 , \34698 );
or \U$34468 ( \34845 , \34843 , \34844 );
not \U$34469 ( \34846 , \34687 );
nand \U$34470 ( \34847 , \34846 , \34694 );
nand \U$34471 ( \34848 , \34845 , \34847 );
not \U$34472 ( \34849 , \34848 );
and \U$34473 ( \34850 , \34842 , \34849 );
not \U$34474 ( \34851 , \34842 );
and \U$34475 ( \34852 , \34851 , \34848 );
nor \U$34476 ( \34853 , \34850 , \34852 );
not \U$34477 ( \34854 , \34853 );
not \U$34478 ( \34855 , \34854 );
not \U$34479 ( \34856 , \34777 );
not \U$34480 ( \34857 , \34723 );
not \U$34481 ( \34858 , \34857 );
or \U$34482 ( \34859 , \34856 , \34858 );
not \U$34483 ( \34860 , \34723 );
not \U$34484 ( \34861 , \34776 );
or \U$34485 ( \34862 , \34860 , \34861 );
nand \U$34486 ( \34863 , \34862 , \34718 );
nand \U$34487 ( \34864 , \34859 , \34863 );
or \U$34488 ( \34865 , \34448 , \34467 );
nand \U$34489 ( \34866 , \34865 , \34444 );
nand \U$34490 ( \34867 , \34448 , \34467 );
nand \U$34491 ( \34868 , \34866 , \34867 );
not \U$34492 ( \34869 , \19009 );
not \U$34493 ( \34870 , \18959 );
not \U$34494 ( \34871 , \34870 );
and \U$34495 ( \34872 , \34869 , \34871 );
and \U$34496 ( \34873 , \19009 , \34870 );
nor \U$34497 ( \34874 , \34872 , \34873 );
not \U$34498 ( \34875 , \34874 );
not \U$34499 ( \34876 , \34668 );
not \U$34500 ( \34877 , \34876 );
not \U$34501 ( \34878 , \34652 );
or \U$34502 ( \34879 , \34877 , \34878 );
not \U$34503 ( \34880 , \34664 );
nand \U$34504 ( \34881 , \34880 , \34658 );
nand \U$34505 ( \34882 , \34879 , \34881 );
not \U$34506 ( \34883 , \34882 );
or \U$34507 ( \34884 , \34875 , \34883 );
or \U$34508 ( \34885 , \34882 , \34874 );
nand \U$34509 ( \34886 , \34884 , \34885 );
not \U$34510 ( \34887 , \34753 );
not \U$34511 ( \34888 , \34765 );
not \U$34512 ( \34889 , \34759 );
or \U$34513 ( \34890 , \34888 , \34889 );
or \U$34514 ( \34891 , \34765 , \34759 );
nand \U$34515 ( \34892 , \34890 , \34891 );
not \U$34516 ( \34893 , \34892 );
or \U$34517 ( \34894 , \34887 , \34893 );
nand \U$34518 ( \34895 , \34758 , \34765 );
nand \U$34519 ( \34896 , \34894 , \34895 );
xor \U$34520 ( \34897 , \34886 , \34896 );
xnor \U$34521 ( \34898 , \19029 , \19058 );
not \U$34522 ( \34899 , \34898 );
not \U$34523 ( \34900 , \34436 );
not \U$34524 ( \34901 , \34431 );
nand \U$34525 ( \34902 , \34900 , \34901 );
not \U$34526 ( \34903 , \34902 );
not \U$34527 ( \34904 , \34443 );
or \U$34528 ( \34905 , \34903 , \34904 );
not \U$34529 ( \34906 , \34901 );
nand \U$34530 ( \34907 , \34906 , \34436 );
nand \U$34531 ( \34908 , \34905 , \34907 );
not \U$34532 ( \34909 , \34908 );
or \U$34533 ( \34910 , \34899 , \34909 );
or \U$34534 ( \34911 , \34908 , \34898 );
nand \U$34535 ( \34912 , \34910 , \34911 );
not \U$34536 ( \34913 , \34912 );
not \U$34537 ( \34914 , \19754 );
not \U$34538 ( \34915 , \19732 );
and \U$34539 ( \34916 , \34914 , \34915 );
and \U$34540 ( \34917 , \19754 , \19732 );
nor \U$34541 ( \34918 , \34916 , \34917 );
xor \U$34542 ( \34919 , \19751 , \34918 );
not \U$34543 ( \34920 , \34919 );
and \U$34544 ( \34921 , \34913 , \34920 );
and \U$34545 ( \34922 , \34912 , \34919 );
nor \U$34546 ( \34923 , \34921 , \34922 );
or \U$34547 ( \34924 , \34897 , \34923 );
nand \U$34548 ( \34925 , \34923 , \34897 );
nand \U$34549 ( \34926 , \34924 , \34925 );
xor \U$34550 ( \34927 , \34868 , \34926 );
xor \U$34551 ( \34928 , \34864 , \34927 );
not \U$34552 ( \34929 , \34559 );
not \U$34553 ( \34930 , \34541 );
or \U$34554 ( \34931 , \34929 , \34930 );
not \U$34555 ( \34932 , \34530 );
nand \U$34556 ( \34933 , \34932 , \34537 );
nand \U$34557 ( \34934 , \34931 , \34933 );
not \U$34558 ( \34935 , \34771 );
nand \U$34559 ( \34936 , \34935 , \34766 );
not \U$34560 ( \34937 , \34936 );
xor \U$34561 ( \34938 , \34736 , \34729 );
xnor \U$34562 ( \34939 , \34938 , \34746 );
not \U$34563 ( \34940 , \34939 );
or \U$34564 ( \34941 , \34937 , \34940 );
not \U$34565 ( \34942 , \34766 );
nand \U$34566 ( \34943 , \34942 , \34771 );
nand \U$34567 ( \34944 , \34941 , \34943 );
xor \U$34568 ( \34945 , \34934 , \34944 );
not \U$34569 ( \34946 , \34508 );
not \U$34570 ( \34947 , \34514 );
or \U$34571 ( \34948 , \34946 , \34947 );
nand \U$34572 ( \34949 , \34948 , \34526 );
nand \U$34573 ( \34950 , \34515 , \34518 );
and \U$34574 ( \34951 , \34949 , \34950 );
xor \U$34575 ( \34952 , \34581 , \34590 );
and \U$34576 ( \34953 , \34952 , \34596 );
and \U$34577 ( \34954 , \34581 , \34590 );
or \U$34578 ( \34955 , \34953 , \34954 );
xor \U$34579 ( \34956 , \34951 , \34955 );
not \U$34580 ( \34957 , \34729 );
not \U$34581 ( \34958 , \34747 );
or \U$34582 ( \34959 , \34957 , \34958 );
not \U$34583 ( \34960 , \34736 );
nand \U$34584 ( \34961 , \34960 , \34746 );
nand \U$34585 ( \34962 , \34959 , \34961 );
xor \U$34586 ( \34963 , \34956 , \34962 );
xor \U$34587 ( \34964 , \34945 , \34963 );
and \U$34588 ( \34965 , \34928 , \34964 );
not \U$34589 ( \34966 , \34928 );
not \U$34590 ( \34967 , \34964 );
and \U$34591 ( \34968 , \34966 , \34967 );
nor \U$34592 ( \34969 , \34965 , \34968 );
not \U$34593 ( \34970 , \34969 );
not \U$34594 ( \34971 , \34970 );
or \U$34595 ( \34972 , \34855 , \34971 );
nand \U$34596 ( \34973 , \34853 , \34969 );
nand \U$34597 ( \34974 , \34972 , \34973 );
not \U$34598 ( \34975 , \34778 );
not \U$34599 ( \34976 , \34975 );
not \U$34600 ( \34977 , \34713 );
or \U$34601 ( \34978 , \34976 , \34977 );
nand \U$34602 ( \34979 , \34702 , \34708 );
nand \U$34603 ( \34980 , \34978 , \34979 );
not \U$34604 ( \34981 , \34980 );
and \U$34605 ( \34982 , \34974 , \34981 );
not \U$34606 ( \34983 , \34974 );
and \U$34607 ( \34984 , \34983 , \34980 );
nor \U$34608 ( \34985 , \34982 , \34984 );
or \U$34609 ( \34986 , \34495 , \34401 );
not \U$34610 ( \34987 , \34986 );
not \U$34611 ( \34988 , \34787 );
or \U$34612 ( \34989 , \34987 , \34988 );
nand \U$34613 ( \34990 , \34495 , \34401 );
nand \U$34614 ( \34991 , \34989 , \34990 );
not \U$34615 ( \34992 , \34991 );
xor \U$34616 ( \34993 , \34985 , \34992 );
not \U$34617 ( \34994 , \34636 );
not \U$34618 ( \34995 , \34783 );
or \U$34619 ( \34996 , \34994 , \34995 );
not \U$34620 ( \34997 , \34630 );
nand \U$34621 ( \34998 , \34997 , \34503 );
nand \U$34622 ( \34999 , \34996 , \34998 );
not \U$34623 ( \35000 , \34999 );
xor \U$34624 ( \35001 , \19766 , \19775 );
xor \U$34625 ( \35002 , \35001 , \19786 );
xnor \U$34626 ( \35003 , \19705 , \19717 );
nor \U$34627 ( \35004 , \35002 , \35003 );
not \U$34628 ( \35005 , \35004 );
nand \U$34629 ( \35006 , \35002 , \35003 );
nand \U$34630 ( \35007 , \35005 , \35006 );
not \U$34631 ( \35008 , \35007 );
not \U$34632 ( \35009 , \34558 );
not \U$34633 ( \35010 , \34546 );
not \U$34634 ( \35011 , \35010 );
not \U$34635 ( \35012 , \34551 );
or \U$34636 ( \35013 , \35011 , \35012 );
or \U$34637 ( \35014 , \34551 , \35010 );
nand \U$34638 ( \35015 , \35013 , \35014 );
not \U$34639 ( \35016 , \35015 );
or \U$34640 ( \35017 , \35009 , \35016 );
not \U$34641 ( \35018 , \35010 );
nand \U$34642 ( \35019 , \35018 , \34551 );
nand \U$34643 ( \35020 , \35017 , \35019 );
not \U$34644 ( \35021 , \35020 );
or \U$34645 ( \35022 , \35008 , \35021 );
or \U$34646 ( \35023 , \35020 , \35007 );
nand \U$34647 ( \35024 , \35022 , \35023 );
buf \U$34648 ( \35025 , \34597 );
or \U$34649 ( \35026 , \35025 , \34627 );
nand \U$34650 ( \35027 , \35026 , \34576 );
nand \U$34651 ( \35028 , \35025 , \34627 );
and \U$34652 ( \35029 , \35027 , \35028 );
xor \U$34653 ( \35030 , \35024 , \35029 );
xor \U$34654 ( \35031 , \19934 , \19922 );
and \U$34655 ( \35032 , \19847 , \19821 );
not \U$34656 ( \35033 , \19847 );
not \U$34657 ( \35034 , \19821 );
and \U$34658 ( \35035 , \35033 , \35034 );
nor \U$34659 ( \35036 , \35032 , \35035 );
xor \U$34660 ( \35037 , \35031 , \35036 );
not \U$34661 ( \35038 , \19885 );
xor \U$34662 ( \35039 , \19881 , \19870 );
not \U$34663 ( \35040 , \35039 );
or \U$34664 ( \35041 , \35038 , \35040 );
not \U$34665 ( \35042 , \35039 );
not \U$34666 ( \35043 , \19885 );
nand \U$34667 ( \35044 , \35042 , \35043 );
nand \U$34668 ( \35045 , \35041 , \35044 );
xor \U$34669 ( \35046 , \35037 , \35045 );
xor \U$34670 ( \35047 , \35030 , \35046 );
not \U$34671 ( \35048 , \35047 );
not \U$34672 ( \35049 , \34629 );
not \U$34673 ( \35050 , \34564 );
or \U$34674 ( \35051 , \35049 , \35050 );
not \U$34675 ( \35052 , \34628 );
not \U$34676 ( \35053 , \34564 );
not \U$34677 ( \35054 , \35053 );
or \U$34678 ( \35055 , \35052 , \35054 );
nand \U$34679 ( \35056 , \35055 , \34569 );
nand \U$34680 ( \35057 , \35051 , \35056 );
not \U$34681 ( \35058 , \34426 );
not \U$34682 ( \35059 , \34468 );
not \U$34683 ( \35060 , \35059 );
or \U$34684 ( \35061 , \35058 , \35060 );
not \U$34685 ( \35062 , \34468 );
not \U$34686 ( \35063 , \34426 );
not \U$34687 ( \35064 , \35063 );
or \U$34688 ( \35065 , \35062 , \35064 );
nand \U$34689 ( \35066 , \35065 , \34493 );
nand \U$34690 ( \35067 , \35061 , \35066 );
and \U$34691 ( \35068 , \35057 , \35067 );
not \U$34692 ( \35069 , \35057 );
not \U$34693 ( \35070 , \35067 );
and \U$34694 ( \35071 , \35069 , \35070 );
nor \U$34695 ( \35072 , \35068 , \35071 );
not \U$34696 ( \35073 , \35072 );
or \U$34697 ( \35074 , \35048 , \35073 );
or \U$34698 ( \35075 , \35072 , \35047 );
nand \U$34699 ( \35076 , \35074 , \35075 );
not \U$34700 ( \35077 , \35076 );
xor \U$34701 ( \35078 , \34408 , \34419 );
and \U$34702 ( \35079 , \35078 , \34494 );
and \U$34703 ( \35080 , \34408 , \34419 );
or \U$34704 ( \35081 , \35079 , \35080 );
not \U$34705 ( \35082 , \35081 );
and \U$34706 ( \35083 , \35077 , \35082 );
and \U$34707 ( \35084 , \35081 , \35076 );
nor \U$34708 ( \35085 , \35083 , \35084 );
not \U$34709 ( \35086 , \35085 );
or \U$34710 ( \35087 , \35000 , \35086 );
or \U$34711 ( \35088 , \34999 , \35085 );
nand \U$34712 ( \35089 , \35087 , \35088 );
xor \U$34713 ( \35090 , \34993 , \35089 );
nand \U$34714 ( \35091 , \34796 , \35090 );
buf \U$34715 ( \35092 , \32026 );
or \U$34716 ( \35093 , \32260 , \35092 );
buf \U$34717 ( \35094 , \32032 );
nand \U$34718 ( \35095 , \35093 , \35094 );
not \U$34719 ( \35096 , \35095 );
not \U$34720 ( \35097 , \34394 );
not \U$34721 ( \35098 , \34792 );
and \U$34722 ( \35099 , \35097 , \35098 );
and \U$34723 ( \35100 , \34394 , \34792 );
nor \U$34724 ( \35101 , \35099 , \35100 );
nand \U$34725 ( \35102 , \35096 , \35101 );
and \U$34726 ( \35103 , \35091 , \35102 );
xor \U$34727 ( \35104 , \19070 , \19063 );
not \U$34728 ( \35105 , \34919 );
not \U$34729 ( \35106 , \35105 );
not \U$34730 ( \35107 , \34912 );
or \U$34731 ( \35108 , \35106 , \35107 );
not \U$34732 ( \35109 , \34898 );
nand \U$34733 ( \35110 , \35109 , \34908 );
nand \U$34734 ( \35111 , \35108 , \35110 );
xor \U$34735 ( \35112 , \35104 , \35111 );
xor \U$34736 ( \35113 , \34951 , \34955 );
and \U$34737 ( \35114 , \35113 , \34962 );
and \U$34738 ( \35115 , \34951 , \34955 );
or \U$34739 ( \35116 , \35114 , \35115 );
and \U$34740 ( \35117 , \35112 , \35116 );
and \U$34741 ( \35118 , \35104 , \35111 );
nor \U$34742 ( \35119 , \35117 , \35118 );
not \U$34743 ( \35120 , \35003 );
not \U$34744 ( \35121 , \35120 );
not \U$34745 ( \35122 , \35020 );
or \U$34746 ( \35123 , \35121 , \35122 );
or \U$34747 ( \35124 , \35020 , \35120 );
nand \U$34748 ( \35125 , \35124 , \35002 );
nand \U$34749 ( \35126 , \35123 , \35125 );
not \U$34750 ( \35127 , \35126 );
and \U$34751 ( \35128 , \19897 , \19904 );
not \U$34752 ( \35129 , \19897 );
and \U$34753 ( \35130 , \35129 , \19903 );
nor \U$34754 ( \35131 , \35128 , \35130 );
not \U$34755 ( \35132 , \35131 );
not \U$34756 ( \35133 , \19939 );
and \U$34757 ( \35134 , \35132 , \35133 );
and \U$34758 ( \35135 , \19939 , \35131 );
nor \U$34759 ( \35136 , \35134 , \35135 );
not \U$34760 ( \35137 , \35136 );
xor \U$34761 ( \35138 , \19721 , \19756 );
xor \U$34762 ( \35139 , \35138 , \19789 );
not \U$34763 ( \35140 , \35139 );
or \U$34764 ( \35141 , \35137 , \35140 );
or \U$34765 ( \35142 , \35139 , \35136 );
nand \U$34766 ( \35143 , \35141 , \35142 );
not \U$34767 ( \35144 , \35143 );
or \U$34768 ( \35145 , \35127 , \35144 );
not \U$34769 ( \35146 , \35136 );
nand \U$34770 ( \35147 , \35146 , \35139 );
nand \U$34771 ( \35148 , \35145 , \35147 );
not \U$34772 ( \35149 , \35148 );
and \U$34773 ( \35150 , \35119 , \35149 );
not \U$34774 ( \35151 , \35119 );
and \U$34775 ( \35152 , \35151 , \35148 );
nor \U$34776 ( \35153 , \35150 , \35152 );
not \U$34777 ( \35154 , \35036 );
not \U$34778 ( \35155 , \35045 );
nand \U$34779 ( \35156 , \35155 , \35031 );
not \U$34780 ( \35157 , \35156 );
or \U$34781 ( \35158 , \35154 , \35157 );
not \U$34782 ( \35159 , \35031 );
nand \U$34783 ( \35160 , \35159 , \35045 );
nand \U$34784 ( \35161 , \35158 , \35160 );
not \U$34785 ( \35162 , \35161 );
xor \U$34786 ( \35163 , \34801 , \34803 );
and \U$34787 ( \35164 , \35163 , \34821 );
and \U$34788 ( \35165 , \34801 , \34803 );
or \U$34789 ( \35166 , \35164 , \35165 );
xor \U$34790 ( \35167 , \19635 , \19632 );
xor \U$34791 ( \35168 , \35167 , \19639 );
xor \U$34792 ( \35169 , \35166 , \35168 );
not \U$34793 ( \35170 , \35169 );
or \U$34794 ( \35171 , \35162 , \35170 );
nand \U$34795 ( \35172 , \35168 , \35166 );
nand \U$34796 ( \35173 , \35171 , \35172 );
xor \U$34797 ( \35174 , \35153 , \35173 );
xor \U$34798 ( \35175 , \35116 , \35112 );
not \U$34799 ( \35176 , \34963 );
not \U$34800 ( \35177 , \34559 );
not \U$34801 ( \35178 , \34541 );
or \U$34802 ( \35179 , \35177 , \35178 );
nand \U$34803 ( \35180 , \35179 , \34933 );
not \U$34804 ( \35181 , \35180 );
not \U$34805 ( \35182 , \35181 );
not \U$34806 ( \35183 , \34944 );
or \U$34807 ( \35184 , \35182 , \35183 );
or \U$34808 ( \35185 , \34944 , \35181 );
nand \U$34809 ( \35186 , \35184 , \35185 );
not \U$34810 ( \35187 , \35186 );
or \U$34811 ( \35188 , \35176 , \35187 );
nand \U$34812 ( \35189 , \34944 , \35180 );
nand \U$34813 ( \35190 , \35188 , \35189 );
xor \U$34814 ( \35191 , \35175 , \35190 );
xor \U$34815 ( \35192 , \35161 , \35169 );
and \U$34816 ( \35193 , \35191 , \35192 );
and \U$34817 ( \35194 , \35175 , \35190 );
or \U$34818 ( \35195 , \35193 , \35194 );
and \U$34819 ( \35196 , \35174 , \35195 );
not \U$34820 ( \35197 , \35174 );
not \U$34821 ( \35198 , \35195 );
and \U$34822 ( \35199 , \35197 , \35198 );
nor \U$34823 ( \35200 , \35196 , \35199 );
not \U$34824 ( \35201 , \19654 );
not \U$34825 ( \35202 , \19793 );
and \U$34826 ( \35203 , \35201 , \35202 );
and \U$34827 ( \35204 , \19654 , \19793 );
nor \U$34828 ( \35205 , \35203 , \35204 );
not \U$34829 ( \35206 , \35205 );
not \U$34830 ( \35207 , \19647 );
and \U$34831 ( \35208 , \35206 , \35207 );
and \U$34832 ( \35209 , \19647 , \35205 );
nor \U$34833 ( \35210 , \35208 , \35209 );
xor \U$34834 ( \35211 , \19354 , \19384 );
xor \U$34835 ( \35212 , \35211 , \19412 );
xor \U$34836 ( \35213 , \19417 , \19452 );
xor \U$34837 ( \35214 , \35213 , \19488 );
xor \U$34838 ( \35215 , \35212 , \35214 );
and \U$34839 ( \35216 , \19148 , \19119 );
not \U$34840 ( \35217 , \19148 );
not \U$34841 ( \35218 , \19119 );
and \U$34842 ( \35219 , \35217 , \35218 );
nor \U$34843 ( \35220 , \35216 , \35219 );
not \U$34844 ( \35221 , \35220 );
not \U$34845 ( \35222 , \34809 );
not \U$34846 ( \35223 , \34819 );
or \U$34847 ( \35224 , \35222 , \35223 );
nand \U$34848 ( \35225 , \34814 , \34818 );
nand \U$34849 ( \35226 , \35224 , \35225 );
not \U$34850 ( \35227 , \35226 );
xor \U$34851 ( \35228 , \19387 , \19396 );
xor \U$34852 ( \35229 , \35228 , \19409 );
xnor \U$34853 ( \35230 , \35227 , \35229 );
not \U$34854 ( \35231 , \35230 );
or \U$34855 ( \35232 , \35221 , \35231 );
not \U$34856 ( \35233 , \35227 );
nand \U$34857 ( \35234 , \35233 , \35229 );
nand \U$34858 ( \35235 , \35232 , \35234 );
xor \U$34859 ( \35236 , \35215 , \35235 );
xor \U$34860 ( \35237 , \35210 , \35236 );
not \U$34861 ( \35238 , \19948 );
not \U$34862 ( \35239 , \19946 );
and \U$34863 ( \35240 , \35238 , \35239 );
and \U$34864 ( \35241 , \19948 , \19946 );
nor \U$34865 ( \35242 , \35240 , \35241 );
xnor \U$34866 ( \35243 , \35237 , \35242 );
and \U$34867 ( \35244 , \35200 , \35243 );
not \U$34868 ( \35245 , \35200 );
not \U$34869 ( \35246 , \35243 );
and \U$34870 ( \35247 , \35245 , \35246 );
nor \U$34871 ( \35248 , \35244 , \35247 );
not \U$34872 ( \35249 , \34854 );
not \U$34873 ( \35250 , \34969 );
or \U$34874 ( \35251 , \35249 , \35250 );
nand \U$34875 ( \35252 , \35251 , \34981 );
nand \U$34876 ( \35253 , \34970 , \34853 );
nand \U$34877 ( \35254 , \35252 , \35253 );
not \U$34878 ( \35255 , \35254 );
not \U$34879 ( \35256 , \35047 );
nand \U$34880 ( \35257 , \35256 , \35057 );
not \U$34881 ( \35258 , \35257 );
not \U$34882 ( \35259 , \35070 );
or \U$34883 ( \35260 , \35258 , \35259 );
not \U$34884 ( \35261 , \35057 );
nand \U$34885 ( \35262 , \35261 , \35047 );
nand \U$34886 ( \35263 , \35260 , \35262 );
not \U$34887 ( \35264 , \35263 );
not \U$34888 ( \35265 , \34848 );
not \U$34889 ( \35266 , \34842 );
or \U$34890 ( \35267 , \35265 , \35266 );
nand \U$34891 ( \35268 , \34841 , \34822 );
nand \U$34892 ( \35269 , \35267 , \35268 );
xor \U$34893 ( \35270 , \35220 , \35227 );
xnor \U$34894 ( \35271 , \35270 , \35229 );
not \U$34895 ( \35272 , \19851 );
and \U$34896 ( \35273 , \19890 , \35272 );
not \U$34897 ( \35274 , \19890 );
and \U$34898 ( \35275 , \35274 , \19851 );
nor \U$34899 ( \35276 , \35273 , \35275 );
not \U$34900 ( \35277 , \35276 );
xor \U$34901 ( \35278 , \19464 , \19484 );
not \U$34902 ( \35279 , \35278 );
xor \U$34903 ( \35280 , \19364 , \19370 );
xor \U$34904 ( \35281 , \35280 , \19381 );
not \U$34905 ( \35282 , \35281 );
nand \U$34906 ( \35283 , \35279 , \35282 );
nand \U$34907 ( \35284 , \35281 , \35278 );
nand \U$34908 ( \35285 , \35283 , \35284 );
not \U$34909 ( \35286 , \34896 );
not \U$34910 ( \35287 , \34886 );
or \U$34911 ( \35288 , \35286 , \35287 );
not \U$34912 ( \35289 , \34874 );
nand \U$34913 ( \35290 , \35289 , \34882 );
nand \U$34914 ( \35291 , \35288 , \35290 );
not \U$34915 ( \35292 , \35291 );
and \U$34916 ( \35293 , \35285 , \35292 );
not \U$34917 ( \35294 , \35285 );
and \U$34918 ( \35295 , \35294 , \35291 );
nor \U$34919 ( \35296 , \35293 , \35295 );
not \U$34920 ( \35297 , \35296 );
or \U$34921 ( \35298 , \35277 , \35297 );
or \U$34922 ( \35299 , \35276 , \35296 );
nand \U$34923 ( \35300 , \35298 , \35299 );
xor \U$34924 ( \35301 , \35271 , \35300 );
not \U$34925 ( \35302 , \35301 );
xor \U$34926 ( \35303 , \35024 , \35029 );
and \U$34927 ( \35304 , \35303 , \35046 );
and \U$34928 ( \35305 , \35024 , \35029 );
or \U$34929 ( \35306 , \35304 , \35305 );
not \U$34930 ( \35307 , \35306 );
and \U$34931 ( \35308 , \35302 , \35307 );
and \U$34932 ( \35309 , \35301 , \35306 );
nor \U$34933 ( \35310 , \35308 , \35309 );
xnor \U$34934 ( \35311 , \35269 , \35310 );
not \U$34935 ( \35312 , \35311 );
or \U$34936 ( \35313 , \35264 , \35312 );
or \U$34937 ( \35314 , \35311 , \35263 );
nand \U$34938 ( \35315 , \35313 , \35314 );
not \U$34939 ( \35316 , \35315 );
or \U$34940 ( \35317 , \35255 , \35316 );
not \U$34941 ( \35318 , \35311 );
nand \U$34942 ( \35319 , \35318 , \35263 );
nand \U$34943 ( \35320 , \35317 , \35319 );
not \U$34944 ( \35321 , \35320 );
xor \U$34945 ( \35322 , \35248 , \35321 );
not \U$34946 ( \35323 , \35126 );
and \U$34947 ( \35324 , \35143 , \35323 );
not \U$34948 ( \35325 , \35143 );
and \U$34949 ( \35326 , \35325 , \35126 );
or \U$34950 ( \35327 , \35324 , \35326 );
not \U$34951 ( \35328 , \35327 );
not \U$34952 ( \35329 , \34868 );
not \U$34953 ( \35330 , \34926 );
or \U$34954 ( \35331 , \35329 , \35330 );
not \U$34955 ( \35332 , \34923 );
nand \U$34956 ( \35333 , \35332 , \34897 );
nand \U$34957 ( \35334 , \35331 , \35333 );
not \U$34958 ( \35335 , \35334 );
nand \U$34959 ( \35336 , \35328 , \35335 );
not \U$34960 ( \35337 , \35336 );
xnor \U$34961 ( \35338 , \34826 , \34831 );
or \U$34962 ( \35339 , \35338 , \34839 );
nand \U$34963 ( \35340 , \34831 , \34826 );
nand \U$34964 ( \35341 , \35339 , \35340 );
not \U$34965 ( \35342 , \35341 );
or \U$34966 ( \35343 , \35337 , \35342 );
nand \U$34967 ( \35344 , \35334 , \35327 );
nand \U$34968 ( \35345 , \35343 , \35344 );
not \U$34969 ( \35346 , \35345 );
buf \U$34970 ( \35347 , \35296 );
or \U$34971 ( \35348 , \35271 , \35347 );
not \U$34972 ( \35349 , \35276 );
nand \U$34973 ( \35350 , \35348 , \35349 );
nand \U$34974 ( \35351 , \35347 , \35271 );
nand \U$34975 ( \35352 , \35350 , \35351 );
not \U$34976 ( \35353 , \35352 );
not \U$34977 ( \35354 , \35291 );
not \U$34978 ( \35355 , \35283 );
or \U$34979 ( \35356 , \35354 , \35355 );
nand \U$34980 ( \35357 , \35356 , \35284 );
not \U$34981 ( \35358 , \19587 );
not \U$34982 ( \35359 , \19584 );
not \U$34983 ( \35360 , \35359 );
or \U$34984 ( \35361 , \35358 , \35360 );
nand \U$34985 ( \35362 , \19584 , \19586 );
nand \U$34986 ( \35363 , \35361 , \35362 );
xor \U$34987 ( \35364 , \35357 , \35363 );
xor \U$34988 ( \35365 , \19074 , \18947 );
xnor \U$34989 ( \35366 , \35365 , \19080 );
xnor \U$34990 ( \35367 , \35364 , \35366 );
not \U$34991 ( \35368 , \35367 );
or \U$34992 ( \35369 , \35353 , \35368 );
or \U$34993 ( \35370 , \35367 , \35352 );
nand \U$34994 ( \35371 , \35369 , \35370 );
not \U$34995 ( \35372 , \35371 );
not \U$34996 ( \35373 , \35372 );
or \U$34997 ( \35374 , \35346 , \35373 );
not \U$34998 ( \35375 , \35345 );
nand \U$34999 ( \35376 , \35371 , \35375 );
nand \U$35000 ( \35377 , \35374 , \35376 );
not \U$35001 ( \35378 , \35377 );
not \U$35002 ( \35379 , \35301 );
nand \U$35003 ( \35380 , \35379 , \35306 );
not \U$35004 ( \35381 , \35380 );
not \U$35005 ( \35382 , \35269 );
or \U$35006 ( \35383 , \35381 , \35382 );
not \U$35007 ( \35384 , \35306 );
nand \U$35008 ( \35385 , \35384 , \35301 );
nand \U$35009 ( \35386 , \35383 , \35385 );
not \U$35010 ( \35387 , \35386 );
nand \U$35011 ( \35388 , \35378 , \35387 );
nand \U$35012 ( \35389 , \35377 , \35386 );
nand \U$35013 ( \35390 , \35388 , \35389 );
not \U$35014 ( \35391 , \34964 );
not \U$35015 ( \35392 , \34928 );
or \U$35016 ( \35393 , \35391 , \35392 );
nand \U$35017 ( \35394 , \34927 , \34864 );
nand \U$35018 ( \35395 , \35393 , \35394 );
not \U$35019 ( \35396 , \35395 );
xor \U$35020 ( \35397 , \35327 , \35335 );
xor \U$35021 ( \35398 , \35397 , \35341 );
not \U$35022 ( \35399 , \35398 );
not \U$35023 ( \35400 , \35399 );
or \U$35024 ( \35401 , \35396 , \35400 );
not \U$35025 ( \35402 , \35398 );
not \U$35026 ( \35403 , \35395 );
not \U$35027 ( \35404 , \35403 );
or \U$35028 ( \35405 , \35402 , \35404 );
xor \U$35029 ( \35406 , \35175 , \35190 );
xor \U$35030 ( \35407 , \35406 , \35192 );
nand \U$35031 ( \35408 , \35405 , \35407 );
nand \U$35032 ( \35409 , \35401 , \35408 );
and \U$35033 ( \35410 , \35390 , \35409 );
not \U$35034 ( \35411 , \35390 );
not \U$35035 ( \35412 , \35409 );
and \U$35036 ( \35413 , \35411 , \35412 );
nor \U$35037 ( \35414 , \35410 , \35413 );
xnor \U$35038 ( \35415 , \35322 , \35414 );
xor \U$35039 ( \35416 , \35254 , \35315 );
not \U$35040 ( \35417 , \35416 );
not \U$35041 ( \35418 , \34999 );
and \U$35042 ( \35419 , \35081 , \35076 );
not \U$35043 ( \35420 , \35419 );
and \U$35044 ( \35421 , \35418 , \35420 );
nor \U$35045 ( \35422 , \35081 , \35076 );
nor \U$35046 ( \35423 , \35421 , \35422 );
not \U$35047 ( \35424 , \35399 );
not \U$35048 ( \35425 , \35403 );
or \U$35049 ( \35426 , \35424 , \35425 );
nand \U$35050 ( \35427 , \35395 , \35398 );
nand \U$35051 ( \35428 , \35426 , \35427 );
not \U$35052 ( \35429 , \35407 );
and \U$35053 ( \35430 , \35428 , \35429 );
not \U$35054 ( \35431 , \35428 );
and \U$35055 ( \35432 , \35431 , \35407 );
nor \U$35056 ( \35433 , \35430 , \35432 );
not \U$35057 ( \35434 , \35433 );
and \U$35058 ( \35435 , \35423 , \35434 );
not \U$35059 ( \35436 , \35423 );
and \U$35060 ( \35437 , \35436 , \35433 );
nor \U$35061 ( \35438 , \35435 , \35437 );
not \U$35062 ( \35439 , \35438 );
or \U$35063 ( \35440 , \35417 , \35439 );
not \U$35064 ( \35441 , \35423 );
nand \U$35065 ( \35442 , \35441 , \35433 );
nand \U$35066 ( \35443 , \35440 , \35442 );
nand \U$35067 ( \35444 , \35415 , \35443 );
xor \U$35068 ( \35445 , \35416 , \35438 );
xor \U$35069 ( \35446 , \34985 , \34992 );
and \U$35070 ( \35447 , \35446 , \35089 );
and \U$35071 ( \35448 , \34985 , \34992 );
or \U$35072 ( \35449 , \35447 , \35448 );
nand \U$35073 ( \35450 , \35445 , \35449 );
nand \U$35074 ( \35451 , \35103 , \35444 , \35450 );
not \U$35075 ( \35452 , \35451 );
nand \U$35076 ( \35453 , \34369 , \35452 );
not \U$35077 ( \35454 , \35453 );
buf \U$35078 ( \35455 , \34795 );
not \U$35079 ( \35456 , \35455 );
not \U$35080 ( \35457 , \35090 );
not \U$35081 ( \35458 , \35457 );
or \U$35082 ( \35459 , \35456 , \35458 );
not \U$35083 ( \35460 , \35101 );
nand \U$35084 ( \35461 , \35460 , \35095 );
nand \U$35085 ( \35462 , \35459 , \35461 );
and \U$35086 ( \35463 , \35444 , \35462 , \35450 );
buf \U$35087 ( \35464 , \35091 );
and \U$35088 ( \35465 , \35463 , \35464 );
not \U$35089 ( \35466 , \35444 );
not \U$35090 ( \35467 , \35445 );
not \U$35091 ( \35468 , \35449 );
nand \U$35092 ( \35469 , \35467 , \35468 );
or \U$35093 ( \35470 , \35466 , \35469 );
nor \U$35094 ( \35471 , \35415 , \35443 );
not \U$35095 ( \35472 , \35471 );
nand \U$35096 ( \35473 , \35470 , \35472 );
nor \U$35097 ( \35474 , \35465 , \35473 );
not \U$35098 ( \35475 , \35474 );
or \U$35099 ( \35476 , \35454 , \35475 );
xor \U$35100 ( \35477 , \19957 , \19963 );
xor \U$35101 ( \35478 , \35477 , \19965 );
not \U$35102 ( \35479 , \35478 );
xor \U$35103 ( \35480 , \19167 , \19164 );
xor \U$35104 ( \35481 , \35480 , \19170 );
xor \U$35105 ( \35482 , \35212 , \35214 );
and \U$35106 ( \35483 , \35482 , \35235 );
and \U$35107 ( \35484 , \35212 , \35214 );
or \U$35108 ( \35485 , \35483 , \35484 );
or \U$35109 ( \35486 , \35481 , \35485 );
not \U$35110 ( \35487 , \35366 );
not \U$35111 ( \35488 , \35364 );
or \U$35112 ( \35489 , \35487 , \35488 );
nand \U$35113 ( \35490 , \35363 , \35357 );
nand \U$35114 ( \35491 , \35489 , \35490 );
nand \U$35115 ( \35492 , \35486 , \35491 );
nand \U$35116 ( \35493 , \35481 , \35485 );
nand \U$35117 ( \35494 , \35492 , \35493 );
not \U$35118 ( \35495 , \35494 );
not \U$35119 ( \35496 , \35495 );
xor \U$35120 ( \35497 , \19181 , \19104 );
xor \U$35121 ( \35498 , \35497 , \19179 );
not \U$35122 ( \35499 , \35498 );
or \U$35123 ( \35500 , \35496 , \35499 );
xor \U$35124 ( \35501 , \19521 , \19523 );
xor \U$35125 ( \35502 , \35501 , \19526 );
not \U$35126 ( \35503 , \35502 );
not \U$35127 ( \35504 , \35498 );
nand \U$35128 ( \35505 , \35504 , \35494 );
nand \U$35129 ( \35506 , \35503 , \35505 );
nand \U$35130 ( \35507 , \35500 , \35506 );
not \U$35131 ( \35508 , \35507 );
not \U$35132 ( \35509 , \35508 );
not \U$35133 ( \35510 , \35498 );
and \U$35134 ( \35511 , \35502 , \35494 );
not \U$35135 ( \35512 , \35502 );
and \U$35136 ( \35513 , \35512 , \35495 );
nor \U$35137 ( \35514 , \35511 , \35513 );
not \U$35138 ( \35515 , \35514 );
or \U$35139 ( \35516 , \35510 , \35515 );
or \U$35140 ( \35517 , \35514 , \35498 );
nand \U$35141 ( \35518 , \35516 , \35517 );
not \U$35142 ( \35519 , \35153 );
not \U$35143 ( \35520 , \35173 );
or \U$35144 ( \35521 , \35519 , \35520 );
not \U$35145 ( \35522 , \35119 );
nand \U$35146 ( \35523 , \35522 , \35148 );
nand \U$35147 ( \35524 , \35521 , \35523 );
not \U$35148 ( \35525 , \35524 );
xnor \U$35149 ( \35526 , \19099 , \19089 );
not \U$35150 ( \35527 , \35526 );
not \U$35151 ( \35528 , \35527 );
xor \U$35152 ( \35529 , \19597 , \19798 );
not \U$35153 ( \35530 , \35529 );
not \U$35154 ( \35531 , \35530 );
or \U$35155 ( \35532 , \35528 , \35531 );
nand \U$35156 ( \35533 , \35529 , \35526 );
nand \U$35157 ( \35534 , \35532 , \35533 );
not \U$35158 ( \35535 , \35534 );
or \U$35159 ( \35536 , \35525 , \35535 );
nand \U$35160 ( \35537 , \35529 , \35527 );
nand \U$35161 ( \35538 , \35536 , \35537 );
not \U$35162 ( \35539 , \35538 );
xor \U$35163 ( \35540 , \19803 , \19805 );
xor \U$35164 ( \35541 , \35540 , \19954 );
not \U$35165 ( \35542 , \35541 );
nand \U$35166 ( \35543 , \35539 , \35542 );
nand \U$35167 ( \35544 , \35518 , \35543 );
nand \U$35168 ( \35545 , \35538 , \35541 );
and \U$35169 ( \35546 , \35544 , \35545 );
not \U$35170 ( \35547 , \35546 );
or \U$35171 ( \35548 , \35509 , \35547 );
not \U$35172 ( \35549 , \35545 );
not \U$35173 ( \35550 , \35544 );
or \U$35174 ( \35551 , \35549 , \35550 );
nand \U$35175 ( \35552 , \35551 , \35507 );
nand \U$35176 ( \35553 , \35548 , \35552 );
not \U$35177 ( \35554 , \35553 );
or \U$35178 ( \35555 , \35479 , \35554 );
or \U$35179 ( \35556 , \35553 , \35478 );
nand \U$35180 ( \35557 , \35555 , \35556 );
nand \U$35181 ( \35558 , \19811 , \19953 );
xor \U$35182 ( \35559 , \19950 , \35558 );
xor \U$35183 ( \35560 , \35491 , \35485 );
xnor \U$35184 ( \35561 , \35560 , \35481 );
xor \U$35185 ( \35562 , \35559 , \35561 );
not \U$35186 ( \35563 , \35242 );
not \U$35187 ( \35564 , \35210 );
and \U$35188 ( \35565 , \35563 , \35564 );
xor \U$35189 ( \35566 , \35210 , \35242 );
and \U$35190 ( \35567 , \35566 , \35236 );
nor \U$35191 ( \35568 , \35565 , \35567 );
and \U$35192 ( \35569 , \35562 , \35568 );
and \U$35193 ( \35570 , \35559 , \35561 );
or \U$35194 ( \35571 , \35569 , \35570 );
not \U$35195 ( \35572 , \35524 );
and \U$35196 ( \35573 , \35534 , \35572 );
not \U$35197 ( \35574 , \35534 );
and \U$35198 ( \35575 , \35574 , \35524 );
or \U$35199 ( \35576 , \35573 , \35575 );
not \U$35200 ( \35577 , \35576 );
not \U$35201 ( \35578 , \35345 );
not \U$35202 ( \35579 , \35371 );
or \U$35203 ( \35580 , \35578 , \35579 );
not \U$35204 ( \35581 , \35367 );
nand \U$35205 ( \35582 , \35581 , \35352 );
nand \U$35206 ( \35583 , \35580 , \35582 );
not \U$35207 ( \35584 , \35583 );
or \U$35208 ( \35585 , \35577 , \35584 );
not \U$35209 ( \35586 , \35583 );
not \U$35210 ( \35587 , \35586 );
not \U$35211 ( \35588 , \35576 );
not \U$35212 ( \35589 , \35588 );
or \U$35213 ( \35590 , \35587 , \35589 );
not \U$35214 ( \35591 , \35174 );
not \U$35215 ( \35592 , \35591 );
not \U$35216 ( \35593 , \35592 );
not \U$35217 ( \35594 , \35246 );
or \U$35218 ( \35595 , \35593 , \35594 );
not \U$35219 ( \35596 , \35591 );
not \U$35220 ( \35597 , \35243 );
or \U$35221 ( \35598 , \35596 , \35597 );
not \U$35222 ( \35599 , \35198 );
nand \U$35223 ( \35600 , \35598 , \35599 );
nand \U$35224 ( \35601 , \35595 , \35600 );
nand \U$35225 ( \35602 , \35590 , \35601 );
nand \U$35226 ( \35603 , \35585 , \35602 );
not \U$35227 ( \35604 , \35603 );
xor \U$35228 ( \35605 , \35571 , \35604 );
not \U$35229 ( \35606 , \35542 );
not \U$35230 ( \35607 , \35539 );
or \U$35231 ( \35608 , \35606 , \35607 );
nand \U$35232 ( \35609 , \35608 , \35545 );
xor \U$35233 ( \35610 , \35609 , \35518 );
and \U$35234 ( \35611 , \35605 , \35610 );
and \U$35235 ( \35612 , \35571 , \35604 );
or \U$35236 ( \35613 , \35611 , \35612 );
nand \U$35237 ( \35614 , \35557 , \35613 );
not \U$35238 ( \35615 , \35320 );
xor \U$35239 ( \35616 , \35248 , \35414 );
not \U$35240 ( \35617 , \35616 );
or \U$35241 ( \35618 , \35615 , \35617 );
nand \U$35242 ( \35619 , \35414 , \35248 );
nand \U$35243 ( \35620 , \35618 , \35619 );
not \U$35244 ( \35621 , \35601 );
not \U$35245 ( \35622 , \35583 );
not \U$35246 ( \35623 , \35588 );
or \U$35247 ( \35624 , \35622 , \35623 );
nand \U$35248 ( \35625 , \35576 , \35586 );
nand \U$35249 ( \35626 , \35624 , \35625 );
not \U$35250 ( \35627 , \35626 );
or \U$35251 ( \35628 , \35621 , \35627 );
or \U$35252 ( \35629 , \35626 , \35601 );
nand \U$35253 ( \35630 , \35628 , \35629 );
not \U$35254 ( \35631 , \35388 );
not \U$35255 ( \35632 , \35409 );
or \U$35256 ( \35633 , \35631 , \35632 );
nand \U$35257 ( \35634 , \35633 , \35389 );
not \U$35258 ( \35635 , \35634 );
xor \U$35259 ( \35636 , \35559 , \35561 );
xor \U$35260 ( \35637 , \35636 , \35568 );
not \U$35261 ( \35638 , \35637 );
or \U$35262 ( \35639 , \35635 , \35638 );
or \U$35263 ( \35640 , \35637 , \35634 );
nand \U$35264 ( \35641 , \35639 , \35640 );
xor \U$35265 ( \35642 , \35630 , \35641 );
nand \U$35266 ( \35643 , \35620 , \35642 );
not \U$35267 ( \35644 , \35478 );
not \U$35268 ( \35645 , \35644 );
not \U$35269 ( \35646 , \35553 );
or \U$35270 ( \35647 , \35645 , \35646 );
nand \U$35271 ( \35648 , \35544 , \35507 , \35545 );
nand \U$35272 ( \35649 , \35647 , \35648 );
xor \U$35273 ( \35650 , \19563 , \19968 );
xnor \U$35274 ( \35651 , \35650 , \19560 );
nand \U$35275 ( \35652 , \35649 , \35651 );
xor \U$35276 ( \35653 , \35571 , \35604 );
xor \U$35277 ( \35654 , \35653 , \35610 );
not \U$35278 ( \35655 , \35630 );
not \U$35279 ( \35656 , \35641 );
or \U$35280 ( \35657 , \35655 , \35656 );
not \U$35281 ( \35658 , \35634 );
nand \U$35282 ( \35659 , \35658 , \35637 );
nand \U$35283 ( \35660 , \35657 , \35659 );
nand \U$35284 ( \35661 , \35654 , \35660 );
and \U$35285 ( \35662 , \35614 , \35643 , \35652 , \35661 );
nand \U$35286 ( \35663 , \35476 , \35662 );
xor \U$35287 ( \35664 , \33669 , \33730 );
xor \U$35288 ( \35665 , \35664 , \33765 );
xor \U$35289 ( \35666 , \33900 , \33926 );
not \U$35290 ( \35667 , \34000 );
not \U$35291 ( \35668 , \35667 );
not \U$35292 ( \35669 , \33990 );
or \U$35293 ( \35670 , \35668 , \35669 );
or \U$35294 ( \35671 , \33990 , \35667 );
nand \U$35295 ( \35672 , \35670 , \35671 );
xor \U$35296 ( \35673 , \35666 , \35672 );
not \U$35297 ( \35674 , \10275 );
not \U$35298 ( \35675 , \33953 );
or \U$35299 ( \35676 , \35674 , \35675 );
not \U$35300 ( \35677 , RIae7a8d0_188);
not \U$35301 ( \35678 , \1789 );
or \U$35302 ( \35679 , \35677 , \35678 );
or \U$35303 ( \35680 , \2577 , RIae7a8d0_188);
nand \U$35304 ( \35681 , \35679 , \35680 );
nand \U$35305 ( \35682 , \35681 , \11205 );
nand \U$35306 ( \35683 , \35676 , \35682 );
not \U$35307 ( \35684 , \35683 );
not \U$35308 ( \35685 , \10519 );
not \U$35309 ( \35686 , \33996 );
or \U$35310 ( \35687 , \35685 , \35686 );
xnor \U$35311 ( \35688 , \3216 , RIae7a7e0_186);
nand \U$35312 ( \35689 , \35688 , \11439 );
nand \U$35313 ( \35690 , \35687 , \35689 );
not \U$35314 ( \35691 , \11422 );
not \U$35315 ( \35692 , \33987 );
or \U$35316 ( \35693 , \35691 , \35692 );
xnor \U$35317 ( \35694 , RIae7a498_179, \13248 );
nand \U$35318 ( \35695 , \35694 , \15382 );
nand \U$35319 ( \35696 , \35693 , \35695 );
xor \U$35320 ( \35697 , \35690 , \35696 );
not \U$35321 ( \35698 , \35697 );
or \U$35322 ( \35699 , \35684 , \35698 );
nand \U$35323 ( \35700 , \35696 , \35690 );
nand \U$35324 ( \35701 , \35699 , \35700 );
and \U$35325 ( \35702 , \35673 , \35701 );
and \U$35326 ( \35703 , \35666 , \35672 );
or \U$35327 ( \35704 , \35702 , \35703 );
xor \U$35328 ( \35705 , \35665 , \35704 );
xnor \U$35329 ( \35706 , \33969 , \34013 );
and \U$35330 ( \35707 , \35705 , \35706 );
and \U$35331 ( \35708 , \35665 , \35704 );
or \U$35332 ( \35709 , \35707 , \35708 );
not \U$35333 ( \35710 , \35709 );
xnor \U$35334 ( \35711 , \33610 , \33611 );
not \U$35335 ( \35712 , \33781 );
not \U$35336 ( \35713 , \33778 );
not \U$35337 ( \35714 , \35713 );
or \U$35338 ( \35715 , \35712 , \35714 );
not \U$35339 ( \35716 , \33781 );
nand \U$35340 ( \35717 , \35716 , \33778 );
nand \U$35341 ( \35718 , \35715 , \35717 );
or \U$35342 ( \35719 , \35711 , \35718 );
nand \U$35343 ( \35720 , \35718 , \35711 );
nand \U$35344 ( \35721 , \35719 , \35720 );
not \U$35345 ( \35722 , \35721 );
or \U$35346 ( \35723 , \35710 , \35722 );
not \U$35347 ( \35724 , \35711 );
nand \U$35348 ( \35725 , \35724 , \35718 );
nand \U$35349 ( \35726 , \35723 , \35725 );
not \U$35350 ( \35727 , \35726 );
xor \U$35351 ( \35728 , \33786 , \33661 );
xnor \U$35352 ( \35729 , \35728 , \33668 );
not \U$35353 ( \35730 , \35729 );
not \U$35354 ( \35731 , \35730 );
or \U$35355 ( \35732 , \35727 , \35731 );
not \U$35356 ( \35733 , \35726 );
nand \U$35357 ( \35734 , \35729 , \35733 );
nand \U$35358 ( \35735 , \35732 , \35734 );
xor \U$35359 ( \35736 , \33800 , \33802 );
xor \U$35360 ( \35737 , \35736 , \33883 );
xor \U$35361 ( \35738 , \33678 , \33726 );
not \U$35362 ( \35739 , \17507 );
not \U$35363 ( \35740 , \33876 );
or \U$35364 ( \35741 , \35739 , \35740 );
and \U$35365 ( \35742 , RIae7a6f0_184, \13008 );
not \U$35366 ( \35743 , RIae7a6f0_184);
and \U$35367 ( \35744 , \35743 , \22917 );
or \U$35368 ( \35745 , \35742 , \35744 );
not \U$35369 ( \35746 , \9473 );
not \U$35370 ( \35747 , \35746 );
nand \U$35371 ( \35748 , \35745 , \35747 );
nand \U$35372 ( \35749 , \35741 , \35748 );
not \U$35373 ( \35750 , \35749 );
not \U$35374 ( \35751 , \10542 );
not \U$35375 ( \35752 , \33963 );
or \U$35376 ( \35753 , \35751 , \35752 );
and \U$35377 ( \35754 , RIae7a060_170, \2402 );
not \U$35378 ( \35755 , RIae7a060_170);
and \U$35379 ( \35756 , \35755 , \5673 );
or \U$35380 ( \35757 , \35754 , \35756 );
nand \U$35381 ( \35758 , \35757 , \9730 );
nand \U$35382 ( \35759 , \35753 , \35758 );
not \U$35383 ( \35760 , \35759 );
not \U$35384 ( \35761 , RIae7aab0_192);
not \U$35385 ( \35762 , \33867 );
or \U$35386 ( \35763 , \35761 , \35762 );
not \U$35387 ( \35764 , \14671 );
not \U$35388 ( \35765 , \1759 );
or \U$35389 ( \35766 , \35764 , \35765 );
or \U$35390 ( \35767 , \30416 , \14671 );
nand \U$35391 ( \35768 , \35766 , \35767 );
nand \U$35392 ( \35769 , \35768 , \16383 );
nand \U$35393 ( \35770 , \35763 , \35769 );
not \U$35394 ( \35771 , \35770 );
not \U$35395 ( \35772 , \35771 );
or \U$35396 ( \35773 , \35760 , \35772 );
or \U$35397 ( \35774 , \35771 , \35759 );
nand \U$35398 ( \35775 , \35773 , \35774 );
not \U$35399 ( \35776 , \35775 );
or \U$35400 ( \35777 , \35750 , \35776 );
not \U$35401 ( \35778 , \35771 );
nand \U$35402 ( \35779 , \35778 , \35759 );
nand \U$35403 ( \35780 , \35777 , \35779 );
xor \U$35404 ( \35781 , \35738 , \35780 );
buf \U$35405 ( \35782 , \35781 );
xor \U$35406 ( \35783 , \33880 , \33870 );
and \U$35407 ( \35784 , \35782 , \35783 );
and \U$35408 ( \35785 , \35738 , \35780 );
nor \U$35409 ( \35786 , \35784 , \35785 );
xor \U$35410 ( \35787 , \33930 , \33939 );
xor \U$35411 ( \35788 , \35787 , \33890 );
or \U$35412 ( \35789 , \35786 , \35788 );
and \U$35413 ( \35790 , \35737 , \35789 );
and \U$35414 ( \35791 , \35788 , \35786 );
nor \U$35415 ( \35792 , \35790 , \35791 );
xor \U$35416 ( \35793 , \34047 , \34272 );
xor \U$35417 ( \35794 , \35792 , \35793 );
xor \U$35418 ( \35795 , \33942 , \33886 );
xnor \U$35419 ( \35796 , \35795 , \34020 );
and \U$35420 ( \35797 , \35794 , \35796 );
and \U$35421 ( \35798 , \35792 , \35793 );
or \U$35422 ( \35799 , \35797 , \35798 );
xnor \U$35423 ( \35800 , \35735 , \35799 );
not \U$35424 ( \35801 , \35800 );
xor \U$35425 ( \35802 , \34277 , \34283 );
xnor \U$35426 ( \35803 , \35802 , \34028 );
not \U$35427 ( \35804 , \35803 );
not \U$35428 ( \35805 , \33812 );
not \U$35429 ( \35806 , \35805 );
not \U$35430 ( \35807 , \33829 );
or \U$35431 ( \35808 , \35806 , \35807 );
or \U$35432 ( \35809 , \33829 , \35805 );
nand \U$35433 ( \35810 , \35808 , \35809 );
not \U$35434 ( \35811 , \2417 );
and \U$35435 ( \35812 , \10740 , \10584 );
not \U$35436 ( \35813 , \10740 );
and \U$35437 ( \35814 , \35813 , RIae79c28_161);
nor \U$35438 ( \35815 , \35812 , \35814 );
not \U$35439 ( \35816 , \35815 );
or \U$35440 ( \35817 , \35811 , \35816 );
nand \U$35441 ( \35818 , \34224 , \2418 );
nand \U$35442 ( \35819 , \35817 , \35818 );
nand \U$35443 ( \35820 , \35810 , \35819 );
not \U$35444 ( \35821 , \35820 );
not \U$35445 ( \35822 , \35819 );
and \U$35446 ( \35823 , \35810 , \35822 );
not \U$35447 ( \35824 , \35810 );
and \U$35448 ( \35825 , \35824 , \35819 );
nor \U$35449 ( \35826 , \35823 , \35825 );
not \U$35450 ( \35827 , \35826 );
not \U$35451 ( \35828 , \19362 );
not \U$35452 ( \35829 , RIae79ef8_167);
not \U$35453 ( \35830 , \19015 );
or \U$35454 ( \35831 , \35829 , \35830 );
not \U$35455 ( \35832 , \10728 );
or \U$35456 ( \35833 , \35832 , RIae79ef8_167);
nand \U$35457 ( \35834 , \35831 , \35833 );
not \U$35458 ( \35835 , \35834 );
or \U$35459 ( \35836 , \35828 , \35835 );
nand \U$35460 ( \35837 , \34055 , \10573 );
nand \U$35461 ( \35838 , \35836 , \35837 );
nand \U$35462 ( \35839 , \35827 , \35838 );
not \U$35463 ( \35840 , \35839 );
or \U$35464 ( \35841 , \35821 , \35840 );
xor \U$35465 ( \35842 , \34217 , \34226 );
xor \U$35466 ( \35843 , \35842 , \34238 );
nand \U$35467 ( \35844 , \35841 , \35843 );
not \U$35468 ( \35845 , \35844 );
xnor \U$35469 ( \35846 , \33855 , \33844 );
not \U$35470 ( \35847 , \35846 );
or \U$35471 ( \35848 , \35845 , \35847 );
not \U$35472 ( \35849 , \35843 );
nand \U$35473 ( \35850 , \35849 , \35839 , \35820 );
nand \U$35474 ( \35851 , \35848 , \35850 );
not \U$35475 ( \35852 , \35851 );
xor \U$35476 ( \35853 , \33948 , \33965 );
xnor \U$35477 ( \35854 , \35853 , \33957 );
xor \U$35478 ( \35855 , \35852 , \35854 );
not \U$35479 ( \35856 , \5039 );
not \U$35480 ( \35857 , \4968 );
not \U$35481 ( \35858 , \10070 );
or \U$35482 ( \35859 , \35857 , \35858 );
or \U$35483 ( \35860 , \10072 , \4968 );
nand \U$35484 ( \35861 , \35859 , \35860 );
not \U$35485 ( \35862 , \35861 );
or \U$35486 ( \35863 , \35856 , \35862 );
nand \U$35487 ( \35864 , \33853 , \5048 );
nand \U$35488 ( \35865 , \35863 , \35864 );
not \U$35489 ( \35866 , \35865 );
not \U$35490 ( \35867 , \4154 );
not \U$35491 ( \35868 , \9875 );
xor \U$35492 ( \35869 , RIae79ca0_162, \35868 );
not \U$35493 ( \35870 , \35869 );
or \U$35494 ( \35871 , \35867 , \35870 );
nand \U$35495 ( \35872 , \34236 , \4853 );
nand \U$35496 ( \35873 , \35871 , \35872 );
and \U$35497 ( \35874 , \35866 , \35873 );
not \U$35498 ( \35875 , \35866 );
not \U$35499 ( \35876 , \35873 );
and \U$35500 ( \35877 , \35875 , \35876 );
nor \U$35501 ( \35878 , \35874 , \35877 );
not \U$35502 ( \35879 , \35878 );
not \U$35503 ( \35880 , \10638 );
not \U$35504 ( \35881 , RIae7a510_180);
not \U$35505 ( \35882 , \17242 );
or \U$35506 ( \35883 , \35881 , \35882 );
or \U$35507 ( \35884 , \22356 , RIae7a510_180);
nand \U$35508 ( \35885 , \35883 , \35884 );
not \U$35509 ( \35886 , \35885 );
or \U$35510 ( \35887 , \35880 , \35886 );
nand \U$35511 ( \35888 , \34201 , \16358 );
nand \U$35512 ( \35889 , \35887 , \35888 );
nand \U$35513 ( \35890 , \35879 , \35889 );
nand \U$35514 ( \35891 , \35865 , \35873 );
and \U$35515 ( \35892 , \35890 , \35891 );
not \U$35516 ( \35893 , \35892 );
not \U$35517 ( \35894 , \9644 );
not \U$35518 ( \35895 , \13165 );
not \U$35519 ( \35896 , \21744 );
or \U$35520 ( \35897 , \35895 , \35896 );
nand \U$35521 ( \35898 , \21747 , RIae7a3a8_177);
nand \U$35522 ( \35899 , \35897 , \35898 );
nor \U$35523 ( \35900 , \35894 , \35899 );
and \U$35524 ( \35901 , \34183 , \9622 );
nor \U$35525 ( \35902 , \35900 , \35901 );
not \U$35526 ( \35903 , \35902 );
not \U$35527 ( \35904 , \9792 );
xor \U$35528 ( \35905 , RIae7a2b8_175, \9395 );
not \U$35529 ( \35906 , \35905 );
or \U$35530 ( \35907 , \35904 , \35906 );
nand \U$35531 ( \35908 , \34143 , \9814 );
nand \U$35532 ( \35909 , \35907 , \35908 );
not \U$35533 ( \35910 , \35909 );
not \U$35534 ( \35911 , \19623 );
not \U$35535 ( \35912 , \9438 );
or \U$35536 ( \35913 , \35911 , \35912 );
not \U$35537 ( \35914 , \14110 );
nand \U$35538 ( \35915 , \35914 , RIae7a240_174);
nand \U$35539 ( \35916 , \35913 , \35915 );
and \U$35540 ( \35917 , \9688 , \35916 );
and \U$35541 ( \35918 , \34157 , \9699 );
nor \U$35542 ( \35919 , \35917 , \35918 );
not \U$35543 ( \35920 , \35919 );
or \U$35544 ( \35921 , \35910 , \35920 );
or \U$35545 ( \35922 , \35919 , \35909 );
nand \U$35546 ( \35923 , \35921 , \35922 );
not \U$35547 ( \35924 , \35923 );
or \U$35548 ( \35925 , \35903 , \35924 );
not \U$35549 ( \35926 , \35909 );
nand \U$35550 ( \35927 , \35926 , \35919 );
nand \U$35551 ( \35928 , \35925 , \35927 );
not \U$35552 ( \35929 , \35928 );
or \U$35553 ( \35930 , \35893 , \35929 );
not \U$35554 ( \35931 , \10709 );
and \U$35555 ( \35932 , \14148 , RIae79fe8_169);
not \U$35556 ( \35933 , \14148 );
and \U$35557 ( \35934 , \35933 , \9504 );
nor \U$35558 ( \35935 , \35932 , \35934 );
not \U$35559 ( \35936 , \35935 );
or \U$35560 ( \35937 , \35931 , \35936 );
not \U$35561 ( \35938 , \34132 );
nand \U$35562 ( \35939 , \35938 , \9518 );
nand \U$35563 ( \35940 , \35937 , \35939 );
not \U$35564 ( \35941 , \35940 );
not \U$35565 ( \35942 , \2007 );
not \U$35566 ( \35943 , \34091 );
or \U$35567 ( \35944 , \35942 , \35943 );
and \U$35568 ( \35945 , RIae797f0_152, \32808 );
not \U$35569 ( \35946 , RIae797f0_152);
and \U$35570 ( \35947 , \35946 , \11318 );
or \U$35571 ( \35948 , \35945 , \35947 );
nand \U$35572 ( \35949 , \35948 , \1988 );
nand \U$35573 ( \35950 , \35944 , \35949 );
not \U$35574 ( \35951 , \35950 );
not \U$35575 ( \35952 , \34072 );
not \U$35576 ( \35953 , \34082 );
or \U$35577 ( \35954 , \35952 , \35953 );
or \U$35578 ( \35955 , \34082 , \34072 );
nand \U$35579 ( \35956 , \35954 , \35955 );
not \U$35580 ( \35957 , \2321 );
not \U$35581 ( \35958 , \33810 );
or \U$35582 ( \35959 , \35957 , \35958 );
and \U$35583 ( \35960 , \16166 , \2981 );
not \U$35584 ( \35961 , \16166 );
and \U$35585 ( \35962 , \35961 , RIae798e0_154);
nor \U$35586 ( \35963 , \35960 , \35962 );
nand \U$35587 ( \35964 , \35963 , \2338 );
nand \U$35588 ( \35965 , \35959 , \35964 );
xor \U$35589 ( \35966 , \35956 , \35965 );
not \U$35590 ( \35967 , \35966 );
or \U$35591 ( \35968 , \35951 , \35967 );
nand \U$35592 ( \35969 , \35965 , \35956 );
nand \U$35593 ( \35970 , \35968 , \35969 );
not \U$35594 ( \35971 , \35970 );
nand \U$35595 ( \35972 , \35941 , \35971 );
not \U$35596 ( \35973 , \35972 );
not \U$35597 ( \35974 , \13158 );
xor \U$35598 ( \35975 , \4972 , RIae7a150_172);
not \U$35599 ( \35976 , \35975 );
or \U$35600 ( \35977 , \35974 , \35976 );
nand \U$35601 ( \35978 , \34113 , \9776 );
nand \U$35602 ( \35979 , \35977 , \35978 );
not \U$35603 ( \35980 , \35979 );
or \U$35604 ( \35981 , \35973 , \35980 );
nand \U$35605 ( \35982 , \35940 , \35970 );
nand \U$35606 ( \35983 , \35981 , \35982 );
nand \U$35607 ( \35984 , \35930 , \35983 );
or \U$35608 ( \35985 , \35928 , \35892 );
nand \U$35609 ( \35986 , \35984 , \35985 );
and \U$35610 ( \35987 , \35855 , \35986 );
and \U$35611 ( \35988 , \35852 , \35854 );
or \U$35612 ( \35989 , \35987 , \35988 );
and \U$35613 ( \35990 , \34176 , \34266 );
not \U$35614 ( \35991 , \34176 );
and \U$35615 ( \35992 , \35991 , \34267 );
or \U$35616 ( \35993 , \35990 , \35992 );
xor \U$35617 ( \35994 , \35989 , \35993 );
not \U$35618 ( \35995 , \12371 );
not \U$35619 ( \35996 , \35694 );
or \U$35620 ( \35997 , \35995 , \35996 );
not \U$35621 ( \35998 , \10625 );
not \U$35622 ( \35999 , \5722 );
or \U$35623 ( \36000 , \35998 , \35999 );
nand \U$35624 ( \36001 , \15207 , RIae7a498_179);
nand \U$35625 ( \36002 , \36000 , \36001 );
nand \U$35626 ( \36003 , \36002 , \11434 );
nand \U$35627 ( \36004 , \35997 , \36003 );
not \U$35628 ( \36005 , \17797 );
xor \U$35629 ( \36006 , RIae7a060_170, \24742 );
not \U$35630 ( \36007 , \36006 );
or \U$35631 ( \36008 , \36005 , \36007 );
nand \U$35632 ( \36009 , \35757 , \11098 );
nand \U$35633 ( \36010 , \36008 , \36009 );
xor \U$35634 ( \36011 , \36004 , \36010 );
not \U$35635 ( \36012 , \10510 );
and \U$35636 ( \36013 , RIae7a7e0_186, \2385 );
not \U$35637 ( \36014 , RIae7a7e0_186);
and \U$35638 ( \36015 , \36014 , \1860 );
nor \U$35639 ( \36016 , \36013 , \36015 );
not \U$35640 ( \36017 , \36016 );
or \U$35641 ( \36018 , \36012 , \36017 );
nand \U$35642 ( \36019 , \35688 , \10519 );
nand \U$35643 ( \36020 , \36018 , \36019 );
and \U$35644 ( \36021 , \36011 , \36020 );
and \U$35645 ( \36022 , \36004 , \36010 );
nor \U$35646 ( \36023 , \36021 , \36022 );
not \U$35647 ( \36024 , \36023 );
not \U$35648 ( \36025 , \36024 );
and \U$35649 ( \36026 , \34193 , \34203 );
not \U$35650 ( \36027 , \34193 );
not \U$35651 ( \36028 , \34203 );
and \U$35652 ( \36029 , \36027 , \36028 );
nor \U$35653 ( \36030 , \36026 , \36029 );
not \U$35654 ( \36031 , \34106 );
not \U$35655 ( \36032 , \34117 );
not \U$35656 ( \36033 , \36032 );
or \U$35657 ( \36034 , \36031 , \36033 );
or \U$35658 ( \36035 , \36032 , \34106 );
nand \U$35659 ( \36036 , \36034 , \36035 );
xor \U$35660 ( \36037 , \36030 , \36036 );
not \U$35661 ( \36038 , \36037 );
or \U$35662 ( \36039 , \36025 , \36038 );
nand \U$35663 ( \36040 , \36036 , \36030 );
nand \U$35664 ( \36041 , \36039 , \36040 );
not \U$35665 ( \36042 , \36041 );
not \U$35666 ( \36043 , \34211 );
not \U$35667 ( \36044 , \36043 );
not \U$35668 ( \36045 , \34252 );
or \U$35669 ( \36046 , \36044 , \36045 );
or \U$35670 ( \36047 , \34252 , \36043 );
nand \U$35671 ( \36048 , \36046 , \36047 );
not \U$35672 ( \36049 , \36048 );
not \U$35673 ( \36050 , \34121 );
not \U$35674 ( \36051 , \36050 );
not \U$35675 ( \36052 , \34172 );
or \U$35676 ( \36053 , \36051 , \36052 );
or \U$35677 ( \36054 , \34172 , \36050 );
nand \U$35678 ( \36055 , \36053 , \36054 );
not \U$35679 ( \36056 , \36055 );
not \U$35680 ( \36057 , \36056 );
or \U$35681 ( \36058 , \36049 , \36057 );
not \U$35682 ( \36059 , \36048 );
nand \U$35683 ( \36060 , \36059 , \36055 );
nand \U$35684 ( \36061 , \36058 , \36060 );
not \U$35685 ( \36062 , \36061 );
or \U$35686 ( \36063 , \36042 , \36062 );
nand \U$35687 ( \36064 , \36055 , \36048 );
nand \U$35688 ( \36065 , \36063 , \36064 );
and \U$35689 ( \36066 , \35994 , \36065 );
and \U$35690 ( \36067 , \35989 , \35993 );
or \U$35691 ( \36068 , \36066 , \36067 );
not \U$35692 ( \36069 , \36068 );
not \U$35693 ( \36070 , \35709 );
not \U$35694 ( \36071 , \36070 );
not \U$35695 ( \36072 , \35721 );
or \U$35696 ( \36073 , \36071 , \36072 );
or \U$35697 ( \36074 , \35721 , \36070 );
nand \U$35698 ( \36075 , \36073 , \36074 );
not \U$35699 ( \36076 , \36075 );
or \U$35700 ( \36077 , \36069 , \36076 );
xor \U$35701 ( \36078 , \35788 , \35786 );
and \U$35702 ( \36079 , \36078 , \35737 );
not \U$35703 ( \36080 , \36078 );
not \U$35704 ( \36081 , \35737 );
and \U$35705 ( \36082 , \36080 , \36081 );
nor \U$35706 ( \36083 , \36079 , \36082 );
not \U$35707 ( \36084 , \36083 );
not \U$35708 ( \36085 , \36084 );
xor \U$35709 ( \36086 , \35781 , \35783 );
not \U$35710 ( \36087 , \34161 );
not \U$35711 ( \36088 , \34146 );
or \U$35712 ( \36089 , \36087 , \36088 );
or \U$35713 ( \36090 , \34161 , \34146 );
nand \U$35714 ( \36091 , \36089 , \36090 );
xor \U$35715 ( \36092 , \34159 , \36091 );
not \U$35716 ( \36093 , \14668 );
and \U$35717 ( \36094 , RIae7aa38_191, \4305 );
not \U$35718 ( \36095 , RIae7aa38_191);
and \U$35719 ( \36096 , \36095 , \3525 );
nor \U$35720 ( \36097 , \36094 , \36096 );
not \U$35721 ( \36098 , \36097 );
or \U$35722 ( \36099 , \36093 , \36098 );
nand \U$35723 ( \36100 , \35768 , RIae7aab0_192);
nand \U$35724 ( \36101 , \36099 , \36100 );
not \U$35725 ( \36102 , \36101 );
xnor \U$35726 ( \36103 , \34069 , \34097 );
not \U$35727 ( \36104 , \36103 );
not \U$35728 ( \36105 , \16594 );
and \U$35729 ( \36106 , RIae7a8d0_188, \15782 );
not \U$35730 ( \36107 , RIae7a8d0_188);
and \U$35731 ( \36108 , \36107 , \19456 );
nor \U$35732 ( \36109 , \36106 , \36108 );
not \U$35733 ( \36110 , \36109 );
or \U$35734 ( \36111 , \36105 , \36110 );
nand \U$35735 ( \36112 , \35681 , \10275 );
nand \U$35736 ( \36113 , \36111 , \36112 );
not \U$35737 ( \36114 , \36113 );
or \U$35738 ( \36115 , \36104 , \36114 );
or \U$35739 ( \36116 , \36113 , \36103 );
nand \U$35740 ( \36117 , \36115 , \36116 );
not \U$35741 ( \36118 , \36117 );
or \U$35742 ( \36119 , \36102 , \36118 );
not \U$35743 ( \36120 , \36103 );
nand \U$35744 ( \36121 , \36120 , \36113 );
nand \U$35745 ( \36122 , \36119 , \36121 );
xor \U$35746 ( \36123 , \36092 , \36122 );
not \U$35747 ( \36124 , \9473 );
and \U$35748 ( \36125 , \5912 , RIae7a6f0_184);
not \U$35749 ( \36126 , \5912 );
and \U$35750 ( \36127 , \36126 , \16101 );
nor \U$35751 ( \36128 , \36125 , \36127 );
not \U$35752 ( \36129 , \36128 );
or \U$35753 ( \36130 , \36124 , \36129 );
not \U$35754 ( \36131 , \35745 );
not \U$35755 ( \36132 , \9705 );
or \U$35756 ( \36133 , \36131 , \36132 );
nand \U$35757 ( \36134 , \36130 , \36133 );
not \U$35758 ( \36135 , \36134 );
not \U$35759 ( \36136 , \15337 );
not \U$35760 ( \36137 , \34064 );
or \U$35761 ( \36138 , \36136 , \36137 );
not \U$35762 ( \36139 , \2442 );
not \U$35763 ( \36140 , \10042 );
or \U$35764 ( \36141 , \36139 , \36140 );
or \U$35765 ( \36142 , \10042 , \2442 );
nand \U$35766 ( \36143 , \36141 , \36142 );
nand \U$35767 ( \36144 , \36143 , \2431 );
nand \U$35768 ( \36145 , \36138 , \36144 );
not \U$35769 ( \36146 , \36145 );
and \U$35770 ( \36147 , \12857 , \1918 );
not \U$35771 ( \36148 , \2321 );
not \U$35772 ( \36149 , \35963 );
or \U$35773 ( \36150 , \36148 , \36149 );
not \U$35774 ( \36151 , RIae798e0_154);
not \U$35775 ( \36152 , \12750 );
or \U$35776 ( \36153 , \36151 , \36152 );
or \U$35777 ( \36154 , \16006 , RIae798e0_154);
nand \U$35778 ( \36155 , \36153 , \36154 );
nand \U$35779 ( \36156 , \36155 , \2338 );
nand \U$35780 ( \36157 , \36150 , \36156 );
xor \U$35781 ( \36158 , \36147 , \36157 );
not \U$35782 ( \36159 , \2007 );
not \U$35783 ( \36160 , \35948 );
or \U$35784 ( \36161 , \36159 , \36160 );
xnor \U$35785 ( \36162 , \10259 , RIae797f0_152);
nand \U$35786 ( \36163 , \36162 , \1987 );
nand \U$35787 ( \36164 , \36161 , \36163 );
and \U$35788 ( \36165 , \36158 , \36164 );
and \U$35789 ( \36166 , \36147 , \36157 );
nor \U$35790 ( \36167 , \36165 , \36166 );
not \U$35791 ( \36168 , \36167 );
and \U$35792 ( \36169 , \36146 , \36168 );
and \U$35793 ( \36170 , \36145 , \36167 );
nor \U$35794 ( \36171 , \36169 , \36170 );
not \U$35795 ( \36172 , \36171 );
not \U$35796 ( \36173 , \36172 );
not \U$35797 ( \36174 , \10573 );
not \U$35798 ( \36175 , \35834 );
or \U$35799 ( \36176 , \36174 , \36175 );
and \U$35800 ( \36177 , \15650 , RIae79ef8_167);
not \U$35801 ( \36178 , \15650 );
and \U$35802 ( \36179 , \36178 , \28303 );
nor \U$35803 ( \36180 , \36177 , \36179 );
nand \U$35804 ( \36181 , \36180 , \14768 );
nand \U$35805 ( \36182 , \36176 , \36181 );
not \U$35806 ( \36183 , \36182 );
or \U$35807 ( \36184 , \36173 , \36183 );
not \U$35808 ( \36185 , \36167 );
nand \U$35809 ( \36186 , \36185 , \36145 );
nand \U$35810 ( \36187 , \36184 , \36186 );
not \U$35811 ( \36188 , \2418 );
not \U$35812 ( \36189 , \35815 );
or \U$35813 ( \36190 , \36188 , \36189 );
not \U$35814 ( \36191 , RIae79c28_161);
not \U$35815 ( \36192 , \10149 );
or \U$35816 ( \36193 , \36191 , \36192 );
or \U$35817 ( \36194 , \10149 , RIae79c28_161);
nand \U$35818 ( \36195 , \36193 , \36194 );
nand \U$35819 ( \36196 , \36195 , \2417 );
nand \U$35820 ( \36197 , \36190 , \36196 );
not \U$35821 ( \36198 , \5049 );
not \U$35822 ( \36199 , \35861 );
or \U$35823 ( \36200 , \36198 , \36199 );
not \U$35824 ( \36201 , \11272 );
and \U$35825 ( \36202 , RIae79d90_164, \36201 );
not \U$35826 ( \36203 , RIae79d90_164);
not \U$35827 ( \36204 , \10168 );
and \U$35828 ( \36205 , \36203 , \36204 );
or \U$35829 ( \36206 , \36202 , \36205 );
nand \U$35830 ( \36207 , \36206 , \6091 );
nand \U$35831 ( \36208 , \36200 , \36207 );
xor \U$35832 ( \36209 , \36197 , \36208 );
not \U$35833 ( \36210 , \4853 );
not \U$35834 ( \36211 , \35869 );
or \U$35835 ( \36212 , \36210 , \36211 );
and \U$35836 ( \36213 , \10007 , RIae79ca0_162);
not \U$35837 ( \36214 , \10007 );
and \U$35838 ( \36215 , \36214 , \6270 );
nor \U$35839 ( \36216 , \36213 , \36215 );
nand \U$35840 ( \36217 , \36216 , \11761 );
nand \U$35841 ( \36218 , \36212 , \36217 );
and \U$35842 ( \36219 , \36209 , \36218 );
and \U$35843 ( \36220 , \36197 , \36208 );
nor \U$35844 ( \36221 , \36219 , \36220 );
xnor \U$35845 ( \36222 , \36187 , \36221 );
not \U$35846 ( \36223 , \36222 );
or \U$35847 ( \36224 , \36135 , \36223 );
not \U$35848 ( \36225 , \36221 );
nand \U$35849 ( \36226 , \36225 , \36187 );
nand \U$35850 ( \36227 , \36224 , \36226 );
and \U$35851 ( \36228 , \36123 , \36227 );
and \U$35852 ( \36229 , \36092 , \36122 );
or \U$35853 ( \36230 , \36228 , \36229 );
xor \U$35854 ( \36231 , \36086 , \36230 );
xor \U$35855 ( \36232 , \35666 , \35672 );
xor \U$35856 ( \36233 , \36232 , \35701 );
and \U$35857 ( \36234 , \36231 , \36233 );
and \U$35858 ( \36235 , \36086 , \36230 );
or \U$35859 ( \36236 , \36234 , \36235 );
not \U$35860 ( \36237 , \36236 );
or \U$35861 ( \36238 , \36085 , \36237 );
not \U$35862 ( \36239 , \36083 );
not \U$35863 ( \36240 , \36236 );
not \U$35864 ( \36241 , \36240 );
or \U$35865 ( \36242 , \36239 , \36241 );
xor \U$35866 ( \36243 , \35665 , \35704 );
xor \U$35867 ( \36244 , \36243 , \35706 );
nand \U$35868 ( \36245 , \36242 , \36244 );
nand \U$35869 ( \36246 , \36238 , \36245 );
not \U$35870 ( \36247 , \36246 );
nand \U$35871 ( \36248 , \36077 , \36247 );
not \U$35872 ( \36249 , \36068 );
not \U$35873 ( \36250 , \36075 );
nand \U$35874 ( \36251 , \36249 , \36250 );
nand \U$35875 ( \36252 , \36248 , \36251 );
not \U$35876 ( \36253 , \36252 );
not \U$35877 ( \36254 , \36253 );
or \U$35878 ( \36255 , \35804 , \36254 );
or \U$35879 ( \36256 , \35803 , \36253 );
nand \U$35880 ( \36257 , \36255 , \36256 );
not \U$35881 ( \36258 , \36257 );
or \U$35882 ( \36259 , \35801 , \36258 );
not \U$35883 ( \36260 , \36253 );
nand \U$35884 ( \36261 , \36260 , \35803 );
nand \U$35885 ( \36262 , \36259 , \36261 );
not \U$35886 ( \36263 , \36262 );
not \U$35887 ( \36264 , \36263 );
and \U$35888 ( \36265 , \33269 , \33279 );
not \U$35889 ( \36266 , \33269 );
not \U$35890 ( \36267 , \33279 );
and \U$35891 ( \36268 , \36266 , \36267 );
nor \U$35892 ( \36269 , \36265 , \36268 );
not \U$35893 ( \36270 , \33300 );
and \U$35894 ( \36271 , \36269 , \36270 );
not \U$35895 ( \36272 , \36269 );
and \U$35896 ( \36273 , \36272 , \33300 );
nor \U$35897 ( \36274 , \36271 , \36273 );
not \U$35898 ( \36275 , \36274 );
not \U$35899 ( \36276 , \36275 );
not \U$35900 ( \36277 , \35733 );
not \U$35901 ( \36278 , \35730 );
or \U$35902 ( \36279 , \36277 , \36278 );
nand \U$35903 ( \36280 , \36279 , \35799 );
nand \U$35904 ( \36281 , \35729 , \35726 );
and \U$35905 ( \36282 , \36280 , \36281 );
not \U$35906 ( \36283 , \36282 );
or \U$35907 ( \36284 , \36276 , \36283 );
not \U$35908 ( \36285 , \36281 );
not \U$35909 ( \36286 , \36280 );
or \U$35910 ( \36287 , \36285 , \36286 );
nand \U$35911 ( \36288 , \36287 , \36274 );
nand \U$35912 ( \36289 , \36284 , \36288 );
not \U$35913 ( \36290 , \36289 );
not \U$35914 ( \36291 , \33797 );
not \U$35915 ( \36292 , \34288 );
or \U$35916 ( \36293 , \36291 , \36292 );
nand \U$35917 ( \36294 , \33796 , \33655 );
nand \U$35918 ( \36295 , \36293 , \36294 );
and \U$35919 ( \36296 , \36295 , \34286 );
not \U$35920 ( \36297 , \36295 );
not \U$35921 ( \36298 , \34286 );
and \U$35922 ( \36299 , \36297 , \36298 );
nor \U$35923 ( \36300 , \36296 , \36299 );
not \U$35924 ( \36301 , \36300 );
or \U$35925 ( \36302 , \36290 , \36301 );
or \U$35926 ( \36303 , \36289 , \36300 );
nand \U$35927 ( \36304 , \36302 , \36303 );
nand \U$35928 ( \36305 , \36264 , \36304 );
not \U$35929 ( \36306 , \36300 );
not \U$35930 ( \36307 , \36306 );
not \U$35931 ( \36308 , \36289 );
or \U$35932 ( \36309 , \36307 , \36308 );
nand \U$35933 ( \36310 , \36280 , \36281 , \36274 );
nand \U$35934 ( \36311 , \36309 , \36310 );
xor \U$35935 ( \36312 , \33654 , \34290 );
xor \U$35936 ( \36313 , \36312 , \34298 );
nand \U$35937 ( \36314 , \36311 , \36313 );
not \U$35938 ( \36315 , \35800 );
not \U$35939 ( \36316 , \36257 );
not \U$35940 ( \36317 , \36316 );
or \U$35941 ( \36318 , \36315 , \36317 );
not \U$35942 ( \36319 , \35800 );
nand \U$35943 ( \36320 , \36319 , \36257 );
nand \U$35944 ( \36321 , \36318 , \36320 );
buf \U$35945 ( \36322 , \36075 );
xor \U$35946 ( \36323 , \36068 , \36322 );
xnor \U$35947 ( \36324 , \36323 , \36246 );
not \U$35948 ( \36325 , \36324 );
xor \U$35949 ( \36326 , \35792 , \35793 );
xor \U$35950 ( \36327 , \36326 , \35796 );
not \U$35951 ( \36328 , \36327 );
not \U$35952 ( \36329 , \36328 );
xnor \U$35953 ( \36330 , \36023 , \36037 );
not \U$35954 ( \36331 , \36330 );
xor \U$35955 ( \36332 , \36092 , \36122 );
xor \U$35956 ( \36333 , \36332 , \36227 );
xor \U$35957 ( \36334 , \36004 , \36010 );
xor \U$35958 ( \36335 , \36334 , \36020 );
not \U$35959 ( \36336 , \36335 );
not \U$35960 ( \36337 , \9517 );
not \U$35961 ( \36338 , \35935 );
or \U$35962 ( \36339 , \36337 , \36338 );
and \U$35963 ( \36340 , RIae79fe8_169, \10461 );
not \U$35964 ( \36341 , RIae79fe8_169);
and \U$35965 ( \36342 , \36341 , \15504 );
or \U$35966 ( \36343 , \36340 , \36342 );
nand \U$35967 ( \36344 , \36343 , \11913 );
nand \U$35968 ( \36345 , \36339 , \36344 );
not \U$35969 ( \36346 , \10696 );
xor \U$35970 ( \36347 , \6347 , RIae7a498_179);
not \U$35971 ( \36348 , \36347 );
or \U$35972 ( \36349 , \36346 , \36348 );
nand \U$35973 ( \36350 , \36002 , \10676 );
nand \U$35974 ( \36351 , \36349 , \36350 );
xor \U$35975 ( \36352 , \36345 , \36351 );
not \U$35976 ( \36353 , \9777 );
not \U$35977 ( \36354 , \35975 );
or \U$35978 ( \36355 , \36353 , \36354 );
xor \U$35979 ( \36356 , RIae7a150_172, \6256 );
nand \U$35980 ( \36357 , \36356 , \10667 );
nand \U$35981 ( \36358 , \36355 , \36357 );
and \U$35982 ( \36359 , \36352 , \36358 );
and \U$35983 ( \36360 , \36345 , \36351 );
nor \U$35984 ( \36361 , \36359 , \36360 );
not \U$35985 ( \36362 , \9622 );
not \U$35986 ( \36363 , \35899 );
not \U$35987 ( \36364 , \36363 );
or \U$35988 ( \36365 , \36362 , \36364 );
and \U$35989 ( \36366 , RIae7a3a8_177, \9367 );
not \U$35990 ( \36367 , RIae7a3a8_177);
and \U$35991 ( \36368 , \36367 , \13287 );
nor \U$35992 ( \36369 , \36366 , \36368 );
nand \U$35993 ( \36370 , \9644 , \36369 );
nand \U$35994 ( \36371 , \36365 , \36370 );
not \U$35995 ( \36372 , \36371 );
not \U$35996 ( \36373 , \35966 );
not \U$35997 ( \36374 , \35950 );
not \U$35998 ( \36375 , \36374 );
and \U$35999 ( \36376 , \36373 , \36375 );
and \U$36000 ( \36377 , \35966 , \36374 );
nor \U$36001 ( \36378 , \36376 , \36377 );
not \U$36002 ( \36379 , \36378 );
not \U$36003 ( \36380 , \10631 );
not \U$36004 ( \36381 , \35885 );
or \U$36005 ( \36382 , \36380 , \36381 );
and \U$36006 ( \36383 , \15102 , RIae7a510_180);
not \U$36007 ( \36384 , \15102 );
and \U$36008 ( \36385 , \36384 , \14931 );
nor \U$36009 ( \36386 , \36383 , \36385 );
nand \U$36010 ( \36387 , \36386 , \10927 );
nand \U$36011 ( \36388 , \36382 , \36387 );
not \U$36012 ( \36389 , \36388 );
or \U$36013 ( \36390 , \36379 , \36389 );
or \U$36014 ( \36391 , \36388 , \36378 );
nand \U$36015 ( \36392 , \36390 , \36391 );
not \U$36016 ( \36393 , \36392 );
or \U$36017 ( \36394 , \36372 , \36393 );
not \U$36018 ( \36395 , \36378 );
nand \U$36019 ( \36396 , \36395 , \36388 );
nand \U$36020 ( \36397 , \36394 , \36396 );
xnor \U$36021 ( \36398 , \36361 , \36397 );
not \U$36022 ( \36399 , \36398 );
or \U$36023 ( \36400 , \36336 , \36399 );
not \U$36024 ( \36401 , \36361 );
nand \U$36025 ( \36402 , \36401 , \36397 );
nand \U$36026 ( \36403 , \36400 , \36402 );
or \U$36027 ( \36404 , \36333 , \36403 );
not \U$36028 ( \36405 , \36404 );
or \U$36029 ( \36406 , \36331 , \36405 );
nand \U$36030 ( \36407 , \36333 , \36403 );
nand \U$36031 ( \36408 , \36406 , \36407 );
not \U$36032 ( \36409 , \36408 );
and \U$36033 ( \36410 , \36061 , \36041 );
not \U$36034 ( \36411 , \36061 );
not \U$36035 ( \36412 , \36041 );
and \U$36036 ( \36413 , \36411 , \36412 );
nor \U$36037 ( \36414 , \36410 , \36413 );
not \U$36038 ( \36415 , \36414 );
or \U$36039 ( \36416 , \36409 , \36415 );
xor \U$36040 ( \36417 , \36086 , \36230 );
xor \U$36041 ( \36418 , \36417 , \36233 );
not \U$36042 ( \36419 , \36418 );
nand \U$36043 ( \36420 , \36416 , \36419 );
or \U$36044 ( \36421 , \36408 , \36414 );
nand \U$36045 ( \36422 , \36420 , \36421 );
not \U$36046 ( \36423 , \36422 );
xor \U$36047 ( \36424 , \35902 , \35923 );
not \U$36048 ( \36425 , \36424 );
and \U$36049 ( \36426 , \35940 , \35970 );
not \U$36050 ( \36427 , \35940 );
and \U$36051 ( \36428 , \36427 , \35971 );
nor \U$36052 ( \36429 , \36426 , \36428 );
and \U$36053 ( \36430 , \35979 , \36429 );
not \U$36054 ( \36431 , \35979 );
not \U$36055 ( \36432 , \36429 );
and \U$36056 ( \36433 , \36431 , \36432 );
nor \U$36057 ( \36434 , \36430 , \36433 );
nand \U$36058 ( \36435 , \36425 , \36434 );
not \U$36059 ( \36436 , \36435 );
not \U$36060 ( \36437 , RIae7aab0_192);
not \U$36061 ( \36438 , \36097 );
or \U$36062 ( \36439 , \36437 , \36438 );
and \U$36063 ( \36440 , \2576 , RIae7aa38_191);
not \U$36064 ( \36441 , \2576 );
and \U$36065 ( \36442 , \36441 , \11326 );
nor \U$36066 ( \36443 , \36440 , \36442 );
nand \U$36067 ( \36444 , \36443 , \14668 );
nand \U$36068 ( \36445 , \36439 , \36444 );
not \U$36069 ( \36446 , \36445 );
not \U$36070 ( \36447 , \36446 );
not \U$36071 ( \36448 , \11098 );
not \U$36072 ( \36449 , \36006 );
or \U$36073 ( \36450 , \36448 , \36449 );
not \U$36074 ( \36451 , RIae7a060_170);
not \U$36075 ( \36452 , \21873 );
or \U$36076 ( \36453 , \36451 , \36452 );
or \U$36077 ( \36454 , \4929 , RIae7a060_170);
nand \U$36078 ( \36455 , \36453 , \36454 );
nand \U$36079 ( \36456 , \36455 , \9730 );
nand \U$36080 ( \36457 , \36450 , \36456 );
not \U$36081 ( \36458 , \36457 );
not \U$36082 ( \36459 , \9527 );
not \U$36083 ( \36460 , \36016 );
or \U$36084 ( \36461 , \36459 , \36460 );
xor \U$36085 ( \36462 , \5673 , RIae7a7e0_186);
nand \U$36086 ( \36463 , \36462 , \11439 );
nand \U$36087 ( \36464 , \36461 , \36463 );
not \U$36088 ( \36465 , \36464 );
and \U$36089 ( \36466 , \36458 , \36465 );
not \U$36090 ( \36467 , \36458 );
and \U$36091 ( \36468 , \36467 , \36464 );
nor \U$36092 ( \36469 , \36466 , \36468 );
not \U$36093 ( \36470 , \36469 );
or \U$36094 ( \36471 , \36447 , \36470 );
nand \U$36095 ( \36472 , \36458 , \36465 );
nand \U$36096 ( \36473 , \36471 , \36472 );
not \U$36097 ( \36474 , \36473 );
or \U$36098 ( \36475 , \36436 , \36474 );
not \U$36099 ( \36476 , \36434 );
nand \U$36100 ( \36477 , \36476 , \36424 );
nand \U$36101 ( \36478 , \36475 , \36477 );
not \U$36102 ( \36479 , \36478 );
nand \U$36103 ( \36480 , \35850 , \35844 );
xor \U$36104 ( \36481 , \36480 , \35846 );
not \U$36105 ( \36482 , \36481 );
xor \U$36106 ( \36483 , \35892 , \35983 );
xnor \U$36107 ( \36484 , \36483 , \35928 );
not \U$36108 ( \36485 , \36484 );
or \U$36109 ( \36486 , \36482 , \36485 );
or \U$36110 ( \36487 , \36484 , \36481 );
nand \U$36111 ( \36488 , \36486 , \36487 );
not \U$36112 ( \36489 , \36488 );
or \U$36113 ( \36490 , \36479 , \36489 );
not \U$36114 ( \36491 , \36481 );
nand \U$36115 ( \36492 , \36491 , \36484 );
nand \U$36116 ( \36493 , \36490 , \36492 );
not \U$36117 ( \36494 , \36493 );
not \U$36118 ( \36495 , \35749 );
and \U$36119 ( \36496 , \35775 , \36495 );
not \U$36120 ( \36497 , \35775 );
and \U$36121 ( \36498 , \36497 , \35749 );
or \U$36122 ( \36499 , \36496 , \36498 );
not \U$36123 ( \36500 , \36499 );
xnor \U$36124 ( \36501 , \35826 , \35838 );
not \U$36125 ( \36502 , \36501 );
not \U$36126 ( \36503 , \35889 );
not \U$36127 ( \36504 , \35878 );
or \U$36128 ( \36505 , \36503 , \36504 );
or \U$36129 ( \36506 , \35889 , \35878 );
nand \U$36130 ( \36507 , \36505 , \36506 );
not \U$36131 ( \36508 , \36507 );
or \U$36132 ( \36509 , \36502 , \36508 );
or \U$36133 ( \36510 , \36507 , \36501 );
not \U$36134 ( \36511 , \13121 );
not \U$36135 ( \36512 , \35916 );
or \U$36136 ( \36513 , \36511 , \36512 );
not \U$36137 ( \36514 , RIae7a240_174);
not \U$36138 ( \36515 , \13301 );
or \U$36139 ( \36516 , \36514 , \36515 );
or \U$36140 ( \36517 , \14657 , RIae7a240_174);
nand \U$36141 ( \36518 , \36516 , \36517 );
nand \U$36142 ( \36519 , \36518 , \9688 );
nand \U$36143 ( \36520 , \36513 , \36519 );
not \U$36144 ( \36521 , \36520 );
not \U$36145 ( \36522 , \9814 );
not \U$36146 ( \36523 , \35905 );
or \U$36147 ( \36524 , \36522 , \36523 );
not \U$36148 ( \36525 , \9412 );
xor \U$36149 ( \36526 , RIae7a2b8_175, \36525 );
nand \U$36150 ( \36527 , \36526 , \9792 );
nand \U$36151 ( \36528 , \36524 , \36527 );
not \U$36152 ( \36529 , \2417 );
xor \U$36153 ( \36530 , \10031 , RIae79c28_161);
not \U$36154 ( \36531 , \36530 );
or \U$36155 ( \36532 , \36529 , \36531 );
nand \U$36156 ( \36533 , \36195 , \2418 );
nand \U$36157 ( \36534 , \36532 , \36533 );
not \U$36158 ( \36535 , \36534 );
or \U$36159 ( \36536 , \16890 , \2320 );
not \U$36160 ( \36537 , \2319 );
nand \U$36161 ( \36538 , \36536 , \36537 , RIae798e0_154);
not \U$36162 ( \36539 , \36538 );
not \U$36163 ( \36540 , \2321 );
not \U$36164 ( \36541 , \36155 );
or \U$36165 ( \36542 , \36540 , \36541 );
and \U$36166 ( \36543 , RIae798e0_154, \12857 );
not \U$36167 ( \36544 , RIae798e0_154);
not \U$36168 ( \36545 , \12858 );
and \U$36169 ( \36546 , \36544 , \36545 );
nor \U$36170 ( \36547 , \36543 , \36546 );
nand \U$36171 ( \36548 , \36547 , \2338 );
nand \U$36172 ( \36549 , \36542 , \36548 );
nand \U$36173 ( \36550 , \36539 , \36549 );
not \U$36174 ( \36551 , \36550 );
not \U$36175 ( \36552 , \2450 );
not \U$36176 ( \36553 , \36143 );
or \U$36177 ( \36554 , \36552 , \36553 );
and \U$36178 ( \36555 , RIae79778_151, \10193 );
not \U$36179 ( \36556 , RIae79778_151);
and \U$36180 ( \36557 , \36556 , \19689 );
nor \U$36181 ( \36558 , \36555 , \36557 );
nand \U$36182 ( \36559 , \36558 , \2431 );
nand \U$36183 ( \36560 , \36554 , \36559 );
not \U$36184 ( \36561 , \36560 );
or \U$36185 ( \36562 , \36551 , \36561 );
or \U$36186 ( \36563 , \36560 , \36550 );
nand \U$36187 ( \36564 , \36562 , \36563 );
not \U$36188 ( \36565 , \36564 );
or \U$36189 ( \36566 , \36535 , \36565 );
not \U$36190 ( \36567 , \36550 );
nand \U$36191 ( \36568 , \36567 , \36560 );
nand \U$36192 ( \36569 , \36566 , \36568 );
and \U$36193 ( \36570 , \36528 , \36569 );
not \U$36194 ( \36571 , \36528 );
not \U$36195 ( \36572 , \36569 );
and \U$36196 ( \36573 , \36571 , \36572 );
nor \U$36197 ( \36574 , \36570 , \36573 );
not \U$36198 ( \36575 , \36574 );
or \U$36199 ( \36576 , \36521 , \36575 );
nand \U$36200 ( \36577 , \36528 , \36569 );
nand \U$36201 ( \36578 , \36576 , \36577 );
nand \U$36202 ( \36579 , \36510 , \36578 );
nand \U$36203 ( \36580 , \36509 , \36579 );
not \U$36204 ( \36581 , \36580 );
or \U$36205 ( \36582 , \36500 , \36581 );
xor \U$36206 ( \36583 , \35683 , \35697 );
not \U$36207 ( \36584 , \36583 );
nand \U$36208 ( \36585 , \36582 , \36584 );
not \U$36209 ( \36586 , \36580 );
not \U$36210 ( \36587 , \36499 );
nand \U$36211 ( \36588 , \36586 , \36587 );
nand \U$36212 ( \36589 , \36585 , \36588 );
not \U$36213 ( \36590 , \36589 );
not \U$36214 ( \36591 , \36590 );
xor \U$36215 ( \36592 , \35852 , \35854 );
xor \U$36216 ( \36593 , \36592 , \35986 );
not \U$36217 ( \36594 , \36593 );
not \U$36218 ( \36595 , \36594 );
or \U$36219 ( \36596 , \36591 , \36595 );
nand \U$36220 ( \36597 , \36593 , \36589 );
nand \U$36221 ( \36598 , \36596 , \36597 );
not \U$36222 ( \36599 , \36598 );
or \U$36223 ( \36600 , \36494 , \36599 );
not \U$36224 ( \36601 , \36593 );
nand \U$36225 ( \36602 , \36601 , \36589 );
nand \U$36226 ( \36603 , \36600 , \36602 );
not \U$36227 ( \36604 , \36603 );
xor \U$36228 ( \36605 , \35989 , \35993 );
xor \U$36229 ( \36606 , \36605 , \36065 );
not \U$36230 ( \36607 , \36606 );
or \U$36231 ( \36608 , \36604 , \36607 );
or \U$36232 ( \36609 , \36606 , \36603 );
nand \U$36233 ( \36610 , \36608 , \36609 );
not \U$36234 ( \36611 , \36610 );
or \U$36235 ( \36612 , \36423 , \36611 );
not \U$36236 ( \36613 , \36606 );
nand \U$36237 ( \36614 , \36613 , \36603 );
nand \U$36238 ( \36615 , \36612 , \36614 );
not \U$36239 ( \36616 , \36615 );
not \U$36240 ( \36617 , \36616 );
or \U$36241 ( \36618 , \36329 , \36617 );
nand \U$36242 ( \36619 , \36615 , \36327 );
nand \U$36243 ( \36620 , \36618 , \36619 );
not \U$36244 ( \36621 , \36620 );
or \U$36245 ( \36622 , \36325 , \36621 );
nand \U$36246 ( \36623 , \36615 , \36328 );
nand \U$36247 ( \36624 , \36622 , \36623 );
nand \U$36248 ( \36625 , \36321 , \36624 );
and \U$36249 ( \36626 , \36620 , \36324 );
not \U$36250 ( \36627 , \36620 );
not \U$36251 ( \36628 , \36324 );
and \U$36252 ( \36629 , \36627 , \36628 );
nor \U$36253 ( \36630 , \36626 , \36629 );
xnor \U$36254 ( \36631 , \36422 , \36610 );
not \U$36255 ( \36632 , \36631 );
not \U$36256 ( \36633 , \36632 );
not \U$36257 ( \36634 , \36240 );
not \U$36258 ( \36635 , \36244 );
or \U$36259 ( \36636 , \36634 , \36635 );
not \U$36260 ( \36637 , \36244 );
nand \U$36261 ( \36638 , \36637 , \36236 );
nand \U$36262 ( \36639 , \36636 , \36638 );
not \U$36263 ( \36640 , \36084 );
xnor \U$36264 ( \36641 , \36639 , \36640 );
not \U$36265 ( \36642 , \36641 );
xor \U$36266 ( \36643 , \36564 , \36534 );
not \U$36267 ( \36644 , \35747 );
and \U$36268 ( \36645 , RIae7a6f0_184, \1860 );
not \U$36269 ( \36646 , RIae7a6f0_184);
and \U$36270 ( \36647 , \36646 , \2385 );
or \U$36271 ( \36648 , \36645 , \36647 );
not \U$36272 ( \36649 , \36648 );
or \U$36273 ( \36650 , \36644 , \36649 );
not \U$36274 ( \36651 , \3216 );
not \U$36275 ( \36652 , RIae7a6f0_184);
and \U$36276 ( \36653 , \36651 , \36652 );
and \U$36277 ( \36654 , \1970 , RIae7a6f0_184);
nor \U$36278 ( \36655 , \36653 , \36654 );
not \U$36279 ( \36656 , \9478 );
or \U$36280 ( \36657 , \36655 , \36656 );
nand \U$36281 ( \36658 , \36650 , \36657 );
xor \U$36282 ( \36659 , \36643 , \36658 );
not \U$36283 ( \36660 , \14668 );
and \U$36284 ( \36661 , RIae7aa38_191, \2564 );
not \U$36285 ( \36662 , RIae7aa38_191);
and \U$36286 ( \36663 , \36662 , \15782 );
or \U$36287 ( \36664 , \36661 , \36663 );
not \U$36288 ( \36665 , \36664 );
or \U$36289 ( \36666 , \36660 , \36665 );
nand \U$36290 ( \36667 , \36443 , RIae7aab0_192);
nand \U$36291 ( \36668 , \36666 , \36667 );
and \U$36292 ( \36669 , \36659 , \36668 );
and \U$36293 ( \36670 , \36643 , \36658 );
or \U$36294 ( \36671 , \36669 , \36670 );
not \U$36295 ( \36672 , \36671 );
not \U$36296 ( \36673 , \14510 );
not \U$36297 ( \36674 , \11207 );
not \U$36298 ( \36675 , \5115 );
or \U$36299 ( \36676 , \36674 , \36675 );
or \U$36300 ( \36677 , \1956 , \11207 );
nand \U$36301 ( \36678 , \36676 , \36677 );
not \U$36302 ( \36679 , \36678 );
or \U$36303 ( \36680 , \36673 , \36679 );
and \U$36304 ( \36681 , RIae7a8d0_188, \13008 );
not \U$36305 ( \36682 , RIae7a8d0_188);
and \U$36306 ( \36683 , \36682 , \2089 );
or \U$36307 ( \36684 , \36681 , \36683 );
nand \U$36308 ( \36685 , \36684 , \10275 );
nand \U$36309 ( \36686 , \36680 , \36685 );
not \U$36310 ( \36687 , \36686 );
not \U$36311 ( \36688 , \36687 );
not \U$36312 ( \36689 , \16564 );
not \U$36313 ( \36690 , RIae7a498_179);
not \U$36314 ( \36691 , \17242 );
or \U$36315 ( \36692 , \36690 , \36691 );
or \U$36316 ( \36693 , \6231 , RIae7a498_179);
nand \U$36317 ( \36694 , \36692 , \36693 );
not \U$36318 ( \36695 , \36694 );
or \U$36319 ( \36696 , \36689 , \36695 );
nand \U$36320 ( \36697 , \36347 , \11422 );
nand \U$36321 ( \36698 , \36696 , \36697 );
not \U$36322 ( \36699 , \36698 );
not \U$36323 ( \36700 , \36699 );
or \U$36324 ( \36701 , \36688 , \36700 );
not \U$36325 ( \36702 , \9776 );
not \U$36326 ( \36703 , \36356 );
or \U$36327 ( \36704 , \36702 , \36703 );
and \U$36328 ( \36705 , RIae7a150_172, \13976 );
not \U$36329 ( \36706 , RIae7a150_172);
and \U$36330 ( \36707 , \36706 , \21732 );
or \U$36331 ( \36708 , \36705 , \36707 );
nand \U$36332 ( \36709 , \36708 , \10667 );
nand \U$36333 ( \36710 , \36704 , \36709 );
nand \U$36334 ( \36711 , \36701 , \36710 );
nand \U$36335 ( \36712 , \36698 , \36686 );
nand \U$36336 ( \36713 , \36711 , \36712 );
xor \U$36337 ( \36714 , \36371 , \36392 );
xor \U$36338 ( \36715 , \36713 , \36714 );
not \U$36339 ( \36716 , \36715 );
or \U$36340 ( \36717 , \36672 , \36716 );
nand \U$36341 ( \36718 , \36714 , \36713 );
nand \U$36342 ( \36719 , \36717 , \36718 );
not \U$36343 ( \36720 , \36134 );
and \U$36344 ( \36721 , \36222 , \36720 );
not \U$36345 ( \36722 , \36222 );
and \U$36346 ( \36723 , \36722 , \36134 );
nor \U$36347 ( \36724 , \36721 , \36723 );
not \U$36348 ( \36725 , \36724 );
or \U$36349 ( \36726 , \36719 , \36725 );
not \U$36350 ( \36727 , \9621 );
not \U$36351 ( \36728 , \36369 );
or \U$36352 ( \36729 , \36727 , \36728 );
not \U$36353 ( \36730 , \13165 );
not \U$36354 ( \36731 , \12614 );
or \U$36355 ( \36732 , \36730 , \36731 );
or \U$36356 ( \36733 , \12614 , \13165 );
nand \U$36357 ( \36734 , \36732 , \36733 );
nand \U$36358 ( \36735 , \36734 , \11013 );
nand \U$36359 ( \36736 , \36729 , \36735 );
not \U$36360 ( \36737 , \36736 );
not \U$36361 ( \36738 , \9687 );
not \U$36362 ( \36739 , RIae7a240_174);
not \U$36363 ( \36740 , \15488 );
or \U$36364 ( \36741 , \36739 , \36740 );
or \U$36365 ( \36742 , \16766 , RIae7a240_174);
nand \U$36366 ( \36743 , \36741 , \36742 );
not \U$36367 ( \36744 , \36743 );
or \U$36368 ( \36745 , \36738 , \36744 );
nand \U$36369 ( \36746 , \36518 , \9699 );
nand \U$36370 ( \36747 , \36745 , \36746 );
not \U$36371 ( \36748 , \36747 );
nand \U$36372 ( \36749 , \36737 , \36748 );
not \U$36373 ( \36750 , \36749 );
not \U$36374 ( \36751 , \10927 );
not \U$36375 ( \36752 , RIae7a510_180);
not \U$36376 ( \36753 , \12707 );
or \U$36377 ( \36754 , \36752 , \36753 );
or \U$36378 ( \36755 , \12707 , RIae7a510_180);
nand \U$36379 ( \36756 , \36754 , \36755 );
not \U$36380 ( \36757 , \36756 );
or \U$36381 ( \36758 , \36751 , \36757 );
nand \U$36382 ( \36759 , \36386 , \16358 );
nand \U$36383 ( \36760 , \36758 , \36759 );
not \U$36384 ( \36761 , \36760 );
or \U$36385 ( \36762 , \36750 , \36761 );
nand \U$36386 ( \36763 , \36747 , \36736 );
nand \U$36387 ( \36764 , \36762 , \36763 );
not \U$36388 ( \36765 , \36764 );
not \U$36389 ( \36766 , \36358 );
not \U$36390 ( \36767 , \36766 );
not \U$36391 ( \36768 , \36352 );
or \U$36392 ( \36769 , \36767 , \36768 );
or \U$36393 ( \36770 , \36352 , \36766 );
nand \U$36394 ( \36771 , \36769 , \36770 );
not \U$36395 ( \36772 , \36771 );
or \U$36396 ( \36773 , \36765 , \36772 );
or \U$36397 ( \36774 , \36771 , \36764 );
not \U$36398 ( \36775 , \9792 );
xor \U$36399 ( \36776 , \12482 , RIae7a2b8_175);
not \U$36400 ( \36777 , \36776 );
or \U$36401 ( \36778 , \36775 , \36777 );
nand \U$36402 ( \36779 , \36526 , \16135 );
nand \U$36403 ( \36780 , \36778 , \36779 );
not \U$36404 ( \36781 , \36780 );
not \U$36405 ( \36782 , \36549 );
not \U$36406 ( \36783 , \36538 );
and \U$36407 ( \36784 , \36782 , \36783 );
and \U$36408 ( \36785 , \36549 , \36538 );
nor \U$36409 ( \36786 , \36784 , \36785 );
not \U$36410 ( \36787 , \2007 );
not \U$36411 ( \36788 , \36162 );
or \U$36412 ( \36789 , \36787 , \36788 );
buf \U$36413 ( \36790 , \10845 );
and \U$36414 ( \36791 , RIae797f0_152, \36790 );
not \U$36415 ( \36792 , RIae797f0_152);
not \U$36416 ( \36793 , \36790 );
and \U$36417 ( \36794 , \36792 , \36793 );
nor \U$36418 ( \36795 , \36791 , \36794 );
nand \U$36419 ( \36796 , \36795 , \1987 );
nand \U$36420 ( \36797 , \36789 , \36796 );
xnor \U$36421 ( \36798 , \36786 , \36797 );
not \U$36422 ( \36799 , \36798 );
not \U$36423 ( \36800 , \2418 );
not \U$36424 ( \36801 , \36530 );
or \U$36425 ( \36802 , \36800 , \36801 );
not \U$36426 ( \36803 , \10584 );
not \U$36427 ( \36804 , \11665 );
or \U$36428 ( \36805 , \36803 , \36804 );
or \U$36429 ( \36806 , \16912 , \10584 );
nand \U$36430 ( \36807 , \36805 , \36806 );
nand \U$36431 ( \36808 , \36807 , \2417 );
nand \U$36432 ( \36809 , \36802 , \36808 );
not \U$36433 ( \36810 , \36809 );
or \U$36434 ( \36811 , \36799 , \36810 );
not \U$36435 ( \36812 , \36786 );
nand \U$36436 ( \36813 , \36812 , \36797 );
nand \U$36437 ( \36814 , \36811 , \36813 );
not \U$36438 ( \36815 , \36814 );
nand \U$36439 ( \36816 , \36781 , \36815 );
not \U$36440 ( \36817 , \36816 );
not \U$36441 ( \36818 , \11439 );
and \U$36442 ( \36819 , \13999 , \9541 );
not \U$36443 ( \36820 , \13999 );
and \U$36444 ( \36821 , \36820 , RIae7a7e0_186);
nor \U$36445 ( \36822 , \36819 , \36821 );
not \U$36446 ( \36823 , \36822 );
or \U$36447 ( \36824 , \36818 , \36823 );
nand \U$36448 ( \36825 , \36462 , \9527 );
nand \U$36449 ( \36826 , \36824 , \36825 );
not \U$36450 ( \36827 , \36826 );
or \U$36451 ( \36828 , \36817 , \36827 );
nand \U$36452 ( \36829 , \36814 , \36780 );
nand \U$36453 ( \36830 , \36828 , \36829 );
nand \U$36454 ( \36831 , \36774 , \36830 );
nand \U$36455 ( \36832 , \36773 , \36831 );
nand \U$36456 ( \36833 , \36726 , \36832 );
nand \U$36457 ( \36834 , \36719 , \36725 );
nand \U$36458 ( \36835 , \36833 , \36834 );
not \U$36459 ( \36836 , \36835 );
not \U$36460 ( \36837 , \10709 );
not \U$36461 ( \36838 , RIae79fe8_169);
not \U$36462 ( \36839 , \33593 );
or \U$36463 ( \36840 , \36838 , \36839 );
nand \U$36464 ( \36841 , \33592 , \9504 );
nand \U$36465 ( \36842 , \36840 , \36841 );
not \U$36466 ( \36843 , \36842 );
or \U$36467 ( \36844 , \36837 , \36843 );
nand \U$36468 ( \36845 , \36343 , \10700 );
nand \U$36469 ( \36846 , \36844 , \36845 );
not \U$36470 ( \36847 , \36846 );
not \U$36471 ( \36848 , \36164 );
and \U$36472 ( \36849 , \36158 , \36848 );
not \U$36473 ( \36850 , \36158 );
and \U$36474 ( \36851 , \36850 , \36164 );
nor \U$36475 ( \36852 , \36849 , \36851 );
not \U$36476 ( \36853 , \36852 );
not \U$36477 ( \36854 , \19362 );
and \U$36478 ( \36855 , RIae79ef8_167, \10070 );
not \U$36479 ( \36856 , RIae79ef8_167);
and \U$36480 ( \36857 , \36856 , \11230 );
nor \U$36481 ( \36858 , \36855 , \36857 );
not \U$36482 ( \36859 , \36858 );
or \U$36483 ( \36860 , \36854 , \36859 );
nand \U$36484 ( \36861 , \36180 , \6212 );
nand \U$36485 ( \36862 , \36860 , \36861 );
not \U$36486 ( \36863 , \36862 );
or \U$36487 ( \36864 , \36853 , \36863 );
or \U$36488 ( \36865 , \36862 , \36852 );
nand \U$36489 ( \36866 , \36864 , \36865 );
not \U$36490 ( \36867 , \36866 );
or \U$36491 ( \36868 , \36847 , \36867 );
not \U$36492 ( \36869 , \36852 );
nand \U$36493 ( \36870 , \36869 , \36862 );
nand \U$36494 ( \36871 , \36868 , \36870 );
xor \U$36495 ( \36872 , \36197 , \36208 );
xor \U$36496 ( \36873 , \36872 , \36218 );
xor \U$36497 ( \36874 , \36871 , \36873 );
not \U$36498 ( \36875 , \5039 );
not \U$36499 ( \36876 , RIae79d90_164);
not \U$36500 ( \36877 , \13896 );
or \U$36501 ( \36878 , \36876 , \36877 );
or \U$36502 ( \36879 , \9875 , RIae79d90_164);
nand \U$36503 ( \36880 , \36878 , \36879 );
not \U$36504 ( \36881 , \36880 );
or \U$36505 ( \36882 , \36875 , \36881 );
nand \U$36506 ( \36883 , \36206 , \5048 );
nand \U$36507 ( \36884 , \36882 , \36883 );
not \U$36508 ( \36885 , \36884 );
not \U$36509 ( \36886 , \4842 );
and \U$36510 ( \36887 , \19035 , \6270 );
not \U$36511 ( \36888 , \19035 );
and \U$36512 ( \36889 , \36888 , RIae79ca0_162);
nor \U$36513 ( \36890 , \36887 , \36889 );
not \U$36514 ( \36891 , \36890 );
or \U$36515 ( \36892 , \36886 , \36891 );
nand \U$36516 ( \36893 , \36216 , \4853 );
nand \U$36517 ( \36894 , \36892 , \36893 );
not \U$36518 ( \36895 , \36894 );
nand \U$36519 ( \36896 , \36885 , \36895 );
not \U$36520 ( \36897 , \36896 );
not \U$36521 ( \36898 , \9745 );
not \U$36522 ( \36899 , \36455 );
or \U$36523 ( \36900 , \36898 , \36899 );
and \U$36524 ( \36901 , \11102 , \17010 );
not \U$36525 ( \36902 , \11102 );
and \U$36526 ( \36903 , \36902 , \12724 );
nor \U$36527 ( \36904 , \36901 , \36903 );
nand \U$36528 ( \36905 , \36904 , \9730 );
nand \U$36529 ( \36906 , \36900 , \36905 );
not \U$36530 ( \36907 , \36906 );
or \U$36531 ( \36908 , \36897 , \36907 );
nand \U$36532 ( \36909 , \36884 , \36894 );
nand \U$36533 ( \36910 , \36908 , \36909 );
and \U$36534 ( \36911 , \36874 , \36910 );
and \U$36535 ( \36912 , \36871 , \36873 );
or \U$36536 ( \36913 , \36911 , \36912 );
not \U$36537 ( \36914 , \9478 );
not \U$36538 ( \36915 , \36128 );
or \U$36539 ( \36916 , \36914 , \36915 );
not \U$36540 ( \36917 , \36655 );
nand \U$36541 ( \36918 , \36917 , \35747 );
nand \U$36542 ( \36919 , \36916 , \36918 );
not \U$36543 ( \36920 , \36919 );
not \U$36544 ( \36921 , \36182 );
not \U$36545 ( \36922 , \36171 );
and \U$36546 ( \36923 , \36921 , \36922 );
and \U$36547 ( \36924 , \36182 , \36171 );
nor \U$36548 ( \36925 , \36923 , \36924 );
not \U$36549 ( \36926 , \36925 );
not \U$36550 ( \36927 , \36926 );
not \U$36551 ( \36928 , \10275 );
not \U$36552 ( \36929 , \36109 );
or \U$36553 ( \36930 , \36928 , \36929 );
nand \U$36554 ( \36931 , \36684 , \11205 );
nand \U$36555 ( \36932 , \36930 , \36931 );
not \U$36556 ( \36933 , \36932 );
not \U$36557 ( \36934 , \36933 );
or \U$36558 ( \36935 , \36927 , \36934 );
nand \U$36559 ( \36936 , \36925 , \36932 );
nand \U$36560 ( \36937 , \36935 , \36936 );
not \U$36561 ( \36938 , \36937 );
or \U$36562 ( \36939 , \36920 , \36938 );
nand \U$36563 ( \36940 , \36932 , \36926 );
nand \U$36564 ( \36941 , \36939 , \36940 );
xor \U$36565 ( \36942 , \36913 , \36941 );
xor \U$36566 ( \36943 , \36117 , \36101 );
and \U$36567 ( \36944 , \36942 , \36943 );
and \U$36568 ( \36945 , \36913 , \36941 );
nor \U$36569 ( \36946 , \36944 , \36945 );
not \U$36570 ( \36947 , \36946 );
xor \U$36571 ( \36948 , \36580 , \36499 );
xor \U$36572 ( \36949 , \36948 , \36583 );
not \U$36573 ( \36950 , \36949 );
or \U$36574 ( \36951 , \36947 , \36950 );
or \U$36575 ( \36952 , \36949 , \36946 );
nand \U$36576 ( \36953 , \36951 , \36952 );
not \U$36577 ( \36954 , \36953 );
or \U$36578 ( \36955 , \36836 , \36954 );
not \U$36579 ( \36956 , \36946 );
nand \U$36580 ( \36957 , \36956 , \36949 );
nand \U$36581 ( \36958 , \36955 , \36957 );
not \U$36582 ( \36959 , \36493 );
and \U$36583 ( \36960 , \36598 , \36959 );
not \U$36584 ( \36961 , \36598 );
and \U$36585 ( \36962 , \36961 , \36493 );
nor \U$36586 ( \36963 , \36960 , \36962 );
nand \U$36587 ( \36964 , \36958 , \36963 );
not \U$36588 ( \36965 , \36964 );
xor \U$36589 ( \36966 , \36330 , \36403 );
xnor \U$36590 ( \36967 , \36966 , \36333 );
not \U$36591 ( \36968 , \36478 );
and \U$36592 ( \36969 , \36488 , \36968 );
not \U$36593 ( \36970 , \36488 );
and \U$36594 ( \36971 , \36970 , \36478 );
nor \U$36595 ( \36972 , \36969 , \36971 );
not \U$36596 ( \36973 , \36972 );
nand \U$36597 ( \36974 , \36967 , \36973 );
not \U$36598 ( \36975 , \36335 );
not \U$36599 ( \36976 , \36398 );
not \U$36600 ( \36977 , \36976 );
or \U$36601 ( \36978 , \36975 , \36977 );
or \U$36602 ( \36979 , \36976 , \36335 );
nand \U$36603 ( \36980 , \36978 , \36979 );
xor \U$36604 ( \36981 , \36507 , \36501 );
xor \U$36605 ( \36982 , \36981 , \36578 );
nor \U$36606 ( \36983 , \36980 , \36982 );
not \U$36607 ( \36984 , \36983 );
not \U$36608 ( \36985 , \36982 );
not \U$36609 ( \36986 , \36980 );
or \U$36610 ( \36987 , \36985 , \36986 );
xor \U$36611 ( \36988 , \36574 , \36520 );
not \U$36612 ( \36989 , \36988 );
not \U$36613 ( \36990 , \36989 );
not \U$36614 ( \36991 , \36919 );
and \U$36615 ( \36992 , \36937 , \36991 );
not \U$36616 ( \36993 , \36937 );
and \U$36617 ( \36994 , \36993 , \36919 );
nor \U$36618 ( \36995 , \36992 , \36994 );
not \U$36619 ( \36996 , \36995 );
or \U$36620 ( \36997 , \36990 , \36996 );
and \U$36621 ( \36998 , \36469 , \36445 );
not \U$36622 ( \36999 , \36469 );
and \U$36623 ( \37000 , \36999 , \36446 );
nor \U$36624 ( \37001 , \36998 , \37000 );
nand \U$36625 ( \37002 , \36997 , \37001 );
not \U$36626 ( \37003 , \36995 );
nand \U$36627 ( \37004 , \37003 , \36988 );
and \U$36628 ( \37005 , \37002 , \37004 );
nand \U$36629 ( \37006 , \36987 , \37005 );
nand \U$36630 ( \37007 , \36984 , \37006 );
not \U$36631 ( \37008 , \37007 );
and \U$36632 ( \37009 , \36974 , \37008 );
nor \U$36633 ( \37010 , \36967 , \36973 );
nor \U$36634 ( \37011 , \37009 , \37010 );
not \U$36635 ( \37012 , \37011 );
or \U$36636 ( \37013 , \36965 , \37012 );
nor \U$36637 ( \37014 , \36958 , \36963 );
not \U$36638 ( \37015 , \37014 );
nand \U$36639 ( \37016 , \37013 , \37015 );
not \U$36640 ( \37017 , \37016 );
or \U$36641 ( \37018 , \36642 , \37017 );
or \U$36642 ( \37019 , \37016 , \36641 );
nand \U$36643 ( \37020 , \37018 , \37019 );
not \U$36644 ( \37021 , \37020 );
or \U$36645 ( \37022 , \36633 , \37021 );
not \U$36646 ( \37023 , \36641 );
nand \U$36647 ( \37024 , \37023 , \37016 );
nand \U$36648 ( \37025 , \37022 , \37024 );
nand \U$36649 ( \37026 , \36630 , \37025 );
and \U$36650 ( \37027 , \36305 , \36314 , \36625 , \37026 );
buf \U$36651 ( \37028 , \37027 );
not \U$36652 ( \37029 , \37028 );
not \U$36653 ( \37030 , \9777 );
not \U$36654 ( \37031 , \36708 );
or \U$36655 ( \37032 , \37030 , \37031 );
and \U$36656 ( \37033 , RIae7a150_172, \9290 );
not \U$36657 ( \37034 , RIae7a150_172);
and \U$36658 ( \37035 , \37034 , \14630 );
nor \U$36659 ( \37036 , \37033 , \37035 );
nand \U$36660 ( \37037 , \37036 , \11087 );
nand \U$36661 ( \37038 , \37032 , \37037 );
not \U$36662 ( \37039 , \37038 );
not \U$36663 ( \37040 , \4154 );
and \U$36664 ( \37041 , \10032 , RIae79ca0_162);
not \U$36665 ( \37042 , \10032 );
and \U$36666 ( \37043 , \37042 , \6270 );
nor \U$36667 ( \37044 , \37041 , \37043 );
not \U$36668 ( \37045 , \37044 );
or \U$36669 ( \37046 , \37040 , \37045 );
not \U$36670 ( \37047 , \4852 );
xnor \U$36671 ( \37048 , \10149 , RIae79ca0_162);
nand \U$36672 ( \37049 , \37047 , \37048 );
nand \U$36673 ( \37050 , \37046 , \37049 );
not \U$36674 ( \37051 , \37050 );
or \U$36675 ( \37052 , RIae79700_150, RIae79778_151);
nand \U$36676 ( \37053 , \37052 , \12857 );
nand \U$36677 ( \37054 , \37053 , \4267 );
not \U$36678 ( \37055 , \37054 );
not \U$36679 ( \37056 , \2007 );
not \U$36680 ( \37057 , \18989 );
and \U$36681 ( \37058 , \37057 , \2521 );
not \U$36682 ( \37059 , \37057 );
and \U$36683 ( \37060 , \37059 , RIae797f0_152);
nor \U$36684 ( \37061 , \37058 , \37060 );
not \U$36685 ( \37062 , \37061 );
or \U$36686 ( \37063 , \37056 , \37062 );
xor \U$36687 ( \37064 , \12857 , RIae797f0_152);
nand \U$36688 ( \37065 , \37064 , \1987 );
nand \U$36689 ( \37066 , \37063 , \37065 );
nand \U$36690 ( \37067 , \37055 , \37066 );
not \U$36691 ( \37068 , \37067 );
not \U$36692 ( \37069 , \2418 );
not \U$36693 ( \37070 , \36807 );
or \U$36694 ( \37071 , \37069 , \37070 );
not \U$36695 ( \37072 , RIae79c28_161);
not \U$36696 ( \37073 , \11240 );
or \U$36697 ( \37074 , \37072 , \37073 );
or \U$36698 ( \37075 , \11240 , RIae79c28_161);
nand \U$36699 ( \37076 , \37074 , \37075 );
nand \U$36700 ( \37077 , \37076 , \2417 );
nand \U$36701 ( \37078 , \37071 , \37077 );
not \U$36702 ( \37079 , \37078 );
or \U$36703 ( \37080 , \37068 , \37079 );
or \U$36704 ( \37081 , \37078 , \37067 );
nand \U$36705 ( \37082 , \37080 , \37081 );
not \U$36706 ( \37083 , \37082 );
or \U$36707 ( \37084 , \37051 , \37083 );
not \U$36708 ( \37085 , \37067 );
nand \U$36709 ( \37086 , \37085 , \37078 );
nand \U$36710 ( \37087 , \37084 , \37086 );
not \U$36711 ( \37088 , \10519 );
not \U$36712 ( \37089 , \36822 );
or \U$36713 ( \37090 , \37088 , \37089 );
and \U$36714 ( \37091 , RIae7a7e0_186, \4169 );
not \U$36715 ( \37092 , RIae7a7e0_186);
and \U$36716 ( \37093 , \37092 , \6242 );
nor \U$36717 ( \37094 , \37091 , \37093 );
nand \U$36718 ( \37095 , \37094 , \9549 );
nand \U$36719 ( \37096 , \37090 , \37095 );
xor \U$36720 ( \37097 , \37087 , \37096 );
not \U$36721 ( \37098 , \37097 );
or \U$36722 ( \37099 , \37039 , \37098 );
nand \U$36723 ( \37100 , \37096 , \37087 );
nand \U$36724 ( \37101 , \37099 , \37100 );
not \U$36725 ( \37102 , \37101 );
not \U$36726 ( \37103 , \9622 );
not \U$36727 ( \37104 , \36734 );
or \U$36728 ( \37105 , \37103 , \37104 );
not \U$36729 ( \37106 , \21948 );
not \U$36730 ( \37107 , RIae7a3a8_177);
and \U$36731 ( \37108 , \37106 , \37107 );
and \U$36732 ( \37109 , \13302 , RIae7a3a8_177);
nor \U$36733 ( \37110 , \37108 , \37109 );
not \U$36734 ( \37111 , \37110 );
nand \U$36735 ( \37112 , \37111 , \9644 );
nand \U$36736 ( \37113 , \37105 , \37112 );
not \U$36737 ( \37114 , \9814 );
not \U$36738 ( \37115 , \36776 );
or \U$36739 ( \37116 , \37114 , \37115 );
not \U$36740 ( \37117 , RIae7a2b8_175);
not \U$36741 ( \37118 , \10461 );
or \U$36742 ( \37119 , \37117 , \37118 );
or \U$36743 ( \37120 , \10461 , RIae7a2b8_175);
nand \U$36744 ( \37121 , \37119 , \37120 );
nand \U$36745 ( \37122 , \37121 , \9792 );
nand \U$36746 ( \37123 , \37116 , \37122 );
nor \U$36747 ( \37124 , \37113 , \37123 );
not \U$36748 ( \37125 , \9699 );
not \U$36749 ( \37126 , \36743 );
or \U$36750 ( \37127 , \37125 , \37126 );
not \U$36751 ( \37128 , \11114 );
not \U$36752 ( \37129 , \11198 );
or \U$36753 ( \37130 , \37128 , \37129 );
nand \U$36754 ( \37131 , \11195 , RIae7a240_174);
nand \U$36755 ( \37132 , \37130 , \37131 );
nand \U$36756 ( \37133 , \37132 , \9688 );
nand \U$36757 ( \37134 , \37127 , \37133 );
not \U$36758 ( \37135 , \37134 );
or \U$36759 ( \37136 , \37124 , \37135 );
nand \U$36760 ( \37137 , \37113 , \37123 );
nand \U$36761 ( \37138 , \37136 , \37137 );
xnor \U$36762 ( \37139 , \36846 , \36866 );
xor \U$36763 ( \37140 , \37138 , \37139 );
not \U$36764 ( \37141 , \37140 );
or \U$36765 ( \37142 , \37102 , \37141 );
or \U$36766 ( \37143 , \37101 , \37140 );
nand \U$36767 ( \37144 , \37142 , \37143 );
not \U$36768 ( \37145 , \36686 );
and \U$36769 ( \37146 , \36710 , \36699 );
not \U$36770 ( \37147 , \36710 );
and \U$36771 ( \37148 , \37147 , \36698 );
or \U$36772 ( \37149 , \37146 , \37148 );
not \U$36773 ( \37150 , \37149 );
or \U$36774 ( \37151 , \37145 , \37150 );
or \U$36775 ( \37152 , \37149 , \36686 );
nand \U$36776 ( \37153 , \37151 , \37152 );
not \U$36777 ( \37154 , \36760 );
not \U$36778 ( \37155 , \36736 );
not \U$36779 ( \37156 , \36748 );
or \U$36780 ( \37157 , \37155 , \37156 );
or \U$36781 ( \37158 , \36736 , \36748 );
nand \U$36782 ( \37159 , \37157 , \37158 );
not \U$36783 ( \37160 , \37159 );
or \U$36784 ( \37161 , \37154 , \37160 );
or \U$36785 ( \37162 , \36760 , \37159 );
nand \U$36786 ( \37163 , \37161 , \37162 );
not \U$36787 ( \37164 , \36884 );
not \U$36788 ( \37165 , \36895 );
and \U$36789 ( \37166 , \37164 , \37165 );
and \U$36790 ( \37167 , \36884 , \36895 );
nor \U$36791 ( \37168 , \37166 , \37167 );
xor \U$36792 ( \37169 , \36906 , \37168 );
or \U$36793 ( \37170 , \37163 , \37169 );
nand \U$36794 ( \37171 , \37163 , \37169 );
nand \U$36795 ( \37172 , \37170 , \37171 );
xor \U$36796 ( \37173 , \37153 , \37172 );
xor \U$36797 ( \37174 , \37144 , \37173 );
not \U$36798 ( \37175 , \4853 );
not \U$36799 ( \37176 , \36890 );
or \U$36800 ( \37177 , \37175 , \37176 );
nand \U$36801 ( \37178 , \37048 , \4154 );
nand \U$36802 ( \37179 , \37177 , \37178 );
not \U$36803 ( \37180 , \6214 );
not \U$36804 ( \37181 , \36858 );
or \U$36805 ( \37182 , \37180 , \37181 );
and \U$36806 ( \37183 , RIae79ef8_167, \36201 );
not \U$36807 ( \37184 , RIae79ef8_167);
and \U$36808 ( \37185 , \37184 , \14546 );
or \U$36809 ( \37186 , \37183 , \37185 );
nand \U$36810 ( \37187 , \37186 , \6200 );
nand \U$36811 ( \37188 , \37182 , \37187 );
xor \U$36812 ( \37189 , \37179 , \37188 );
not \U$36813 ( \37190 , \5048 );
not \U$36814 ( \37191 , \36880 );
or \U$36815 ( \37192 , \37190 , \37191 );
and \U$36816 ( \37193 , \10007 , RIae79d90_164);
not \U$36817 ( \37194 , \10007 );
and \U$36818 ( \37195 , \37194 , \4968 );
nor \U$36819 ( \37196 , \37193 , \37195 );
nand \U$36820 ( \37197 , \37196 , \5039 );
nand \U$36821 ( \37198 , \37192 , \37197 );
xor \U$36822 ( \37199 , \37189 , \37198 );
xnor \U$36823 ( \37200 , \36809 , \36798 );
not \U$36824 ( \37201 , \10542 );
not \U$36825 ( \37202 , \36904 );
or \U$36826 ( \37203 , \37201 , \37202 );
and \U$36827 ( \37204 , RIae7a060_170, \24679 );
not \U$36828 ( \37205 , RIae7a060_170);
and \U$36829 ( \37206 , \37205 , \15128 );
nor \U$36830 ( \37207 , \37204 , \37206 );
nand \U$36831 ( \37208 , \37207 , \9730 );
nand \U$36832 ( \37209 , \37203 , \37208 );
xor \U$36833 ( \37210 , \37200 , \37209 );
not \U$36834 ( \37211 , \10631 );
not \U$36835 ( \37212 , \36756 );
or \U$36836 ( \37213 , \37211 , \37212 );
not \U$36837 ( \37214 , \17324 );
not \U$36838 ( \37215 , \15088 );
or \U$36839 ( \37216 , \37214 , \37215 );
not \U$36840 ( \37217 , \15091 );
nand \U$36841 ( \37218 , \37217 , RIae7a510_180);
nand \U$36842 ( \37219 , \37216 , \37218 );
nand \U$36843 ( \37220 , \37219 , \10638 );
nand \U$36844 ( \37221 , \37213 , \37220 );
xnor \U$36845 ( \37222 , \37210 , \37221 );
xor \U$36846 ( \37223 , \37199 , \37222 );
not \U$36847 ( \37224 , \11205 );
and \U$36848 ( \37225 , RIae7a8d0_188, \1860 );
not \U$36849 ( \37226 , RIae7a8d0_188);
and \U$36850 ( \37227 , \37226 , \17596 );
or \U$36851 ( \37228 , \37225 , \37227 );
not \U$36852 ( \37229 , \37228 );
or \U$36853 ( \37230 , \37224 , \37229 );
not \U$36854 ( \37231 , RIae7a8d0_188);
not \U$36855 ( \37232 , \1969 );
or \U$36856 ( \37233 , \37231 , \37232 );
or \U$36857 ( \37234 , \12997 , RIae7a8d0_188);
nand \U$36858 ( \37235 , \37233 , \37234 );
nand \U$36859 ( \37236 , \37235 , \10275 );
nand \U$36860 ( \37237 , \37230 , \37236 );
not \U$36861 ( \37238 , \37237 );
not \U$36862 ( \37239 , RIae7a150_172);
not \U$36863 ( \37240 , \14120 );
or \U$36864 ( \37241 , \37239 , \37240 );
or \U$36865 ( \37242 , \12687 , RIae7a150_172);
nand \U$36866 ( \37243 , \37241 , \37242 );
and \U$36867 ( \37244 , \11087 , \37243 );
and \U$36868 ( \37245 , \37036 , \9776 );
nor \U$36869 ( \37246 , \37244 , \37245 );
not \U$36870 ( \37247 , \37246 );
not \U$36871 ( \37248 , \16564 );
and \U$36872 ( \37249 , RIae7a498_179, \17387 );
not \U$36873 ( \37250 , RIae7a498_179);
and \U$36874 ( \37251 , \37250 , \15519 );
or \U$36875 ( \37252 , \37249 , \37251 );
not \U$36876 ( \37253 , \37252 );
or \U$36877 ( \37254 , \37248 , \37253 );
not \U$36878 ( \37255 , \10625 );
not \U$36879 ( \37256 , \15102 );
or \U$36880 ( \37257 , \37255 , \37256 );
nand \U$36881 ( \37258 , \9313 , RIae7a498_179);
nand \U$36882 ( \37259 , \37257 , \37258 );
nand \U$36883 ( \37260 , \37259 , \10675 );
nand \U$36884 ( \37261 , \37254 , \37260 );
not \U$36885 ( \37262 , \37261 );
or \U$36886 ( \37263 , \37247 , \37262 );
or \U$36887 ( \37264 , \37261 , \37246 );
nand \U$36888 ( \37265 , \37263 , \37264 );
not \U$36889 ( \37266 , \37265 );
or \U$36890 ( \37267 , \37238 , \37266 );
not \U$36891 ( \37268 , \37246 );
nand \U$36892 ( \37269 , \37268 , \37261 );
nand \U$36893 ( \37270 , \37267 , \37269 );
and \U$36894 ( \37271 , \37223 , \37270 );
and \U$36895 ( \37272 , \37199 , \37222 );
or \U$36896 ( \37273 , \37271 , \37272 );
and \U$36897 ( \37274 , \37174 , \37273 );
and \U$36898 ( \37275 , \37144 , \37173 );
or \U$36899 ( \37276 , \37274 , \37275 );
not \U$36900 ( \37277 , \2431 );
not \U$36901 ( \37278 , \2504 );
not \U$36902 ( \37279 , \10272 );
or \U$36903 ( \37280 , \37278 , \37279 );
or \U$36904 ( \37281 , \11321 , \2447 );
nand \U$36905 ( \37282 , \37280 , \37281 );
not \U$36906 ( \37283 , \37282 );
or \U$36907 ( \37284 , \37277 , \37283 );
not \U$36908 ( \37285 , \36558 );
or \U$36909 ( \37286 , \37285 , \18314 );
nand \U$36910 ( \37287 , \37284 , \37286 );
not \U$36911 ( \37288 , \2450 );
not \U$36912 ( \37289 , \37282 );
or \U$36913 ( \37290 , \37288 , \37289 );
and \U$36914 ( \37291 , \10259 , \2504 );
not \U$36915 ( \37292 , \10259 );
and \U$36916 ( \37293 , \37292 , RIae79778_151);
nor \U$36917 ( \37294 , \37291 , \37293 );
nand \U$36918 ( \37295 , \37294 , \2431 );
nand \U$36919 ( \37296 , \37290 , \37295 );
not \U$36920 ( \37297 , \37296 );
and \U$36921 ( \37298 , \12857 , \2321 );
not \U$36922 ( \37299 , \2007 );
not \U$36923 ( \37300 , \36795 );
or \U$36924 ( \37301 , \37299 , \37300 );
nand \U$36925 ( \37302 , \37061 , \1987 );
nand \U$36926 ( \37303 , \37301 , \37302 );
xor \U$36927 ( \37304 , \37298 , \37303 );
not \U$36928 ( \37305 , \37304 );
or \U$36929 ( \37306 , \37297 , \37305 );
nand \U$36930 ( \37307 , \37303 , \37298 );
nand \U$36931 ( \37308 , \37306 , \37307 );
xor \U$36932 ( \37309 , \37287 , \37308 );
not \U$36933 ( \37310 , \37309 );
not \U$36934 ( \37311 , \9518 );
not \U$36935 ( \37312 , \36842 );
or \U$36936 ( \37313 , \37311 , \37312 );
not \U$36937 ( \37314 , RIae79fe8_169);
not \U$36938 ( \37315 , \11387 );
or \U$36939 ( \37316 , \37314 , \37315 );
or \U$36940 ( \37317 , \15653 , RIae79fe8_169);
nand \U$36941 ( \37318 , \37316 , \37317 );
nand \U$36942 ( \37319 , \37318 , \9499 );
nand \U$36943 ( \37320 , \37313 , \37319 );
not \U$36944 ( \37321 , \37320 );
or \U$36945 ( \37322 , \37310 , \37321 );
nand \U$36946 ( \37323 , \37308 , \37287 );
nand \U$36947 ( \37324 , \37322 , \37323 );
not \U$36948 ( \37325 , \37324 );
xor \U$36949 ( \37326 , \37179 , \37188 );
and \U$36950 ( \37327 , \37326 , \37198 );
and \U$36951 ( \37328 , \37179 , \37188 );
or \U$36952 ( \37329 , \37327 , \37328 );
not \U$36953 ( \37330 , \37329 );
nand \U$36954 ( \37331 , \37325 , \37330 );
not \U$36955 ( \37332 , \37331 );
not \U$36956 ( \37333 , \37200 );
not \U$36957 ( \37334 , \37333 );
not \U$36958 ( \37335 , \37221 );
or \U$36959 ( \37336 , \37334 , \37335 );
not \U$36960 ( \37337 , \37209 );
nand \U$36961 ( \37338 , \37336 , \37337 );
not \U$36962 ( \37339 , \37221 );
nand \U$36963 ( \37340 , \37339 , \37200 );
nand \U$36964 ( \37341 , \37338 , \37340 );
not \U$36965 ( \37342 , \37341 );
not \U$36966 ( \37343 , \37342 );
or \U$36967 ( \37344 , \37332 , \37343 );
nand \U$36968 ( \37345 , \37324 , \37329 );
nand \U$36969 ( \37346 , \37344 , \37345 );
xnor \U$36970 ( \37347 , \36906 , \37168 );
not \U$36971 ( \37348 , \37347 );
not \U$36972 ( \37349 , \37163 );
not \U$36973 ( \37350 , \37349 );
or \U$36974 ( \37351 , \37348 , \37350 );
nand \U$36975 ( \37352 , \37351 , \37153 );
and \U$36976 ( \37353 , \37352 , \37171 );
xor \U$36977 ( \37354 , \37346 , \37353 );
not \U$36978 ( \37355 , \37140 );
not \U$36979 ( \37356 , \37355 );
not \U$36980 ( \37357 , \37101 );
or \U$36981 ( \37358 , \37356 , \37357 );
not \U$36982 ( \37359 , \37139 );
nand \U$36983 ( \37360 , \37359 , \37138 );
nand \U$36984 ( \37361 , \37358 , \37360 );
xor \U$36985 ( \37362 , \37354 , \37361 );
xor \U$36986 ( \37363 , \37276 , \37362 );
not \U$36987 ( \37364 , \36671 );
and \U$36988 ( \37365 , \36715 , \37364 );
not \U$36989 ( \37366 , \36715 );
and \U$36990 ( \37367 , \37366 , \36671 );
nor \U$36991 ( \37368 , \37365 , \37367 );
not \U$36992 ( \37369 , \37368 );
xor \U$36993 ( \37370 , \36871 , \36873 );
xor \U$36994 ( \37371 , \37370 , \36910 );
xor \U$36995 ( \37372 , \36764 , \36830 );
not \U$36996 ( \37373 , \36771 );
and \U$36997 ( \37374 , \37372 , \37373 );
not \U$36998 ( \37375 , \37372 );
and \U$36999 ( \37376 , \37375 , \36771 );
nor \U$37000 ( \37377 , \37374 , \37376 );
xnor \U$37001 ( \37378 , \37371 , \37377 );
not \U$37002 ( \37379 , \37378 );
or \U$37003 ( \37380 , \37369 , \37379 );
or \U$37004 ( \37381 , \37378 , \37368 );
nand \U$37005 ( \37382 , \37380 , \37381 );
and \U$37006 ( \37383 , \37363 , \37382 );
and \U$37007 ( \37384 , \37276 , \37362 );
or \U$37008 ( \37385 , \37383 , \37384 );
not \U$37009 ( \37386 , \37385 );
not \U$37010 ( \37387 , \36473 );
and \U$37011 ( \37388 , \36424 , \36476 );
not \U$37012 ( \37389 , \36424 );
and \U$37013 ( \37390 , \37389 , \36434 );
nor \U$37014 ( \37391 , \37388 , \37390 );
not \U$37015 ( \37392 , \37391 );
or \U$37016 ( \37393 , \37387 , \37392 );
or \U$37017 ( \37394 , \37391 , \36473 );
nand \U$37018 ( \37395 , \37393 , \37394 );
and \U$37019 ( \37396 , \36942 , \36943 );
not \U$37020 ( \37397 , \36942 );
not \U$37021 ( \37398 , \36943 );
and \U$37022 ( \37399 , \37397 , \37398 );
nor \U$37023 ( \37400 , \37396 , \37399 );
xor \U$37024 ( \37401 , \37395 , \37400 );
xor \U$37025 ( \37402 , \37346 , \37353 );
and \U$37026 ( \37403 , \37402 , \37361 );
and \U$37027 ( \37404 , \37346 , \37353 );
or \U$37028 ( \37405 , \37403 , \37404 );
xor \U$37029 ( \37406 , \37401 , \37405 );
not \U$37030 ( \37407 , \36780 );
not \U$37031 ( \37408 , \36815 );
or \U$37032 ( \37409 , \37407 , \37408 );
or \U$37033 ( \37410 , \36780 , \36815 );
nand \U$37034 ( \37411 , \37409 , \37410 );
xnor \U$37035 ( \37412 , \36826 , \37411 );
not \U$37036 ( \37413 , \10275 );
not \U$37037 ( \37414 , \36678 );
or \U$37038 ( \37415 , \37413 , \37414 );
nand \U$37039 ( \37416 , \37235 , \16594 );
nand \U$37040 ( \37417 , \37415 , \37416 );
not \U$37041 ( \37418 , \37417 );
not \U$37042 ( \37419 , RIae7aab0_192);
not \U$37043 ( \37420 , \36664 );
or \U$37044 ( \37421 , \37419 , \37420 );
and \U$37045 ( \37422 , RIae7aa38_191, \14439 );
not \U$37046 ( \37423 , RIae7aa38_191);
and \U$37047 ( \37424 , \37423 , \5891 );
or \U$37048 ( \37425 , \37422 , \37424 );
nand \U$37049 ( \37426 , \37425 , \14668 );
nand \U$37050 ( \37427 , \37421 , \37426 );
not \U$37051 ( \37428 , \37427 );
or \U$37052 ( \37429 , \37418 , \37428 );
or \U$37053 ( \37430 , \37427 , \37417 );
not \U$37054 ( \37431 , \11422 );
not \U$37055 ( \37432 , \36694 );
or \U$37056 ( \37433 , \37431 , \37432 );
nand \U$37057 ( \37434 , \37259 , \16564 );
nand \U$37058 ( \37435 , \37433 , \37434 );
nand \U$37059 ( \37436 , \37430 , \37435 );
nand \U$37060 ( \37437 , \37429 , \37436 );
not \U$37061 ( \37438 , \37437 );
xor \U$37062 ( \37439 , \37412 , \37438 );
not \U$37063 ( \37440 , \37320 );
not \U$37064 ( \37441 , \37440 );
not \U$37065 ( \37442 , \37309 );
and \U$37066 ( \37443 , \37441 , \37442 );
and \U$37067 ( \37444 , \37440 , \37309 );
nor \U$37068 ( \37445 , \37443 , \37444 );
not \U$37069 ( \37446 , \17507 );
not \U$37070 ( \37447 , \36648 );
or \U$37071 ( \37448 , \37446 , \37447 );
and \U$37072 ( \37449 , \16101 , \10492 );
not \U$37073 ( \37450 , \16101 );
and \U$37074 ( \37451 , \37450 , \21866 );
nor \U$37075 ( \37452 , \37449 , \37451 );
nand \U$37076 ( \37453 , \37452 , \9473 );
nand \U$37077 ( \37454 , \37448 , \37453 );
not \U$37078 ( \37455 , \37454 );
nand \U$37079 ( \37456 , \37445 , \37455 );
not \U$37080 ( \37457 , \19362 );
and \U$37081 ( \37458 , \10749 , \9560 );
not \U$37082 ( \37459 , \10749 );
and \U$37083 ( \37460 , \37459 , RIae79ef8_167);
nor \U$37084 ( \37461 , \37458 , \37460 );
not \U$37085 ( \37462 , \37461 );
or \U$37086 ( \37463 , \37457 , \37462 );
nand \U$37087 ( \37464 , \37186 , \6212 );
nand \U$37088 ( \37465 , \37463 , \37464 );
not \U$37089 ( \37466 , \37465 );
xnor \U$37090 ( \37467 , \37304 , \37296 );
not \U$37091 ( \37468 , \37467 );
and \U$37092 ( \37469 , \37466 , \37468 );
and \U$37093 ( \37470 , \37465 , \37467 );
nor \U$37094 ( \37471 , \37469 , \37470 );
not \U$37095 ( \37472 , \9792 );
not \U$37096 ( \37473 , \29995 );
not \U$37097 ( \37474 , \16829 );
or \U$37098 ( \37475 , \37473 , \37474 );
or \U$37099 ( \37476 , \12644 , \9799 );
nand \U$37100 ( \37477 , \37475 , \37476 );
not \U$37101 ( \37478 , \37477 );
or \U$37102 ( \37479 , \37472 , \37478 );
nand \U$37103 ( \37480 , \37121 , \9814 );
nand \U$37104 ( \37481 , \37479 , \37480 );
not \U$37105 ( \37482 , \37481 );
or \U$37106 ( \37483 , \37471 , \37482 );
not \U$37107 ( \37484 , \37467 );
nand \U$37108 ( \37485 , \37484 , \37465 );
nand \U$37109 ( \37486 , \37483 , \37485 );
and \U$37110 ( \37487 , \37456 , \37486 );
nor \U$37111 ( \37488 , \37445 , \37455 );
nor \U$37112 ( \37489 , \37487 , \37488 );
and \U$37113 ( \37490 , \37439 , \37489 );
and \U$37114 ( \37491 , \37412 , \37438 );
or \U$37115 ( \37492 , \37490 , \37491 );
not \U$37116 ( \37493 , \37492 );
xor \U$37117 ( \37494 , \36988 , \36995 );
xnor \U$37118 ( \37495 , \37494 , \37001 );
xor \U$37119 ( \37496 , \37493 , \37495 );
not \U$37120 ( \37497 , \37324 );
not \U$37121 ( \37498 , \37330 );
and \U$37122 ( \37499 , \37497 , \37498 );
and \U$37123 ( \37500 , \37324 , \37330 );
nor \U$37124 ( \37501 , \37499 , \37500 );
and \U$37125 ( \37502 , \37341 , \37501 );
not \U$37126 ( \37503 , \37341 );
not \U$37127 ( \37504 , \37501 );
and \U$37128 ( \37505 , \37503 , \37504 );
nor \U$37129 ( \37506 , \37502 , \37505 );
xor \U$37130 ( \37507 , \36643 , \36658 );
xor \U$37131 ( \37508 , \37507 , \36668 );
xor \U$37132 ( \37509 , \37506 , \37508 );
not \U$37133 ( \37510 , \9699 );
not \U$37134 ( \37511 , \37132 );
or \U$37135 ( \37512 , \37510 , \37511 );
not \U$37136 ( \37513 , RIae7a240_174);
not \U$37137 ( \37514 , \12483 );
or \U$37138 ( \37515 , \37513 , \37514 );
or \U$37139 ( \37516 , \29247 , RIae7a240_174);
nand \U$37140 ( \37517 , \37515 , \37516 );
nand \U$37141 ( \37518 , \37517 , \19466 );
nand \U$37142 ( \37519 , \37512 , \37518 );
not \U$37143 ( \37520 , \37519 );
not \U$37144 ( \37521 , \9744 );
not \U$37145 ( \37522 , \37207 );
or \U$37146 ( \37523 , \37521 , \37522 );
not \U$37147 ( \37524 , RIae7a060_170);
not \U$37148 ( \37525 , \12700 );
or \U$37149 ( \37526 , \37524 , \37525 );
or \U$37150 ( \37527 , \13976 , RIae7a060_170);
nand \U$37151 ( \37528 , \37526 , \37527 );
nand \U$37152 ( \37529 , \37528 , \9730 );
nand \U$37153 ( \37530 , \37523 , \37529 );
not \U$37154 ( \37531 , \37530 );
not \U$37155 ( \37532 , \4853 );
not \U$37156 ( \37533 , \37044 );
or \U$37157 ( \37534 , \37532 , \37533 );
not \U$37158 ( \37535 , \10042 );
not \U$37159 ( \37536 , \4844 );
or \U$37160 ( \37537 , \37535 , \37536 );
or \U$37161 ( \37538 , \10042 , \2406 );
nand \U$37162 ( \37539 , \37537 , \37538 );
nand \U$37163 ( \37540 , \37539 , \4842 );
nand \U$37164 ( \37541 , \37534 , \37540 );
xnor \U$37165 ( \37542 , \37054 , \37066 );
not \U$37166 ( \37543 , \2450 );
not \U$37167 ( \37544 , \37294 );
or \U$37168 ( \37545 , \37543 , \37544 );
not \U$37169 ( \37546 , RIae79778_151);
not \U$37170 ( \37547 , \16651 );
or \U$37171 ( \37548 , \37546 , \37547 );
or \U$37172 ( \37549 , \16651 , RIae79778_151);
nand \U$37173 ( \37550 , \37548 , \37549 );
not \U$37174 ( \37551 , \37550 );
or \U$37175 ( \37552 , \37551 , \2430 );
nand \U$37176 ( \37553 , \37545 , \37552 );
xor \U$37177 ( \37554 , \37542 , \37553 );
and \U$37178 ( \37555 , \37541 , \37554 );
and \U$37179 ( \37556 , \37542 , \37553 );
nor \U$37180 ( \37557 , \37555 , \37556 );
nand \U$37181 ( \37558 , \37531 , \37557 );
not \U$37182 ( \37559 , \37558 );
or \U$37183 ( \37560 , \37520 , \37559 );
not \U$37184 ( \37561 , \37557 );
nand \U$37185 ( \37562 , \37561 , \37530 );
nand \U$37186 ( \37563 , \37560 , \37562 );
not \U$37187 ( \37564 , \10631 );
not \U$37188 ( \37565 , \37219 );
or \U$37189 ( \37566 , \37564 , \37565 );
not \U$37190 ( \37567 , \10633 );
not \U$37191 ( \37568 , \12614 );
or \U$37192 ( \37569 , \37567 , \37568 );
or \U$37193 ( \37570 , \12614 , \17324 );
nand \U$37194 ( \37571 , \37569 , \37570 );
nand \U$37195 ( \37572 , \37571 , \11400 );
nand \U$37196 ( \37573 , \37566 , \37572 );
not \U$37197 ( \37574 , \9517 );
not \U$37198 ( \37575 , \37318 );
or \U$37199 ( \37576 , \37574 , \37575 );
not \U$37200 ( \37577 , \11918 );
not \U$37201 ( \37578 , \33735 );
or \U$37202 ( \37579 , \37577 , \37578 );
or \U$37203 ( \37580 , \10066 , \11918 );
nand \U$37204 ( \37581 , \37579 , \37580 );
nand \U$37205 ( \37582 , \37581 , \9499 );
nand \U$37206 ( \37583 , \37576 , \37582 );
not \U$37207 ( \37584 , \37583 );
not \U$37208 ( \37585 , \6091 );
not \U$37209 ( \37586 , RIae79d90_164);
buf \U$37210 ( \37587 , \16193 );
not \U$37211 ( \37588 , \37587 );
or \U$37212 ( \37589 , \37586 , \37588 );
nand \U$37213 ( \37590 , \16194 , \10900 );
nand \U$37214 ( \37591 , \37589 , \37590 );
not \U$37215 ( \37592 , \37591 );
or \U$37216 ( \37593 , \37585 , \37592 );
nand \U$37217 ( \37594 , \37196 , \5048 );
nand \U$37218 ( \37595 , \37593 , \37594 );
not \U$37219 ( \37596 , \37595 );
not \U$37220 ( \37597 , \37596 );
and \U$37221 ( \37598 , \37584 , \37597 );
and \U$37222 ( \37599 , \37583 , \37596 );
nor \U$37223 ( \37600 , \37598 , \37599 );
not \U$37224 ( \37601 , \37600 );
and \U$37225 ( \37602 , \37573 , \37601 );
and \U$37226 ( \37603 , \37583 , \37595 );
nor \U$37227 ( \37604 , \37602 , \37603 );
not \U$37228 ( \37605 , \37604 );
or \U$37229 ( \37606 , \37563 , \37605 );
not \U$37230 ( \37607 , \9473 );
and \U$37231 ( \37608 , RIae7a6f0_184, \5860 );
not \U$37232 ( \37609 , RIae7a6f0_184);
and \U$37233 ( \37610 , \37609 , \24742 );
or \U$37234 ( \37611 , \37608 , \37610 );
not \U$37235 ( \37612 , \37611 );
or \U$37236 ( \37613 , \37607 , \37612 );
nand \U$37237 ( \37614 , \37452 , \17507 );
nand \U$37238 ( \37615 , \37613 , \37614 );
not \U$37239 ( \37616 , \37615 );
not \U$37240 ( \37617 , \37110 );
not \U$37241 ( \37618 , \9621 );
not \U$37242 ( \37619 , \37618 );
and \U$37243 ( \37620 , \37617 , \37619 );
not \U$37244 ( \37621 , RIae7a3a8_177);
not \U$37245 ( \37622 , \29286 );
or \U$37246 ( \37623 , \37621 , \37622 );
or \U$37247 ( \37624 , \9398 , RIae7a3a8_177);
nand \U$37248 ( \37625 , \37623 , \37624 );
and \U$37249 ( \37626 , \37625 , \9644 );
nor \U$37250 ( \37627 , \37620 , \37626 );
not \U$37251 ( \37628 , \37627 );
not \U$37252 ( \37629 , \9549 );
not \U$37253 ( \37630 , RIae7a7e0_186);
not \U$37254 ( \37631 , \10829 );
or \U$37255 ( \37632 , \37630 , \37631 );
or \U$37256 ( \37633 , \10829 , RIae7a7e0_186);
nand \U$37257 ( \37634 , \37632 , \37633 );
not \U$37258 ( \37635 , \37634 );
or \U$37259 ( \37636 , \37629 , \37635 );
nand \U$37260 ( \37637 , \37094 , \29519 );
nand \U$37261 ( \37638 , \37636 , \37637 );
not \U$37262 ( \37639 , \37638 );
or \U$37263 ( \37640 , \37628 , \37639 );
or \U$37264 ( \37641 , \37638 , \37627 );
nand \U$37265 ( \37642 , \37640 , \37641 );
not \U$37266 ( \37643 , \37642 );
or \U$37267 ( \37644 , \37616 , \37643 );
not \U$37268 ( \37645 , \37627 );
nand \U$37269 ( \37646 , \37645 , \37638 );
nand \U$37270 ( \37647 , \37644 , \37646 );
nand \U$37271 ( \37648 , \37606 , \37647 );
nand \U$37272 ( \37649 , \37563 , \37605 );
nand \U$37273 ( \37650 , \37648 , \37649 );
and \U$37274 ( \37651 , \37509 , \37650 );
and \U$37275 ( \37652 , \37506 , \37508 );
or \U$37276 ( \37653 , \37651 , \37652 );
and \U$37277 ( \37654 , \37496 , \37653 );
and \U$37278 ( \37655 , \37493 , \37495 );
or \U$37279 ( \37656 , \37654 , \37655 );
nand \U$37280 ( \37657 , \37406 , \37656 );
not \U$37281 ( \37658 , \37657 );
not \U$37282 ( \37659 , \37658 );
and \U$37283 ( \37660 , \37386 , \37659 );
not \U$37284 ( \37661 , \37406 );
not \U$37285 ( \37662 , \37656 );
nand \U$37286 ( \37663 , \37661 , \37662 );
not \U$37287 ( \37664 , \37663 );
nor \U$37288 ( \37665 , \37660 , \37664 );
not \U$37289 ( \37666 , \37665 );
not \U$37290 ( \37667 , \37666 );
xnor \U$37291 ( \37668 , \36972 , \37007 );
not \U$37292 ( \37669 , \37668 );
not \U$37293 ( \37670 , \36967 );
not \U$37294 ( \37671 , \37670 );
and \U$37295 ( \37672 , \37669 , \37671 );
and \U$37296 ( \37673 , \37668 , \37670 );
nor \U$37297 ( \37674 , \37672 , \37673 );
xor \U$37298 ( \37675 , \37395 , \37400 );
and \U$37299 ( \37676 , \37675 , \37405 );
and \U$37300 ( \37677 , \37395 , \37400 );
or \U$37301 ( \37678 , \37676 , \37677 );
not \U$37302 ( \37679 , \37678 );
not \U$37303 ( \37680 , \36835 );
not \U$37304 ( \37681 , \36953 );
not \U$37305 ( \37682 , \37681 );
or \U$37306 ( \37683 , \37680 , \37682 );
not \U$37307 ( \37684 , \36835 );
nand \U$37308 ( \37685 , \36953 , \37684 );
nand \U$37309 ( \37686 , \37683 , \37685 );
not \U$37310 ( \37687 , \37686 );
not \U$37311 ( \37688 , \37687 );
or \U$37312 ( \37689 , \37679 , \37688 );
not \U$37313 ( \37690 , \37678 );
nand \U$37314 ( \37691 , \37686 , \37690 );
nand \U$37315 ( \37692 , \37689 , \37691 );
not \U$37316 ( \37693 , \37368 );
not \U$37317 ( \37694 , \37693 );
not \U$37318 ( \37695 , \37378 );
or \U$37319 ( \37696 , \37694 , \37695 );
not \U$37320 ( \37697 , \37377 );
nand \U$37321 ( \37698 , \37697 , \37371 );
nand \U$37322 ( \37699 , \37696 , \37698 );
not \U$37323 ( \37700 , \37699 );
xor \U$37324 ( \37701 , \36724 , \36832 );
xor \U$37325 ( \37702 , \37701 , \36719 );
not \U$37326 ( \37703 , \37702 );
not \U$37327 ( \37704 , \37703 );
or \U$37328 ( \37705 , \37700 , \37704 );
not \U$37329 ( \37706 , \37702 );
not \U$37330 ( \37707 , \37699 );
not \U$37331 ( \37708 , \37707 );
or \U$37332 ( \37709 , \37706 , \37708 );
not \U$37333 ( \37710 , \37005 );
not \U$37334 ( \37711 , \37710 );
not \U$37335 ( \37712 , \36983 );
nand \U$37336 ( \37713 , \36980 , \36982 );
nand \U$37337 ( \37714 , \37712 , \37713 );
not \U$37338 ( \37715 , \37714 );
or \U$37339 ( \37716 , \37711 , \37715 );
or \U$37340 ( \37717 , \37714 , \37710 );
nand \U$37341 ( \37718 , \37716 , \37717 );
nand \U$37342 ( \37719 , \37709 , \37718 );
nand \U$37343 ( \37720 , \37705 , \37719 );
and \U$37344 ( \37721 , \37692 , \37720 );
not \U$37345 ( \37722 , \37692 );
not \U$37346 ( \37723 , \37720 );
and \U$37347 ( \37724 , \37722 , \37723 );
nor \U$37348 ( \37725 , \37721 , \37724 );
and \U$37349 ( \37726 , \37674 , \37725 );
not \U$37350 ( \37727 , \37674 );
not \U$37351 ( \37728 , \37725 );
and \U$37352 ( \37729 , \37727 , \37728 );
nor \U$37353 ( \37730 , \37726 , \37729 );
not \U$37354 ( \37731 , \37730 );
or \U$37355 ( \37732 , \37667 , \37731 );
not \U$37356 ( \37733 , \37674 );
nand \U$37357 ( \37734 , \37733 , \37728 );
nand \U$37358 ( \37735 , \37732 , \37734 );
xor \U$37359 ( \37736 , \36414 , \36408 );
xnor \U$37360 ( \37737 , \37736 , \36418 );
not \U$37361 ( \37738 , \37690 );
not \U$37362 ( \37739 , \37687 );
or \U$37363 ( \37740 , \37738 , \37739 );
nand \U$37364 ( \37741 , \37740 , \37720 );
nand \U$37365 ( \37742 , \37686 , \37678 );
and \U$37366 ( \37743 , \37741 , \37742 );
xor \U$37367 ( \37744 , \37737 , \37743 );
not \U$37368 ( \37745 , \37014 );
nand \U$37369 ( \37746 , \37745 , \36964 );
not \U$37370 ( \37747 , \37011 );
and \U$37371 ( \37748 , \37746 , \37747 );
not \U$37372 ( \37749 , \37746 );
and \U$37373 ( \37750 , \37749 , \37011 );
nor \U$37374 ( \37751 , \37748 , \37750 );
xor \U$37375 ( \37752 , \37744 , \37751 );
nand \U$37376 ( \37753 , \37735 , \37752 );
not \U$37377 ( \37754 , \36631 );
not \U$37378 ( \37755 , \37020 );
or \U$37379 ( \37756 , \37754 , \37755 );
or \U$37380 ( \37757 , \37020 , \36631 );
nand \U$37381 ( \37758 , \37756 , \37757 );
xor \U$37382 ( \37759 , \37737 , \37743 );
and \U$37383 ( \37760 , \37759 , \37751 );
and \U$37384 ( \37761 , \37737 , \37743 );
or \U$37385 ( \37762 , \37760 , \37761 );
nand \U$37386 ( \37763 , \37758 , \37762 );
xor \U$37387 ( \37764 , \37674 , \37665 );
xnor \U$37388 ( \37765 , \37764 , \37725 );
and \U$37389 ( \37766 , \37707 , \37702 );
not \U$37390 ( \37767 , \37707 );
and \U$37391 ( \37768 , \37767 , \37703 );
nor \U$37392 ( \37769 , \37766 , \37768 );
not \U$37393 ( \37770 , \37718 );
and \U$37394 ( \37771 , \37769 , \37770 );
not \U$37395 ( \37772 , \37769 );
and \U$37396 ( \37773 , \37772 , \37718 );
nor \U$37397 ( \37774 , \37771 , \37773 );
nand \U$37398 ( \37775 , \37657 , \37663 );
not \U$37399 ( \37776 , \37775 );
not \U$37400 ( \37777 , \37385 );
and \U$37401 ( \37778 , \37776 , \37777 );
and \U$37402 ( \37779 , \37775 , \37385 );
nor \U$37403 ( \37780 , \37778 , \37779 );
xor \U$37404 ( \37781 , \37774 , \37780 );
xor \U$37405 ( \37782 , \37493 , \37495 );
xor \U$37406 ( \37783 , \37782 , \37653 );
not \U$37407 ( \37784 , \37783 );
xor \U$37408 ( \37785 , \37435 , \37417 );
xnor \U$37409 ( \37786 , \37785 , \37427 );
not \U$37410 ( \37787 , \37786 );
not \U$37411 ( \37788 , \37787 );
not \U$37412 ( \37789 , \37124 );
nand \U$37413 ( \37790 , \37789 , \37137 );
and \U$37414 ( \37791 , \37790 , \37134 );
not \U$37415 ( \37792 , \37790 );
and \U$37416 ( \37793 , \37792 , \37135 );
nor \U$37417 ( \37794 , \37791 , \37793 );
not \U$37418 ( \37795 , \37794 );
not \U$37419 ( \37796 , \37795 );
or \U$37420 ( \37797 , \37788 , \37796 );
not \U$37421 ( \37798 , \37786 );
not \U$37422 ( \37799 , \37794 );
or \U$37423 ( \37800 , \37798 , \37799 );
xor \U$37424 ( \37801 , \37087 , \37038 );
xor \U$37425 ( \37802 , \37801 , \37096 );
nand \U$37426 ( \37803 , \37800 , \37802 );
nand \U$37427 ( \37804 , \37797 , \37803 );
not \U$37428 ( \37805 , \37804 );
xor \U$37429 ( \37806 , \37412 , \37438 );
xor \U$37430 ( \37807 , \37806 , \37489 );
nand \U$37431 ( \37808 , \37805 , \37807 );
not \U$37432 ( \37809 , \37808 );
not \U$37433 ( \37810 , \6091 );
and \U$37434 ( \37811 , \33414 , \4968 );
not \U$37435 ( \37812 , \33414 );
and \U$37436 ( \37813 , \37812 , RIae79d90_164);
nor \U$37437 ( \37814 , \37811 , \37813 );
not \U$37438 ( \37815 , \37814 );
or \U$37439 ( \37816 , \37810 , \37815 );
not \U$37440 ( \37817 , \10142 );
not \U$37441 ( \37818 , RIae79d90_164);
and \U$37442 ( \37819 , \37817 , \37818 );
and \U$37443 ( \37820 , \10142 , RIae79d90_164);
nor \U$37444 ( \37821 , \37819 , \37820 );
nand \U$37445 ( \37822 , \37821 , \5048 );
nand \U$37446 ( \37823 , \37816 , \37822 );
not \U$37447 ( \37824 , \37823 );
or \U$37448 ( \37825 , RIae79bb0_160, RIae79c28_161);
nand \U$37449 ( \37826 , \37825 , \12857 );
nand \U$37450 ( \37827 , \37826 , \2505 );
not \U$37451 ( \37828 , \37827 );
not \U$37452 ( \37829 , \2450 );
not \U$37453 ( \37830 , RIae79778_151);
not \U$37454 ( \37831 , \16005 );
or \U$37455 ( \37832 , \37830 , \37831 );
or \U$37456 ( \37833 , \12750 , RIae79778_151);
nand \U$37457 ( \37834 , \37832 , \37833 );
not \U$37458 ( \37835 , \37834 );
or \U$37459 ( \37836 , \37829 , \37835 );
not \U$37460 ( \37837 , RIae79778_151);
not \U$37461 ( \37838 , \14601 );
or \U$37462 ( \37839 , \37837 , \37838 );
or \U$37463 ( \37840 , \17971 , RIae79778_151);
nand \U$37464 ( \37841 , \37839 , \37840 );
nand \U$37465 ( \37842 , \37841 , \2431 );
nand \U$37466 ( \37843 , \37836 , \37842 );
nand \U$37467 ( \37844 , \37828 , \37843 );
not \U$37468 ( \37845 , \37844 );
not \U$37469 ( \37846 , \4155 );
not \U$37470 ( \37847 , \37539 );
or \U$37471 ( \37848 , \37846 , \37847 );
and \U$37472 ( \37849 , RIae79ca0_162, \11581 );
not \U$37473 ( \37850 , RIae79ca0_162);
and \U$37474 ( \37851 , \37850 , \32565 );
or \U$37475 ( \37852 , \37849 , \37851 );
nand \U$37476 ( \37853 , \37852 , \4154 );
nand \U$37477 ( \37854 , \37848 , \37853 );
not \U$37478 ( \37855 , \37854 );
or \U$37479 ( \37856 , \37845 , \37855 );
or \U$37480 ( \37857 , \37854 , \37844 );
nand \U$37481 ( \37858 , \37856 , \37857 );
not \U$37482 ( \37859 , \37858 );
or \U$37483 ( \37860 , \37824 , \37859 );
not \U$37484 ( \37861 , \37844 );
nand \U$37485 ( \37862 , \37861 , \37854 );
nand \U$37486 ( \37863 , \37860 , \37862 );
not \U$37487 ( \37864 , \37863 );
not \U$37488 ( \37865 , \37864 );
not \U$37489 ( \37866 , \9730 );
not \U$37490 ( \37867 , RIae7a060_170);
not \U$37491 ( \37868 , \9286 );
or \U$37492 ( \37869 , \37867 , \37868 );
nand \U$37493 ( \37870 , \6345 , \9749 );
nand \U$37494 ( \37871 , \37869 , \37870 );
not \U$37495 ( \37872 , \37871 );
or \U$37496 ( \37873 , \37866 , \37872 );
nand \U$37497 ( \37874 , \37528 , \10542 );
nand \U$37498 ( \37875 , \37873 , \37874 );
not \U$37499 ( \37876 , \37875 );
not \U$37500 ( \37877 , \37876 );
or \U$37501 ( \37878 , \37865 , \37877 );
not \U$37502 ( \37879 , \9776 );
not \U$37503 ( \37880 , \37243 );
or \U$37504 ( \37881 , \37879 , \37880 );
and \U$37505 ( \37882 , \15102 , RIae7a150_172);
not \U$37506 ( \37883 , \15102 );
and \U$37507 ( \37884 , \37883 , \10672 );
nor \U$37508 ( \37885 , \37882 , \37884 );
nand \U$37509 ( \37886 , \37885 , \10667 );
nand \U$37510 ( \37887 , \37881 , \37886 );
nand \U$37511 ( \37888 , \37878 , \37887 );
nand \U$37512 ( \37889 , \37875 , \37863 );
nand \U$37513 ( \37890 , \37888 , \37889 );
not \U$37514 ( \37891 , \37890 );
and \U$37515 ( \37892 , \37471 , \37481 );
not \U$37516 ( \37893 , \37471 );
and \U$37517 ( \37894 , \37893 , \37482 );
nor \U$37518 ( \37895 , \37892 , \37894 );
not \U$37519 ( \37896 , \37895 );
not \U$37520 ( \37897 , \37600 );
not \U$37521 ( \37898 , \37573 );
or \U$37522 ( \37899 , \37897 , \37898 );
or \U$37523 ( \37900 , \37573 , \37600 );
nand \U$37524 ( \37901 , \37899 , \37900 );
not \U$37525 ( \37902 , \37901 );
or \U$37526 ( \37903 , \37896 , \37902 );
or \U$37527 ( \37904 , \37901 , \37895 );
nand \U$37528 ( \37905 , \37903 , \37904 );
not \U$37529 ( \37906 , \37905 );
or \U$37530 ( \37907 , \37891 , \37906 );
not \U$37531 ( \37908 , \37895 );
nand \U$37532 ( \37909 , \37908 , \37901 );
nand \U$37533 ( \37910 , \37907 , \37909 );
not \U$37534 ( \37911 , \37910 );
not \U$37535 ( \37912 , \16383 );
and \U$37536 ( \37913 , \5115 , RIae7aa38_191);
not \U$37537 ( \37914 , \5115 );
and \U$37538 ( \37915 , \37914 , \11326 );
nor \U$37539 ( \37916 , \37913 , \37915 );
not \U$37540 ( \37917 , \37916 );
or \U$37541 ( \37918 , \37912 , \37917 );
nand \U$37542 ( \37919 , \37425 , RIae7aab0_192);
nand \U$37543 ( \37920 , \37918 , \37919 );
not \U$37544 ( \37921 , \37920 );
not \U$37545 ( \37922 , \37050 );
not \U$37546 ( \37923 , \37922 );
not \U$37547 ( \37924 , \37082 );
or \U$37548 ( \37925 , \37923 , \37924 );
or \U$37549 ( \37926 , \37082 , \37922 );
nand \U$37550 ( \37927 , \37925 , \37926 );
not \U$37551 ( \37928 , \37927 );
not \U$37552 ( \37929 , \2418 );
not \U$37553 ( \37930 , \37076 );
or \U$37554 ( \37931 , \37929 , \37930 );
not \U$37555 ( \37932 , \10584 );
not \U$37556 ( \37933 , \11321 );
or \U$37557 ( \37934 , \37932 , \37933 );
or \U$37558 ( \37935 , \28259 , \10584 );
nand \U$37559 ( \37936 , \37934 , \37935 );
nand \U$37560 ( \37937 , \37936 , \2417 );
nand \U$37561 ( \37938 , \37931 , \37937 );
not \U$37562 ( \37939 , \37938 );
and \U$37563 ( \37940 , \12857 , \2007 );
not \U$37564 ( \37941 , \2431 );
not \U$37565 ( \37942 , \37834 );
or \U$37566 ( \37943 , \37941 , \37942 );
nand \U$37567 ( \37944 , \37550 , \2450 );
nand \U$37568 ( \37945 , \37943 , \37944 );
xor \U$37569 ( \37946 , \37940 , \37945 );
not \U$37570 ( \37947 , \2418 );
not \U$37571 ( \37948 , \37936 );
or \U$37572 ( \37949 , \37947 , \37948 );
not \U$37573 ( \37950 , RIae79c28_161);
not \U$37574 ( \37951 , \10259 );
or \U$37575 ( \37952 , \37950 , \37951 );
or \U$37576 ( \37953 , \10259 , RIae79c28_161);
nand \U$37577 ( \37954 , \37952 , \37953 );
nand \U$37578 ( \37955 , \37954 , \2417 );
nand \U$37579 ( \37956 , \37949 , \37955 );
and \U$37580 ( \37957 , \37946 , \37956 );
and \U$37581 ( \37958 , \37940 , \37945 );
nor \U$37582 ( \37959 , \37957 , \37958 );
not \U$37583 ( \37960 , \37959 );
or \U$37584 ( \37961 , \37939 , \37960 );
or \U$37585 ( \37962 , \37938 , \37959 );
nand \U$37586 ( \37963 , \37961 , \37962 );
not \U$37587 ( \37964 , \16135 );
not \U$37588 ( \37965 , \37477 );
or \U$37589 ( \37966 , \37964 , \37965 );
and \U$37590 ( \37967 , RIae7a2b8_175, \19025 );
not \U$37591 ( \37968 , RIae7a2b8_175);
and \U$37592 ( \37969 , \37968 , \10084 );
nor \U$37593 ( \37970 , \37967 , \37969 );
nand \U$37594 ( \37971 , \37970 , \9792 );
nand \U$37595 ( \37972 , \37966 , \37971 );
and \U$37596 ( \37973 , \37963 , \37972 );
not \U$37597 ( \37974 , \37938 );
nor \U$37598 ( \37975 , \37974 , \37959 );
nor \U$37599 ( \37976 , \37973 , \37975 );
not \U$37600 ( \37977 , \37976 );
or \U$37601 ( \37978 , \37928 , \37977 );
or \U$37602 ( \37979 , \37976 , \37927 );
nand \U$37603 ( \37980 , \37978 , \37979 );
not \U$37604 ( \37981 , \37980 );
or \U$37605 ( \37982 , \37921 , \37981 );
not \U$37606 ( \37983 , \37976 );
nand \U$37607 ( \37984 , \37983 , \37927 );
nand \U$37608 ( \37985 , \37982 , \37984 );
not \U$37609 ( \37986 , \37985 );
not \U$37610 ( \37987 , \37986 );
xnor \U$37611 ( \37988 , \37554 , \37541 );
not \U$37612 ( \37989 , \37988 );
not \U$37613 ( \37990 , \12233 );
not \U$37614 ( \37991 , \37571 );
or \U$37615 ( \37992 , \37990 , \37991 );
and \U$37616 ( \37993 , RIae7a510_180, \14657 );
not \U$37617 ( \37994 , RIae7a510_180);
and \U$37618 ( \37995 , \37994 , \19736 );
or \U$37619 ( \37996 , \37993 , \37995 );
nand \U$37620 ( \37997 , \37996 , \10638 );
nand \U$37621 ( \37998 , \37992 , \37997 );
not \U$37622 ( \37999 , \37998 );
or \U$37623 ( \38000 , \37989 , \37999 );
or \U$37624 ( \38001 , \37998 , \37988 );
nand \U$37625 ( \38002 , \38000 , \38001 );
not \U$37626 ( \38003 , \38002 );
not \U$37627 ( \38004 , \9705 );
not \U$37628 ( \38005 , \37611 );
or \U$37629 ( \38006 , \38004 , \38005 );
not \U$37630 ( \38007 , \16101 );
not \U$37631 ( \38008 , \4169 );
or \U$37632 ( \38009 , \38007 , \38008 );
nand \U$37633 ( \38010 , \21873 , RIae7a6f0_184);
nand \U$37634 ( \38011 , \38009 , \38010 );
nand \U$37635 ( \38012 , \38011 , \9473 );
nand \U$37636 ( \38013 , \38006 , \38012 );
not \U$37637 ( \38014 , \38013 );
or \U$37638 ( \38015 , \38003 , \38014 );
not \U$37639 ( \38016 , \37988 );
nand \U$37640 ( \38017 , \38016 , \37998 );
nand \U$37641 ( \38018 , \38015 , \38017 );
not \U$37642 ( \38019 , \38018 );
and \U$37643 ( \38020 , \37591 , \5048 );
and \U$37644 ( \38021 , \37821 , \6091 );
nor \U$37645 ( \38022 , \38020 , \38021 );
not \U$37646 ( \38023 , \38022 );
not \U$37647 ( \38024 , \38023 );
not \U$37648 ( \38025 , \9517 );
not \U$37649 ( \38026 , \37581 );
or \U$37650 ( \38027 , \38025 , \38026 );
not \U$37651 ( \38028 , RIae79fe8_169);
not \U$37652 ( \38029 , \9897 );
or \U$37653 ( \38030 , \38028 , \38029 );
or \U$37654 ( \38031 , \9897 , RIae79fe8_169);
nand \U$37655 ( \38032 , \38030 , \38031 );
nand \U$37656 ( \38033 , \38032 , \9499 );
nand \U$37657 ( \38034 , \38027 , \38033 );
not \U$37658 ( \38035 , \6212 );
not \U$37659 ( \38036 , \37461 );
or \U$37660 ( \38037 , \38035 , \38036 );
xnor \U$37661 ( \38038 , \10000 , RIae79ef8_167);
nand \U$37662 ( \38039 , \38038 , \19362 );
nand \U$37663 ( \38040 , \38037 , \38039 );
xor \U$37664 ( \38041 , \38034 , \38040 );
not \U$37665 ( \38042 , \38041 );
or \U$37666 ( \38043 , \38024 , \38042 );
nand \U$37667 ( \38044 , \38040 , \38034 );
nand \U$37668 ( \38045 , \38043 , \38044 );
not \U$37669 ( \38046 , \38045 );
not \U$37670 ( \38047 , \9621 );
not \U$37671 ( \38048 , \37625 );
or \U$37672 ( \38049 , \38047 , \38048 );
not \U$37673 ( \38050 , RIae7a3a8_177);
not \U$37674 ( \38051 , \9412 );
or \U$37675 ( \38052 , \38050 , \38051 );
or \U$37676 ( \38053 , \9417 , RIae7a3a8_177);
nand \U$37677 ( \38054 , \38052 , \38053 );
nand \U$37678 ( \38055 , \11013 , \38054 );
nand \U$37679 ( \38056 , \38049 , \38055 );
not \U$37680 ( \38057 , \38056 );
not \U$37681 ( \38058 , \9699 );
not \U$37682 ( \38059 , \37517 );
or \U$37683 ( \38060 , \38058 , \38059 );
not \U$37684 ( \38061 , RIae7a240_174);
not \U$37685 ( \38062 , \9941 );
or \U$37686 ( \38063 , \38061 , \38062 );
not \U$37687 ( \38064 , RIae7a240_174);
nand \U$37688 ( \38065 , \11186 , \38064 );
nand \U$37689 ( \38066 , \38063 , \38065 );
nand \U$37690 ( \38067 , \38066 , \19466 );
nand \U$37691 ( \38068 , \38060 , \38067 );
not \U$37692 ( \38069 , \38068 );
nand \U$37693 ( \38070 , \38057 , \38069 );
not \U$37694 ( \38071 , \29519 );
not \U$37695 ( \38072 , \37634 );
or \U$37696 ( \38073 , \38071 , \38072 );
and \U$37697 ( \38074 , RIae7a7e0_186, \5108 );
not \U$37698 ( \38075 , RIae7a7e0_186);
and \U$37699 ( \38076 , \38075 , \6256 );
or \U$37700 ( \38077 , \38074 , \38076 );
nand \U$37701 ( \38078 , \38077 , \9549 );
nand \U$37702 ( \38079 , \38073 , \38078 );
nand \U$37703 ( \38080 , \38070 , \38079 );
nand \U$37704 ( \38081 , \38056 , \38068 );
and \U$37705 ( \38082 , \38080 , \38081 );
not \U$37706 ( \38083 , \38082 );
or \U$37707 ( \38084 , \38046 , \38083 );
not \U$37708 ( \38085 , \38081 );
not \U$37709 ( \38086 , \38080 );
or \U$37710 ( \38087 , \38085 , \38086 );
not \U$37711 ( \38088 , \38045 );
nand \U$37712 ( \38089 , \38087 , \38088 );
nand \U$37713 ( \38090 , \38084 , \38089 );
not \U$37714 ( \38091 , \38090 );
or \U$37715 ( \38092 , \38019 , \38091 );
not \U$37716 ( \38093 , \38081 );
not \U$37717 ( \38094 , \38080 );
or \U$37718 ( \38095 , \38093 , \38094 );
nand \U$37719 ( \38096 , \38095 , \38045 );
nand \U$37720 ( \38097 , \38092 , \38096 );
not \U$37721 ( \38098 , \38097 );
or \U$37722 ( \38099 , \37987 , \38098 );
or \U$37723 ( \38100 , \38097 , \37986 );
nand \U$37724 ( \38101 , \38099 , \38100 );
not \U$37725 ( \38102 , \38101 );
or \U$37726 ( \38103 , \37911 , \38102 );
buf \U$37727 ( \38104 , \38097 );
nand \U$37728 ( \38105 , \38104 , \37985 );
nand \U$37729 ( \38106 , \38103 , \38105 );
not \U$37730 ( \38107 , \38106 );
or \U$37731 ( \38108 , \37809 , \38107 );
not \U$37732 ( \38109 , \37807 );
nand \U$37733 ( \38110 , \38109 , \37804 );
nand \U$37734 ( \38111 , \38108 , \38110 );
not \U$37735 ( \38112 , \38111 );
not \U$37736 ( \38113 , \38112 );
and \U$37737 ( \38114 , \37784 , \38113 );
and \U$37738 ( \38115 , \37783 , \38112 );
nor \U$37739 ( \38116 , \38114 , \38115 );
not \U$37740 ( \38117 , \38116 );
xor \U$37741 ( \38118 , \37506 , \37508 );
xor \U$37742 ( \38119 , \38118 , \37650 );
xor \U$37743 ( \38120 , \37144 , \37173 );
xor \U$37744 ( \38121 , \38120 , \37273 );
xor \U$37745 ( \38122 , \38119 , \38121 );
not \U$37746 ( \38123 , \10275 );
not \U$37747 ( \38124 , \37228 );
or \U$37748 ( \38125 , \38123 , \38124 );
and \U$37749 ( \38126 , RIae7a8d0_188, \2403 );
not \U$37750 ( \38127 , RIae7a8d0_188);
and \U$37751 ( \38128 , \38127 , \5673 );
or \U$37752 ( \38129 , \38126 , \38128 );
nand \U$37753 ( \38130 , \38129 , \17847 );
nand \U$37754 ( \38131 , \38125 , \38130 );
not \U$37755 ( \38132 , \38131 );
not \U$37756 ( \38133 , \10676 );
not \U$37757 ( \38134 , \37252 );
or \U$37758 ( \38135 , \38133 , \38134 );
xor \U$37759 ( \38136 , RIae7a498_179, \15088 );
nand \U$37760 ( \38137 , \38136 , \16564 );
nand \U$37761 ( \38138 , \38135 , \38137 );
not \U$37762 ( \38139 , \38138 );
not \U$37763 ( \38140 , \38139 );
or \U$37764 ( \38141 , \38132 , \38140 );
or \U$37765 ( \38142 , \38139 , \38131 );
nand \U$37766 ( \38143 , \38141 , \38142 );
not \U$37767 ( \38144 , RIae7aab0_192);
not \U$37768 ( \38145 , \37916 );
or \U$37769 ( \38146 , \38144 , \38145 );
and \U$37770 ( \38147 , \23255 , \11326 );
not \U$37771 ( \38148 , \23255 );
and \U$37772 ( \38149 , \38148 , RIae7aa38_191);
nor \U$37773 ( \38150 , \38147 , \38149 );
nand \U$37774 ( \38151 , \38150 , \14668 );
nand \U$37775 ( \38152 , \38146 , \38151 );
and \U$37776 ( \38153 , \38143 , \38152 );
and \U$37777 ( \38154 , \38138 , \38131 );
nor \U$37778 ( \38155 , \38153 , \38154 );
not \U$37779 ( \38156 , \38155 );
not \U$37780 ( \38157 , \38156 );
not \U$37781 ( \38158 , \37615 );
not \U$37782 ( \38159 , \38158 );
not \U$37783 ( \38160 , \37642 );
or \U$37784 ( \38161 , \38159 , \38160 );
or \U$37785 ( \38162 , \37642 , \38158 );
nand \U$37786 ( \38163 , \38161 , \38162 );
not \U$37787 ( \38164 , \37237 );
not \U$37788 ( \38165 , \38164 );
not \U$37789 ( \38166 , \37265 );
or \U$37790 ( \38167 , \38165 , \38166 );
or \U$37791 ( \38168 , \37265 , \38164 );
nand \U$37792 ( \38169 , \38167 , \38168 );
xor \U$37793 ( \38170 , \38163 , \38169 );
not \U$37794 ( \38171 , \38170 );
or \U$37795 ( \38172 , \38157 , \38171 );
nand \U$37796 ( \38173 , \38163 , \38169 );
nand \U$37797 ( \38174 , \38172 , \38173 );
xor \U$37798 ( \38175 , \37454 , \37445 );
xnor \U$37799 ( \38176 , \38175 , \37486 );
xor \U$37800 ( \38177 , \38174 , \38176 );
xor \U$37801 ( \38178 , \37604 , \37563 );
xor \U$37802 ( \38179 , \38178 , \37647 );
not \U$37803 ( \38180 , \38179 );
and \U$37804 ( \38181 , \38177 , \38180 );
and \U$37805 ( \38182 , \38174 , \38176 );
or \U$37806 ( \38183 , \38181 , \38182 );
and \U$37807 ( \38184 , \38122 , \38183 );
and \U$37808 ( \38185 , \38119 , \38121 );
or \U$37809 ( \38186 , \38184 , \38185 );
and \U$37810 ( \38187 , \38117 , \38186 );
not \U$37811 ( \38188 , \37783 );
nor \U$37812 ( \38189 , \38188 , \38112 );
nor \U$37813 ( \38190 , \38187 , \38189 );
and \U$37814 ( \38191 , \37781 , \38190 );
and \U$37815 ( \38192 , \37774 , \37780 );
or \U$37816 ( \38193 , \38191 , \38192 );
nand \U$37817 ( \38194 , \37765 , \38193 );
xor \U$37818 ( \38195 , \37774 , \37780 );
xor \U$37819 ( \38196 , \38195 , \38190 );
xor \U$37820 ( \38197 , \37276 , \37362 );
xor \U$37821 ( \38198 , \38197 , \37382 );
not \U$37822 ( \38199 , \38106 );
not \U$37823 ( \38200 , \37804 );
not \U$37824 ( \38201 , \37807 );
or \U$37825 ( \38202 , \38200 , \38201 );
or \U$37826 ( \38203 , \37807 , \37804 );
nand \U$37827 ( \38204 , \38202 , \38203 );
not \U$37828 ( \38205 , \38204 );
and \U$37829 ( \38206 , \38199 , \38205 );
and \U$37830 ( \38207 , \38106 , \38204 );
nor \U$37831 ( \38208 , \38206 , \38207 );
not \U$37832 ( \38209 , \38208 );
xor \U$37833 ( \38210 , \37795 , \37787 );
xor \U$37834 ( \38211 , \38210 , \37802 );
not \U$37835 ( \38212 , \38211 );
xor \U$37836 ( \38213 , \37199 , \37222 );
xor \U$37837 ( \38214 , \38213 , \37270 );
not \U$37838 ( \38215 , \37920 );
not \U$37839 ( \38216 , \38215 );
not \U$37840 ( \38217 , \37980 );
or \U$37841 ( \38218 , \38216 , \38217 );
or \U$37842 ( \38219 , \37980 , \38215 );
nand \U$37843 ( \38220 , \38218 , \38219 );
not \U$37844 ( \38221 , \38220 );
xor \U$37845 ( \38222 , \37557 , \37519 );
xor \U$37846 ( \38223 , \38222 , \37530 );
not \U$37847 ( \38224 , \38223 );
or \U$37848 ( \38225 , \38221 , \38224 );
or \U$37849 ( \38226 , \38223 , \38220 );
nand \U$37850 ( \38227 , \38225 , \38226 );
xor \U$37851 ( \38228 , \37940 , \37945 );
xor \U$37852 ( \38229 , \38228 , \37956 );
not \U$37853 ( \38230 , \6212 );
not \U$37854 ( \38231 , \38038 );
or \U$37855 ( \38232 , \38230 , \38231 );
and \U$37856 ( \38233 , \16194 , RIae79ef8_167);
not \U$37857 ( \38234 , \16194 );
and \U$37858 ( \38235 , \38234 , \9560 );
nor \U$37859 ( \38236 , \38233 , \38235 );
nand \U$37860 ( \38237 , \38236 , \6200 );
nand \U$37861 ( \38238 , \38232 , \38237 );
xor \U$37862 ( \38239 , \38229 , \38238 );
not \U$37863 ( \38240 , \37970 );
not \U$37864 ( \38241 , \9814 );
or \U$37865 ( \38242 , \38240 , \38241 );
and \U$37866 ( \38243 , RIae7a2b8_175, \10071 );
not \U$37867 ( \38244 , RIae7a2b8_175);
and \U$37868 ( \38245 , \38244 , \10072 );
nor \U$37869 ( \38246 , \38243 , \38245 );
not \U$37870 ( \38247 , \9792 );
or \U$37871 ( \38248 , \38246 , \38247 );
nand \U$37872 ( \38249 , \38242 , \38248 );
and \U$37873 ( \38250 , \38239 , \38249 );
and \U$37874 ( \38251 , \38229 , \38238 );
or \U$37875 ( \38252 , \38250 , \38251 );
not \U$37876 ( \38253 , \38252 );
xnor \U$37877 ( \38254 , \37972 , \37963 );
not \U$37878 ( \38255 , \38254 );
or \U$37879 ( \38256 , \38253 , \38255 );
or \U$37880 ( \38257 , \38252 , \38254 );
nand \U$37881 ( \38258 , \38256 , \38257 );
not \U$37882 ( \38259 , \38258 );
not \U$37883 ( \38260 , \10667 );
and \U$37884 ( \38261 , \24815 , RIae7a150_172);
not \U$37885 ( \38262 , \24815 );
and \U$37886 ( \38263 , \38262 , \10672 );
nor \U$37887 ( \38264 , \38261 , \38263 );
not \U$37888 ( \38265 , \38264 );
or \U$37889 ( \38266 , \38260 , \38265 );
nand \U$37890 ( \38267 , \37885 , \9777 );
nand \U$37891 ( \38268 , \38266 , \38267 );
not \U$37892 ( \38269 , \38268 );
not \U$37893 ( \38270 , \37827 );
not \U$37894 ( \38271 , \37843 );
or \U$37895 ( \38272 , \38270 , \38271 );
or \U$37896 ( \38273 , \37843 , \37827 );
nand \U$37897 ( \38274 , \38272 , \38273 );
not \U$37898 ( \38275 , \2417 );
not \U$37899 ( \38276 , RIae79c28_161);
not \U$37900 ( \38277 , \10844 );
or \U$37901 ( \38278 , \38276 , \38277 );
or \U$37902 ( \38279 , \17166 , RIae79c28_161);
nand \U$37903 ( \38280 , \38278 , \38279 );
not \U$37904 ( \38281 , \38280 );
or \U$37905 ( \38282 , \38275 , \38281 );
nand \U$37906 ( \38283 , \37954 , \2418 );
nand \U$37907 ( \38284 , \38282 , \38283 );
xor \U$37908 ( \38285 , \38274 , \38284 );
not \U$37909 ( \38286 , \38285 );
not \U$37910 ( \38287 , \5048 );
not \U$37911 ( \38288 , \37814 );
or \U$37912 ( \38289 , \38287 , \38288 );
and \U$37913 ( \38290 , \10042 , \4968 );
not \U$37914 ( \38291 , \10042 );
and \U$37915 ( \38292 , \38291 , RIae79d90_164);
or \U$37916 ( \38293 , \38290 , \38292 );
nand \U$37917 ( \38294 , \38293 , \5039 );
nand \U$37918 ( \38295 , \38289 , \38294 );
not \U$37919 ( \38296 , \38295 );
or \U$37920 ( \38297 , \38286 , \38296 );
nand \U$37921 ( \38298 , \38284 , \38274 );
nand \U$37922 ( \38299 , \38297 , \38298 );
not \U$37923 ( \38300 , \10519 );
not \U$37924 ( \38301 , \38077 );
or \U$37925 ( \38302 , \38300 , \38301 );
not \U$37926 ( \38303 , \9529 );
not \U$37927 ( \38304 , \5722 );
or \U$37928 ( \38305 , \38303 , \38304 );
or \U$37929 ( \38306 , \9280 , \9529 );
nand \U$37930 ( \38307 , \38305 , \38306 );
nand \U$37931 ( \38308 , \38307 , \9549 );
nand \U$37932 ( \38309 , \38302 , \38308 );
xor \U$37933 ( \38310 , \38299 , \38309 );
not \U$37934 ( \38311 , \38310 );
or \U$37935 ( \38312 , \38269 , \38311 );
nand \U$37936 ( \38313 , \38309 , \38299 );
nand \U$37937 ( \38314 , \38312 , \38313 );
not \U$37938 ( \38315 , \38314 );
or \U$37939 ( \38316 , \38259 , \38315 );
not \U$37940 ( \38317 , \38254 );
nand \U$37941 ( \38318 , \38317 , \38252 );
nand \U$37942 ( \38319 , \38316 , \38318 );
nand \U$37943 ( \38320 , \38227 , \38319 );
not \U$37944 ( \38321 , \38223 );
nand \U$37945 ( \38322 , \38321 , \38220 );
nand \U$37946 ( \38323 , \38214 , \38320 , \38322 );
not \U$37947 ( \38324 , \38322 );
not \U$37948 ( \38325 , \38320 );
or \U$37949 ( \38326 , \38324 , \38325 );
not \U$37950 ( \38327 , \38214 );
nand \U$37951 ( \38328 , \38326 , \38327 );
nand \U$37952 ( \38329 , \38323 , \38328 );
not \U$37953 ( \38330 , \38329 );
or \U$37954 ( \38331 , \38212 , \38330 );
not \U$37955 ( \38332 , \38322 );
not \U$37956 ( \38333 , \38320 );
or \U$37957 ( \38334 , \38332 , \38333 );
nand \U$37958 ( \38335 , \38334 , \38214 );
nand \U$37959 ( \38336 , \38331 , \38335 );
not \U$37960 ( \38337 , \38336 );
nand \U$37961 ( \38338 , \38209 , \38337 );
not \U$37962 ( \38339 , \38338 );
not \U$37963 ( \38340 , \37910 );
xor \U$37964 ( \38341 , \37985 , \38340 );
xnor \U$37965 ( \38342 , \38341 , \38104 );
not \U$37966 ( \38343 , \38342 );
xor \U$37967 ( \38344 , \37890 , \37905 );
not \U$37968 ( \38345 , \38344 );
xor \U$37969 ( \38346 , \38069 , \38056 );
xnor \U$37970 ( \38347 , \38346 , \38079 );
not \U$37971 ( \38348 , \38347 );
xor \U$37972 ( \38349 , \37863 , \37887 );
xor \U$37973 ( \38350 , \38349 , \37876 );
not \U$37974 ( \38351 , \38350 );
not \U$37975 ( \38352 , \38351 );
or \U$37976 ( \38353 , \38348 , \38352 );
not \U$37977 ( \38354 , \38002 );
not \U$37978 ( \38355 , \38013 );
not \U$37979 ( \38356 , \38355 );
or \U$37980 ( \38357 , \38354 , \38356 );
or \U$37981 ( \38358 , \38355 , \38002 );
nand \U$37982 ( \38359 , \38357 , \38358 );
not \U$37983 ( \38360 , \38347 );
nand \U$37984 ( \38361 , \38350 , \38360 );
nand \U$37985 ( \38362 , \38359 , \38361 );
nand \U$37986 ( \38363 , \38353 , \38362 );
not \U$37987 ( \38364 , \38363 );
not \U$37988 ( \38365 , \11014 );
not \U$37989 ( \38366 , \11690 );
not \U$37990 ( \38367 , \12484 );
or \U$37991 ( \38368 , \38366 , \38367 );
or \U$37992 ( \38369 , \9609 , \11690 );
nand \U$37993 ( \38370 , \38368 , \38369 );
not \U$37994 ( \38371 , \38370 );
or \U$37995 ( \38372 , \38365 , \38371 );
nand \U$37996 ( \38373 , \38054 , \9622 );
nand \U$37997 ( \38374 , \38372 , \38373 );
not \U$37998 ( \38375 , \11098 );
not \U$37999 ( \38376 , \37871 );
or \U$38000 ( \38377 , \38375 , \38376 );
and \U$38001 ( \38378 , RIae7a060_170, \9298 );
not \U$38002 ( \38379 , RIae7a060_170);
and \U$38003 ( \38380 , \38379 , \9299 );
nor \U$38004 ( \38381 , \38378 , \38380 );
nand \U$38005 ( \38382 , \38381 , \17797 );
nand \U$38006 ( \38383 , \38377 , \38382 );
xor \U$38007 ( \38384 , \38374 , \38383 );
not \U$38008 ( \38385 , \14510 );
and \U$38009 ( \38386 , RIae7a8d0_188, \19325 );
not \U$38010 ( \38387 , RIae7a8d0_188);
and \U$38011 ( \38388 , \38387 , \24742 );
or \U$38012 ( \38389 , \38386 , \38388 );
not \U$38013 ( \38390 , \38389 );
or \U$38014 ( \38391 , \38385 , \38390 );
nand \U$38015 ( \38392 , \38129 , \10275 );
nand \U$38016 ( \38393 , \38391 , \38392 );
and \U$38017 ( \38394 , \38384 , \38393 );
and \U$38018 ( \38395 , \38374 , \38383 );
or \U$38019 ( \38396 , \38394 , \38395 );
not \U$38020 ( \38397 , \38396 );
not \U$38021 ( \38398 , \38041 );
not \U$38022 ( \38399 , \38022 );
and \U$38023 ( \38400 , \38398 , \38399 );
and \U$38024 ( \38401 , \38041 , \38022 );
nor \U$38025 ( \38402 , \38400 , \38401 );
not \U$38026 ( \38403 , \38402 );
not \U$38027 ( \38404 , \10709 );
not \U$38028 ( \38405 , RIae79fe8_169);
not \U$38029 ( \38406 , \10750 );
or \U$38030 ( \38407 , \38405 , \38406 );
or \U$38031 ( \38408 , \9875 , RIae79fe8_169);
nand \U$38032 ( \38409 , \38407 , \38408 );
not \U$38033 ( \38410 , \38409 );
or \U$38034 ( \38411 , \38404 , \38410 );
nand \U$38035 ( \38412 , \38032 , \9517 );
nand \U$38036 ( \38413 , \38411 , \38412 );
not \U$38037 ( \38414 , \19466 );
not \U$38038 ( \38415 , \11114 );
not \U$38039 ( \38416 , \10725 );
not \U$38040 ( \38417 , \38416 );
or \U$38041 ( \38418 , \38415 , \38417 );
nand \U$38042 ( \38419 , \13657 , RIae7a240_174);
nand \U$38043 ( \38420 , \38418 , \38419 );
not \U$38044 ( \38421 , \38420 );
or \U$38045 ( \38422 , \38414 , \38421 );
nand \U$38046 ( \38423 , \38066 , \9699 );
nand \U$38047 ( \38424 , \38422 , \38423 );
xor \U$38048 ( \38425 , \38413 , \38424 );
not \U$38049 ( \38426 , \10927 );
not \U$38050 ( \38427 , \17324 );
not \U$38051 ( \38428 , \10938 );
or \U$38052 ( \38429 , \38427 , \38428 );
nand \U$38053 ( \38430 , \19422 , RIae7a510_180);
nand \U$38054 ( \38431 , \38429 , \38430 );
not \U$38055 ( \38432 , \38431 );
or \U$38056 ( \38433 , \38426 , \38432 );
nand \U$38057 ( \38434 , \37996 , \16358 );
nand \U$38058 ( \38435 , \38433 , \38434 );
and \U$38059 ( \38436 , \38425 , \38435 );
and \U$38060 ( \38437 , \38413 , \38424 );
or \U$38061 ( \38438 , \38436 , \38437 );
not \U$38062 ( \38439 , \38438 );
or \U$38063 ( \38440 , \38403 , \38439 );
or \U$38064 ( \38441 , \38438 , \38402 );
nand \U$38065 ( \38442 , \38440 , \38441 );
not \U$38066 ( \38443 , \38442 );
or \U$38067 ( \38444 , \38397 , \38443 );
not \U$38068 ( \38445 , \38402 );
nand \U$38069 ( \38446 , \38445 , \38438 );
nand \U$38070 ( \38447 , \38444 , \38446 );
not \U$38071 ( \38448 , \38447 );
not \U$38072 ( \38449 , \38448 );
or \U$38073 ( \38450 , \38364 , \38449 );
or \U$38074 ( \38451 , \38363 , \38448 );
nand \U$38075 ( \38452 , \38450 , \38451 );
not \U$38076 ( \38453 , \38452 );
or \U$38077 ( \38454 , \38345 , \38453 );
not \U$38078 ( \38455 , \38448 );
nand \U$38079 ( \38456 , \38455 , \38363 );
nand \U$38080 ( \38457 , \38454 , \38456 );
not \U$38081 ( \38458 , \38457 );
nand \U$38082 ( \38459 , \38343 , \38458 );
not \U$38083 ( \38460 , \38459 );
not \U$38084 ( \38461 , \38152 );
not \U$38085 ( \38462 , \38461 );
not \U$38086 ( \38463 , \38143 );
or \U$38087 ( \38464 , \38462 , \38463 );
or \U$38088 ( \38465 , \38461 , \38143 );
nand \U$38089 ( \38466 , \38464 , \38465 );
not \U$38090 ( \38467 , \38466 );
not \U$38091 ( \38468 , \14668 );
and \U$38092 ( \38469 , \1860 , \14671 );
not \U$38093 ( \38470 , \1860 );
and \U$38094 ( \38471 , \38470 , RIae7aa38_191);
nor \U$38095 ( \38472 , \38469 , \38471 );
not \U$38096 ( \38473 , \38472 );
or \U$38097 ( \38474 , \38468 , \38473 );
nand \U$38098 ( \38475 , \38150 , RIae7aab0_192);
nand \U$38099 ( \38476 , \38474 , \38475 );
not \U$38100 ( \38477 , \38476 );
not \U$38101 ( \38478 , \9473 );
xor \U$38102 ( \38479 , \4972 , RIae7a6f0_184);
not \U$38103 ( \38480 , \38479 );
or \U$38104 ( \38481 , \38478 , \38480 );
nand \U$38105 ( \38482 , \38011 , \9478 );
nand \U$38106 ( \38483 , \38481 , \38482 );
not \U$38107 ( \38484 , \38483 );
not \U$38108 ( \38485 , \10696 );
not \U$38109 ( \38486 , \10625 );
not \U$38110 ( \38487 , \9438 );
or \U$38111 ( \38488 , \38486 , \38487 );
not \U$38112 ( \38489 , \14110 );
nand \U$38113 ( \38490 , \38489 , RIae7a498_179);
nand \U$38114 ( \38491 , \38488 , \38490 );
not \U$38115 ( \38492 , \38491 );
or \U$38116 ( \38493 , \38485 , \38492 );
nand \U$38117 ( \38494 , \38136 , \10677 );
nand \U$38118 ( \38495 , \38493 , \38494 );
not \U$38119 ( \38496 , \38495 );
nand \U$38120 ( \38497 , \38484 , \38496 );
not \U$38121 ( \38498 , \38497 );
or \U$38122 ( \38499 , \38477 , \38498 );
nand \U$38123 ( \38500 , \38483 , \38495 );
nand \U$38124 ( \38501 , \38499 , \38500 );
not \U$38125 ( \38502 , \38501 );
xnor \U$38126 ( \38503 , \37858 , \37823 );
not \U$38127 ( \38504 , \38503 );
not \U$38128 ( \38505 , RIae7a2b8_175);
not \U$38129 ( \38506 , \10171 );
or \U$38130 ( \38507 , \38505 , \38506 );
or \U$38131 ( \38508 , \10171 , RIae7a2b8_175);
nand \U$38132 ( \38509 , \38507 , \38508 );
not \U$38133 ( \38510 , \38509 );
not \U$38134 ( \38511 , \9792 );
or \U$38135 ( \38512 , \38510 , \38511 );
not \U$38136 ( \38513 , \38246 );
nand \U$38137 ( \38514 , \38513 , \9814 );
nand \U$38138 ( \38515 , \38512 , \38514 );
not \U$38139 ( \38516 , \38515 );
not \U$38140 ( \38517 , \37852 );
or \U$38141 ( \38518 , \38517 , \4852 );
not \U$38142 ( \38519 , \2406 );
not \U$38143 ( \38520 , \10272 );
or \U$38144 ( \38521 , \38519 , \38520 );
or \U$38145 ( \38522 , \12842 , \26312 );
nand \U$38146 ( \38523 , \38521 , \38522 );
not \U$38147 ( \38524 , \38523 );
or \U$38148 ( \38525 , \38524 , \11760 );
nand \U$38149 ( \38526 , \38518 , \38525 );
and \U$38150 ( \38527 , \12857 , \2450 );
not \U$38151 ( \38528 , \2418 );
not \U$38152 ( \38529 , \38280 );
or \U$38153 ( \38530 , \38528 , \38529 );
not \U$38154 ( \38531 , \12750 );
not \U$38155 ( \38532 , RIae79c28_161);
and \U$38156 ( \38533 , \38531 , \38532 );
and \U$38157 ( \38534 , \16006 , RIae79c28_161);
nor \U$38158 ( \38535 , \38533 , \38534 );
not \U$38159 ( \38536 , \38535 );
nand \U$38160 ( \38537 , \38536 , \2417 );
nand \U$38161 ( \38538 , \38530 , \38537 );
xor \U$38162 ( \38539 , \38527 , \38538 );
not \U$38163 ( \38540 , \4155 );
not \U$38164 ( \38541 , \38523 );
or \U$38165 ( \38542 , \38540 , \38541 );
not \U$38166 ( \38543 , \11755 );
not \U$38167 ( \38544 , \18971 );
or \U$38168 ( \38545 , \38543 , \38544 );
nand \U$38169 ( \38546 , \10259 , RIae79ca0_162);
nand \U$38170 ( \38547 , \38545 , \38546 );
nand \U$38171 ( \38548 , \38547 , \4154 );
nand \U$38172 ( \38549 , \38542 , \38548 );
and \U$38173 ( \38550 , \38539 , \38549 );
and \U$38174 ( \38551 , \38527 , \38538 );
nor \U$38175 ( \38552 , \38550 , \38551 );
not \U$38176 ( \38553 , \38552 );
xor \U$38177 ( \38554 , \38526 , \38553 );
not \U$38178 ( \38555 , \38554 );
or \U$38179 ( \38556 , \38516 , \38555 );
not \U$38180 ( \38557 , \38552 );
nand \U$38181 ( \38558 , \38557 , \38526 );
nand \U$38182 ( \38559 , \38556 , \38558 );
not \U$38183 ( \38560 , \38559 );
not \U$38184 ( \38561 , \38560 );
or \U$38185 ( \38562 , \38504 , \38561 );
not \U$38186 ( \38563 , \38420 );
not \U$38187 ( \38564 , \9699 );
or \U$38188 ( \38565 , \38563 , \38564 );
not \U$38189 ( \38566 , \11114 );
not \U$38190 ( \38567 , \11386 );
or \U$38191 ( \38568 , \38566 , \38567 );
or \U$38192 ( \38569 , \10087 , \12312 );
nand \U$38193 ( \38570 , \38568 , \38569 );
nand \U$38194 ( \38571 , \38570 , \13720 );
nand \U$38195 ( \38572 , \38565 , \38571 );
not \U$38196 ( \38573 , \38572 );
not \U$38197 ( \38574 , \38236 );
or \U$38198 ( \38575 , \38574 , \6213 );
not \U$38199 ( \38576 , \10149 );
not \U$38200 ( \38577 , RIae79ef8_167);
and \U$38201 ( \38578 , \38576 , \38577 );
and \U$38202 ( \38579 , \10149 , RIae79ef8_167);
nor \U$38203 ( \38580 , \38578 , \38579 );
or \U$38204 ( \38581 , \38580 , \19868 );
nand \U$38205 ( \38582 , \38575 , \38581 );
not \U$38206 ( \38583 , \38582 );
not \U$38207 ( \38584 , \9518 );
not \U$38208 ( \38585 , \38409 );
or \U$38209 ( \38586 , \38584 , \38585 );
and \U$38210 ( \38587 , \16719 , \11069 );
not \U$38211 ( \38588 , \16719 );
and \U$38212 ( \38589 , \38588 , RIae79fe8_169);
nor \U$38213 ( \38590 , \38587 , \38589 );
nand \U$38214 ( \38591 , \38590 , \10709 );
nand \U$38215 ( \38592 , \38586 , \38591 );
not \U$38216 ( \38593 , \38592 );
nand \U$38217 ( \38594 , \38583 , \38593 );
not \U$38218 ( \38595 , \38594 );
or \U$38219 ( \38596 , \38573 , \38595 );
nand \U$38220 ( \38597 , \38592 , \38582 );
nand \U$38221 ( \38598 , \38596 , \38597 );
nand \U$38222 ( \38599 , \38562 , \38598 );
not \U$38223 ( \38600 , \38503 );
nand \U$38224 ( \38601 , \38600 , \38559 );
and \U$38225 ( \38602 , \38599 , \38601 );
nand \U$38226 ( \38603 , \38502 , \38602 );
not \U$38227 ( \38604 , \38603 );
or \U$38228 ( \38605 , \38467 , \38604 );
not \U$38229 ( \38606 , \38602 );
nand \U$38230 ( \38607 , \38606 , \38501 );
nand \U$38231 ( \38608 , \38605 , \38607 );
not \U$38232 ( \38609 , \38608 );
and \U$38233 ( \38610 , \38090 , \38018 );
not \U$38234 ( \38611 , \38090 );
not \U$38235 ( \38612 , \38018 );
and \U$38236 ( \38613 , \38611 , \38612 );
nor \U$38237 ( \38614 , \38610 , \38613 );
xor \U$38238 ( \38615 , \38155 , \38614 );
xnor \U$38239 ( \38616 , \38615 , \38170 );
not \U$38240 ( \38617 , \38616 );
or \U$38241 ( \38618 , \38609 , \38617 );
nand \U$38242 ( \38619 , \38155 , \38170 );
not \U$38243 ( \38620 , \38619 );
not \U$38244 ( \38621 , \38170 );
nand \U$38245 ( \38622 , \38621 , \38156 );
not \U$38246 ( \38623 , \38622 );
or \U$38247 ( \38624 , \38620 , \38623 );
nand \U$38248 ( \38625 , \38624 , \38614 );
nand \U$38249 ( \38626 , \38618 , \38625 );
not \U$38250 ( \38627 , \38626 );
or \U$38251 ( \38628 , \38460 , \38627 );
not \U$38252 ( \38629 , \38343 );
nand \U$38253 ( \38630 , \38629 , \38457 );
nand \U$38254 ( \38631 , \38628 , \38630 );
not \U$38255 ( \38632 , \38631 );
or \U$38256 ( \38633 , \38339 , \38632 );
nand \U$38257 ( \38634 , \38208 , \38336 );
nand \U$38258 ( \38635 , \38633 , \38634 );
xor \U$38259 ( \38636 , \38198 , \38635 );
not \U$38260 ( \38637 , \38186 );
not \U$38261 ( \38638 , \38116 );
or \U$38262 ( \38639 , \38637 , \38638 );
or \U$38263 ( \38640 , \38116 , \38186 );
nand \U$38264 ( \38641 , \38639 , \38640 );
and \U$38265 ( \38642 , \38636 , \38641 );
and \U$38266 ( \38643 , \38198 , \38635 );
or \U$38267 ( \38644 , \38642 , \38643 );
not \U$38268 ( \38645 , \38644 );
nand \U$38269 ( \38646 , \38196 , \38645 );
nand \U$38270 ( \38647 , \37753 , \37763 , \38194 , \38646 );
not \U$38271 ( \38648 , \38647 );
not \U$38272 ( \38649 , \38648 );
not \U$38273 ( \38650 , RIae7aab0_192);
not \U$38274 ( \38651 , \38472 );
or \U$38275 ( \38652 , \38650 , \38651 );
and \U$38276 ( \38653 , \2403 , \11326 );
not \U$38277 ( \38654 , \2403 );
and \U$38278 ( \38655 , \38654 , RIae7aa38_191);
nor \U$38279 ( \38656 , \38653 , \38655 );
nand \U$38280 ( \38657 , \38656 , \14669 );
nand \U$38281 ( \38658 , \38652 , \38657 );
not \U$38282 ( \38659 , \38658 );
not \U$38283 ( \38660 , \9792 );
not \U$38284 ( \38661 , \11054 );
not \U$38285 ( \38662 , \9868 );
or \U$38286 ( \38663 , \38661 , \38662 );
or \U$38287 ( \38664 , \9868 , \9804 );
nand \U$38288 ( \38665 , \38663 , \38664 );
not \U$38289 ( \38666 , \38665 );
or \U$38290 ( \38667 , \38660 , \38666 );
nand \U$38291 ( \38668 , \38509 , \9814 );
nand \U$38292 ( \38669 , \38667 , \38668 );
not \U$38293 ( \38670 , \38669 );
xnor \U$38294 ( \38671 , \38549 , \38539 );
not \U$38295 ( \38672 , \38671 );
not \U$38296 ( \38673 , \9687 );
not \U$38297 ( \38674 , \11114 );
not \U$38298 ( \38675 , \10070 );
or \U$38299 ( \38676 , \38674 , \38675 );
or \U$38300 ( \38677 , \10066 , \11114 );
nand \U$38301 ( \38678 , \38676 , \38677 );
not \U$38302 ( \38679 , \38678 );
or \U$38303 ( \38680 , \38673 , \38679 );
not \U$38304 ( \38681 , \30532 );
nand \U$38305 ( \38682 , \38681 , \38570 );
nand \U$38306 ( \38683 , \38680 , \38682 );
not \U$38307 ( \38684 , \38683 );
or \U$38308 ( \38685 , \38672 , \38684 );
or \U$38309 ( \38686 , \38683 , \38671 );
nand \U$38310 ( \38687 , \38685 , \38686 );
not \U$38311 ( \38688 , \38687 );
or \U$38312 ( \38689 , \38670 , \38688 );
not \U$38313 ( \38690 , \38671 );
nand \U$38314 ( \38691 , \38690 , \38683 );
nand \U$38315 ( \38692 , \38689 , \38691 );
not \U$38316 ( \38693 , \10676 );
not \U$38317 ( \38694 , \38491 );
or \U$38318 ( \38695 , \38693 , \38694 );
and \U$38319 ( \38696 , RIae7a498_179, \14657 );
not \U$38320 ( \38697 , RIae7a498_179);
and \U$38321 ( \38698 , \38697 , \16786 );
or \U$38322 ( \38699 , \38696 , \38698 );
nand \U$38323 ( \38700 , \38699 , \10696 );
nand \U$38324 ( \38701 , \38695 , \38700 );
xor \U$38325 ( \38702 , \38692 , \38701 );
not \U$38326 ( \38703 , \38702 );
or \U$38327 ( \38704 , \38659 , \38703 );
nand \U$38328 ( \38705 , \38692 , \38701 );
nand \U$38329 ( \38706 , \38704 , \38705 );
and \U$38330 ( \38707 , \38310 , \38268 );
not \U$38331 ( \38708 , \38310 );
not \U$38332 ( \38709 , \38268 );
and \U$38333 ( \38710 , \38708 , \38709 );
nor \U$38334 ( \38711 , \38707 , \38710 );
xor \U$38335 ( \38712 , \38706 , \38711 );
not \U$38336 ( \38713 , \38712 );
xor \U$38337 ( \38714 , \38496 , \38476 );
xnor \U$38338 ( \38715 , \38714 , \38483 );
not \U$38339 ( \38716 , \38715 );
not \U$38340 ( \38717 , \38716 );
and \U$38341 ( \38718 , \38713 , \38717 );
and \U$38342 ( \38719 , \38712 , \38716 );
nor \U$38343 ( \38720 , \38718 , \38719 );
not \U$38344 ( \38721 , \38720 );
xor \U$38345 ( \38722 , \38658 , \38702 );
not \U$38346 ( \38723 , \5048 );
xor \U$38347 ( \38724 , RIae79d90_164, \10193 );
not \U$38348 ( \38725 , \38724 );
or \U$38349 ( \38726 , \38723 , \38725 );
not \U$38350 ( \38727 , \4968 );
not \U$38351 ( \38728 , \10272 );
or \U$38352 ( \38729 , \38727 , \38728 );
or \U$38353 ( \38730 , \11318 , \4968 );
nand \U$38354 ( \38731 , \38729 , \38730 );
nand \U$38355 ( \38732 , \38731 , \5039 );
nand \U$38356 ( \38733 , \38726 , \38732 );
not \U$38357 ( \38734 , \5048 );
not \U$38358 ( \38735 , \38731 );
or \U$38359 ( \38736 , \38734 , \38735 );
and \U$38360 ( \38737 , \10259 , \13059 );
not \U$38361 ( \38738 , \10259 );
and \U$38362 ( \38739 , \38738 , RIae79d90_164);
nor \U$38363 ( \38740 , \38737 , \38739 );
nand \U$38364 ( \38741 , \38740 , \5039 );
nand \U$38365 ( \38742 , \38736 , \38741 );
not \U$38366 ( \38743 , \38742 );
nand \U$38367 ( \38744 , \12857 , \2411 );
not \U$38368 ( \38745 , \38744 );
not \U$38369 ( \38746 , \4155 );
not \U$38370 ( \38747 , \2406 );
not \U$38371 ( \38748 , \10845 );
or \U$38372 ( \38749 , \38747 , \38748 );
nand \U$38373 ( \38750 , \16651 , RIae79ca0_162);
nand \U$38374 ( \38751 , \38749 , \38750 );
not \U$38375 ( \38752 , \38751 );
or \U$38376 ( \38753 , \38746 , \38752 );
and \U$38377 ( \38754 , RIae79ca0_162, \12750 );
not \U$38378 ( \38755 , RIae79ca0_162);
and \U$38379 ( \38756 , \38755 , \12751 );
or \U$38380 ( \38757 , \38754 , \38756 );
nand \U$38381 ( \38758 , \38757 , \4154 );
nand \U$38382 ( \38759 , \38753 , \38758 );
not \U$38383 ( \38760 , \38759 );
or \U$38384 ( \38761 , \38745 , \38760 );
or \U$38385 ( \38762 , \38759 , \38744 );
nand \U$38386 ( \38763 , \38761 , \38762 );
not \U$38387 ( \38764 , \38763 );
or \U$38388 ( \38765 , \38743 , \38764 );
not \U$38389 ( \38766 , \38744 );
nand \U$38390 ( \38767 , \38766 , \38759 );
nand \U$38391 ( \38768 , \38765 , \38767 );
xor \U$38392 ( \38769 , \38733 , \38768 );
not \U$38393 ( \38770 , \9699 );
not \U$38394 ( \38771 , \38678 );
or \U$38395 ( \38772 , \38770 , \38771 );
and \U$38396 ( \38773 , RIae7a240_174, \11272 );
not \U$38397 ( \38774 , RIae7a240_174);
and \U$38398 ( \38775 , \38774 , \9897 );
nor \U$38399 ( \38776 , \38773 , \38775 );
nand \U$38400 ( \38777 , \38776 , \19466 );
nand \U$38401 ( \38778 , \38772 , \38777 );
and \U$38402 ( \38779 , \38769 , \38778 );
and \U$38403 ( \38780 , \38733 , \38768 );
nor \U$38404 ( \38781 , \38779 , \38780 );
not \U$38405 ( \38782 , \38781 );
not \U$38406 ( \38783 , \9504 );
not \U$38407 ( \38784 , \27671 );
or \U$38408 ( \38785 , \38783 , \38784 );
or \U$38409 ( \38786 , \27671 , \11069 );
nand \U$38410 ( \38787 , \38785 , \38786 );
and \U$38411 ( \38788 , \38787 , \9517 );
and \U$38412 ( \38789 , RIae79fe8_169, \10149 );
not \U$38413 ( \38790 , RIae79fe8_169);
and \U$38414 ( \38791 , \38790 , \10141 );
or \U$38415 ( \38792 , \38789 , \38791 );
and \U$38416 ( \38793 , \38792 , \9499 );
nor \U$38417 ( \38794 , \38788 , \38793 );
not \U$38418 ( \38795 , \38794 );
not \U$38419 ( \38796 , \16135 );
not \U$38420 ( \38797 , \38665 );
or \U$38421 ( \38798 , \38796 , \38797 );
xor \U$38422 ( \38799 , \10007 , RIae7a2b8_175);
nand \U$38423 ( \38800 , \38799 , \9792 );
nand \U$38424 ( \38801 , \38798 , \38800 );
not \U$38425 ( \38802 , \38801 );
or \U$38426 ( \38803 , \38795 , \38802 );
or \U$38427 ( \38804 , \38801 , \38794 );
nand \U$38428 ( \38805 , \38803 , \38804 );
not \U$38429 ( \38806 , \38805 );
not \U$38430 ( \38807 , \9621 );
not \U$38431 ( \38808 , RIae7a3a8_177);
not \U$38432 ( \38809 , \17400 );
or \U$38433 ( \38810 , \38808 , \38809 );
or \U$38434 ( \38811 , \10729 , RIae7a3a8_177);
nand \U$38435 ( \38812 , \38810 , \38811 );
not \U$38436 ( \38813 , \38812 );
or \U$38437 ( \38814 , \38807 , \38813 );
not \U$38438 ( \38815 , \16469 );
not \U$38439 ( \38816 , \15653 );
not \U$38440 ( \38817 , \38816 );
or \U$38441 ( \38818 , \38815 , \38817 );
nand \U$38442 ( \38819 , \17406 , RIae7a3a8_177);
nand \U$38443 ( \38820 , \38818 , \38819 );
nand \U$38444 ( \38821 , \38820 , \11013 );
nand \U$38445 ( \38822 , \38814 , \38821 );
not \U$38446 ( \38823 , \38822 );
or \U$38447 ( \38824 , \38806 , \38823 );
not \U$38448 ( \38825 , \38794 );
nand \U$38449 ( \38826 , \38825 , \38801 );
nand \U$38450 ( \38827 , \38824 , \38826 );
not \U$38451 ( \38828 , \38827 );
or \U$38452 ( \38829 , \38782 , \38828 );
or \U$38453 ( \38830 , \38827 , \38781 );
nand \U$38454 ( \38831 , \38829 , \38830 );
not \U$38455 ( \38832 , \38831 );
not \U$38456 ( \38833 , \10631 );
not \U$38457 ( \38834 , \9412 );
not \U$38458 ( \38835 , RIae7a510_180);
and \U$38459 ( \38836 , \38834 , \38835 );
and \U$38460 ( \38837 , \11804 , RIae7a510_180);
nor \U$38461 ( \38838 , \38836 , \38837 );
not \U$38462 ( \38839 , \38838 );
not \U$38463 ( \38840 , \38839 );
or \U$38464 ( \38841 , \38833 , \38840 );
xor \U$38465 ( \38842 , RIae7a510_180, \12482 );
nand \U$38466 ( \38843 , \38842 , \10637 );
nand \U$38467 ( \38844 , \38841 , \38843 );
not \U$38468 ( \38845 , \38844 );
not \U$38469 ( \38846 , \9643 );
not \U$38470 ( \38847 , \38812 );
or \U$38471 ( \38848 , \38846 , \38847 );
not \U$38472 ( \38849 , RIae7a3a8_177);
not \U$38473 ( \38850 , \11187 );
or \U$38474 ( \38851 , \38849 , \38850 );
or \U$38475 ( \38852 , \11187 , RIae7a3a8_177);
nand \U$38476 ( \38853 , \38851 , \38852 );
nand \U$38477 ( \38854 , \38853 , \9622 );
nand \U$38478 ( \38855 , \38848 , \38854 );
not \U$38479 ( \38856 , \38855 );
not \U$38480 ( \38857 , \9517 );
not \U$38481 ( \38858 , \38590 );
or \U$38482 ( \38859 , \38857 , \38858 );
nand \U$38483 ( \38860 , \38787 , \9499 );
nand \U$38484 ( \38861 , \38859 , \38860 );
not \U$38485 ( \38862 , \38861 );
not \U$38486 ( \38863 , \38862 );
and \U$38487 ( \38864 , \38856 , \38863 );
and \U$38488 ( \38865 , \38855 , \38862 );
nor \U$38489 ( \38866 , \38864 , \38865 );
not \U$38490 ( \38867 , \38866 );
or \U$38491 ( \38868 , \38845 , \38867 );
or \U$38492 ( \38869 , \38866 , \38844 );
nand \U$38493 ( \38870 , \38868 , \38869 );
not \U$38494 ( \38871 , \38870 );
or \U$38495 ( \38872 , \38832 , \38871 );
not \U$38496 ( \38873 , \38781 );
nand \U$38497 ( \38874 , \38873 , \38827 );
nand \U$38498 ( \38875 , \38872 , \38874 );
xor \U$38499 ( \38876 , \38722 , \38875 );
not \U$38500 ( \38877 , \38876 );
xor \U$38501 ( \38878 , \38687 , \38669 );
not \U$38502 ( \38879 , \9776 );
not \U$38503 ( \38880 , \10672 );
not \U$38504 ( \38881 , \9438 );
or \U$38505 ( \38882 , \38880 , \38881 );
or \U$38506 ( \38883 , \12614 , \10658 );
nand \U$38507 ( \38884 , \38882 , \38883 );
not \U$38508 ( \38885 , \38884 );
or \U$38509 ( \38886 , \38879 , \38885 );
not \U$38510 ( \38887 , RIae7a150_172);
not \U$38511 ( \38888 , \32526 );
or \U$38512 ( \38889 , \38887 , \38888 );
nand \U$38513 ( \38890 , \9455 , \10658 );
nand \U$38514 ( \38891 , \38889 , \38890 );
nand \U$38515 ( \38892 , \38891 , \9758 );
nand \U$38516 ( \38893 , \38886 , \38892 );
not \U$38517 ( \38894 , \9705 );
and \U$38518 ( \38895 , RIae7a6f0_184, \5722 );
not \U$38519 ( \38896 , RIae7a6f0_184);
and \U$38520 ( \38897 , \38896 , \28338 );
nor \U$38521 ( \38898 , \38895 , \38897 );
not \U$38522 ( \38899 , \38898 );
or \U$38523 ( \38900 , \38894 , \38899 );
and \U$38524 ( \38901 , RIae7a6f0_184, \9286 );
not \U$38525 ( \38902 , RIae7a6f0_184);
and \U$38526 ( \38903 , \38902 , \6345 );
or \U$38527 ( \38904 , \38901 , \38903 );
nand \U$38528 ( \38905 , \38904 , \9473 );
nand \U$38529 ( \38906 , \38900 , \38905 );
xor \U$38530 ( \38907 , \38893 , \38906 );
not \U$38531 ( \38908 , \14668 );
not \U$38532 ( \38909 , RIae7aa38_191);
not \U$38533 ( \38910 , \21873 );
or \U$38534 ( \38911 , \38909 , \38910 );
or \U$38535 ( \38912 , \6244 , RIae7aa38_191);
nand \U$38536 ( \38913 , \38911 , \38912 );
not \U$38537 ( \38914 , \38913 );
or \U$38538 ( \38915 , \38908 , \38914 );
not \U$38539 ( \38916 , RIae7aa38_191);
not \U$38540 ( \38917 , \29061 );
or \U$38541 ( \38918 , \38916 , \38917 );
or \U$38542 ( \38919 , \10809 , RIae7aa38_191);
nand \U$38543 ( \38920 , \38918 , \38919 );
nand \U$38544 ( \38921 , \38920 , RIae7aab0_192);
nand \U$38545 ( \38922 , \38915 , \38921 );
and \U$38546 ( \38923 , \38907 , \38922 );
and \U$38547 ( \38924 , \38893 , \38906 );
or \U$38548 ( \38925 , \38923 , \38924 );
xor \U$38549 ( \38926 , \38878 , \38925 );
not \U$38550 ( \38927 , \9499 );
and \U$38551 ( \38928 , RIae79fe8_169, \11589 );
not \U$38552 ( \38929 , RIae79fe8_169);
and \U$38553 ( \38930 , \38929 , \10856 );
or \U$38554 ( \38931 , \38928 , \38930 );
not \U$38555 ( \38932 , \38931 );
or \U$38556 ( \38933 , \38927 , \38932 );
nand \U$38557 ( \38934 , \38792 , \9517 );
nand \U$38558 ( \38935 , \38933 , \38934 );
not \U$38559 ( \38936 , \38935 );
not \U$38560 ( \38937 , \4155 );
not \U$38561 ( \38938 , \38757 );
or \U$38562 ( \38939 , \38937 , \38938 );
not \U$38563 ( \38940 , \4844 );
not \U$38564 ( \38941 , \12857 );
or \U$38565 ( \38942 , \38940 , \38941 );
or \U$38566 ( \38943 , \12857 , \11755 );
nand \U$38567 ( \38944 , \38942 , \38943 );
nand \U$38568 ( \38945 , \38944 , \4154 );
nand \U$38569 ( \38946 , \38939 , \38945 );
not \U$38570 ( \38947 , \4146 );
nand \U$38571 ( \38948 , \38947 , \12857 );
nand \U$38572 ( \38949 , \38948 , \4144 , RIae79ca0_162);
not \U$38573 ( \38950 , \38949 );
and \U$38574 ( \38951 , \38946 , \38950 );
not \U$38575 ( \38952 , \6212 );
and \U$38576 ( \38953 , RIae79ef8_167, \10042 );
not \U$38577 ( \38954 , RIae79ef8_167);
and \U$38578 ( \38955 , \38954 , \10046 );
nor \U$38579 ( \38956 , \38953 , \38955 );
not \U$38580 ( \38957 , \38956 );
or \U$38581 ( \38958 , \38952 , \38957 );
not \U$38582 ( \38959 , RIae79ef8_167);
not \U$38583 ( \38960 , \16036 );
or \U$38584 ( \38961 , \38959 , \38960 );
or \U$38585 ( \38962 , \11581 , RIae79ef8_167);
nand \U$38586 ( \38963 , \38961 , \38962 );
nand \U$38587 ( \38964 , \38963 , \6199 );
nand \U$38588 ( \38965 , \38958 , \38964 );
xor \U$38589 ( \38966 , \38951 , \38965 );
not \U$38590 ( \38967 , \38966 );
or \U$38591 ( \38968 , \38936 , \38967 );
nand \U$38592 ( \38969 , \38965 , \38951 );
nand \U$38593 ( \38970 , \38968 , \38969 );
not \U$38594 ( \38971 , \10519 );
and \U$38595 ( \38972 , RIae7a7e0_186, \12684 );
not \U$38596 ( \38973 , RIae7a7e0_186);
and \U$38597 ( \38974 , \38973 , \6232 );
or \U$38598 ( \38975 , \38972 , \38974 );
not \U$38599 ( \38976 , \38975 );
or \U$38600 ( \38977 , \38971 , \38976 );
and \U$38601 ( \38978 , \9316 , \9537 );
not \U$38602 ( \38979 , \9316 );
and \U$38603 ( \38980 , \38979 , RIae7a7e0_186);
nor \U$38604 ( \38981 , \38978 , \38980 );
nand \U$38605 ( \38982 , \38981 , \9549 );
nand \U$38606 ( \38983 , \38977 , \38982 );
xor \U$38607 ( \38984 , \38970 , \38983 );
not \U$38608 ( \38985 , \9745 );
not \U$38609 ( \38986 , RIae7a060_170);
not \U$38610 ( \38987 , \17387 );
or \U$38611 ( \38988 , \38986 , \38987 );
or \U$38612 ( \38989 , \15520 , RIae7a060_170);
nand \U$38613 ( \38990 , \38988 , \38989 );
not \U$38614 ( \38991 , \38990 );
or \U$38615 ( \38992 , \38985 , \38991 );
and \U$38616 ( \38993 , \11102 , \15091 );
not \U$38617 ( \38994 , \11102 );
and \U$38618 ( \38995 , \38994 , \29050 );
or \U$38619 ( \38996 , \38993 , \38995 );
nand \U$38620 ( \38997 , \38996 , \9729 );
nand \U$38621 ( \38998 , \38992 , \38997 );
and \U$38622 ( \38999 , \38984 , \38998 );
and \U$38623 ( \39000 , \38970 , \38983 );
or \U$38624 ( \39001 , \38999 , \39000 );
and \U$38625 ( \39002 , \38926 , \39001 );
and \U$38626 ( \39003 , \38878 , \38925 );
or \U$38627 ( \39004 , \39002 , \39003 );
not \U$38628 ( \39005 , \39004 );
or \U$38629 ( \39006 , \38877 , \39005 );
nand \U$38630 ( \39007 , \38875 , \38722 );
nand \U$38631 ( \39008 , \39006 , \39007 );
not \U$38632 ( \39009 , \39008 );
and \U$38633 ( \39010 , \38721 , \39009 );
and \U$38634 ( \39011 , \39008 , \38720 );
nor \U$38635 ( \39012 , \39010 , \39011 );
not \U$38636 ( \39013 , \39012 );
not \U$38637 ( \39014 , \39013 );
xor \U$38638 ( \39015 , \38582 , \38593 );
xor \U$38639 ( \39016 , \39015 , \38572 );
not \U$38640 ( \39017 , \9622 );
not \U$38641 ( \39018 , \38370 );
or \U$38642 ( \39019 , \39017 , \39018 );
nand \U$38643 ( \39020 , \38853 , \9643 );
nand \U$38644 ( \39021 , \39019 , \39020 );
xor \U$38645 ( \39022 , \38295 , \38285 );
xor \U$38646 ( \39023 , \39021 , \39022 );
and \U$38647 ( \39024 , \38431 , \10631 );
not \U$38648 ( \39025 , \10927 );
nor \U$38649 ( \39026 , \39025 , \38838 );
nor \U$38650 ( \39027 , \39024 , \39026 );
xnor \U$38651 ( \39028 , \39023 , \39027 );
xor \U$38652 ( \39029 , \39016 , \39028 );
not \U$38653 ( \39030 , \9776 );
and \U$38654 ( \39031 , RIae7a150_172, \13287 );
not \U$38655 ( \39032 , RIae7a150_172);
and \U$38656 ( \39033 , \39032 , \15091 );
or \U$38657 ( \39034 , \39031 , \39033 );
not \U$38658 ( \39035 , \39034 );
or \U$38659 ( \39036 , \39030 , \39035 );
nand \U$38660 ( \39037 , \38884 , \9758 );
nand \U$38661 ( \39038 , \39036 , \39037 );
not \U$38662 ( \39039 , \9730 );
not \U$38663 ( \39040 , \38990 );
or \U$38664 ( \39041 , \39039 , \39040 );
and \U$38665 ( \39042 , RIae7a060_170, \14644 );
not \U$38666 ( \39043 , RIae7a060_170);
and \U$38667 ( \39044 , \39043 , \9313 );
nor \U$38668 ( \39045 , \39042 , \39044 );
nand \U$38669 ( \39046 , \39045 , \9745 );
nand \U$38670 ( \39047 , \39041 , \39046 );
xor \U$38671 ( \39048 , \39038 , \39047 );
not \U$38672 ( \39049 , \16383 );
not \U$38673 ( \39050 , \38920 );
or \U$38674 ( \39051 , \39049 , \39050 );
nand \U$38675 ( \39052 , \38656 , RIae7aab0_192);
nand \U$38676 ( \39053 , \39051 , \39052 );
and \U$38677 ( \39054 , \39048 , \39053 );
and \U$38678 ( \39055 , \39038 , \39047 );
or \U$38679 ( \39056 , \39054 , \39055 );
xnor \U$38680 ( \39057 , \39029 , \39056 );
buf \U$38681 ( \39058 , \39057 );
not \U$38682 ( \39059 , \39058 );
not \U$38683 ( \39060 , \10519 );
and \U$38684 ( \39061 , RIae7a7e0_186, \14630 );
not \U$38685 ( \39062 , RIae7a7e0_186);
and \U$38686 ( \39063 , \39062 , \9290 );
or \U$38687 ( \39064 , \39061 , \39063 );
not \U$38688 ( \39065 , \39064 );
or \U$38689 ( \39066 , \39060 , \39065 );
nand \U$38690 ( \39067 , \38975 , \11851 );
nand \U$38691 ( \39068 , \39066 , \39067 );
not \U$38692 ( \39069 , \39068 );
not \U$38693 ( \39070 , \4155 );
not \U$38694 ( \39071 , \38547 );
or \U$38695 ( \39072 , \39070 , \39071 );
nand \U$38696 ( \39073 , \38751 , \4154 );
nand \U$38697 ( \39074 , \39072 , \39073 );
not \U$38698 ( \39075 , \39074 );
not \U$38699 ( \39076 , \10584 );
not \U$38700 ( \39077 , \12857 );
or \U$38701 ( \39078 , \39076 , \39077 );
or \U$38702 ( \39079 , \12857 , \10584 );
nand \U$38703 ( \39080 , \39078 , \39079 );
not \U$38704 ( \39081 , \39080 );
not \U$38705 ( \39082 , \2416 );
or \U$38706 ( \39083 , \39081 , \39082 );
or \U$38707 ( \39084 , \38535 , \2410 );
nand \U$38708 ( \39085 , \39083 , \39084 );
not \U$38709 ( \39086 , \39085 );
nand \U$38710 ( \39087 , \12857 , \2408 );
nand \U$38711 ( \39088 , \39087 , \2409 , RIae79c28_161);
not \U$38712 ( \39089 , \39088 );
and \U$38713 ( \39090 , \39086 , \39089 );
and \U$38714 ( \39091 , \39085 , \39088 );
nor \U$38715 ( \39092 , \39090 , \39091 );
nand \U$38716 ( \39093 , \39075 , \39092 );
not \U$38717 ( \39094 , \39093 );
not \U$38718 ( \39095 , \6212 );
not \U$38719 ( \39096 , RIae79ef8_167);
not \U$38720 ( \39097 , \33414 );
or \U$38721 ( \39098 , \39096 , \39097 );
or \U$38722 ( \39099 , \11589 , RIae79ef8_167);
nand \U$38723 ( \39100 , \39098 , \39099 );
not \U$38724 ( \39101 , \39100 );
or \U$38725 ( \39102 , \39095 , \39101 );
nand \U$38726 ( \39103 , \38956 , \6199 );
nand \U$38727 ( \39104 , \39102 , \39103 );
not \U$38728 ( \39105 , \39104 );
or \U$38729 ( \39106 , \39094 , \39105 );
not \U$38730 ( \39107 , \39092 );
nand \U$38731 ( \39108 , \39107 , \39074 );
nand \U$38732 ( \39109 , \39106 , \39108 );
not \U$38733 ( \39110 , \39109 );
not \U$38734 ( \39111 , \39110 );
not \U$38735 ( \39112 , \10275 );
not \U$38736 ( \39113 , RIae7a8d0_188);
not \U$38737 ( \39114 , \6238 );
or \U$38738 ( \39115 , \39113 , \39114 );
or \U$38739 ( \39116 , \6244 , RIae7a8d0_188);
nand \U$38740 ( \39117 , \39115 , \39116 );
not \U$38741 ( \39118 , \39117 );
or \U$38742 ( \39119 , \39112 , \39118 );
not \U$38743 ( \39120 , RIae7a8d0_188);
not \U$38744 ( \39121 , \10829 );
or \U$38745 ( \39122 , \39120 , \39121 );
or \U$38746 ( \39123 , \10226 , RIae7a8d0_188);
nand \U$38747 ( \39124 , \39122 , \39123 );
nand \U$38748 ( \39125 , \39124 , \14510 );
nand \U$38749 ( \39126 , \39119 , \39125 );
not \U$38750 ( \39127 , \39126 );
or \U$38751 ( \39128 , \39111 , \39127 );
or \U$38752 ( \39129 , \39126 , \39110 );
nand \U$38753 ( \39130 , \39128 , \39129 );
not \U$38754 ( \39131 , \39130 );
or \U$38755 ( \39132 , \39069 , \39131 );
nand \U$38756 ( \39133 , \39126 , \39109 );
nand \U$38757 ( \39134 , \39132 , \39133 );
not \U$38758 ( \39135 , \39134 );
not \U$38759 ( \39136 , \38844 );
or \U$38760 ( \39137 , \38866 , \39136 );
nand \U$38761 ( \39138 , \38855 , \38861 );
nand \U$38762 ( \39139 , \39137 , \39138 );
not \U$38763 ( \39140 , \39139 );
xnor \U$38764 ( \39141 , \38554 , \38515 );
not \U$38765 ( \39142 , \39141 );
and \U$38766 ( \39143 , \39140 , \39142 );
and \U$38767 ( \39144 , \39139 , \39141 );
nor \U$38768 ( \39145 , \39143 , \39144 );
not \U$38769 ( \39146 , \39145 );
and \U$38770 ( \39147 , \39135 , \39146 );
and \U$38771 ( \39148 , \39134 , \39145 );
nor \U$38772 ( \39149 , \39147 , \39148 );
not \U$38773 ( \39150 , \39149 );
not \U$38774 ( \39151 , \39150 );
not \U$38775 ( \39152 , \39104 );
not \U$38776 ( \39153 , \39092 );
not \U$38777 ( \39154 , \39074 );
or \U$38778 ( \39155 , \39153 , \39154 );
or \U$38779 ( \39156 , \39074 , \39092 );
nand \U$38780 ( \39157 , \39155 , \39156 );
not \U$38781 ( \39158 , \39157 );
and \U$38782 ( \39159 , \39152 , \39158 );
and \U$38783 ( \39160 , \39104 , \39157 );
nor \U$38784 ( \39161 , \39159 , \39160 );
not \U$38785 ( \39162 , \10631 );
not \U$38786 ( \39163 , \38842 );
or \U$38787 ( \39164 , \39162 , \39163 );
and \U$38788 ( \39165 , RIae7a510_180, \9941 );
not \U$38789 ( \39166 , RIae7a510_180);
and \U$38790 ( \39167 , \39166 , \10465 );
or \U$38791 ( \39168 , \39165 , \39167 );
nand \U$38792 ( \39169 , \39168 , \10637 );
nand \U$38793 ( \39170 , \39164 , \39169 );
nor \U$38794 ( \39171 , \39161 , \39170 );
not \U$38795 ( \39172 , \39171 );
not \U$38796 ( \39173 , \39172 );
not \U$38797 ( \39174 , \10275 );
not \U$38798 ( \39175 , \39124 );
or \U$38799 ( \39176 , \39174 , \39175 );
not \U$38800 ( \39177 , RIae7a8d0_188);
not \U$38801 ( \39178 , \5108 );
or \U$38802 ( \39179 , \39177 , \39178 );
or \U$38803 ( \39180 , \27827 , RIae7a8d0_188);
nand \U$38804 ( \39181 , \39179 , \39180 );
nand \U$38805 ( \39182 , \39181 , \17847 );
nand \U$38806 ( \39183 , \39176 , \39182 );
not \U$38807 ( \39184 , \39183 );
or \U$38808 ( \39185 , \39173 , \39184 );
nand \U$38809 ( \39186 , \39161 , \39170 );
nand \U$38810 ( \39187 , \39185 , \39186 );
not \U$38811 ( \39188 , \39085 );
nor \U$38812 ( \39189 , \39188 , \39088 );
not \U$38813 ( \39190 , \5048 );
not \U$38814 ( \39191 , \38293 );
or \U$38815 ( \39192 , \39190 , \39191 );
nand \U$38816 ( \39193 , \38724 , \5039 );
nand \U$38817 ( \39194 , \39192 , \39193 );
xor \U$38818 ( \39195 , \39189 , \39194 );
not \U$38819 ( \39196 , \19362 );
not \U$38820 ( \39197 , \39100 );
or \U$38821 ( \39198 , \39196 , \39197 );
or \U$38822 ( \39199 , \38580 , \6213 );
nand \U$38823 ( \39200 , \39198 , \39199 );
xor \U$38824 ( \39201 , \39195 , \39200 );
not \U$38825 ( \39202 , \9478 );
not \U$38826 ( \39203 , RIae7a6f0_184);
not \U$38827 ( \39204 , \15128 );
or \U$38828 ( \39205 , \39203 , \39204 );
or \U$38829 ( \39206 , \16310 , RIae7a6f0_184);
nand \U$38830 ( \39207 , \39205 , \39206 );
not \U$38831 ( \39208 , \39207 );
or \U$38832 ( \39209 , \39202 , \39208 );
nand \U$38833 ( \39210 , \38898 , \9473 );
nand \U$38834 ( \39211 , \39209 , \39210 );
xor \U$38835 ( \39212 , \39201 , \39211 );
not \U$38836 ( \39213 , \11434 );
and \U$38837 ( \39214 , \16766 , \10625 );
not \U$38838 ( \39215 , \16766 );
and \U$38839 ( \39216 , \39215 , RIae7a498_179);
nor \U$38840 ( \39217 , \39214 , \39216 );
not \U$38841 ( \39218 , \39217 );
or \U$38842 ( \39219 , \39213 , \39218 );
nand \U$38843 ( \39220 , \38699 , \11422 );
nand \U$38844 ( \39221 , \39219 , \39220 );
xor \U$38845 ( \39222 , \39212 , \39221 );
xor \U$38846 ( \39223 , \39187 , \39222 );
xor \U$38847 ( \39224 , \39109 , \39068 );
xor \U$38848 ( \39225 , \39224 , \39126 );
and \U$38849 ( \39226 , \39223 , \39225 );
and \U$38850 ( \39227 , \39187 , \39222 );
or \U$38851 ( \39228 , \39226 , \39227 );
not \U$38852 ( \39229 , \39228 );
not \U$38853 ( \39230 , \39229 );
or \U$38854 ( \39231 , \39151 , \39230 );
nand \U$38855 ( \39232 , \39149 , \39228 );
nand \U$38856 ( \39233 , \39231 , \39232 );
not \U$38857 ( \39234 , \39233 );
or \U$38858 ( \39235 , \39059 , \39234 );
nand \U$38859 ( \39236 , \39150 , \39228 );
nand \U$38860 ( \39237 , \39235 , \39236 );
not \U$38861 ( \39238 , \39237 );
or \U$38862 ( \39239 , \39014 , \39238 );
not \U$38863 ( \39240 , \38720 );
nand \U$38864 ( \39241 , \39240 , \39008 );
nand \U$38865 ( \39242 , \39239 , \39241 );
xor \U$38866 ( \39243 , \38374 , \38383 );
xor \U$38867 ( \39244 , \39243 , \38393 );
not \U$38868 ( \39245 , \39244 );
xor \U$38869 ( \39246 , \38229 , \38238 );
xor \U$38870 ( \39247 , \39246 , \38249 );
not \U$38871 ( \39248 , \39247 );
and \U$38872 ( \39249 , \39245 , \39248 );
and \U$38873 ( \39250 , \39247 , \39244 );
not \U$38874 ( \39251 , \9549 );
not \U$38875 ( \39252 , \39064 );
or \U$38876 ( \39253 , \39251 , \39252 );
nand \U$38877 ( \39254 , \38307 , \29519 );
nand \U$38878 ( \39255 , \39253 , \39254 );
not \U$38879 ( \39256 , \39255 );
not \U$38880 ( \39257 , \9777 );
not \U$38881 ( \39258 , \38264 );
or \U$38882 ( \39259 , \39257 , \39258 );
nand \U$38883 ( \39260 , \39034 , \11087 );
nand \U$38884 ( \39261 , \39259 , \39260 );
not \U$38885 ( \39262 , \39261 );
or \U$38886 ( \39263 , \39256 , \39262 );
or \U$38887 ( \39264 , \39261 , \39255 );
not \U$38888 ( \39265 , \9705 );
not \U$38889 ( \39266 , \38479 );
or \U$38890 ( \39267 , \39265 , \39266 );
nand \U$38891 ( \39268 , \39207 , \35747 );
nand \U$38892 ( \39269 , \39267 , \39268 );
nand \U$38893 ( \39270 , \39264 , \39269 );
nand \U$38894 ( \39271 , \39263 , \39270 );
nor \U$38895 ( \39272 , \39250 , \39271 );
nor \U$38896 ( \39273 , \39249 , \39272 );
xor \U$38897 ( \39274 , \38347 , \38351 );
xor \U$38898 ( \39275 , \39274 , \38359 );
xor \U$38899 ( \39276 , \39273 , \39275 );
not \U$38900 ( \39277 , \38715 );
not \U$38901 ( \39278 , \38712 );
or \U$38902 ( \39279 , \39277 , \39278 );
nand \U$38903 ( \39280 , \38706 , \38711 );
nand \U$38904 ( \39281 , \39279 , \39280 );
xor \U$38905 ( \39282 , \39276 , \39281 );
not \U$38906 ( \39283 , \39282 );
nand \U$38907 ( \39284 , \39021 , \39022 );
and \U$38908 ( \39285 , \39027 , \39284 );
nor \U$38909 ( \39286 , \39021 , \39022 );
nor \U$38910 ( \39287 , \39285 , \39286 );
xor \U$38911 ( \39288 , \38413 , \38424 );
xor \U$38912 ( \39289 , \39288 , \38435 );
xor \U$38913 ( \39290 , \39287 , \39289 );
not \U$38914 ( \39291 , \39200 );
not \U$38915 ( \39292 , \39195 );
or \U$38916 ( \39293 , \39291 , \39292 );
nand \U$38917 ( \39294 , \39194 , \39189 );
nand \U$38918 ( \39295 , \39293 , \39294 );
not \U$38919 ( \39296 , \9744 );
not \U$38920 ( \39297 , \38381 );
or \U$38921 ( \39298 , \39296 , \39297 );
nand \U$38922 ( \39299 , \39045 , \9729 );
nand \U$38923 ( \39300 , \39298 , \39299 );
xor \U$38924 ( \39301 , \39295 , \39300 );
not \U$38925 ( \39302 , \39301 );
not \U$38926 ( \39303 , \14510 );
not \U$38927 ( \39304 , \39117 );
or \U$38928 ( \39305 , \39303 , \39304 );
nand \U$38929 ( \39306 , \38389 , \10275 );
nand \U$38930 ( \39307 , \39305 , \39306 );
not \U$38931 ( \39308 , \39307 );
or \U$38932 ( \39309 , \39302 , \39308 );
nand \U$38933 ( \39310 , \39300 , \39295 );
nand \U$38934 ( \39311 , \39309 , \39310 );
xor \U$38935 ( \39312 , \39290 , \39311 );
not \U$38936 ( \39313 , \39312 );
not \U$38937 ( \39314 , \39145 );
not \U$38938 ( \39315 , \39314 );
not \U$38939 ( \39316 , \39134 );
or \U$38940 ( \39317 , \39315 , \39316 );
not \U$38941 ( \39318 , \39141 );
nand \U$38942 ( \39319 , \39318 , \39139 );
nand \U$38943 ( \39320 , \39317 , \39319 );
not \U$38944 ( \39321 , \38503 );
not \U$38945 ( \39322 , \38559 );
or \U$38946 ( \39323 , \39321 , \39322 );
or \U$38947 ( \39324 , \38559 , \38503 );
nand \U$38948 ( \39325 , \39323 , \39324 );
xor \U$38949 ( \39326 , \38598 , \39325 );
xor \U$38950 ( \39327 , \39320 , \39326 );
not \U$38951 ( \39328 , \39327 );
or \U$38952 ( \39329 , \39313 , \39328 );
nand \U$38953 ( \39330 , \39320 , \39326 );
nand \U$38954 ( \39331 , \39329 , \39330 );
not \U$38955 ( \39332 , \39331 );
not \U$38956 ( \39333 , \39332 );
or \U$38957 ( \39334 , \39283 , \39333 );
or \U$38958 ( \39335 , \39332 , \39282 );
nand \U$38959 ( \39336 , \39334 , \39335 );
xor \U$38960 ( \39337 , \39242 , \39336 );
not \U$38961 ( \39338 , \39337 );
xor \U$38962 ( \39339 , \38602 , \38466 );
xnor \U$38963 ( \39340 , \39339 , \38501 );
not \U$38964 ( \39341 , \38258 );
not \U$38965 ( \39342 , \38314 );
not \U$38966 ( \39343 , \39342 );
or \U$38967 ( \39344 , \39341 , \39343 );
or \U$38968 ( \39345 , \39342 , \38258 );
nand \U$38969 ( \39346 , \39344 , \39345 );
xor \U$38970 ( \39347 , \39287 , \39289 );
and \U$38971 ( \39348 , \39347 , \39311 );
and \U$38972 ( \39349 , \39287 , \39289 );
or \U$38973 ( \39350 , \39348 , \39349 );
xor \U$38974 ( \39351 , \39346 , \39350 );
buf \U$38975 ( \39352 , \38442 );
and \U$38976 ( \39353 , \39352 , \38396 );
not \U$38977 ( \39354 , \39352 );
not \U$38978 ( \39355 , \38396 );
and \U$38979 ( \39356 , \39354 , \39355 );
nor \U$38980 ( \39357 , \39353 , \39356 );
and \U$38981 ( \39358 , \39351 , \39357 );
not \U$38982 ( \39359 , \39351 );
not \U$38983 ( \39360 , \39357 );
and \U$38984 ( \39361 , \39359 , \39360 );
nor \U$38985 ( \39362 , \39358 , \39361 );
xor \U$38986 ( \39363 , \39340 , \39362 );
not \U$38987 ( \39364 , \39301 );
and \U$38988 ( \39365 , \39307 , \39364 );
not \U$38989 ( \39366 , \39307 );
and \U$38990 ( \39367 , \39366 , \39301 );
nor \U$38991 ( \39368 , \39365 , \39367 );
xor \U$38992 ( \39369 , \39201 , \39211 );
and \U$38993 ( \39370 , \39369 , \39221 );
and \U$38994 ( \39371 , \39201 , \39211 );
nor \U$38995 ( \39372 , \39370 , \39371 );
xor \U$38996 ( \39373 , \39368 , \39372 );
xor \U$38997 ( \39374 , \39255 , \39261 );
xnor \U$38998 ( \39375 , \39374 , \39269 );
and \U$38999 ( \39376 , \39373 , \39375 );
and \U$39000 ( \39377 , \39368 , \39372 );
or \U$39001 ( \39378 , \39376 , \39377 );
not \U$39002 ( \39379 , \39378 );
xor \U$39003 ( \39380 , \39247 , \39271 );
xnor \U$39004 ( \39381 , \39380 , \39244 );
not \U$39005 ( \39382 , \39381 );
or \U$39006 ( \39383 , \39379 , \39382 );
not \U$39007 ( \39384 , \39028 );
not \U$39008 ( \39385 , \39016 );
not \U$39009 ( \39386 , \39056 );
or \U$39010 ( \39387 , \39385 , \39386 );
or \U$39011 ( \39388 , \39056 , \39016 );
nand \U$39012 ( \39389 , \39387 , \39388 );
not \U$39013 ( \39390 , \39389 );
or \U$39014 ( \39391 , \39384 , \39390 );
not \U$39015 ( \39392 , \39016 );
nand \U$39016 ( \39393 , \39392 , \39056 );
nand \U$39017 ( \39394 , \39391 , \39393 );
nand \U$39018 ( \39395 , \39383 , \39394 );
not \U$39019 ( \39396 , \39378 );
not \U$39020 ( \39397 , \39381 );
nand \U$39021 ( \39398 , \39396 , \39397 );
nand \U$39022 ( \39399 , \39395 , \39398 );
xnor \U$39023 ( \39400 , \39363 , \39399 );
not \U$39024 ( \39401 , \39400 );
not \U$39025 ( \39402 , \39401 );
xor \U$39026 ( \39403 , \39326 , \39312 );
xnor \U$39027 ( \39404 , \39403 , \39320 );
xor \U$39028 ( \39405 , \39378 , \39397 );
not \U$39029 ( \39406 , \39394 );
xnor \U$39030 ( \39407 , \39405 , \39406 );
nand \U$39031 ( \39408 , \39404 , \39407 );
not \U$39032 ( \39409 , \39408 );
not \U$39033 ( \39410 , \39012 );
not \U$39034 ( \39411 , \39237 );
or \U$39035 ( \39412 , \39410 , \39411 );
or \U$39036 ( \39413 , \39237 , \39012 );
nand \U$39037 ( \39414 , \39412 , \39413 );
not \U$39038 ( \39415 , \39414 );
or \U$39039 ( \39416 , \39409 , \39415 );
not \U$39040 ( \39417 , \39404 );
not \U$39041 ( \39418 , \39407 );
nand \U$39042 ( \39419 , \39417 , \39418 );
nand \U$39043 ( \39420 , \39416 , \39419 );
not \U$39044 ( \39421 , \39420 );
not \U$39045 ( \39422 , \39421 );
or \U$39046 ( \39423 , \39402 , \39422 );
nand \U$39047 ( \39424 , \39420 , \39400 );
nand \U$39048 ( \39425 , \39423 , \39424 );
not \U$39049 ( \39426 , \39425 );
or \U$39050 ( \39427 , \39338 , \39426 );
nand \U$39051 ( \39428 , \39420 , \39401 );
nand \U$39052 ( \39429 , \39427 , \39428 );
not \U$39053 ( \39430 , \39429 );
xor \U$39054 ( \39431 , \38319 , \38227 );
not \U$39055 ( \39432 , \39357 );
not \U$39056 ( \39433 , \39351 );
or \U$39057 ( \39434 , \39432 , \39433 );
nand \U$39058 ( \39435 , \39350 , \39346 );
nand \U$39059 ( \39436 , \39434 , \39435 );
xor \U$39060 ( \39437 , \39431 , \39436 );
xor \U$39061 ( \39438 , \39273 , \39275 );
and \U$39062 ( \39439 , \39438 , \39281 );
and \U$39063 ( \39440 , \39273 , \39275 );
or \U$39064 ( \39441 , \39439 , \39440 );
and \U$39065 ( \39442 , \39437 , \39441 );
not \U$39066 ( \39443 , \39437 );
not \U$39067 ( \39444 , \39441 );
and \U$39068 ( \39445 , \39443 , \39444 );
nor \U$39069 ( \39446 , \39442 , \39445 );
not \U$39070 ( \39447 , \39242 );
not \U$39071 ( \39448 , \39336 );
or \U$39072 ( \39449 , \39447 , \39448 );
nand \U$39073 ( \39450 , \39331 , \39282 );
nand \U$39074 ( \39451 , \39449 , \39450 );
xor \U$39075 ( \39452 , \39446 , \39451 );
buf \U$39076 ( \39453 , \38452 );
and \U$39077 ( \39454 , \39453 , \38344 );
not \U$39078 ( \39455 , \39453 );
not \U$39079 ( \39456 , \38344 );
and \U$39080 ( \39457 , \39455 , \39456 );
nor \U$39081 ( \39458 , \39454 , \39457 );
not \U$39082 ( \39459 , \39340 );
not \U$39083 ( \39460 , \39399 );
or \U$39084 ( \39461 , \39459 , \39460 );
or \U$39085 ( \39462 , \39399 , \39340 );
nand \U$39086 ( \39463 , \39462 , \39362 );
nand \U$39087 ( \39464 , \39461 , \39463 );
xor \U$39088 ( \39465 , \39458 , \39464 );
not \U$39089 ( \39466 , \38608 );
and \U$39090 ( \39467 , \38616 , \39466 );
not \U$39091 ( \39468 , \38616 );
and \U$39092 ( \39469 , \39468 , \38608 );
nor \U$39093 ( \39470 , \39467 , \39469 );
not \U$39094 ( \39471 , \39470 );
xnor \U$39095 ( \39472 , \39465 , \39471 );
xnor \U$39096 ( \39473 , \39452 , \39472 );
not \U$39097 ( \39474 , \39473 );
nand \U$39098 ( \39475 , \39430 , \39474 );
not \U$39099 ( \39476 , \39470 );
not \U$39100 ( \39477 , \39458 );
not \U$39101 ( \39478 , \39477 );
or \U$39102 ( \39479 , \39476 , \39478 );
nand \U$39103 ( \39480 , \39479 , \39464 );
not \U$39104 ( \39481 , \38457 );
not \U$39105 ( \39482 , \38343 );
or \U$39106 ( \39483 , \39481 , \39482 );
nand \U$39107 ( \39484 , \38342 , \38458 );
nand \U$39108 ( \39485 , \39483 , \39484 );
not \U$39109 ( \39486 , \39485 );
not \U$39110 ( \39487 , \38626 );
or \U$39111 ( \39488 , \39486 , \39487 );
or \U$39112 ( \39489 , \38626 , \39485 );
nand \U$39113 ( \39490 , \39488 , \39489 );
not \U$39114 ( \39491 , \39477 );
nand \U$39115 ( \39492 , \39491 , \39471 );
and \U$39116 ( \39493 , \39480 , \39490 , \39492 );
not \U$39117 ( \39494 , \39493 );
not \U$39118 ( \39495 , \39480 );
not \U$39119 ( \39496 , \39492 );
or \U$39120 ( \39497 , \39495 , \39496 );
not \U$39121 ( \39498 , \39490 );
nand \U$39122 ( \39499 , \39497 , \39498 );
nand \U$39123 ( \39500 , \39494 , \39499 );
xor \U$39124 ( \39501 , \38329 , \38211 );
not \U$39125 ( \39502 , \39501 );
xor \U$39126 ( \39503 , \38176 , \38179 );
xnor \U$39127 ( \39504 , \39503 , \38174 );
not \U$39128 ( \39505 , \39504 );
not \U$39129 ( \39506 , \39505 );
or \U$39130 ( \39507 , \39502 , \39506 );
not \U$39131 ( \39508 , \39501 );
nand \U$39132 ( \39509 , \39508 , \39504 );
nand \U$39133 ( \39510 , \39507 , \39509 );
not \U$39134 ( \39511 , \39441 );
not \U$39135 ( \39512 , \39437 );
or \U$39136 ( \39513 , \39511 , \39512 );
nand \U$39137 ( \39514 , \39436 , \39431 );
nand \U$39138 ( \39515 , \39513 , \39514 );
not \U$39139 ( \39516 , \39515 );
and \U$39140 ( \39517 , \39510 , \39516 );
not \U$39141 ( \39518 , \39510 );
and \U$39142 ( \39519 , \39518 , \39515 );
nor \U$39143 ( \39520 , \39517 , \39519 );
not \U$39144 ( \39521 , \39520 );
and \U$39145 ( \39522 , \39500 , \39521 );
not \U$39146 ( \39523 , \39500 );
and \U$39147 ( \39524 , \39523 , \39520 );
nor \U$39148 ( \39525 , \39522 , \39524 );
not \U$39149 ( \39526 , \39446 );
nand \U$39150 ( \39527 , \39472 , \39526 );
buf \U$39151 ( \39528 , \39451 );
and \U$39152 ( \39529 , \39527 , \39528 );
nor \U$39153 ( \39530 , \39472 , \39526 );
nor \U$39154 ( \39531 , \39529 , \39530 );
nand \U$39155 ( \39532 , \39525 , \39531 );
and \U$39156 ( \39533 , \39475 , \39532 );
not \U$39157 ( \39534 , \39533 );
buf \U$39158 ( \39535 , \39414 );
not \U$39159 ( \39536 , \39535 );
nand \U$39160 ( \39537 , \39419 , \39408 );
not \U$39161 ( \39538 , \39537 );
and \U$39162 ( \39539 , \39536 , \39538 );
and \U$39163 ( \39540 , \39535 , \39537 );
nor \U$39164 ( \39541 , \39539 , \39540 );
not \U$39165 ( \39542 , \39541 );
xor \U$39166 ( \39543 , \38970 , \38983 );
xor \U$39167 ( \39544 , \39543 , \38998 );
buf \U$39168 ( \39545 , \38805 );
xor \U$39169 ( \39546 , \38822 , \39545 );
or \U$39170 ( \39547 , \39544 , \39546 );
xor \U$39171 ( \39548 , \38893 , \38906 );
xor \U$39172 ( \39549 , \39548 , \38922 );
nand \U$39173 ( \39550 , \39547 , \39549 );
nand \U$39174 ( \39551 , \39544 , \39546 );
nand \U$39175 ( \39552 , \39550 , \39551 );
not \U$39176 ( \39553 , \39552 );
not \U$39177 ( \39554 , \10637 );
and \U$39178 ( \39555 , RIae7a510_180, \33592 );
not \U$39179 ( \39556 , RIae7a510_180);
and \U$39180 ( \39557 , \39556 , \13660 );
nor \U$39181 ( \39558 , \39555 , \39557 );
not \U$39182 ( \39559 , \39558 );
or \U$39183 ( \39560 , \39554 , \39559 );
nand \U$39184 ( \39561 , \39168 , \16358 );
nand \U$39185 ( \39562 , \39560 , \39561 );
not \U$39186 ( \39563 , \9792 );
and \U$39187 ( \39564 , \16193 , \29995 );
not \U$39188 ( \39565 , \16193 );
and \U$39189 ( \39566 , \39565 , RIae7a2b8_175);
nor \U$39190 ( \39567 , \39564 , \39566 );
not \U$39191 ( \39568 , \39567 );
or \U$39192 ( \39569 , \39563 , \39568 );
nand \U$39193 ( \39570 , \38799 , \9813 );
nand \U$39194 ( \39571 , \39569 , \39570 );
nor \U$39195 ( \39572 , \39562 , \39571 );
not \U$39196 ( \39573 , \39572 );
not \U$39197 ( \39574 , \39573 );
not \U$39198 ( \39575 , \11851 );
not \U$39199 ( \39576 , RIae7a7e0_186);
not \U$39200 ( \39577 , \21744 );
or \U$39201 ( \39578 , \39576 , \39577 );
nand \U$39202 ( \39579 , \15519 , \9529 );
nand \U$39203 ( \39580 , \39578 , \39579 );
not \U$39204 ( \39581 , \39580 );
or \U$39205 ( \39582 , \39575 , \39581 );
nand \U$39206 ( \39583 , \38981 , \9527 );
nand \U$39207 ( \39584 , \39582 , \39583 );
not \U$39208 ( \39585 , \39584 );
or \U$39209 ( \39586 , \39574 , \39585 );
nand \U$39210 ( \39587 , \39562 , \39571 );
nand \U$39211 ( \39588 , \39586 , \39587 );
not \U$39212 ( \39589 , \10667 );
not \U$39213 ( \39590 , RIae7a150_172);
not \U$39214 ( \39591 , \22560 );
or \U$39215 ( \39592 , \39590 , \39591 );
or \U$39216 ( \39593 , \16766 , RIae7a150_172);
nand \U$39217 ( \39594 , \39592 , \39593 );
not \U$39218 ( \39595 , \39594 );
or \U$39219 ( \39596 , \39589 , \39595 );
nand \U$39220 ( \39597 , \38891 , \9776 );
nand \U$39221 ( \39598 , \39596 , \39597 );
not \U$39222 ( \39599 , \39598 );
not \U$39223 ( \39600 , \11098 );
not \U$39224 ( \39601 , \38996 );
or \U$39225 ( \39602 , \39600 , \39601 );
not \U$39226 ( \39603 , \11102 );
not \U$39227 ( \39604 , \12614 );
or \U$39228 ( \39605 , \39603 , \39604 );
or \U$39229 ( \39606 , \14110 , \9749 );
nand \U$39230 ( \39607 , \39605 , \39606 );
nand \U$39231 ( \39608 , \39607 , \9730 );
nand \U$39232 ( \39609 , \39602 , \39608 );
not \U$39233 ( \39610 , \9705 );
not \U$39234 ( \39611 , \38904 );
or \U$39235 ( \39612 , \39610 , \39611 );
and \U$39236 ( \39613 , RIae7a6f0_184, \12683 );
not \U$39237 ( \39614 , RIae7a6f0_184);
and \U$39238 ( \39615 , \39614 , \9298 );
or \U$39239 ( \39616 , \39613 , \39615 );
nand \U$39240 ( \39617 , \39616 , \9473 );
nand \U$39241 ( \39618 , \39612 , \39617 );
nand \U$39242 ( \39619 , \39609 , \39618 );
nand \U$39243 ( \39620 , \39599 , \39619 );
or \U$39244 ( \39621 , \39609 , \39618 );
and \U$39245 ( \39622 , \39620 , \39621 );
nor \U$39246 ( \39623 , \39588 , \39622 );
not \U$39247 ( \39624 , \38946 );
not \U$39248 ( \39625 , \38949 );
and \U$39249 ( \39626 , \39624 , \39625 );
and \U$39250 ( \39627 , \38946 , \38949 );
nor \U$39251 ( \39628 , \39626 , \39627 );
not \U$39252 ( \39629 , \39628 );
not \U$39253 ( \39630 , \5048 );
not \U$39254 ( \39631 , \38740 );
or \U$39255 ( \39632 , \39630 , \39631 );
and \U$39256 ( \39633 , \16651 , \13059 );
not \U$39257 ( \39634 , \16651 );
and \U$39258 ( \39635 , \39634 , RIae79d90_164);
nor \U$39259 ( \39636 , \39633 , \39635 );
nand \U$39260 ( \39637 , \39636 , \5039 );
nand \U$39261 ( \39638 , \39632 , \39637 );
not \U$39262 ( \39639 , \39638 );
or \U$39263 ( \39640 , \39629 , \39639 );
or \U$39264 ( \39641 , \39638 , \39628 );
nand \U$39265 ( \39642 , \39640 , \39641 );
not \U$39266 ( \39643 , \39642 );
not \U$39267 ( \39644 , \9517 );
not \U$39268 ( \39645 , \38931 );
or \U$39269 ( \39646 , \39644 , \39645 );
not \U$39270 ( \39647 , \18027 );
not \U$39271 ( \39648 , \10042 );
or \U$39272 ( \39649 , \39647 , \39648 );
or \U$39273 ( \39650 , \10042 , \11069 );
nand \U$39274 ( \39651 , \39649 , \39650 );
nand \U$39275 ( \39652 , \39651 , \9499 );
nand \U$39276 ( \39653 , \39646 , \39652 );
not \U$39277 ( \39654 , \39653 );
or \U$39278 ( \39655 , \39643 , \39654 );
not \U$39279 ( \39656 , \39628 );
nand \U$39280 ( \39657 , \39656 , \39638 );
nand \U$39281 ( \39658 , \39655 , \39657 );
not \U$39282 ( \39659 , \10275 );
not \U$39283 ( \39660 , \39181 );
or \U$39284 ( \39661 , \39659 , \39660 );
not \U$39285 ( \39662 , \18088 );
not \U$39286 ( \39663 , \9279 );
or \U$39287 ( \39664 , \39662 , \39663 );
or \U$39288 ( \39665 , \5722 , \11207 );
nand \U$39289 ( \39666 , \39664 , \39665 );
nand \U$39290 ( \39667 , \39666 , \16594 );
nand \U$39291 ( \39668 , \39661 , \39667 );
xor \U$39292 ( \39669 , \39658 , \39668 );
not \U$39293 ( \39670 , RIae7aab0_192);
not \U$39294 ( \39671 , \38913 );
or \U$39295 ( \39672 , \39670 , \39671 );
and \U$39296 ( \39673 , RIae7aa38_191, \10226 );
not \U$39297 ( \39674 , RIae7aa38_191);
and \U$39298 ( \39675 , \39674 , \12724 );
or \U$39299 ( \39676 , \39673 , \39675 );
nand \U$39300 ( \39677 , \39676 , \14669 );
nand \U$39301 ( \39678 , \39672 , \39677 );
and \U$39302 ( \39679 , \39669 , \39678 );
and \U$39303 ( \39680 , \39658 , \39668 );
nor \U$39304 ( \39681 , \39679 , \39680 );
or \U$39305 ( \39682 , \39623 , \39681 );
nand \U$39306 ( \39683 , \39588 , \39622 );
nand \U$39307 ( \39684 , \39682 , \39683 );
xor \U$39308 ( \39685 , \38878 , \39001 );
xnor \U$39309 ( \39686 , \39685 , \38925 );
not \U$39310 ( \39687 , \39686 );
xor \U$39311 ( \39688 , \39684 , \39687 );
not \U$39312 ( \39689 , \39688 );
or \U$39313 ( \39690 , \39553 , \39689 );
not \U$39314 ( \39691 , \39686 );
nand \U$39315 ( \39692 , \39691 , \39684 );
nand \U$39316 ( \39693 , \39690 , \39692 );
not \U$39317 ( \39694 , \39693 );
xor \U$39318 ( \39695 , \39368 , \39372 );
xor \U$39319 ( \39696 , \39695 , \39375 );
not \U$39320 ( \39697 , \39696 );
buf \U$39321 ( \39698 , \38870 );
buf \U$39322 ( \39699 , \38831 );
not \U$39323 ( \39700 , \39699 );
and \U$39324 ( \39701 , \39698 , \39700 );
not \U$39325 ( \39702 , \39698 );
and \U$39326 ( \39703 , \39702 , \39699 );
nor \U$39327 ( \39704 , \39701 , \39703 );
not \U$39328 ( \39705 , \39704 );
not \U$39329 ( \39706 , \39705 );
xor \U$39330 ( \39707 , \38733 , \38768 );
xor \U$39331 ( \39708 , \39707 , \38778 );
not \U$39332 ( \39709 , \10676 );
not \U$39333 ( \39710 , \39217 );
or \U$39334 ( \39711 , \39709 , \39710 );
not \U$39335 ( \39712 , \10625 );
not \U$39336 ( \39713 , \15947 );
or \U$39337 ( \39714 , \39712 , \39713 );
or \U$39338 ( \39715 , \11803 , \10625 );
nand \U$39339 ( \39716 , \39714 , \39715 );
nand \U$39340 ( \39717 , \39716 , \16564 );
nand \U$39341 ( \39718 , \39711 , \39717 );
xor \U$39342 ( \39719 , \39708 , \39718 );
not \U$39343 ( \39720 , \9644 );
and \U$39344 ( \39721 , \13905 , RIae7a3a8_177);
not \U$39345 ( \39722 , \13905 );
and \U$39346 ( \39723 , \39722 , \16469 );
nor \U$39347 ( \39724 , \39721 , \39723 );
not \U$39348 ( \39725 , \39724 );
or \U$39349 ( \39726 , \39720 , \39725 );
nand \U$39350 ( \39727 , \38820 , \9622 );
nand \U$39351 ( \39728 , \39726 , \39727 );
not \U$39352 ( \39729 , \39728 );
not \U$39353 ( \39730 , \38742 );
and \U$39354 ( \39731 , \38763 , \39730 );
not \U$39355 ( \39732 , \38763 );
and \U$39356 ( \39733 , \39732 , \38742 );
nor \U$39357 ( \39734 , \39731 , \39733 );
not \U$39358 ( \39735 , \39734 );
not \U$39359 ( \39736 , \9687 );
not \U$39360 ( \39737 , RIae7a240_174);
not \U$39361 ( \39738 , \9875 );
or \U$39362 ( \39739 , \39737 , \39738 );
or \U$39363 ( \39740 , \9875 , RIae7a240_174);
nand \U$39364 ( \39741 , \39739 , \39740 );
not \U$39365 ( \39742 , \39741 );
or \U$39366 ( \39743 , \39736 , \39742 );
nand \U$39367 ( \39744 , \38776 , \9699 );
nand \U$39368 ( \39745 , \39743 , \39744 );
not \U$39369 ( \39746 , \39745 );
or \U$39370 ( \39747 , \39735 , \39746 );
or \U$39371 ( \39748 , \39745 , \39734 );
nand \U$39372 ( \39749 , \39747 , \39748 );
not \U$39373 ( \39750 , \39749 );
or \U$39374 ( \39751 , \39729 , \39750 );
not \U$39375 ( \39752 , \39734 );
nand \U$39376 ( \39753 , \39752 , \39745 );
nand \U$39377 ( \39754 , \39751 , \39753 );
and \U$39378 ( \39755 , \39719 , \39754 );
and \U$39379 ( \39756 , \39708 , \39718 );
or \U$39380 ( \39757 , \39755 , \39756 );
xor \U$39381 ( \39758 , \39038 , \39047 );
xor \U$39382 ( \39759 , \39758 , \39053 );
xor \U$39383 ( \39760 , \39757 , \39759 );
not \U$39384 ( \39761 , \39760 );
or \U$39385 ( \39762 , \39706 , \39761 );
nand \U$39386 ( \39763 , \39759 , \39757 );
nand \U$39387 ( \39764 , \39762 , \39763 );
not \U$39388 ( \39765 , \39764 );
or \U$39389 ( \39766 , \39697 , \39765 );
or \U$39390 ( \39767 , \39764 , \39696 );
nand \U$39391 ( \39768 , \39766 , \39767 );
not \U$39392 ( \39769 , \39768 );
or \U$39393 ( \39770 , \39694 , \39769 );
not \U$39394 ( \39771 , \39696 );
nand \U$39395 ( \39772 , \39771 , \39764 );
nand \U$39396 ( \39773 , \39770 , \39772 );
not \U$39397 ( \39774 , \39773 );
xor \U$39398 ( \39775 , \38876 , \39004 );
xor \U$39399 ( \39776 , \39057 , \39775 );
xnor \U$39400 ( \39777 , \39776 , \39233 );
not \U$39401 ( \39778 , \9621 );
not \U$39402 ( \39779 , \39724 );
or \U$39403 ( \39780 , \39778 , \39779 );
not \U$39404 ( \39781 , \11690 );
not \U$39405 ( \39782 , \36204 );
or \U$39406 ( \39783 , \39781 , \39782 );
nand \U$39407 ( \39784 , \10171 , RIae7a3a8_177);
nand \U$39408 ( \39785 , \39783 , \39784 );
nand \U$39409 ( \39786 , \39785 , \9643 );
nand \U$39410 ( \39787 , \39780 , \39786 );
not \U$39411 ( \39788 , \39787 );
not \U$39412 ( \39789 , \38963 );
or \U$39413 ( \39790 , \39789 , \6213 );
not \U$39414 ( \39791 , \6203 );
not \U$39415 ( \39792 , \11321 );
or \U$39416 ( \39793 , \39791 , \39792 );
or \U$39417 ( \39794 , \11318 , \6207 );
nand \U$39418 ( \39795 , \39793 , \39794 );
not \U$39419 ( \39796 , \39795 );
not \U$39420 ( \39797 , \6200 );
or \U$39421 ( \39798 , \39796 , \39797 );
nand \U$39422 ( \39799 , \39790 , \39798 );
not \U$39423 ( \39800 , \6212 );
not \U$39424 ( \39801 , \39795 );
or \U$39425 ( \39802 , \39800 , \39801 );
not \U$39426 ( \39803 , \6207 );
not \U$39427 ( \39804 , \18971 );
or \U$39428 ( \39805 , \39803 , \39804 );
buf \U$39429 ( \39806 , \10259 );
nand \U$39430 ( \39807 , \39806 , RIae79ef8_167);
nand \U$39431 ( \39808 , \39805 , \39807 );
nand \U$39432 ( \39809 , \39808 , \6199 );
nand \U$39433 ( \39810 , \39802 , \39809 );
not \U$39434 ( \39811 , \39810 );
nand \U$39435 ( \39812 , \12857 , \4155 );
not \U$39436 ( \39813 , \39812 );
not \U$39437 ( \39814 , \5048 );
not \U$39438 ( \39815 , \39636 );
or \U$39439 ( \39816 , \39814 , \39815 );
not \U$39440 ( \39817 , RIae79d90_164);
not \U$39441 ( \39818 , \12750 );
or \U$39442 ( \39819 , \39817 , \39818 );
or \U$39443 ( \39820 , \16006 , RIae79d90_164);
nand \U$39444 ( \39821 , \39819 , \39820 );
nand \U$39445 ( \39822 , \39821 , \5039 );
nand \U$39446 ( \39823 , \39816 , \39822 );
not \U$39447 ( \39824 , \39823 );
or \U$39448 ( \39825 , \39813 , \39824 );
or \U$39449 ( \39826 , \39823 , \39812 );
nand \U$39450 ( \39827 , \39825 , \39826 );
not \U$39451 ( \39828 , \39827 );
or \U$39452 ( \39829 , \39811 , \39828 );
not \U$39453 ( \39830 , \39812 );
nand \U$39454 ( \39831 , \39830 , \39823 );
nand \U$39455 ( \39832 , \39829 , \39831 );
xor \U$39456 ( \39833 , \39799 , \39832 );
not \U$39457 ( \39834 , \39833 );
or \U$39458 ( \39835 , \39788 , \39834 );
nand \U$39459 ( \39836 , \39832 , \39799 );
nand \U$39460 ( \39837 , \39835 , \39836 );
not \U$39461 ( \39838 , \39837 );
not \U$39462 ( \39839 , \10695 );
and \U$39463 ( \39840 , RIae7a498_179, \9607 );
not \U$39464 ( \39841 , RIae7a498_179);
and \U$39465 ( \39842 , \39841 , \12483 );
nor \U$39466 ( \39843 , \39840 , \39842 );
not \U$39467 ( \39844 , \39843 );
or \U$39468 ( \39845 , \39839 , \39844 );
nand \U$39469 ( \39846 , \39716 , \10675 );
nand \U$39470 ( \39847 , \39845 , \39846 );
not \U$39471 ( \39848 , \39847 );
not \U$39472 ( \39849 , \38935 );
not \U$39473 ( \39850 , \39849 );
not \U$39474 ( \39851 , \38966 );
or \U$39475 ( \39852 , \39850 , \39851 );
or \U$39476 ( \39853 , \38966 , \39849 );
nand \U$39477 ( \39854 , \39852 , \39853 );
not \U$39478 ( \39855 , \39854 );
not \U$39479 ( \39856 , \39855 );
or \U$39480 ( \39857 , \39848 , \39856 );
not \U$39481 ( \39858 , \39847 );
nand \U$39482 ( \39859 , \39858 , \39854 );
nand \U$39483 ( \39860 , \39857 , \39859 );
not \U$39484 ( \39861 , \39860 );
or \U$39485 ( \39862 , \39838 , \39861 );
nand \U$39486 ( \39863 , \39854 , \39847 );
nand \U$39487 ( \39864 , \39862 , \39863 );
not \U$39488 ( \39865 , \39864 );
not \U$39489 ( \39866 , \39865 );
not \U$39490 ( \39867 , \39866 );
not \U$39491 ( \39868 , \39171 );
nand \U$39492 ( \39869 , \39868 , \39186 );
xnor \U$39493 ( \39870 , \39183 , \39869 );
not \U$39494 ( \39871 , \39870 );
or \U$39495 ( \39872 , \39867 , \39871 );
or \U$39496 ( \39873 , \39870 , \39866 );
xor \U$39497 ( \39874 , \39749 , \39728 );
not \U$39498 ( \39875 , \39874 );
not \U$39499 ( \39876 , \10542 );
not \U$39500 ( \39877 , \39607 );
or \U$39501 ( \39878 , \39876 , \39877 );
and \U$39502 ( \39879 , \9455 , RIae7a060_170);
not \U$39503 ( \39880 , \9455 );
and \U$39504 ( \39881 , \39880 , \9749 );
nor \U$39505 ( \39882 , \39879 , \39881 );
nand \U$39506 ( \39883 , \39882 , \9729 );
nand \U$39507 ( \39884 , \39878 , \39883 );
not \U$39508 ( \39885 , \39884 );
xor \U$39509 ( \39886 , RIae7a2b8_175, \10141 );
not \U$39510 ( \39887 , \39886 );
not \U$39511 ( \39888 , \9813 );
or \U$39512 ( \39889 , \39887 , \39888 );
not \U$39513 ( \39890 , \10031 );
not \U$39514 ( \39891 , \39890 );
not \U$39515 ( \39892 , RIae7a2b8_175);
and \U$39516 ( \39893 , \39891 , \39892 );
and \U$39517 ( \39894 , \16922 , RIae7a2b8_175);
nor \U$39518 ( \39895 , \39893 , \39894 );
or \U$39519 ( \39896 , \39895 , \38247 );
nand \U$39520 ( \39897 , \39889 , \39896 );
not \U$39521 ( \39898 , \39897 );
or \U$39522 ( \39899 , RIae79e80_166, RIae79ef8_167);
nand \U$39523 ( \39900 , \39899 , \12857 );
and \U$39524 ( \39901 , \39900 , \4969 );
not \U$39525 ( \39902 , \5048 );
not \U$39526 ( \39903 , \39821 );
or \U$39527 ( \39904 , \39902 , \39903 );
not \U$39528 ( \39905 , \4968 );
not \U$39529 ( \39906 , \12857 );
or \U$39530 ( \39907 , \39905 , \39906 );
or \U$39531 ( \39908 , \12857 , \6084 );
nand \U$39532 ( \39909 , \39907 , \39908 );
nand \U$39533 ( \39910 , \39909 , \5039 );
nand \U$39534 ( \39911 , \39904 , \39910 );
and \U$39535 ( \39912 , \39901 , \39911 );
not \U$39536 ( \39913 , \39912 );
not \U$39537 ( \39914 , \9516 );
not \U$39538 ( \39915 , \39651 );
or \U$39539 ( \39916 , \39914 , \39915 );
buf \U$39540 ( \39917 , \16035 );
and \U$39541 ( \39918 , RIae79fe8_169, \39917 );
not \U$39542 ( \39919 , RIae79fe8_169);
and \U$39543 ( \39920 , \39919 , \16036 );
nor \U$39544 ( \39921 , \39918 , \39920 );
nand \U$39545 ( \39922 , \39921 , \9499 );
nand \U$39546 ( \39923 , \39916 , \39922 );
not \U$39547 ( \39924 , \39923 );
not \U$39548 ( \39925 , \39924 );
or \U$39549 ( \39926 , \39913 , \39925 );
or \U$39550 ( \39927 , \39924 , \39912 );
nand \U$39551 ( \39928 , \39926 , \39927 );
not \U$39552 ( \39929 , \39928 );
or \U$39553 ( \39930 , \39898 , \39929 );
nand \U$39554 ( \39931 , \39923 , \39912 );
nand \U$39555 ( \39932 , \39930 , \39931 );
not \U$39556 ( \39933 , \10275 );
not \U$39557 ( \39934 , \39666 );
or \U$39558 ( \39935 , \39933 , \39934 );
xor \U$39559 ( \39936 , RIae7a8d0_188, \6345 );
nand \U$39560 ( \39937 , \39936 , \11204 );
nand \U$39561 ( \39938 , \39935 , \39937 );
xor \U$39562 ( \39939 , \39932 , \39938 );
not \U$39563 ( \39940 , \39939 );
or \U$39564 ( \39941 , \39885 , \39940 );
nand \U$39565 ( \39942 , \39938 , \39932 );
nand \U$39566 ( \39943 , \39941 , \39942 );
not \U$39567 ( \39944 , \39943 );
or \U$39568 ( \39945 , \39875 , \39944 );
or \U$39569 ( \39946 , \39943 , \39874 );
not \U$39570 ( \39947 , \9776 );
not \U$39571 ( \39948 , \39594 );
or \U$39572 ( \39949 , \39947 , \39948 );
xnor \U$39573 ( \39950 , \9412 , RIae7a150_172);
nand \U$39574 ( \39951 , \39950 , \9758 );
nand \U$39575 ( \39952 , \39949 , \39951 );
not \U$39576 ( \39953 , \39952 );
not \U$39577 ( \39954 , \11422 );
not \U$39578 ( \39955 , \39843 );
or \U$39579 ( \39956 , \39954 , \39955 );
xor \U$39580 ( \39957 , \16837 , RIae7a498_179);
nand \U$39581 ( \39958 , \39957 , \10695 );
nand \U$39582 ( \39959 , \39956 , \39958 );
not \U$39583 ( \39960 , \39959 );
not \U$39584 ( \39961 , \9478 );
not \U$39585 ( \39962 , \39616 );
or \U$39586 ( \39963 , \39961 , \39962 );
and \U$39587 ( \39964 , RIae7a6f0_184, \16274 );
not \U$39588 ( \39965 , RIae7a6f0_184);
and \U$39589 ( \39966 , \39965 , \16271 );
nor \U$39590 ( \39967 , \39964 , \39966 );
nand \U$39591 ( \39968 , \39967 , \9473 );
nand \U$39592 ( \39969 , \39963 , \39968 );
not \U$39593 ( \39970 , \39969 );
not \U$39594 ( \39971 , \39970 );
or \U$39595 ( \39972 , \39960 , \39971 );
or \U$39596 ( \39973 , \39970 , \39959 );
nand \U$39597 ( \39974 , \39972 , \39973 );
not \U$39598 ( \39975 , \39974 );
or \U$39599 ( \39976 , \39953 , \39975 );
nand \U$39600 ( \39977 , \39969 , \39959 );
nand \U$39601 ( \39978 , \39976 , \39977 );
nand \U$39602 ( \39979 , \39946 , \39978 );
nand \U$39603 ( \39980 , \39945 , \39979 );
nand \U$39604 ( \39981 , \39873 , \39980 );
nand \U$39605 ( \39982 , \39872 , \39981 );
not \U$39606 ( \39983 , \39982 );
not \U$39607 ( \39984 , \39704 );
not \U$39608 ( \39985 , \39760 );
and \U$39609 ( \39986 , \39984 , \39985 );
and \U$39610 ( \39987 , \39760 , \39704 );
nor \U$39611 ( \39988 , \39986 , \39987 );
not \U$39612 ( \39989 , \39988 );
xor \U$39613 ( \39990 , \39187 , \39222 );
xor \U$39614 ( \39991 , \39990 , \39225 );
not \U$39615 ( \39992 , \39991 );
or \U$39616 ( \39993 , \39989 , \39992 );
or \U$39617 ( \39994 , \39991 , \39988 );
nand \U$39618 ( \39995 , \39993 , \39994 );
not \U$39619 ( \39996 , \39995 );
or \U$39620 ( \39997 , \39983 , \39996 );
not \U$39621 ( \39998 , \39988 );
nand \U$39622 ( \39999 , \39998 , \39991 );
nand \U$39623 ( \40000 , \39997 , \39999 );
not \U$39624 ( \40001 , \40000 );
nor \U$39625 ( \40002 , \39777 , \40001 );
xor \U$39626 ( \40003 , \39058 , \39233 );
nand \U$39627 ( \40004 , \40003 , \39775 );
not \U$39628 ( \40005 , \40004 );
nor \U$39629 ( \40006 , \40002 , \40005 );
not \U$39630 ( \40007 , \40006 );
or \U$39631 ( \40008 , \39774 , \40007 );
not \U$39632 ( \40009 , \40004 );
not \U$39633 ( \40010 , \40002 );
not \U$39634 ( \40011 , \40010 );
or \U$39635 ( \40012 , \40009 , \40011 );
not \U$39636 ( \40013 , \39773 );
nand \U$39637 ( \40014 , \40012 , \40013 );
nand \U$39638 ( \40015 , \40008 , \40014 );
not \U$39639 ( \40016 , \40015 );
or \U$39640 ( \40017 , \39542 , \40016 );
or \U$39641 ( \40018 , \40015 , \39541 );
nand \U$39642 ( \40019 , \40017 , \40018 );
not \U$39643 ( \40020 , \40019 );
xor \U$39644 ( \40021 , \39546 , \39544 );
xnor \U$39645 ( \40022 , \40021 , \39549 );
not \U$39646 ( \40023 , \40022 );
and \U$39647 ( \40024 , \39870 , \39864 );
not \U$39648 ( \40025 , \39870 );
and \U$39649 ( \40026 , \40025 , \39865 );
nor \U$39650 ( \40027 , \40024 , \40026 );
not \U$39651 ( \40028 , \39980 );
and \U$39652 ( \40029 , \40027 , \40028 );
not \U$39653 ( \40030 , \40027 );
and \U$39654 ( \40031 , \40030 , \39980 );
nor \U$39655 ( \40032 , \40029 , \40031 );
not \U$39656 ( \40033 , \40032 );
or \U$39657 ( \40034 , \40023 , \40033 );
and \U$39658 ( \40035 , \39621 , \39619 );
xor \U$39659 ( \40036 , \40035 , \39598 );
not \U$39660 ( \40037 , \40036 );
not \U$39661 ( \40038 , \39837 );
not \U$39662 ( \40039 , \40038 );
not \U$39663 ( \40040 , \39860 );
or \U$39664 ( \40041 , \40039 , \40040 );
or \U$39665 ( \40042 , \39860 , \40038 );
nand \U$39666 ( \40043 , \40041 , \40042 );
not \U$39667 ( \40044 , \40043 );
xor \U$39668 ( \40045 , \39658 , \39668 );
xor \U$39669 ( \40046 , \40045 , \39678 );
not \U$39670 ( \40047 , \40046 );
not \U$39671 ( \40048 , \40047 );
or \U$39672 ( \40049 , \40044 , \40048 );
not \U$39673 ( \40050 , \40043 );
nand \U$39674 ( \40051 , \40050 , \40046 );
nand \U$39675 ( \40052 , \40049 , \40051 );
not \U$39676 ( \40053 , \40052 );
or \U$39677 ( \40054 , \40037 , \40053 );
not \U$39678 ( \40055 , \40047 );
nand \U$39679 ( \40056 , \40055 , \40043 );
nand \U$39680 ( \40057 , \40054 , \40056 );
nand \U$39681 ( \40058 , \40034 , \40057 );
not \U$39682 ( \40059 , \40032 );
not \U$39683 ( \40060 , \40022 );
nand \U$39684 ( \40061 , \40059 , \40060 );
nand \U$39685 ( \40062 , \40058 , \40061 );
not \U$39686 ( \40063 , RIae7aab0_192);
not \U$39687 ( \40064 , \39676 );
or \U$39688 ( \40065 , \40063 , \40064 );
not \U$39689 ( \40066 , \14671 );
not \U$39690 ( \40067 , \16311 );
or \U$39691 ( \40068 , \40066 , \40067 );
nand \U$39692 ( \40069 , \15128 , RIae7aa38_191);
nand \U$39693 ( \40070 , \40068 , \40069 );
nand \U$39694 ( \40071 , \40070 , \16383 );
nand \U$39695 ( \40072 , \40065 , \40071 );
not \U$39696 ( \40073 , \40072 );
xnor \U$39697 ( \40074 , \39653 , \39642 );
not \U$39698 ( \40075 , \40074 );
not \U$39699 ( \40076 , \10519 );
not \U$39700 ( \40077 , \39580 );
or \U$39701 ( \40078 , \40076 , \40077 );
and \U$39702 ( \40079 , RIae7a7e0_186, \29050 );
not \U$39703 ( \40080 , RIae7a7e0_186);
and \U$39704 ( \40081 , \40080 , \15091 );
or \U$39705 ( \40082 , \40079 , \40081 );
nand \U$39706 ( \40083 , \40082 , \11439 );
nand \U$39707 ( \40084 , \40078 , \40083 );
nand \U$39708 ( \40085 , \40075 , \40084 );
nand \U$39709 ( \40086 , \40073 , \40085 );
not \U$39710 ( \40087 , \40084 );
nand \U$39711 ( \40088 , \40087 , \40074 );
nand \U$39712 ( \40089 , \40086 , \40088 );
not \U$39713 ( \40090 , \40089 );
not \U$39714 ( \40091 , \9699 );
not \U$39715 ( \40092 , \39741 );
or \U$39716 ( \40093 , \40091 , \40092 );
and \U$39717 ( \40094 , RIae7a240_174, \10000 );
not \U$39718 ( \40095 , RIae7a240_174);
and \U$39719 ( \40096 , \40095 , \10007 );
or \U$39720 ( \40097 , \40094 , \40096 );
nand \U$39721 ( \40098 , \40097 , \9687 );
nand \U$39722 ( \40099 , \40093 , \40098 );
not \U$39723 ( \40100 , \9813 );
not \U$39724 ( \40101 , \39567 );
or \U$39725 ( \40102 , \40100 , \40101 );
nand \U$39726 ( \40103 , \39886 , \9792 );
nand \U$39727 ( \40104 , \40102 , \40103 );
nand \U$39728 ( \40105 , \40099 , \40104 );
not \U$39729 ( \40106 , \40105 );
not \U$39730 ( \40107 , \10631 );
not \U$39731 ( \40108 , \39558 );
or \U$39732 ( \40109 , \40107 , \40108 );
not \U$39733 ( \40110 , RIae7a510_180);
not \U$39734 ( \40111 , \11387 );
or \U$39735 ( \40112 , \40110 , \40111 );
or \U$39736 ( \40113 , \10084 , RIae7a510_180);
nand \U$39737 ( \40114 , \40112 , \40113 );
nand \U$39738 ( \40115 , \40114 , \11400 );
nand \U$39739 ( \40116 , \40109 , \40115 );
not \U$39740 ( \40117 , \40116 );
not \U$39741 ( \40118 , \40117 );
or \U$39742 ( \40119 , \40106 , \40118 );
not \U$39743 ( \40120 , \40099 );
not \U$39744 ( \40121 , \40104 );
nand \U$39745 ( \40122 , \40120 , \40121 );
nand \U$39746 ( \40123 , \40119 , \40122 );
not \U$39747 ( \40124 , \40123 );
not \U$39748 ( \40125 , \39584 );
not \U$39749 ( \40126 , \39587 );
nor \U$39750 ( \40127 , \40126 , \39572 );
not \U$39751 ( \40128 , \40127 );
and \U$39752 ( \40129 , \40125 , \40128 );
and \U$39753 ( \40130 , \39584 , \40127 );
nor \U$39754 ( \40131 , \40129 , \40130 );
not \U$39755 ( \40132 , \40131 );
or \U$39756 ( \40133 , \40124 , \40132 );
or \U$39757 ( \40134 , \40131 , \40123 );
nand \U$39758 ( \40135 , \40133 , \40134 );
not \U$39759 ( \40136 , \40135 );
or \U$39760 ( \40137 , \40090 , \40136 );
not \U$39761 ( \40138 , \40131 );
nand \U$39762 ( \40139 , \40138 , \40123 );
nand \U$39763 ( \40140 , \40137 , \40139 );
xor \U$39764 ( \40141 , \39708 , \39718 );
xor \U$39765 ( \40142 , \40141 , \39754 );
not \U$39766 ( \40143 , \40142 );
nand \U$39767 ( \40144 , \40140 , \40143 );
not \U$39768 ( \40145 , \40144 );
not \U$39769 ( \40146 , \40140 );
not \U$39770 ( \40147 , \40143 );
and \U$39771 ( \40148 , \40146 , \40147 );
not \U$39772 ( \40149 , \39623 );
nand \U$39773 ( \40150 , \40149 , \39683 );
not \U$39774 ( \40151 , \40150 );
not \U$39775 ( \40152 , \39681 );
and \U$39776 ( \40153 , \40151 , \40152 );
and \U$39777 ( \40154 , \40150 , \39681 );
nor \U$39778 ( \40155 , \40153 , \40154 );
nor \U$39779 ( \40156 , \40148 , \40155 );
nor \U$39780 ( \40157 , \40145 , \40156 );
xor \U$39781 ( \40158 , \40062 , \40157 );
xor \U$39782 ( \40159 , \39552 , \39688 );
and \U$39783 ( \40160 , \40158 , \40159 );
and \U$39784 ( \40161 , \40062 , \40157 );
or \U$39785 ( \40162 , \40160 , \40161 );
xor \U$39786 ( \40163 , \39768 , \39693 );
xor \U$39787 ( \40164 , \40162 , \40163 );
not \U$39788 ( \40165 , \40164 );
not \U$39789 ( \40166 , \39777 );
not \U$39790 ( \40167 , \40000 );
and \U$39791 ( \40168 , \40166 , \40167 );
and \U$39792 ( \40169 , \39777 , \40000 );
nor \U$39793 ( \40170 , \40168 , \40169 );
not \U$39794 ( \40171 , \40170 );
not \U$39795 ( \40172 , \40171 );
or \U$39796 ( \40173 , \40165 , \40172 );
nand \U$39797 ( \40174 , \40162 , \40163 );
nand \U$39798 ( \40175 , \40173 , \40174 );
not \U$39799 ( \40176 , \40175 );
nand \U$39800 ( \40177 , \40020 , \40176 );
not \U$39801 ( \40178 , \39541 );
not \U$39802 ( \40179 , \40178 );
not \U$39803 ( \40180 , \40015 );
or \U$39804 ( \40181 , \40179 , \40180 );
not \U$39805 ( \40182 , \40004 );
not \U$39806 ( \40183 , \40010 );
or \U$39807 ( \40184 , \40182 , \40183 );
nand \U$39808 ( \40185 , \40184 , \39773 );
nand \U$39809 ( \40186 , \40181 , \40185 );
not \U$39810 ( \40187 , \40186 );
xnor \U$39811 ( \40188 , \39425 , \39337 );
nand \U$39812 ( \40189 , \40187 , \40188 );
nand \U$39813 ( \40190 , \40177 , \40189 );
nand \U$39814 ( \40191 , \40019 , \40175 );
not \U$39815 ( \40192 , \11434 );
not \U$39816 ( \40193 , RIae7a498_179);
buf \U$39817 ( \40194 , \16829 );
not \U$39818 ( \40195 , \40194 );
not \U$39819 ( \40196 , \40195 );
or \U$39820 ( \40197 , \40193 , \40196 );
buf \U$39821 ( \40198 , \13657 );
or \U$39822 ( \40199 , \40198 , RIae7a498_179);
nand \U$39823 ( \40200 , \40197 , \40199 );
not \U$39824 ( \40201 , \40200 );
or \U$39825 ( \40202 , \40192 , \40201 );
nand \U$39826 ( \40203 , \39957 , \10676 );
nand \U$39827 ( \40204 , \40202 , \40203 );
not \U$39828 ( \40205 , \40204 );
xor \U$39829 ( \40206 , \39827 , \39810 );
not \U$39830 ( \40207 , \11013 );
and \U$39831 ( \40208 , RIae7a3a8_177, \9868 );
not \U$39832 ( \40209 , RIae7a3a8_177);
and \U$39833 ( \40210 , \40209 , \13896 );
nor \U$39834 ( \40211 , \40208 , \40210 );
not \U$39835 ( \40212 , \40211 );
or \U$39836 ( \40213 , \40207 , \40212 );
nand \U$39837 ( \40214 , \39785 , \9622 );
nand \U$39838 ( \40215 , \40213 , \40214 );
xor \U$39839 ( \40216 , \40206 , \40215 );
not \U$39840 ( \40217 , \40216 );
or \U$39841 ( \40218 , \40205 , \40217 );
nand \U$39842 ( \40219 , \40215 , \40206 );
nand \U$39843 ( \40220 , \40218 , \40219 );
not \U$39844 ( \40221 , \40220 );
xnor \U$39845 ( \40222 , \39787 , \39833 );
nand \U$39846 ( \40223 , \40221 , \40222 );
not \U$39847 ( \40224 , \40223 );
not \U$39848 ( \40225 , \9730 );
not \U$39849 ( \40226 , RIae7a060_170);
not \U$39850 ( \40227 , \10937 );
or \U$39851 ( \40228 , \40226 , \40227 );
or \U$39852 ( \40229 , \12603 , RIae7a060_170);
nand \U$39853 ( \40230 , \40228 , \40229 );
not \U$39854 ( \40231 , \40230 );
or \U$39855 ( \40232 , \40225 , \40231 );
nand \U$39856 ( \40233 , \39882 , \10542 );
nand \U$39857 ( \40234 , \40232 , \40233 );
not \U$39858 ( \40235 , \40234 );
not \U$39859 ( \40236 , \11205 );
not \U$39860 ( \40237 , RIae7a8d0_188);
not \U$39861 ( \40238 , \22353 );
or \U$39862 ( \40239 , \40237 , \40238 );
or \U$39863 ( \40240 , \12684 , RIae7a8d0_188);
nand \U$39864 ( \40241 , \40239 , \40240 );
not \U$39865 ( \40242 , \40241 );
or \U$39866 ( \40243 , \40236 , \40242 );
nand \U$39867 ( \40244 , \39936 , \10275 );
nand \U$39868 ( \40245 , \40243 , \40244 );
xor \U$39869 ( \40246 , \39901 , \39911 );
not \U$39870 ( \40247 , \39808 );
or \U$39871 ( \40248 , \40247 , \6193 );
not \U$39872 ( \40249 , \6207 );
not \U$39873 ( \40250 , \36790 );
or \U$39874 ( \40251 , \40249 , \40250 );
nand \U$39875 ( \40252 , \10844 , RIae79ef8_167);
nand \U$39876 ( \40253 , \40251 , \40252 );
not \U$39877 ( \40254 , \40253 );
or \U$39878 ( \40255 , \40254 , \6198 );
nand \U$39879 ( \40256 , \40248 , \40255 );
xor \U$39880 ( \40257 , \40246 , \40256 );
not \U$39881 ( \40258 , \39921 );
not \U$39882 ( \40259 , \9517 );
or \U$39883 ( \40260 , \40258 , \40259 );
xor \U$39884 ( \40261 , RIae79fe8_169, \11321 );
not \U$39885 ( \40262 , \40261 );
not \U$39886 ( \40263 , \9499 );
or \U$39887 ( \40264 , \40262 , \40263 );
nand \U$39888 ( \40265 , \40260 , \40264 );
and \U$39889 ( \40266 , \40257 , \40265 );
and \U$39890 ( \40267 , \40246 , \40256 );
nor \U$39891 ( \40268 , \40266 , \40267 );
and \U$39892 ( \40269 , \40245 , \40268 );
not \U$39893 ( \40270 , \40245 );
not \U$39894 ( \40271 , \40268 );
and \U$39895 ( \40272 , \40270 , \40271 );
or \U$39896 ( \40273 , \40269 , \40272 );
not \U$39897 ( \40274 , \40273 );
or \U$39898 ( \40275 , \40235 , \40274 );
nand \U$39899 ( \40276 , \40245 , \40271 );
nand \U$39900 ( \40277 , \40275 , \40276 );
not \U$39901 ( \40278 , \40277 );
or \U$39902 ( \40279 , \40224 , \40278 );
not \U$39903 ( \40280 , \40222 );
nand \U$39904 ( \40281 , \40280 , \40220 );
nand \U$39905 ( \40282 , \40279 , \40281 );
and \U$39906 ( \40283 , \39943 , \39874 );
not \U$39907 ( \40284 , \39943 );
not \U$39908 ( \40285 , \39874 );
and \U$39909 ( \40286 , \40284 , \40285 );
nor \U$39910 ( \40287 , \40283 , \40286 );
xor \U$39911 ( \40288 , \40287 , \39978 );
xor \U$39912 ( \40289 , \40282 , \40288 );
not \U$39913 ( \40290 , \40116 );
not \U$39914 ( \40291 , \40099 );
not \U$39915 ( \40292 , \40121 );
and \U$39916 ( \40293 , \40291 , \40292 );
and \U$39917 ( \40294 , \40099 , \40121 );
nor \U$39918 ( \40295 , \40293 , \40294 );
not \U$39919 ( \40296 , \40295 );
or \U$39920 ( \40297 , \40290 , \40296 );
or \U$39921 ( \40298 , \40295 , \40116 );
nand \U$39922 ( \40299 , \40297 , \40298 );
not \U$39923 ( \40300 , \40299 );
not \U$39924 ( \40301 , \11400 );
xor \U$39925 ( \40302 , RIae7a510_180, \10066 );
not \U$39926 ( \40303 , \40302 );
or \U$39927 ( \40304 , \40301 , \40303 );
nand \U$39928 ( \40305 , \40114 , \10631 );
nand \U$39929 ( \40306 , \40304 , \40305 );
not \U$39930 ( \40307 , \9687 );
not \U$39931 ( \40308 , RIae7a240_174);
not \U$39932 ( \40309 , \10740 );
or \U$39933 ( \40310 , \40308 , \40309 );
or \U$39934 ( \40311 , \19035 , RIae7a240_174);
nand \U$39935 ( \40312 , \40310 , \40311 );
not \U$39936 ( \40313 , \40312 );
or \U$39937 ( \40314 , \40307 , \40313 );
nand \U$39938 ( \40315 , \40097 , \9699 );
nand \U$39939 ( \40316 , \40314 , \40315 );
xnor \U$39940 ( \40317 , \40306 , \40316 );
not \U$39941 ( \40318 , \40317 );
not \U$39942 ( \40319 , \40318 );
not \U$39943 ( \40320 , \11439 );
not \U$39944 ( \40321 , \9529 );
not \U$39945 ( \40322 , \12614 );
or \U$39946 ( \40323 , \40321 , \40322 );
not \U$39947 ( \40324 , \9442 );
or \U$39948 ( \40325 , \40324 , \17112 );
nand \U$39949 ( \40326 , \40323 , \40325 );
not \U$39950 ( \40327 , \40326 );
or \U$39951 ( \40328 , \40320 , \40327 );
nand \U$39952 ( \40329 , \40082 , \10519 );
nand \U$39953 ( \40330 , \40328 , \40329 );
not \U$39954 ( \40331 , \40330 );
or \U$39955 ( \40332 , \40319 , \40331 );
nand \U$39956 ( \40333 , \40306 , \40316 );
nand \U$39957 ( \40334 , \40332 , \40333 );
not \U$39958 ( \40335 , \40334 );
or \U$39959 ( \40336 , \40300 , \40335 );
not \U$39960 ( \40337 , \9777 );
not \U$39961 ( \40338 , \39950 );
or \U$39962 ( \40339 , \40337 , \40338 );
and \U$39963 ( \40340 , RIae7a150_172, \9607 );
not \U$39964 ( \40341 , RIae7a150_172);
and \U$39965 ( \40342 , \40341 , \29247 );
nor \U$39966 ( \40343 , \40340 , \40342 );
nand \U$39967 ( \40344 , \40343 , \10667 );
nand \U$39968 ( \40345 , \40339 , \40344 );
not \U$39969 ( \40346 , \40345 );
not \U$39970 ( \40347 , \9473 );
and \U$39971 ( \40348 , \17387 , \16101 );
not \U$39972 ( \40349 , \17387 );
and \U$39973 ( \40350 , \40349 , RIae7a6f0_184);
nor \U$39974 ( \40351 , \40348 , \40350 );
not \U$39975 ( \40352 , \40351 );
or \U$39976 ( \40353 , \40347 , \40352 );
nand \U$39977 ( \40354 , \39967 , \9478 );
nand \U$39978 ( \40355 , \40353 , \40354 );
not \U$39979 ( \40356 , \40355 );
or \U$39980 ( \40357 , \40346 , \40356 );
or \U$39981 ( \40358 , \40355 , \40345 );
not \U$39982 ( \40359 , RIae7aab0_192);
not \U$39983 ( \40360 , \40070 );
or \U$39984 ( \40361 , \40359 , \40360 );
and \U$39985 ( \40362 , RIae7aa38_191, \13976 );
not \U$39986 ( \40363 , RIae7aa38_191);
and \U$39987 ( \40364 , \40363 , \21732 );
or \U$39988 ( \40365 , \40362 , \40364 );
nand \U$39989 ( \40366 , \40365 , \14668 );
nand \U$39990 ( \40367 , \40361 , \40366 );
nand \U$39991 ( \40368 , \40358 , \40367 );
nand \U$39992 ( \40369 , \40357 , \40368 );
not \U$39993 ( \40370 , \40299 );
not \U$39994 ( \40371 , \40334 );
nand \U$39995 ( \40372 , \40370 , \40371 );
nand \U$39996 ( \40373 , \40369 , \40372 );
nand \U$39997 ( \40374 , \40336 , \40373 );
and \U$39998 ( \40375 , \40289 , \40374 );
and \U$39999 ( \40376 , \40282 , \40288 );
or \U$40000 ( \40377 , \40375 , \40376 );
not \U$40001 ( \40378 , \40052 );
not \U$40002 ( \40379 , \40036 );
not \U$40003 ( \40380 , \40379 );
and \U$40004 ( \40381 , \40378 , \40380 );
and \U$40005 ( \40382 , \40052 , \40379 );
nor \U$40006 ( \40383 , \40381 , \40382 );
not \U$40007 ( \40384 , \40383 );
not \U$40008 ( \40385 , \40384 );
not \U$40009 ( \40386 , \40089 );
not \U$40010 ( \40387 , \40135 );
not \U$40011 ( \40388 , \40387 );
or \U$40012 ( \40389 , \40386 , \40388 );
not \U$40013 ( \40390 , \40089 );
nand \U$40014 ( \40391 , \40390 , \40135 );
nand \U$40015 ( \40392 , \40389 , \40391 );
not \U$40016 ( \40393 , \40392 );
not \U$40017 ( \40394 , \40393 );
or \U$40018 ( \40395 , \40385 , \40394 );
not \U$40019 ( \40396 , \40392 );
not \U$40020 ( \40397 , \40383 );
or \U$40021 ( \40398 , \40396 , \40397 );
xor \U$40022 ( \40399 , \40074 , \40084 );
xnor \U$40023 ( \40400 , \40399 , \40072 );
not \U$40024 ( \40401 , \40400 );
and \U$40025 ( \40402 , \39939 , \39884 );
not \U$40026 ( \40403 , \39939 );
not \U$40027 ( \40404 , \39884 );
and \U$40028 ( \40405 , \40403 , \40404 );
nor \U$40029 ( \40406 , \40402 , \40405 );
xor \U$40030 ( \40407 , \39974 , \39952 );
and \U$40031 ( \40408 , \40406 , \40407 );
not \U$40032 ( \40409 , \40408 );
and \U$40033 ( \40410 , \40401 , \40409 );
nor \U$40034 ( \40411 , \40407 , \40406 );
nor \U$40035 ( \40412 , \40410 , \40411 );
nand \U$40036 ( \40413 , \40398 , \40412 );
nand \U$40037 ( \40414 , \40395 , \40413 );
xor \U$40038 ( \40415 , \40377 , \40414 );
xor \U$40039 ( \40416 , \40142 , \40155 );
xnor \U$40040 ( \40417 , \40416 , \40140 );
and \U$40041 ( \40418 , \40415 , \40417 );
and \U$40042 ( \40419 , \40377 , \40414 );
or \U$40043 ( \40420 , \40418 , \40419 );
xor \U$40044 ( \40421 , \39995 , \39982 );
or \U$40045 ( \40422 , \40420 , \40421 );
xor \U$40046 ( \40423 , \40062 , \40157 );
xor \U$40047 ( \40424 , \40423 , \40159 );
and \U$40048 ( \40425 , \40422 , \40424 );
and \U$40049 ( \40426 , \40421 , \40420 );
nor \U$40050 ( \40427 , \40425 , \40426 );
not \U$40051 ( \40428 , \40427 );
not \U$40052 ( \40429 , \40170 );
not \U$40053 ( \40430 , \40164 );
or \U$40054 ( \40431 , \40429 , \40430 );
or \U$40055 ( \40432 , \40164 , \40170 );
nand \U$40056 ( \40433 , \40431 , \40432 );
nand \U$40057 ( \40434 , \40428 , \40433 );
not \U$40058 ( \40435 , \40434 );
not \U$40059 ( \40436 , \40369 );
and \U$40060 ( \40437 , \40299 , \40371 );
not \U$40061 ( \40438 , \40299 );
and \U$40062 ( \40439 , \40438 , \40334 );
or \U$40063 ( \40440 , \40437 , \40439 );
not \U$40064 ( \40441 , \40440 );
or \U$40065 ( \40442 , \40436 , \40441 );
or \U$40066 ( \40443 , \40440 , \40369 );
nand \U$40067 ( \40444 , \40442 , \40443 );
not \U$40068 ( \40445 , \40444 );
xor \U$40069 ( \40446 , \40273 , \40234 );
not \U$40070 ( \40447 , \40446 );
not \U$40071 ( \40448 , \40447 );
xor \U$40072 ( \40449 , \40216 , \40204 );
not \U$40073 ( \40450 , \40449 );
not \U$40074 ( \40451 , \40450 );
or \U$40075 ( \40452 , \40448 , \40451 );
not \U$40076 ( \40453 , \40449 );
not \U$40077 ( \40454 , \40446 );
or \U$40078 ( \40455 , \40453 , \40454 );
xor \U$40079 ( \40456 , \40345 , \40367 );
xnor \U$40080 ( \40457 , \40456 , \40355 );
nand \U$40081 ( \40458 , \40455 , \40457 );
nand \U$40082 ( \40459 , \40452 , \40458 );
not \U$40083 ( \40460 , \40459 );
or \U$40084 ( \40461 , \40445 , \40460 );
xor \U$40085 ( \40462 , \40406 , \40407 );
xor \U$40086 ( \40463 , \40400 , \40462 );
nand \U$40087 ( \40464 , \40461 , \40463 );
not \U$40088 ( \40465 , \40444 );
not \U$40089 ( \40466 , \40459 );
nand \U$40090 ( \40467 , \40465 , \40466 );
nand \U$40091 ( \40468 , \40464 , \40467 );
xor \U$40092 ( \40469 , \40282 , \40288 );
xor \U$40093 ( \40470 , \40469 , \40374 );
xor \U$40094 ( \40471 , \40468 , \40470 );
not \U$40095 ( \40472 , \10275 );
not \U$40096 ( \40473 , \40241 );
or \U$40097 ( \40474 , \40472 , \40473 );
xor \U$40098 ( \40475 , RIae7a8d0_188, \15102 );
nand \U$40099 ( \40476 , \40475 , \11205 );
nand \U$40100 ( \40477 , \40474 , \40476 );
not \U$40101 ( \40478 , \40477 );
not \U$40102 ( \40479 , \9687 );
not \U$40103 ( \40480 , \19623 );
not \U$40104 ( \40481 , \33415 );
or \U$40105 ( \40482 , \40480 , \40481 );
nand \U$40106 ( \40483 , \16922 , RIae7a240_174);
nand \U$40107 ( \40484 , \40482 , \40483 );
not \U$40108 ( \40485 , \40484 );
or \U$40109 ( \40486 , \40479 , \40485 );
not \U$40110 ( \40487 , RIae7a240_174);
not \U$40111 ( \40488 , \10149 );
or \U$40112 ( \40489 , \40487 , \40488 );
buf \U$40113 ( \40490 , \10149 );
or \U$40114 ( \40491 , \40490 , RIae7a240_174);
nand \U$40115 ( \40492 , \40489 , \40491 );
nand \U$40116 ( \40493 , \40492 , \9699 );
nand \U$40117 ( \40494 , \40486 , \40493 );
not \U$40118 ( \40495 , \40494 );
not \U$40119 ( \40496 , \5870 );
or \U$40120 ( \40497 , RIae79f70_168, RIae79fe8_169);
nand \U$40121 ( \40498 , \40497 , \12857 );
nand \U$40122 ( \40499 , \40496 , \40498 );
not \U$40123 ( \40500 , \40499 );
not \U$40124 ( \40501 , \6212 );
and \U$40125 ( \40502 , RIae79ef8_167, \18989 );
not \U$40126 ( \40503 , RIae79ef8_167);
and \U$40127 ( \40504 , \40503 , \37057 );
nor \U$40128 ( \40505 , \40502 , \40504 );
not \U$40129 ( \40506 , \40505 );
or \U$40130 ( \40507 , \40501 , \40506 );
not \U$40131 ( \40508 , \6203 );
not \U$40132 ( \40509 , \12857 );
or \U$40133 ( \40510 , \40508 , \40509 );
or \U$40134 ( \40511 , \12858 , \28303 );
nand \U$40135 ( \40512 , \40510 , \40511 );
nand \U$40136 ( \40513 , \40512 , \6199 );
nand \U$40137 ( \40514 , \40507 , \40513 );
nand \U$40138 ( \40515 , \40500 , \40514 );
not \U$40139 ( \40516 , \40515 );
not \U$40140 ( \40517 , \9813 );
not \U$40141 ( \40518 , \11054 );
not \U$40142 ( \40519 , \16912 );
or \U$40143 ( \40520 , \40518 , \40519 );
or \U$40144 ( \40521 , \11665 , \9799 );
nand \U$40145 ( \40522 , \40520 , \40521 );
not \U$40146 ( \40523 , \40522 );
or \U$40147 ( \40524 , \40517 , \40523 );
and \U$40148 ( \40525 , \39917 , RIae7a2b8_175);
not \U$40149 ( \40526 , \39917 );
and \U$40150 ( \40527 , \40526 , \28198 );
nor \U$40151 ( \40528 , \40525 , \40527 );
nand \U$40152 ( \40529 , \40528 , \9791 );
nand \U$40153 ( \40530 , \40524 , \40529 );
not \U$40154 ( \40531 , \40530 );
or \U$40155 ( \40532 , \40516 , \40531 );
or \U$40156 ( \40533 , \40530 , \40515 );
nand \U$40157 ( \40534 , \40532 , \40533 );
not \U$40158 ( \40535 , \40534 );
or \U$40159 ( \40536 , \40495 , \40535 );
not \U$40160 ( \40537 , \40515 );
nand \U$40161 ( \40538 , \40537 , \40530 );
nand \U$40162 ( \40539 , \40536 , \40538 );
not \U$40163 ( \40540 , \29519 );
not \U$40164 ( \40541 , \40326 );
or \U$40165 ( \40542 , \40540 , \40541 );
not \U$40166 ( \40543 , \9529 );
not \U$40167 ( \40544 , \9459 );
or \U$40168 ( \40545 , \40543 , \40544 );
nand \U$40169 ( \40546 , \9456 , RIae7a7e0_186);
nand \U$40170 ( \40547 , \40545 , \40546 );
nand \U$40171 ( \40548 , \40547 , \9549 );
nand \U$40172 ( \40549 , \40542 , \40548 );
xor \U$40173 ( \40550 , \40539 , \40549 );
not \U$40174 ( \40551 , \40550 );
or \U$40175 ( \40552 , \40478 , \40551 );
nand \U$40176 ( \40553 , \40549 , \40539 );
nand \U$40177 ( \40554 , \40552 , \40553 );
not \U$40178 ( \40555 , \40554 );
not \U$40179 ( \40556 , \9744 );
not \U$40180 ( \40557 , \40230 );
or \U$40181 ( \40558 , \40556 , \40557 );
not \U$40182 ( \40559 , RIae7a060_170);
not \U$40183 ( \40560 , \9412 );
or \U$40184 ( \40561 , \40559 , \40560 );
or \U$40185 ( \40562 , \9412 , RIae7a060_170);
nand \U$40186 ( \40563 , \40561 , \40562 );
nand \U$40187 ( \40564 , \40563 , \9729 );
nand \U$40188 ( \40565 , \40558 , \40564 );
not \U$40189 ( \40566 , \9776 );
not \U$40190 ( \40567 , \40343 );
or \U$40191 ( \40568 , \40566 , \40567 );
and \U$40192 ( \40569 , RIae7a150_172, \15501 );
not \U$40193 ( \40570 , RIae7a150_172);
and \U$40194 ( \40571 , \40570 , \15504 );
or \U$40195 ( \40572 , \40569 , \40571 );
nand \U$40196 ( \40573 , \40572 , \9758 );
nand \U$40197 ( \40574 , \40568 , \40573 );
or \U$40198 ( \40575 , \40565 , \40574 );
not \U$40199 ( \40576 , \14668 );
and \U$40200 ( \40577 , RIae7aa38_191, \9291 );
not \U$40201 ( \40578 , RIae7aa38_191);
and \U$40202 ( \40579 , \40578 , \6345 );
or \U$40203 ( \40580 , \40577 , \40579 );
not \U$40204 ( \40581 , \40580 );
or \U$40205 ( \40582 , \40576 , \40581 );
nand \U$40206 ( \40583 , \40365 , RIae7aab0_192);
nand \U$40207 ( \40584 , \40582 , \40583 );
nand \U$40208 ( \40585 , \40575 , \40584 );
nand \U$40209 ( \40586 , \40565 , \40574 );
nand \U$40210 ( \40587 , \40585 , \40586 );
not \U$40211 ( \40588 , \40587 );
not \U$40212 ( \40589 , \40588 );
and \U$40213 ( \40590 , \40330 , \40317 );
not \U$40214 ( \40591 , \40330 );
and \U$40215 ( \40592 , \40591 , \40318 );
or \U$40216 ( \40593 , \40590 , \40592 );
not \U$40217 ( \40594 , \40593 );
or \U$40218 ( \40595 , \40589 , \40594 );
or \U$40219 ( \40596 , \40593 , \40588 );
nand \U$40220 ( \40597 , \40595 , \40596 );
not \U$40221 ( \40598 , \40597 );
or \U$40222 ( \40599 , \40555 , \40598 );
nand \U$40223 ( \40600 , \40593 , \40587 );
nand \U$40224 ( \40601 , \40599 , \40600 );
not \U$40225 ( \40602 , \40601 );
not \U$40226 ( \40603 , \9621 );
not \U$40227 ( \40604 , \40211 );
or \U$40228 ( \40605 , \40603 , \40604 );
and \U$40229 ( \40606 , \10000 , \11690 );
not \U$40230 ( \40607 , \10000 );
and \U$40231 ( \40608 , \40607 , RIae7a3a8_177);
nor \U$40232 ( \40609 , \40606 , \40608 );
nand \U$40233 ( \40610 , \40609 , \9643 );
nand \U$40234 ( \40611 , \40605 , \40610 );
not \U$40235 ( \40612 , \40611 );
not \U$40236 ( \40613 , \9699 );
not \U$40237 ( \40614 , \40312 );
or \U$40238 ( \40615 , \40613 , \40614 );
nand \U$40239 ( \40616 , \40492 , \9687 );
nand \U$40240 ( \40617 , \40615 , \40616 );
not \U$40241 ( \40618 , \10631 );
not \U$40242 ( \40619 , \40302 );
or \U$40243 ( \40620 , \40618 , \40619 );
not \U$40244 ( \40621 , \36204 );
and \U$40245 ( \40622 , \10633 , \40621 );
not \U$40246 ( \40623 , \10633 );
and \U$40247 ( \40624 , \40623 , \11272 );
nor \U$40248 ( \40625 , \40622 , \40624 );
nand \U$40249 ( \40626 , \40625 , \11400 );
nand \U$40250 ( \40627 , \40620 , \40626 );
xor \U$40251 ( \40628 , \40617 , \40627 );
not \U$40252 ( \40629 , \40628 );
or \U$40253 ( \40630 , \40612 , \40629 );
nand \U$40254 ( \40631 , \40627 , \40617 );
nand \U$40255 ( \40632 , \40630 , \40631 );
not \U$40256 ( \40633 , \40632 );
xnor \U$40257 ( \40634 , \39897 , \39928 );
not \U$40258 ( \40635 , \40634 );
and \U$40259 ( \40636 , \12857 , \5048 );
not \U$40260 ( \40637 , \6212 );
not \U$40261 ( \40638 , \40253 );
or \U$40262 ( \40639 , \40637 , \40638 );
nand \U$40263 ( \40640 , \40505 , \6199 );
nand \U$40264 ( \40641 , \40639 , \40640 );
xor \U$40265 ( \40642 , \40636 , \40641 );
not \U$40266 ( \40643 , \9516 );
not \U$40267 ( \40644 , \40261 );
or \U$40268 ( \40645 , \40643 , \40644 );
and \U$40269 ( \40646 , RIae79fe8_169, \39806 );
not \U$40270 ( \40647 , RIae79fe8_169);
and \U$40271 ( \40648 , \40647 , \28267 );
or \U$40272 ( \40649 , \40646 , \40648 );
nand \U$40273 ( \40650 , \40649 , \9499 );
nand \U$40274 ( \40651 , \40645 , \40650 );
and \U$40275 ( \40652 , \40642 , \40651 );
and \U$40276 ( \40653 , \40636 , \40641 );
nor \U$40277 ( \40654 , \40652 , \40653 );
not \U$40278 ( \40655 , \40654 );
not \U$40279 ( \40656 , \9792 );
not \U$40280 ( \40657 , \40522 );
or \U$40281 ( \40658 , \40656 , \40657 );
not \U$40282 ( \40659 , \39895 );
nand \U$40283 ( \40660 , \40659 , \9813 );
nand \U$40284 ( \40661 , \40658 , \40660 );
not \U$40285 ( \40662 , \40661 );
or \U$40286 ( \40663 , \40655 , \40662 );
or \U$40287 ( \40664 , \40661 , \40654 );
nand \U$40288 ( \40665 , \40663 , \40664 );
not \U$40289 ( \40666 , \40665 );
not \U$40290 ( \40667 , \11422 );
not \U$40291 ( \40668 , \40200 );
or \U$40292 ( \40669 , \40667 , \40668 );
not \U$40293 ( \40670 , \10625 );
not \U$40294 ( \40671 , \38816 );
or \U$40295 ( \40672 , \40670 , \40671 );
nand \U$40296 ( \40673 , \10084 , RIae7a498_179);
nand \U$40297 ( \40674 , \40672 , \40673 );
nand \U$40298 ( \40675 , \40674 , \10695 );
nand \U$40299 ( \40676 , \40669 , \40675 );
not \U$40300 ( \40677 , \40676 );
or \U$40301 ( \40678 , \40666 , \40677 );
not \U$40302 ( \40679 , \40654 );
nand \U$40303 ( \40680 , \40679 , \40661 );
nand \U$40304 ( \40681 , \40678 , \40680 );
not \U$40305 ( \40682 , \40681 );
or \U$40306 ( \40683 , \40635 , \40682 );
or \U$40307 ( \40684 , \40681 , \40634 );
nand \U$40308 ( \40685 , \40683 , \40684 );
not \U$40309 ( \40686 , \40685 );
or \U$40310 ( \40687 , \40633 , \40686 );
not \U$40311 ( \40688 , \40634 );
nand \U$40312 ( \40689 , \40688 , \40681 );
nand \U$40313 ( \40690 , \40687 , \40689 );
not \U$40314 ( \40691 , \40690 );
or \U$40315 ( \40692 , \40602 , \40691 );
not \U$40316 ( \40693 , \40601 );
not \U$40317 ( \40694 , \40690 );
not \U$40318 ( \40695 , \40694 );
and \U$40319 ( \40696 , \40693 , \40695 );
and \U$40320 ( \40697 , \40601 , \40694 );
nor \U$40321 ( \40698 , \40696 , \40697 );
xor \U$40322 ( \40699 , \40220 , \40222 );
xor \U$40323 ( \40700 , \40699 , \40277 );
or \U$40324 ( \40701 , \40698 , \40700 );
nand \U$40325 ( \40702 , \40692 , \40701 );
and \U$40326 ( \40703 , \40471 , \40702 );
and \U$40327 ( \40704 , \40468 , \40470 );
or \U$40328 ( \40705 , \40703 , \40704 );
xor \U$40329 ( \40706 , \40057 , \40060 );
xor \U$40330 ( \40707 , \40706 , \40059 );
or \U$40331 ( \40708 , \40705 , \40707 );
xor \U$40332 ( \40709 , \40377 , \40414 );
xor \U$40333 ( \40710 , \40709 , \40417 );
and \U$40334 ( \40711 , \40708 , \40710 );
and \U$40335 ( \40712 , \40707 , \40705 );
nor \U$40336 ( \40713 , \40711 , \40712 );
not \U$40337 ( \40714 , \40713 );
xor \U$40338 ( \40715 , \40421 , \40420 );
and \U$40339 ( \40716 , \40715 , \40424 );
not \U$40340 ( \40717 , \40715 );
not \U$40341 ( \40718 , \40424 );
and \U$40342 ( \40719 , \40717 , \40718 );
nor \U$40343 ( \40720 , \40716 , \40719 );
nand \U$40344 ( \40721 , \40714 , \40720 );
not \U$40345 ( \40722 , \40721 );
or \U$40346 ( \40723 , \40435 , \40722 );
not \U$40347 ( \40724 , \40433 );
buf \U$40348 ( \40725 , \40427 );
nand \U$40349 ( \40726 , \40724 , \40725 );
nand \U$40350 ( \40727 , \40723 , \40726 );
nand \U$40351 ( \40728 , \40191 , \40727 );
not \U$40352 ( \40729 , \40728 );
or \U$40353 ( \40730 , \40190 , \40729 );
not \U$40354 ( \40731 , \40188 );
nand \U$40355 ( \40732 , \40731 , \40186 );
nand \U$40356 ( \40733 , \40730 , \40732 );
not \U$40357 ( \40734 , \40733 );
or \U$40358 ( \40735 , \39534 , \40734 );
nand \U$40359 ( \40736 , \39473 , \39429 );
not \U$40360 ( \40737 , \40736 );
nand \U$40361 ( \40738 , \40737 , \39532 );
xor \U$40362 ( \40739 , \38119 , \38121 );
xor \U$40363 ( \40740 , \40739 , \38183 );
not \U$40364 ( \40741 , \40740 );
not \U$40365 ( \40742 , \39515 );
not \U$40366 ( \40743 , \39510 );
or \U$40367 ( \40744 , \40742 , \40743 );
nand \U$40368 ( \40745 , \39504 , \39501 );
nand \U$40369 ( \40746 , \40744 , \40745 );
not \U$40370 ( \40747 , \40746 );
not \U$40371 ( \40748 , \40747 );
or \U$40372 ( \40749 , \40741 , \40748 );
or \U$40373 ( \40750 , \40747 , \40740 );
nand \U$40374 ( \40751 , \40749 , \40750 );
not \U$40375 ( \40752 , \38337 );
not \U$40376 ( \40753 , \38208 );
or \U$40377 ( \40754 , \40752 , \40753 );
or \U$40378 ( \40755 , \38208 , \38337 );
nand \U$40379 ( \40756 , \40754 , \40755 );
not \U$40380 ( \40757 , \40756 );
not \U$40381 ( \40758 , \38631 );
or \U$40382 ( \40759 , \40757 , \40758 );
or \U$40383 ( \40760 , \38631 , \40756 );
nand \U$40384 ( \40761 , \40759 , \40760 );
nand \U$40385 ( \40762 , \40751 , \40761 );
xor \U$40386 ( \40763 , \38198 , \38635 );
xor \U$40387 ( \40764 , \40763 , \38641 );
not \U$40388 ( \40765 , \40740 );
nand \U$40389 ( \40766 , \40765 , \40747 );
nand \U$40390 ( \40767 , \40762 , \40764 , \40766 );
xor \U$40391 ( \40768 , \40740 , \40761 );
xor \U$40392 ( \40769 , \40768 , \40747 );
and \U$40393 ( \40770 , \39520 , \39499 );
buf \U$40394 ( \40771 , \39493 );
nor \U$40395 ( \40772 , \40770 , \40771 );
nand \U$40396 ( \40773 , \40769 , \40772 );
not \U$40397 ( \40774 , \39525 );
not \U$40398 ( \40775 , \39531 );
nand \U$40399 ( \40776 , \40774 , \40775 );
and \U$40400 ( \40777 , \40738 , \40767 , \40773 , \40776 );
nand \U$40401 ( \40778 , \40735 , \40777 );
not \U$40402 ( \40779 , \40764 );
nand \U$40403 ( \40780 , \40762 , \40766 );
nand \U$40404 ( \40781 , \40779 , \40780 );
not \U$40405 ( \40782 , \40769 );
not \U$40406 ( \40783 , \40772 );
nand \U$40407 ( \40784 , \40782 , \40783 );
nand \U$40408 ( \40785 , \40781 , \40784 );
not \U$40409 ( \40786 , \40785 );
nand \U$40410 ( \40787 , \40778 , \40786 );
not \U$40411 ( \40788 , \40777 );
not \U$40412 ( \40789 , \40767 );
nand \U$40413 ( \40790 , \40788 , \40789 );
nand \U$40414 ( \40791 , \40787 , \40790 );
not \U$40415 ( \40792 , \40791 );
or \U$40416 ( \40793 , \38649 , \40792 );
buf \U$40417 ( \40794 , \37753 );
not \U$40418 ( \40795 , \40794 );
not \U$40419 ( \40796 , \38194 );
nor \U$40420 ( \40797 , \38196 , \38645 );
not \U$40421 ( \40798 , \40797 );
or \U$40422 ( \40799 , \40796 , \40798 );
not \U$40423 ( \40800 , \37765 );
not \U$40424 ( \40801 , \38193 );
nand \U$40425 ( \40802 , \40800 , \40801 );
nand \U$40426 ( \40803 , \40799 , \40802 );
not \U$40427 ( \40804 , \40803 );
or \U$40428 ( \40805 , \40795 , \40804 );
nor \U$40429 ( \40806 , \37758 , \37762 );
nor \U$40430 ( \40807 , \37735 , \37752 );
nor \U$40431 ( \40808 , \40806 , \40807 );
nand \U$40432 ( \40809 , \40805 , \40808 );
buf \U$40433 ( \40810 , \37763 );
nand \U$40434 ( \40811 , \40809 , \40810 );
nand \U$40435 ( \40812 , \40793 , \40811 );
not \U$40436 ( \40813 , \40812 );
or \U$40437 ( \40814 , \37029 , \40813 );
nand \U$40438 ( \40815 , \36305 , \36314 , \36625 );
nor \U$40439 ( \40816 , \36624 , \36321 );
nor \U$40440 ( \40817 , \36630 , \37025 );
nor \U$40441 ( \40818 , \40816 , \40817 );
or \U$40442 ( \40819 , \40815 , \40818 );
not \U$40443 ( \40820 , \36304 );
nand \U$40444 ( \40821 , \40820 , \36263 );
not \U$40445 ( \40822 , \36314 );
or \U$40446 ( \40823 , \40821 , \40822 );
or \U$40447 ( \40824 , \36311 , \36313 );
nand \U$40448 ( \40825 , \40823 , \40824 );
not \U$40449 ( \40826 , \40825 );
nand \U$40450 ( \40827 , \40819 , \40826 );
not \U$40451 ( \40828 , \40726 );
not \U$40452 ( \40829 , \40828 );
not \U$40453 ( \40830 , \40713 );
nor \U$40454 ( \40831 , \40830 , \40720 );
not \U$40455 ( \40832 , \40831 );
nand \U$40456 ( \40833 , \40829 , \40832 , \40189 , \40177 );
not \U$40457 ( \40834 , \39533 );
nor \U$40458 ( \40835 , \38647 , \40833 , \40785 , \40834 );
not \U$40459 ( \40836 , \29519 );
and \U$40460 ( \40837 , \10750 , \9541 );
not \U$40461 ( \40838 , \10750 );
and \U$40462 ( \40839 , \40838 , RIae7a7e0_186);
nor \U$40463 ( \40840 , \40837 , \40839 );
not \U$40464 ( \40841 , \40840 );
or \U$40465 ( \40842 , \40836 , \40841 );
not \U$40466 ( \40843 , \9529 );
not \U$40467 ( \40844 , \10007 );
or \U$40468 ( \40845 , \40843 , \40844 );
or \U$40469 ( \40846 , \10007 , \9541 );
nand \U$40470 ( \40847 , \40845 , \40846 );
nand \U$40471 ( \40848 , \40847 , \9549 );
nand \U$40472 ( \40849 , \40842 , \40848 );
not \U$40473 ( \40850 , \40849 );
not \U$40474 ( \40851 , \40850 );
not \U$40475 ( \40852 , \10676 );
and \U$40476 ( \40853 , RIae7a498_179, \11240 );
not \U$40477 ( \40854 , RIae7a498_179);
and \U$40478 ( \40855 , \40854 , \32565 );
or \U$40479 ( \40856 , \40853 , \40855 );
not \U$40480 ( \40857 , \40856 );
or \U$40481 ( \40858 , \40852 , \40857 );
xor \U$40482 ( \40859 , RIae7a498_179, \11321 );
nand \U$40483 ( \40860 , \40859 , \10695 );
nand \U$40484 ( \40861 , \40858 , \40860 );
not \U$40485 ( \40862 , \40861 );
not \U$40486 ( \40863 , \10631 );
not \U$40487 ( \40864 , \16164 );
not \U$40488 ( \40865 , RIae7a510_180);
and \U$40489 ( \40866 , \40864 , \40865 );
and \U$40490 ( \40867 , \16652 , RIae7a510_180);
nor \U$40491 ( \40868 , \40866 , \40867 );
not \U$40492 ( \40869 , \40868 );
or \U$40493 ( \40870 , \40863 , \40869 );
not \U$40494 ( \40871 , \17324 );
not \U$40495 ( \40872 , \18989 );
or \U$40496 ( \40873 , \40871 , \40872 );
not \U$40497 ( \40874 , \14931 );
nand \U$40498 ( \40875 , \40874 , \12750 );
nand \U$40499 ( \40876 , \40873 , \40875 );
nand \U$40500 ( \40877 , \40876 , \10637 );
nand \U$40501 ( \40878 , \40870 , \40877 );
not \U$40502 ( \40879 , \40878 );
nand \U$40503 ( \40880 , \12857 , \9620 );
not \U$40504 ( \40881 , \40880 );
and \U$40505 ( \40882 , \40879 , \40881 );
and \U$40506 ( \40883 , \40878 , \40880 );
nor \U$40507 ( \40884 , \40882 , \40883 );
not \U$40508 ( \40885 , \40884 );
not \U$40509 ( \40886 , \10675 );
not \U$40510 ( \40887 , \40859 );
or \U$40511 ( \40888 , \40886 , \40887 );
xnor \U$40512 ( \40889 , RIae7a498_179, \17155 );
nand \U$40513 ( \40890 , \40889 , \10695 );
nand \U$40514 ( \40891 , \40888 , \40890 );
and \U$40515 ( \40892 , \40885 , \40891 );
not \U$40516 ( \40893 , \40878 );
nor \U$40517 ( \40894 , \40893 , \40880 );
nor \U$40518 ( \40895 , \40892 , \40894 );
not \U$40519 ( \40896 , \40895 );
or \U$40520 ( \40897 , \40862 , \40896 );
or \U$40521 ( \40898 , \40895 , \40861 );
nand \U$40522 ( \40899 , \40897 , \40898 );
not \U$40523 ( \40900 , \40899 );
or \U$40524 ( \40901 , \40851 , \40900 );
or \U$40525 ( \40902 , \40899 , \40850 );
nand \U$40526 ( \40903 , \40901 , \40902 );
not \U$40527 ( \40904 , \40903 );
not \U$40528 ( \40905 , \10275 );
and \U$40529 ( \40906 , RIae7a8d0_188, \10084 );
not \U$40530 ( \40907 , RIae7a8d0_188);
and \U$40531 ( \40908 , \40907 , \38816 );
or \U$40532 ( \40909 , \40906 , \40908 );
not \U$40533 ( \40910 , \40909 );
or \U$40534 ( \40911 , \40905 , \40910 );
and \U$40535 ( \40912 , \10070 , RIae7a8d0_188);
not \U$40536 ( \40913 , \10070 );
and \U$40537 ( \40914 , \40913 , \18088 );
nor \U$40538 ( \40915 , \40912 , \40914 );
nand \U$40539 ( \40916 , \40915 , \11205 );
nand \U$40540 ( \40917 , \40911 , \40916 );
not \U$40541 ( \40918 , \40917 );
not \U$40542 ( \40919 , \9472 );
not \U$40543 ( \40920 , RIae7a6f0_184);
not \U$40544 ( \40921 , \9875 );
or \U$40545 ( \40922 , \40920 , \40921 );
or \U$40546 ( \40923 , \10750 , RIae7a6f0_184);
nand \U$40547 ( \40924 , \40922 , \40923 );
not \U$40548 ( \40925 , \40924 );
or \U$40549 ( \40926 , \40919 , \40925 );
and \U$40550 ( \40927 , RIae7a6f0_184, \10171 );
not \U$40551 ( \40928 , RIae7a6f0_184);
and \U$40552 ( \40929 , \40928 , \14546 );
or \U$40553 ( \40930 , \40927 , \40929 );
nand \U$40554 ( \40931 , \40930 , \9478 );
nand \U$40555 ( \40932 , \40926 , \40931 );
not \U$40556 ( \40933 , \10630 );
not \U$40557 ( \40934 , \40876 );
or \U$40558 ( \40935 , \40933 , \40934 );
not \U$40559 ( \40936 , \10636 );
not \U$40560 ( \40937 , \10633 );
not \U$40561 ( \40938 , \12857 );
or \U$40562 ( \40939 , \40937 , \40938 );
or \U$40563 ( \40940 , \12857 , \10633 );
nand \U$40564 ( \40941 , \40939 , \40940 );
nand \U$40565 ( \40942 , \40936 , \40941 );
nand \U$40566 ( \40943 , \40935 , \40942 );
not \U$40567 ( \40944 , \40943 );
not \U$40568 ( \40945 , \10628 );
not \U$40569 ( \40946 , \10625 );
or \U$40570 ( \40947 , \40945 , \40946 );
nand \U$40571 ( \40948 , \40947 , \12857 );
nand \U$40572 ( \40949 , \40948 , \24527 );
not \U$40573 ( \40950 , \40949 );
and \U$40574 ( \40951 , \40944 , \40950 );
and \U$40575 ( \40952 , \40943 , \40949 );
nor \U$40576 ( \40953 , \40951 , \40952 );
not \U$40577 ( \40954 , \40953 );
not \U$40578 ( \40955 , \10675 );
not \U$40579 ( \40956 , \40889 );
or \U$40580 ( \40957 , \40955 , \40956 );
not \U$40581 ( \40958 , \10625 );
not \U$40582 ( \40959 , \16652 );
or \U$40583 ( \40960 , \40958 , \40959 );
nand \U$40584 ( \40961 , \16651 , RIae7a498_179);
nand \U$40585 ( \40962 , \40960 , \40961 );
nand \U$40586 ( \40963 , \40962 , \10695 );
nand \U$40587 ( \40964 , \40957 , \40963 );
not \U$40588 ( \40965 , \40964 );
or \U$40589 ( \40966 , \40954 , \40965 );
or \U$40590 ( \40967 , \40964 , \40953 );
nand \U$40591 ( \40968 , \40966 , \40967 );
not \U$40592 ( \40969 , \40968 );
not \U$40593 ( \40970 , \9776 );
not \U$40594 ( \40971 , \10658 );
not \U$40595 ( \40972 , \10193 );
or \U$40596 ( \40973 , \40971 , \40972 );
nand \U$40597 ( \40974 , \11577 , RIae7a150_172);
nand \U$40598 ( \40975 , \40973 , \40974 );
not \U$40599 ( \40976 , \40975 );
or \U$40600 ( \40977 , \40970 , \40976 );
not \U$40601 ( \40978 , \10658 );
not \U$40602 ( \40979 , \12842 );
or \U$40603 ( \40980 , \40978 , \40979 );
or \U$40604 ( \40981 , \28259 , \10672 );
nand \U$40605 ( \40982 , \40980 , \40981 );
nand \U$40606 ( \40983 , \40982 , \9757 );
nand \U$40607 ( \40984 , \40977 , \40983 );
not \U$40608 ( \40985 , \40984 );
or \U$40609 ( \40986 , \40969 , \40985 );
not \U$40610 ( \40987 , \40953 );
nand \U$40611 ( \40988 , \40987 , \40964 );
nand \U$40612 ( \40989 , \40986 , \40988 );
xor \U$40613 ( \40990 , \40932 , \40989 );
not \U$40614 ( \40991 , \40990 );
or \U$40615 ( \40992 , \40918 , \40991 );
nand \U$40616 ( \40993 , \40932 , \40989 );
nand \U$40617 ( \40994 , \40992 , \40993 );
not \U$40618 ( \40995 , \40994 );
not \U$40619 ( \40996 , \40995 );
or \U$40620 ( \40997 , \40904 , \40996 );
or \U$40621 ( \40998 , \40995 , \40903 );
nand \U$40622 ( \40999 , \40997 , \40998 );
not \U$40623 ( \41000 , \40999 );
and \U$40624 ( \41001 , \40884 , \40891 );
nor \U$40625 ( \41002 , \40884 , \40891 );
nor \U$40626 ( \41003 , \41001 , \41002 );
not \U$40627 ( \41004 , \41003 );
not \U$40628 ( \41005 , \9549 );
and \U$40629 ( \41006 , RIae7a7e0_186, \37587 );
not \U$40630 ( \41007 , RIae7a7e0_186);
and \U$40631 ( \41008 , \41007 , \10743 );
or \U$40632 ( \41009 , \41006 , \41008 );
not \U$40633 ( \41010 , \41009 );
or \U$40634 ( \41011 , \41005 , \41010 );
nand \U$40635 ( \41012 , \40847 , \29518 );
nand \U$40636 ( \41013 , \41011 , \41012 );
not \U$40637 ( \41014 , \41013 );
and \U$40638 ( \41015 , \41004 , \41014 );
and \U$40639 ( \41016 , \41003 , \41013 );
nor \U$40640 ( \41017 , \41015 , \41016 );
not \U$40641 ( \41018 , \41017 );
not \U$40642 ( \41019 , \41018 );
not \U$40643 ( \41020 , \14667 );
not \U$40644 ( \41021 , RIae7aa38_191);
not \U$40645 ( \41022 , \10725 );
or \U$40646 ( \41023 , \41021 , \41022 );
not \U$40647 ( \41024 , \40194 );
or \U$40648 ( \41025 , \41024 , RIae7aa38_191);
nand \U$40649 ( \41026 , \41023 , \41025 );
not \U$40650 ( \41027 , \41026 );
or \U$40651 ( \41028 , \41020 , \41027 );
not \U$40652 ( \41029 , RIae7aa38_191);
not \U$40653 ( \41030 , \15501 );
or \U$40654 ( \41031 , \41029 , \41030 );
or \U$40655 ( \41032 , \10464 , RIae7aa38_191);
nand \U$40656 ( \41033 , \41031 , \41032 );
nand \U$40657 ( \41034 , \41033 , RIae7aab0_192);
nand \U$40658 ( \41035 , \41028 , \41034 );
not \U$40659 ( \41036 , \41035 );
or \U$40660 ( \41037 , \41019 , \41036 );
not \U$40661 ( \41038 , \41003 );
nand \U$40662 ( \41039 , \41038 , \41013 );
nand \U$40663 ( \41040 , \41037 , \41039 );
not \U$40664 ( \41041 , \41040 );
not \U$40665 ( \41042 , \41041 );
and \U$40666 ( \41043 , \41000 , \41042 );
and \U$40667 ( \41044 , \40999 , \41041 );
nor \U$40668 ( \41045 , \41043 , \41044 );
not \U$40669 ( \41046 , \41045 );
not \U$40670 ( \41047 , \11204 );
and \U$40671 ( \41048 , \9875 , \11207 );
not \U$40672 ( \41049 , \9875 );
and \U$40673 ( \41050 , \41049 , RIae7a8d0_188);
nor \U$40674 ( \41051 , \41048 , \41050 );
not \U$40675 ( \41052 , \41051 );
or \U$40676 ( \41053 , \41047 , \41052 );
xnor \U$40677 ( \41054 , \10171 , RIae7a8d0_188);
nand \U$40678 ( \41055 , \41054 , \10275 );
nand \U$40679 ( \41056 , \41053 , \41055 );
not \U$40680 ( \41057 , \41056 );
nand \U$40681 ( \41058 , \12857 , \10630 );
not \U$40682 ( \41059 , \41058 );
not \U$40683 ( \41060 , \10675 );
not \U$40684 ( \41061 , \40962 );
or \U$40685 ( \41062 , \41060 , \41061 );
not \U$40686 ( \41063 , RIae7a498_179);
not \U$40687 ( \41064 , \16006 );
or \U$40688 ( \41065 , \41063 , \41064 );
or \U$40689 ( \41066 , \16006 , RIae7a498_179);
nand \U$40690 ( \41067 , \41065 , \41066 );
nand \U$40691 ( \41068 , \41067 , \10695 );
nand \U$40692 ( \41069 , \41062 , \41068 );
not \U$40693 ( \41070 , \41069 );
or \U$40694 ( \41071 , \41059 , \41070 );
or \U$40695 ( \41072 , \41069 , \41058 );
nand \U$40696 ( \41073 , \41071 , \41072 );
not \U$40697 ( \41074 , \9776 );
not \U$40698 ( \41075 , \40982 );
or \U$40699 ( \41076 , \41074 , \41075 );
and \U$40700 ( \41077 , RIae7a150_172, \39806 );
not \U$40701 ( \41078 , RIae7a150_172);
and \U$40702 ( \41079 , \41078 , \28267 );
or \U$40703 ( \41080 , \41077 , \41079 );
nand \U$40704 ( \41081 , \41080 , \9757 );
nand \U$40705 ( \41082 , \41076 , \41081 );
xnor \U$40706 ( \41083 , \41073 , \41082 );
not \U$40707 ( \41084 , \41083 );
not \U$40708 ( \41085 , \41084 );
not \U$40709 ( \41086 , \9478 );
xor \U$40710 ( \41087 , RIae7a6f0_184, \10007 );
not \U$40711 ( \41088 , \41087 );
or \U$40712 ( \41089 , \41086 , \41088 );
not \U$40713 ( \41090 , RIae7a6f0_184);
not \U$40714 ( \41091 , \16193 );
or \U$40715 ( \41092 , \41090 , \41091 );
or \U$40716 ( \41093 , \10740 , RIae7a6f0_184);
nand \U$40717 ( \41094 , \41092 , \41093 );
nand \U$40718 ( \41095 , \41094 , \9472 );
nand \U$40719 ( \41096 , \41089 , \41095 );
not \U$40720 ( \41097 , \41096 );
not \U$40721 ( \41098 , \41097 );
or \U$40722 ( \41099 , \41085 , \41098 );
nand \U$40723 ( \41100 , \41096 , \41083 );
nand \U$40724 ( \41101 , \41099 , \41100 );
not \U$40725 ( \41102 , \41101 );
or \U$40726 ( \41103 , \41057 , \41102 );
nand \U$40727 ( \41104 , \41096 , \41084 );
nand \U$40728 ( \41105 , \41103 , \41104 );
not \U$40729 ( \41106 , \41105 );
xor \U$40730 ( \41107 , \40968 , \40984 );
not \U$40731 ( \41108 , \41107 );
or \U$40732 ( \41109 , RIae7a150_172, RIae7a420_178);
nand \U$40733 ( \41110 , \41109 , \12857 );
and \U$40734 ( \41111 , \41110 , \22054 );
not \U$40735 ( \41112 , \10675 );
not \U$40736 ( \41113 , \41067 );
or \U$40737 ( \41114 , \41112 , \41113 );
and \U$40738 ( \41115 , RIae7a498_179, \12857 );
not \U$40739 ( \41116 , RIae7a498_179);
and \U$40740 ( \41117 , \41116 , \17971 );
nor \U$40741 ( \41118 , \41115 , \41117 );
nand \U$40742 ( \41119 , \41118 , \10695 );
nand \U$40743 ( \41120 , \41114 , \41119 );
and \U$40744 ( \41121 , \41111 , \41120 );
not \U$40745 ( \41122 , \9744 );
not \U$40746 ( \41123 , \16912 );
not \U$40747 ( \41124 , \9749 );
or \U$40748 ( \41125 , \41123 , \41124 );
or \U$40749 ( \41126 , \10043 , \11102 );
nand \U$40750 ( \41127 , \41125 , \41126 );
not \U$40751 ( \41128 , \41127 );
or \U$40752 ( \41129 , \41122 , \41128 );
and \U$40753 ( \41130 , RIae7a060_170, \11240 );
not \U$40754 ( \41131 , RIae7a060_170);
and \U$40755 ( \41132 , \41131 , \11578 );
or \U$40756 ( \41133 , \41130 , \41132 );
nand \U$40757 ( \41134 , \41133 , \9728 );
nand \U$40758 ( \41135 , \41129 , \41134 );
xor \U$40759 ( \41136 , \41121 , \41135 );
not \U$40760 ( \41137 , \9549 );
not \U$40761 ( \41138 , RIae7a7e0_186);
not \U$40762 ( \41139 , \16922 );
or \U$40763 ( \41140 , \41138 , \41139 );
or \U$40764 ( \41141 , \16922 , RIae7a7e0_186);
nand \U$40765 ( \41142 , \41140 , \41141 );
not \U$40766 ( \41143 , \41142 );
or \U$40767 ( \41144 , \41137 , \41143 );
xor \U$40768 ( \41145 , \10142 , RIae7a7e0_186);
nand \U$40769 ( \41146 , \41145 , \29518 );
nand \U$40770 ( \41147 , \41144 , \41146 );
and \U$40771 ( \41148 , \41136 , \41147 );
and \U$40772 ( \41149 , \41121 , \41135 );
nor \U$40773 ( \41150 , \41148 , \41149 );
not \U$40774 ( \41151 , \41150 );
or \U$40775 ( \41152 , \41108 , \41151 );
or \U$40776 ( \41153 , \41150 , \41107 );
nand \U$40777 ( \41154 , \41152 , \41153 );
not \U$40778 ( \41155 , \41154 );
or \U$40779 ( \41156 , \41106 , \41155 );
not \U$40780 ( \41157 , \41150 );
nand \U$40781 ( \41158 , \41157 , \41107 );
nand \U$40782 ( \41159 , \41156 , \41158 );
not \U$40783 ( \41160 , \41159 );
not \U$40784 ( \41161 , \41035 );
not \U$40785 ( \41162 , \41017 );
and \U$40786 ( \41163 , \41161 , \41162 );
and \U$40787 ( \41164 , \41035 , \41017 );
nor \U$40788 ( \41165 , \41163 , \41164 );
not \U$40789 ( \41166 , \41165 );
not \U$40790 ( \41167 , \40917 );
not \U$40791 ( \41168 , \41167 );
not \U$40792 ( \41169 , \40990 );
or \U$40793 ( \41170 , \41168 , \41169 );
or \U$40794 ( \41171 , \40990 , \41167 );
nand \U$40795 ( \41172 , \41170 , \41171 );
not \U$40796 ( \41173 , \41172 );
or \U$40797 ( \41174 , \41166 , \41173 );
or \U$40798 ( \41175 , \41172 , \41165 );
nand \U$40799 ( \41176 , \41174 , \41175 );
not \U$40800 ( \41177 , \41176 );
or \U$40801 ( \41178 , \41160 , \41177 );
not \U$40802 ( \41179 , \41165 );
nand \U$40803 ( \41180 , \41179 , \41172 );
nand \U$40804 ( \41181 , \41178 , \41180 );
nand \U$40805 ( \41182 , \41046 , \41181 );
not \U$40806 ( \41183 , \41181 );
nand \U$40807 ( \41184 , \41045 , \41183 );
nand \U$40808 ( \41185 , \41182 , \41184 );
not \U$40809 ( \41186 , \10542 );
not \U$40810 ( \41187 , RIae7a060_170);
not \U$40811 ( \41188 , \27672 );
or \U$40812 ( \41189 , \41187 , \41188 );
or \U$40813 ( \41190 , \37587 , RIae7a060_170);
nand \U$40814 ( \41191 , \41189 , \41190 );
not \U$40815 ( \41192 , \41191 );
or \U$40816 ( \41193 , \41186 , \41192 );
and \U$40817 ( \41194 , RIae7a060_170, \10149 );
not \U$40818 ( \41195 , RIae7a060_170);
and \U$40819 ( \41196 , \41195 , \10142 );
or \U$40820 ( \41197 , \41194 , \41196 );
not \U$40821 ( \41198 , \41197 );
not \U$40822 ( \41199 , \9728 );
or \U$40823 ( \41200 , \41198 , \41199 );
nand \U$40824 ( \41201 , \41193 , \41200 );
not \U$40825 ( \41202 , \9478 );
xor \U$40826 ( \41203 , \10072 , RIae7a6f0_184);
not \U$40827 ( \41204 , \41203 );
or \U$40828 ( \41205 , \41202 , \41204 );
nand \U$40829 ( \41206 , \40930 , \9473 );
nand \U$40830 ( \41207 , \41205 , \41206 );
xor \U$40831 ( \41208 , \41201 , \41207 );
not \U$40832 ( \41209 , \10275 );
not \U$40833 ( \41210 , \40194 );
and \U$40834 ( \41211 , \41210 , RIae7a8d0_188);
not \U$40835 ( \41212 , \41210 );
and \U$40836 ( \41213 , \41212 , \11207 );
or \U$40837 ( \41214 , \41211 , \41213 );
not \U$40838 ( \41215 , \41214 );
or \U$40839 ( \41216 , \41209 , \41215 );
nand \U$40840 ( \41217 , \40909 , \11205 );
nand \U$40841 ( \41218 , \41216 , \41217 );
xor \U$40842 ( \41219 , \41208 , \41218 );
not \U$40843 ( \41220 , \41219 );
not \U$40844 ( \41221 , \41220 );
not \U$40845 ( \41222 , RIae7aab0_192);
and \U$40846 ( \41223 , \16752 , RIae7aa38_191);
not \U$40847 ( \41224 , \16752 );
and \U$40848 ( \41225 , \41224 , \11326 );
nor \U$40849 ( \41226 , \41223 , \41225 );
not \U$40850 ( \41227 , \41226 );
or \U$40851 ( \41228 , \41222 , \41227 );
nand \U$40852 ( \41229 , \41033 , \14668 );
nand \U$40853 ( \41230 , \41228 , \41229 );
not \U$40854 ( \41231 , \9776 );
and \U$40855 ( \41232 , \17955 , \10672 );
not \U$40856 ( \41233 , \17955 );
and \U$40857 ( \41234 , \41233 , RIae7a150_172);
nor \U$40858 ( \41235 , \41232 , \41234 );
not \U$40859 ( \41236 , \41235 );
or \U$40860 ( \41237 , \41231 , \41236 );
not \U$40861 ( \41238 , \10043 );
not \U$40862 ( \41239 , \10672 );
or \U$40863 ( \41240 , \41238 , \41239 );
or \U$40864 ( \41241 , \16912 , \9750 );
nand \U$40865 ( \41242 , \41240 , \41241 );
nand \U$40866 ( \41243 , \9758 , \41242 );
nand \U$40867 ( \41244 , \41237 , \41243 );
not \U$40868 ( \41245 , \10631 );
not \U$40869 ( \41246 , RIae7a510_180);
not \U$40870 ( \41247 , \11309 );
not \U$40871 ( \41248 , \41247 );
or \U$40872 ( \41249 , \41246 , \41248 );
or \U$40873 ( \41250 , RIae7a510_180, \39806 );
nand \U$40874 ( \41251 , \41249 , \41250 );
not \U$40875 ( \41252 , \41251 );
or \U$40876 ( \41253 , \41245 , \41252 );
nand \U$40877 ( \41254 , \40868 , \10637 );
nand \U$40878 ( \41255 , \41253 , \41254 );
not \U$40879 ( \41256 , \41255 );
not \U$40880 ( \41257 , \13165 );
not \U$40881 ( \41258 , \16009 );
or \U$40882 ( \41259 , \41257 , \41258 );
nand \U$40883 ( \41260 , \12750 , RIae7a3a8_177);
nand \U$40884 ( \41261 , \41259 , \41260 );
not \U$40885 ( \41262 , \41261 );
or \U$40886 ( \41263 , \41262 , \9637 );
and \U$40887 ( \41264 , RIae7a3a8_177, \17971 );
not \U$40888 ( \41265 , RIae7a3a8_177);
and \U$40889 ( \41266 , \41265 , \12857 );
nor \U$40890 ( \41267 , \41264 , \41266 );
not \U$40891 ( \41268 , \9643 );
or \U$40892 ( \41269 , \41267 , \41268 );
nand \U$40893 ( \41270 , \41263 , \41269 );
not \U$40894 ( \41271 , \41270 );
not \U$40895 ( \41272 , \25344 );
or \U$40896 ( \41273 , RIae7a510_180, RIae7a600_182);
nand \U$40897 ( \41274 , \41273 , \12857 );
nand \U$40898 ( \41275 , \41272 , \41274 );
not \U$40899 ( \41276 , \41275 );
and \U$40900 ( \41277 , \41271 , \41276 );
and \U$40901 ( \41278 , \41270 , \41275 );
nor \U$40902 ( \41279 , \41277 , \41278 );
not \U$40903 ( \41280 , \41279 );
and \U$40904 ( \41281 , \41256 , \41280 );
and \U$40905 ( \41282 , \41255 , \41279 );
nor \U$40906 ( \41283 , \41281 , \41282 );
and \U$40907 ( \41284 , \41244 , \41283 );
not \U$40908 ( \41285 , \41244 );
not \U$40909 ( \41286 , \41283 );
and \U$40910 ( \41287 , \41285 , \41286 );
or \U$40911 ( \41288 , \41284 , \41287 );
not \U$40912 ( \41289 , \41288 );
not \U$40913 ( \41290 , \9728 );
not \U$40914 ( \41291 , \9749 );
not \U$40915 ( \41292 , \16922 );
not \U$40916 ( \41293 , \41292 );
or \U$40917 ( \41294 , \41291 , \41293 );
nand \U$40918 ( \41295 , \16922 , RIae7a060_170);
nand \U$40919 ( \41296 , \41294 , \41295 );
not \U$40920 ( \41297 , \41296 );
or \U$40921 ( \41298 , \41290 , \41297 );
nand \U$40922 ( \41299 , \41197 , \9744 );
nand \U$40923 ( \41300 , \41298 , \41299 );
not \U$40924 ( \41301 , \41300 );
not \U$40925 ( \41302 , \40949 );
nand \U$40926 ( \41303 , \41302 , \40943 );
not \U$40927 ( \41304 , \41303 );
not \U$40928 ( \41305 , \9776 );
not \U$40929 ( \41306 , \41242 );
or \U$40930 ( \41307 , \41305 , \41306 );
nand \U$40931 ( \41308 , \40975 , \9757 );
nand \U$40932 ( \41309 , \41307 , \41308 );
not \U$40933 ( \41310 , \41309 );
or \U$40934 ( \41311 , \41304 , \41310 );
or \U$40935 ( \41312 , \41309 , \41303 );
nand \U$40936 ( \41313 , \41311 , \41312 );
not \U$40937 ( \41314 , \41313 );
or \U$40938 ( \41315 , \41301 , \41314 );
not \U$40939 ( \41316 , \41303 );
nand \U$40940 ( \41317 , \41316 , \41309 );
nand \U$40941 ( \41318 , \41315 , \41317 );
not \U$40942 ( \41319 , \41318 );
not \U$40943 ( \41320 , \41319 );
or \U$40944 ( \41321 , \41289 , \41320 );
or \U$40945 ( \41322 , \41319 , \41288 );
nand \U$40946 ( \41323 , \41321 , \41322 );
xor \U$40947 ( \41324 , \41230 , \41323 );
not \U$40948 ( \41325 , \41324 );
or \U$40949 ( \41326 , \41221 , \41325 );
not \U$40950 ( \41327 , \41324 );
nand \U$40951 ( \41328 , \41327 , \41219 );
nand \U$40952 ( \41329 , \41326 , \41328 );
not \U$40953 ( \41330 , \9478 );
not \U$40954 ( \41331 , \40924 );
or \U$40955 ( \41332 , \41330 , \41331 );
nand \U$40956 ( \41333 , \41087 , \9473 );
nand \U$40957 ( \41334 , \41332 , \41333 );
not \U$40958 ( \41335 , \10275 );
not \U$40959 ( \41336 , \40915 );
or \U$40960 ( \41337 , \41335 , \41336 );
nand \U$40961 ( \41338 , \41054 , \11205 );
nand \U$40962 ( \41339 , \41337 , \41338 );
xor \U$40963 ( \41340 , \41334 , \41339 );
not \U$40964 ( \41341 , RIae7aab0_192);
not \U$40965 ( \41342 , \41026 );
or \U$40966 ( \41343 , \41341 , \41342 );
not \U$40967 ( \41344 , \11326 );
not \U$40968 ( \41345 , \19025 );
or \U$40969 ( \41346 , \41344 , \41345 );
nand \U$40970 ( \41347 , \10084 , RIae7aa38_191);
nand \U$40971 ( \41348 , \41346 , \41347 );
nand \U$40972 ( \41349 , \41348 , \14667 );
nand \U$40973 ( \41350 , \41343 , \41349 );
and \U$40974 ( \41351 , \41340 , \41350 );
and \U$40975 ( \41352 , \41334 , \41339 );
or \U$40976 ( \41353 , \41351 , \41352 );
not \U$40977 ( \41354 , \41353 );
not \U$40978 ( \41355 , \41300 );
not \U$40979 ( \41356 , \41355 );
buf \U$40980 ( \41357 , \41313 );
not \U$40981 ( \41358 , \41357 );
or \U$40982 ( \41359 , \41356 , \41358 );
or \U$40983 ( \41360 , \41357 , \41355 );
nand \U$40984 ( \41361 , \41359 , \41360 );
not \U$40985 ( \41362 , \41361 );
not \U$40986 ( \41363 , \9527 );
not \U$40987 ( \41364 , \41009 );
or \U$40988 ( \41365 , \41363 , \41364 );
nand \U$40989 ( \41366 , \41145 , \9549 );
nand \U$40990 ( \41367 , \41365 , \41366 );
not \U$40991 ( \41368 , \41367 );
not \U$40992 ( \41369 , \41082 );
not \U$40993 ( \41370 , \41073 );
or \U$40994 ( \41371 , \41369 , \41370 );
not \U$40995 ( \41372 , \41058 );
nand \U$40996 ( \41373 , \41372 , \41069 );
nand \U$40997 ( \41374 , \41371 , \41373 );
not \U$40998 ( \41375 , \9744 );
not \U$40999 ( \41376 , \41296 );
or \U$41000 ( \41377 , \41375 , \41376 );
nand \U$41001 ( \41378 , \41127 , \9728 );
nand \U$41002 ( \41379 , \41377 , \41378 );
xor \U$41003 ( \41380 , \41374 , \41379 );
not \U$41004 ( \41381 , \41380 );
or \U$41005 ( \41382 , \41368 , \41381 );
nand \U$41006 ( \41383 , \41379 , \41374 );
nand \U$41007 ( \41384 , \41382 , \41383 );
not \U$41008 ( \41385 , \41384 );
not \U$41009 ( \41386 , \41385 );
or \U$41010 ( \41387 , \41362 , \41386 );
not \U$41011 ( \41388 , \41361 );
nand \U$41012 ( \41389 , \41388 , \41384 );
nand \U$41013 ( \41390 , \41387 , \41389 );
not \U$41014 ( \41391 , \41390 );
or \U$41015 ( \41392 , \41354 , \41391 );
nand \U$41016 ( \41393 , \41384 , \41361 );
nand \U$41017 ( \41394 , \41392 , \41393 );
not \U$41018 ( \41395 , \41394 );
and \U$41019 ( \41396 , \41329 , \41395 );
not \U$41020 ( \41397 , \41329 );
and \U$41021 ( \41398 , \41397 , \41394 );
nor \U$41022 ( \41399 , \41396 , \41398 );
xor \U$41023 ( \41400 , \41185 , \41399 );
not \U$41024 ( \41401 , \41159 );
and \U$41025 ( \41402 , \41176 , \41401 );
not \U$41026 ( \41403 , \41176 );
and \U$41027 ( \41404 , \41403 , \41159 );
nor \U$41028 ( \41405 , \41402 , \41404 );
not \U$41029 ( \41406 , \41405 );
not \U$41030 ( \41407 , \41406 );
not \U$41031 ( \41408 , \41353 );
and \U$41032 ( \41409 , \41390 , \41408 );
not \U$41033 ( \41410 , \41390 );
and \U$41034 ( \41411 , \41410 , \41353 );
nor \U$41035 ( \41412 , \41409 , \41411 );
not \U$41036 ( \41413 , \41412 );
not \U$41037 ( \41414 , \41367 );
not \U$41038 ( \41415 , \41414 );
not \U$41039 ( \41416 , \41380 );
or \U$41040 ( \41417 , \41415 , \41416 );
or \U$41041 ( \41418 , \41380 , \41414 );
nand \U$41042 ( \41419 , \41417 , \41418 );
xor \U$41043 ( \41420 , \41121 , \41135 );
xor \U$41044 ( \41421 , \41420 , \41147 );
not \U$41045 ( \41422 , \41421 );
not \U$41046 ( \41423 , \9744 );
not \U$41047 ( \41424 , \41133 );
or \U$41048 ( \41425 , \41423 , \41424 );
not \U$41049 ( \41426 , \9749 );
not \U$41050 ( \41427 , \10272 );
or \U$41051 ( \41428 , \41426 , \41427 );
or \U$41052 ( \41429 , \11318 , \9749 );
nand \U$41053 ( \41430 , \41428 , \41429 );
nand \U$41054 ( \41431 , \41430 , \9728 );
nand \U$41055 ( \41432 , \41425 , \41431 );
not \U$41056 ( \41433 , \41432 );
xor \U$41057 ( \41434 , \41111 , \41120 );
not \U$41058 ( \41435 , \9776 );
not \U$41059 ( \41436 , \41080 );
or \U$41060 ( \41437 , \41435 , \41436 );
not \U$41061 ( \41438 , \10672 );
not \U$41062 ( \41439 , \36790 );
or \U$41063 ( \41440 , \41438 , \41439 );
nand \U$41064 ( \41441 , \17166 , RIae7a150_172);
nand \U$41065 ( \41442 , \41440 , \41441 );
nand \U$41066 ( \41443 , \41442 , \9757 );
nand \U$41067 ( \41444 , \41437 , \41443 );
xor \U$41068 ( \41445 , \41434 , \41444 );
not \U$41069 ( \41446 , \41445 );
or \U$41070 ( \41447 , \41433 , \41446 );
nand \U$41071 ( \41448 , \41444 , \41434 );
nand \U$41072 ( \41449 , \41447 , \41448 );
not \U$41073 ( \41450 , \14667 );
and \U$41074 ( \41451 , RIae7aa38_191, \10071 );
not \U$41075 ( \41452 , RIae7aa38_191);
and \U$41076 ( \41453 , \41452 , \10072 );
or \U$41077 ( \41454 , \41451 , \41453 );
not \U$41078 ( \41455 , \41454 );
or \U$41079 ( \41456 , \41450 , \41455 );
nand \U$41080 ( \41457 , \41348 , RIae7aab0_192);
nand \U$41081 ( \41458 , \41456 , \41457 );
xor \U$41082 ( \41459 , \41449 , \41458 );
not \U$41083 ( \41460 , \41459 );
or \U$41084 ( \41461 , \41422 , \41460 );
nand \U$41085 ( \41462 , \41458 , \41449 );
nand \U$41086 ( \41463 , \41461 , \41462 );
xor \U$41087 ( \41464 , \41419 , \41463 );
xor \U$41088 ( \41465 , \41334 , \41339 );
xor \U$41089 ( \41466 , \41465 , \41350 );
and \U$41090 ( \41467 , \41464 , \41466 );
and \U$41091 ( \41468 , \41419 , \41463 );
or \U$41092 ( \41469 , \41467 , \41468 );
not \U$41093 ( \41470 , \41469 );
or \U$41094 ( \41471 , \41413 , \41470 );
or \U$41095 ( \41472 , \41469 , \41412 );
nand \U$41096 ( \41473 , \41471 , \41472 );
not \U$41097 ( \41474 , \41473 );
or \U$41098 ( \41475 , \41407 , \41474 );
not \U$41099 ( \41476 , \41412 );
nand \U$41100 ( \41477 , \41476 , \41469 );
nand \U$41101 ( \41478 , \41475 , \41477 );
nand \U$41102 ( \41479 , \41400 , \41478 );
not \U$41103 ( \41480 , \41479 );
not \U$41104 ( \41481 , \41406 );
not \U$41105 ( \41482 , \41473 );
not \U$41106 ( \41483 , \41482 );
or \U$41107 ( \41484 , \41481 , \41483 );
nand \U$41108 ( \41485 , \41473 , \41405 );
nand \U$41109 ( \41486 , \41484 , \41485 );
xnor \U$41110 ( \41487 , \41154 , \41105 );
not \U$41111 ( \41488 , \41487 );
not \U$41112 ( \41489 , RIae7aab0_192);
not \U$41113 ( \41490 , \41454 );
or \U$41114 ( \41491 , \41489 , \41490 );
xnor \U$41115 ( \41492 , \10171 , RIae7aa38_191);
nand \U$41116 ( \41493 , \41492 , \14667 );
nand \U$41117 ( \41494 , \41491 , \41493 );
not \U$41118 ( \41495 , \41494 );
not \U$41119 ( \41496 , \9478 );
not \U$41120 ( \41497 , \41094 );
or \U$41121 ( \41498 , \41496 , \41497 );
and \U$41122 ( \41499 , \40490 , \16101 );
not \U$41123 ( \41500 , \40490 );
and \U$41124 ( \41501 , \41500 , RIae7a6f0_184);
nor \U$41125 ( \41502 , \41499 , \41501 );
nand \U$41126 ( \41503 , \41502 , \9473 );
nand \U$41127 ( \41504 , \41498 , \41503 );
not \U$41128 ( \41505 , \41432 );
not \U$41129 ( \41506 , \41505 );
not \U$41130 ( \41507 , \41445 );
or \U$41131 ( \41508 , \41506 , \41507 );
or \U$41132 ( \41509 , \41445 , \41505 );
nand \U$41133 ( \41510 , \41508 , \41509 );
xor \U$41134 ( \41511 , \41504 , \41510 );
not \U$41135 ( \41512 , \41511 );
or \U$41136 ( \41513 , \41495 , \41512 );
nand \U$41137 ( \41514 , \41510 , \41504 );
nand \U$41138 ( \41515 , \41513 , \41514 );
not \U$41139 ( \41516 , \41515 );
not \U$41140 ( \41517 , \41056 );
not \U$41141 ( \41518 , \41517 );
not \U$41142 ( \41519 , \41101 );
or \U$41143 ( \41520 , \41518 , \41519 );
or \U$41144 ( \41521 , \41101 , \41517 );
nand \U$41145 ( \41522 , \41520 , \41521 );
not \U$41146 ( \41523 , \41522 );
not \U$41147 ( \41524 , \10275 );
not \U$41148 ( \41525 , \41051 );
or \U$41149 ( \41526 , \41524 , \41525 );
and \U$41150 ( \41527 , RIae7a8d0_188, \10000 );
not \U$41151 ( \41528 , RIae7a8d0_188);
and \U$41152 ( \41529 , \41528 , \10007 );
or \U$41153 ( \41530 , \41527 , \41529 );
nand \U$41154 ( \41531 , \41530 , \11204 );
nand \U$41155 ( \41532 , \41526 , \41531 );
not \U$41156 ( \41533 , \41532 );
and \U$41157 ( \41534 , \12857 , \10675 );
not \U$41158 ( \41535 , \9775 );
not \U$41159 ( \41536 , \41442 );
or \U$41160 ( \41537 , \41535 , \41536 );
and \U$41161 ( \41538 , \16006 , RIae7a150_172);
and \U$41162 ( \41539 , \16009 , \10658 );
nor \U$41163 ( \41540 , \41538 , \41539 );
or \U$41164 ( \41541 , \41540 , \9756 );
nand \U$41165 ( \41542 , \41537 , \41541 );
xor \U$41166 ( \41543 , \41534 , \41542 );
not \U$41167 ( \41544 , \9744 );
not \U$41168 ( \41545 , \41430 );
or \U$41169 ( \41546 , \41544 , \41545 );
and \U$41170 ( \41547 , RIae7a060_170, \39806 );
not \U$41171 ( \41548 , RIae7a060_170);
and \U$41172 ( \41549 , \41548 , \18971 );
or \U$41173 ( \41550 , \41547 , \41549 );
nand \U$41174 ( \41551 , \41550 , \9728 );
nand \U$41175 ( \41552 , \41546 , \41551 );
and \U$41176 ( \41553 , \41543 , \41552 );
and \U$41177 ( \41554 , \41534 , \41542 );
nor \U$41178 ( \41555 , \41553 , \41554 );
not \U$41179 ( \41556 , \41555 );
not \U$41180 ( \41557 , \29518 );
not \U$41181 ( \41558 , \41142 );
or \U$41182 ( \41559 , \41557 , \41558 );
not \U$41183 ( \41560 , \11665 );
not \U$41184 ( \41561 , \9537 );
or \U$41185 ( \41562 , \41560 , \41561 );
or \U$41186 ( \41563 , \16912 , \17112 );
nand \U$41187 ( \41564 , \41562 , \41563 );
nand \U$41188 ( \41565 , \41564 , \9549 );
nand \U$41189 ( \41566 , \41559 , \41565 );
not \U$41190 ( \41567 , \41566 );
or \U$41191 ( \41568 , \41556 , \41567 );
or \U$41192 ( \41569 , \41566 , \41555 );
nand \U$41193 ( \41570 , \41568 , \41569 );
not \U$41194 ( \41571 , \41570 );
or \U$41195 ( \41572 , \41533 , \41571 );
not \U$41196 ( \41573 , \41555 );
nand \U$41197 ( \41574 , \41573 , \41566 );
nand \U$41198 ( \41575 , \41572 , \41574 );
not \U$41199 ( \41576 , \41575 );
not \U$41200 ( \41577 , \41576 );
or \U$41201 ( \41578 , \41523 , \41577 );
not \U$41202 ( \41579 , \41522 );
nand \U$41203 ( \41580 , \41579 , \41575 );
nand \U$41204 ( \41581 , \41578 , \41580 );
not \U$41205 ( \41582 , \41581 );
or \U$41206 ( \41583 , \41516 , \41582 );
nand \U$41207 ( \41584 , \41575 , \41522 );
nand \U$41208 ( \41585 , \41583 , \41584 );
not \U$41209 ( \41586 , \41585 );
not \U$41210 ( \41587 , \41586 );
or \U$41211 ( \41588 , \41488 , \41587 );
xor \U$41212 ( \41589 , \41419 , \41463 );
xor \U$41213 ( \41590 , \41589 , \41466 );
nand \U$41214 ( \41591 , \41588 , \41590 );
not \U$41215 ( \41592 , \41487 );
nand \U$41216 ( \41593 , \41592 , \41585 );
nand \U$41217 ( \41594 , \41591 , \41593 );
nand \U$41218 ( \41595 , \41486 , \41594 );
not \U$41219 ( \41596 , \41595 );
or \U$41220 ( \41597 , \41480 , \41596 );
not \U$41221 ( \41598 , \41400 );
not \U$41222 ( \41599 , \41478 );
nand \U$41223 ( \41600 , \41598 , \41599 );
nand \U$41224 ( \41601 , \41597 , \41600 );
not \U$41225 ( \41602 , \41601 );
and \U$41226 ( \41603 , \12857 , \9699 );
not \U$41227 ( \41604 , \9620 );
not \U$41228 ( \41605 , \11690 );
not \U$41229 ( \41606 , \16652 );
or \U$41230 ( \41607 , \41605 , \41606 );
nand \U$41231 ( \41608 , \16651 , RIae7a3a8_177);
nand \U$41232 ( \41609 , \41607 , \41608 );
not \U$41233 ( \41610 , \41609 );
or \U$41234 ( \41611 , \41604 , \41610 );
nand \U$41235 ( \41612 , \41261 , \9643 );
nand \U$41236 ( \41613 , \41611 , \41612 );
xor \U$41237 ( \41614 , \41603 , \41613 );
not \U$41238 ( \41615 , \10631 );
not \U$41239 ( \41616 , \10633 );
not \U$41240 ( \41617 , \10272 );
or \U$41241 ( \41618 , \41616 , \41617 );
or \U$41242 ( \41619 , \11318 , \14931 );
nand \U$41243 ( \41620 , \41618 , \41619 );
not \U$41244 ( \41621 , \41620 );
or \U$41245 ( \41622 , \41615 , \41621 );
nand \U$41246 ( \41623 , \41251 , \10637 );
nand \U$41247 ( \41624 , \41622 , \41623 );
xnor \U$41248 ( \41625 , \41614 , \41624 );
not \U$41249 ( \41626 , \41625 );
not \U$41250 ( \41627 , \9549 );
not \U$41251 ( \41628 , \40840 );
or \U$41252 ( \41629 , \41627 , \41628 );
and \U$41253 ( \41630 , RIae7a7e0_186, \10171 );
not \U$41254 ( \41631 , RIae7a7e0_186);
and \U$41255 ( \41632 , \41631 , \13544 );
or \U$41256 ( \41633 , \41630 , \41632 );
nand \U$41257 ( \41634 , \41633 , \29519 );
nand \U$41258 ( \41635 , \41629 , \41634 );
not \U$41259 ( \41636 , \41635 );
or \U$41260 ( \41637 , \41626 , \41636 );
or \U$41261 ( \41638 , \41635 , \41625 );
nand \U$41262 ( \41639 , \41637 , \41638 );
not \U$41263 ( \41640 , \9728 );
not \U$41264 ( \41641 , \41191 );
or \U$41265 ( \41642 , \41640 , \41641 );
and \U$41266 ( \41643 , \11102 , \10000 );
not \U$41267 ( \41644 , \11102 );
and \U$41268 ( \41645 , \41644 , \10007 );
nor \U$41269 ( \41646 , \41643 , \41645 );
nand \U$41270 ( \41647 , \41646 , \9745 );
nand \U$41271 ( \41648 , \41642 , \41647 );
xor \U$41272 ( \41649 , \41639 , \41648 );
not \U$41273 ( \41650 , \40849 );
not \U$41274 ( \41651 , \40899 );
or \U$41275 ( \41652 , \41650 , \41651 );
not \U$41276 ( \41653 , \40895 );
nand \U$41277 ( \41654 , \41653 , \40861 );
nand \U$41278 ( \41655 , \41652 , \41654 );
not \U$41279 ( \41656 , \41286 );
not \U$41280 ( \41657 , \41244 );
or \U$41281 ( \41658 , \41656 , \41657 );
not \U$41282 ( \41659 , \41279 );
nand \U$41283 ( \41660 , \41659 , \41255 );
nand \U$41284 ( \41661 , \41658 , \41660 );
not \U$41285 ( \41662 , \41661 );
not \U$41286 ( \41663 , \41662 );
not \U$41287 ( \41664 , \41275 );
nand \U$41288 ( \41665 , \41664 , \41270 );
not \U$41289 ( \41666 , \41665 );
not \U$41290 ( \41667 , \10675 );
not \U$41291 ( \41668 , \10625 );
not \U$41292 ( \41669 , \10043 );
or \U$41293 ( \41670 , \41668 , \41669 );
or \U$41294 ( \41671 , \16912 , \10625 );
nand \U$41295 ( \41672 , \41670 , \41671 );
not \U$41296 ( \41673 , \41672 );
or \U$41297 ( \41674 , \41667 , \41673 );
nand \U$41298 ( \41675 , \40856 , \10695 );
nand \U$41299 ( \41676 , \41674 , \41675 );
not \U$41300 ( \41677 , \41676 );
or \U$41301 ( \41678 , \41666 , \41677 );
or \U$41302 ( \41679 , \41676 , \41665 );
nand \U$41303 ( \41680 , \41678 , \41679 );
buf \U$41304 ( \41681 , \41680 );
not \U$41305 ( \41682 , \10667 );
not \U$41306 ( \41683 , \41235 );
or \U$41307 ( \41684 , \41682 , \41683 );
not \U$41308 ( \41685 , RIae7a150_172);
not \U$41309 ( \41686 , \10149 );
or \U$41310 ( \41687 , \41685 , \41686 );
or \U$41311 ( \41688 , \10149 , RIae7a150_172);
nand \U$41312 ( \41689 , \41687 , \41688 );
nand \U$41313 ( \41690 , \41689 , \9776 );
nand \U$41314 ( \41691 , \41684 , \41690 );
and \U$41315 ( \41692 , \41681 , \41691 );
not \U$41316 ( \41693 , \41681 );
not \U$41317 ( \41694 , \41691 );
and \U$41318 ( \41695 , \41693 , \41694 );
nor \U$41319 ( \41696 , \41692 , \41695 );
not \U$41320 ( \41697 , \41696 );
or \U$41321 ( \41698 , \41663 , \41697 );
or \U$41322 ( \41699 , \41696 , \41662 );
nand \U$41323 ( \41700 , \41698 , \41699 );
xor \U$41324 ( \41701 , \41655 , \41700 );
xor \U$41325 ( \41702 , \41649 , \41701 );
not \U$41326 ( \41703 , \41040 );
not \U$41327 ( \41704 , \40999 );
or \U$41328 ( \41705 , \41703 , \41704 );
nand \U$41329 ( \41706 , \40994 , \40903 );
nand \U$41330 ( \41707 , \41705 , \41706 );
xor \U$41331 ( \41708 , \41702 , \41707 );
not \U$41332 ( \41709 , \41708 );
xor \U$41333 ( \41710 , \41201 , \41207 );
and \U$41334 ( \41711 , \41710 , \41218 );
and \U$41335 ( \41712 , \41201 , \41207 );
or \U$41336 ( \41713 , \41711 , \41712 );
not \U$41337 ( \41714 , \41230 );
not \U$41338 ( \41715 , \41323 );
or \U$41339 ( \41716 , \41714 , \41715 );
not \U$41340 ( \41717 , \41319 );
nand \U$41341 ( \41718 , \41717 , \41288 );
nand \U$41342 ( \41719 , \41716 , \41718 );
xor \U$41343 ( \41720 , \41713 , \41719 );
not \U$41344 ( \41721 , \14668 );
not \U$41345 ( \41722 , \41226 );
or \U$41346 ( \41723 , \41721 , \41722 );
and \U$41347 ( \41724 , \11195 , \11326 );
not \U$41348 ( \41725 , \11195 );
and \U$41349 ( \41726 , \41725 , RIae7aa38_191);
nor \U$41350 ( \41727 , \41724 , \41726 );
not \U$41351 ( \41728 , \41727 );
or \U$41352 ( \41729 , \41728 , \14666 );
nand \U$41353 ( \41730 , \41723 , \41729 );
not \U$41354 ( \41731 , \9478 );
and \U$41355 ( \41732 , RIae7a6f0_184, \10084 );
not \U$41356 ( \41733 , RIae7a6f0_184);
and \U$41357 ( \41734 , \41733 , \19025 );
or \U$41358 ( \41735 , \41732 , \41734 );
not \U$41359 ( \41736 , \41735 );
or \U$41360 ( \41737 , \41731 , \41736 );
nand \U$41361 ( \41738 , \41203 , \9473 );
nand \U$41362 ( \41739 , \41737 , \41738 );
not \U$41363 ( \41740 , \16594 );
not \U$41364 ( \41741 , \41214 );
or \U$41365 ( \41742 , \41740 , \41741 );
and \U$41366 ( \41743 , RIae7a8d0_188, \10461 );
not \U$41367 ( \41744 , RIae7a8d0_188);
and \U$41368 ( \41745 , \41744 , \10465 );
or \U$41369 ( \41746 , \41743 , \41745 );
nand \U$41370 ( \41747 , \41746 , \10275 );
nand \U$41371 ( \41748 , \41742 , \41747 );
xor \U$41372 ( \41749 , \41739 , \41748 );
xor \U$41373 ( \41750 , \41730 , \41749 );
xnor \U$41374 ( \41751 , \41720 , \41750 );
not \U$41375 ( \41752 , \41394 );
not \U$41376 ( \41753 , \41329 );
or \U$41377 ( \41754 , \41752 , \41753 );
nand \U$41378 ( \41755 , \41324 , \41219 );
nand \U$41379 ( \41756 , \41754 , \41755 );
or \U$41380 ( \41757 , \41751 , \41756 );
nand \U$41381 ( \41758 , \41756 , \41751 );
nand \U$41382 ( \41759 , \41757 , \41758 );
not \U$41383 ( \41760 , \41759 );
or \U$41384 ( \41761 , \41709 , \41760 );
or \U$41385 ( \41762 , \41759 , \41708 );
nand \U$41386 ( \41763 , \41761 , \41762 );
not \U$41387 ( \41764 , \41182 );
not \U$41388 ( \41765 , \41399 );
or \U$41389 ( \41766 , \41764 , \41765 );
nand \U$41390 ( \41767 , \41766 , \41184 );
nand \U$41391 ( \41768 , \41763 , \41767 );
nand \U$41392 ( \41769 , \41602 , \41768 );
or \U$41393 ( \41770 , \41763 , \41767 );
nand \U$41394 ( \41771 , \41769 , \41770 );
or \U$41395 ( \41772 , \41719 , \41713 );
nand \U$41396 ( \41773 , \41772 , \41750 );
nand \U$41397 ( \41774 , \41719 , \41713 );
nand \U$41398 ( \41775 , \41773 , \41774 );
not \U$41399 ( \41776 , \41775 );
not \U$41400 ( \41777 , \41776 );
not \U$41401 ( \41778 , RIae7aab0_192);
and \U$41402 ( \41779 , \19422 , \11326 );
not \U$41403 ( \41780 , \19422 );
and \U$41404 ( \41781 , \41780 , RIae7aa38_191);
nor \U$41405 ( \41782 , \41779 , \41781 );
not \U$41406 ( \41783 , \41782 );
or \U$41407 ( \41784 , \41778 , \41783 );
nand \U$41408 ( \41785 , \41727 , \14667 );
nand \U$41409 ( \41786 , \41784 , \41785 );
not \U$41410 ( \41787 , \41624 );
not \U$41411 ( \41788 , \41614 );
or \U$41412 ( \41789 , \41787 , \41788 );
nand \U$41413 ( \41790 , \41613 , \41603 );
nand \U$41414 ( \41791 , \41789 , \41790 );
not \U$41415 ( \41792 , \10675 );
not \U$41416 ( \41793 , \11427 );
not \U$41417 ( \41794 , \41292 );
or \U$41418 ( \41795 , \41793 , \41794 );
nand \U$41419 ( \41796 , \11589 , RIae7a498_179);
nand \U$41420 ( \41797 , \41795 , \41796 );
not \U$41421 ( \41798 , \41797 );
or \U$41422 ( \41799 , \41792 , \41798 );
nand \U$41423 ( \41800 , \41672 , \10695 );
nand \U$41424 ( \41801 , \41799 , \41800 );
xor \U$41425 ( \41802 , \41791 , \41801 );
not \U$41426 ( \41803 , \29519 );
and \U$41427 ( \41804 , RIae7a7e0_186, \11230 );
not \U$41428 ( \41805 , RIae7a7e0_186);
and \U$41429 ( \41806 , \41805 , \10072 );
or \U$41430 ( \41807 , \41804 , \41806 );
not \U$41431 ( \41808 , \41807 );
or \U$41432 ( \41809 , \41803 , \41808 );
nand \U$41433 ( \41810 , \41633 , \9549 );
nand \U$41434 ( \41811 , \41809 , \41810 );
not \U$41435 ( \41812 , \41811 );
and \U$41436 ( \41813 , \41802 , \41812 );
not \U$41437 ( \41814 , \41802 );
and \U$41438 ( \41815 , \41814 , \41811 );
nor \U$41439 ( \41816 , \41813 , \41815 );
xor \U$41440 ( \41817 , \41786 , \41816 );
not \U$41441 ( \41818 , \41648 );
not \U$41442 ( \41819 , \41639 );
or \U$41443 ( \41820 , \41818 , \41819 );
not \U$41444 ( \41821 , \41625 );
nand \U$41445 ( \41822 , \41821 , \41635 );
nand \U$41446 ( \41823 , \41820 , \41822 );
xor \U$41447 ( \41824 , \41817 , \41823 );
not \U$41448 ( \41825 , \41655 );
not \U$41449 ( \41826 , \41700 );
or \U$41450 ( \41827 , \41825 , \41826 );
not \U$41451 ( \41828 , \41662 );
nand \U$41452 ( \41829 , \41828 , \41696 );
nand \U$41453 ( \41830 , \41827 , \41829 );
xnor \U$41454 ( \41831 , \41824 , \41830 );
not \U$41455 ( \41832 , \41831 );
or \U$41456 ( \41833 , \41777 , \41832 );
or \U$41457 ( \41834 , \41831 , \41776 );
nand \U$41458 ( \41835 , \41833 , \41834 );
not \U$41459 ( \41836 , \41835 );
xor \U$41460 ( \41837 , \41649 , \41701 );
and \U$41461 ( \41838 , \41837 , \41707 );
and \U$41462 ( \41839 , \41649 , \41701 );
or \U$41463 ( \41840 , \41838 , \41839 );
not \U$41464 ( \41841 , \41840 );
not \U$41465 ( \41842 , \41841 );
not \U$41466 ( \41843 , \41730 );
not \U$41467 ( \41844 , \41749 );
or \U$41468 ( \41845 , \41843 , \41844 );
nand \U$41469 ( \41846 , \41748 , \41739 );
nand \U$41470 ( \41847 , \41845 , \41846 );
not \U$41471 ( \41848 , \9744 );
not \U$41472 ( \41849 , RIae7a060_170);
not \U$41473 ( \41850 , \9875 );
or \U$41474 ( \41851 , \41849 , \41850 );
or \U$41475 ( \41852 , \13896 , RIae7a060_170);
nand \U$41476 ( \41853 , \41851 , \41852 );
not \U$41477 ( \41854 , \41853 );
or \U$41478 ( \41855 , \41848 , \41854 );
nand \U$41479 ( \41856 , \41646 , \9728 );
nand \U$41480 ( \41857 , \41855 , \41856 );
not \U$41481 ( \41858 , \9776 );
xnor \U$41482 ( \41859 , \10740 , RIae7a150_172);
not \U$41483 ( \41860 , \41859 );
or \U$41484 ( \41861 , \41858 , \41860 );
nand \U$41485 ( \41862 , \41689 , \10667 );
nand \U$41486 ( \41863 , \41861 , \41862 );
or \U$41487 ( \41864 , \41857 , \41863 );
nand \U$41488 ( \41865 , \41857 , \41863 );
nand \U$41489 ( \41866 , \41864 , \41865 );
not \U$41490 ( \41867 , \9478 );
not \U$41491 ( \41868 , RIae7a6f0_184);
not \U$41492 ( \41869 , \10725 );
or \U$41493 ( \41870 , \41868 , \41869 );
not \U$41494 ( \41871 , \35832 );
nand \U$41495 ( \41872 , \41871 , \16104 );
nand \U$41496 ( \41873 , \41870 , \41872 );
not \U$41497 ( \41874 , \41873 );
or \U$41498 ( \41875 , \41867 , \41874 );
nand \U$41499 ( \41876 , \41735 , \9473 );
nand \U$41500 ( \41877 , \41875 , \41876 );
xor \U$41501 ( \41878 , \41866 , \41877 );
not \U$41502 ( \41879 , \41878 );
not \U$41503 ( \41880 , \41879 );
not \U$41504 ( \41881 , \10275 );
and \U$41505 ( \41882 , \16752 , RIae7a8d0_188);
not \U$41506 ( \41883 , \16752 );
and \U$41507 ( \41884 , \41883 , \18088 );
nor \U$41508 ( \41885 , \41882 , \41884 );
not \U$41509 ( \41886 , \41885 );
or \U$41510 ( \41887 , \41881 , \41886 );
nand \U$41511 ( \41888 , \41746 , \16594 );
nand \U$41512 ( \41889 , \41887 , \41888 );
not \U$41513 ( \41890 , \41889 );
not \U$41514 ( \41891 , \41890 );
not \U$41515 ( \41892 , \10631 );
and \U$41516 ( \41893 , RIae7a510_180, \11240 );
not \U$41517 ( \41894 , RIae7a510_180);
and \U$41518 ( \41895 , \41894 , \30081 );
or \U$41519 ( \41896 , \41893 , \41895 );
not \U$41520 ( \41897 , \41896 );
or \U$41521 ( \41898 , \41892 , \41897 );
nand \U$41522 ( \41899 , \41620 , \10637 );
nand \U$41523 ( \41900 , \41898 , \41899 );
or \U$41524 ( \41901 , RIae7a330_176, RIae7a3a8_177);
nand \U$41525 ( \41902 , \41901 , \12857 );
and \U$41526 ( \41903 , RIae7a330_176, RIae7a3a8_177);
nor \U$41527 ( \41904 , \41903 , \38064 );
and \U$41528 ( \41905 , \41902 , \41904 );
not \U$41529 ( \41906 , \9699 );
buf \U$41530 ( \41907 , \12750 );
and \U$41531 ( \41908 , \11114 , \41907 );
not \U$41532 ( \41909 , \11114 );
and \U$41533 ( \41910 , \41909 , \16009 );
nor \U$41534 ( \41911 , \41908 , \41910 );
not \U$41535 ( \41912 , \41911 );
or \U$41536 ( \41913 , \41906 , \41912 );
xnor \U$41537 ( \41914 , \36545 , RIae7a240_174);
nand \U$41538 ( \41915 , \41914 , \9687 );
nand \U$41539 ( \41916 , \41913 , \41915 );
xor \U$41540 ( \41917 , \41905 , \41916 );
not \U$41541 ( \41918 , \41917 );
not \U$41542 ( \41919 , \13165 );
not \U$41543 ( \41920 , \39806 );
not \U$41544 ( \41921 , \41920 );
or \U$41545 ( \41922 , \41919 , \41921 );
nand \U$41546 ( \41923 , \41247 , RIae7a3a8_177);
nand \U$41547 ( \41924 , \41922 , \41923 );
and \U$41548 ( \41925 , \9621 , \41924 );
and \U$41549 ( \41926 , \41609 , \9643 );
nor \U$41550 ( \41927 , \41925 , \41926 );
not \U$41551 ( \41928 , \41927 );
or \U$41552 ( \41929 , \41918 , \41928 );
or \U$41553 ( \41930 , \41927 , \41917 );
nand \U$41554 ( \41931 , \41929 , \41930 );
xor \U$41555 ( \41932 , \41900 , \41931 );
not \U$41556 ( \41933 , \41691 );
not \U$41557 ( \41934 , \41680 );
or \U$41558 ( \41935 , \41933 , \41934 );
not \U$41559 ( \41936 , \41665 );
nand \U$41560 ( \41937 , \41936 , \41676 );
nand \U$41561 ( \41938 , \41935 , \41937 );
xor \U$41562 ( \41939 , \41932 , \41938 );
not \U$41563 ( \41940 , \41939 );
or \U$41564 ( \41941 , \41891 , \41940 );
or \U$41565 ( \41942 , \41939 , \41890 );
nand \U$41566 ( \41943 , \41941 , \41942 );
not \U$41567 ( \41944 , \41943 );
not \U$41568 ( \41945 , \41944 );
or \U$41569 ( \41946 , \41880 , \41945 );
nand \U$41570 ( \41947 , \41943 , \41878 );
nand \U$41571 ( \41948 , \41946 , \41947 );
not \U$41572 ( \41949 , \41948 );
and \U$41573 ( \41950 , \41847 , \41949 );
not \U$41574 ( \41951 , \41847 );
and \U$41575 ( \41952 , \41951 , \41948 );
or \U$41576 ( \41953 , \41950 , \41952 );
not \U$41577 ( \41954 , \41953 );
or \U$41578 ( \41955 , \41842 , \41954 );
or \U$41579 ( \41956 , \41953 , \41841 );
nand \U$41580 ( \41957 , \41955 , \41956 );
not \U$41581 ( \41958 , \41957 );
or \U$41582 ( \41959 , \41836 , \41958 );
or \U$41583 ( \41960 , \41957 , \41835 );
nand \U$41584 ( \41961 , \41959 , \41960 );
not \U$41585 ( \41962 , \41708 );
not \U$41586 ( \41963 , \41962 );
not \U$41587 ( \41964 , \41759 );
or \U$41588 ( \41965 , \41963 , \41964 );
not \U$41589 ( \41966 , \41756 );
nand \U$41590 ( \41967 , \41966 , \41751 );
nand \U$41591 ( \41968 , \41965 , \41967 );
nand \U$41592 ( \41969 , \41961 , \41968 );
nand \U$41593 ( \41970 , \41771 , \41969 );
xor \U$41594 ( \41971 , \41552 , \41543 );
not \U$41595 ( \41972 , \11204 );
not \U$41596 ( \41973 , RIae7a8d0_188);
not \U$41597 ( \41974 , \27672 );
or \U$41598 ( \41975 , \41973 , \41974 );
or \U$41599 ( \41976 , \37587 , RIae7a8d0_188);
nand \U$41600 ( \41977 , \41975 , \41976 );
not \U$41601 ( \41978 , \41977 );
or \U$41602 ( \41979 , \41972 , \41978 );
nand \U$41603 ( \41980 , \41530 , \10275 );
nand \U$41604 ( \41981 , \41979 , \41980 );
xor \U$41605 ( \41982 , \41971 , \41981 );
not \U$41606 ( \41983 , \14667 );
and \U$41607 ( \41984 , RIae7aa38_191, \9868 );
not \U$41608 ( \41985 , RIae7aa38_191);
and \U$41609 ( \41986 , \41985 , \10750 );
nor \U$41610 ( \41987 , \41984 , \41986 );
not \U$41611 ( \41988 , \41987 );
or \U$41612 ( \41989 , \41983 , \41988 );
nand \U$41613 ( \41990 , \41492 , RIae7aab0_192);
nand \U$41614 ( \41991 , \41989 , \41990 );
and \U$41615 ( \41992 , \41982 , \41991 );
and \U$41616 ( \41993 , \41971 , \41981 );
or \U$41617 ( \41994 , \41992 , \41993 );
not \U$41618 ( \41995 , \41994 );
not \U$41619 ( \41996 , \41995 );
not \U$41620 ( \41997 , \9775 );
or \U$41621 ( \41998 , \41540 , \41997 );
and \U$41622 ( \41999 , \16890 , RIae7a150_172);
and \U$41623 ( \42000 , \12858 , \10658 );
nor \U$41624 ( \42001 , \41999 , \42000 );
or \U$41625 ( \42002 , \42001 , \9756 );
nand \U$41626 ( \42003 , \41998 , \42002 );
and \U$41627 ( \42004 , \12857 , \9773 );
nor \U$41628 ( \42005 , \42004 , \21099 );
and \U$41629 ( \42006 , \42003 , \42005 );
not \U$41630 ( \42007 , \29518 );
not \U$41631 ( \42008 , \41564 );
or \U$41632 ( \42009 , \42007 , \42008 );
not \U$41633 ( \42010 , RIae7a7e0_186);
not \U$41634 ( \42011 , \11577 );
or \U$41635 ( \42012 , \42010 , \42011 );
or \U$41636 ( \42013 , \10194 , RIae7a7e0_186);
nand \U$41637 ( \42014 , \42012 , \42013 );
nand \U$41638 ( \42015 , \42014 , \9549 );
nand \U$41639 ( \42016 , \42009 , \42015 );
xor \U$41640 ( \42017 , \42006 , \42016 );
not \U$41641 ( \42018 , \9473 );
and \U$41642 ( \42019 , \32534 , RIae7a6f0_184);
not \U$41643 ( \42020 , \32534 );
and \U$41644 ( \42021 , \42020 , \16101 );
nor \U$41645 ( \42022 , \42019 , \42021 );
not \U$41646 ( \42023 , \42022 );
or \U$41647 ( \42024 , \42018 , \42023 );
nand \U$41648 ( \42025 , \41502 , \9478 );
nand \U$41649 ( \42026 , \42024 , \42025 );
and \U$41650 ( \42027 , \42017 , \42026 );
and \U$41651 ( \42028 , \42006 , \42016 );
nor \U$41652 ( \42029 , \42027 , \42028 );
not \U$41653 ( \42030 , \42029 );
not \U$41654 ( \42031 , \41570 );
not \U$41655 ( \42032 , \41532 );
not \U$41656 ( \42033 , \42032 );
and \U$41657 ( \42034 , \42031 , \42033 );
and \U$41658 ( \42035 , \41570 , \42032 );
nor \U$41659 ( \42036 , \42034 , \42035 );
not \U$41660 ( \42037 , \42036 );
not \U$41661 ( \42038 , \42037 );
or \U$41662 ( \42039 , \42030 , \42038 );
not \U$41663 ( \42040 , \42029 );
nand \U$41664 ( \42041 , \42040 , \42036 );
nand \U$41665 ( \42042 , \42039 , \42041 );
not \U$41666 ( \42043 , \42042 );
or \U$41667 ( \42044 , \41996 , \42043 );
or \U$41668 ( \42045 , \42042 , \41995 );
nand \U$41669 ( \42046 , \42044 , \42045 );
not \U$41670 ( \42047 , \42046 );
not \U$41671 ( \42048 , \42047 );
xnor \U$41672 ( \42049 , \41511 , \41494 );
not \U$41673 ( \42050 , \42049 );
not \U$41674 ( \42051 , \10275 );
not \U$41675 ( \42052 , \41977 );
or \U$41676 ( \42053 , \42051 , \42052 );
not \U$41677 ( \42054 , \40490 );
not \U$41678 ( \42055 , RIae7a8d0_188);
and \U$41679 ( \42056 , \42054 , \42055 );
and \U$41680 ( \42057 , \40490 , RIae7a8d0_188);
nor \U$41681 ( \42058 , \42056 , \42057 );
not \U$41682 ( \42059 , \11204 );
or \U$41683 ( \42060 , \42058 , \42059 );
nand \U$41684 ( \42061 , \42053 , \42060 );
not \U$41685 ( \42062 , \42061 );
not \U$41686 ( \42063 , \9744 );
not \U$41687 ( \42064 , \16652 );
not \U$41688 ( \42065 , RIae7a060_170);
and \U$41689 ( \42066 , \42064 , \42065 );
and \U$41690 ( \42067 , \36790 , RIae7a060_170);
nor \U$41691 ( \42068 , \42066 , \42067 );
not \U$41692 ( \42069 , \42068 );
or \U$41693 ( \42070 , \42063 , \42069 );
not \U$41694 ( \42071 , RIae7a060_170);
not \U$41695 ( \42072 , \16006 );
or \U$41696 ( \42073 , \42071 , \42072 );
or \U$41697 ( \42074 , \16006 , RIae7a060_170);
nand \U$41698 ( \42075 , \42073 , \42074 );
nand \U$41699 ( \42076 , \42075 , \9728 );
nand \U$41700 ( \42077 , \42070 , \42076 );
and \U$41701 ( \42078 , \12857 , \9775 );
xor \U$41702 ( \42079 , \42077 , \42078 );
not \U$41703 ( \42080 , \42079 );
not \U$41704 ( \42081 , \29518 );
not \U$41705 ( \42082 , \10272 );
not \U$41706 ( \42083 , RIae7a7e0_186);
and \U$41707 ( \42084 , \42082 , \42083 );
and \U$41708 ( \42085 , \11321 , RIae7a7e0_186);
nor \U$41709 ( \42086 , \42084 , \42085 );
not \U$41710 ( \42087 , \42086 );
or \U$41711 ( \42088 , \42081 , \42087 );
and \U$41712 ( \42089 , RIae7a7e0_186, \39806 );
not \U$41713 ( \42090 , RIae7a7e0_186);
and \U$41714 ( \42091 , \42090 , \18971 );
or \U$41715 ( \42092 , \42089 , \42091 );
nand \U$41716 ( \42093 , \42092 , \9549 );
nand \U$41717 ( \42094 , \42088 , \42093 );
not \U$41718 ( \42095 , \42094 );
or \U$41719 ( \42096 , \42080 , \42095 );
nand \U$41720 ( \42097 , \42077 , \42078 );
nand \U$41721 ( \42098 , \42096 , \42097 );
not \U$41722 ( \42099 , \9478 );
not \U$41723 ( \42100 , \42022 );
or \U$41724 ( \42101 , \42099 , \42100 );
not \U$41725 ( \42102 , \11665 );
and \U$41726 ( \42103 , RIae7a6f0_184, \42102 );
not \U$41727 ( \42104 , RIae7a6f0_184);
and \U$41728 ( \42105 , \42104 , \10043 );
or \U$41729 ( \42106 , \42103 , \42105 );
nand \U$41730 ( \42107 , \42106 , \9473 );
nand \U$41731 ( \42108 , \42101 , \42107 );
xor \U$41732 ( \42109 , \42098 , \42108 );
not \U$41733 ( \42110 , \42109 );
or \U$41734 ( \42111 , \42062 , \42110 );
nand \U$41735 ( \42112 , \42108 , \42098 );
nand \U$41736 ( \42113 , \42111 , \42112 );
not \U$41737 ( \42114 , \42113 );
not \U$41738 ( \42115 , \9744 );
not \U$41739 ( \42116 , \41550 );
or \U$41740 ( \42117 , \42115 , \42116 );
nand \U$41741 ( \42118 , \42068 , \9728 );
nand \U$41742 ( \42119 , \42117 , \42118 );
xnor \U$41743 ( \42120 , \42003 , \42005 );
xor \U$41744 ( \42121 , \42119 , \42120 );
not \U$41745 ( \42122 , \42014 );
not \U$41746 ( \42123 , \42122 );
not \U$41747 ( \42124 , \9526 );
and \U$41748 ( \42125 , \42123 , \42124 );
and \U$41749 ( \42126 , \42086 , \9549 );
nor \U$41750 ( \42127 , \42125 , \42126 );
or \U$41751 ( \42128 , \42121 , \42127 );
not \U$41752 ( \42129 , \42119 );
or \U$41753 ( \42130 , \42129 , \42120 );
nand \U$41754 ( \42131 , \42128 , \42130 );
not \U$41755 ( \42132 , \42131 );
not \U$41756 ( \42133 , \42017 );
not \U$41757 ( \42134 , \42026 );
not \U$41758 ( \42135 , \42134 );
and \U$41759 ( \42136 , \42133 , \42135 );
and \U$41760 ( \42137 , \42017 , \42134 );
nor \U$41761 ( \42138 , \42136 , \42137 );
not \U$41762 ( \42139 , \42138 );
or \U$41763 ( \42140 , \42132 , \42139 );
or \U$41764 ( \42141 , \42138 , \42131 );
nand \U$41765 ( \42142 , \42140 , \42141 );
not \U$41766 ( \42143 , \42142 );
or \U$41767 ( \42144 , \42114 , \42143 );
not \U$41768 ( \42145 , \42138 );
nand \U$41769 ( \42146 , \42145 , \42131 );
nand \U$41770 ( \42147 , \42144 , \42146 );
not \U$41771 ( \42148 , \42147 );
or \U$41772 ( \42149 , \42050 , \42148 );
or \U$41773 ( \42150 , \42147 , \42049 );
nand \U$41774 ( \42151 , \42149 , \42150 );
not \U$41775 ( \42152 , \42151 );
or \U$41776 ( \42153 , \42048 , \42152 );
not \U$41777 ( \42154 , \42046 );
or \U$41778 ( \42155 , \42154 , \42151 );
nand \U$41779 ( \42156 , \42153 , \42155 );
buf \U$41780 ( \42157 , \42142 );
not \U$41781 ( \42158 , \42113 );
and \U$41782 ( \42159 , \42157 , \42158 );
not \U$41783 ( \42160 , \42157 );
and \U$41784 ( \42161 , \42160 , \42113 );
nor \U$41785 ( \42162 , \42159 , \42161 );
not \U$41786 ( \42163 , \42162 );
not \U$41787 ( \42164 , \42163 );
and \U$41788 ( \42165 , \42121 , \42127 );
not \U$41789 ( \42166 , \42121 );
not \U$41790 ( \42167 , \42127 );
and \U$41791 ( \42168 , \42166 , \42167 );
nor \U$41792 ( \42169 , \42165 , \42168 );
not \U$41793 ( \42170 , \42169 );
not \U$41794 ( \42171 , RIae7aab0_192);
not \U$41795 ( \42172 , \41987 );
or \U$41796 ( \42173 , \42171 , \42172 );
not \U$41797 ( \42174 , \11326 );
not \U$41798 ( \42175 , \10007 );
or \U$41799 ( \42176 , \42174 , \42175 );
or \U$41800 ( \42177 , \10007 , \11326 );
nand \U$41801 ( \42178 , \42176 , \42177 );
nand \U$41802 ( \42179 , \42178 , \14667 );
nand \U$41803 ( \42180 , \42173 , \42179 );
not \U$41804 ( \42181 , \42180 );
nand \U$41805 ( \42182 , \9537 , \9725 );
and \U$41806 ( \42183 , \12857 , \42182 );
nor \U$41807 ( \42184 , \42183 , \15731 );
not \U$41808 ( \42185 , \9744 );
not \U$41809 ( \42186 , \42075 );
or \U$41810 ( \42187 , \42185 , \42186 );
and \U$41811 ( \42188 , RIae7a060_170, \12857 );
not \U$41812 ( \42189 , RIae7a060_170);
and \U$41813 ( \42190 , \42189 , \16890 );
nor \U$41814 ( \42191 , \42188 , \42190 );
nand \U$41815 ( \42192 , \42191 , \9728 );
nand \U$41816 ( \42193 , \42187 , \42192 );
and \U$41817 ( \42194 , \42184 , \42193 );
not \U$41818 ( \42195 , \9478 );
not \U$41819 ( \42196 , \42106 );
or \U$41820 ( \42197 , \42195 , \42196 );
not \U$41821 ( \42198 , \16101 );
not \U$41822 ( \42199 , \30081 );
or \U$41823 ( \42200 , \42198 , \42199 );
nand \U$41824 ( \42201 , \11240 , RIae7a6f0_184);
nand \U$41825 ( \42202 , \42200 , \42201 );
nand \U$41826 ( \42203 , \42202 , \9472 );
nand \U$41827 ( \42204 , \42197 , \42203 );
xor \U$41828 ( \42205 , \42194 , \42204 );
or \U$41829 ( \42206 , \42058 , \10276 );
not \U$41830 ( \42207 , \42059 );
not \U$41831 ( \42208 , \18088 );
not \U$41832 ( \42209 , \33415 );
or \U$41833 ( \42210 , \42208 , \42209 );
nand \U$41834 ( \42211 , \11589 , RIae7a8d0_188);
nand \U$41835 ( \42212 , \42210 , \42211 );
nand \U$41836 ( \42213 , \42207 , \42212 );
nand \U$41837 ( \42214 , \42206 , \42213 );
and \U$41838 ( \42215 , \42205 , \42214 );
and \U$41839 ( \42216 , \42194 , \42204 );
nor \U$41840 ( \42217 , \42215 , \42216 );
not \U$41841 ( \42218 , \42217 );
or \U$41842 ( \42219 , \42181 , \42218 );
or \U$41843 ( \42220 , \42217 , \42180 );
nand \U$41844 ( \42221 , \42219 , \42220 );
not \U$41845 ( \42222 , \42221 );
or \U$41846 ( \42223 , \42170 , \42222 );
not \U$41847 ( \42224 , \42217 );
nand \U$41848 ( \42225 , \42224 , \42180 );
nand \U$41849 ( \42226 , \42223 , \42225 );
xor \U$41850 ( \42227 , \41971 , \41981 );
xor \U$41851 ( \42228 , \42227 , \41991 );
xor \U$41852 ( \42229 , \42226 , \42228 );
not \U$41853 ( \42230 , \42229 );
or \U$41854 ( \42231 , \42164 , \42230 );
nand \U$41855 ( \42232 , \42226 , \42228 );
nand \U$41856 ( \42233 , \42231 , \42232 );
nor \U$41857 ( \42234 , \42156 , \42233 );
and \U$41858 ( \42235 , \42109 , \42061 );
not \U$41859 ( \42236 , \42109 );
not \U$41860 ( \42237 , \42061 );
and \U$41861 ( \42238 , \42236 , \42237 );
nor \U$41862 ( \42239 , \42235 , \42238 );
not \U$41863 ( \42240 , \42178 );
or \U$41864 ( \42241 , \42240 , \14666 );
and \U$41865 ( \42242 , RIae7aa38_191, \27672 );
not \U$41866 ( \42243 , RIae7aa38_191);
and \U$41867 ( \42244 , \42243 , \27671 );
nor \U$41868 ( \42245 , \42242 , \42244 );
or \U$41869 ( \42246 , \42245 , \18053 );
nand \U$41870 ( \42247 , \42241 , \42246 );
not \U$41871 ( \42248 , \42247 );
xor \U$41872 ( \42249 , \42079 , \42094 );
not \U$41873 ( \42250 , \42249 );
xor \U$41874 ( \42251 , \42184 , \42193 );
not \U$41875 ( \42252 , \29518 );
not \U$41876 ( \42253 , \42092 );
or \U$41877 ( \42254 , \42252 , \42253 );
and \U$41878 ( \42255 , RIae7a7e0_186, \16652 );
not \U$41879 ( \42256 , RIae7a7e0_186);
and \U$41880 ( \42257 , \42256 , \16651 );
nor \U$41881 ( \42258 , \42255 , \42257 );
nand \U$41882 ( \42259 , \42258 , \9549 );
nand \U$41883 ( \42260 , \42254 , \42259 );
xor \U$41884 ( \42261 , \42251 , \42260 );
not \U$41885 ( \42262 , \42261 );
not \U$41886 ( \42263 , \10275 );
not \U$41887 ( \42264 , \42212 );
or \U$41888 ( \42265 , \42263 , \42264 );
not \U$41889 ( \42266 , \11207 );
not \U$41890 ( \42267 , \16912 );
or \U$41891 ( \42268 , \42266 , \42267 );
or \U$41892 ( \42269 , \10043 , \18088 );
nand \U$41893 ( \42270 , \42268 , \42269 );
nand \U$41894 ( \42271 , \42270 , \11204 );
nand \U$41895 ( \42272 , \42265 , \42271 );
not \U$41896 ( \42273 , \42272 );
or \U$41897 ( \42274 , \42262 , \42273 );
nand \U$41898 ( \42275 , \42260 , \42251 );
nand \U$41899 ( \42276 , \42274 , \42275 );
not \U$41900 ( \42277 , \42276 );
not \U$41901 ( \42278 , \42277 );
or \U$41902 ( \42279 , \42250 , \42278 );
or \U$41903 ( \42280 , \42277 , \42249 );
nand \U$41904 ( \42281 , \42279 , \42280 );
not \U$41905 ( \42282 , \42281 );
or \U$41906 ( \42283 , \42248 , \42282 );
not \U$41907 ( \42284 , \42277 );
nand \U$41908 ( \42285 , \42284 , \42249 );
nand \U$41909 ( \42286 , \42283 , \42285 );
xor \U$41910 ( \42287 , \42239 , \42286 );
xor \U$41911 ( \42288 , \42221 , \42169 );
and \U$41912 ( \42289 , \42287 , \42288 );
and \U$41913 ( \42290 , \42239 , \42286 );
nor \U$41914 ( \42291 , \42289 , \42290 );
not \U$41915 ( \42292 , \42291 );
not \U$41916 ( \42293 , \42162 );
not \U$41917 ( \42294 , \42229 );
or \U$41918 ( \42295 , \42293 , \42294 );
or \U$41919 ( \42296 , \42229 , \42162 );
nand \U$41920 ( \42297 , \42295 , \42296 );
nand \U$41921 ( \42298 , \42292 , \42297 );
or \U$41922 ( \42299 , \42234 , \42298 );
nand \U$41923 ( \42300 , \42156 , \42233 );
nand \U$41924 ( \42301 , \42299 , \42300 );
not \U$41925 ( \42302 , \42301 );
not \U$41926 ( \42303 , \41421 );
and \U$41927 ( \42304 , \41459 , \42303 );
not \U$41928 ( \42305 , \41459 );
and \U$41929 ( \42306 , \42305 , \41421 );
nor \U$41930 ( \42307 , \42304 , \42306 );
not \U$41931 ( \42308 , \41994 );
not \U$41932 ( \42309 , \42042 );
or \U$41933 ( \42310 , \42308 , \42309 );
not \U$41934 ( \42311 , \42029 );
nand \U$41935 ( \42312 , \42311 , \42037 );
nand \U$41936 ( \42313 , \42310 , \42312 );
xor \U$41937 ( \42314 , \42307 , \42313 );
not \U$41938 ( \42315 , \41581 );
not \U$41939 ( \42316 , \41515 );
not \U$41940 ( \42317 , \42316 );
and \U$41941 ( \42318 , \42315 , \42317 );
and \U$41942 ( \42319 , \41581 , \42316 );
nor \U$41943 ( \42320 , \42318 , \42319 );
xnor \U$41944 ( \42321 , \42314 , \42320 );
not \U$41945 ( \42322 , \42049 );
nand \U$41946 ( \42323 , \42322 , \42147 );
not \U$41947 ( \42324 , \42323 );
not \U$41948 ( \42325 , \42154 );
or \U$41949 ( \42326 , \42324 , \42325 );
not \U$41950 ( \42327 , \42147 );
nand \U$41951 ( \42328 , \42327 , \42049 );
nand \U$41952 ( \42329 , \42326 , \42328 );
nand \U$41953 ( \42330 , \42321 , \42329 );
not \U$41954 ( \42331 , \42330 );
or \U$41955 ( \42332 , \42302 , \42331 );
or \U$41956 ( \42333 , \42321 , \42329 );
nand \U$41957 ( \42334 , \42332 , \42333 );
not \U$41958 ( \42335 , \41590 );
not \U$41959 ( \42336 , \41487 );
not \U$41960 ( \42337 , \41585 );
or \U$41961 ( \42338 , \42336 , \42337 );
or \U$41962 ( \42339 , \41585 , \41487 );
nand \U$41963 ( \42340 , \42338 , \42339 );
not \U$41964 ( \42341 , \42340 );
or \U$41965 ( \42342 , \42335 , \42341 );
or \U$41966 ( \42343 , \42340 , \41590 );
nand \U$41967 ( \42344 , \42342 , \42343 );
not \U$41968 ( \42345 , \42307 );
not \U$41969 ( \42346 , \42320 );
or \U$41970 ( \42347 , \42345 , \42346 );
nand \U$41971 ( \42348 , \42347 , \42313 );
or \U$41972 ( \42349 , \42307 , \42320 );
and \U$41973 ( \42350 , \42348 , \42349 );
nand \U$41974 ( \42351 , \42344 , \42350 );
nand \U$41975 ( \42352 , \42334 , \42351 );
not \U$41976 ( \42353 , \42291 );
nor \U$41977 ( \42354 , \42297 , \42353 );
nor \U$41978 ( \42355 , \42234 , \42354 );
or \U$41979 ( \42356 , \42245 , \14666 );
and \U$41980 ( \42357 , RIae7aa38_191, \40490 );
not \U$41981 ( \42358 , RIae7aa38_191);
and \U$41982 ( \42359 , \42358 , \10142 );
nor \U$41983 ( \42360 , \42357 , \42359 );
not \U$41984 ( \42361 , \14667 );
or \U$41985 ( \42362 , \42360 , \42361 );
nand \U$41986 ( \42363 , \42356 , \42362 );
not \U$41987 ( \42364 , \42202 );
or \U$41988 ( \42365 , \42364 , \36656 );
not \U$41989 ( \42366 , \16101 );
not \U$41990 ( \42367 , \11318 );
or \U$41991 ( \42368 , \42366 , \42367 );
or \U$41992 ( \42369 , \11318 , \27644 );
nand \U$41993 ( \42370 , \42368 , \42369 );
not \U$41994 ( \42371 , \42370 );
not \U$41995 ( \42372 , \9472 );
or \U$41996 ( \42373 , \42371 , \42372 );
nand \U$41997 ( \42374 , \42365 , \42373 );
not \U$41998 ( \42375 , \42374 );
not \U$41999 ( \42376 , \42375 );
not \U$42000 ( \42377 , \29518 );
not \U$42001 ( \42378 , \42258 );
or \U$42002 ( \42379 , \42377 , \42378 );
not \U$42003 ( \42380 , RIae7a7e0_186);
not \U$42004 ( \42381 , \18986 );
or \U$42005 ( \42382 , \42380 , \42381 );
or \U$42006 ( \42383 , \12750 , RIae7a7e0_186);
nand \U$42007 ( \42384 , \42382 , \42383 );
nand \U$42008 ( \42385 , \42384 , \9549 );
nand \U$42009 ( \42386 , \42379 , \42385 );
and \U$42010 ( \42387 , \12857 , \9744 );
nor \U$42011 ( \42388 , \42386 , \42387 );
not \U$42012 ( \42389 , \42388 );
not \U$42013 ( \42390 , \42389 );
not \U$42014 ( \42391 , \9470 );
not \U$42015 ( \42392 , \42370 );
or \U$42016 ( \42393 , \42391 , \42392 );
and \U$42017 ( \42394 , RIae7a6f0_184, \39806 );
not \U$42018 ( \42395 , RIae7a6f0_184);
and \U$42019 ( \42396 , \42395 , \41920 );
or \U$42020 ( \42397 , \42394 , \42396 );
nand \U$42021 ( \42398 , \42397 , \9472 );
nand \U$42022 ( \42399 , \42393 , \42398 );
not \U$42023 ( \42400 , \42399 );
or \U$42024 ( \42401 , \42390 , \42400 );
nand \U$42025 ( \42402 , \42386 , \42387 );
nand \U$42026 ( \42403 , \42401 , \42402 );
not \U$42027 ( \42404 , \42403 );
or \U$42028 ( \42405 , \42376 , \42404 );
or \U$42029 ( \42406 , \42403 , \42375 );
nand \U$42030 ( \42407 , \42405 , \42406 );
xor \U$42031 ( \42408 , \42363 , \42407 );
not \U$42032 ( \42409 , \42408 );
not \U$42033 ( \42410 , \14667 );
and \U$42034 ( \42411 , \33415 , RIae7aa38_191);
not \U$42035 ( \42412 , \33415 );
and \U$42036 ( \42413 , \42412 , \11326 );
nor \U$42037 ( \42414 , \42411 , \42413 );
not \U$42038 ( \42415 , \42414 );
or \U$42039 ( \42416 , \42410 , \42415 );
not \U$42040 ( \42417 , \42360 );
nand \U$42041 ( \42418 , \42417 , RIae7aab0_192);
nand \U$42042 ( \42419 , \42416 , \42418 );
not \U$42043 ( \42420 , \42419 );
not \U$42044 ( \42421 , \10275 );
not \U$42045 ( \42422 , \42270 );
or \U$42046 ( \42423 , \42421 , \42422 );
not \U$42047 ( \42424 , RIae7a8d0_188);
not \U$42048 ( \42425 , \11240 );
or \U$42049 ( \42426 , \42424 , \42425 );
or \U$42050 ( \42427 , \10194 , RIae7a8d0_188);
nand \U$42051 ( \42428 , \42426 , \42427 );
nand \U$42052 ( \42429 , \42428 , \11204 );
nand \U$42053 ( \42430 , \42423 , \42429 );
nand \U$42054 ( \42431 , \16101 , \9522 );
and \U$42055 ( \42432 , \12857 , \42431 );
nor \U$42056 ( \42433 , \42432 , \13415 );
not \U$42057 ( \42434 , \29518 );
not \U$42058 ( \42435 , \42384 );
or \U$42059 ( \42436 , \42434 , \42435 );
xor \U$42060 ( \42437 , \12857 , RIae7a7e0_186);
nand \U$42061 ( \42438 , \42437 , \9549 );
nand \U$42062 ( \42439 , \42436 , \42438 );
and \U$42063 ( \42440 , \42433 , \42439 );
nor \U$42064 ( \42441 , \42430 , \42440 );
buf \U$42065 ( \42442 , \42441 );
or \U$42066 ( \42443 , \42420 , \42442 );
nand \U$42067 ( \42444 , \42430 , \42440 );
nand \U$42068 ( \42445 , \42443 , \42444 );
xor \U$42069 ( \42446 , \42272 , \42261 );
nor \U$42070 ( \42447 , \42445 , \42446 );
not \U$42071 ( \42448 , \42447 );
not \U$42072 ( \42449 , \42448 );
or \U$42073 ( \42450 , \42409 , \42449 );
nand \U$42074 ( \42451 , \42445 , \42446 );
nand \U$42075 ( \42452 , \42450 , \42451 );
not \U$42076 ( \42453 , \42452 );
xnor \U$42077 ( \42454 , \42205 , \42214 );
nand \U$42078 ( \42455 , \42407 , \42363 );
nand \U$42079 ( \42456 , \42403 , \42374 );
and \U$42080 ( \42457 , \42455 , \42456 );
xor \U$42081 ( \42458 , \42454 , \42457 );
not \U$42082 ( \42459 , \42247 );
and \U$42083 ( \42460 , \42281 , \42459 );
not \U$42084 ( \42461 , \42281 );
and \U$42085 ( \42462 , \42461 , \42247 );
nor \U$42086 ( \42463 , \42460 , \42462 );
xor \U$42087 ( \42464 , \42458 , \42463 );
nand \U$42088 ( \42465 , \42453 , \42464 );
not \U$42089 ( \42466 , \42465 );
not \U$42090 ( \42467 , \42447 );
nand \U$42091 ( \42468 , \42467 , \42451 );
xor \U$42092 ( \42469 , \42468 , \42408 );
xor \U$42093 ( \42470 , \42433 , \42439 );
not \U$42094 ( \42471 , \9470 );
not \U$42095 ( \42472 , \42397 );
or \U$42096 ( \42473 , \42471 , \42472 );
and \U$42097 ( \42474 , RIae7a6f0_184, \16651 );
not \U$42098 ( \42475 , RIae7a6f0_184);
and \U$42099 ( \42476 , \42475 , \16652 );
or \U$42100 ( \42477 , \42474 , \42476 );
nand \U$42101 ( \42478 , \42477 , \9472 );
nand \U$42102 ( \42479 , \42473 , \42478 );
xor \U$42103 ( \42480 , \42470 , \42479 );
not \U$42104 ( \42481 , \11204 );
not \U$42105 ( \42482 , \11207 );
not \U$42106 ( \42483 , \10272 );
or \U$42107 ( \42484 , \42482 , \42483 );
or \U$42108 ( \42485 , \10272 , \18088 );
nand \U$42109 ( \42486 , \42484 , \42485 );
not \U$42110 ( \42487 , \42486 );
or \U$42111 ( \42488 , \42481 , \42487 );
not \U$42112 ( \42489 , \42428 );
or \U$42113 ( \42490 , \42489 , \10276 );
nand \U$42114 ( \42491 , \42488 , \42490 );
and \U$42115 ( \42492 , \42480 , \42491 );
and \U$42116 ( \42493 , \42470 , \42479 );
or \U$42117 ( \42494 , \42492 , \42493 );
not \U$42118 ( \42495 , \42388 );
nand \U$42119 ( \42496 , \42495 , \42402 );
xor \U$42120 ( \42497 , \42496 , \42399 );
not \U$42121 ( \42498 , \42497 );
or \U$42122 ( \42499 , \42494 , \42498 );
not \U$42123 ( \42500 , \42420 );
not \U$42124 ( \42501 , \42441 );
nand \U$42125 ( \42502 , \42501 , \42444 );
not \U$42126 ( \42503 , \42502 );
or \U$42127 ( \42504 , \42500 , \42503 );
or \U$42128 ( \42505 , \42502 , \42420 );
nand \U$42129 ( \42506 , \42504 , \42505 );
not \U$42130 ( \42507 , \42497 );
not \U$42131 ( \42508 , \42494 );
or \U$42132 ( \42509 , \42507 , \42508 );
or \U$42133 ( \42510 , \42494 , \42497 );
nand \U$42134 ( \42511 , \42509 , \42510 );
nand \U$42135 ( \42512 , \42506 , \42511 );
nand \U$42136 ( \42513 , \42499 , \42512 );
nand \U$42137 ( \42514 , \42469 , \42513 );
not \U$42138 ( \42515 , \42514 );
or \U$42139 ( \42516 , \42506 , \42511 );
nand \U$42140 ( \42517 , \42516 , \42512 );
not \U$42141 ( \42518 , \10275 );
not \U$42142 ( \42519 , \42486 );
or \U$42143 ( \42520 , \42518 , \42519 );
and \U$42144 ( \42521 , RIae7a8d0_188, \39806 );
not \U$42145 ( \42522 , RIae7a8d0_188);
not \U$42146 ( \42523 , \39806 );
and \U$42147 ( \42524 , \42522 , \42523 );
or \U$42148 ( \42525 , \42521 , \42524 );
nand \U$42149 ( \42526 , \42525 , \11204 );
nand \U$42150 ( \42527 , \42520 , \42526 );
not \U$42151 ( \42528 , \42527 );
not \U$42152 ( \42529 , \9470 );
not \U$42153 ( \42530 , \42477 );
or \U$42154 ( \42531 , \42529 , \42530 );
not \U$42155 ( \42532 , RIae7a6f0_184);
not \U$42156 ( \42533 , \18986 );
or \U$42157 ( \42534 , \42532 , \42533 );
or \U$42158 ( \42535 , \41907 , RIae7a6f0_184);
nand \U$42159 ( \42536 , \42534 , \42535 );
nand \U$42160 ( \42537 , \42536 , \9472 );
nand \U$42161 ( \42538 , \42531 , \42537 );
and \U$42162 ( \42539 , \12857 , \29518 );
xor \U$42163 ( \42540 , \42538 , \42539 );
not \U$42164 ( \42541 , \42540 );
or \U$42165 ( \42542 , \42528 , \42541 );
nand \U$42166 ( \42543 , \42538 , \42539 );
nand \U$42167 ( \42544 , \42542 , \42543 );
not \U$42168 ( \42545 , RIae7aab0_192);
not \U$42169 ( \42546 , \42414 );
or \U$42170 ( \42547 , \42545 , \42546 );
not \U$42171 ( \42548 , \14671 );
not \U$42172 ( \42549 , \10043 );
or \U$42173 ( \42550 , \42548 , \42549 );
or \U$42174 ( \42551 , \10043 , \14671 );
nand \U$42175 ( \42552 , \42550 , \42551 );
nand \U$42176 ( \42553 , \42552 , \14667 );
nand \U$42177 ( \42554 , \42547 , \42553 );
xor \U$42178 ( \42555 , \42544 , \42554 );
xor \U$42179 ( \42556 , \42470 , \42479 );
xor \U$42180 ( \42557 , \42556 , \42491 );
and \U$42181 ( \42558 , \42555 , \42557 );
and \U$42182 ( \42559 , \42544 , \42554 );
or \U$42183 ( \42560 , \42558 , \42559 );
or \U$42184 ( \42561 , \42517 , \42560 );
or \U$42185 ( \42562 , RIae7a858_187, RIae7a8d0_188);
nand \U$42186 ( \42563 , \42562 , \12857 );
nand \U$42187 ( \42564 , \42563 , \11668 );
not \U$42188 ( \42565 , \42564 );
not \U$42189 ( \42566 , \9470 );
not \U$42190 ( \42567 , \42536 );
or \U$42191 ( \42568 , \42566 , \42567 );
and \U$42192 ( \42569 , RIae7a6f0_184, \12857 );
not \U$42193 ( \42570 , RIae7a6f0_184);
and \U$42194 ( \42571 , \42570 , \14601 );
nor \U$42195 ( \42572 , \42569 , \42571 );
nand \U$42196 ( \42573 , \42572 , \9471 );
nand \U$42197 ( \42574 , \42568 , \42573 );
not \U$42198 ( \42575 , \42574 );
or \U$42199 ( \42576 , \42565 , \42575 );
or \U$42200 ( \42577 , \42574 , \42564 );
nand \U$42201 ( \42578 , \42576 , \42577 );
not \U$42202 ( \42579 , \10275 );
not \U$42203 ( \42580 , \42525 );
or \U$42204 ( \42581 , \42579 , \42580 );
and \U$42205 ( \42582 , \10844 , \11207 );
not \U$42206 ( \42583 , \10844 );
and \U$42207 ( \42584 , \42583 , RIae7a8d0_188);
nor \U$42208 ( \42585 , \42582 , \42584 );
nand \U$42209 ( \42586 , \42585 , \11204 );
nand \U$42210 ( \42587 , \42581 , \42586 );
xor \U$42211 ( \42588 , \42578 , \42587 );
not \U$42212 ( \42589 , RIae7aab0_192);
and \U$42213 ( \42590 , RIae7aa38_191, \10195 );
not \U$42214 ( \42591 , RIae7aa38_191);
and \U$42215 ( \42592 , \42591 , \10194 );
nor \U$42216 ( \42593 , \42590 , \42592 );
not \U$42217 ( \42594 , \42593 );
or \U$42218 ( \42595 , \42589 , \42594 );
not \U$42219 ( \42596 , \14671 );
not \U$42220 ( \42597 , \10272 );
or \U$42221 ( \42598 , \42596 , \42597 );
or \U$42222 ( \42599 , \10272 , \14671 );
nand \U$42223 ( \42600 , \42598 , \42599 );
nand \U$42224 ( \42601 , \42600 , \14667 );
nand \U$42225 ( \42602 , \42595 , \42601 );
and \U$42226 ( \42603 , \42588 , \42602 );
and \U$42227 ( \42604 , \42587 , \42578 );
nor \U$42228 ( \42605 , \42603 , \42604 );
not \U$42229 ( \42606 , \42605 );
xor \U$42230 ( \42607 , \42527 , \42540 );
not \U$42231 ( \42608 , RIae7aab0_192);
not \U$42232 ( \42609 , \42552 );
or \U$42233 ( \42610 , \42608 , \42609 );
nand \U$42234 ( \42611 , \42593 , \14667 );
nand \U$42235 ( \42612 , \42610 , \42611 );
not \U$42236 ( \42613 , \42612 );
not \U$42237 ( \42614 , \42564 );
nand \U$42238 ( \42615 , \42614 , \42574 );
not \U$42239 ( \42616 , \42615 );
and \U$42240 ( \42617 , \42613 , \42616 );
and \U$42241 ( \42618 , \42612 , \42615 );
nor \U$42242 ( \42619 , \42617 , \42618 );
and \U$42243 ( \42620 , \42607 , \42619 );
not \U$42244 ( \42621 , \42607 );
not \U$42245 ( \42622 , \42619 );
and \U$42246 ( \42623 , \42621 , \42622 );
nor \U$42247 ( \42624 , \42620 , \42623 );
not \U$42248 ( \42625 , \42624 );
or \U$42249 ( \42626 , \42606 , \42625 );
not \U$42250 ( \42627 , \42588 );
and \U$42251 ( \42628 , \42602 , \42627 );
not \U$42252 ( \42629 , \42602 );
and \U$42253 ( \42630 , \42629 , \42588 );
nor \U$42254 ( \42631 , \42628 , \42630 );
not \U$42255 ( \42632 , \10275 );
not \U$42256 ( \42633 , \42585 );
or \U$42257 ( \42634 , \42632 , \42633 );
not \U$42258 ( \42635 , RIae7a8d0_188);
not \U$42259 ( \42636 , \16006 );
or \U$42260 ( \42637 , \42635 , \42636 );
or \U$42261 ( \42638 , \16006 , RIae7a8d0_188);
nand \U$42262 ( \42639 , \42637 , \42638 );
nand \U$42263 ( \42640 , \42639 , \11204 );
nand \U$42264 ( \42641 , \42634 , \42640 );
nand \U$42265 ( \42642 , \12857 , \9470 );
not \U$42266 ( \42643 , \42642 );
and \U$42267 ( \42644 , \42641 , \42643 );
not \U$42268 ( \42645 , RIae7aab0_192);
not \U$42269 ( \42646 , \42600 );
or \U$42270 ( \42647 , \42645 , \42646 );
xor \U$42271 ( \42648 , RIae7aa38_191, \39806 );
or \U$42272 ( \42649 , \42648 , \42361 );
nand \U$42273 ( \42650 , \42647 , \42649 );
not \U$42274 ( \42651 , \42642 );
not \U$42275 ( \42652 , \42641 );
or \U$42276 ( \42653 , \42651 , \42652 );
or \U$42277 ( \42654 , \42641 , \42642 );
nand \U$42278 ( \42655 , \42653 , \42654 );
and \U$42279 ( \42656 , \42650 , \42655 );
nor \U$42280 ( \42657 , \42644 , \42656 );
nand \U$42281 ( \42658 , \42631 , \42657 );
not \U$42282 ( \42659 , RIae7a9c0_190);
nand \U$42283 ( \42660 , \16890 , \14671 );
not \U$42284 ( \42661 , \42660 );
or \U$42285 ( \42662 , \42659 , \42661 );
and \U$42286 ( \42663 , \12857 , RIae7aa38_191);
nor \U$42287 ( \42664 , \42663 , \11207 );
nand \U$42288 ( \42665 , \42662 , \42664 );
not \U$42289 ( \42666 , \42665 );
not \U$42290 ( \42667 , \10275 );
not \U$42291 ( \42668 , \42639 );
or \U$42292 ( \42669 , \42667 , \42668 );
not \U$42293 ( \42670 , \18088 );
not \U$42294 ( \42671 , \12857 );
or \U$42295 ( \42672 , \42670 , \42671 );
or \U$42296 ( \42673 , \12857 , \18088 );
nand \U$42297 ( \42674 , \42672 , \42673 );
nand \U$42298 ( \42675 , \42674 , \10280 );
nand \U$42299 ( \42676 , \42669 , \42675 );
not \U$42300 ( \42677 , \42676 );
or \U$42301 ( \42678 , \42666 , \42677 );
or \U$42302 ( \42679 , \42676 , \42665 );
nand \U$42303 ( \42680 , \42678 , \42679 );
not \U$42304 ( \42681 , \42680 );
not \U$42305 ( \42682 , \42681 );
not \U$42306 ( \42683 , \11326 );
not \U$42307 ( \42684 , \16651 );
or \U$42308 ( \42685 , \42683 , \42684 );
nand \U$42309 ( \42686 , \16164 , RIae7aa38_191);
nand \U$42310 ( \42687 , \42685 , \42686 );
nor \U$42311 ( \42688 , \42687 , \14666 );
or \U$42312 ( \42689 , \42688 , \14667 );
and \U$42313 ( \42690 , \12857 , \10276 );
not \U$42314 ( \42691 , \42660 );
nor \U$42315 ( \42692 , \42690 , \42691 );
not \U$42316 ( \42693 , \12857 );
not \U$42317 ( \42694 , \42688 );
or \U$42318 ( \42695 , \42693 , \42694 );
not \U$42319 ( \42696 , \41907 );
nand \U$42320 ( \42697 , \42695 , \42696 );
nand \U$42321 ( \42698 , \42689 , \42692 , \42697 );
not \U$42322 ( \42699 , \42698 );
or \U$42323 ( \42700 , \42682 , \42699 );
or \U$42324 ( \42701 , \42648 , \14666 );
or \U$42325 ( \42702 , \42687 , \42361 );
nand \U$42326 ( \42703 , \42701 , \42702 );
nand \U$42327 ( \42704 , \42700 , \42703 );
not \U$42328 ( \42705 , \42698 );
nand \U$42329 ( \42706 , \42705 , \42680 );
nand \U$42330 ( \42707 , \42704 , \42706 );
not \U$42331 ( \42708 , \42707 );
xor \U$42332 ( \42709 , \42650 , \42655 );
not \U$42333 ( \42710 , \42709 );
or \U$42334 ( \42711 , \42708 , \42710 );
not \U$42335 ( \42712 , \42665 );
nand \U$42336 ( \42713 , \42712 , \42676 );
nand \U$42337 ( \42714 , \42711 , \42713 );
or \U$42338 ( \42715 , \42707 , \42709 );
nand \U$42339 ( \42716 , \42658 , \42714 , \42715 );
or \U$42340 ( \42717 , \42657 , \42631 );
nand \U$42341 ( \42718 , \42716 , \42717 );
nand \U$42342 ( \42719 , \42626 , \42718 );
xor \U$42343 ( \42720 , \42544 , \42554 );
xor \U$42344 ( \42721 , \42720 , \42557 );
not \U$42345 ( \42722 , \42607 );
not \U$42346 ( \42723 , \42622 );
or \U$42347 ( \42724 , \42722 , \42723 );
not \U$42348 ( \42725 , \42615 );
nand \U$42349 ( \42726 , \42725 , \42612 );
nand \U$42350 ( \42727 , \42724 , \42726 );
nand \U$42351 ( \42728 , \42721 , \42727 );
or \U$42352 ( \42729 , \42605 , \42624 );
nand \U$42353 ( \42730 , \42719 , \42728 , \42729 );
or \U$42354 ( \42731 , \42721 , \42727 );
nand \U$42355 ( \42732 , \42561 , \42730 , \42731 );
nand \U$42356 ( \42733 , \42517 , \42560 );
nand \U$42357 ( \42734 , \42732 , \42733 );
not \U$42358 ( \42735 , \42734 );
or \U$42359 ( \42736 , \42515 , \42735 );
not \U$42360 ( \42737 , \42469 );
not \U$42361 ( \42738 , \42513 );
nand \U$42362 ( \42739 , \42737 , \42738 );
nand \U$42363 ( \42740 , \42736 , \42739 );
not \U$42364 ( \42741 , \42740 );
or \U$42365 ( \42742 , \42466 , \42741 );
not \U$42366 ( \42743 , \42464 );
nand \U$42367 ( \42744 , \42743 , \42452 );
nand \U$42368 ( \42745 , \42742 , \42744 );
not \U$42369 ( \42746 , \42745 );
xor \U$42370 ( \42747 , \42454 , \42457 );
and \U$42371 ( \42748 , \42747 , \42463 );
and \U$42372 ( \42749 , \42454 , \42457 );
or \U$42373 ( \42750 , \42748 , \42749 );
not \U$42374 ( \42751 , \42750 );
xor \U$42375 ( \42752 , \42239 , \42286 );
xor \U$42376 ( \42753 , \42752 , \42288 );
not \U$42377 ( \42754 , \42753 );
or \U$42378 ( \42755 , \42751 , \42754 );
or \U$42379 ( \42756 , \42753 , \42750 );
nand \U$42380 ( \42757 , \42755 , \42756 );
not \U$42381 ( \42758 , \42757 );
or \U$42382 ( \42759 , \42746 , \42758 );
not \U$42383 ( \42760 , \42750 );
nand \U$42384 ( \42761 , \42760 , \42753 );
nand \U$42385 ( \42762 , \42759 , \42761 );
nand \U$42386 ( \42763 , \42351 , \42355 , \42330 , \42762 );
or \U$42387 ( \42764 , \42344 , \42350 );
nand \U$42388 ( \42765 , \42352 , \42763 , \42764 );
not \U$42389 ( \42766 , \41594 );
not \U$42390 ( \42767 , \41486 );
nand \U$42391 ( \42768 , \42766 , \42767 );
and \U$42392 ( \42769 , \41600 , \42768 );
nand \U$42393 ( \42770 , \42765 , \41969 , \41768 , \42769 );
or \U$42394 ( \42771 , \41961 , \41968 );
nand \U$42395 ( \42772 , \41970 , \42770 , \42771 );
not \U$42396 ( \42773 , \41775 );
not \U$42397 ( \42774 , \41831 );
or \U$42398 ( \42775 , \42773 , \42774 );
not \U$42399 ( \42776 , \41824 );
nand \U$42400 ( \42777 , \42776 , \41830 );
nand \U$42401 ( \42778 , \42775 , \42777 );
not \U$42402 ( \42779 , \42778 );
not \U$42403 ( \42780 , \10667 );
not \U$42404 ( \42781 , \41859 );
or \U$42405 ( \42782 , \42780 , \42781 );
and \U$42406 ( \42783 , \10658 , \11260 );
not \U$42407 ( \42784 , \10658 );
and \U$42408 ( \42785 , \42784 , \10007 );
nor \U$42409 ( \42786 , \42783 , \42785 );
nand \U$42410 ( \42787 , \42786 , \9776 );
nand \U$42411 ( \42788 , \42782 , \42787 );
not \U$42412 ( \42789 , \42788 );
not \U$42413 ( \42790 , \9473 );
not \U$42414 ( \42791 , \41873 );
or \U$42415 ( \42792 , \42790 , \42791 );
and \U$42416 ( \42793 , \10465 , RIae7a6f0_184);
not \U$42417 ( \42794 , \10465 );
and \U$42418 ( \42795 , \42794 , \16101 );
nor \U$42419 ( \42796 , \42793 , \42795 );
nand \U$42420 ( \42797 , \42796 , \9478 );
nand \U$42421 ( \42798 , \42792 , \42797 );
not \U$42422 ( \42799 , \42798 );
not \U$42423 ( \42800 , \42799 );
or \U$42424 ( \42801 , \42789 , \42800 );
or \U$42425 ( \42802 , \42799 , \42788 );
nand \U$42426 ( \42803 , \42801 , \42802 );
not \U$42427 ( \42804 , \11205 );
not \U$42428 ( \42805 , \41885 );
or \U$42429 ( \42806 , \42804 , \42805 );
and \U$42430 ( \42807 , RIae7a8d0_188, \9412 );
not \U$42431 ( \42808 , RIae7a8d0_188);
and \U$42432 ( \42809 , \42808 , \11198 );
or \U$42433 ( \42810 , \42807 , \42809 );
nand \U$42434 ( \42811 , \42810 , \10275 );
nand \U$42435 ( \42812 , \42806 , \42811 );
xor \U$42436 ( \42813 , \42803 , \42812 );
not \U$42437 ( \42814 , \41889 );
not \U$42438 ( \42815 , \41939 );
or \U$42439 ( \42816 , \42814 , \42815 );
nand \U$42440 ( \42817 , \41938 , \41932 );
nand \U$42441 ( \42818 , \42816 , \42817 );
nand \U$42442 ( \42819 , \41931 , \41900 );
not \U$42443 ( \42820 , \41927 );
nand \U$42444 ( \42821 , \42820 , \41917 );
and \U$42445 ( \42822 , \42819 , \42821 );
not \U$42446 ( \42823 , \42822 );
and \U$42447 ( \42824 , \41905 , \41916 );
not \U$42448 ( \42825 , \16358 );
not \U$42449 ( \42826 , \10633 );
not \U$42450 ( \42827 , \10043 );
or \U$42451 ( \42828 , \42826 , \42827 );
or \U$42452 ( \42829 , \11665 , \10633 );
nand \U$42453 ( \42830 , \42828 , \42829 );
not \U$42454 ( \42831 , \42830 );
or \U$42455 ( \42832 , \42825 , \42831 );
nand \U$42456 ( \42833 , \41896 , \10637 );
nand \U$42457 ( \42834 , \42832 , \42833 );
xor \U$42458 ( \42835 , \42824 , \42834 );
not \U$42459 ( \42836 , \10695 );
not \U$42460 ( \42837 , \41797 );
or \U$42461 ( \42838 , \42836 , \42837 );
and \U$42462 ( \42839 , RIae7a498_179, \10149 );
not \U$42463 ( \42840 , RIae7a498_179);
and \U$42464 ( \42841 , \42840 , \10142 );
or \U$42465 ( \42842 , \42839 , \42841 );
nand \U$42466 ( \42843 , \42842 , \10676 );
nand \U$42467 ( \42844 , \42838 , \42843 );
xor \U$42468 ( \42845 , \42835 , \42844 );
not \U$42469 ( \42846 , \42845 );
or \U$42470 ( \42847 , \42823 , \42846 );
or \U$42471 ( \42848 , \42845 , \42822 );
nand \U$42472 ( \42849 , \42847 , \42848 );
not \U$42473 ( \42850 , \16383 );
not \U$42474 ( \42851 , \41782 );
or \U$42475 ( \42852 , \42850 , \42851 );
and \U$42476 ( \42853 , RIae7aa38_191, \9455 );
not \U$42477 ( \42854 , RIae7aa38_191);
and \U$42478 ( \42855 , \42854 , \21948 );
nor \U$42479 ( \42856 , \42853 , \42855 );
nand \U$42480 ( \42857 , \42856 , RIae7aab0_192);
nand \U$42481 ( \42858 , \42852 , \42857 );
xor \U$42482 ( \42859 , \42849 , \42858 );
xor \U$42483 ( \42860 , \42818 , \42859 );
xor \U$42484 ( \42861 , \42813 , \42860 );
not \U$42485 ( \42862 , \42861 );
and \U$42486 ( \42863 , \12857 , \9813 );
not \U$42487 ( \42864 , \9699 );
and \U$42488 ( \42865 , RIae7a240_174, \16652 );
not \U$42489 ( \42866 , RIae7a240_174);
and \U$42490 ( \42867 , \42866 , \28243 );
nor \U$42491 ( \42868 , \42865 , \42867 );
not \U$42492 ( \42869 , \42868 );
or \U$42493 ( \42870 , \42864 , \42869 );
nand \U$42494 ( \42871 , \41911 , \9687 );
nand \U$42495 ( \42872 , \42870 , \42871 );
xor \U$42496 ( \42873 , \42863 , \42872 );
not \U$42497 ( \42874 , \9621 );
and \U$42498 ( \42875 , RIae7a3a8_177, \32808 );
not \U$42499 ( \42876 , RIae7a3a8_177);
and \U$42500 ( \42877 , \42876 , \11318 );
or \U$42501 ( \42878 , \42875 , \42877 );
not \U$42502 ( \42879 , \42878 );
or \U$42503 ( \42880 , \42874 , \42879 );
nand \U$42504 ( \42881 , \41924 , \9643 );
nand \U$42505 ( \42882 , \42880 , \42881 );
xnor \U$42506 ( \42883 , \42873 , \42882 );
not \U$42507 ( \42884 , \42883 );
not \U$42508 ( \42885 , \9728 );
not \U$42509 ( \42886 , \41853 );
or \U$42510 ( \42887 , \42885 , \42886 );
and \U$42511 ( \42888 , RIae7a060_170, \13544 );
not \U$42512 ( \42889 , RIae7a060_170);
and \U$42513 ( \42890 , \42889 , \10171 );
nor \U$42514 ( \42891 , \42888 , \42890 );
nand \U$42515 ( \42892 , \42891 , \9745 );
nand \U$42516 ( \42893 , \42887 , \42892 );
not \U$42517 ( \42894 , \42893 );
or \U$42518 ( \42895 , \42884 , \42894 );
or \U$42519 ( \42896 , \42893 , \42883 );
nand \U$42520 ( \42897 , \42895 , \42896 );
not \U$42521 ( \42898 , \42897 );
not \U$42522 ( \42899 , \10519 );
and \U$42523 ( \42900 , RIae7a7e0_186, \10084 );
not \U$42524 ( \42901 , RIae7a7e0_186);
and \U$42525 ( \42902 , \42901 , \21106 );
or \U$42526 ( \42903 , \42900 , \42902 );
not \U$42527 ( \42904 , \42903 );
or \U$42528 ( \42905 , \42899 , \42904 );
nand \U$42529 ( \42906 , \41807 , \11439 );
nand \U$42530 ( \42907 , \42905 , \42906 );
not \U$42531 ( \42908 , \42907 );
not \U$42532 ( \42909 , \42908 );
and \U$42533 ( \42910 , \42898 , \42909 );
and \U$42534 ( \42911 , \42897 , \42908 );
nor \U$42535 ( \42912 , \42910 , \42911 );
not \U$42536 ( \42913 , \42912 );
not \U$42537 ( \42914 , \42913 );
and \U$42538 ( \42915 , \41802 , \41811 );
and \U$42539 ( \42916 , \41791 , \41801 );
nor \U$42540 ( \42917 , \42915 , \42916 );
not \U$42541 ( \42918 , \42917 );
not \U$42542 ( \42919 , \41877 );
not \U$42543 ( \42920 , \41864 );
or \U$42544 ( \42921 , \42919 , \42920 );
nand \U$42545 ( \42922 , \42921 , \41865 );
not \U$42546 ( \42923 , \42922 );
or \U$42547 ( \42924 , \42918 , \42923 );
or \U$42548 ( \42925 , \42922 , \42917 );
nand \U$42549 ( \42926 , \42924 , \42925 );
not \U$42550 ( \42927 , \42926 );
not \U$42551 ( \42928 , \42927 );
or \U$42552 ( \42929 , \42914 , \42928 );
nand \U$42553 ( \42930 , \42926 , \42912 );
nand \U$42554 ( \42931 , \42929 , \42930 );
not \U$42555 ( \42932 , \42931 );
not \U$42556 ( \42933 , \41823 );
not \U$42557 ( \42934 , \41786 );
nand \U$42558 ( \42935 , \42934 , \41816 );
not \U$42559 ( \42936 , \42935 );
or \U$42560 ( \42937 , \42933 , \42936 );
not \U$42561 ( \42938 , \41816 );
nand \U$42562 ( \42939 , \42938 , \41786 );
nand \U$42563 ( \42940 , \42937 , \42939 );
not \U$42564 ( \42941 , \42940 );
not \U$42565 ( \42942 , \42941 );
and \U$42566 ( \42943 , \42932 , \42942 );
and \U$42567 ( \42944 , \42931 , \42941 );
nor \U$42568 ( \42945 , \42943 , \42944 );
not \U$42569 ( \42946 , \42945 );
not \U$42570 ( \42947 , \41847 );
not \U$42571 ( \42948 , \41948 );
or \U$42572 ( \42949 , \42947 , \42948 );
nand \U$42573 ( \42950 , \41943 , \41879 );
nand \U$42574 ( \42951 , \42949 , \42950 );
not \U$42575 ( \42952 , \42951 );
or \U$42576 ( \42953 , \42946 , \42952 );
or \U$42577 ( \42954 , \42951 , \42945 );
nand \U$42578 ( \42955 , \42953 , \42954 );
not \U$42579 ( \42956 , \42955 );
not \U$42580 ( \42957 , \42956 );
or \U$42581 ( \42958 , \42862 , \42957 );
not \U$42582 ( \42959 , \42861 );
nand \U$42583 ( \42960 , \42959 , \42955 );
nand \U$42584 ( \42961 , \42958 , \42960 );
not \U$42585 ( \42962 , \42961 );
or \U$42586 ( \42963 , \42779 , \42962 );
nand \U$42587 ( \42964 , \42955 , \42861 );
nand \U$42588 ( \42965 , \42963 , \42964 );
not \U$42589 ( \42966 , \42965 );
not \U$42590 ( \42967 , \42913 );
not \U$42591 ( \42968 , \42926 );
or \U$42592 ( \42969 , \42967 , \42968 );
not \U$42593 ( \42970 , \42917 );
nand \U$42594 ( \42971 , \42970 , \42922 );
nand \U$42595 ( \42972 , \42969 , \42971 );
not \U$42596 ( \42973 , \10675 );
not \U$42597 ( \42974 , RIae7a498_179);
not \U$42598 ( \42975 , \27672 );
or \U$42599 ( \42976 , \42974 , \42975 );
nand \U$42600 ( \42977 , \10743 , \10625 );
nand \U$42601 ( \42978 , \42976 , \42977 );
not \U$42602 ( \42979 , \42978 );
or \U$42603 ( \42980 , \42973 , \42979 );
nand \U$42604 ( \42981 , \42842 , \10695 );
nand \U$42605 ( \42982 , \42980 , \42981 );
not \U$42606 ( \42983 , \10542 );
and \U$42607 ( \42984 , RIae7a060_170, \11562 );
not \U$42608 ( \42985 , RIae7a060_170);
and \U$42609 ( \42986 , \42985 , \10072 );
or \U$42610 ( \42987 , \42984 , \42986 );
not \U$42611 ( \42988 , \42987 );
or \U$42612 ( \42989 , \42983 , \42988 );
nand \U$42613 ( \42990 , \42891 , \9728 );
nand \U$42614 ( \42991 , \42989 , \42990 );
xor \U$42615 ( \42992 , \42982 , \42991 );
not \U$42616 ( \42993 , \9776 );
not \U$42617 ( \42994 , \10672 );
not \U$42618 ( \42995 , \9868 );
or \U$42619 ( \42996 , \42994 , \42995 );
nand \U$42620 ( \42997 , \10750 , RIae7a150_172);
nand \U$42621 ( \42998 , \42996 , \42997 );
not \U$42622 ( \42999 , \42998 );
or \U$42623 ( \43000 , \42993 , \42999 );
nand \U$42624 ( \43001 , \42786 , \9758 );
nand \U$42625 ( \43002 , \43000 , \43001 );
xor \U$42626 ( \43003 , \42992 , \43002 );
not \U$42627 ( \43004 , \43003 );
not \U$42628 ( \43005 , \43004 );
not \U$42629 ( \43006 , \42812 );
not \U$42630 ( \43007 , \42803 );
or \U$42631 ( \43008 , \43006 , \43007 );
not \U$42632 ( \43009 , \42799 );
nand \U$42633 ( \43010 , \43009 , \42788 );
nand \U$42634 ( \43011 , \43008 , \43010 );
not \U$42635 ( \43012 , \42907 );
not \U$42636 ( \43013 , \42897 );
or \U$42637 ( \43014 , \43012 , \43013 );
not \U$42638 ( \43015 , \42883 );
nand \U$42639 ( \43016 , \43015 , \42893 );
nand \U$42640 ( \43017 , \43014 , \43016 );
xor \U$42641 ( \43018 , \43011 , \43017 );
not \U$42642 ( \43019 , \43018 );
or \U$42643 ( \43020 , \43005 , \43019 );
or \U$42644 ( \43021 , \43018 , \43004 );
nand \U$42645 ( \43022 , \43020 , \43021 );
xor \U$42646 ( \43023 , \42972 , \43022 );
or \U$42647 ( \43024 , \42859 , \42818 );
and \U$42648 ( \43025 , \43024 , \42813 );
and \U$42649 ( \43026 , \42818 , \42859 );
nor \U$42650 ( \43027 , \43025 , \43026 );
xor \U$42651 ( \43028 , \43023 , \43027 );
not \U$42652 ( \43029 , \43028 );
not \U$42653 ( \43030 , \42858 );
not \U$42654 ( \43031 , \42849 );
or \U$42655 ( \43032 , \43030 , \43031 );
not \U$42656 ( \43033 , \42822 );
nand \U$42657 ( \43034 , \43033 , \42845 );
nand \U$42658 ( \43035 , \43032 , \43034 );
not \U$42659 ( \43036 , \43035 );
and \U$42660 ( \43037 , RIae7a2b8_175, \18989 );
not \U$42661 ( \43038 , RIae7a2b8_175);
and \U$42662 ( \43039 , \43038 , \16006 );
or \U$42663 ( \43040 , \43037 , \43039 );
or \U$42664 ( \43041 , \43040 , \9786 );
xnor \U$42665 ( \43042 , \12857 , RIae7a2b8_175);
not \U$42666 ( \43043 , \9791 );
or \U$42667 ( \43044 , \43042 , \43043 );
nand \U$42668 ( \43045 , \43041 , \43044 );
not \U$42669 ( \43046 , \43045 );
not \U$42670 ( \43047 , \23809 );
or \U$42671 ( \43048 , RIae7a1c8_173, RIae7a240_174);
nand \U$42672 ( \43049 , \43048 , \12857 );
nand \U$42673 ( \43050 , \43047 , \43049 );
not \U$42674 ( \43051 , \43050 );
and \U$42675 ( \43052 , \43046 , \43051 );
and \U$42676 ( \43053 , \43045 , \43050 );
nor \U$42677 ( \43054 , \43052 , \43053 );
not \U$42678 ( \43055 , \9699 );
and \U$42679 ( \43056 , RIae7a240_174, \39806 );
not \U$42680 ( \43057 , RIae7a240_174);
and \U$42681 ( \43058 , \43057 , \42523 );
or \U$42682 ( \43059 , \43056 , \43058 );
not \U$42683 ( \43060 , \43059 );
or \U$42684 ( \43061 , \43055 , \43060 );
nand \U$42685 ( \43062 , \42868 , \9687 );
nand \U$42686 ( \43063 , \43061 , \43062 );
xnor \U$42687 ( \43064 , \43054 , \43063 );
not \U$42688 ( \43065 , \10631 );
not \U$42689 ( \43066 , RIae7a510_180);
not \U$42690 ( \43067 , \10337 );
or \U$42691 ( \43068 , \43066 , \43067 );
or \U$42692 ( \43069 , \16922 , RIae7a510_180);
nand \U$42693 ( \43070 , \43068 , \43069 );
not \U$42694 ( \43071 , \43070 );
or \U$42695 ( \43072 , \43065 , \43071 );
nand \U$42696 ( \43073 , \11400 , \42830 );
nand \U$42697 ( \43074 , \43072 , \43073 );
xor \U$42698 ( \43075 , \43064 , \43074 );
not \U$42699 ( \43076 , RIae7aab0_192);
not \U$42700 ( \43077 , \14671 );
not \U$42701 ( \43078 , \14110 );
or \U$42702 ( \43079 , \43077 , \43078 );
nand \U$42703 ( \43080 , \38489 , RIae7aa38_191);
nand \U$42704 ( \43081 , \43079 , \43080 );
not \U$42705 ( \43082 , \43081 );
or \U$42706 ( \43083 , \43076 , \43082 );
nand \U$42707 ( \43084 , \42856 , \14667 );
nand \U$42708 ( \43085 , \43083 , \43084 );
xor \U$42709 ( \43086 , \43075 , \43085 );
not \U$42710 ( \43087 , \10275 );
and \U$42711 ( \43088 , RIae7a8d0_188, \9398 );
not \U$42712 ( \43089 , RIae7a8d0_188);
and \U$42713 ( \43090 , \43089 , \10936 );
or \U$42714 ( \43091 , \43088 , \43090 );
not \U$42715 ( \43092 , \43091 );
or \U$42716 ( \43093 , \43087 , \43092 );
nand \U$42717 ( \43094 , \42810 , \17847 );
nand \U$42718 ( \43095 , \43093 , \43094 );
xnor \U$42719 ( \43096 , \43086 , \43095 );
nand \U$42720 ( \43097 , \43036 , \43096 );
not \U$42721 ( \43098 , \43096 );
nand \U$42722 ( \43099 , \43098 , \43035 );
nand \U$42723 ( \43100 , \43097 , \43099 );
xor \U$42724 ( \43101 , \42824 , \42834 );
and \U$42725 ( \43102 , \43101 , \42844 );
and \U$42726 ( \43103 , \42824 , \42834 );
or \U$42727 ( \43104 , \43102 , \43103 );
not \U$42728 ( \43105 , \10519 );
not \U$42729 ( \43106 , RIae7a7e0_186);
not \U$42730 ( \43107 , \40195 );
or \U$42731 ( \43108 , \43106 , \43107 );
or \U$42732 ( \43109 , \40198 , RIae7a7e0_186);
nand \U$42733 ( \43110 , \43108 , \43109 );
not \U$42734 ( \43111 , \43110 );
or \U$42735 ( \43112 , \43105 , \43111 );
nand \U$42736 ( \43113 , \42903 , \9549 );
nand \U$42737 ( \43114 , \43112 , \43113 );
not \U$42738 ( \43115 , \43114 );
not \U$42739 ( \43116 , \9621 );
and \U$42740 ( \43117 , RIae7a3a8_177, \11576 );
not \U$42741 ( \43118 , RIae7a3a8_177);
and \U$42742 ( \43119 , \43118 , \11240 );
nor \U$42743 ( \43120 , \43117 , \43119 );
not \U$42744 ( \43121 , \43120 );
or \U$42745 ( \43122 , \43116 , \43121 );
nand \U$42746 ( \43123 , \42878 , \9643 );
nand \U$42747 ( \43124 , \43122 , \43123 );
not \U$42748 ( \43125 , \43124 );
not \U$42749 ( \43126 , \43125 );
not \U$42750 ( \43127 , \42882 );
not \U$42751 ( \43128 , \42873 );
or \U$42752 ( \43129 , \43127 , \43128 );
nand \U$42753 ( \43130 , \42872 , \42863 );
nand \U$42754 ( \43131 , \43129 , \43130 );
not \U$42755 ( \43132 , \43131 );
or \U$42756 ( \43133 , \43126 , \43132 );
or \U$42757 ( \43134 , \43131 , \43125 );
nand \U$42758 ( \43135 , \43133 , \43134 );
not \U$42759 ( \43136 , \43135 );
and \U$42760 ( \43137 , \43115 , \43136 );
and \U$42761 ( \43138 , \43114 , \43135 );
nor \U$42762 ( \43139 , \43137 , \43138 );
xor \U$42763 ( \43140 , \43104 , \43139 );
not \U$42764 ( \43141 , \9478 );
xor \U$42765 ( \43142 , RIae7a6f0_184, \14148 );
not \U$42766 ( \43143 , \43142 );
or \U$42767 ( \43144 , \43141 , \43143 );
not \U$42768 ( \43145 , \42796 );
or \U$42769 ( \43146 , \43145 , \35746 );
nand \U$42770 ( \43147 , \43144 , \43146 );
and \U$42771 ( \43148 , \43140 , \43147 );
not \U$42772 ( \43149 , \43140 );
not \U$42773 ( \43150 , \43147 );
and \U$42774 ( \43151 , \43149 , \43150 );
nor \U$42775 ( \43152 , \43148 , \43151 );
not \U$42776 ( \43153 , \43152 );
and \U$42777 ( \43154 , \43100 , \43153 );
not \U$42778 ( \43155 , \43100 );
and \U$42779 ( \43156 , \43155 , \43152 );
nor \U$42780 ( \43157 , \43154 , \43156 );
not \U$42781 ( \43158 , \42945 );
not \U$42782 ( \43159 , \43158 );
not \U$42783 ( \43160 , \42951 );
or \U$42784 ( \43161 , \43159 , \43160 );
not \U$42785 ( \43162 , \42941 );
nand \U$42786 ( \43163 , \43162 , \42931 );
nand \U$42787 ( \43164 , \43161 , \43163 );
xor \U$42788 ( \43165 , \43157 , \43164 );
not \U$42789 ( \43166 , \43165 );
or \U$42790 ( \43167 , \43029 , \43166 );
or \U$42791 ( \43168 , \43165 , \43028 );
nand \U$42792 ( \43169 , \43167 , \43168 );
not \U$42793 ( \43170 , \43169 );
nand \U$42794 ( \43171 , \42966 , \43170 );
not \U$42795 ( \43172 , \42778 );
not \U$42796 ( \43173 , \43172 );
not \U$42797 ( \43174 , \42961 );
or \U$42798 ( \43175 , \43173 , \43174 );
or \U$42799 ( \43176 , \42961 , \43172 );
nand \U$42800 ( \43177 , \43175 , \43176 );
not \U$42801 ( \43178 , \41840 );
not \U$42802 ( \43179 , \41953 );
or \U$42803 ( \43180 , \43178 , \43179 );
not \U$42804 ( \43181 , \41953 );
nand \U$42805 ( \43182 , \43181 , \41841 );
nand \U$42806 ( \43183 , \41835 , \43182 );
nand \U$42807 ( \43184 , \43180 , \43183 );
or \U$42808 ( \43185 , \43177 , \43184 );
and \U$42809 ( \43186 , \42772 , \43171 , \43185 );
not \U$42810 ( \43187 , \43003 );
not \U$42811 ( \43188 , \43018 );
or \U$42812 ( \43189 , \43187 , \43188 );
nand \U$42813 ( \43190 , \43011 , \43017 );
nand \U$42814 ( \43191 , \43189 , \43190 );
and \U$42815 ( \43192 , RIae7a6f0_184, \11198 );
not \U$42816 ( \43193 , RIae7a6f0_184);
and \U$42817 ( \43194 , \43193 , \11804 );
or \U$42818 ( \43195 , \43192 , \43194 );
not \U$42819 ( \43196 , \43195 );
not \U$42820 ( \43197 , \36656 );
and \U$42821 ( \43198 , \43196 , \43197 );
and \U$42822 ( \43199 , \43142 , \9473 );
nor \U$42823 ( \43200 , \43198 , \43199 );
not \U$42824 ( \43201 , \43200 );
not \U$42825 ( \43202 , RIae7aab0_192);
and \U$42826 ( \43203 , RIae7aa38_191, \25333 );
not \U$42827 ( \43204 , RIae7aa38_191);
and \U$42828 ( \43205 , \43204 , \14691 );
or \U$42829 ( \43206 , \43203 , \43205 );
not \U$42830 ( \43207 , \43206 );
or \U$42831 ( \43208 , \43202 , \43207 );
nand \U$42832 ( \43209 , \43081 , \14668 );
nand \U$42833 ( \43210 , \43208 , \43209 );
not \U$42834 ( \43211 , \43210 );
or \U$42835 ( \43212 , \43201 , \43211 );
or \U$42836 ( \43213 , \43210 , \43200 );
nand \U$42837 ( \43214 , \43212 , \43213 );
nand \U$42838 ( \43215 , \43074 , \43064 );
not \U$42839 ( \43216 , \43054 );
nand \U$42840 ( \43217 , \43216 , \43063 );
and \U$42841 ( \43218 , \43215 , \43217 );
and \U$42842 ( \43219 , \43214 , \43218 );
not \U$42843 ( \43220 , \43214 );
not \U$42844 ( \43221 , \43218 );
and \U$42845 ( \43222 , \43220 , \43221 );
nor \U$42846 ( \43223 , \43219 , \43222 );
not \U$42847 ( \43224 , \43223 );
not \U$42848 ( \43225 , \43224 );
not \U$42849 ( \43226 , \43150 );
not \U$42850 ( \43227 , \43140 );
or \U$42851 ( \43228 , \43226 , \43227 );
or \U$42852 ( \43229 , \43139 , \43104 );
nand \U$42853 ( \43230 , \43228 , \43229 );
not \U$42854 ( \43231 , \43230 );
or \U$42855 ( \43232 , \43225 , \43231 );
or \U$42856 ( \43233 , \43230 , \43224 );
nand \U$42857 ( \43234 , \43232 , \43233 );
not \U$42858 ( \43235 , \43234 );
xor \U$42859 ( \43236 , \43191 , \43235 );
not \U$42860 ( \43237 , \9621 );
not \U$42861 ( \43238 , \11690 );
not \U$42862 ( \43239 , \16912 );
or \U$42863 ( \43240 , \43238 , \43239 );
or \U$42864 ( \43241 , \11665 , \11690 );
nand \U$42865 ( \43242 , \43240 , \43241 );
not \U$42866 ( \43243 , \43242 );
or \U$42867 ( \43244 , \43237 , \43243 );
nand \U$42868 ( \43245 , \43120 , \9643 );
nand \U$42869 ( \43246 , \43244 , \43245 );
buf \U$42870 ( \43247 , \43246 );
not \U$42871 ( \43248 , \43247 );
not \U$42872 ( \43249 , \43050 );
nand \U$42873 ( \43250 , \43249 , \43045 );
not \U$42874 ( \43251 , \43250 );
and \U$42875 ( \43252 , \43248 , \43251 );
and \U$42876 ( \43253 , \43247 , \43250 );
nor \U$42877 ( \43254 , \43252 , \43253 );
not \U$42878 ( \43255 , \10637 );
not \U$42879 ( \43256 , \43070 );
or \U$42880 ( \43257 , \43255 , \43256 );
not \U$42881 ( \43258 , RIae7a510_180);
not \U$42882 ( \43259 , \40490 );
or \U$42883 ( \43260 , \43258 , \43259 );
or \U$42884 ( \43261 , \40490 , RIae7a510_180);
nand \U$42885 ( \43262 , \43260 , \43261 );
nand \U$42886 ( \43263 , \43262 , \10631 );
nand \U$42887 ( \43264 , \43257 , \43263 );
xnor \U$42888 ( \43265 , \43254 , \43264 );
not \U$42889 ( \43266 , \43265 );
not \U$42890 ( \43267 , \43131 );
nand \U$42891 ( \43268 , \43267 , \43125 );
not \U$42892 ( \43269 , \43268 );
not \U$42893 ( \43270 , \43114 );
or \U$42894 ( \43271 , \43269 , \43270 );
nand \U$42895 ( \43272 , \43131 , \43124 );
nand \U$42896 ( \43273 , \43271 , \43272 );
not \U$42897 ( \43274 , \42991 );
not \U$42898 ( \43275 , \42982 );
and \U$42899 ( \43276 , \43274 , \43275 );
and \U$42900 ( \43277 , \42982 , \42991 );
nor \U$42901 ( \43278 , \43277 , \43002 );
nor \U$42902 ( \43279 , \43276 , \43278 );
nor \U$42903 ( \43280 , \43273 , \43279 );
not \U$42904 ( \43281 , \43280 );
nand \U$42905 ( \43282 , \43273 , \43279 );
nand \U$42906 ( \43283 , \43281 , \43282 );
not \U$42907 ( \43284 , \43283 );
or \U$42908 ( \43285 , \43266 , \43284 );
or \U$42909 ( \43286 , \43283 , \43265 );
nand \U$42910 ( \43287 , \43285 , \43286 );
not \U$42911 ( \43288 , \43097 );
not \U$42912 ( \43289 , \43152 );
or \U$42913 ( \43290 , \43288 , \43289 );
nand \U$42914 ( \43291 , \43290 , \43099 );
xor \U$42915 ( \43292 , \43287 , \43291 );
not \U$42916 ( \43293 , \10695 );
not \U$42917 ( \43294 , \42978 );
or \U$42918 ( \43295 , \43293 , \43294 );
not \U$42919 ( \43296 , \10625 );
not \U$42920 ( \43297 , \10007 );
or \U$42921 ( \43298 , \43296 , \43297 );
nand \U$42922 ( \43299 , \11260 , RIae7a498_179);
nand \U$42923 ( \43300 , \43298 , \43299 );
nand \U$42924 ( \43301 , \43300 , \10675 );
nand \U$42925 ( \43302 , \43295 , \43301 );
not \U$42926 ( \43303 , \9758 );
not \U$42927 ( \43304 , \42998 );
or \U$42928 ( \43305 , \43303 , \43304 );
not \U$42929 ( \43306 , \10658 );
not \U$42930 ( \43307 , \36204 );
or \U$42931 ( \43308 , \43306 , \43307 );
nand \U$42932 ( \43309 , \10171 , RIae7a150_172);
nand \U$42933 ( \43310 , \43308 , \43309 );
nand \U$42934 ( \43311 , \43310 , \9776 );
nand \U$42935 ( \43312 , \43305 , \43311 );
xor \U$42936 ( \43313 , \43302 , \43312 );
not \U$42937 ( \43314 , \11205 );
not \U$42938 ( \43315 , \43091 );
or \U$42939 ( \43316 , \43314 , \43315 );
and \U$42940 ( \43317 , RIae7a8d0_188, \14657 );
not \U$42941 ( \43318 , RIae7a8d0_188);
and \U$42942 ( \43319 , \43318 , \19736 );
or \U$42943 ( \43320 , \43317 , \43319 );
nand \U$42944 ( \43321 , \43320 , \10275 );
nand \U$42945 ( \43322 , \43316 , \43321 );
xor \U$42946 ( \43323 , \43313 , \43322 );
or \U$42947 ( \43324 , \43085 , \43075 );
nand \U$42948 ( \43325 , \43324 , \43095 );
nand \U$42949 ( \43326 , \43085 , \43075 );
nand \U$42950 ( \43327 , \43325 , \43326 );
xor \U$42951 ( \43328 , \43323 , \43327 );
not \U$42952 ( \43329 , \10542 );
xor \U$42953 ( \43330 , \19025 , RIae7a060_170);
not \U$42954 ( \43331 , \43330 );
or \U$42955 ( \43332 , \43329 , \43331 );
nand \U$42956 ( \43333 , \42987 , \9728 );
nand \U$42957 ( \43334 , \43332 , \43333 );
nand \U$42958 ( \43335 , \12857 , \9493 );
not \U$42959 ( \43336 , \43335 );
not \U$42960 ( \43337 , \9813 );
not \U$42961 ( \43338 , \9799 );
not \U$42962 ( \43339 , \36790 );
or \U$42963 ( \43340 , \43338 , \43339 );
nand \U$42964 ( \43341 , \36793 , RIae7a2b8_175);
nand \U$42965 ( \43342 , \43340 , \43341 );
not \U$42966 ( \43343 , \43342 );
or \U$42967 ( \43344 , \43337 , \43343 );
or \U$42968 ( \43345 , \43040 , \43043 );
nand \U$42969 ( \43346 , \43344 , \43345 );
not \U$42970 ( \43347 , \43346 );
or \U$42971 ( \43348 , \43336 , \43347 );
or \U$42972 ( \43349 , \43346 , \43335 );
nand \U$42973 ( \43350 , \43348 , \43349 );
not \U$42974 ( \43351 , \9699 );
not \U$42975 ( \43352 , \11114 );
not \U$42976 ( \43353 , \11318 );
or \U$42977 ( \43354 , \43352 , \43353 );
or \U$42978 ( \43355 , \10272 , \11114 );
nand \U$42979 ( \43356 , \43354 , \43355 );
not \U$42980 ( \43357 , \43356 );
or \U$42981 ( \43358 , \43351 , \43357 );
nand \U$42982 ( \43359 , \43059 , \9687 );
nand \U$42983 ( \43360 , \43358 , \43359 );
xor \U$42984 ( \43361 , \43350 , \43360 );
not \U$42985 ( \43362 , \43361 );
not \U$42986 ( \43363 , \9549 );
not \U$42987 ( \43364 , \43110 );
or \U$42988 ( \43365 , \43363 , \43364 );
and \U$42989 ( \43366 , RIae7a7e0_186, \10461 );
not \U$42990 ( \43367 , RIae7a7e0_186);
and \U$42991 ( \43368 , \43367 , \10465 );
or \U$42992 ( \43369 , \43366 , \43368 );
nand \U$42993 ( \43370 , \43369 , \10519 );
nand \U$42994 ( \43371 , \43365 , \43370 );
not \U$42995 ( \43372 , \43371 );
not \U$42996 ( \43373 , \43372 );
or \U$42997 ( \43374 , \43362 , \43373 );
or \U$42998 ( \43375 , \43372 , \43361 );
nand \U$42999 ( \43376 , \43374 , \43375 );
xor \U$43000 ( \43377 , \43334 , \43376 );
xor \U$43001 ( \43378 , \43328 , \43377 );
xnor \U$43002 ( \43379 , \43292 , \43378 );
xor \U$43003 ( \43380 , \43236 , \43379 );
not \U$43004 ( \43381 , \43027 );
and \U$43005 ( \43382 , \43023 , \43381 );
and \U$43006 ( \43383 , \42972 , \43022 );
nor \U$43007 ( \43384 , \43382 , \43383 );
xor \U$43008 ( \43385 , \43380 , \43384 );
not \U$43009 ( \43386 , \43028 );
and \U$43010 ( \43387 , \43165 , \43386 );
and \U$43011 ( \43388 , \43157 , \43164 );
nor \U$43012 ( \43389 , \43387 , \43388 );
nand \U$43013 ( \43390 , \43385 , \43389 );
not \U$43014 ( \43391 , \10275 );
and \U$43015 ( \43392 , RIae7a8d0_188, \14110 );
not \U$43016 ( \43393 , RIae7a8d0_188);
and \U$43017 ( \43394 , \43393 , \12615 );
nor \U$43018 ( \43395 , \43392 , \43394 );
not \U$43019 ( \43396 , \43395 );
or \U$43020 ( \43397 , \43391 , \43396 );
nand \U$43021 ( \43398 , \43320 , \14510 );
nand \U$43022 ( \43399 , \43397 , \43398 );
not \U$43023 ( \43400 , \10519 );
and \U$43024 ( \43401 , \16752 , RIae7a7e0_186);
not \U$43025 ( \43402 , \16752 );
and \U$43026 ( \43403 , \43402 , \9541 );
nor \U$43027 ( \43404 , \43401 , \43403 );
not \U$43028 ( \43405 , \43404 );
or \U$43029 ( \43406 , \43400 , \43405 );
nand \U$43030 ( \43407 , \43369 , \9549 );
nand \U$43031 ( \43408 , \43406 , \43407 );
nand \U$43032 ( \43409 , \43399 , \43408 );
or \U$43033 ( \43410 , \43399 , \43408 );
nand \U$43034 ( \43411 , \43409 , \43410 );
not \U$43035 ( \43412 , RIae7aab0_192);
and \U$43036 ( \43413 , RIae7aa38_191, \17387 );
not \U$43037 ( \43414 , RIae7aa38_191);
and \U$43038 ( \43415 , \43414 , \23180 );
or \U$43039 ( \43416 , \43413 , \43415 );
not \U$43040 ( \43417 , \43416 );
or \U$43041 ( \43418 , \43412 , \43417 );
nand \U$43042 ( \43419 , \43206 , \14667 );
nand \U$43043 ( \43420 , \43418 , \43419 );
xor \U$43044 ( \43421 , \43411 , \43420 );
not \U$43045 ( \43422 , \43280 );
not \U$43046 ( \43423 , \43265 );
nand \U$43047 ( \43424 , \43282 , \43423 );
nand \U$43048 ( \43425 , \43422 , \43424 );
or \U$43049 ( \43426 , \43421 , \43425 );
nand \U$43050 ( \43427 , \43421 , \43425 );
nand \U$43051 ( \43428 , \43426 , \43427 );
xor \U$43052 ( \43429 , \43323 , \43327 );
and \U$43053 ( \43430 , \43429 , \43377 );
and \U$43054 ( \43431 , \43323 , \43327 );
or \U$43055 ( \43432 , \43430 , \43431 );
and \U$43056 ( \43433 , \43428 , \43432 );
not \U$43057 ( \43434 , \43428 );
not \U$43058 ( \43435 , \43432 );
and \U$43059 ( \43436 , \43434 , \43435 );
nor \U$43060 ( \43437 , \43433 , \43436 );
or \U$43061 ( \43438 , \43287 , \43378 );
nand \U$43062 ( \43439 , \43438 , \43291 );
nand \U$43063 ( \43440 , \43378 , \43287 );
and \U$43064 ( \43441 , \43439 , \43440 );
xor \U$43065 ( \43442 , \43437 , \43441 );
not \U$43066 ( \43443 , \11114 );
not \U$43067 ( \43444 , \10195 );
or \U$43068 ( \43445 , \43443 , \43444 );
nand \U$43069 ( \43446 , \19689 , RIae7a240_174);
nand \U$43070 ( \43447 , \43445 , \43446 );
not \U$43071 ( \43448 , \43447 );
or \U$43072 ( \43449 , \43448 , \30532 );
not \U$43073 ( \43450 , \43356 );
not \U$43074 ( \43451 , \9687 );
or \U$43075 ( \43452 , \43450 , \43451 );
nand \U$43076 ( \43453 , \43449 , \43452 );
not \U$43077 ( \43454 , \43360 );
not \U$43078 ( \43455 , \43350 );
or \U$43079 ( \43456 , \43454 , \43455 );
not \U$43080 ( \43457 , \43335 );
nand \U$43081 ( \43458 , \43457 , \43346 );
nand \U$43082 ( \43459 , \43456 , \43458 );
xor \U$43083 ( \43460 , \43453 , \43459 );
not \U$43084 ( \43461 , RIae7a510_180);
and \U$43085 ( \43462 , \27672 , \43461 );
not \U$43086 ( \43463 , \27672 );
and \U$43087 ( \43464 , \43463 , RIae7a510_180);
nor \U$43088 ( \43465 , \43462 , \43464 );
not \U$43089 ( \43466 , \43465 );
or \U$43090 ( \43467 , \43466 , \12232 );
not \U$43091 ( \43468 , \43262 );
not \U$43092 ( \43469 , \11400 );
or \U$43093 ( \43470 , \43468 , \43469 );
nand \U$43094 ( \43471 , \43467 , \43470 );
xor \U$43095 ( \43472 , \43460 , \43471 );
not \U$43096 ( \43473 , \9776 );
and \U$43097 ( \43474 , RIae7a150_172, \10067 );
not \U$43098 ( \43475 , RIae7a150_172);
and \U$43099 ( \43476 , \43475 , \10066 );
or \U$43100 ( \43477 , \43474 , \43476 );
not \U$43101 ( \43478 , \43477 );
or \U$43102 ( \43479 , \43473 , \43478 );
nand \U$43103 ( \43480 , \43310 , \9758 );
nand \U$43104 ( \43481 , \43479 , \43480 );
not \U$43105 ( \43482 , \10676 );
not \U$43106 ( \43483 , RIae7a498_179);
not \U$43107 ( \43484 , \9875 );
or \U$43108 ( \43485 , \43483 , \43484 );
or \U$43109 ( \43486 , \13896 , RIae7a498_179);
nand \U$43110 ( \43487 , \43485 , \43486 );
not \U$43111 ( \43488 , \43487 );
or \U$43112 ( \43489 , \43482 , \43488 );
nand \U$43113 ( \43490 , \43300 , \10695 );
nand \U$43114 ( \43491 , \43489 , \43490 );
not \U$43115 ( \43492 , \43491 );
xor \U$43116 ( \43493 , \43481 , \43492 );
not \U$43117 ( \43494 , \9745 );
and \U$43118 ( \43495 , RIae7a060_170, \41210 );
not \U$43119 ( \43496 , RIae7a060_170);
not \U$43120 ( \43497 , \40195 );
and \U$43121 ( \43498 , \43496 , \43497 );
or \U$43122 ( \43499 , \43495 , \43498 );
not \U$43123 ( \43500 , \43499 );
or \U$43124 ( \43501 , \43494 , \43500 );
nand \U$43125 ( \43502 , \43330 , \9730 );
nand \U$43126 ( \43503 , \43501 , \43502 );
and \U$43127 ( \43504 , \43493 , \43503 );
not \U$43128 ( \43505 , \43493 );
not \U$43129 ( \43506 , \43503 );
and \U$43130 ( \43507 , \43505 , \43506 );
nor \U$43131 ( \43508 , \43504 , \43507 );
not \U$43132 ( \43509 , \43508 );
xor \U$43133 ( \43510 , \43472 , \43509 );
not \U$43134 ( \43511 , \43334 );
not \U$43135 ( \43512 , \43376 );
or \U$43136 ( \43513 , \43511 , \43512 );
not \U$43137 ( \43514 , \43372 );
nand \U$43138 ( \43515 , \43514 , \43361 );
nand \U$43139 ( \43516 , \43513 , \43515 );
xnor \U$43140 ( \43517 , \43510 , \43516 );
xor \U$43141 ( \43518 , \43302 , \43312 );
and \U$43142 ( \43519 , \43518 , \43322 );
and \U$43143 ( \43520 , \43302 , \43312 );
or \U$43144 ( \43521 , \43519 , \43520 );
not \U$43145 ( \43522 , \43250 );
not \U$43146 ( \43523 , \43246 );
not \U$43147 ( \43524 , \43523 );
or \U$43148 ( \43525 , \43522 , \43524 );
nand \U$43149 ( \43526 , \43525 , \43264 );
not \U$43150 ( \43527 , \43250 );
nand \U$43151 ( \43528 , \43527 , \43246 );
nand \U$43152 ( \43529 , \43526 , \43528 );
not \U$43153 ( \43530 , \43529 );
or \U$43154 ( \43531 , RIae7a2b8_175, RIae7a678_183);
nand \U$43155 ( \43532 , \43531 , \12857 );
and \U$43156 ( \43533 , \43532 , \22947 );
not \U$43157 ( \43534 , \9493 );
and \U$43158 ( \43535 , \12750 , \11069 );
not \U$43159 ( \43536 , \12750 );
and \U$43160 ( \43537 , \43536 , RIae79fe8_169);
nor \U$43161 ( \43538 , \43535 , \43537 );
not \U$43162 ( \43539 , \43538 );
or \U$43163 ( \43540 , \43534 , \43539 );
xnor \U$43164 ( \43541 , \16890 , RIae79fe8_169);
nand \U$43165 ( \43542 , \43541 , \9499 );
nand \U$43166 ( \43543 , \43540 , \43542 );
xor \U$43167 ( \43544 , \43533 , \43543 );
not \U$43168 ( \43545 , \9813 );
not \U$43169 ( \43546 , RIae7a2b8_175);
not \U$43170 ( \43547 , \39806 );
or \U$43171 ( \43548 , \43546 , \43547 );
nand \U$43172 ( \43549 , \42523 , \29995 );
nand \U$43173 ( \43550 , \43548 , \43549 );
not \U$43174 ( \43551 , \43550 );
or \U$43175 ( \43552 , \43545 , \43551 );
nand \U$43176 ( \43553 , \43342 , \9791 );
nand \U$43177 ( \43554 , \43552 , \43553 );
xor \U$43178 ( \43555 , \43544 , \43554 );
not \U$43179 ( \43556 , \9621 );
not \U$43180 ( \43557 , \11690 );
not \U$43181 ( \43558 , \33415 );
or \U$43182 ( \43559 , \43557 , \43558 );
nand \U$43183 ( \43560 , \17955 , RIae7a3a8_177);
nand \U$43184 ( \43561 , \43559 , \43560 );
not \U$43185 ( \43562 , \43561 );
or \U$43186 ( \43563 , \43556 , \43562 );
nand \U$43187 ( \43564 , \43242 , \9643 );
nand \U$43188 ( \43565 , \43563 , \43564 );
xor \U$43189 ( \43566 , \43555 , \43565 );
not \U$43190 ( \43567 , \43566 );
not \U$43191 ( \43568 , \43567 );
or \U$43192 ( \43569 , \43530 , \43568 );
not \U$43193 ( \43570 , \43529 );
nand \U$43194 ( \43571 , \43570 , \43566 );
nand \U$43195 ( \43572 , \43569 , \43571 );
not \U$43196 ( \43573 , \43572 );
not \U$43197 ( \43574 , \9478 );
not \U$43198 ( \43575 , \27644 );
not \U$43199 ( \43576 , \22557 );
or \U$43200 ( \43577 , \43575 , \43576 );
nand \U$43201 ( \43578 , \22560 , RIae7a6f0_184);
nand \U$43202 ( \43579 , \43577 , \43578 );
not \U$43203 ( \43580 , \43579 );
or \U$43204 ( \43581 , \43574 , \43580 );
not \U$43205 ( \43582 , \43195 );
nand \U$43206 ( \43583 , \43582 , \9473 );
nand \U$43207 ( \43584 , \43581 , \43583 );
not \U$43208 ( \43585 , \43584 );
not \U$43209 ( \43586 , \43585 );
and \U$43210 ( \43587 , \43573 , \43586 );
and \U$43211 ( \43588 , \43572 , \43585 );
nor \U$43212 ( \43589 , \43587 , \43588 );
not \U$43213 ( \43590 , \43589 );
xor \U$43214 ( \43591 , \43521 , \43590 );
not \U$43215 ( \43592 , \43221 );
not \U$43216 ( \43593 , \43214 );
or \U$43217 ( \43594 , \43592 , \43593 );
not \U$43218 ( \43595 , \43200 );
nand \U$43219 ( \43596 , \43595 , \43210 );
nand \U$43220 ( \43597 , \43594 , \43596 );
xnor \U$43221 ( \43598 , \43591 , \43597 );
xor \U$43222 ( \43599 , \43517 , \43598 );
nand \U$43223 ( \43600 , \43230 , \43223 );
not \U$43224 ( \43601 , \43600 );
not \U$43225 ( \43602 , \43191 );
or \U$43226 ( \43603 , \43601 , \43602 );
not \U$43227 ( \43604 , \43230 );
nand \U$43228 ( \43605 , \43604 , \43224 );
nand \U$43229 ( \43606 , \43603 , \43605 );
not \U$43230 ( \43607 , \43606 );
xor \U$43231 ( \43608 , \43599 , \43607 );
xor \U$43232 ( \43609 , \43442 , \43608 );
xor \U$43233 ( \43610 , \43236 , \43379 );
and \U$43234 ( \43611 , \43610 , \43384 );
and \U$43235 ( \43612 , \43236 , \43379 );
or \U$43236 ( \43613 , \43611 , \43612 );
nand \U$43237 ( \43614 , \43609 , \43613 );
and \U$43238 ( \43615 , \43390 , \43614 );
nand \U$43239 ( \43616 , \43186 , \43615 );
nand \U$43240 ( \43617 , \43177 , \43184 );
nand \U$43241 ( \43618 , \42965 , \43169 );
nand \U$43242 ( \43619 , \43617 , \43618 );
nand \U$43243 ( \43620 , \43171 , \43619 );
not \U$43244 ( \43621 , \43390 );
or \U$43245 ( \43622 , \43620 , \43621 );
or \U$43246 ( \43623 , \43385 , \43389 );
nand \U$43247 ( \43624 , \43622 , \43623 );
nand \U$43248 ( \43625 , \43624 , \43614 );
or \U$43249 ( \43626 , \43609 , \43613 );
nand \U$43250 ( \43627 , \43616 , \43625 , \43626 );
not \U$43251 ( \43628 , \40665 );
and \U$43252 ( \43629 , \40676 , \43628 );
not \U$43253 ( \43630 , \40676 );
and \U$43254 ( \43631 , \43630 , \40665 );
nor \U$43255 ( \43632 , \43629 , \43631 );
not \U$43256 ( \43633 , \43632 );
xor \U$43257 ( \43634 , \40611 , \40628 );
not \U$43258 ( \43635 , \43634 );
or \U$43259 ( \43636 , \43633 , \43635 );
or \U$43260 ( \43637 , \43634 , \43632 );
nand \U$43261 ( \43638 , \43636 , \43637 );
not \U$43262 ( \43639 , \40499 );
not \U$43263 ( \43640 , \40514 );
or \U$43264 ( \43641 , \43639 , \43640 );
or \U$43265 ( \43642 , \40514 , \40499 );
nand \U$43266 ( \43643 , \43641 , \43642 );
not \U$43267 ( \43644 , \43643 );
not \U$43268 ( \43645 , \9516 );
not \U$43269 ( \43646 , \40649 );
or \U$43270 ( \43647 , \43645 , \43646 );
not \U$43271 ( \43648 , \18027 );
not \U$43272 ( \43649 , \10845 );
or \U$43273 ( \43650 , \43648 , \43649 );
nand \U$43274 ( \43651 , \16651 , RIae79fe8_169);
nand \U$43275 ( \43652 , \43650 , \43651 );
nand \U$43276 ( \43653 , \43652 , \9499 );
nand \U$43277 ( \43654 , \43647 , \43653 );
not \U$43278 ( \43655 , \43654 );
or \U$43279 ( \43656 , \43644 , \43655 );
not \U$43280 ( \43657 , \43643 );
not \U$43281 ( \43658 , \43654 );
not \U$43282 ( \43659 , \43658 );
or \U$43283 ( \43660 , \43657 , \43659 );
or \U$43284 ( \43661 , \43658 , \43643 );
nand \U$43285 ( \43662 , \43660 , \43661 );
not \U$43286 ( \43663 , \16135 );
not \U$43287 ( \43664 , \40528 );
or \U$43288 ( \43665 , \43663 , \43664 );
not \U$43289 ( \43666 , RIae7a2b8_175);
not \U$43290 ( \43667 , \28259 );
or \U$43291 ( \43668 , \43666 , \43667 );
or \U$43292 ( \43669 , \11318 , RIae7a2b8_175);
nand \U$43293 ( \43670 , \43668 , \43669 );
not \U$43294 ( \43671 , \43670 );
nand \U$43295 ( \43672 , \43671 , \9792 );
nand \U$43296 ( \43673 , \43665 , \43672 );
nand \U$43297 ( \43674 , \43662 , \43673 );
nand \U$43298 ( \43675 , \43656 , \43674 );
not \U$43299 ( \43676 , \10510 );
not \U$43300 ( \43677 , RIae7a7e0_186);
not \U$43301 ( \43678 , \19422 );
or \U$43302 ( \43679 , \43677 , \43678 );
or \U$43303 ( \43680 , \16766 , RIae7a7e0_186);
nand \U$43304 ( \43681 , \43679 , \43680 );
not \U$43305 ( \43682 , \43681 );
or \U$43306 ( \43683 , \43676 , \43682 );
nand \U$43307 ( \43684 , \40547 , \29519 );
nand \U$43308 ( \43685 , \43683 , \43684 );
xor \U$43309 ( \43686 , \43675 , \43685 );
not \U$43310 ( \43687 , RIae7a8d0_188);
not \U$43311 ( \43688 , \17387 );
or \U$43312 ( \43689 , \43687 , \43688 );
nand \U$43313 ( \43690 , \21747 , \18088 );
nand \U$43314 ( \43691 , \43689 , \43690 );
not \U$43315 ( \43692 , \43691 );
not \U$43316 ( \43693 , \14510 );
or \U$43317 ( \43694 , \43692 , \43693 );
nand \U$43318 ( \43695 , \40475 , \10275 );
nand \U$43319 ( \43696 , \43694 , \43695 );
and \U$43320 ( \43697 , \43686 , \43696 );
and \U$43321 ( \43698 , \43675 , \43685 );
or \U$43322 ( \43699 , \43697 , \43698 );
xnor \U$43323 ( \43700 , \43638 , \43699 );
not \U$43324 ( \43701 , \43700 );
not \U$43325 ( \43702 , \9729 );
and \U$43326 ( \43703 , RIae7a060_170, \9608 );
not \U$43327 ( \43704 , RIae7a060_170);
and \U$43328 ( \43705 , \43704 , \12077 );
or \U$43329 ( \43706 , \43703 , \43705 );
not \U$43330 ( \43707 , \43706 );
or \U$43331 ( \43708 , \43702 , \43707 );
nand \U$43332 ( \43709 , \40563 , \9744 );
nand \U$43333 ( \43710 , \43708 , \43709 );
not \U$43334 ( \43711 , \43710 );
not \U$43335 ( \43712 , \43711 );
not \U$43336 ( \43713 , \40494 );
and \U$43337 ( \43714 , \40534 , \43713 );
not \U$43338 ( \43715 , \40534 );
and \U$43339 ( \43716 , \43715 , \40494 );
nor \U$43340 ( \43717 , \43714 , \43716 );
not \U$43341 ( \43718 , \43717 );
not \U$43342 ( \43719 , \43718 );
or \U$43343 ( \43720 , \43712 , \43719 );
nand \U$43344 ( \43721 , \43710 , \43717 );
nand \U$43345 ( \43722 , \43720 , \43721 );
not \U$43346 ( \43723 , \14667 );
and \U$43347 ( \43724 , RIae7aa38_191, \12687 );
not \U$43348 ( \43725 , RIae7aa38_191);
and \U$43349 ( \43726 , \43725 , \6230 );
or \U$43350 ( \43727 , \43724 , \43726 );
not \U$43351 ( \43728 , \43727 );
or \U$43352 ( \43729 , \43723 , \43728 );
nand \U$43353 ( \43730 , \40580 , RIae7aab0_192);
nand \U$43354 ( \43731 , \43729 , \43730 );
and \U$43355 ( \43732 , \43722 , \43731 );
not \U$43356 ( \43733 , \43722 );
not \U$43357 ( \43734 , \43731 );
and \U$43358 ( \43735 , \43733 , \43734 );
nor \U$43359 ( \43736 , \43732 , \43735 );
not \U$43360 ( \43737 , \10631 );
and \U$43361 ( \43738 , \11260 , \43461 );
not \U$43362 ( \43739 , \11260 );
and \U$43363 ( \43740 , \43739 , RIae7a510_180);
nor \U$43364 ( \43741 , \43738 , \43740 );
not \U$43365 ( \43742 , \43741 );
or \U$43366 ( \43743 , \43737 , \43742 );
nand \U$43367 ( \43744 , \43465 , \10637 );
nand \U$43368 ( \43745 , \43743 , \43744 );
and \U$43369 ( \43746 , \12857 , \6212 );
not \U$43370 ( \43747 , \43746 );
not \U$43371 ( \43748 , \9493 );
not \U$43372 ( \43749 , \43652 );
or \U$43373 ( \43750 , \43748 , \43749 );
nand \U$43374 ( \43751 , \43538 , \9499 );
nand \U$43375 ( \43752 , \43750 , \43751 );
not \U$43376 ( \43753 , \43752 );
not \U$43377 ( \43754 , \43753 );
or \U$43378 ( \43755 , \43747 , \43754 );
or \U$43379 ( \43756 , \43753 , \43746 );
nand \U$43380 ( \43757 , \43755 , \43756 );
not \U$43381 ( \43758 , \9791 );
not \U$43382 ( \43759 , \43550 );
or \U$43383 ( \43760 , \43758 , \43759 );
or \U$43384 ( \43761 , \43670 , \9786 );
nand \U$43385 ( \43762 , \43760 , \43761 );
xor \U$43386 ( \43763 , \43757 , \43762 );
xor \U$43387 ( \43764 , \43745 , \43763 );
not \U$43388 ( \43765 , \43764 );
not \U$43389 ( \43766 , \9730 );
not \U$43390 ( \43767 , \43499 );
or \U$43391 ( \43768 , \43766 , \43767 );
and \U$43392 ( \43769 , RIae7a060_170, \10465 );
not \U$43393 ( \43770 , RIae7a060_170);
and \U$43394 ( \43771 , \43770 , \10464 );
nor \U$43395 ( \43772 , \43769 , \43771 );
nand \U$43396 ( \43773 , \43772 , \10542 );
nand \U$43397 ( \43774 , \43768 , \43773 );
not \U$43398 ( \43775 , \43774 );
or \U$43399 ( \43776 , \43765 , \43775 );
nand \U$43400 ( \43777 , \43745 , \43763 );
nand \U$43401 ( \43778 , \43776 , \43777 );
not \U$43402 ( \43779 , \43778 );
not \U$43403 ( \43780 , RIae7aab0_192);
not \U$43404 ( \43781 , \43727 );
or \U$43405 ( \43782 , \43780 , \43781 );
and \U$43406 ( \43783 , \9316 , \11326 );
not \U$43407 ( \43784 , \9316 );
and \U$43408 ( \43785 , \43784 , RIae7aa38_191);
nor \U$43409 ( \43786 , \43783 , \43785 );
nand \U$43410 ( \43787 , \43786 , \14667 );
nand \U$43411 ( \43788 , \43782 , \43787 );
not \U$43412 ( \43789 , \43788 );
not \U$43413 ( \43790 , \43789 );
not \U$43414 ( \43791 , \9621 );
and \U$43415 ( \43792 , \19035 , \11690 );
not \U$43416 ( \43793 , \19035 );
and \U$43417 ( \43794 , \43793 , RIae7a3a8_177);
nor \U$43418 ( \43795 , \43792 , \43794 );
not \U$43419 ( \43796 , \43795 );
or \U$43420 ( \43797 , \43791 , \43796 );
and \U$43421 ( \43798 , RIae7a3a8_177, \10142 );
not \U$43422 ( \43799 , RIae7a3a8_177);
and \U$43423 ( \43800 , \43799 , \40490 );
nor \U$43424 ( \43801 , \43798 , \43800 );
nand \U$43425 ( \43802 , \43801 , \9643 );
nand \U$43426 ( \43803 , \43797 , \43802 );
not \U$43427 ( \43804 , \43762 );
not \U$43428 ( \43805 , \43757 );
or \U$43429 ( \43806 , \43804 , \43805 );
nand \U$43430 ( \43807 , \43752 , \43746 );
nand \U$43431 ( \43808 , \43806 , \43807 );
not \U$43432 ( \43809 , \43808 );
not \U$43433 ( \43810 , \9699 );
not \U$43434 ( \43811 , \40484 );
or \U$43435 ( \43812 , \43810 , \43811 );
not \U$43436 ( \43813 , \11114 );
not \U$43437 ( \43814 , \16912 );
or \U$43438 ( \43815 , \43813 , \43814 );
or \U$43439 ( \43816 , \10043 , \19623 );
nand \U$43440 ( \43817 , \43815 , \43816 );
nand \U$43441 ( \43818 , \43817 , \9687 );
nand \U$43442 ( \43819 , \43812 , \43818 );
not \U$43443 ( \43820 , \43819 );
not \U$43444 ( \43821 , \43820 );
or \U$43445 ( \43822 , \43809 , \43821 );
or \U$43446 ( \43823 , \43820 , \43808 );
nand \U$43447 ( \43824 , \43822 , \43823 );
xor \U$43448 ( \43825 , \43803 , \43824 );
not \U$43449 ( \43826 , \43825 );
or \U$43450 ( \43827 , \43790 , \43826 );
or \U$43451 ( \43828 , \43825 , \43789 );
nand \U$43452 ( \43829 , \43827 , \43828 );
not \U$43453 ( \43830 , \43829 );
or \U$43454 ( \43831 , \43779 , \43830 );
nand \U$43455 ( \43832 , \43825 , \43788 );
nand \U$43456 ( \43833 , \43831 , \43832 );
xor \U$43457 ( \43834 , \43736 , \43833 );
xor \U$43458 ( \43835 , \43675 , \43685 );
xor \U$43459 ( \43836 , \43835 , \43696 );
and \U$43460 ( \43837 , \43834 , \43836 );
and \U$43461 ( \43838 , \43736 , \43833 );
or \U$43462 ( \43839 , \43837 , \43838 );
not \U$43463 ( \43840 , \43839 );
or \U$43464 ( \43841 , \43701 , \43840 );
or \U$43465 ( \43842 , \43839 , \43700 );
nand \U$43466 ( \43843 , \43841 , \43842 );
not \U$43467 ( \43844 , \43662 );
not \U$43468 ( \43845 , \43673 );
not \U$43469 ( \43846 , \43845 );
and \U$43470 ( \43847 , \43844 , \43846 );
and \U$43471 ( \43848 , \43662 , \43845 );
nor \U$43472 ( \43849 , \43847 , \43848 );
not \U$43473 ( \43850 , \9745 );
not \U$43474 ( \43851 , \43706 );
or \U$43475 ( \43852 , \43850 , \43851 );
nand \U$43476 ( \43853 , \43772 , \9730 );
nand \U$43477 ( \43854 , \43852 , \43853 );
xnor \U$43478 ( \43855 , \43849 , \43854 );
xor \U$43479 ( \43856 , RIae7a6f0_184, \12614 );
not \U$43480 ( \43857 , \43856 );
or \U$43481 ( \43858 , \43857 , \36656 );
and \U$43482 ( \43859 , RIae7a6f0_184, \13302 );
not \U$43483 ( \43860 , RIae7a6f0_184);
and \U$43484 ( \43861 , \43860 , \16786 );
or \U$43485 ( \43862 , \43859 , \43861 );
not \U$43486 ( \43863 , \43862 );
or \U$43487 ( \43864 , \43863 , \35746 );
nand \U$43488 ( \43865 , \43858 , \43864 );
nand \U$43489 ( \43866 , \43855 , \43865 );
not \U$43490 ( \43867 , \43849 );
nand \U$43491 ( \43868 , \43867 , \43854 );
and \U$43492 ( \43869 , \43866 , \43868 );
not \U$43493 ( \43870 , \43869 );
not \U$43494 ( \43871 , \43870 );
not \U$43495 ( \43872 , \10519 );
not \U$43496 ( \43873 , \43681 );
or \U$43497 ( \43874 , \43872 , \43873 );
xnor \U$43498 ( \43875 , \9412 , RIae7a7e0_186);
nand \U$43499 ( \43876 , \43875 , \10510 );
nand \U$43500 ( \43877 , \43874 , \43876 );
not \U$43501 ( \43878 , \43877 );
and \U$43502 ( \43879 , \43533 , \43543 );
not \U$43503 ( \43880 , \9699 );
not \U$43504 ( \43881 , \43817 );
or \U$43505 ( \43882 , \43880 , \43881 );
nand \U$43506 ( \43883 , \43447 , \9687 );
nand \U$43507 ( \43884 , \43882 , \43883 );
xor \U$43508 ( \43885 , \43879 , \43884 );
not \U$43509 ( \43886 , \9643 );
not \U$43510 ( \43887 , \43561 );
or \U$43511 ( \43888 , \43886 , \43887 );
nand \U$43512 ( \43889 , \43801 , \9621 );
nand \U$43513 ( \43890 , \43888 , \43889 );
and \U$43514 ( \43891 , \43885 , \43890 );
and \U$43515 ( \43892 , \43879 , \43884 );
nor \U$43516 ( \43893 , \43891 , \43892 );
not \U$43517 ( \43894 , \43893 );
not \U$43518 ( \43895 , \43691 );
not \U$43519 ( \43896 , \10275 );
or \U$43520 ( \43897 , \43895 , \43896 );
and \U$43521 ( \43898 , RIae7a8d0_188, \25333 );
not \U$43522 ( \43899 , RIae7a8d0_188);
and \U$43523 ( \43900 , \43899 , \14691 );
or \U$43524 ( \43901 , \43898 , \43900 );
nand \U$43525 ( \43902 , \43901 , \11205 );
nand \U$43526 ( \43903 , \43897 , \43902 );
not \U$43527 ( \43904 , \43903 );
or \U$43528 ( \43905 , \43894 , \43904 );
or \U$43529 ( \43906 , \43903 , \43893 );
nand \U$43530 ( \43907 , \43905 , \43906 );
not \U$43531 ( \43908 , \43907 );
or \U$43532 ( \43909 , \43878 , \43908 );
not \U$43533 ( \43910 , \43893 );
nand \U$43534 ( \43911 , \43910 , \43903 );
nand \U$43535 ( \43912 , \43909 , \43911 );
not \U$43536 ( \43913 , \11087 );
not \U$43537 ( \43914 , \10658 );
not \U$43538 ( \43915 , \43497 );
or \U$43539 ( \43916 , \43914 , \43915 );
nand \U$43540 ( \43917 , \41024 , RIae7a150_172);
nand \U$43541 ( \43918 , \43916 , \43917 );
not \U$43542 ( \43919 , \43918 );
or \U$43543 ( \43920 , \43913 , \43919 );
nand \U$43544 ( \43921 , \40572 , \9776 );
nand \U$43545 ( \43922 , \43920 , \43921 );
xor \U$43546 ( \43923 , \40636 , \40641 );
xor \U$43547 ( \43924 , \43923 , \40651 );
not \U$43548 ( \43925 , \43924 );
not \U$43549 ( \43926 , \9643 );
not \U$43550 ( \43927 , \43795 );
or \U$43551 ( \43928 , \43926 , \43927 );
nand \U$43552 ( \43929 , \40609 , \9621 );
nand \U$43553 ( \43930 , \43928 , \43929 );
not \U$43554 ( \43931 , \43930 );
not \U$43555 ( \43932 , \43931 );
or \U$43556 ( \43933 , \43925 , \43932 );
or \U$43557 ( \43934 , \43931 , \43924 );
nand \U$43558 ( \43935 , \43933 , \43934 );
xor \U$43559 ( \43936 , \43922 , \43935 );
xor \U$43560 ( \43937 , \43912 , \43936 );
not \U$43561 ( \43938 , \43937 );
or \U$43562 ( \43939 , \43871 , \43938 );
nand \U$43563 ( \43940 , \43912 , \43936 );
nand \U$43564 ( \43941 , \43939 , \43940 );
not \U$43565 ( \43942 , \43941 );
and \U$43566 ( \43943 , \43843 , \43942 );
not \U$43567 ( \43944 , \43843 );
and \U$43568 ( \43945 , \43944 , \43941 );
nor \U$43569 ( \43946 , \43943 , \43945 );
not \U$43570 ( \43947 , \43946 );
xor \U$43571 ( \43948 , \43736 , \43833 );
xor \U$43572 ( \43949 , \43948 , \43836 );
not \U$43573 ( \43950 , \14668 );
not \U$43574 ( \43951 , \43416 );
or \U$43575 ( \43952 , \43950 , \43951 );
nand \U$43576 ( \43953 , \43786 , RIae7aab0_192);
nand \U$43577 ( \43954 , \43952 , \43953 );
not \U$43578 ( \43955 , \43954 );
not \U$43579 ( \43956 , \9473 );
not \U$43580 ( \43957 , \43579 );
or \U$43581 ( \43958 , \43956 , \43957 );
nand \U$43582 ( \43959 , \43862 , \9705 );
nand \U$43583 ( \43960 , \43958 , \43959 );
not \U$43584 ( \43961 , \43960 );
not \U$43585 ( \43962 , \43961 );
not \U$43586 ( \43963 , \17847 );
not \U$43587 ( \43964 , \43395 );
or \U$43588 ( \43965 , \43963 , \43964 );
nand \U$43589 ( \43966 , \43901 , \10275 );
nand \U$43590 ( \43967 , \43965 , \43966 );
not \U$43591 ( \43968 , \43967 );
and \U$43592 ( \43969 , \43962 , \43968 );
and \U$43593 ( \43970 , \43967 , \43961 );
nor \U$43594 ( \43971 , \43969 , \43970 );
not \U$43595 ( \43972 , \43971 );
or \U$43596 ( \43973 , \43955 , \43972 );
or \U$43597 ( \43974 , \43971 , \43954 );
nand \U$43598 ( \43975 , \43973 , \43974 );
not \U$43599 ( \43976 , \43975 );
xnor \U$43600 ( \43977 , \43774 , \43764 );
not \U$43601 ( \43978 , \43977 );
not \U$43602 ( \43979 , \43420 );
not \U$43603 ( \43980 , \43410 );
or \U$43604 ( \43981 , \43979 , \43980 );
nand \U$43605 ( \43982 , \43981 , \43409 );
not \U$43606 ( \43983 , \43982 );
or \U$43607 ( \43984 , \43978 , \43983 );
or \U$43608 ( \43985 , \43982 , \43977 );
nand \U$43609 ( \43986 , \43984 , \43985 );
not \U$43610 ( \43987 , \43986 );
or \U$43611 ( \43988 , \43976 , \43987 );
not \U$43612 ( \43989 , \43977 );
nand \U$43613 ( \43990 , \43989 , \43982 );
nand \U$43614 ( \43991 , \43988 , \43990 );
not \U$43615 ( \43992 , \43991 );
not \U$43616 ( \43993 , \43778 );
and \U$43617 ( \43994 , \43829 , \43993 );
not \U$43618 ( \43995 , \43829 );
and \U$43619 ( \43996 , \43995 , \43778 );
nor \U$43620 ( \43997 , \43994 , \43996 );
not \U$43621 ( \43998 , \43997 );
xor \U$43622 ( \43999 , \43453 , \43459 );
and \U$43623 ( \44000 , \43999 , \43471 );
and \U$43624 ( \44001 , \43453 , \43459 );
or \U$43625 ( \44002 , \44000 , \44001 );
not \U$43626 ( \44003 , \44002 );
not \U$43627 ( \44004 , \10519 );
not \U$43628 ( \44005 , \43875 );
or \U$43629 ( \44006 , \44004 , \44005 );
nand \U$43630 ( \44007 , \43404 , \11439 );
nand \U$43631 ( \44008 , \44006 , \44007 );
not \U$43632 ( \44009 , \10695 );
not \U$43633 ( \44010 , \43487 );
or \U$43634 ( \44011 , \44009 , \44010 );
not \U$43635 ( \44012 , \10625 );
not \U$43636 ( \44013 , \36204 );
or \U$43637 ( \44014 , \44012 , \44013 );
nand \U$43638 ( \44015 , \10171 , RIae7a498_179);
nand \U$43639 ( \44016 , \44014 , \44015 );
nand \U$43640 ( \44017 , \44016 , \10675 );
nand \U$43641 ( \44018 , \44011 , \44017 );
not \U$43642 ( \44019 , \44018 );
not \U$43643 ( \44020 , \10667 );
not \U$43644 ( \44021 , \43477 );
or \U$43645 ( \44022 , \44020 , \44021 );
not \U$43646 ( \44023 , RIae7a150_172);
not \U$43647 ( \44024 , \10084 );
or \U$43648 ( \44025 , \44023 , \44024 );
nand \U$43649 ( \44026 , \38816 , \10672 );
nand \U$43650 ( \44027 , \44025 , \44026 );
nand \U$43651 ( \44028 , \44027 , \9776 );
nand \U$43652 ( \44029 , \44022 , \44028 );
not \U$43653 ( \44030 , \44029 );
not \U$43654 ( \44031 , \44030 );
or \U$43655 ( \44032 , \44019 , \44031 );
or \U$43656 ( \44033 , \44018 , \44030 );
nand \U$43657 ( \44034 , \44032 , \44033 );
xor \U$43658 ( \44035 , \44008 , \44034 );
not \U$43659 ( \44036 , \44035 );
or \U$43660 ( \44037 , \44003 , \44036 );
or \U$43661 ( \44038 , \44035 , \44002 );
not \U$43662 ( \44039 , \43584 );
not \U$43663 ( \44040 , \43572 );
or \U$43664 ( \44041 , \44039 , \44040 );
not \U$43665 ( \44042 , \43567 );
nand \U$43666 ( \44043 , \44042 , \43529 );
nand \U$43667 ( \44044 , \44041 , \44043 );
nand \U$43668 ( \44045 , \44038 , \44044 );
nand \U$43669 ( \44046 , \44037 , \44045 );
not \U$43670 ( \44047 , \44046 );
or \U$43671 ( \44048 , \43998 , \44047 );
or \U$43672 ( \44049 , \43997 , \44046 );
nand \U$43673 ( \44050 , \44048 , \44049 );
not \U$43674 ( \44051 , \44050 );
or \U$43675 ( \44052 , \43992 , \44051 );
not \U$43676 ( \44053 , \43997 );
nand \U$43677 ( \44054 , \44053 , \44046 );
nand \U$43678 ( \44055 , \44052 , \44054 );
xor \U$43679 ( \44056 , \43949 , \44055 );
not \U$43680 ( \44057 , \43555 );
not \U$43681 ( \44058 , \43565 );
or \U$43682 ( \44059 , \44057 , \44058 );
nand \U$43683 ( \44060 , \43554 , \43544 );
nand \U$43684 ( \44061 , \44059 , \44060 );
not \U$43685 ( \44062 , \44061 );
not \U$43686 ( \44063 , \44062 );
xor \U$43687 ( \44064 , \43879 , \43884 );
xor \U$43688 ( \44065 , \44064 , \43890 );
not \U$43689 ( \44066 , \44065 );
not \U$43690 ( \44067 , \44066 );
or \U$43691 ( \44068 , \44063 , \44067 );
not \U$43692 ( \44069 , \43481 );
not \U$43693 ( \44070 , \43491 );
or \U$43694 ( \44071 , \44069 , \44070 );
not \U$43695 ( \44072 , \43481 );
nand \U$43696 ( \44073 , \44072 , \43492 );
nand \U$43697 ( \44074 , \43503 , \44073 );
nand \U$43698 ( \44075 , \44071 , \44074 );
nand \U$43699 ( \44076 , \44068 , \44075 );
nand \U$43700 ( \44077 , \44065 , \44061 );
and \U$43701 ( \44078 , \44076 , \44077 );
not \U$43702 ( \44079 , \44078 );
not \U$43703 ( \44080 , \44079 );
xor \U$43704 ( \44081 , \43877 , \43907 );
not \U$43705 ( \44082 , \44081 );
or \U$43706 ( \44083 , \44080 , \44082 );
xor \U$43707 ( \44084 , \43877 , \44078 );
xnor \U$43708 ( \44085 , \44084 , \43907 );
xor \U$43709 ( \44086 , \43855 , \43865 );
nand \U$43710 ( \44087 , \44085 , \44086 );
nand \U$43711 ( \44088 , \44083 , \44087 );
and \U$43712 ( \44089 , \44056 , \44088 );
and \U$43713 ( \44090 , \43949 , \44055 );
or \U$43714 ( \44091 , \44089 , \44090 );
not \U$43715 ( \44092 , \44091 );
or \U$43716 ( \44093 , \43947 , \44092 );
or \U$43717 ( \44094 , \44091 , \43946 );
nand \U$43718 ( \44095 , \44093 , \44094 );
not \U$43719 ( \44096 , \9776 );
not \U$43720 ( \44097 , \43918 );
or \U$43721 ( \44098 , \44096 , \44097 );
nand \U$43722 ( \44099 , \44027 , \9758 );
nand \U$43723 ( \44100 , \44098 , \44099 );
not \U$43724 ( \44101 , \44100 );
not \U$43725 ( \44102 , \10676 );
and \U$43726 ( \44103 , RIae7a498_179, \10066 );
not \U$43727 ( \44104 , RIae7a498_179);
and \U$43728 ( \44105 , \44104 , \11230 );
nor \U$43729 ( \44106 , \44103 , \44105 );
not \U$43730 ( \44107 , \44106 );
or \U$43731 ( \44108 , \44102 , \44107 );
nand \U$43732 ( \44109 , \44016 , \10695 );
nand \U$43733 ( \44110 , \44108 , \44109 );
not \U$43734 ( \44111 , \44110 );
not \U$43735 ( \44112 , \16358 );
and \U$43736 ( \44113 , RIae7a510_180, \10750 );
not \U$43737 ( \44114 , RIae7a510_180);
and \U$43738 ( \44115 , \44114 , \9868 );
or \U$43739 ( \44116 , \44113 , \44115 );
not \U$43740 ( \44117 , \44116 );
or \U$43741 ( \44118 , \44112 , \44117 );
nand \U$43742 ( \44119 , \43741 , \10637 );
nand \U$43743 ( \44120 , \44118 , \44119 );
not \U$43744 ( \44121 , \44120 );
not \U$43745 ( \44122 , \44121 );
or \U$43746 ( \44123 , \44111 , \44122 );
or \U$43747 ( \44124 , \44121 , \44110 );
nand \U$43748 ( \44125 , \44123 , \44124 );
not \U$43749 ( \44126 , \44125 );
or \U$43750 ( \44127 , \44101 , \44126 );
nand \U$43751 ( \44128 , \44120 , \44110 );
nand \U$43752 ( \44129 , \44127 , \44128 );
not \U$43753 ( \44130 , \44129 );
not \U$43754 ( \44131 , \43803 );
not \U$43755 ( \44132 , \43824 );
or \U$43756 ( \44133 , \44131 , \44132 );
nand \U$43757 ( \44134 , \43819 , \43808 );
nand \U$43758 ( \44135 , \44133 , \44134 );
not \U$43759 ( \44136 , \44135 );
and \U$43760 ( \44137 , \44130 , \44136 );
not \U$43761 ( \44138 , \44130 );
and \U$43762 ( \44139 , \44138 , \44135 );
nor \U$43763 ( \44140 , \44137 , \44139 );
not \U$43764 ( \44141 , \44140 );
not \U$43765 ( \44142 , \11400 );
not \U$43766 ( \44143 , \44116 );
or \U$43767 ( \44144 , \44142 , \44143 );
nand \U$43768 ( \44145 , \40625 , \10631 );
nand \U$43769 ( \44146 , \44144 , \44145 );
not \U$43770 ( \44147 , \44146 );
not \U$43771 ( \44148 , \16564 );
not \U$43772 ( \44149 , \44106 );
or \U$43773 ( \44150 , \44148 , \44149 );
nand \U$43774 ( \44151 , \40674 , \11422 );
nand \U$43775 ( \44152 , \44150 , \44151 );
not \U$43776 ( \44153 , \44152 );
not \U$43777 ( \44154 , \44153 );
or \U$43778 ( \44155 , \44147 , \44154 );
or \U$43779 ( \44156 , \44153 , \44146 );
nand \U$43780 ( \44157 , \44155 , \44156 );
not \U$43781 ( \44158 , \9478 );
xnor \U$43782 ( \44159 , RIae7a6f0_184, \25333 );
not \U$43783 ( \44160 , \44159 );
or \U$43784 ( \44161 , \44158 , \44160 );
nand \U$43785 ( \44162 , \43856 , \9473 );
nand \U$43786 ( \44163 , \44161 , \44162 );
xor \U$43787 ( \44164 , \44157 , \44163 );
not \U$43788 ( \44165 , \44164 );
or \U$43789 ( \44166 , \44141 , \44165 );
nand \U$43790 ( \44167 , \44129 , \44135 );
nand \U$43791 ( \44168 , \44166 , \44167 );
not \U$43792 ( \44169 , \43717 );
not \U$43793 ( \44170 , \43711 );
or \U$43794 ( \44171 , \44169 , \44170 );
not \U$43795 ( \44172 , \43718 );
not \U$43796 ( \44173 , \43710 );
or \U$43797 ( \44174 , \44172 , \44173 );
nand \U$43798 ( \44175 , \44174 , \43734 );
nand \U$43799 ( \44176 , \44171 , \44175 );
not \U$43800 ( \44177 , \44176 );
not \U$43801 ( \44178 , \44157 );
not \U$43802 ( \44179 , \44163 );
or \U$43803 ( \44180 , \44178 , \44179 );
nand \U$43804 ( \44181 , \44152 , \44146 );
nand \U$43805 ( \44182 , \44180 , \44181 );
and \U$43806 ( \44183 , \44177 , \44182 );
not \U$43807 ( \44184 , \44177 );
not \U$43808 ( \44185 , \44182 );
and \U$43809 ( \44186 , \44184 , \44185 );
nor \U$43810 ( \44187 , \44183 , \44186 );
not \U$43811 ( \44188 , \44187 );
xnor \U$43812 ( \44189 , \40550 , \40477 );
not \U$43813 ( \44190 , \44189 );
and \U$43814 ( \44191 , \44188 , \44190 );
and \U$43815 ( \44192 , \44187 , \44189 );
nor \U$43816 ( \44193 , \44191 , \44192 );
xor \U$43817 ( \44194 , \44168 , \44193 );
and \U$43818 ( \44195 , \43922 , \43935 );
and \U$43819 ( \44196 , \43930 , \43924 );
nor \U$43820 ( \44197 , \44195 , \44196 );
not \U$43821 ( \44198 , \40574 );
and \U$43822 ( \44199 , \40565 , \44198 );
not \U$43823 ( \44200 , \40565 );
and \U$43824 ( \44201 , \44200 , \40574 );
nor \U$43825 ( \44202 , \44199 , \44201 );
xnor \U$43826 ( \44203 , \40584 , \44202 );
xor \U$43827 ( \44204 , \44197 , \44203 );
xor \U$43828 ( \44205 , \40246 , \40256 );
xor \U$43829 ( \44206 , \44205 , \40265 );
not \U$43830 ( \44207 , \44206 );
not \U$43831 ( \44208 , \17507 );
not \U$43832 ( \44209 , \40351 );
or \U$43833 ( \44210 , \44208 , \44209 );
nand \U$43834 ( \44211 , \44159 , \9473 );
nand \U$43835 ( \44212 , \44210 , \44211 );
and \U$43836 ( \44213 , \44207 , \44212 );
not \U$43837 ( \44214 , \44207 );
not \U$43838 ( \44215 , \44212 );
and \U$43839 ( \44216 , \44214 , \44215 );
or \U$43840 ( \44217 , \44213 , \44216 );
xnor \U$43841 ( \44218 , \44204 , \44217 );
buf \U$43842 ( \44219 , \44218 );
xnor \U$43843 ( \44220 , \44194 , \44219 );
not \U$43844 ( \44221 , \44008 );
not \U$43845 ( \44222 , \44034 );
or \U$43846 ( \44223 , \44221 , \44222 );
nand \U$43847 ( \44224 , \44029 , \44018 );
nand \U$43848 ( \44225 , \44223 , \44224 );
xor \U$43849 ( \44226 , \44125 , \44100 );
xor \U$43850 ( \44227 , \44225 , \44226 );
not \U$43851 ( \44228 , \44227 );
not \U$43852 ( \44229 , \43954 );
not \U$43853 ( \44230 , \43971 );
not \U$43854 ( \44231 , \44230 );
or \U$43855 ( \44232 , \44229 , \44231 );
nand \U$43856 ( \44233 , \43960 , \43967 );
nand \U$43857 ( \44234 , \44232 , \44233 );
not \U$43858 ( \44235 , \44234 );
or \U$43859 ( \44236 , \44228 , \44235 );
nand \U$43860 ( \44237 , \44225 , \44226 );
nand \U$43861 ( \44238 , \44236 , \44237 );
not \U$43862 ( \44239 , \44238 );
and \U$43863 ( \44240 , \44140 , \44164 );
not \U$43864 ( \44241 , \44140 );
not \U$43865 ( \44242 , \44164 );
and \U$43866 ( \44243 , \44241 , \44242 );
nor \U$43867 ( \44244 , \44240 , \44243 );
not \U$43868 ( \44245 , \44244 );
nand \U$43869 ( \44246 , \44239 , \44245 );
not \U$43870 ( \44247 , \44246 );
xor \U$43871 ( \44248 , \43936 , \43869 );
xnor \U$43872 ( \44249 , \44248 , \43912 );
not \U$43873 ( \44250 , \44249 );
or \U$43874 ( \44251 , \44247 , \44250 );
nand \U$43875 ( \44252 , \44238 , \44244 );
nand \U$43876 ( \44253 , \44251 , \44252 );
not \U$43877 ( \44254 , \44253 );
and \U$43878 ( \44255 , \44220 , \44254 );
not \U$43879 ( \44256 , \44220 );
and \U$43880 ( \44257 , \44256 , \44253 );
nor \U$43881 ( \44258 , \44255 , \44257 );
xnor \U$43882 ( \44259 , \44095 , \44258 );
not \U$43883 ( \44260 , \44259 );
xnor \U$43884 ( \44261 , \44234 , \44227 );
xnor \U$43885 ( \44262 , \43991 , \44050 );
xor \U$43886 ( \44263 , \44261 , \44262 );
not \U$43887 ( \44264 , \44086 );
and \U$43888 ( \44265 , \44085 , \44264 );
not \U$43889 ( \44266 , \44085 );
and \U$43890 ( \44267 , \44266 , \44086 );
nor \U$43891 ( \44268 , \44265 , \44267 );
and \U$43892 ( \44269 , \44263 , \44268 );
and \U$43893 ( \44270 , \44261 , \44262 );
or \U$43894 ( \44271 , \44269 , \44270 );
not \U$43895 ( \44272 , \44271 );
and \U$43896 ( \44273 , \44238 , \44244 );
not \U$43897 ( \44274 , \44238 );
and \U$43898 ( \44275 , \44274 , \44245 );
nor \U$43899 ( \44276 , \44273 , \44275 );
xor \U$43900 ( \44277 , \44249 , \44276 );
xor \U$43901 ( \44278 , \43949 , \44055 );
xor \U$43902 ( \44279 , \44278 , \44088 );
xor \U$43903 ( \44280 , \44277 , \44279 );
not \U$43904 ( \44281 , \44280 );
or \U$43905 ( \44282 , \44272 , \44281 );
or \U$43906 ( \44283 , \44279 , \44277 );
nand \U$43907 ( \44284 , \44282 , \44283 );
nand \U$43908 ( \44285 , \44260 , \44284 );
not \U$43909 ( \44286 , \44271 );
xor \U$43910 ( \44287 , \44277 , \44286 );
xnor \U$43911 ( \44288 , \44287 , \44279 );
not \U$43912 ( \44289 , \43472 );
nand \U$43913 ( \44290 , \44289 , \43508 );
not \U$43914 ( \44291 , \44290 );
not \U$43915 ( \44292 , \43516 );
or \U$43916 ( \44293 , \44291 , \44292 );
nand \U$43917 ( \44294 , \43509 , \43472 );
nand \U$43918 ( \44295 , \44293 , \44294 );
not \U$43919 ( \44296 , \44061 );
not \U$43920 ( \44297 , \44066 );
or \U$43921 ( \44298 , \44296 , \44297 );
nand \U$43922 ( \44299 , \44065 , \44062 );
nand \U$43923 ( \44300 , \44298 , \44299 );
xor \U$43924 ( \44301 , \44075 , \44300 );
nand \U$43925 ( \44302 , \44295 , \44301 );
not \U$43926 ( \44303 , \44302 );
not \U$43927 ( \44304 , \43986 );
not \U$43928 ( \44305 , \43975 );
not \U$43929 ( \44306 , \44305 );
and \U$43930 ( \44307 , \44304 , \44306 );
and \U$43931 ( \44308 , \43986 , \44305 );
nor \U$43932 ( \44309 , \44307 , \44308 );
not \U$43933 ( \44310 , \44309 );
or \U$43934 ( \44311 , \44303 , \44310 );
nor \U$43935 ( \44312 , \44295 , \44301 );
not \U$43936 ( \44313 , \44312 );
nand \U$43937 ( \44314 , \44311 , \44313 );
not \U$43938 ( \44315 , \43597 );
not \U$43939 ( \44316 , \43521 );
nand \U$43940 ( \44317 , \44316 , \43589 );
not \U$43941 ( \44318 , \44317 );
or \U$43942 ( \44319 , \44315 , \44318 );
nand \U$43943 ( \44320 , \43590 , \43521 );
nand \U$43944 ( \44321 , \44319 , \44320 );
not \U$43945 ( \44322 , \44321 );
xor \U$43946 ( \44323 , \44002 , \44035 );
xnor \U$43947 ( \44324 , \44323 , \44044 );
not \U$43948 ( \44325 , \44324 );
not \U$43949 ( \44326 , \44325 );
or \U$43950 ( \44327 , \44322 , \44326 );
not \U$43951 ( \44328 , \44324 );
not \U$43952 ( \44329 , \44321 );
not \U$43953 ( \44330 , \44329 );
or \U$43954 ( \44331 , \44328 , \44330 );
not \U$43955 ( \44332 , \43427 );
not \U$43956 ( \44333 , \43432 );
or \U$43957 ( \44334 , \44332 , \44333 );
nand \U$43958 ( \44335 , \44334 , \43426 );
nand \U$43959 ( \44336 , \44331 , \44335 );
nand \U$43960 ( \44337 , \44327 , \44336 );
not \U$43961 ( \44338 , \44337 );
nor \U$43962 ( \44339 , \44314 , \44338 );
not \U$43963 ( \44340 , \44339 );
not \U$43964 ( \44341 , \44340 );
xor \U$43965 ( \44342 , \44261 , \44262 );
xor \U$43966 ( \44343 , \44342 , \44268 );
not \U$43967 ( \44344 , \44343 );
or \U$43968 ( \44345 , \44341 , \44344 );
nand \U$43969 ( \44346 , \44314 , \44338 );
nand \U$43970 ( \44347 , \44345 , \44346 );
nand \U$43971 ( \44348 , \44288 , \44347 );
not \U$43972 ( \44349 , \44339 );
nand \U$43973 ( \44350 , \44349 , \44346 );
not \U$43974 ( \44351 , \44350 );
not \U$43975 ( \44352 , \44343 );
or \U$43976 ( \44353 , \44351 , \44352 );
or \U$43977 ( \44354 , \44343 , \44350 );
nand \U$43978 ( \44355 , \44353 , \44354 );
xor \U$43979 ( \44356 , \43517 , \43598 );
and \U$43980 ( \44357 , \44356 , \43607 );
and \U$43981 ( \44358 , \43517 , \43598 );
or \U$43982 ( \44359 , \44357 , \44358 );
not \U$43983 ( \44360 , \44359 );
not \U$43984 ( \44361 , \44312 );
nand \U$43985 ( \44362 , \44361 , \44302 );
not \U$43986 ( \44363 , \44362 );
not \U$43987 ( \44364 , \44309 );
and \U$43988 ( \44365 , \44363 , \44364 );
and \U$43989 ( \44366 , \44309 , \44362 );
nor \U$43990 ( \44367 , \44365 , \44366 );
not \U$43991 ( \44368 , \44367 );
not \U$43992 ( \44369 , \44321 );
not \U$43993 ( \44370 , \44324 );
or \U$43994 ( \44371 , \44369 , \44370 );
or \U$43995 ( \44372 , \44321 , \44324 );
nand \U$43996 ( \44373 , \44371 , \44372 );
not \U$43997 ( \44374 , \44335 );
and \U$43998 ( \44375 , \44373 , \44374 );
not \U$43999 ( \44376 , \44373 );
and \U$44000 ( \44377 , \44376 , \44335 );
nor \U$44001 ( \44378 , \44375 , \44377 );
not \U$44002 ( \44379 , \44378 );
or \U$44003 ( \44380 , \44368 , \44379 );
or \U$44004 ( \44381 , \44378 , \44367 );
nand \U$44005 ( \44382 , \44380 , \44381 );
not \U$44006 ( \44383 , \44382 );
or \U$44007 ( \44384 , \44360 , \44383 );
not \U$44008 ( \44385 , \44367 );
nand \U$44009 ( \44386 , \44385 , \44378 );
nand \U$44010 ( \44387 , \44384 , \44386 );
nand \U$44011 ( \44388 , \44355 , \44387 );
not \U$44012 ( \44389 , \44359 );
not \U$44013 ( \44390 , \44382 );
not \U$44014 ( \44391 , \44390 );
or \U$44015 ( \44392 , \44389 , \44391 );
or \U$44016 ( \44393 , \44390 , \44359 );
nand \U$44017 ( \44394 , \44392 , \44393 );
xor \U$44018 ( \44395 , \43437 , \43441 );
and \U$44019 ( \44396 , \44395 , \43608 );
and \U$44020 ( \44397 , \43437 , \43441 );
or \U$44021 ( \44398 , \44396 , \44397 );
nand \U$44022 ( \44399 , \44394 , \44398 );
and \U$44023 ( \44400 , \44388 , \44399 );
and \U$44024 ( \44401 , \44285 , \44348 , \44400 );
nand \U$44025 ( \44402 , \43627 , \44401 );
not \U$44026 ( \44403 , \44348 );
not \U$44027 ( \44404 , \44388 );
nor \U$44028 ( \44405 , \44394 , \44398 );
not \U$44029 ( \44406 , \44405 );
or \U$44030 ( \44407 , \44404 , \44406 );
not \U$44031 ( \44408 , \44355 );
not \U$44032 ( \44409 , \44387 );
nand \U$44033 ( \44410 , \44408 , \44409 );
nand \U$44034 ( \44411 , \44407 , \44410 );
not \U$44035 ( \44412 , \44411 );
or \U$44036 ( \44413 , \44403 , \44412 );
not \U$44037 ( \44414 , \44288 );
not \U$44038 ( \44415 , \44347 );
nand \U$44039 ( \44416 , \44414 , \44415 );
nand \U$44040 ( \44417 , \44413 , \44416 );
nand \U$44041 ( \44418 , \44417 , \44285 );
not \U$44042 ( \44419 , \44284 );
nand \U$44043 ( \44420 , \44419 , \44259 );
nand \U$44044 ( \44421 , \44402 , \44418 , \44420 );
xor \U$44045 ( \44422 , \40468 , \40470 );
xor \U$44046 ( \44423 , \44422 , \40702 );
not \U$44047 ( \44424 , \40685 );
not \U$44048 ( \44425 , \40632 );
not \U$44049 ( \44426 , \44425 );
and \U$44050 ( \44427 , \44424 , \44426 );
and \U$44051 ( \44428 , \40685 , \44425 );
nor \U$44052 ( \44429 , \44427 , \44428 );
not \U$44053 ( \44430 , \43699 );
not \U$44054 ( \44431 , \43638 );
or \U$44055 ( \44432 , \44430 , \44431 );
not \U$44056 ( \44433 , \43632 );
nand \U$44057 ( \44434 , \44433 , \43634 );
nand \U$44058 ( \44435 , \44432 , \44434 );
not \U$44059 ( \44436 , \44435 );
xor \U$44060 ( \44437 , \44429 , \44436 );
not \U$44061 ( \44438 , \44215 );
not \U$44062 ( \44439 , \44207 );
and \U$44063 ( \44440 , \44438 , \44439 );
not \U$44064 ( \44441 , \44197 );
and \U$44065 ( \44442 , \44217 , \44441 );
nor \U$44066 ( \44443 , \44440 , \44442 );
and \U$44067 ( \44444 , \44437 , \44443 );
and \U$44068 ( \44445 , \44429 , \44436 );
or \U$44069 ( \44446 , \44444 , \44445 );
not \U$44070 ( \44447 , \44446 );
not \U$44071 ( \44448 , \40700 );
and \U$44072 ( \44449 , \40698 , \44448 );
not \U$44073 ( \44450 , \40698 );
and \U$44074 ( \44451 , \44450 , \40700 );
nor \U$44075 ( \44452 , \44449 , \44451 );
not \U$44076 ( \44453 , \44452 );
or \U$44077 ( \44454 , \44447 , \44453 );
xor \U$44078 ( \44455 , \40444 , \40466 );
xnor \U$44079 ( \44456 , \44455 , \40463 );
nand \U$44080 ( \44457 , \44454 , \44456 );
not \U$44081 ( \44458 , \44446 );
not \U$44082 ( \44459 , \44452 );
nand \U$44083 ( \44460 , \44458 , \44459 );
and \U$44084 ( \44461 , \44457 , \44460 );
not \U$44085 ( \44462 , \40412 );
not \U$44086 ( \44463 , \40392 );
or \U$44087 ( \44464 , \44462 , \44463 );
or \U$44088 ( \44465 , \40392 , \40412 );
nand \U$44089 ( \44466 , \44464 , \44465 );
and \U$44090 ( \44467 , \44466 , \40384 );
not \U$44091 ( \44468 , \44466 );
and \U$44092 ( \44469 , \44468 , \40383 );
nor \U$44093 ( \44470 , \44467 , \44469 );
not \U$44094 ( \44471 , \44470 );
and \U$44095 ( \44472 , \44461 , \44471 );
not \U$44096 ( \44473 , \44461 );
and \U$44097 ( \44474 , \44473 , \44470 );
nor \U$44098 ( \44475 , \44472 , \44474 );
xnor \U$44099 ( \44476 , \44423 , \44475 );
not \U$44100 ( \44477 , \44189 );
nand \U$44101 ( \44478 , \44477 , \44182 );
not \U$44102 ( \44479 , \44185 );
not \U$44103 ( \44480 , \44189 );
or \U$44104 ( \44481 , \44479 , \44480 );
nand \U$44105 ( \44482 , \44481 , \44177 );
nand \U$44106 ( \44483 , \44478 , \44482 );
not \U$44107 ( \44484 , \40554 );
not \U$44108 ( \44485 , \44484 );
not \U$44109 ( \44486 , \40597 );
or \U$44110 ( \44487 , \44485 , \44486 );
or \U$44111 ( \44488 , \40597 , \44484 );
nand \U$44112 ( \44489 , \44487 , \44488 );
xor \U$44113 ( \44490 , \44483 , \44489 );
not \U$44114 ( \44491 , \40446 );
not \U$44115 ( \44492 , \40450 );
or \U$44116 ( \44493 , \44491 , \44492 );
nand \U$44117 ( \44494 , \40447 , \40449 );
nand \U$44118 ( \44495 , \44493 , \44494 );
xnor \U$44119 ( \44496 , \44495 , \40457 );
and \U$44120 ( \44497 , \44490 , \44496 );
and \U$44121 ( \44498 , \44483 , \44489 );
or \U$44122 ( \44499 , \44497 , \44498 );
not \U$44123 ( \44500 , \44499 );
not \U$44124 ( \44501 , \43700 );
not \U$44125 ( \44502 , \44501 );
not \U$44126 ( \44503 , \43839 );
or \U$44127 ( \44504 , \44502 , \44503 );
nand \U$44128 ( \44505 , \43843 , \43941 );
nand \U$44129 ( \44506 , \44504 , \44505 );
not \U$44130 ( \44507 , \44506 );
xor \U$44131 ( \44508 , \44429 , \44436 );
xor \U$44132 ( \44509 , \44508 , \44443 );
not \U$44133 ( \44510 , \44509 );
not \U$44134 ( \44511 , \44168 );
not \U$44135 ( \44512 , \44218 );
or \U$44136 ( \44513 , \44511 , \44512 );
and \U$44137 ( \44514 , \44217 , \44197 );
not \U$44138 ( \44515 , \44217 );
and \U$44139 ( \44516 , \44515 , \44441 );
or \U$44140 ( \44517 , \44514 , \44516 );
nand \U$44141 ( \44518 , \44517 , \44203 );
nand \U$44142 ( \44519 , \44513 , \44518 );
not \U$44143 ( \44520 , \44519 );
or \U$44144 ( \44521 , \44510 , \44520 );
or \U$44145 ( \44522 , \44519 , \44509 );
nand \U$44146 ( \44523 , \44521 , \44522 );
not \U$44147 ( \44524 , \44523 );
or \U$44148 ( \44525 , \44507 , \44524 );
not \U$44149 ( \44526 , \44509 );
nand \U$44150 ( \44527 , \44526 , \44519 );
nand \U$44151 ( \44528 , \44525 , \44527 );
not \U$44152 ( \44529 , \44528 );
or \U$44153 ( \44530 , \44500 , \44529 );
xor \U$44154 ( \44531 , \44446 , \44459 );
xnor \U$44155 ( \44532 , \44531 , \44456 );
not \U$44156 ( \44533 , \44532 );
nand \U$44157 ( \44534 , \44530 , \44533 );
or \U$44158 ( \44535 , \44528 , \44499 );
nand \U$44159 ( \44536 , \44534 , \44535 );
nand \U$44160 ( \44537 , \44476 , \44536 );
not \U$44161 ( \44538 , \44423 );
nand \U$44162 ( \44539 , \44538 , \44475 );
not \U$44163 ( \44540 , \44539 );
nand \U$44164 ( \44541 , \44461 , \44471 );
not \U$44165 ( \44542 , \44541 );
or \U$44166 ( \44543 , \44540 , \44542 );
xor \U$44167 ( \44544 , \40707 , \40705 );
not \U$44168 ( \44545 , \44544 );
not \U$44169 ( \44546 , \40710 );
or \U$44170 ( \44547 , \44545 , \44546 );
or \U$44171 ( \44548 , \40710 , \44544 );
nand \U$44172 ( \44549 , \44547 , \44548 );
nand \U$44173 ( \44550 , \44543 , \44549 );
and \U$44174 ( \44551 , \44537 , \44550 );
xor \U$44175 ( \44552 , \44483 , \44489 );
xor \U$44176 ( \44553 , \44552 , \44496 );
nand \U$44177 ( \44554 , \44220 , \44253 );
not \U$44178 ( \44555 , \44168 );
buf \U$44179 ( \44556 , \44219 );
nand \U$44180 ( \44557 , \44555 , \44556 );
not \U$44181 ( \44558 , \44557 );
not \U$44182 ( \44559 , \44556 );
nand \U$44183 ( \44560 , \44559 , \44168 );
not \U$44184 ( \44561 , \44560 );
or \U$44185 ( \44562 , \44558 , \44561 );
not \U$44186 ( \44563 , \44193 );
nand \U$44187 ( \44564 , \44562 , \44563 );
nand \U$44188 ( \44565 , \44554 , \44564 );
xor \U$44189 ( \44566 , \44553 , \44565 );
not \U$44190 ( \44567 , \44506 );
and \U$44191 ( \44568 , \44523 , \44567 );
not \U$44192 ( \44569 , \44523 );
and \U$44193 ( \44570 , \44569 , \44506 );
nor \U$44194 ( \44571 , \44568 , \44570 );
xnor \U$44195 ( \44572 , \44566 , \44571 );
not \U$44196 ( \44573 , \44572 );
nand \U$44197 ( \44574 , \44258 , \43946 );
and \U$44198 ( \44575 , \44574 , \44091 );
nor \U$44199 ( \44576 , \44258 , \43946 );
nor \U$44200 ( \44577 , \44575 , \44576 );
nand \U$44201 ( \44578 , \44573 , \44577 );
xor \U$44202 ( \44579 , \44499 , \44528 );
xor \U$44203 ( \44580 , \44579 , \44532 );
not \U$44204 ( \44581 , \44553 );
not \U$44205 ( \44582 , \44565 );
or \U$44206 ( \44583 , \44581 , \44582 );
nand \U$44207 ( \44584 , \44583 , \44571 );
not \U$44208 ( \44585 , \44553 );
nand \U$44209 ( \44586 , \44585 , \44564 , \44554 );
and \U$44210 ( \44587 , \44584 , \44586 );
nor \U$44211 ( \44588 , \44580 , \44587 );
not \U$44212 ( \44589 , \44588 );
and \U$44213 ( \44590 , \44551 , \44578 , \44589 );
nand \U$44214 ( \44591 , \44421 , \44590 );
buf \U$44215 ( \44592 , \44537 );
not \U$44216 ( \44593 , \44592 );
not \U$44217 ( \44594 , \44577 );
nand \U$44218 ( \44595 , \44594 , \44572 );
or \U$44219 ( \44596 , \44595 , \44588 );
nand \U$44220 ( \44597 , \44580 , \44587 );
nand \U$44221 ( \44598 , \44596 , \44597 );
not \U$44222 ( \44599 , \44598 );
or \U$44223 ( \44600 , \44593 , \44599 );
or \U$44224 ( \44601 , \44536 , \44476 );
nand \U$44225 ( \44602 , \44600 , \44601 );
nand \U$44226 ( \44603 , \44602 , \44550 );
not \U$44227 ( \44604 , \44549 );
nand \U$44228 ( \44605 , \44539 , \44604 , \44541 );
nand \U$44229 ( \44606 , \44591 , \44603 , \44605 );
and \U$44230 ( \44607 , \37027 , \40835 , \44606 );
nor \U$44231 ( \44608 , \40827 , \44607 );
nand \U$44232 ( \44609 , \40814 , \44608 );
nand \U$44233 ( \44610 , \34302 , \34301 );
not \U$44234 ( \44611 , \44610 );
nor \U$44235 ( \44612 , \34340 , \34312 );
nor \U$44236 ( \44613 , \44611 , \44612 );
and \U$44237 ( \44614 , \44613 , \34366 , \34305 );
and \U$44238 ( \44615 , \32278 , \32280 );
nand \U$44239 ( \44616 , \44614 , \44615 , \32287 );
nor \U$44240 ( \44617 , \44616 , \35451 );
nand \U$44241 ( \44618 , \44609 , \44617 , \35662 );
nor \U$44242 ( \44619 , \35620 , \35642 );
not \U$44243 ( \44620 , \44619 );
not \U$44244 ( \44621 , \35661 );
or \U$44245 ( \44622 , \44620 , \44621 );
not \U$44246 ( \44623 , \35660 );
not \U$44247 ( \44624 , \35654 );
nand \U$44248 ( \44625 , \44623 , \44624 );
nand \U$44249 ( \44626 , \44622 , \44625 );
nor \U$44250 ( \44627 , \35557 , \35613 );
or \U$44251 ( \44628 , \44626 , \44627 );
and \U$44252 ( \44629 , \35614 , \35652 );
nand \U$44253 ( \44630 , \44628 , \44629 );
or \U$44254 ( \44631 , \35649 , \35651 );
nand \U$44255 ( \44632 , \44630 , \44631 );
not \U$44256 ( \44633 , \44632 );
nand \U$44257 ( \44634 , \35663 , \44618 , \44633 );
nand \U$44258 ( \44635 , \22818 , \27525 , \44634 );
nand \U$44259 ( \44636 , \20771 , \20691 );
nor \U$44260 ( \44637 , \44636 , \20760 );
not \U$44261 ( \44638 , \44637 );
not \U$44262 ( \44639 , \20569 );
nor \U$44263 ( \44640 , \20265 , \20587 );
not \U$44264 ( \44641 , \44640 );
nand \U$44265 ( \44642 , \19549 , \19970 );
nand \U$44266 ( \44643 , \20264 , \20257 );
nand \U$44267 ( \44644 , \44642 , \44643 );
not \U$44268 ( \44645 , \44644 );
or \U$44269 ( \44646 , \44641 , \44645 );
buf \U$44270 ( \44647 , \20579 );
buf \U$44271 ( \44648 , \20586 );
nand \U$44272 ( \44649 , \44647 , \44648 );
nand \U$44273 ( \44650 , \44646 , \44649 );
not \U$44274 ( \44651 , \44650 );
or \U$44275 ( \44652 , \44639 , \44651 );
or \U$44276 ( \44653 , \20546 , \20568 );
nand \U$44277 ( \44654 , \44652 , \44653 );
not \U$44278 ( \44655 , \44654 );
or \U$44279 ( \44656 , \44638 , \44655 );
not \U$44280 ( \44657 , \20591 );
not \U$44281 ( \44658 , \20690 );
and \U$44282 ( \44659 , \44657 , \44658 );
nor \U$44283 ( \44660 , \20763 , \20770 );
nor \U$44284 ( \44661 , \44659 , \44660 );
not \U$44285 ( \44662 , \20691 );
nor \U$44286 ( \44663 , \44661 , \44662 );
nor \U$44287 ( \44664 , \20723 , \20727 );
not \U$44288 ( \44665 , \44664 );
not \U$44289 ( \44666 , \20759 );
or \U$44290 ( \44667 , \44665 , \44666 );
not \U$44291 ( \44668 , \20751 );
not \U$44292 ( \44669 , \20758 );
nand \U$44293 ( \44670 , \44668 , \44669 );
nand \U$44294 ( \44671 , \44667 , \44670 );
not \U$44295 ( \44672 , \44671 );
nor \U$44296 ( \44673 , \44672 , \44636 );
nor \U$44297 ( \44674 , \44663 , \44673 );
nand \U$44298 ( \44675 , \44656 , \44674 );
not \U$44299 ( \44676 , \44675 );
nor \U$44300 ( \44677 , \22815 , \15930 );
not \U$44301 ( \44678 , \44677 );
or \U$44302 ( \44679 , \44676 , \44678 );
not \U$44303 ( \44680 , \22803 );
not \U$44304 ( \44681 , \22813 );
buf \U$44305 ( \44682 , \20780 );
not \U$44306 ( \44683 , \21305 );
nand \U$44307 ( \44684 , \44682 , \44683 );
or \U$44308 ( \44685 , \44681 , \44684 );
or \U$44309 ( \44686 , \22811 , \22812 );
buf \U$44310 ( \44687 , \21824 );
buf \U$44311 ( \44688 , \22304 );
nand \U$44312 ( \44689 , \44687 , \44688 );
nand \U$44313 ( \44690 , \44685 , \44686 , \44689 );
not \U$44314 ( \44691 , \44690 );
or \U$44315 ( \44692 , \44680 , \44691 );
and \U$44316 ( \44693 , \15919 , \15929 );
nand \U$44317 ( \44694 , \14222 , \14882 );
nand \U$44318 ( \44695 , \13617 , \14219 );
and \U$44319 ( \44696 , \44694 , \44695 );
nor \U$44320 ( \44697 , \44696 , \14220 );
nand \U$44321 ( \44698 , \22814 , \44693 , \44697 );
nand \U$44322 ( \44699 , \44692 , \44698 );
not \U$44323 ( \44700 , \15919 );
not \U$44324 ( \44701 , \15925 );
nor \U$44325 ( \44702 , \44701 , \15928 );
not \U$44326 ( \44703 , \44702 );
or \U$44327 ( \44704 , \44700 , \44703 );
or \U$44328 ( \44705 , \15905 , \15918 );
nand \U$44329 ( \44706 , \44704 , \44705 );
not \U$44330 ( \44707 , \44706 );
not \U$44331 ( \44708 , \22814 );
or \U$44332 ( \44709 , \44707 , \44708 );
not \U$44333 ( \44710 , \22794 );
nand \U$44334 ( \44711 , \22294 , \22299 );
nand \U$44335 ( \44712 , \44710 , \44711 , \22799 );
nand \U$44336 ( \44713 , \44709 , \44712 );
nor \U$44337 ( \44714 , \44699 , \44713 );
nand \U$44338 ( \44715 , \44679 , \44714 );
nand \U$44339 ( \44716 , \44715 , \27525 );
and \U$44340 ( \44717 , \24218 , \24175 );
and \U$44341 ( \44718 , \44717 , \27524 , \24246 , \24260 );
not \U$44342 ( \44719 , \44718 );
nor \U$44343 ( \44720 , \25677 , \26086 );
nand \U$44344 ( \44721 , \26907 , \27287 , \44720 );
or \U$44345 ( \44722 , \27128 , \27276 );
nand \U$44346 ( \44723 , \44721 , \44722 );
not \U$44347 ( \44724 , \26864 );
not \U$44348 ( \44725 , \26893 );
or \U$44349 ( \44726 , \44724 , \44725 );
nor \U$44350 ( \44727 , \26900 , \26904 );
nand \U$44351 ( \44728 , \44726 , \44727 );
not \U$44352 ( \44729 , \26893 );
not \U$44353 ( \44730 , \26864 );
nand \U$44354 ( \44731 , \44729 , \44730 );
nand \U$44355 ( \44732 , \44728 , \44731 );
not \U$44356 ( \44733 , \44732 );
not \U$44357 ( \44734 , \27287 );
or \U$44358 ( \44735 , \44733 , \44734 );
buf \U$44359 ( \44736 , \27284 );
nor \U$44360 ( \44737 , \44736 , \27281 );
buf \U$44361 ( \44738 , \27277 );
nand \U$44362 ( \44739 , \44737 , \44738 );
nand \U$44363 ( \44740 , \44735 , \44739 );
nor \U$44364 ( \44741 , \44723 , \44740 );
not \U$44365 ( \44742 , \25648 );
nand \U$44366 ( \44743 , \26098 , \26091 );
not \U$44367 ( \44744 , \44743 );
nand \U$44368 ( \44745 , \44744 , \25671 );
not \U$44369 ( \44746 , \25649 );
not \U$44370 ( \44747 , \25670 );
nand \U$44371 ( \44748 , \44746 , \25651 , \44747 );
nand \U$44372 ( \44749 , \44745 , \44748 );
not \U$44373 ( \44750 , \44749 );
or \U$44374 ( \44751 , \44742 , \44750 );
or \U$44375 ( \44752 , \25647 , \25203 );
nand \U$44376 ( \44753 , \44751 , \44752 );
nor \U$44377 ( \44754 , \26906 , \27286 );
buf \U$44378 ( \44755 , \26087 );
nand \U$44379 ( \44756 , \44753 , \44754 , \44755 );
nand \U$44380 ( \44757 , \44741 , \44756 );
not \U$44381 ( \44758 , \44757 );
or \U$44382 ( \44759 , \44719 , \44758 );
not \U$44383 ( \44760 , \27459 );
nor \U$44384 ( \44761 , \27466 , \27465 );
not \U$44385 ( \44762 , \44761 );
or \U$44386 ( \44763 , \44760 , \44762 );
or \U$44387 ( \44764 , \27432 , \27458 );
nand \U$44388 ( \44765 , \44763 , \44764 );
nor \U$44389 ( \44766 , \27514 , \27521 );
nor \U$44390 ( \44767 , \44765 , \44766 );
not \U$44391 ( \44768 , \27502 );
not \U$44392 ( \44769 , \27506 );
or \U$44393 ( \44770 , \44768 , \44769 );
nand \U$44394 ( \44771 , \44770 , \27522 );
or \U$44395 ( \44772 , \44767 , \44771 );
or \U$44396 ( \44773 , \27502 , \27506 );
nand \U$44397 ( \44774 , \44772 , \44773 );
and \U$44398 ( \44775 , \44774 , \24261 );
not \U$44399 ( \44776 , \24260 );
not \U$44400 ( \44777 , \24246 );
nor \U$44401 ( \44778 , \24060 , \24173 );
not \U$44402 ( \44779 , \44778 );
not \U$44403 ( \44780 , \24217 );
or \U$44404 ( \44781 , \44779 , \44780 );
not \U$44405 ( \44782 , \24216 );
nand \U$44406 ( \44783 , \44782 , \24184 , \24182 );
nand \U$44407 ( \44784 , \44781 , \44783 );
not \U$44408 ( \44785 , \44784 );
or \U$44409 ( \44786 , \44777 , \44785 );
or \U$44410 ( \44787 , \24245 , \24235 );
nand \U$44411 ( \44788 , \44786 , \44787 );
not \U$44412 ( \44789 , \44788 );
or \U$44413 ( \44790 , \44776 , \44789 );
not \U$44414 ( \44791 , \24259 );
nand \U$44415 ( \44792 , \44791 , \24255 , \24248 );
nand \U$44416 ( \44793 , \44790 , \44792 );
nor \U$44417 ( \44794 , \44775 , \44793 );
nand \U$44418 ( \44795 , \44759 , \44794 );
not \U$44419 ( \44796 , \44795 );
nand \U$44420 ( \44797 , \44635 , \44716 , \44796 );
not \U$44421 ( \44798 , \44797 );
or \U$44422 ( \44799 , \9274 , \44798 );
not \U$44423 ( \44800 , \9271 );
not \U$44424 ( \44801 , \8410 );
not \U$44425 ( \44802 , \8563 );
and \U$44426 ( \44803 , \4528 , \4249 , \4810 , \6823 );
not \U$44427 ( \44804 , \6574 );
not \U$44428 ( \44805 , \6529 );
nor \U$44429 ( \44806 , \6467 , \5843 );
not \U$44430 ( \44807 , \44806 );
or \U$44431 ( \44808 , \44805 , \44807 );
not \U$44432 ( \44809 , \6524 );
not \U$44433 ( \44810 , \6528 );
nand \U$44434 ( \44811 , \44809 , \44810 );
nand \U$44435 ( \44812 , \44808 , \44811 );
nand \U$44436 ( \44813 , \6565 , \44812 );
or \U$44437 ( \44814 , \6557 , \6564 );
nand \U$44438 ( \44815 , \44813 , \44814 );
not \U$44439 ( \44816 , \44815 );
or \U$44440 ( \44817 , \44804 , \44816 );
not \U$44441 ( \44818 , \6573 );
nand \U$44442 ( \44819 , \44818 , \6569 , \6567 );
nand \U$44443 ( \44820 , \44817 , \44819 );
nand \U$44444 ( \44821 , \44803 , \44820 );
not \U$44445 ( \44822 , \4810 );
nand \U$44446 ( \44823 , \4248 , \3872 );
or \U$44447 ( \44824 , \44823 , \4527 );
nand \U$44448 ( \44825 , \4255 , \4526 );
nand \U$44449 ( \44826 , \44824 , \44825 );
not \U$44450 ( \44827 , \44826 );
or \U$44451 ( \44828 , \44822 , \44827 );
or \U$44452 ( \44829 , \4800 , \4809 );
nand \U$44453 ( \44830 , \44828 , \44829 );
nand \U$44454 ( \44831 , \44830 , \6824 );
not \U$44455 ( \44832 , \6822 );
nand \U$44456 ( \44833 , \44832 , \6579 , \6577 );
nand \U$44457 ( \44834 , \44821 , \44831 , \44833 );
not \U$44458 ( \44835 , \44834 );
or \U$44459 ( \44836 , \44802 , \44835 );
not \U$44460 ( \44837 , \8515 );
not \U$44461 ( \44838 , \8561 );
nor \U$44462 ( \44839 , \8540 , \8545 );
not \U$44463 ( \44840 , \44839 );
or \U$44464 ( \44841 , \44838 , \44840 );
not \U$44465 ( \44842 , \8558 );
xor \U$44466 ( \44843 , \8494 , \8511 );
xnor \U$44467 ( \44844 , \44843 , \8508 );
nand \U$44468 ( \44845 , \44842 , \44844 );
nand \U$44469 ( \44846 , \44841 , \44845 );
not \U$44470 ( \44847 , \44846 );
or \U$44471 ( \44848 , \44837 , \44847 );
or \U$44472 ( \44849 , \8492 , \8514 );
nand \U$44473 ( \44850 , \44848 , \44849 );
buf \U$44474 ( \44851 , \8524 );
nand \U$44475 ( \44852 , \44850 , \44851 );
or \U$44476 ( \44853 , \8523 , \8517 );
nand \U$44477 ( \44854 , \44852 , \44853 );
not \U$44478 ( \44855 , \44854 );
nand \U$44479 ( \44856 , \44836 , \44855 );
not \U$44480 ( \44857 , \44856 );
or \U$44481 ( \44858 , \44801 , \44857 );
not \U$44482 ( \44859 , \8230 );
nand \U$44483 ( \44860 , \7970 , \8037 );
or \U$44484 ( \44861 , \7968 , \44860 );
nand \U$44485 ( \44862 , \7967 , \7787 );
nand \U$44486 ( \44863 , \44861 , \44862 );
not \U$44487 ( \44864 , \44863 );
or \U$44488 ( \44865 , \44859 , \44864 );
nand \U$44489 ( \44866 , \8228 , \8229 );
nand \U$44490 ( \44867 , \44866 , \8225 );
nand \U$44491 ( \44868 , \44865 , \44867 );
and \U$44492 ( \44869 , \44868 , \8409 );
or \U$44493 ( \44870 , \8221 , \8231 );
nand \U$44494 ( \44871 , \44870 , \8408 );
not \U$44495 ( \44872 , \44871 );
nor \U$44496 ( \44873 , \44872 , \8406 );
nor \U$44497 ( \44874 , \44869 , \44873 );
nand \U$44498 ( \44875 , \44858 , \44874 );
not \U$44499 ( \44876 , \44875 );
or \U$44500 ( \44877 , \44800 , \44876 );
not \U$44501 ( \44878 , \9270 );
not \U$44502 ( \44879 , \9259 );
not \U$44503 ( \44880 , \9014 );
nand \U$44504 ( \44881 , \8866 , \8859 );
or \U$44505 ( \44882 , \8853 , \44881 );
nand \U$44506 ( \44883 , \8852 , \8717 );
nand \U$44507 ( \44884 , \44882 , \44883 );
not \U$44508 ( \44885 , \44884 );
or \U$44509 ( \44886 , \44880 , \44885 );
or \U$44510 ( \44887 , \8871 , \9013 );
nand \U$44511 ( \44888 , \44886 , \44887 );
nand \U$44512 ( \44889 , \44888 , \9122 );
not \U$44513 ( \44890 , \9121 );
buf \U$44514 ( \44891 , \9021 );
nand \U$44515 ( \44892 , \44890 , \44891 );
nand \U$44516 ( \44893 , \44889 , \44892 );
not \U$44517 ( \44894 , \44893 );
or \U$44518 ( \44895 , \44879 , \44894 );
not \U$44519 ( \44896 , \9258 );
not \U$44520 ( \44897 , \9195 );
nand \U$44521 ( \44898 , \44897 , \9130 );
or \U$44522 ( \44899 , \9233 , \44898 );
nand \U$44523 ( \44900 , \9232 , \9225 );
nand \U$44524 ( \44901 , \44899 , \44900 );
not \U$44525 ( \44902 , \44901 );
or \U$44526 ( \44903 , \44896 , \44902 );
nand \U$44527 ( \44904 , \9241 , \9257 );
nand \U$44528 ( \44905 , \44903 , \44904 );
not \U$44529 ( \44906 , \44905 );
nand \U$44530 ( \44907 , \44895 , \44906 );
not \U$44531 ( \44908 , \44907 );
or \U$44532 ( \44909 , \44878 , \44908 );
nand \U$44533 ( \44910 , \9265 , \9269 );
nand \U$44534 ( \44911 , \44909 , \44910 );
not \U$44535 ( \44912 , \44911 );
nand \U$44536 ( \44913 , \44877 , \44912 );
not \U$44537 ( \44914 , \44913 );
nand \U$44538 ( \44915 , \44799 , \44914 );
not \U$44539 ( \44916 , \44915 );
or \U$44540 ( \44917 , \1720 , \44916 );
nor \U$44541 ( \44918 , \1540 , \1539 );
and \U$44542 ( \44919 , \44918 , \1390 );
nor \U$44543 ( \44920 , \1389 , \1339 );
nor \U$44544 ( \44921 , \44919 , \44920 );
not \U$44545 ( \44922 , \1581 );
or \U$44546 ( \44923 , \44921 , \44922 );
or \U$44547 ( \44924 , \1546 , \1580 );
nand \U$44548 ( \44925 , \44923 , \44924 );
and \U$44549 ( \44926 , \44925 , \1624 );
nor \U$44550 ( \44927 , \1619 , \1623 );
nor \U$44551 ( \44928 , \44926 , \44927 );
not \U$44552 ( \44929 , \1698 );
or \U$44553 ( \44930 , \44928 , \44929 );
or \U$44554 ( \44931 , \1655 , \1659 );
not \U$44555 ( \44932 , \44931 );
not \U$44556 ( \44933 , \1697 );
and \U$44557 ( \44934 , \44932 , \44933 );
not \U$44558 ( \44935 , \1696 );
nor \U$44559 ( \44936 , \44935 , \1665 );
nor \U$44560 ( \44937 , \44934 , \44936 );
nand \U$44561 ( \44938 , \44930 , \44937 );
and \U$44562 ( \44939 , \44938 , \1718 );
nor \U$44563 ( \44940 , \1704 , \1717 );
nor \U$44564 ( \44941 , \44939 , \44940 );
nand \U$44565 ( \44942 , \44917 , \44941 );
not \U$44566 ( \44943 , \44942 );
xor \U$44567 ( \44944 , \1631 , \1706 );
xor \U$44568 ( \44945 , \44944 , \1711 );
and \U$44569 ( \44946 , \1669 , \44945 );
xor \U$44570 ( \44947 , \1631 , \1706 );
xor \U$44571 ( \44948 , \44947 , \1711 );
and \U$44572 ( \44949 , \1715 , \44948 );
and \U$44573 ( \44950 , \1669 , \1715 );
or \U$44574 ( \44951 , \44946 , \44949 , \44950 );
xor \U$44575 ( \44952 , \1631 , \1706 );
and \U$44576 ( \44953 , \44952 , \1711 );
and \U$44577 ( \44954 , \1631 , \1706 );
or \U$44578 ( \44955 , \44953 , \44954 );
not \U$44579 ( \44956 , \44955 );
not \U$44580 ( \44957 , \1673 );
and \U$44581 ( \44958 , \1709 , \1129 );
and \U$44582 ( \44959 , \1122 , RIae78b48_125);
nor \U$44583 ( \44960 , \44958 , \44959 );
not \U$44584 ( \44961 , \44960 );
or \U$44585 ( \44962 , \44957 , \44961 );
or \U$44586 ( \44963 , \44960 , \1673 );
nand \U$44587 ( \44964 , \44962 , \44963 );
not \U$44588 ( \44965 , \44964 );
and \U$44589 ( \44966 , \44956 , \44965 );
and \U$44590 ( \44967 , \44955 , \44964 );
nor \U$44591 ( \44968 , \44966 , \44967 );
xnor \U$44592 ( \44969 , \44951 , \44968 );
not \U$44593 ( \44970 , \44969 );
and \U$44594 ( \44971 , \44943 , \44970 );
and \U$44595 ( \44972 , \44942 , \44969 );
nor \U$44596 ( \44973 , \44971 , \44972 );
not \U$44597 ( \44974 , RIae7aee8_201);
not \U$44598 ( \44975 , RIae7af60_202);
and \U$44599 ( \44976 , \44974 , \44975 );
and \U$44600 ( \44977 , RIae7aee8_201, RIae7af60_202);
nor \U$44601 ( \44978 , \44976 , \44977 );
not \U$44602 ( \44979 , \44978 );
xor \U$44603 ( \44980 , RIae7afd8_203, RIae7b050_204);
not \U$44604 ( \44981 , \44980 );
and \U$44605 ( \44982 , \44979 , \44981 );
and \U$44606 ( \44983 , \44978 , \44980 );
nor \U$44607 ( \44984 , \44982 , \44983 );
not \U$44608 ( \44985 , \44984 );
xor \U$44609 ( \44986 , RIae7b0c8_205, RIae7b140_206);
not \U$44610 ( \44987 , \44986 );
not \U$44611 ( \44988 , RIae7b230_208);
not \U$44612 ( \44989 , RIae7b1b8_207);
or \U$44613 ( \44990 , \44988 , \44989 );
or \U$44614 ( \44991 , RIae7b1b8_207, RIae7b230_208);
nand \U$44615 ( \44992 , \44990 , \44991 );
not \U$44616 ( \44993 , \44992 );
or \U$44617 ( \44994 , \44987 , \44993 );
or \U$44618 ( \44995 , \44992 , \44986 );
nand \U$44619 ( \44996 , \44994 , \44995 );
not \U$44620 ( \44997 , \44996 );
and \U$44621 ( \44998 , \44985 , \44997 );
and \U$44622 ( \44999 , \44984 , \44996 );
nor \U$44623 ( \45000 , \44998 , \44999 );
not \U$44624 ( \45001 , \45000 );
xor \U$44625 ( \45002 , RIae7ab28_193, RIae7aba0_194);
not \U$44626 ( \45003 , \45002 );
not \U$44627 ( \45004 , RIae7ac90_196);
not \U$44628 ( \45005 , RIae7ac18_195);
or \U$44629 ( \45006 , \45004 , \45005 );
or \U$44630 ( \45007 , RIae7ac18_195, RIae7ac90_196);
nand \U$44631 ( \45008 , \45006 , \45007 );
not \U$44632 ( \45009 , \45008 );
or \U$44633 ( \45010 , \45003 , \45009 );
or \U$44634 ( \45011 , \45008 , \45002 );
nand \U$44635 ( \45012 , \45010 , \45011 );
not \U$44636 ( \45013 , \45012 );
xnor \U$44637 ( \45014 , RIae7ad08_197, RIae7ad80_198);
not \U$44638 ( \45015 , \45014 );
xor \U$44639 ( \45016 , RIae7adf8_199, RIae7ae70_200);
not \U$44640 ( \45017 , \45016 );
and \U$44641 ( \45018 , \45015 , \45017 );
and \U$44642 ( \45019 , \45014 , \45016 );
nor \U$44643 ( \45020 , \45018 , \45019 );
not \U$44644 ( \45021 , \45020 );
or \U$44645 ( \45022 , \45013 , \45021 );
or \U$44646 ( \45023 , \45020 , \45012 );
nand \U$44647 ( \45024 , \45022 , \45023 );
not \U$44648 ( \45025 , \45024 );
and \U$44649 ( \45026 , \45001 , \45025 );
and \U$44650 ( \45027 , \45000 , \45024 );
nor \U$44651 ( \45028 , \45026 , \45027 );
not \U$44652 ( \45029 , \45028 );
not \U$44653 ( \45030 , RIae7ba28_225);
not \U$44654 ( \45031 , RIae7baa0_226);
and \U$44655 ( \45032 , \45030 , \45031 );
and \U$44656 ( \45033 , RIae7ba28_225, RIae7baa0_226);
nor \U$44657 ( \45034 , \45032 , \45033 );
not \U$44658 ( \45035 , \45034 );
xor \U$44659 ( \45036 , RIae7bb18_227, RIae7bb90_228);
not \U$44660 ( \45037 , \45036 );
and \U$44661 ( \45038 , \45035 , \45037 );
and \U$44662 ( \45039 , \45034 , \45036 );
nor \U$44663 ( \45040 , \45038 , \45039 );
not \U$44664 ( \45041 , \45040 );
xor \U$44665 ( \45042 , RIae7bed8_235, RIae7bf50_236);
not \U$44666 ( \45043 , \45042 );
xnor \U$44667 ( \45044 , RIae7bde8_233, RIae7be60_234);
not \U$44668 ( \45045 , \45044 );
or \U$44669 ( \45046 , \45043 , \45045 );
or \U$44670 ( \45047 , \45044 , \45042 );
nand \U$44671 ( \45048 , \45046 , \45047 );
not \U$44672 ( \45049 , \45048 );
and \U$44673 ( \45050 , \45041 , \45049 );
and \U$44674 ( \45051 , \45040 , \45048 );
nor \U$44675 ( \45052 , \45050 , \45051 );
not \U$44676 ( \45053 , \45052 );
xor \U$44677 ( \45054 , RIae7b848_221, RIae7b8c0_222);
not \U$44678 ( \45055 , \45054 );
not \U$44679 ( \45056 , RIae7b9b0_224);
not \U$44680 ( \45057 , RIae7b938_223);
or \U$44681 ( \45058 , \45056 , \45057 );
or \U$44682 ( \45059 , RIae7b938_223, RIae7b9b0_224);
nand \U$44683 ( \45060 , \45058 , \45059 );
not \U$44684 ( \45061 , \45060 );
or \U$44685 ( \45062 , \45055 , \45061 );
or \U$44686 ( \45063 , \45060 , \45054 );
nand \U$44687 ( \45064 , \45062 , \45063 );
not \U$44688 ( \45065 , \45064 );
xnor \U$44689 ( \45066 , RIae7b668_217, RIae7b6e0_218);
not \U$44690 ( \45067 , \45066 );
xor \U$44691 ( \45068 , RIae7b758_219, RIae7b7d0_220);
not \U$44692 ( \45069 , \45068 );
and \U$44693 ( \45070 , \45067 , \45069 );
and \U$44694 ( \45071 , \45066 , \45068 );
nor \U$44695 ( \45072 , \45070 , \45071 );
not \U$44696 ( \45073 , \45072 );
or \U$44697 ( \45074 , \45065 , \45073 );
or \U$44698 ( \45075 , \45072 , \45064 );
nand \U$44699 ( \45076 , \45074 , \45075 );
not \U$44700 ( \45077 , \45076 );
or \U$44701 ( \45078 , \45053 , \45077 );
or \U$44702 ( \45079 , \45052 , \45076 );
nand \U$44703 ( \45080 , \45078 , \45079 );
not \U$44704 ( \45081 , \45080 );
and \U$44705 ( \45082 , \45029 , \45081 );
and \U$44706 ( \45083 , \45028 , \45080 );
nor \U$44707 ( \45084 , \45082 , \45083 );
not \U$44708 ( \45085 , \45084 );
not \U$44709 ( \45086 , RIae7bfc8_237);
not \U$44710 ( \45087 , RIae7c040_238);
and \U$44711 ( \45088 , \45086 , \45087 );
and \U$44712 ( \45089 , RIae7bfc8_237, RIae7c040_238);
nor \U$44713 ( \45090 , \45088 , \45089 );
not \U$44714 ( \45091 , \45090 );
xor \U$44715 ( \45092 , RIae7c0b8_239, RIae7c130_240);
not \U$44716 ( \45093 , \45092 );
and \U$44717 ( \45094 , \45091 , \45093 );
and \U$44718 ( \45095 , \45090 , \45092 );
nor \U$44719 ( \45096 , \45094 , \45095 );
not \U$44720 ( \45097 , \45096 );
not \U$44721 ( \45098 , RIae7c658_251);
not \U$44722 ( \45099 , RIae7c6d0_252);
and \U$44723 ( \45100 , \45098 , \45099 );
and \U$44724 ( \45101 , RIae7c658_251, RIae7c6d0_252);
nor \U$44725 ( \45102 , \45100 , \45101 );
not \U$44726 ( \45103 , \45102 );
xor \U$44727 ( \45104 , RIae7bc08_229, RIae7bc80_230);
not \U$44728 ( \45105 , \45104 );
and \U$44729 ( \45106 , \45103 , \45105 );
and \U$44730 ( \45107 , \45102 , \45104 );
nor \U$44731 ( \45108 , \45106 , \45107 );
not \U$44732 ( \45109 , \45108 );
and \U$44733 ( \45110 , \45097 , \45109 );
and \U$44734 ( \45111 , \45108 , \45096 );
nor \U$44735 ( \45112 , \45110 , \45111 );
not \U$44736 ( \45113 , \45112 );
xor \U$44737 ( \45114 , RIae7c748_253, RIae7c7c0_254);
not \U$44738 ( \45115 , \45114 );
not \U$44739 ( \45116 , RIae7c8b0_256);
not \U$44740 ( \45117 , RIae7c838_255);
or \U$44741 ( \45118 , \45116 , \45117 );
or \U$44742 ( \45119 , RIae7c838_255, RIae7c8b0_256);
nand \U$44743 ( \45120 , \45118 , \45119 );
not \U$44744 ( \45121 , \45120 );
or \U$44745 ( \45122 , \45115 , \45121 );
or \U$44746 ( \45123 , \45120 , \45114 );
nand \U$44747 ( \45124 , \45122 , \45123 );
not \U$44748 ( \45125 , \45124 );
xnor \U$44749 ( \45126 , RIae7bcf8_231, RIae7bd70_232);
not \U$44750 ( \45127 , \45126 );
xor \U$44751 ( \45128 , RIae7c568_249, RIae7c5e0_250);
not \U$44752 ( \45129 , \45128 );
and \U$44753 ( \45130 , \45127 , \45129 );
and \U$44754 ( \45131 , \45126 , \45128 );
nor \U$44755 ( \45132 , \45130 , \45131 );
not \U$44756 ( \45133 , \45132 );
or \U$44757 ( \45134 , \45125 , \45133 );
or \U$44758 ( \45135 , \45132 , \45124 );
nand \U$44759 ( \45136 , \45134 , \45135 );
not \U$44760 ( \45137 , \45136 );
and \U$44761 ( \45138 , \45113 , \45137 );
and \U$44762 ( \45139 , \45112 , \45136 );
nor \U$44763 ( \45140 , \45138 , \45139 );
not \U$44764 ( \45141 , \45140 );
xnor \U$44765 ( \45142 , RIae7c388_245, RIae7c400_246);
not \U$44766 ( \45143 , \45142 );
xor \U$44767 ( \45144 , RIae7c478_247, RIae7c4f0_248);
not \U$44768 ( \45145 , \45144 );
and \U$44769 ( \45146 , \45143 , \45145 );
and \U$44770 ( \45147 , \45142 , \45144 );
nor \U$44771 ( \45148 , \45146 , \45147 );
not \U$44772 ( \45149 , \45148 );
not \U$44773 ( \45150 , RIae7c1a8_241);
not \U$44774 ( \45151 , RIae7c220_242);
and \U$44775 ( \45152 , \45150 , \45151 );
and \U$44776 ( \45153 , RIae7c1a8_241, RIae7c220_242);
nor \U$44777 ( \45154 , \45152 , \45153 );
not \U$44778 ( \45155 , \45154 );
xor \U$44779 ( \45156 , RIae7c298_243, RIae7c310_244);
not \U$44780 ( \45157 , \45156 );
and \U$44781 ( \45158 , \45155 , \45157 );
and \U$44782 ( \45159 , \45154 , \45156 );
nor \U$44783 ( \45160 , \45158 , \45159 );
not \U$44784 ( \45161 , \45160 );
and \U$44785 ( \45162 , \45149 , \45161 );
and \U$44786 ( \45163 , \45148 , \45160 );
nor \U$44787 ( \45164 , \45162 , \45163 );
not \U$44788 ( \45165 , \45164 );
xor \U$44789 ( \45166 , RIae7b488_213, RIae7b500_214);
not \U$44790 ( \45167 , \45166 );
not \U$44791 ( \45168 , RIae7b5f0_216);
not \U$44792 ( \45169 , RIae7b578_215);
or \U$44793 ( \45170 , \45168 , \45169 );
or \U$44794 ( \45171 , RIae7b578_215, RIae7b5f0_216);
nand \U$44795 ( \45172 , \45170 , \45171 );
not \U$44796 ( \45173 , \45172 );
or \U$44797 ( \45174 , \45167 , \45173 );
or \U$44798 ( \45175 , \45172 , \45166 );
nand \U$44799 ( \45176 , \45174 , \45175 );
not \U$44800 ( \45177 , \45176 );
xor \U$44801 ( \45178 , RIae7b398_211, RIae7b410_212);
not \U$44802 ( \45179 , \45178 );
xor \U$44803 ( \45180 , RIae7b2a8_209, RIae7b320_210);
not \U$44804 ( \45181 , \45180 );
or \U$44805 ( \45182 , \45179 , \45181 );
or \U$44806 ( \45183 , \45180 , \45178 );
nand \U$44807 ( \45184 , \45182 , \45183 );
not \U$44808 ( \45185 , \45184 );
or \U$44809 ( \45186 , \45177 , \45185 );
or \U$44810 ( \45187 , \45184 , \45176 );
nand \U$44811 ( \45188 , \45186 , \45187 );
not \U$44812 ( \45189 , \45188 );
or \U$44813 ( \45190 , \45165 , \45189 );
or \U$44814 ( \45191 , \45164 , \45188 );
nand \U$44815 ( \45192 , \45190 , \45191 );
not \U$44816 ( \45193 , \45192 );
or \U$44817 ( \45194 , \45141 , \45193 );
or \U$44818 ( \45195 , \45140 , \45192 );
nand \U$44819 ( \45196 , \45194 , \45195 );
not \U$44820 ( \45197 , \45196 );
and \U$44821 ( \45198 , \45085 , \45197 );
and \U$44822 ( \45199 , \45084 , \45196 );
nor \U$44823 ( \45200 , \45198 , \45199 );
buf \U$44824 ( \45201 , \45200 );
not \U$44825 ( \45202 , \45201 );
not \U$44826 ( \45203 , \45202 );
not \U$44827 ( \45204 , \45203 );
nor \U$44828 ( \45205 , \44973 , \45204 );
buf \U$44829 ( \45206 , \45205 );
not \U$44830 ( \45207 , \9271 );
nand \U$44831 ( \45208 , \1625 , \1698 );
nor \U$44832 ( \45209 , \45207 , \45208 );
not \U$44833 ( \45210 , \45209 );
not \U$44834 ( \45211 , \6825 );
nor \U$44835 ( \45212 , \45211 , \8564 );
not \U$44836 ( \45213 , \45212 );
nand \U$44837 ( \45214 , \44635 , \44716 , \44796 );
not \U$44838 ( \45215 , \45214 );
or \U$44839 ( \45216 , \45213 , \45215 );
not \U$44840 ( \45217 , \44875 );
nand \U$44841 ( \45218 , \45216 , \45217 );
not \U$44842 ( \45219 , \45218 );
or \U$44843 ( \45220 , \45210 , \45219 );
not \U$44844 ( \45221 , \1698 );
not \U$44845 ( \45222 , \1625 );
not \U$44846 ( \45223 , \44911 );
or \U$44847 ( \45224 , \45222 , \45223 );
buf \U$44848 ( \45225 , \44928 );
nand \U$44849 ( \45226 , \45224 , \45225 );
not \U$44850 ( \45227 , \45226 );
or \U$44851 ( \45228 , \45221 , \45227 );
nand \U$44852 ( \45229 , \45228 , \44937 );
not \U$44853 ( \45230 , \45229 );
nand \U$44854 ( \45231 , \45220 , \45230 );
not \U$44855 ( \45232 , \45231 );
not \U$44856 ( \45233 , \44940 );
nand \U$44857 ( \45234 , \45233 , \1718 );
not \U$44858 ( \45235 , \45234 );
and \U$44859 ( \45236 , \45232 , \45235 );
and \U$44860 ( \45237 , \45231 , \45234 );
nor \U$44861 ( \45238 , \45236 , \45237 );
nor \U$44862 ( \45239 , \45238 , \45204 );
buf \U$44863 ( \45240 , \45239 );
nand \U$44864 ( \45241 , \1625 , \1660 );
nor \U$44865 ( \45242 , \45207 , \45241 );
not \U$44866 ( \45243 , \45242 );
not \U$44867 ( \45244 , \45218 );
or \U$44868 ( \45245 , \45243 , \45244 );
not \U$44869 ( \45246 , \1660 );
not \U$44870 ( \45247 , \45226 );
or \U$44871 ( \45248 , \45246 , \45247 );
nand \U$44872 ( \45249 , \45248 , \44931 );
not \U$44873 ( \45250 , \45249 );
nand \U$44874 ( \45251 , \45245 , \45250 );
or \U$44875 ( \45252 , \44936 , \1697 );
xor \U$44876 ( \45253 , \45251 , \45252 );
nor \U$44877 ( \45254 , \45253 , \45204 );
buf \U$44878 ( \45255 , \45254 );
not \U$44879 ( \45256 , \1625 );
not \U$44880 ( \45257 , \44915 );
or \U$44881 ( \45258 , \45256 , \45257 );
nand \U$44882 ( \45259 , \45258 , \45225 );
not \U$44883 ( \45260 , \45259 );
nand \U$44884 ( \45261 , \44931 , \1660 );
not \U$44885 ( \45262 , \45261 );
and \U$44886 ( \45263 , \45260 , \45262 );
and \U$44887 ( \45264 , \45259 , \45261 );
nor \U$44888 ( \45265 , \45263 , \45264 );
nor \U$44889 ( \45266 , \45265 , \45204 );
buf \U$44890 ( \45267 , \45266 );
not \U$44891 ( \45268 , \1582 );
not \U$44892 ( \45269 , \45214 );
or \U$44893 ( \45270 , \45269 , \9272 );
nand \U$44894 ( \45271 , \45270 , \44914 );
not \U$44895 ( \45272 , \45271 );
or \U$44896 ( \45273 , \45268 , \45272 );
not \U$44897 ( \45274 , \44925 );
nand \U$44898 ( \45275 , \45273 , \45274 );
not \U$44899 ( \45276 , \45275 );
not \U$44900 ( \45277 , \44927 );
nand \U$44901 ( \45278 , \45277 , \1624 );
not \U$44902 ( \45279 , \45278 );
and \U$44903 ( \45280 , \45276 , \45279 );
and \U$44904 ( \45281 , \45275 , \45278 );
nor \U$44905 ( \45282 , \45280 , \45281 );
nor \U$44906 ( \45283 , \45282 , \45204 );
buf \U$44907 ( \45284 , \45283 );
not \U$44908 ( \45285 , \1542 );
not \U$44909 ( \45286 , \44915 );
or \U$44910 ( \45287 , \45285 , \45286 );
nand \U$44911 ( \45288 , \45287 , \44921 );
not \U$44912 ( \45289 , \45288 );
nand \U$44913 ( \45290 , \1581 , \44924 );
not \U$44914 ( \45291 , \45290 );
and \U$44915 ( \45292 , \45289 , \45291 );
and \U$44916 ( \45293 , \45288 , \45290 );
nor \U$44917 ( \45294 , \45292 , \45293 );
nor \U$44918 ( \45295 , \45294 , \45204 );
buf \U$44919 ( \45296 , \45295 );
not \U$44920 ( \45297 , \1541 );
not \U$44921 ( \45298 , \44915 );
or \U$44922 ( \45299 , \45297 , \45298 );
not \U$44923 ( \45300 , \44918 );
nand \U$44924 ( \45301 , \45299 , \45300 );
not \U$44925 ( \45302 , \45301 );
not \U$44926 ( \45303 , \44920 );
nand \U$44927 ( \45304 , \45303 , \1390 );
not \U$44928 ( \45305 , \45304 );
and \U$44929 ( \45306 , \45302 , \45305 );
and \U$44930 ( \45307 , \45301 , \45304 );
nor \U$44931 ( \45308 , \45306 , \45307 );
nor \U$44932 ( \45309 , \45308 , \45204 );
buf \U$44933 ( \45310 , \45309 );
nand \U$44934 ( \45311 , \45300 , \1541 );
xor \U$44935 ( \45312 , \44915 , \45311 );
nor \U$44936 ( \45313 , \45312 , \45204 );
buf \U$44937 ( \45314 , \45313 );
buf \U$44938 ( \45315 , \9124 );
and \U$44939 ( \45316 , \45315 , \9259 );
not \U$44940 ( \45317 , \45316 );
not \U$44941 ( \45318 , \45218 );
or \U$44942 ( \45319 , \45317 , \45318 );
not \U$44943 ( \45320 , \44907 );
nand \U$44944 ( \45321 , \45319 , \45320 );
nand \U$44945 ( \45322 , \9270 , \44910 );
xor \U$44946 ( \45323 , \45321 , \45322 );
nor \U$44947 ( \45324 , \45323 , \45204 );
buf \U$44948 ( \45325 , \45324 );
and \U$44949 ( \45326 , \9234 , \9196 );
not \U$44950 ( \45327 , \45326 );
and \U$44951 ( \45328 , \6825 , \8565 , \45315 );
not \U$44952 ( \45329 , \45328 );
not \U$44953 ( \45330 , \44795 );
nand \U$44954 ( \45331 , \44635 , \44716 , \45330 );
not \U$44955 ( \45332 , \45331 );
or \U$44956 ( \45333 , \45329 , \45332 );
not \U$44957 ( \45334 , \45217 );
and \U$44958 ( \45335 , \45334 , \45315 );
not \U$44959 ( \45336 , \9122 );
not \U$44960 ( \45337 , \44888 );
or \U$44961 ( \45338 , \45336 , \45337 );
nand \U$44962 ( \45339 , \45338 , \44892 );
nor \U$44963 ( \45340 , \45335 , \45339 );
nand \U$44964 ( \45341 , \45333 , \45340 );
not \U$44965 ( \45342 , \45341 );
or \U$44966 ( \45343 , \45327 , \45342 );
not \U$44967 ( \45344 , \44901 );
nand \U$44968 ( \45345 , \45343 , \45344 );
not \U$44969 ( \45346 , \45345 );
nand \U$44970 ( \45347 , \9258 , \44904 );
not \U$44971 ( \45348 , \45347 );
and \U$44972 ( \45349 , \45346 , \45348 );
and \U$44973 ( \45350 , \45345 , \45347 );
nor \U$44974 ( \45351 , \45349 , \45350 );
nor \U$44975 ( \45352 , \45351 , \45204 );
buf \U$44976 ( \45353 , \45352 );
not \U$44977 ( \45354 , \9196 );
not \U$44978 ( \45355 , \45341 );
or \U$44979 ( \45356 , \45354 , \45355 );
not \U$44980 ( \45357 , \9195 );
nand \U$44981 ( \45358 , \45357 , \9130 );
nand \U$44982 ( \45359 , \45356 , \45358 );
not \U$44983 ( \45360 , \45359 );
nand \U$44984 ( \45361 , \9234 , \44900 );
not \U$44985 ( \45362 , \45361 );
and \U$44986 ( \45363 , \45360 , \45362 );
and \U$44987 ( \45364 , \45359 , \45361 );
nor \U$44988 ( \45365 , \45363 , \45364 );
nor \U$44989 ( \45366 , \45365 , \45204 );
buf \U$44990 ( \45367 , \45366 );
buf \U$44991 ( \45368 , \45341 );
not \U$44992 ( \45369 , \45368 );
nand \U$44993 ( \45370 , \9196 , \44898 );
not \U$44994 ( \45371 , \45370 );
and \U$44995 ( \45372 , \45369 , \45371 );
and \U$44996 ( \45373 , \45368 , \45370 );
nor \U$44997 ( \45374 , \45372 , \45373 );
nor \U$44998 ( \45375 , \45374 , \45204 );
buf \U$44999 ( \45376 , \45375 );
not \U$45000 ( \45377 , \45203 );
not \U$45001 ( \45378 , \8868 );
not \U$45002 ( \45379 , \45378 );
not \U$45003 ( \45380 , \45218 );
or \U$45004 ( \45381 , \45379 , \45380 );
buf \U$45005 ( \45382 , \44884 );
not \U$45006 ( \45383 , \45382 );
nand \U$45007 ( \45384 , \45381 , \45383 );
nand \U$45008 ( \45385 , \9122 , \44892 );
and \U$45009 ( \45386 , \45385 , \9014 );
and \U$45010 ( \45387 , \45384 , \45386 );
not \U$45011 ( \45388 , \44887 );
nor \U$45012 ( \45389 , \45382 , \45385 , \45388 );
not \U$45013 ( \45390 , \45389 );
nand \U$45014 ( \45391 , \45218 , \45378 );
not \U$45015 ( \45392 , \45391 );
or \U$45016 ( \45393 , \45390 , \45392 );
not \U$45017 ( \45394 , \45385 );
not \U$45018 ( \45395 , \9014 );
and \U$45019 ( \45396 , \45394 , \45395 );
and \U$45020 ( \45397 , \45385 , \45388 );
nor \U$45021 ( \45398 , \45396 , \45397 );
nand \U$45022 ( \45399 , \45393 , \45398 );
nor \U$45023 ( \45400 , \45387 , \45399 );
nor \U$45024 ( \45401 , \45377 , \45400 );
buf \U$45025 ( \45402 , \45401 );
nand \U$45026 ( \45403 , \9014 , \44887 );
xor \U$45027 ( \45404 , \45384 , \45403 );
nor \U$45028 ( \45405 , \45404 , \45204 );
buf \U$45029 ( \45406 , \45405 );
not \U$45030 ( \45407 , \8867 );
not \U$45031 ( \45408 , \45218 );
or \U$45032 ( \45409 , \45407 , \45408 );
nand \U$45033 ( \45410 , \45409 , \44881 );
nand \U$45034 ( \45411 , \8854 , \44883 );
xor \U$45035 ( \45412 , \45410 , \45411 );
nor \U$45036 ( \45413 , \45412 , \45204 );
buf \U$45037 ( \45414 , \45413 );
or \U$45038 ( \45415 , \8859 , \8866 );
nand \U$45039 ( \45416 , \45415 , \44881 );
xor \U$45040 ( \45417 , \45416 , \45218 );
nor \U$45041 ( \45418 , \45417 , \45204 );
buf \U$45042 ( \45419 , \45418 );
and \U$45043 ( \45420 , \8038 , \7969 , \8230 );
nor \U$45044 ( \45421 , \45420 , \44868 );
not \U$45045 ( \45422 , \8409 );
nor \U$45046 ( \45423 , \45422 , \44873 );
nor \U$45047 ( \45424 , \45421 , \45423 , \45202 );
not \U$45048 ( \45425 , \45424 );
not \U$45049 ( \45426 , \6825 );
not \U$45050 ( \45427 , \44797 );
or \U$45051 ( \45428 , \45426 , \45427 );
not \U$45052 ( \45429 , \44834 );
nand \U$45053 ( \45430 , \45428 , \45429 );
nand \U$45054 ( \45431 , \8563 , \45430 );
or \U$45055 ( \45432 , \45425 , \45431 );
not \U$45056 ( \45433 , \44868 );
not \U$45057 ( \45434 , \45433 );
nand \U$45058 ( \45435 , \45423 , \45203 );
nor \U$45059 ( \45436 , \45434 , \45435 , \44854 );
nand \U$45060 ( \45437 , \45431 , \45436 );
not \U$45061 ( \45438 , \45421 );
not \U$45062 ( \45439 , \45438 );
not \U$45063 ( \45440 , \45435 );
and \U$45064 ( \45441 , \45439 , \45440 );
nand \U$45065 ( \45442 , \44852 , \45433 , \44853 );
and \U$45066 ( \45443 , \45442 , \45424 );
nor \U$45067 ( \45444 , \45441 , \45443 );
nand \U$45068 ( \45445 , \45432 , \45437 , \45444 );
buf \U$45069 ( \45446 , \45445 );
not \U$45070 ( \45447 , \8038 );
nor \U$45071 ( \45448 , \45447 , \7968 );
not \U$45072 ( \45449 , \45448 );
not \U$45073 ( \45450 , \44856 );
not \U$45074 ( \45451 , \44716 );
not \U$45075 ( \45452 , \44635 );
or \U$45076 ( \45453 , \45451 , \45452 );
and \U$45077 ( \45454 , \6825 , \8563 );
nand \U$45078 ( \45455 , \45453 , \45454 );
not \U$45079 ( \45456 , \45330 );
nand \U$45080 ( \45457 , \45456 , \45454 );
nand \U$45081 ( \45458 , \45450 , \45455 , \45457 );
not \U$45082 ( \45459 , \45458 );
or \U$45083 ( \45460 , \45449 , \45459 );
not \U$45084 ( \45461 , \44863 );
nand \U$45085 ( \45462 , \45460 , \45461 );
nand \U$45086 ( \45463 , \8230 , \44867 );
xor \U$45087 ( \45464 , \45462 , \45463 );
nor \U$45088 ( \45465 , \45464 , \45204 );
buf \U$45089 ( \45466 , \45465 );
not \U$45090 ( \45467 , \8038 );
not \U$45091 ( \45468 , \45458 );
or \U$45092 ( \45469 , \45467 , \45468 );
nand \U$45093 ( \45470 , \45469 , \44860 );
nand \U$45094 ( \45471 , \7969 , \44862 );
xor \U$45095 ( \45472 , \45470 , \45471 );
nor \U$45096 ( \45473 , \45472 , \45204 );
buf \U$45097 ( \45474 , \45473 );
not \U$45098 ( \45475 , \45458 );
nand \U$45099 ( \45476 , \8038 , \44860 );
not \U$45100 ( \45477 , \45476 );
and \U$45101 ( \45478 , \45475 , \45477 );
and \U$45102 ( \45479 , \45458 , \45476 );
nor \U$45103 ( \45480 , \45478 , \45479 );
nor \U$45104 ( \45481 , \45480 , \45204 );
buf \U$45105 ( \45482 , \45481 );
and \U$45106 ( \45483 , \44853 , \44851 );
not \U$45107 ( \45484 , \8515 );
nor \U$45108 ( \45485 , \45483 , \45484 );
and \U$45109 ( \45486 , \8546 , \8562 );
not \U$45110 ( \45487 , \45486 );
not \U$45111 ( \45488 , \45430 );
or \U$45112 ( \45489 , \45487 , \45488 );
not \U$45113 ( \45490 , \44846 );
nand \U$45114 ( \45491 , \45489 , \45490 );
and \U$45115 ( \45492 , \45485 , \45491 );
and \U$45116 ( \45493 , \45490 , \45483 , \44849 );
not \U$45117 ( \45494 , \45493 );
nand \U$45118 ( \45495 , \45430 , \45486 );
not \U$45119 ( \45496 , \45495 );
or \U$45120 ( \45497 , \45494 , \45496 );
not \U$45121 ( \45498 , \45483 );
not \U$45122 ( \45499 , \44849 );
and \U$45123 ( \45500 , \45498 , \45499 );
and \U$45124 ( \45501 , \45483 , \45484 );
nor \U$45125 ( \45502 , \45500 , \45501 );
nand \U$45126 ( \45503 , \45497 , \45502 );
nor \U$45127 ( \45504 , \45492 , \45503 );
nor \U$45128 ( \45505 , \45204 , \45504 );
buf \U$45129 ( \45506 , \45505 );
nand \U$45130 ( \45507 , \8515 , \44849 );
xor \U$45131 ( \45508 , \45491 , \45507 );
nor \U$45132 ( \45509 , \45508 , \45204 );
buf \U$45133 ( \45510 , \45509 );
not \U$45134 ( \45511 , \8546 );
not \U$45135 ( \45512 , \45430 );
or \U$45136 ( \45513 , \45511 , \45512 );
not \U$45137 ( \45514 , \44839 );
nand \U$45138 ( \45515 , \45513 , \45514 );
nand \U$45139 ( \45516 , \44845 , \8562 );
xor \U$45140 ( \45517 , \45515 , \45516 );
nor \U$45141 ( \45518 , \45517 , \45204 );
buf \U$45142 ( \45519 , \45518 );
nand \U$45143 ( \45520 , \45514 , \8546 );
xor \U$45144 ( \45521 , \45430 , \45520 );
nor \U$45145 ( \45522 , \45521 , \45204 );
buf \U$45146 ( \45523 , \45522 );
not \U$45147 ( \45524 , \6575 );
not \U$45148 ( \45525 , \44797 );
or \U$45149 ( \45526 , \45524 , \45525 );
not \U$45150 ( \45527 , \44820 );
nand \U$45151 ( \45528 , \45526 , \45527 );
not \U$45152 ( \45529 , \45528 );
not \U$45153 ( \45530 , \4811 );
or \U$45154 ( \45531 , \45529 , \45530 );
not \U$45155 ( \45532 , \44830 );
nand \U$45156 ( \45533 , \45531 , \45532 );
nand \U$45157 ( \45534 , \6824 , \44833 );
xor \U$45158 ( \45535 , \45533 , \45534 );
nor \U$45159 ( \45536 , \45535 , \45204 );
buf \U$45160 ( \45537 , \45536 );
buf \U$45161 ( \45538 , \4250 );
and \U$45162 ( \45539 , \4528 , \45538 );
not \U$45163 ( \45540 , \45539 );
not \U$45164 ( \45541 , \45528 );
or \U$45165 ( \45542 , \45540 , \45541 );
not \U$45166 ( \45543 , \44826 );
nand \U$45167 ( \45544 , \45542 , \45543 );
nand \U$45168 ( \45545 , \4810 , \44829 );
xor \U$45169 ( \45546 , \45544 , \45545 );
nor \U$45170 ( \45547 , \45546 , \45204 );
buf \U$45171 ( \45548 , \45547 );
not \U$45172 ( \45549 , \45538 );
not \U$45173 ( \45550 , \45528 );
or \U$45174 ( \45551 , \45549 , \45550 );
nand \U$45175 ( \45552 , \45551 , \44823 );
nand \U$45176 ( \45553 , \4528 , \44825 );
xor \U$45177 ( \45554 , \45552 , \45553 );
nor \U$45178 ( \45555 , \45554 , \45204 );
buf \U$45179 ( \45556 , \45555 );
nand \U$45180 ( \45557 , \44823 , \45538 );
xor \U$45181 ( \45558 , \45528 , \45557 );
nor \U$45182 ( \45559 , \45558 , \45204 );
buf \U$45183 ( \45560 , \45559 );
and \U$45184 ( \45561 , \6530 , \6565 );
not \U$45185 ( \45562 , \45561 );
not \U$45186 ( \45563 , \44797 );
or \U$45187 ( \45564 , \45562 , \45563 );
not \U$45188 ( \45565 , \44815 );
nand \U$45189 ( \45566 , \45564 , \45565 );
not \U$45190 ( \45567 , \45566 );
nand \U$45191 ( \45568 , \44819 , \6574 );
not \U$45192 ( \45569 , \45568 );
and \U$45193 ( \45570 , \45567 , \45569 );
and \U$45194 ( \45571 , \45566 , \45568 );
nor \U$45195 ( \45572 , \45570 , \45571 );
nor \U$45196 ( \45573 , \45572 , \45202 );
buf \U$45197 ( \45574 , \45573 );
not \U$45198 ( \45575 , \6530 );
not \U$45199 ( \45576 , \45331 );
or \U$45200 ( \45577 , \45575 , \45576 );
not \U$45201 ( \45578 , \44812 );
nand \U$45202 ( \45579 , \45577 , \45578 );
nand \U$45203 ( \45580 , \44814 , \6565 );
xor \U$45204 ( \45581 , \45579 , \45580 );
nor \U$45205 ( \45582 , \45581 , \45202 );
buf \U$45206 ( \45583 , \45582 );
not \U$45207 ( \45584 , \6468 );
not \U$45208 ( \45585 , \45331 );
or \U$45209 ( \45586 , \45584 , \45585 );
not \U$45210 ( \45587 , \44806 );
nand \U$45211 ( \45588 , \45586 , \45587 );
nand \U$45212 ( \45589 , \6529 , \44811 );
xor \U$45213 ( \45590 , \45588 , \45589 );
nor \U$45214 ( \45591 , \45590 , \45202 );
buf \U$45215 ( \45592 , \45591 );
nand \U$45216 ( \45593 , \45587 , \6468 );
xor \U$45217 ( \45594 , \45331 , \45593 );
nor \U$45218 ( \45595 , \45594 , \45202 );
buf \U$45219 ( \45596 , \45595 );
and \U$45220 ( \45597 , \44717 , \24246 );
not \U$45221 ( \45598 , \45597 );
not \U$45222 ( \45599 , \27524 );
not \U$45223 ( \45600 , \27288 );
not \U$45224 ( \45601 , \44715 );
not \U$45225 ( \45602 , \44632 );
nand \U$45226 ( \45603 , \45602 , \35663 , \44618 );
buf \U$45227 ( \45604 , \15931 );
buf \U$45228 ( \45605 , \20772 );
buf \U$45229 ( \45606 , \22816 );
nand \U$45230 ( \45607 , \45603 , \45604 , \45605 , \45606 );
nand \U$45231 ( \45608 , \45601 , \45607 );
not \U$45232 ( \45609 , \45608 );
or \U$45233 ( \45610 , \45600 , \45609 );
not \U$45234 ( \45611 , \44757 );
nand \U$45235 ( \45612 , \45610 , \45611 );
not \U$45236 ( \45613 , \45612 );
or \U$45237 ( \45614 , \45599 , \45613 );
not \U$45238 ( \45615 , \44774 );
nand \U$45239 ( \45616 , \45614 , \45615 );
not \U$45240 ( \45617 , \45616 );
or \U$45241 ( \45618 , \45598 , \45617 );
not \U$45242 ( \45619 , \44788 );
nand \U$45243 ( \45620 , \45618 , \45619 );
not \U$45244 ( \45621 , \45620 );
nand \U$45245 ( \45622 , \44792 , \24260 );
not \U$45246 ( \45623 , \45622 );
and \U$45247 ( \45624 , \45621 , \45623 );
and \U$45248 ( \45625 , \45620 , \45622 );
nor \U$45249 ( \45626 , \45624 , \45625 );
nor \U$45250 ( \45627 , \45626 , \45204 );
buf \U$45251 ( \45628 , \45627 );
not \U$45252 ( \45629 , \44717 );
not \U$45253 ( \45630 , \45616 );
or \U$45254 ( \45631 , \45629 , \45630 );
not \U$45255 ( \45632 , \44784 );
nand \U$45256 ( \45633 , \45631 , \45632 );
not \U$45257 ( \45634 , \45633 );
nand \U$45258 ( \45635 , \44787 , \24246 );
not \U$45259 ( \45636 , \45635 );
and \U$45260 ( \45637 , \45634 , \45636 );
and \U$45261 ( \45638 , \45633 , \45635 );
nor \U$45262 ( \45639 , \45637 , \45638 );
nor \U$45263 ( \45640 , \45639 , \45204 );
buf \U$45264 ( \45641 , \45640 );
buf \U$45265 ( \45642 , \24175 );
not \U$45266 ( \45643 , \45642 );
not \U$45267 ( \45644 , \45616 );
or \U$45268 ( \45645 , \45643 , \45644 );
not \U$45269 ( \45646 , \44778 );
nand \U$45270 ( \45647 , \45645 , \45646 );
not \U$45271 ( \45648 , \45647 );
nand \U$45272 ( \45649 , \24218 , \44783 );
not \U$45273 ( \45650 , \45649 );
and \U$45274 ( \45651 , \45648 , \45650 );
and \U$45275 ( \45652 , \45647 , \45649 );
nor \U$45276 ( \45653 , \45651 , \45652 );
nor \U$45277 ( \45654 , \45653 , \45204 );
buf \U$45278 ( \45655 , \45654 );
nand \U$45279 ( \45656 , \45646 , \45642 );
xor \U$45280 ( \45657 , \45616 , \45656 );
nor \U$45281 ( \45658 , \45657 , \45204 );
buf \U$45282 ( \45659 , \45658 );
buf \U$45283 ( \45660 , \27522 );
not \U$45284 ( \45661 , \45660 );
not \U$45285 ( \45662 , \27468 );
not \U$45286 ( \45663 , \45662 );
not \U$45287 ( \45664 , \45612 );
or \U$45288 ( \45665 , \45663 , \45664 );
not \U$45289 ( \45666 , \44765 );
nand \U$45290 ( \45667 , \45665 , \45666 );
not \U$45291 ( \45668 , \45667 );
or \U$45292 ( \45669 , \45661 , \45668 );
not \U$45293 ( \45670 , \44766 );
nand \U$45294 ( \45671 , \45669 , \45670 );
not \U$45295 ( \45672 , \45671 );
not \U$45296 ( \45673 , \27502 );
not \U$45297 ( \45674 , \27506 );
or \U$45298 ( \45675 , \45673 , \45674 );
or \U$45299 ( \45676 , \27506 , \27502 );
nand \U$45300 ( \45677 , \45675 , \45676 );
not \U$45301 ( \45678 , \45677 );
and \U$45302 ( \45679 , \45672 , \45678 );
and \U$45303 ( \45680 , \45671 , \45677 );
nor \U$45304 ( \45681 , \45679 , \45680 );
nor \U$45305 ( \45682 , \45681 , \45204 );
buf \U$45306 ( \45683 , \45682 );
not \U$45307 ( \45684 , \45667 );
nand \U$45308 ( \45685 , \45670 , \45660 );
not \U$45309 ( \45686 , \45685 );
and \U$45310 ( \45687 , \45684 , \45686 );
and \U$45311 ( \45688 , \45667 , \45685 );
nor \U$45312 ( \45689 , \45687 , \45688 );
nor \U$45313 ( \45690 , \45689 , \45204 );
buf \U$45314 ( \45691 , \45690 );
not \U$45315 ( \45692 , \27467 );
buf \U$45316 ( \45693 , \45612 );
not \U$45317 ( \45694 , \45693 );
or \U$45318 ( \45695 , \45692 , \45694 );
not \U$45319 ( \45696 , \44761 );
nand \U$45320 ( \45697 , \45695 , \45696 );
not \U$45321 ( \45698 , \45697 );
nand \U$45322 ( \45699 , \44764 , \27459 );
not \U$45323 ( \45700 , \45699 );
and \U$45324 ( \45701 , \45698 , \45700 );
and \U$45325 ( \45702 , \45697 , \45699 );
nor \U$45326 ( \45703 , \45701 , \45702 );
nor \U$45327 ( \45704 , \45703 , \45204 );
buf \U$45328 ( \45705 , \45704 );
not \U$45329 ( \45706 , \44761 );
nand \U$45330 ( \45707 , \45706 , \27467 );
xor \U$45331 ( \45708 , \45693 , \45707 );
nor \U$45332 ( \45709 , \45708 , \45202 );
buf \U$45333 ( \45710 , \45709 );
buf \U$45334 ( \45711 , \27285 );
not \U$45335 ( \45712 , \45711 );
not \U$45336 ( \45713 , \26907 );
not \U$45337 ( \45714 , \26101 );
not \U$45338 ( \45715 , \45608 );
or \U$45339 ( \45716 , \45714 , \45715 );
not \U$45340 ( \45717 , \44755 );
buf \U$45341 ( \45718 , \44753 );
not \U$45342 ( \45719 , \45718 );
or \U$45343 ( \45720 , \45717 , \45719 );
not \U$45344 ( \45721 , \44720 );
nand \U$45345 ( \45722 , \45720 , \45721 );
not \U$45346 ( \45723 , \45722 );
nand \U$45347 ( \45724 , \45716 , \45723 );
not \U$45348 ( \45725 , \45724 );
or \U$45349 ( \45726 , \45713 , \45725 );
not \U$45350 ( \45727 , \44732 );
nand \U$45351 ( \45728 , \45726 , \45727 );
not \U$45352 ( \45729 , \45728 );
or \U$45353 ( \45730 , \45712 , \45729 );
not \U$45354 ( \45731 , \44737 );
nand \U$45355 ( \45732 , \45730 , \45731 );
not \U$45356 ( \45733 , \45732 );
nand \U$45357 ( \45734 , \44722 , \44738 );
not \U$45358 ( \45735 , \45734 );
and \U$45359 ( \45736 , \45733 , \45735 );
and \U$45360 ( \45737 , \45732 , \45734 );
nor \U$45361 ( \45738 , \45736 , \45737 );
nor \U$45362 ( \45739 , \45738 , \45204 );
buf \U$45363 ( \45740 , \45739 );
not \U$45364 ( \45741 , \45728 );
nand \U$45365 ( \45742 , \45731 , \45711 );
not \U$45366 ( \45743 , \45742 );
and \U$45367 ( \45744 , \45741 , \45743 );
and \U$45368 ( \45745 , \45728 , \45742 );
nor \U$45369 ( \45746 , \45744 , \45745 );
nor \U$45370 ( \45747 , \45746 , \45204 );
buf \U$45371 ( \45748 , \45747 );
buf \U$45372 ( \45749 , \26905 );
not \U$45373 ( \45750 , \45749 );
not \U$45374 ( \45751 , \45724 );
or \U$45375 ( \45752 , \45750 , \45751 );
not \U$45376 ( \45753 , \44727 );
nand \U$45377 ( \45754 , \45752 , \45753 );
not \U$45378 ( \45755 , \45754 );
nor \U$45379 ( \45756 , \44730 , \44729 );
not \U$45380 ( \45757 , \45756 );
nand \U$45381 ( \45758 , \45757 , \44731 );
not \U$45382 ( \45759 , \45758 );
and \U$45383 ( \45760 , \45755 , \45759 );
and \U$45384 ( \45761 , \45754 , \45758 );
nor \U$45385 ( \45762 , \45760 , \45761 );
nor \U$45386 ( \45763 , \45762 , \45204 );
buf \U$45387 ( \45764 , \45763 );
nand \U$45388 ( \45765 , \45749 , \45753 );
xor \U$45389 ( \45766 , \45724 , \45765 );
nor \U$45390 ( \45767 , \45766 , \45202 );
buf \U$45391 ( \45768 , \45767 );
buf \U$45392 ( \45769 , \25648 );
not \U$45393 ( \45770 , \45769 );
buf \U$45394 ( \45771 , \45608 );
not \U$45395 ( \45772 , \45771 );
buf \U$45396 ( \45773 , \25671 );
buf \U$45397 ( \45774 , \26100 );
nand \U$45398 ( \45775 , \45773 , \45774 );
nor \U$45399 ( \45776 , \45772 , \45775 );
not \U$45400 ( \45777 , \45776 );
or \U$45401 ( \45778 , \45770 , \45777 );
not \U$45402 ( \45779 , \45718 );
nand \U$45403 ( \45780 , \45778 , \45779 );
not \U$45404 ( \45781 , \45780 );
not \U$45405 ( \45782 , \44720 );
nand \U$45406 ( \45783 , \45782 , \44755 );
not \U$45407 ( \45784 , \45783 );
and \U$45408 ( \45785 , \45781 , \45784 );
and \U$45409 ( \45786 , \45780 , \45783 );
nor \U$45410 ( \45787 , \45785 , \45786 );
nor \U$45411 ( \45788 , \45787 , \45204 );
buf \U$45412 ( \45789 , \45788 );
not \U$45413 ( \45790 , \45775 );
not \U$45414 ( \45791 , \45790 );
not \U$45415 ( \45792 , \45771 );
or \U$45416 ( \45793 , \45791 , \45792 );
not \U$45417 ( \45794 , \44749 );
nand \U$45418 ( \45795 , \45793 , \45794 );
nand \U$45419 ( \45796 , \44752 , \45769 );
and \U$45420 ( \45797 , \45795 , \45796 );
not \U$45421 ( \45798 , \45795 );
not \U$45422 ( \45799 , \45796 );
and \U$45423 ( \45800 , \45798 , \45799 );
nor \U$45424 ( \45801 , \45797 , \45800 );
nor \U$45425 ( \45802 , \45801 , \45204 );
buf \U$45426 ( \45803 , \45802 );
not \U$45427 ( \45804 , \45774 );
or \U$45428 ( \45805 , \45772 , \45804 );
buf \U$45429 ( \45806 , \44743 );
nand \U$45430 ( \45807 , \45805 , \45806 );
not \U$45431 ( \45808 , \45807 );
nand \U$45432 ( \45809 , \44748 , \45773 );
not \U$45433 ( \45810 , \45809 );
and \U$45434 ( \45811 , \45808 , \45810 );
and \U$45435 ( \45812 , \45807 , \45809 );
nor \U$45436 ( \45813 , \45811 , \45812 );
nor \U$45437 ( \45814 , \45813 , \45202 );
buf \U$45438 ( \45815 , \45814 );
nand \U$45439 ( \45816 , \45806 , \45774 );
not \U$45440 ( \45817 , \45816 );
and \U$45441 ( \45818 , \45772 , \45817 );
not \U$45442 ( \45819 , \45772 );
and \U$45443 ( \45820 , \45819 , \45816 );
nor \U$45444 ( \45821 , \45818 , \45820 );
nor \U$45445 ( \45822 , \45821 , \45202 );
buf \U$45446 ( \45823 , \45822 );
buf \U$45447 ( \45824 , \22305 );
not \U$45448 ( \45825 , \45824 );
not \U$45449 ( \45826 , \45825 );
not \U$45450 ( \45827 , \21306 );
buf \U$45451 ( \45828 , \44681 );
nor \U$45452 ( \45829 , \45827 , \45828 );
not \U$45453 ( \45830 , \45829 );
not \U$45454 ( \45831 , \45604 );
not \U$45455 ( \45832 , \45605 );
not \U$45456 ( \45833 , \44634 );
or \U$45457 ( \45834 , \45832 , \45833 );
not \U$45458 ( \45835 , \44675 );
nand \U$45459 ( \45836 , \45834 , \45835 );
not \U$45460 ( \45837 , \45836 );
or \U$45461 ( \45838 , \45831 , \45837 );
buf \U$45462 ( \45839 , \15919 );
not \U$45463 ( \45840 , \45839 );
not \U$45464 ( \45841 , \44697 );
buf \U$45465 ( \45842 , \15929 );
not \U$45466 ( \45843 , \45842 );
or \U$45467 ( \45844 , \45841 , \45843 );
not \U$45468 ( \45845 , \44702 );
nand \U$45469 ( \45846 , \45844 , \45845 );
not \U$45470 ( \45847 , \45846 );
or \U$45471 ( \45848 , \45840 , \45847 );
nand \U$45472 ( \45849 , \45848 , \44705 );
not \U$45473 ( \45850 , \45849 );
nand \U$45474 ( \45851 , \45838 , \45850 );
not \U$45475 ( \45852 , \45851 );
or \U$45476 ( \45853 , \45830 , \45852 );
buf \U$45477 ( \45854 , \44684 );
nor \U$45478 ( \45855 , \45828 , \45854 );
not \U$45479 ( \45856 , \44686 );
nor \U$45480 ( \45857 , \45855 , \45856 );
nand \U$45481 ( \45858 , \45853 , \45857 );
not \U$45482 ( \45859 , \45858 );
or \U$45483 ( \45860 , \45826 , \45859 );
buf \U$45484 ( \45861 , \44689 );
nand \U$45485 ( \45862 , \45860 , \45861 );
not \U$45486 ( \45863 , \45862 );
not \U$45487 ( \45864 , \22802 );
nand \U$45488 ( \45865 , \45864 , \44712 );
not \U$45489 ( \45866 , \45865 );
and \U$45490 ( \45867 , \45863 , \45866 );
and \U$45491 ( \45868 , \45862 , \45865 );
nor \U$45492 ( \45869 , \45867 , \45868 );
nor \U$45493 ( \45870 , \45869 , \45204 );
buf \U$45494 ( \45871 , \45870 );
not \U$45495 ( \45872 , \45824 );
nand \U$45496 ( \45873 , \45872 , \45861 );
xor \U$45497 ( \45874 , \45858 , \45873 );
nor \U$45498 ( \45875 , \45874 , \45204 );
buf \U$45499 ( \45876 , \45875 );
not \U$45500 ( \45877 , \21306 );
not \U$45501 ( \45878 , \45851 );
or \U$45502 ( \45879 , \45877 , \45878 );
nand \U$45503 ( \45880 , \45879 , \45854 );
not \U$45504 ( \45881 , \45880 );
or \U$45505 ( \45882 , \45856 , \45828 );
not \U$45506 ( \45883 , \45882 );
and \U$45507 ( \45884 , \45881 , \45883 );
and \U$45508 ( \45885 , \45880 , \45882 );
nor \U$45509 ( \45886 , \45884 , \45885 );
nor \U$45510 ( \45887 , \45886 , \45204 );
buf \U$45511 ( \45888 , \45887 );
not \U$45512 ( \45889 , \45827 );
nand \U$45513 ( \45890 , \45889 , \45854 );
and \U$45514 ( \45891 , \45851 , \45890 );
not \U$45515 ( \45892 , \45851 );
not \U$45516 ( \45893 , \45890 );
and \U$45517 ( \45894 , \45892 , \45893 );
nor \U$45518 ( \45895 , \45891 , \45894 );
nor \U$45519 ( \45896 , \45895 , \45204 );
buf \U$45520 ( \45897 , \45896 );
buf \U$45521 ( \45898 , \14884 );
not \U$45522 ( \45899 , \45898 );
not \U$45523 ( \45900 , \45842 );
nor \U$45524 ( \45901 , \45899 , \45900 );
not \U$45525 ( \45902 , \45901 );
not \U$45526 ( \45903 , \45836 );
or \U$45527 ( \45904 , \45902 , \45903 );
not \U$45528 ( \45905 , \45846 );
nand \U$45529 ( \45906 , \45904 , \45905 );
nand \U$45530 ( \45907 , \44705 , \45839 );
and \U$45531 ( \45908 , \45906 , \45907 );
not \U$45532 ( \45909 , \45906 );
not \U$45533 ( \45910 , \45907 );
and \U$45534 ( \45911 , \45909 , \45910 );
nor \U$45535 ( \45912 , \45908 , \45911 );
nor \U$45536 ( \45913 , \45912 , \45204 );
buf \U$45537 ( \45914 , \45913 );
not \U$45538 ( \45915 , \45898 );
not \U$45539 ( \45916 , \45836 );
or \U$45540 ( \45917 , \45915 , \45916 );
nand \U$45541 ( \45918 , \45917 , \45841 );
not \U$45542 ( \45919 , \45900 );
nand \U$45543 ( \45920 , \45919 , \45845 );
and \U$45544 ( \45921 , \45918 , \45920 );
not \U$45545 ( \45922 , \45918 );
not \U$45546 ( \45923 , \45920 );
and \U$45547 ( \45924 , \45922 , \45923 );
nor \U$45548 ( \45925 , \45921 , \45924 );
nor \U$45549 ( \45926 , \45925 , \45204 );
buf \U$45550 ( \45927 , \45926 );
not \U$45551 ( \45928 , \14883 );
not \U$45552 ( \45929 , \45928 );
not \U$45553 ( \45930 , \45836 );
or \U$45554 ( \45931 , \45929 , \45930 );
buf \U$45555 ( \45932 , \44694 );
nand \U$45556 ( \45933 , \45931 , \45932 );
not \U$45557 ( \45934 , \14220 );
nand \U$45558 ( \45935 , \45934 , \44695 );
and \U$45559 ( \45936 , \45933 , \45935 );
not \U$45560 ( \45937 , \45933 );
not \U$45561 ( \45938 , \45935 );
and \U$45562 ( \45939 , \45937 , \45938 );
nor \U$45563 ( \45940 , \45936 , \45939 );
nor \U$45564 ( \45941 , \45940 , \45204 );
buf \U$45565 ( \45942 , \45941 );
nand \U$45566 ( \45943 , \45932 , \45928 );
xor \U$45567 ( \45944 , \45836 , \45943 );
nor \U$45568 ( \45945 , \45944 , \45202 );
buf \U$45569 ( \45946 , \45945 );
buf \U$45570 ( \45947 , \20771 );
not \U$45571 ( \45948 , \45947 );
not \U$45572 ( \45949 , \20761 );
not \U$45573 ( \45950 , \20589 );
buf \U$45574 ( \45951 , \44634 );
not \U$45575 ( \45952 , \45951 );
or \U$45576 ( \45953 , \45950 , \45952 );
not \U$45577 ( \45954 , \44654 );
nand \U$45578 ( \45955 , \45953 , \45954 );
not \U$45579 ( \45956 , \45955 );
or \U$45580 ( \45957 , \45949 , \45956 );
nand \U$45581 ( \45958 , \45957 , \44672 );
not \U$45582 ( \45959 , \45958 );
or \U$45583 ( \45960 , \45948 , \45959 );
not \U$45584 ( \45961 , \44660 );
nand \U$45585 ( \45962 , \45960 , \45961 );
not \U$45586 ( \45963 , \45962 );
not \U$45587 ( \45964 , \44662 );
nand \U$45588 ( \45965 , \44657 , \44658 );
nand \U$45589 ( \45966 , \45964 , \45965 );
not \U$45590 ( \45967 , \45966 );
and \U$45591 ( \45968 , \45963 , \45967 );
and \U$45592 ( \45969 , \45962 , \45966 );
nor \U$45593 ( \45970 , \45968 , \45969 );
nor \U$45594 ( \45971 , \45970 , \45204 );
buf \U$45595 ( \45972 , \45971 );
nand \U$45596 ( \45973 , \45947 , \45961 );
and \U$45597 ( \45974 , \45958 , \45973 );
not \U$45598 ( \45975 , \45958 );
not \U$45599 ( \45976 , \45973 );
and \U$45600 ( \45977 , \45975 , \45976 );
nor \U$45601 ( \45978 , \45974 , \45977 );
nor \U$45602 ( \45979 , \45978 , \45204 );
buf \U$45603 ( \45980 , \45979 );
buf \U$45604 ( \45981 , \20728 );
not \U$45605 ( \45982 , \45981 );
not \U$45606 ( \45983 , \45955 );
or \U$45607 ( \45984 , \45982 , \45983 );
not \U$45608 ( \45985 , \44664 );
nand \U$45609 ( \45986 , \45984 , \45985 );
nand \U$45610 ( \45987 , \44670 , \20759 );
and \U$45611 ( \45988 , \45986 , \45987 );
not \U$45612 ( \45989 , \45986 );
not \U$45613 ( \45990 , \45987 );
and \U$45614 ( \45991 , \45989 , \45990 );
nor \U$45615 ( \45992 , \45988 , \45991 );
nor \U$45616 ( \45993 , \45992 , \45202 );
buf \U$45617 ( \45994 , \45993 );
nand \U$45618 ( \45995 , \45981 , \45985 );
and \U$45619 ( \45996 , \45955 , \45995 );
not \U$45620 ( \45997 , \45955 );
not \U$45621 ( \45998 , \45995 );
and \U$45622 ( \45999 , \45997 , \45998 );
nor \U$45623 ( \46000 , \45996 , \45999 );
nor \U$45624 ( \46001 , \46000 , \45202 );
buf \U$45625 ( \46002 , \46001 );
not \U$45626 ( \46003 , \44644 );
not \U$45627 ( \46004 , \46003 );
buf \U$45628 ( \46005 , \19971 );
nand \U$45629 ( \46006 , \45951 , \46005 );
not \U$45630 ( \46007 , \46006 );
or \U$45631 ( \46008 , \46004 , \46007 );
buf \U$45632 ( \46009 , \20266 );
nand \U$45633 ( \46010 , \46008 , \46009 );
not \U$45634 ( \46011 , \20588 );
or \U$45635 ( \46012 , \46010 , \46011 );
nand \U$45636 ( \46013 , \46012 , \44649 );
not \U$45637 ( \46014 , \46013 );
nand \U$45638 ( \46015 , \44653 , \20569 );
not \U$45639 ( \46016 , \46015 );
and \U$45640 ( \46017 , \46014 , \46016 );
and \U$45641 ( \46018 , \46013 , \46015 );
nor \U$45642 ( \46019 , \46017 , \46018 );
nor \U$45643 ( \46020 , \46019 , \45202 );
buf \U$45644 ( \46021 , \46020 );
and \U$45645 ( \46022 , \44649 , \20588 );
xor \U$45646 ( \46023 , \46010 , \46022 );
nor \U$45647 ( \46024 , \46023 , \45204 );
buf \U$45648 ( \46025 , \46024 );
not \U$45649 ( \46026 , \46005 );
buf \U$45650 ( \46027 , \45951 );
not \U$45651 ( \46028 , \46027 );
or \U$45652 ( \46029 , \46026 , \46028 );
nand \U$45653 ( \46030 , \46029 , \44642 );
nand \U$45654 ( \46031 , \46009 , \44643 );
xor \U$45655 ( \46032 , \46030 , \46031 );
nor \U$45656 ( \46033 , \46032 , \45202 );
buf \U$45657 ( \46034 , \46033 );
and \U$45658 ( \46035 , \44642 , \46005 );
not \U$45659 ( \46036 , \46027 );
and \U$45660 ( \46037 , \46035 , \46036 );
not \U$45661 ( \46038 , \46035 );
and \U$45662 ( \46039 , \46038 , \46027 );
nor \U$45663 ( \46040 , \46037 , \46039 );
nor \U$45664 ( \46041 , \46040 , \45204 );
buf \U$45665 ( \46042 , \46041 );
buf \U$45666 ( \46043 , \35614 );
not \U$45667 ( \46044 , \46043 );
buf \U$45668 ( \46045 , \35643 );
and \U$45669 ( \46046 , \46045 , \35661 );
not \U$45670 ( \46047 , \46046 );
not \U$45671 ( \46048 , \35452 );
not \U$45672 ( \46049 , \44616 );
not \U$45673 ( \46050 , \46049 );
not \U$45674 ( \46051 , \44609 );
or \U$45675 ( \46052 , \46050 , \46051 );
not \U$45676 ( \46053 , \34369 );
nand \U$45677 ( \46054 , \46052 , \46053 );
not \U$45678 ( \46055 , \46054 );
or \U$45679 ( \46056 , \46048 , \46055 );
buf \U$45680 ( \46057 , \35474 );
nand \U$45681 ( \46058 , \46056 , \46057 );
not \U$45682 ( \46059 , \46058 );
or \U$45683 ( \46060 , \46047 , \46059 );
not \U$45684 ( \46061 , \44626 );
nand \U$45685 ( \46062 , \46060 , \46061 );
not \U$45686 ( \46063 , \46062 );
or \U$45687 ( \46064 , \46044 , \46063 );
not \U$45688 ( \46065 , \44627 );
nand \U$45689 ( \46066 , \46064 , \46065 );
not \U$45690 ( \46067 , \46066 );
nand \U$45691 ( \46068 , \44631 , \35652 );
not \U$45692 ( \46069 , \46068 );
and \U$45693 ( \46070 , \46067 , \46069 );
and \U$45694 ( \46071 , \46066 , \46068 );
nor \U$45695 ( \46072 , \46070 , \46071 );
or \U$45696 ( \46073 , \46072 , \45202 );
or \U$45697 ( \46074 , \45203 , \860 );
nand \U$45698 ( \46075 , \46073 , \46074 );
buf \U$45699 ( \46076 , \46075 );
nand \U$45700 ( \46077 , \46043 , \46065 );
xor \U$45701 ( \46078 , \46062 , \46077 );
or \U$45702 ( \46079 , \46078 , \45202 );
or \U$45703 ( \46080 , \45203 , \888 );
nand \U$45704 ( \46081 , \46079 , \46080 );
buf \U$45705 ( \46082 , \46081 );
not \U$45706 ( \46083 , \46045 );
not \U$45707 ( \46084 , \46058 );
or \U$45708 ( \46085 , \46083 , \46084 );
not \U$45709 ( \46086 , \44619 );
nand \U$45710 ( \46087 , \46085 , \46086 );
not \U$45711 ( \46088 , \46087 );
nand \U$45712 ( \46089 , \44625 , \35661 );
not \U$45713 ( \46090 , \46089 );
and \U$45714 ( \46091 , \46088 , \46090 );
and \U$45715 ( \46092 , \46087 , \46089 );
nor \U$45716 ( \46093 , \46091 , \46092 );
or \U$45717 ( \46094 , \46093 , \45202 );
or \U$45718 ( \46095 , \45203 , \1286 );
nand \U$45719 ( \46096 , \46094 , \46095 );
buf \U$45720 ( \46097 , \46096 );
not \U$45721 ( \46098 , \44619 );
nand \U$45722 ( \46099 , \46098 , \46045 );
xor \U$45723 ( \46100 , \46058 , \46099 );
or \U$45724 ( \46101 , \46100 , \45204 );
or \U$45725 ( \46102 , \45203 , \922 );
nand \U$45726 ( \46103 , \46101 , \46102 );
buf \U$45727 ( \46104 , \46103 );
and \U$45728 ( \46105 , \45204 , \1066 );
not \U$45729 ( \46106 , \45204 );
not \U$45730 ( \46107 , \35450 );
not \U$45731 ( \46108 , \35103 );
not \U$45732 ( \46109 , \46054 );
or \U$45733 ( \46110 , \46108 , \46109 );
nand \U$45734 ( \46111 , \35462 , \35464 );
nand \U$45735 ( \46112 , \46110 , \46111 );
not \U$45736 ( \46113 , \46112 );
or \U$45737 ( \46114 , \46107 , \46113 );
nand \U$45738 ( \46115 , \46114 , \35469 );
not \U$45739 ( \46116 , \46115 );
or \U$45740 ( \46117 , \35471 , \35466 );
not \U$45741 ( \46118 , \46117 );
and \U$45742 ( \46119 , \46116 , \46118 );
and \U$45743 ( \46120 , \46115 , \46117 );
nor \U$45744 ( \46121 , \46119 , \46120 );
and \U$45745 ( \46122 , \46106 , \46121 );
nor \U$45746 ( \46123 , \46105 , \46122 );
buf \U$45747 ( \46124 , \46123 );
and \U$45748 ( \46125 , \45202 , \1083 );
not \U$45749 ( \46126 , \45202 );
not \U$45750 ( \46127 , \46112 );
nand \U$45751 ( \46128 , \35469 , \35450 );
not \U$45752 ( \46129 , \46128 );
and \U$45753 ( \46130 , \46127 , \46129 );
and \U$45754 ( \46131 , \46112 , \46128 );
nor \U$45755 ( \46132 , \46130 , \46131 );
and \U$45756 ( \46133 , \46126 , \46132 );
nor \U$45757 ( \46134 , \46125 , \46133 );
buf \U$45758 ( \46135 , \46134 );
not \U$45759 ( \46136 , \35102 );
not \U$45760 ( \46137 , \46054 );
or \U$45761 ( \46138 , \46136 , \46137 );
buf \U$45762 ( \46139 , \35461 );
nand \U$45763 ( \46140 , \46138 , \46139 );
not \U$45764 ( \46141 , \35457 );
not \U$45765 ( \46142 , \35455 );
or \U$45766 ( \46143 , \46141 , \46142 );
nand \U$45767 ( \46144 , \46143 , \35464 );
xor \U$45768 ( \46145 , \46140 , \46144 );
or \U$45769 ( \46146 , \46145 , \45202 );
or \U$45770 ( \46147 , \45203 , \1132 );
nand \U$45771 ( \46148 , \46146 , \46147 );
buf \U$45772 ( \46149 , \46148 );
not \U$45773 ( \46150 , \46054 );
nand \U$45774 ( \46151 , \46139 , \35102 );
not \U$45775 ( \46152 , \46151 );
and \U$45776 ( \46153 , \46150 , \46152 );
and \U$45777 ( \46154 , \46054 , \46151 );
nor \U$45778 ( \46155 , \46153 , \46154 );
or \U$45779 ( \46156 , \46155 , \45202 );
or \U$45780 ( \46157 , \45203 , \793 );
nand \U$45781 ( \46158 , \46156 , \46157 );
buf \U$45782 ( \46159 , \46158 );
buf \U$45783 ( \46160 , \32278 );
not \U$45784 ( \46161 , \46160 );
not \U$45785 ( \46162 , \32287 );
not \U$45786 ( \46163 , \44614 );
not \U$45787 ( \46164 , \37028 );
not \U$45788 ( \46165 , \40812 );
or \U$45789 ( \46166 , \46164 , \46165 );
buf \U$45790 ( \46167 , \44608 );
nand \U$45791 ( \46168 , \46166 , \46167 );
not \U$45792 ( \46169 , \46168 );
or \U$45793 ( \46170 , \46163 , \46169 );
buf \U$45794 ( \46171 , \34366 );
nand \U$45795 ( \46172 , \34363 , \46171 );
nand \U$45796 ( \46173 , \46170 , \46172 );
not \U$45797 ( \46174 , \46173 );
or \U$45798 ( \46175 , \46162 , \46174 );
buf \U$45799 ( \46176 , \31214 );
and \U$45800 ( \46177 , \31210 , \46176 );
nand \U$45801 ( \46178 , \46175 , \46177 );
not \U$45802 ( \46179 , \46178 );
or \U$45803 ( \46180 , \46161 , \46179 );
not \U$45804 ( \46181 , \31759 );
not \U$45805 ( \46182 , \46181 );
nand \U$45806 ( \46183 , \46180 , \46182 );
nand \U$45807 ( \46184 , \32280 , \32283 );
xor \U$45808 ( \46185 , \46183 , \46184 );
or \U$45809 ( \46186 , \46185 , \45202 );
or \U$45810 ( \46187 , \45203 , \1039 );
nand \U$45811 ( \46188 , \46186 , \46187 );
buf \U$45812 ( \46189 , \46188 );
not \U$45813 ( \46190 , \46178 );
not \U$45814 ( \46191 , \46181 );
nand \U$45815 ( \46192 , \46191 , \46160 );
not \U$45816 ( \46193 , \46192 );
and \U$45817 ( \46194 , \46190 , \46193 );
and \U$45818 ( \46195 , \46178 , \46192 );
nor \U$45819 ( \46196 , \46194 , \46195 );
or \U$45820 ( \46197 , \46196 , \45202 );
or \U$45821 ( \46198 , \45203 , \1046 );
nand \U$45822 ( \46199 , \46197 , \46198 );
buf \U$45823 ( \46200 , \46199 );
buf \U$45824 ( \46201 , \32286 );
not \U$45825 ( \46202 , \46201 );
not \U$45826 ( \46203 , \46173 );
or \U$45827 ( \46204 , \46202 , \46203 );
not \U$45828 ( \46205 , \31209 );
nand \U$45829 ( \46206 , \46204 , \46205 );
not \U$45830 ( \46207 , \46206 );
nand \U$45831 ( \46208 , \46176 , \31177 );
not \U$45832 ( \46209 , \46208 );
and \U$45833 ( \46210 , \46207 , \46209 );
and \U$45834 ( \46211 , \46206 , \46208 );
nor \U$45835 ( \46212 , \46210 , \46211 );
or \U$45836 ( \46213 , \46212 , \45202 );
or \U$45837 ( \46214 , \45203 , \997 );
nand \U$45838 ( \46215 , \46213 , \46214 );
buf \U$45839 ( \46216 , \46215 );
not \U$45840 ( \46217 , \46173 );
nand \U$45841 ( \46218 , \46201 , \46205 );
not \U$45842 ( \46219 , \46218 );
and \U$45843 ( \46220 , \46217 , \46219 );
and \U$45844 ( \46221 , \46173 , \46218 );
nor \U$45845 ( \46222 , \46220 , \46221 );
or \U$45846 ( \46223 , \46222 , \45204 );
or \U$45847 ( \46224 , \45203 , \1004 );
nand \U$45848 ( \46225 , \46223 , \46224 );
buf \U$45849 ( \46226 , \46225 );
not \U$45850 ( \46227 , \34341 );
not \U$45851 ( \46228 , \46227 );
buf \U$45852 ( \46229 , \44610 );
nand \U$45853 ( \46230 , \46168 , \46229 );
not \U$45854 ( \46231 , \34305 );
or \U$45855 ( \46232 , \46230 , \46231 );
buf \U$45856 ( \46233 , \34306 );
nand \U$45857 ( \46234 , \46232 , \46233 );
not \U$45858 ( \46235 , \46234 );
or \U$45859 ( \46236 , \46228 , \46235 );
buf \U$45860 ( \46237 , \34361 );
nand \U$45861 ( \46238 , \46236 , \46237 );
not \U$45862 ( \46239 , \46238 );
nand \U$45863 ( \46240 , \34360 , \46171 );
not \U$45864 ( \46241 , \46240 );
and \U$45865 ( \46242 , \46239 , \46241 );
and \U$45866 ( \46243 , \46238 , \46240 );
nor \U$45867 ( \46244 , \46242 , \46243 );
or \U$45868 ( \46245 , \46244 , \45204 );
or \U$45869 ( \46246 , \45203 , \1503 );
nand \U$45870 ( \46247 , \46245 , \46246 );
buf \U$45871 ( \46248 , \46247 );
not \U$45872 ( \46249 , \46234 );
not \U$45873 ( \46250 , \34341 );
nand \U$45874 ( \46251 , \46250 , \46237 );
not \U$45875 ( \46252 , \46251 );
and \U$45876 ( \46253 , \46249 , \46252 );
and \U$45877 ( \46254 , \46234 , \46251 );
nor \U$45878 ( \46255 , \46253 , \46254 );
or \U$45879 ( \46256 , \46255 , \45202 );
or \U$45880 ( \46257 , \45203 , \1493 );
nand \U$45881 ( \46258 , \46256 , \46257 );
buf \U$45882 ( \46259 , \46258 );
not \U$45883 ( \46260 , \46229 );
not \U$45884 ( \46261 , \46168 );
or \U$45885 ( \46262 , \46260 , \46261 );
not \U$45886 ( \46263 , \34303 );
nand \U$45887 ( \46264 , \46262 , \46263 );
not \U$45888 ( \46265 , \33647 );
nand \U$45889 ( \46266 , \46265 , \34305 );
xor \U$45890 ( \46267 , \46264 , \46266 );
or \U$45891 ( \46268 , \46267 , \45202 );
or \U$45892 ( \46269 , \45203 , \1902 );
nand \U$45893 ( \46270 , \46268 , \46269 );
buf \U$45894 ( \46271 , \46270 );
nand \U$45895 ( \46272 , \46263 , \46229 );
xor \U$45896 ( \46273 , \46168 , \46272 );
or \U$45897 ( \46274 , \46273 , \45202 );
or \U$45898 ( \46275 , \45203 , \1905 );
nand \U$45899 ( \46276 , \46274 , \46275 );
buf \U$45900 ( \46277 , \46276 );
buf \U$45901 ( \46278 , \36305 );
not \U$45902 ( \46279 , \46278 );
not \U$45903 ( \46280 , \36625 );
not \U$45904 ( \46281 , \37026 );
not \U$45905 ( \46282 , \38648 );
not \U$45906 ( \46283 , \40833 );
nand \U$45907 ( \46284 , \44606 , \46283 , \40786 , \39533 );
nand \U$45908 ( \46285 , \46284 , \40787 , \40790 );
not \U$45909 ( \46286 , \46285 );
or \U$45910 ( \46287 , \46282 , \46286 );
nand \U$45911 ( \46288 , \46287 , \40811 );
not \U$45912 ( \46289 , \46288 );
or \U$45913 ( \46290 , \46281 , \46289 );
not \U$45914 ( \46291 , \40817 );
nand \U$45915 ( \46292 , \46290 , \46291 );
not \U$45916 ( \46293 , \46292 );
or \U$45917 ( \46294 , \46280 , \46293 );
buf \U$45918 ( \46295 , \40816 );
not \U$45919 ( \46296 , \46295 );
nand \U$45920 ( \46297 , \46294 , \46296 );
not \U$45921 ( \46298 , \46297 );
or \U$45922 ( \46299 , \46279 , \46298 );
nand \U$45923 ( \46300 , \46299 , \40821 );
nand \U$45924 ( \46301 , \40824 , \36314 );
xor \U$45925 ( \46302 , \46300 , \46301 );
or \U$45926 ( \46303 , \46302 , \45202 );
or \U$45927 ( \46304 , \45203 , \2056 );
nand \U$45928 ( \46305 , \46303 , \46304 );
buf \U$45929 ( \46306 , \46305 );
nand \U$45930 ( \46307 , \46278 , \40821 );
xor \U$45931 ( \46308 , \46297 , \46307 );
or \U$45932 ( \46309 , \46308 , \45202 );
or \U$45933 ( \46310 , \45203 , \2057 );
nand \U$45934 ( \46311 , \46309 , \46310 );
buf \U$45935 ( \46312 , \46311 );
not \U$45936 ( \46313 , \46295 );
nand \U$45937 ( \46314 , \46313 , \36625 );
xor \U$45938 ( \46315 , \46292 , \46314 );
or \U$45939 ( \46316 , \46315 , \45202 );
or \U$45940 ( \46317 , \45203 , \3147 );
nand \U$45941 ( \46318 , \46316 , \46317 );
buf \U$45942 ( \46319 , \46318 );
not \U$45943 ( \46320 , \40817 );
nand \U$45944 ( \46321 , \46320 , \37026 );
xor \U$45945 ( \46322 , \46288 , \46321 );
or \U$45946 ( \46323 , \46322 , \45202 );
or \U$45947 ( \46324 , \45203 , \1816 );
nand \U$45948 ( \46325 , \46323 , \46324 );
buf \U$45949 ( \46326 , \46325 );
buf \U$45950 ( \46327 , \40794 );
not \U$45951 ( \46328 , \46327 );
buf \U$45952 ( \46329 , \38194 );
not \U$45953 ( \46330 , \46329 );
not \U$45954 ( \46331 , \46285 );
not \U$45955 ( \46332 , \38646 );
nor \U$45956 ( \46333 , \46331 , \46332 );
not \U$45957 ( \46334 , \46333 );
or \U$45958 ( \46335 , \46330 , \46334 );
not \U$45959 ( \46336 , \40803 );
nand \U$45960 ( \46337 , \46335 , \46336 );
not \U$45961 ( \46338 , \46337 );
or \U$45962 ( \46339 , \46328 , \46338 );
not \U$45963 ( \46340 , \40807 );
nand \U$45964 ( \46341 , \46339 , \46340 );
not \U$45965 ( \46342 , \46341 );
not \U$45966 ( \46343 , \40806 );
nand \U$45967 ( \46344 , \46343 , \40810 );
not \U$45968 ( \46345 , \46344 );
and \U$45969 ( \46346 , \46342 , \46345 );
and \U$45970 ( \46347 , \46341 , \46344 );
nor \U$45971 ( \46348 , \46346 , \46347 );
or \U$45972 ( \46349 , \46348 , \45202 );
or \U$45973 ( \46350 , \45203 , \2268 );
nand \U$45974 ( \46351 , \46349 , \46350 );
buf \U$45975 ( \46352 , \46351 );
not \U$45976 ( \46353 , \46337 );
not \U$45977 ( \46354 , \40807 );
nand \U$45978 ( \46355 , \46354 , \46327 );
not \U$45979 ( \46356 , \46355 );
and \U$45980 ( \46357 , \46353 , \46356 );
and \U$45981 ( \46358 , \46337 , \46355 );
nor \U$45982 ( \46359 , \46357 , \46358 );
or \U$45983 ( \46360 , \46359 , \45202 );
or \U$45984 ( \46361 , \45203 , \2246 );
nand \U$45985 ( \46362 , \46360 , \46361 );
buf \U$45986 ( \46363 , \46362 );
not \U$45987 ( \46364 , \38646 );
not \U$45988 ( \46365 , \46331 );
not \U$45989 ( \46366 , \46365 );
or \U$45990 ( \46367 , \46364 , \46366 );
not \U$45991 ( \46368 , \40797 );
nand \U$45992 ( \46369 , \46367 , \46368 );
nand \U$45993 ( \46370 , \40802 , \46329 );
and \U$45994 ( \46371 , \46369 , \46370 );
not \U$45995 ( \46372 , \46369 );
not \U$45996 ( \46373 , \46370 );
and \U$45997 ( \46374 , \46372 , \46373 );
nor \U$45998 ( \46375 , \46371 , \46374 );
or \U$45999 ( \46376 , \46375 , \45202 );
or \U$46000 ( \46377 , \45203 , \4653 );
nand \U$46001 ( \46378 , \46376 , \46377 );
buf \U$46002 ( \46379 , \46378 );
not \U$46003 ( \46380 , \40797 );
nand \U$46004 ( \46381 , \46380 , \38646 );
xor \U$46005 ( \46382 , \46365 , \46381 );
or \U$46006 ( \46383 , \46382 , \45202 );
or \U$46007 ( \46384 , \45203 , \2184 );
nand \U$46008 ( \46385 , \46383 , \46384 );
buf \U$46009 ( \46386 , \46385 );
not \U$46010 ( \46387 , \40784 );
not \U$46011 ( \46388 , \39533 );
not \U$46012 ( \46389 , \46283 );
not \U$46013 ( \46390 , \44606 );
or \U$46014 ( \46391 , \46389 , \46390 );
not \U$46015 ( \46392 , \40733 );
nand \U$46016 ( \46393 , \46391 , \46392 );
not \U$46017 ( \46394 , \46393 );
or \U$46018 ( \46395 , \46388 , \46394 );
and \U$46019 ( \46396 , \40738 , \40776 );
nand \U$46020 ( \46397 , \46395 , \46396 );
not \U$46021 ( \46398 , \46397 );
or \U$46022 ( \46399 , \46387 , \46398 );
buf \U$46023 ( \46400 , \40773 );
nand \U$46024 ( \46401 , \46399 , \46400 );
not \U$46025 ( \46402 , \46401 );
not \U$46026 ( \46403 , \40789 );
nand \U$46027 ( \46404 , \46403 , \40781 );
not \U$46028 ( \46405 , \46404 );
and \U$46029 ( \46406 , \46402 , \46405 );
and \U$46030 ( \46407 , \46401 , \46404 );
nor \U$46031 ( \46408 , \46406 , \46407 );
or \U$46032 ( \46409 , \46408 , \45202 );
or \U$46033 ( \46410 , \45203 , \3039 );
nand \U$46034 ( \46411 , \46409 , \46410 );
buf \U$46035 ( \46412 , \46411 );
not \U$46036 ( \46413 , \46397 );
nand \U$46037 ( \46414 , \40784 , \46400 );
not \U$46038 ( \46415 , \46414 );
and \U$46039 ( \46416 , \46413 , \46415 );
and \U$46040 ( \46417 , \46397 , \46414 );
nor \U$46041 ( \46418 , \46416 , \46417 );
or \U$46042 ( \46419 , \46418 , \45202 );
or \U$46043 ( \46420 , \45203 , \1926 );
nand \U$46044 ( \46421 , \46419 , \46420 );
buf \U$46045 ( \46422 , \46421 );
not \U$46046 ( \46423 , \39475 );
not \U$46047 ( \46424 , \46393 );
or \U$46048 ( \46425 , \46423 , \46424 );
buf \U$46049 ( \46426 , \40736 );
nand \U$46050 ( \46427 , \46425 , \46426 );
not \U$46051 ( \46428 , \46427 );
nand \U$46052 ( \46429 , \40776 , \39532 );
not \U$46053 ( \46430 , \46429 );
and \U$46054 ( \46431 , \46428 , \46430 );
and \U$46055 ( \46432 , \46427 , \46429 );
nor \U$46056 ( \46433 , \46431 , \46432 );
or \U$46057 ( \46434 , \46433 , \45202 );
or \U$46058 ( \46435 , \45203 , \21036 );
nand \U$46059 ( \46436 , \46434 , \46435 );
buf \U$46060 ( \46437 , \46436 );
nand \U$46061 ( \46438 , \39475 , \46426 );
and \U$46062 ( \46439 , \46393 , \46438 );
not \U$46063 ( \46440 , \46393 );
not \U$46064 ( \46441 , \46438 );
and \U$46065 ( \46442 , \46440 , \46441 );
nor \U$46066 ( \46443 , \46439 , \46442 );
or \U$46067 ( \46444 , \46443 , \45202 );
or \U$46068 ( \46445 , \45203 , \2335 );
nand \U$46069 ( \46446 , \46444 , \46445 );
buf \U$46070 ( \46447 , \46446 );
not \U$46071 ( \46448 , \40177 );
not \U$46072 ( \46449 , \40831 );
nand \U$46073 ( \46450 , \44606 , \46449 );
or \U$46074 ( \46451 , \46450 , \40828 );
buf \U$46075 ( \46452 , \40727 );
nand \U$46076 ( \46453 , \46451 , \46452 );
not \U$46077 ( \46454 , \46453 );
or \U$46078 ( \46455 , \46448 , \46454 );
buf \U$46079 ( \46456 , \40191 );
nand \U$46080 ( \46457 , \46455 , \46456 );
not \U$46081 ( \46458 , \46457 );
nand \U$46082 ( \46459 , \40189 , \40732 );
not \U$46083 ( \46460 , \46459 );
and \U$46084 ( \46461 , \46458 , \46460 );
and \U$46085 ( \46462 , \46457 , \46459 );
nor \U$46086 ( \46463 , \46461 , \46462 );
or \U$46087 ( \46464 , \46463 , \45202 );
or \U$46088 ( \46465 , \45203 , \1997 );
nand \U$46089 ( \46466 , \46464 , \46465 );
buf \U$46090 ( \46467 , \46466 );
not \U$46091 ( \46468 , \46453 );
nand \U$46092 ( \46469 , \46456 , \40177 );
not \U$46093 ( \46470 , \46469 );
and \U$46094 ( \46471 , \46468 , \46470 );
and \U$46095 ( \46472 , \46453 , \46469 );
nor \U$46096 ( \46473 , \46471 , \46472 );
or \U$46097 ( \46474 , \46473 , \45202 );
or \U$46098 ( \46475 , \45203 , \1981 );
nand \U$46099 ( \46476 , \46474 , \46475 );
buf \U$46100 ( \46477 , \46476 );
nand \U$46101 ( \46478 , \46450 , \40721 );
nand \U$46102 ( \46479 , \40726 , \40434 );
and \U$46103 ( \46480 , \46478 , \46479 );
not \U$46104 ( \46481 , \46478 );
not \U$46105 ( \46482 , \46479 );
and \U$46106 ( \46483 , \46481 , \46482 );
nor \U$46107 ( \46484 , \46480 , \46483 );
or \U$46108 ( \46485 , \46484 , \45202 );
or \U$46109 ( \46486 , \45203 , \2504 );
nand \U$46110 ( \46487 , \46485 , \46486 );
buf \U$46111 ( \46488 , \46487 );
nand \U$46112 ( \46489 , \40721 , \46449 );
xor \U$46113 ( \46490 , \44606 , \46489 );
or \U$46114 ( \46491 , \46490 , \45202 );
or \U$46115 ( \46492 , \45203 , \2427 );
nand \U$46116 ( \46493 , \46491 , \46492 );
buf \U$46117 ( \46494 , \46493 );
not \U$46118 ( \46495 , \44578 );
nor \U$46119 ( \46496 , \46495 , \44588 );
not \U$46120 ( \46497 , \46496 );
buf \U$46121 ( \46498 , \44421 );
not \U$46122 ( \46499 , \46498 );
or \U$46123 ( \46500 , \46497 , \46499 );
not \U$46124 ( \46501 , \44598 );
nand \U$46125 ( \46502 , \46500 , \46501 );
not \U$46126 ( \46503 , \46502 );
not \U$46127 ( \46504 , \44592 );
or \U$46128 ( \46505 , \46503 , \46504 );
nand \U$46129 ( \46506 , \46505 , \44601 );
not \U$46130 ( \46507 , \46506 );
not \U$46131 ( \46508 , \44605 );
not \U$46132 ( \46509 , \46508 );
nand \U$46133 ( \46510 , \46509 , \44550 );
not \U$46134 ( \46511 , \46510 );
and \U$46135 ( \46512 , \46507 , \46511 );
and \U$46136 ( \46513 , \46506 , \46510 );
nor \U$46137 ( \46514 , \46512 , \46513 );
or \U$46138 ( \46515 , \46514 , \45202 );
or \U$46139 ( \46516 , \45203 , \10584 );
nand \U$46140 ( \46517 , \46515 , \46516 );
buf \U$46141 ( \46518 , \46517 );
nand \U$46142 ( \46519 , \44601 , \44592 );
and \U$46143 ( \46520 , \46502 , \46519 );
not \U$46144 ( \46521 , \46502 );
not \U$46145 ( \46522 , \46519 );
and \U$46146 ( \46523 , \46521 , \46522 );
nor \U$46147 ( \46524 , \46520 , \46523 );
or \U$46148 ( \46525 , \46524 , \45202 );
or \U$46149 ( \46526 , \45203 , \2407 );
nand \U$46150 ( \46527 , \46525 , \46526 );
buf \U$46151 ( \46528 , \46527 );
not \U$46152 ( \46529 , \44578 );
not \U$46153 ( \46530 , \46498 );
or \U$46154 ( \46531 , \46529 , \46530 );
nand \U$46155 ( \46532 , \46531 , \44595 );
nand \U$46156 ( \46533 , \44597 , \44589 );
and \U$46157 ( \46534 , \46532 , \46533 );
not \U$46158 ( \46535 , \46532 );
not \U$46159 ( \46536 , \46533 );
and \U$46160 ( \46537 , \46535 , \46536 );
nor \U$46161 ( \46538 , \46534 , \46537 );
or \U$46162 ( \46539 , \46538 , \45202 );
or \U$46163 ( \46540 , \45203 , \11755 );
nand \U$46164 ( \46541 , \46539 , \46540 );
buf \U$46165 ( \46542 , \46541 );
nand \U$46166 ( \46543 , \44595 , \44578 );
and \U$46167 ( \46544 , \46498 , \46543 );
not \U$46168 ( \46545 , \46498 );
not \U$46169 ( \46546 , \46543 );
and \U$46170 ( \46547 , \46545 , \46546 );
nor \U$46171 ( \46548 , \46544 , \46547 );
or \U$46172 ( \46549 , \46548 , \45202 );
or \U$46173 ( \46550 , \45203 , \4151 );
nand \U$46174 ( \46551 , \46549 , \46550 );
buf \U$46175 ( \46552 , \46551 );
not \U$46176 ( \46553 , \44348 );
not \U$46177 ( \46554 , \44400 );
buf \U$46178 ( \46555 , \43627 );
not \U$46179 ( \46556 , \46555 );
or \U$46180 ( \46557 , \46554 , \46556 );
not \U$46181 ( \46558 , \44411 );
nand \U$46182 ( \46559 , \46557 , \46558 );
not \U$46183 ( \46560 , \46559 );
or \U$46184 ( \46561 , \46553 , \46560 );
buf \U$46185 ( \46562 , \44416 );
nand \U$46186 ( \46563 , \46561 , \46562 );
not \U$46187 ( \46564 , \46563 );
not \U$46188 ( \46565 , \44420 );
not \U$46189 ( \46566 , \46565 );
nand \U$46190 ( \46567 , \46566 , \44285 );
not \U$46191 ( \46568 , \46567 );
and \U$46192 ( \46569 , \46564 , \46568 );
and \U$46193 ( \46570 , \46563 , \46567 );
nor \U$46194 ( \46571 , \46569 , \46570 );
or \U$46195 ( \46572 , \46571 , \45202 );
or \U$46196 ( \46573 , \45203 , \4968 );
nand \U$46197 ( \46574 , \46572 , \46573 );
buf \U$46198 ( \46575 , \46574 );
nand \U$46199 ( \46576 , \46562 , \44348 );
and \U$46200 ( \46577 , \46559 , \46576 );
not \U$46201 ( \46578 , \46559 );
not \U$46202 ( \46579 , \46576 );
and \U$46203 ( \46580 , \46578 , \46579 );
nor \U$46204 ( \46581 , \46577 , \46580 );
or \U$46205 ( \46582 , \46581 , \45202 );
or \U$46206 ( \46583 , \45203 , \5030 );
nand \U$46207 ( \46584 , \46582 , \46583 );
buf \U$46208 ( \46585 , \46584 );
not \U$46209 ( \46586 , \44399 );
not \U$46210 ( \46587 , \46555 );
or \U$46211 ( \46588 , \46586 , \46587 );
not \U$46212 ( \46589 , \44405 );
nand \U$46213 ( \46590 , \46588 , \46589 );
not \U$46214 ( \46591 , \46590 );
nand \U$46215 ( \46592 , \44388 , \44410 );
not \U$46216 ( \46593 , \46592 );
and \U$46217 ( \46594 , \46591 , \46593 );
and \U$46218 ( \46595 , \46590 , \46592 );
nor \U$46219 ( \46596 , \46594 , \46595 );
or \U$46220 ( \46597 , \46596 , \45202 );
or \U$46221 ( \46598 , \45203 , \12209 );
nand \U$46222 ( \46599 , \46597 , \46598 );
buf \U$46223 ( \46600 , \46599 );
xor \U$46224 ( \46601 , \44394 , \44398 );
not \U$46225 ( \46602 , \46601 );
and \U$46226 ( \46603 , \46555 , \46602 );
not \U$46227 ( \46604 , \46555 );
and \U$46228 ( \46605 , \46604 , \46601 );
nor \U$46229 ( \46606 , \46603 , \46605 );
or \U$46230 ( \46607 , \46606 , \45202 );
or \U$46231 ( \46608 , \45203 , \6189 );
nand \U$46232 ( \46609 , \46607 , \46608 );
buf \U$46233 ( \46610 , \46609 );
not \U$46234 ( \46611 , \43390 );
not \U$46235 ( \46612 , \43186 );
nand \U$46236 ( \46613 , \46612 , \43620 );
not \U$46237 ( \46614 , \46613 );
or \U$46238 ( \46615 , \46611 , \46614 );
not \U$46239 ( \46616 , \43623 );
not \U$46240 ( \46617 , \46616 );
nand \U$46241 ( \46618 , \46615 , \46617 );
nand \U$46242 ( \46619 , \43626 , \43614 );
and \U$46243 ( \46620 , \46618 , \46619 );
not \U$46244 ( \46621 , \46618 );
not \U$46245 ( \46622 , \46619 );
and \U$46246 ( \46623 , \46621 , \46622 );
nor \U$46247 ( \46624 , \46620 , \46623 );
or \U$46248 ( \46625 , \46624 , \45202 );
or \U$46249 ( \46626 , \45203 , \18027 );
nand \U$46250 ( \46627 , \46625 , \46626 );
buf \U$46251 ( \46628 , \46627 );
not \U$46252 ( \46629 , \46616 );
nand \U$46253 ( \46630 , \46629 , \43390 );
and \U$46254 ( \46631 , \46613 , \46630 );
not \U$46255 ( \46632 , \46613 );
not \U$46256 ( \46633 , \46630 );
and \U$46257 ( \46634 , \46632 , \46633 );
nor \U$46258 ( \46635 , \46631 , \46634 );
or \U$46259 ( \46636 , \46635 , \45202 );
or \U$46260 ( \46637 , \45203 , \9491 );
nand \U$46261 ( \46638 , \46636 , \46637 );
buf \U$46262 ( \46639 , \46638 );
not \U$46263 ( \46640 , \43185 );
buf \U$46264 ( \46641 , \42772 );
not \U$46265 ( \46642 , \46641 );
or \U$46266 ( \46643 , \46640 , \46642 );
buf \U$46267 ( \46644 , \43617 );
nand \U$46268 ( \46645 , \46643 , \46644 );
nand \U$46269 ( \46646 , \43171 , \43618 );
and \U$46270 ( \46647 , \46645 , \46646 );
not \U$46271 ( \46648 , \46645 );
not \U$46272 ( \46649 , \46646 );
and \U$46273 ( \46650 , \46648 , \46649 );
nor \U$46274 ( \46651 , \46647 , \46650 );
or \U$46275 ( \46652 , \46651 , \45202 );
or \U$46276 ( \46653 , \45203 , \12184 );
nand \U$46277 ( \46654 , \46652 , \46653 );
buf \U$46278 ( \46655 , \46654 );
nand \U$46279 ( \46656 , \46644 , \43185 );
and \U$46280 ( \46657 , \46656 , \46641 );
not \U$46281 ( \46658 , \46656 );
not \U$46282 ( \46659 , \46641 );
and \U$46283 ( \46660 , \46658 , \46659 );
nor \U$46284 ( \46661 , \46657 , \46660 );
or \U$46285 ( \46662 , \46661 , \45202 );
or \U$46286 ( \46663 , \45201 , \9782 );
nand \U$46287 ( \46664 , \46662 , \46663 );
buf \U$46288 ( \46665 , \46664 );
not \U$46289 ( \46666 , \41768 );
not \U$46290 ( \46667 , \42769 );
not \U$46291 ( \46668 , \42765 );
or \U$46292 ( \46669 , \46667 , \46668 );
nand \U$46293 ( \46670 , \46669 , \41601 );
not \U$46294 ( \46671 , \46670 );
or \U$46295 ( \46672 , \46666 , \46671 );
nand \U$46296 ( \46673 , \46672 , \41770 );
not \U$46297 ( \46674 , \42771 );
not \U$46298 ( \46675 , \46674 );
nand \U$46299 ( \46676 , \46675 , \41969 );
xor \U$46300 ( \46677 , \46673 , \46676 );
or \U$46301 ( \46678 , \46677 , \45202 );
or \U$46302 ( \46679 , \45201 , \11114 );
nand \U$46303 ( \46680 , \46678 , \46679 );
buf \U$46304 ( \46681 , \46680 );
not \U$46305 ( \46682 , \46670 );
nand \U$46306 ( \46683 , \41770 , \41768 );
not \U$46307 ( \46684 , \46683 );
and \U$46308 ( \46685 , \46682 , \46684 );
and \U$46309 ( \46686 , \46670 , \46683 );
nor \U$46310 ( \46687 , \46685 , \46686 );
or \U$46311 ( \46688 , \46687 , \45202 );
or \U$46312 ( \46689 , \45201 , \9680 );
nand \U$46313 ( \46690 , \46688 , \46689 );
buf \U$46314 ( \46691 , \46690 );
not \U$46315 ( \46692 , \42768 );
not \U$46316 ( \46693 , \42765 );
or \U$46317 ( \46694 , \46692 , \46693 );
nand \U$46318 ( \46695 , \46694 , \41595 );
not \U$46319 ( \46696 , \41479 );
not \U$46320 ( \46697 , \46696 );
nand \U$46321 ( \46698 , \46697 , \41600 );
xor \U$46322 ( \46699 , \46695 , \46698 );
or \U$46323 ( \46700 , \46699 , \45202 );
or \U$46324 ( \46701 , \45201 , \16469 );
nand \U$46325 ( \46702 , \46700 , \46701 );
buf \U$46326 ( \46703 , \46702 );
and \U$46327 ( \46704 , \45202 , \9640 );
not \U$46328 ( \46705 , \45202 );
nand \U$46329 ( \46706 , \42768 , \41595 );
xor \U$46330 ( \46707 , \42765 , \46706 );
and \U$46331 ( \46708 , \46705 , \46707 );
nor \U$46332 ( \46709 , \46704 , \46708 );
buf \U$46333 ( \46710 , \46709 );
buf \U$46334 ( \46711 , \42330 );
not \U$46335 ( \46712 , \46711 );
not \U$46336 ( \46713 , \42355 );
not \U$46337 ( \46714 , \42762 );
or \U$46338 ( \46715 , \46713 , \46714 );
not \U$46339 ( \46716 , \42301 );
nand \U$46340 ( \46717 , \46715 , \46716 );
not \U$46341 ( \46718 , \46717 );
or \U$46342 ( \46719 , \46712 , \46718 );
nand \U$46343 ( \46720 , \46719 , \42333 );
not \U$46344 ( \46721 , \42764 );
not \U$46345 ( \46722 , \46721 );
nand \U$46346 ( \46723 , \46722 , \42351 );
and \U$46347 ( \46724 , \46720 , \46723 );
not \U$46348 ( \46725 , \46720 );
not \U$46349 ( \46726 , \46723 );
and \U$46350 ( \46727 , \46725 , \46726 );
nor \U$46351 ( \46728 , \46724 , \46727 );
or \U$46352 ( \46729 , \46728 , \45202 );
or \U$46353 ( \46730 , \45201 , \10633 );
nand \U$46354 ( \46731 , \46729 , \46730 );
buf \U$46355 ( \46732 , \46731 );
nand \U$46356 ( \46733 , \46711 , \42333 );
and \U$46357 ( \46734 , \46717 , \46733 );
not \U$46358 ( \46735 , \46717 );
not \U$46359 ( \46736 , \46733 );
and \U$46360 ( \46737 , \46735 , \46736 );
nor \U$46361 ( \46738 , \46734 , \46737 );
or \U$46362 ( \46739 , \46738 , \45202 );
or \U$46363 ( \46740 , \45201 , \10628 );
nand \U$46364 ( \46741 , \46739 , \46740 );
buf \U$46365 ( \46742 , \46741 );
not \U$46366 ( \46743 , \42354 );
not \U$46367 ( \46744 , \46743 );
not \U$46368 ( \46745 , \42762 );
or \U$46369 ( \46746 , \46744 , \46745 );
nand \U$46370 ( \46747 , \46746 , \42298 );
not \U$46371 ( \46748 , \42234 );
nand \U$46372 ( \46749 , \46748 , \42300 );
and \U$46373 ( \46750 , \46747 , \46749 );
not \U$46374 ( \46751 , \46747 );
not \U$46375 ( \46752 , \46749 );
and \U$46376 ( \46753 , \46751 , \46752 );
nor \U$46377 ( \46754 , \46750 , \46753 );
or \U$46378 ( \46755 , \46754 , \45202 );
or \U$46379 ( \46756 , \45201 , \27628 );
nand \U$46380 ( \46757 , \46755 , \46756 );
buf \U$46381 ( \46758 , \46757 );
nand \U$46382 ( \46759 , \46743 , \42298 );
xor \U$46383 ( \46760 , \42762 , \46759 );
or \U$46384 ( \46761 , \46760 , \45202 );
or \U$46385 ( \46762 , \45201 , \10670 );
nand \U$46386 ( \46763 , \46761 , \46762 );
buf \U$46387 ( \46764 , \46763 );
not \U$46388 ( \46765 , \42757 );
and \U$46389 ( \46766 , \42745 , \46765 );
not \U$46390 ( \46767 , \42745 );
and \U$46391 ( \46768 , \46767 , \42757 );
nor \U$46392 ( \46769 , \46766 , \46768 );
or \U$46393 ( \46770 , \46769 , \45202 );
or \U$46394 ( \46771 , \45201 , \10658 );
nand \U$46395 ( \46772 , \46770 , \46771 );
buf \U$46396 ( \46773 , \46772 );
nand \U$46397 ( \46774 , \42744 , \42465 );
xor \U$46398 ( \46775 , \46774 , \42740 );
not \U$46399 ( \46776 , \45200 );
or \U$46400 ( \46777 , \46775 , \46776 );
or \U$46401 ( \46778 , \45201 , \9752 );
nand \U$46402 ( \46779 , \46777 , \46778 );
buf \U$46403 ( \46780 , \46779 );
nand \U$46404 ( \46781 , \42739 , \42514 );
xor \U$46405 ( \46782 , \46781 , \42734 );
or \U$46406 ( \46783 , \46782 , \46776 );
or \U$46407 ( \46784 , \45200 , \9749 );
nand \U$46408 ( \46785 , \46783 , \46784 );
buf \U$46409 ( \46786 , \46785 );
endmodule

