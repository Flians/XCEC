//
// Conformal-LEC Version 20.10-d213 (02-Sep-2020)
//
module top(RIbe29380_53,RIbe27d78_6,RIbe27ee0_9,RIbe286d8_26,RIbe28570_23,RIbe28e58_42,RIbe28de0_41,RIbe28840_29,RIbe28750_27,
        RIbe29920_65,RIbe27b98_2,RIbe284f8_22,RIbe28318_18,RIbe28048_12,RIbe27d00_5,RIbe29a88_68,RIbe27c10_3,RIbe290b0_47,RIbe28c78_38,
        RIbe28c00_37,RIbe29308_52,RIbe293f8_54,RIbe29038_46,RIbe28fc0_45,RIbe29650_59,RIbe288b8_30,RIbe28a98_34,RIbe296c8_60,RIbe29830_63,
        RIbe291a0_49,RIbe295d8_58,RIbe29740_61,RIbe282a0_17,RIbe28138_14,RIbe29470_55,RIbe297b8_62,RIbe294e8_56,RIbe280c0_13,RIbe28228_16,
        RIbe281b0_15,RIbe29290_51,RIbe28930_31,RIbe29560_57,RIbe28a20_33,RIbe289a8_32,RIbe29b00_69,RIbe29128_48,RIbe28b88_36,RIbe28b10_35,
        RIbe29218_50,RIbe29a10_67,RIbe28408_20,RIbe28390_19,RIbe28480_21,RIbe27c88_4,RIbe27df0_7,RIbe287c8_28,RIbe28d68_40,RIbe29998_66,
        RIbe285e8_24,RIbe28660_25,RIbe27e68_8,RIbe298a8_64,RIbe28cf0_39,RIbe27f58_10,RIbe27b20_1,RIbe29b78_70,RIbe27fd0_11,RIbe28ed0_43,
        RIbe29ce0_73,RIbe29d58_74,RIbe28f48_44,RIbe2a2f8_86,RIbe29bf0_71,RIbe29dd0_75,RIbe29c68_72,RIbe29fb0_79,RIbe29e48_76,RIbe29f38_78,
        RIbe29ec0_77,RIbe2aa00_101,RIbe2a898_98,RIbe2aa78_102,RIbe2b6a8_128,RIbe2b5b8_126,RIbe2a3e8_88,RIbe2a370_87,RIbe2acd0_107,RIbe2a028_80,
        RIbe2a118_82,RIbe2a0a0_81,RIbe2b360_121,RIbe2a820_97,RIbe2b2e8_120,RIbe2a4d8_90,RIbe2a910_99,RIbe2a988_100,RIbe2a550_91,RIbe2a460_89,
        RIbe2adc0_109,RIbe2a5c8_92,RIbe2ad48_108,RIbe2b540_125,RIbe2a190_83,RIbe2a640_93,RIbe2ac58_106,RIbe2a6b8_94,RIbe2abe0_105,RIbe2a7a8_96,
        RIbe2b4c8_124,RIbe2b450_123,RIbe2b3d8_122,RIbe2aeb0_111,RIbe2ae38_110,RIbe2a730_95,RIbe2a208_84,RIbe2b180_117,RIbe2b270_119,RIbe2af28_112,
        RIbe2b1f8_118,RIbe2b018_114,RIbe2afa0_113,RIbe2a280_85,RIbe2b108_116,RIbe2b090_115,RIbe2ab68_104,RIbe2aaf0_103,RIbe2b630_127,R_81_9fc6f08,
        R_82_9fc5ea0,R_83_90f04e0,R_84_90effa0,R_85_90e8ad0,R_86_90e3e08,R_87_90f1a88,R_88_90e8638,R_89_90f1200,R_8a_90f12a8,R_8b_90f0cc0,
        R_8c_90ef088,R_8d_90f1158,R_8e_90e49d8,R_8f_90e3eb0,R_90_9fc69c8,R_91_90e9c88,R_92_90f0588,R_93_90eacf0,R_94_90ebb60,R_95_90e66b8,
        R_96_9fc6d10,R_97_90ead98,R_98_90e90b8,R_99_90eb038,R_9a_90e9d30,R_9b_90e7bb8,R_9c_9fc7b80,R_9d_90ebd58,R_9e_90e9a90,R_9f_90efb08,
        R_a0_90e6e98,R_a1_90f0780,R_a2_90e2da0,R_a3_90f0240,R_a4_9fc7ad8,R_a5_9fc73a0,R_a6_9fc6680,R_a7_90e4f18,R_a8_90e3388,R_a9_9fc67d0,
        R_aa_90f17e8,R_ab_90e4888,R_ac_90e9010,R_ad_90eee90,R_ae_90e53b0,R_af_90ebc08,R_b0_90e8440,R_b1_90ea900,R_b2_90e9400,R_b3_9fc6bc0,
        R_b4_90e4690,R_b5_90e3778,R_b6_90e9160,R_b7_90e29b0,R_b8_90e2278,R_b9_9fc6a70,R_ba_90ebf50,R_bb_90f0e10,R_bc_9fc7640,R_bd_90f1dd0,
        R_be_90f0630,R_bf_90f0eb8,R_c0_90e34d8,R_c1_90e9f28,R_c2_90f0d68,R_c3_90ea7b0,R_c4_9fc7448,R_c5_90eb428,R_c6_90e81a0,R_c7_90f0a20,
        R_c8_90efda8,R_c9_90e2c50,R_ca_90e88d8,R_cb_9fc6530,R_cc_90f06d8,R_cd_90efa60,R_ce_90e2b00,R_cf_9fc6920,R_d0_90f1f20,R_d1_90e7678,
        R_d2_90efd00,R_d3_90e7e58,R_d4_90e7d08,R_d5_90eaa50,R_d6_90e3040,R_d7_90efe50,R_d8_90f1350,R_d9_9fc71a8,R_da_9fc9cf8,R_db_90ef9b8,
        R_dc_90e4540,R_dd_90f0ac8,R_de_90e30e8,R_df_9fc6290,R_e0_9fc78e0,R_e1_90e5500,R_e2_90e68b0,R_e3_90eede8,R_e4_90e64c0,R_e5_9fc7100,
        R_e6_90e2470,R_e7_90ebea8,R_e8_90e4a80,R_e9_90ef910,R_ea_9fc7c28,R_eb_90eb4d0,R_ec_90f14a0,R_ed_90ef5c8,R_ee_90e4498,R_ef_90e4000,
        R_f0_90f0048,R_f1_90ea3c0,R_f2_90f1e78,R_f3_90f00f0);
input RIbe29380_53,RIbe27d78_6,RIbe27ee0_9,RIbe286d8_26,RIbe28570_23,RIbe28e58_42,RIbe28de0_41,RIbe28840_29,RIbe28750_27,
        RIbe29920_65,RIbe27b98_2,RIbe284f8_22,RIbe28318_18,RIbe28048_12,RIbe27d00_5,RIbe29a88_68,RIbe27c10_3,RIbe290b0_47,RIbe28c78_38,
        RIbe28c00_37,RIbe29308_52,RIbe293f8_54,RIbe29038_46,RIbe28fc0_45,RIbe29650_59,RIbe288b8_30,RIbe28a98_34,RIbe296c8_60,RIbe29830_63,
        RIbe291a0_49,RIbe295d8_58,RIbe29740_61,RIbe282a0_17,RIbe28138_14,RIbe29470_55,RIbe297b8_62,RIbe294e8_56,RIbe280c0_13,RIbe28228_16,
        RIbe281b0_15,RIbe29290_51,RIbe28930_31,RIbe29560_57,RIbe28a20_33,RIbe289a8_32,RIbe29b00_69,RIbe29128_48,RIbe28b88_36,RIbe28b10_35,
        RIbe29218_50,RIbe29a10_67,RIbe28408_20,RIbe28390_19,RIbe28480_21,RIbe27c88_4,RIbe27df0_7,RIbe287c8_28,RIbe28d68_40,RIbe29998_66,
        RIbe285e8_24,RIbe28660_25,RIbe27e68_8,RIbe298a8_64,RIbe28cf0_39,RIbe27f58_10,RIbe27b20_1,RIbe29b78_70,RIbe27fd0_11,RIbe28ed0_43,
        RIbe29ce0_73,RIbe29d58_74,RIbe28f48_44,RIbe2a2f8_86,RIbe29bf0_71,RIbe29dd0_75,RIbe29c68_72,RIbe29fb0_79,RIbe29e48_76,RIbe29f38_78,
        RIbe29ec0_77,RIbe2aa00_101,RIbe2a898_98,RIbe2aa78_102,RIbe2b6a8_128,RIbe2b5b8_126,RIbe2a3e8_88,RIbe2a370_87,RIbe2acd0_107,RIbe2a028_80,
        RIbe2a118_82,RIbe2a0a0_81,RIbe2b360_121,RIbe2a820_97,RIbe2b2e8_120,RIbe2a4d8_90,RIbe2a910_99,RIbe2a988_100,RIbe2a550_91,RIbe2a460_89,
        RIbe2adc0_109,RIbe2a5c8_92,RIbe2ad48_108,RIbe2b540_125,RIbe2a190_83,RIbe2a640_93,RIbe2ac58_106,RIbe2a6b8_94,RIbe2abe0_105,RIbe2a7a8_96,
        RIbe2b4c8_124,RIbe2b450_123,RIbe2b3d8_122,RIbe2aeb0_111,RIbe2ae38_110,RIbe2a730_95,RIbe2a208_84,RIbe2b180_117,RIbe2b270_119,RIbe2af28_112,
        RIbe2b1f8_118,RIbe2b018_114,RIbe2afa0_113,RIbe2a280_85,RIbe2b108_116,RIbe2b090_115,RIbe2ab68_104,RIbe2aaf0_103,RIbe2b630_127;
output R_81_9fc6f08,R_82_9fc5ea0,R_83_90f04e0,R_84_90effa0,R_85_90e8ad0,R_86_90e3e08,R_87_90f1a88,R_88_90e8638,R_89_90f1200,
        R_8a_90f12a8,R_8b_90f0cc0,R_8c_90ef088,R_8d_90f1158,R_8e_90e49d8,R_8f_90e3eb0,R_90_9fc69c8,R_91_90e9c88,R_92_90f0588,R_93_90eacf0,
        R_94_90ebb60,R_95_90e66b8,R_96_9fc6d10,R_97_90ead98,R_98_90e90b8,R_99_90eb038,R_9a_90e9d30,R_9b_90e7bb8,R_9c_9fc7b80,R_9d_90ebd58,
        R_9e_90e9a90,R_9f_90efb08,R_a0_90e6e98,R_a1_90f0780,R_a2_90e2da0,R_a3_90f0240,R_a4_9fc7ad8,R_a5_9fc73a0,R_a6_9fc6680,R_a7_90e4f18,
        R_a8_90e3388,R_a9_9fc67d0,R_aa_90f17e8,R_ab_90e4888,R_ac_90e9010,R_ad_90eee90,R_ae_90e53b0,R_af_90ebc08,R_b0_90e8440,R_b1_90ea900,
        R_b2_90e9400,R_b3_9fc6bc0,R_b4_90e4690,R_b5_90e3778,R_b6_90e9160,R_b7_90e29b0,R_b8_90e2278,R_b9_9fc6a70,R_ba_90ebf50,R_bb_90f0e10,
        R_bc_9fc7640,R_bd_90f1dd0,R_be_90f0630,R_bf_90f0eb8,R_c0_90e34d8,R_c1_90e9f28,R_c2_90f0d68,R_c3_90ea7b0,R_c4_9fc7448,R_c5_90eb428,
        R_c6_90e81a0,R_c7_90f0a20,R_c8_90efda8,R_c9_90e2c50,R_ca_90e88d8,R_cb_9fc6530,R_cc_90f06d8,R_cd_90efa60,R_ce_90e2b00,R_cf_9fc6920,
        R_d0_90f1f20,R_d1_90e7678,R_d2_90efd00,R_d3_90e7e58,R_d4_90e7d08,R_d5_90eaa50,R_d6_90e3040,R_d7_90efe50,R_d8_90f1350,R_d9_9fc71a8,
        R_da_9fc9cf8,R_db_90ef9b8,R_dc_90e4540,R_dd_90f0ac8,R_de_90e30e8,R_df_9fc6290,R_e0_9fc78e0,R_e1_90e5500,R_e2_90e68b0,R_e3_90eede8,
        R_e4_90e64c0,R_e5_9fc7100,R_e6_90e2470,R_e7_90ebea8,R_e8_90e4a80,R_e9_90ef910,R_ea_9fc7c28,R_eb_90eb4d0,R_ec_90f14a0,R_ed_90ef5c8,
        R_ee_90e4498,R_ef_90e4000,R_f0_90f0048,R_f1_90ea3c0,R_f2_90f1e78,R_f3_90f00f0;

wire \244 , \245 , \246_N$2 , \247_N$4 , \248_ZERO , \249 , \250 , \251_N$1 , \252_N$3 ,
         \253_ONE , \254 , \255 , \256 , \257 , \258 , \259 , \260 , \261 , \262 ,
         \263 , \264 , \265 , \266 , \267 , \268 , \269 , \270 , \271 , \272 ,
         \273 , \274 , \275 , \276 , \277 , \278 , \279 , \280 , \281 , \282 ,
         \283 , \284 , \285 , \286 , \287 , \288 , \289 , \290 , \291 , \292 ,
         \293 , \294 , \295 , \296 , \297 , \298 , \299 , \300 , \301 , \302 ,
         \303 , \304 , \305 , \306 , \307 , \308 , \309 , \310 , \311 , \312 ,
         \313 , \314 , \315 , \316 , \317 , \318 , \319 , \320 , \321 , \322 ,
         \323 , \324 , \325 , \326 , \327 , \328 , \329 , \330 , \331 , \332 ,
         \333 , \334 , \335 , \336 , \337 , \338 , \339 , \340 , \341 , \342 ,
         \343 , \344 , \345 , \346 , \347 , \348 , \349 , \350 , \351 , \352 ,
         \353 , \354 , \355 , \356 , \357 , \358 , \359 , \360 , \361 , \362 ,
         \363 , \364 , \365 , \366 , \367 , \368 , \369 , \370 , \371 , \372 ,
         \373 , \374 , \375 , \376 , \377 , \378 , \379 , \380 , \381 , \382 ,
         \383 , \384 , \385 , \386 , \387 , \388 , \389 , \390 , \391 , \392 ,
         \393 , \394 , \395 , \396 , \397 , \398 , \399 , \400 , \401 , \402 ,
         \403 , \404 , \405 , \406 , \407 , \408 , \409 , \410 , \411 , \412 ,
         \413 , \414 , \415 , \416 , \417 , \418 , \419 , \420 , \421 , \422 ,
         \423 , \424 , \425 , \426 , \427 , \428 , \429 , \430 , \431 , \432 ,
         \433 , \434 , \435 , \436 , \437 , \438 , \439 , \440 , \441 , \442 ,
         \443 , \444 , \445 , \446 , \447 , \448 , \449 , \450 , \451 , \452 ,
         \453 , \454 , \455 , \456 , \457 , \458 , \459 , \460 , \461 , \462 ,
         \463 , \464 , \465 , \466 , \467 , \468 , \469 , \470 , \471 , \472 ,
         \473 , \474 , \475 , \476 , \477 , \478 , \479 , \480 , \481 , \482 ,
         \483 , \484 , \485 , \486 , \487 , \488 , \489 , \490 , \491 , \492 ,
         \493 , \494 , \495 , \496 , \497 , \498 , \499 , \500 , \501 , \502 ,
         \503 , \504 , \505 , \506 , \507 , \508 , \509 , \510 , \511 , \512 ,
         \513 , \514 , \515 , \516 , \517 , \518 , \519 , \520 , \521 , \522 ,
         \523 , \524 , \525 , \526 , \527 , \528 , \529 , \530 , \531 , \532 ,
         \533 , \534 , \535 , \536 , \537 , \538 , \539 , \540 , \541 , \542 ,
         \543 , \544 , \545 , \546 , \547 , \548 , \549 , \550 , \551 , \552 ,
         \553 , \554 , \555 , \556 , \557 , \558 , \559 , \560 , \561 , \562 ,
         \563 , \564 , \565 , \566 , \567 , \568 , \569 , \570 , \571 , \572 ,
         \573 , \574 , \575 , \576 , \577 , \578 , \579 , \580 , \581 , \582 ,
         \583 , \584 , \585 , \586 , \587 , \588 , \589 , \590 , \591 , \592 ,
         \593 , \594 , \595 , \596 , \597 , \598 , \599 , \600 , \601 , \602 ,
         \603 , \604 , \605 , \606 , \607 , \608 , \609 , \610 , \611 , \612 ,
         \613 , \614 , \615 , \616 , \617 , \618 , \619 , \620 , \621 , \622 ,
         \623 , \624 , \625 , \626 , \627 , \628 , \629 , \630 , \631 , \632 ,
         \633 , \634 , \635 , \636 , \637 , \638 , \639 , \640 , \641 , \642 ,
         \643 , \644 , \645 , \646 , \647 , \648 , \649 , \650 , \651 , \652 ,
         \653 , \654 , \655 , \656 , \657 , \658 , \659 , \660 , \661 , \662 ,
         \663 , \664 , \665 , \666 , \667 , \668 , \669 , \670 , \671 , \672 ,
         \673 , \674 , \675 , \676 , \677 , \678 , \679 , \680 , \681 , \682 ,
         \683 , \684 , \685 , \686 , \687 , \688 , \689 , \690 , \691 , \692 ,
         \693 , \694 , \695 , \696 , \697 , \698 , \699 , \700 , \701 , \702 ,
         \703 , \704 , \705 , \706 , \707 , \708 , \709 , \710 , \711 , \712 ,
         \713 , \714 , \715 , \716 , \717 , \718 , \719 , \720 , \721 , \722 ,
         \723 , \724 , \725 , \726 , \727 , \728 , \729 , \730 , \731 , \732 ,
         \733 , \734 , \735 , \736 , \737 , \738 , \739 , \740 , \741 , \742 ,
         \743 , \744 , \745 , \746 , \747 , \748 , \749 , \750 , \751 , \752 ,
         \753 , \754 , \755 , \756 , \757 , \758 , \759 , \760 , \761 , \762 ,
         \763 , \764 , \765 , \766 , \767 , \768 , \769 , \770 , \771 , \772 ,
         \773 , \774 , \775 , \776 , \777 , \778 , \779 , \780 , \781 , \782 ,
         \783 , \784 , \785 , \786 , \787 , \788 , \789 , \790 , \791 , \792 ,
         \793 , \794 , \795 , \796 , \797 , \798 , \799 , \800 , \801 , \802 ,
         \803 , \804 , \805 , \806 , \807 , \808 , \809 , \810 , \811 , \812 ,
         \813 , \814 , \815 , \816 , \817 , \818 , \819 , \820 , \821 , \822 ,
         \823 , \824 , \825 , \826 , \827 , \828 , \829 , \830 , \831 , \832 ,
         \833 , \834 , \835 , \836 , \837 , \838 , \839 , \840 , \841 , \842 ,
         \843 , \844 , \845 , \846 , \847 , \848 , \849 , \850 , \851 , \852 ,
         \853 , \854 , \855 , \856 , \857 , \858 , \859 , \860 , \861 , \862 ,
         \863 , \864 , \865 , \866 , \867 , \868 , \869 , \870 , \871 , \872 ,
         \873 , \874 , \875 , \876 , \877 , \878 , \879 , \880 , \881 , \882 ,
         \883 , \884 , \885 , \886 , \887 , \888 , \889 , \890 , \891 , \892 ,
         \893 , \894 , \895 , \896 , \897 , \898 , \899 , \900 , \901 , \902 ,
         \903 , \904 , \905 , \906 , \907 , \908 , \909 , \910 , \911 , \912 ,
         \913 , \914 , \915 , \916 , \917 , \918 , \919 , \920 , \921 , \922 ,
         \923 , \924 , \925 , \926 , \927 , \928 , \929 , \930 , \931 , \932 ,
         \933 , \934 , \935 , \936 , \937 , \938 , \939 , \940 , \941 , \942 ,
         \943 , \944 , \945 , \946 , \947 , \948 , \949 , \950 , \951 , \952 ,
         \953 , \954 , \955 , \956 , \957 , \958 , \959 , \960 , \961 , \962 ,
         \963 , \964 , \965 , \966 , \967 , \968 , \969 , \970 , \971 , \972 ,
         \973 , \974 , \975 , \976 , \977 , \978 , \979 , \980 , \981 , \982 ,
         \983 , \984 , \985 , \986 , \987 , \988 , \989 , \990 , \991 , \992 ,
         \993 , \994 , \995 , \996 , \997 , \998 , \999 , \1000 , \1001 , \1002 ,
         \1003 , \1004 , \1005 , \1006 , \1007 , \1008 , \1009 , \1010 , \1011 , \1012 ,
         \1013 , \1014 , \1015 , \1016 , \1017 , \1018 , \1019 , \1020 , \1021 , \1022 ,
         \1023 , \1024 , \1025 , \1026 , \1027 , \1028 , \1029 , \1030 , \1031 , \1032 ,
         \1033 , \1034 , \1035 , \1036 , \1037 , \1038 , \1039 , \1040 , \1041 , \1042 ,
         \1043 , \1044 , \1045 , \1046 , \1047 , \1048 , \1049 , \1050 , \1051 , \1052 ,
         \1053 , \1054 , \1055 , \1056 , \1057 , \1058 , \1059 , \1060 , \1061 , \1062 ,
         \1063 , \1064 , \1065 , \1066 , \1067 , \1068 , \1069 , \1070 , \1071 , \1072 ,
         \1073 , \1074 , \1075 , \1076 , \1077 , \1078 , \1079 , \1080 , \1081 , \1082 ,
         \1083 , \1084 , \1085 , \1086 , \1087 , \1088 , \1089 , \1090 , \1091 , \1092 ,
         \1093 , \1094 , \1095 , \1096 , \1097 , \1098 , \1099 , \1100 , \1101 , \1102 ,
         \1103 , \1104 , \1105 , \1106 , \1107 , \1108 , \1109 , \1110 , \1111 , \1112 ,
         \1113 , \1114 , \1115 , \1116 , \1117 , \1118 , \1119 , \1120 , \1121 , \1122 ,
         \1123 , \1124 , \1125 , \1126 , \1127 , \1128 , \1129 , \1130 , \1131 , \1132 ,
         \1133 , \1134 , \1135 , \1136 , \1137 , \1138 , \1139 , \1140 , \1141 , \1142 ,
         \1143 , \1144 , \1145 , \1146 , \1147 , \1148 , \1149 , \1150 , \1151 , \1152 ,
         \1153 , \1154 , \1155 , \1156 , \1157 , \1158 , \1159 , \1160 , \1161 , \1162 ,
         \1163 , \1164 , \1165 , \1166 , \1167 , \1168 , \1169 , \1170 , \1171 , \1172 ,
         \1173 , \1174 , \1175 , \1176 , \1177 , \1178 , \1179 , \1180 , \1181 , \1182 ,
         \1183 , \1184 , \1185 , \1186 , \1187 , \1188 , \1189 , \1190 , \1191 , \1192 ,
         \1193 , \1194 , \1195 , \1196 , \1197 , \1198 , \1199 , \1200 , \1201 , \1202 ,
         \1203 , \1204 , \1205 , \1206 , \1207 , \1208 , \1209 , \1210 , \1211 , \1212 ,
         \1213 , \1214 , \1215 , \1216 , \1217 , \1218 , \1219 , \1220 , \1221 , \1222 ,
         \1223 , \1224 , \1225 , \1226 , \1227 , \1228 , \1229 , \1230 , \1231 , \1232 ,
         \1233 , \1234 , \1235 , \1236 , \1237 , \1238 , \1239 , \1240 , \1241 , \1242 ,
         \1243 , \1244 , \1245 , \1246 , \1247 , \1248 , \1249 , \1250 , \1251 , \1252 ,
         \1253 , \1254 , \1255 , \1256 , \1257 , \1258 , \1259 , \1260 , \1261 , \1262 ,
         \1263 , \1264 , \1265 , \1266 , \1267 , \1268 , \1269 , \1270 , \1271 , \1272 ,
         \1273 , \1274 , \1275 , \1276 , \1277 , \1278 , \1279 , \1280 , \1281 , \1282 ,
         \1283 , \1284 , \1285 , \1286 , \1287 , \1288 , \1289 , \1290 , \1291 , \1292 ,
         \1293 , \1294 , \1295 , \1296 , \1297 , \1298 , \1299 , \1300 , \1301 , \1302 ,
         \1303 , \1304 , \1305 , \1306 , \1307 , \1308 , \1309 , \1310 , \1311 , \1312 ,
         \1313 , \1314 , \1315 , \1316 , \1317 , \1318 , \1319 , \1320 , \1321 , \1322 ,
         \1323 , \1324 , \1325 , \1326 , \1327 , \1328 , \1329 , \1330 , \1331 , \1332 ,
         \1333 , \1334 , \1335 , \1336 , \1337 , \1338 , \1339 , \1340 , \1341 , \1342 ,
         \1343 , \1344 , \1345 , \1346 , \1347 , \1348 , \1349 , \1350 , \1351 , \1352 ,
         \1353 , \1354 , \1355 , \1356 , \1357 , \1358 , \1359 , \1360 , \1361 , \1362 ,
         \1363 , \1364 , \1365 , \1366 , \1367 , \1368 , \1369 , \1370 , \1371 , \1372 ,
         \1373 , \1374 , \1375 , \1376 , \1377 , \1378 , \1379 , \1380 , \1381 , \1382 ,
         \1383 , \1384 , \1385 , \1386 , \1387 , \1388 , \1389 , \1390 , \1391 , \1392 ,
         \1393 , \1394 , \1395 , \1396 , \1397 , \1398 , \1399 , \1400 , \1401 , \1402 ,
         \1403 , \1404 , \1405 , \1406 , \1407 , \1408 , \1409 , \1410 , \1411 , \1412 ,
         \1413 , \1414 , \1415 , \1416 , \1417 , \1418 , \1419 , \1420 , \1421 , \1422 ,
         \1423 , \1424 , \1425 , \1426 , \1427 , \1428 , \1429 , \1430 , \1431 , \1432 ,
         \1433 , \1434 , \1435 , \1436 , \1437 , \1438 , \1439 , \1440 , \1441 , \1442 ,
         \1443 , \1444 , \1445 , \1446 , \1447 , \1448 , \1449 , \1450 , \1451 , \1452 ,
         \1453 , \1454 , \1455 , \1456 , \1457 , \1458 , \1459 , \1460 , \1461 , \1462 ,
         \1463 , \1464 , \1465 , \1466 , \1467 , \1468 , \1469 , \1470 , \1471 , \1472 ,
         \1473 , \1474 , \1475 , \1476 , \1477 , \1478 , \1479 , \1480 , \1481 , \1482 ,
         \1483 , \1484 , \1485 , \1486 , \1487 , \1488 , \1489 , \1490 , \1491 , \1492 ,
         \1493 , \1494 , \1495 , \1496 , \1497 , \1498 , \1499 , \1500 , \1501 , \1502 ,
         \1503 , \1504 , \1505 , \1506 , \1507 , \1508 , \1509 , \1510 , \1511 , \1512 ,
         \1513 , \1514 , \1515 , \1516 , \1517 , \1518 , \1519 , \1520 , \1521 , \1522 ,
         \1523 , \1524 , \1525 , \1526 , \1527 , \1528 , \1529 , \1530 , \1531 , \1532 ,
         \1533 , \1534 , \1535 , \1536 , \1537 , \1538 , \1539 , \1540 , \1541 , \1542 ,
         \1543 , \1544 , \1545 , \1546 , \1547 , \1548 , \1549 , \1550 , \1551 , \1552 ,
         \1553 , \1554 , \1555 , \1556 , \1557 , \1558 , \1559 , \1560 , \1561 , \1562 ,
         \1563 , \1564 , \1565 , \1566 , \1567 , \1568 , \1569 , \1570 , \1571 , \1572 ,
         \1573 , \1574 , \1575 , \1576 , \1577 , \1578 , \1579 , \1580 , \1581 , \1582 ,
         \1583 , \1584 , \1585 , \1586 , \1587 , \1588 , \1589 , \1590 , \1591 , \1592 ,
         \1593 , \1594 , \1595 , \1596 , \1597 , \1598 , \1599 , \1600 , \1601 , \1602 ,
         \1603 , \1604 , \1605 , \1606 , \1607 , \1608 , \1609 , \1610 , \1611 , \1612 ,
         \1613 , \1614 , \1615 , \1616 , \1617 , \1618 , \1619 , \1620 , \1621 , \1622 ,
         \1623 , \1624 , \1625 , \1626 , \1627 , \1628 , \1629 , \1630 , \1631 , \1632 ,
         \1633 , \1634 , \1635 , \1636 , \1637 , \1638 , \1639 , \1640 , \1641 , \1642 ,
         \1643 , \1644 , \1645 , \1646 , \1647 , \1648 , \1649 , \1650 , \1651 , \1652 ,
         \1653 , \1654 , \1655 , \1656 , \1657 , \1658 , \1659 , \1660 , \1661 , \1662 ,
         \1663 , \1664 , \1665 , \1666 , \1667 , \1668 , \1669 , \1670 , \1671 , \1672 ,
         \1673 , \1674 , \1675 , \1676 , \1677 , \1678 , \1679 , \1680 , \1681 , \1682 ,
         \1683 , \1684 , \1685 , \1686 , \1687 , \1688 , \1689 , \1690 , \1691 , \1692 ,
         \1693 , \1694 , \1695 , \1696 , \1697 , \1698 , \1699 , \1700 , \1701 , \1702 ,
         \1703 , \1704 , \1705 , \1706 , \1707 , \1708 , \1709 , \1710 , \1711 , \1712 ,
         \1713 , \1714 , \1715 , \1716 , \1717 , \1718 , \1719 , \1720 , \1721 , \1722 ,
         \1723 , \1724 , \1725 , \1726 , \1727 , \1728 , \1729 , \1730 , \1731 , \1732 ,
         \1733 , \1734 , \1735 , \1736 , \1737 , \1738 , \1739 , \1740 , \1741 , \1742 ,
         \1743 , \1744 , \1745 , \1746 , \1747 , \1748 , \1749 , \1750 , \1751 , \1752 ,
         \1753 , \1754 , \1755 , \1756 , \1757 , \1758 , \1759 , \1760 , \1761 , \1762 ,
         \1763 , \1764 , \1765 , \1766 , \1767 , \1768 , \1769 , \1770 , \1771 , \1772 ,
         \1773 , \1774 , \1775 , \1776 , \1777 , \1778 , \1779 , \1780 , \1781 , \1782 ,
         \1783 , \1784 , \1785 , \1786 , \1787 , \1788 , \1789 , \1790 , \1791 , \1792 ,
         \1793 , \1794 , \1795 , \1796 , \1797 , \1798 , \1799 , \1800 , \1801 , \1802 ,
         \1803 , \1804 , \1805 , \1806 , \1807 , \1808 , \1809 , \1810 , \1811 , \1812 ,
         \1813 , \1814 , \1815 , \1816 , \1817 , \1818 , \1819 , \1820 , \1821 , \1822 ,
         \1823 , \1824 , \1825 , \1826 , \1827 , \1828 , \1829 , \1830 , \1831 , \1832 ,
         \1833 , \1834 , \1835 , \1836 , \1837 , \1838 , \1839 , \1840 , \1841 , \1842 ,
         \1843 , \1844 , \1845 , \1846 , \1847 , \1848 , \1849 , \1850 , \1851 , \1852 ,
         \1853 , \1854 , \1855 , \1856 , \1857 , \1858 , \1859 , \1860 , \1861 , \1862 ,
         \1863 , \1864 , \1865 , \1866 , \1867 , \1868 , \1869 , \1870 , \1871 , \1872 ,
         \1873 , \1874 , \1875 , \1876 , \1877 , \1878 , \1879 , \1880 , \1881 , \1882 ,
         \1883 , \1884 , \1885 , \1886 , \1887 , \1888 , \1889 , \1890 , \1891 , \1892 ,
         \1893 , \1894 , \1895 , \1896 , \1897 , \1898 , \1899 , \1900 , \1901 , \1902 ,
         \1903 , \1904 , \1905 , \1906 , \1907 , \1908 , \1909 , \1910 , \1911 , \1912 ,
         \1913 , \1914 , \1915 , \1916 , \1917 , \1918 , \1919 , \1920 , \1921 , \1922 ,
         \1923 , \1924 , \1925 , \1926 , \1927 , \1928 , \1929 , \1930 , \1931 , \1932 ,
         \1933 , \1934 , \1935 , \1936 , \1937 , \1938 , \1939 , \1940 , \1941 , \1942 ,
         \1943 , \1944 , \1945 , \1946 , \1947 , \1948 , \1949 , \1950 , \1951 , \1952 ,
         \1953 , \1954 , \1955 , \1956 , \1957 , \1958 , \1959 , \1960 , \1961 , \1962 ,
         \1963 , \1964 , \1965 , \1966 , \1967 , \1968 , \1969 , \1970 , \1971 , \1972 ,
         \1973 , \1974 , \1975 , \1976 , \1977 , \1978 , \1979 , \1980 , \1981 , \1982 ,
         \1983 , \1984 , \1985 , \1986 , \1987 , \1988 , \1989 , \1990 , \1991 , \1992 ,
         \1993 , \1994 , \1995 , \1996 , \1997 , \1998 , \1999 , \2000 , \2001 , \2002 ,
         \2003 , \2004 , \2005 , \2006 , \2007 , \2008 , \2009 , \2010 , \2011 , \2012 ,
         \2013 , \2014 , \2015 , \2016 , \2017 , \2018 , \2019 , \2020 , \2021 , \2022 ,
         \2023 , \2024 , \2025 , \2026 , \2027 , \2028 , \2029 , \2030 , \2031 , \2032 ,
         \2033 , \2034 , \2035 , \2036 , \2037 , \2038 , \2039 , \2040 , \2041 , \2042 ,
         \2043 , \2044 , \2045 , \2046 , \2047 , \2048 , \2049 , \2050 , \2051 , \2052 ,
         \2053 , \2054 , \2055 , \2056 , \2057 , \2058 , \2059 , \2060 , \2061 , \2062 ,
         \2063 , \2064 , \2065 , \2066 , \2067 , \2068 , \2069 , \2070 , \2071 , \2072 ,
         \2073 , \2074 , \2075 , \2076 , \2077 , \2078 , \2079 , \2080 , \2081 , \2082 ,
         \2083 , \2084 , \2085 , \2086 , \2087 , \2088 , \2089 , \2090 , \2091 , \2092 ,
         \2093 , \2094 , \2095 , \2096 , \2097 , \2098 , \2099 , \2100 , \2101 , \2102 ,
         \2103 , \2104 , \2105 , \2106 , \2107 , \2108 , \2109 , \2110 , \2111 , \2112 ,
         \2113 , \2114 , \2115 , \2116 , \2117 , \2118 , \2119 , \2120 , \2121 , \2122 ,
         \2123 , \2124 , \2125 , \2126 , \2127 , \2128 , \2129 , \2130 , \2131 , \2132 ,
         \2133 , \2134 , \2135 , \2136 , \2137 , \2138 , \2139 , \2140 , \2141 , \2142 ,
         \2143 , \2144 , \2145 , \2146 , \2147 , \2148 , \2149 , \2150 , \2151 , \2152 ,
         \2153 , \2154 , \2155 , \2156 , \2157 , \2158 , \2159 , \2160 , \2161 , \2162 ,
         \2163 , \2164 , \2165 , \2166 , \2167 , \2168 , \2169 , \2170 , \2171 , \2172 ,
         \2173 , \2174 , \2175 , \2176 , \2177 , \2178 , \2179 , \2180 , \2181 , \2182 ,
         \2183 , \2184 , \2185 , \2186 , \2187 , \2188 , \2189 , \2190 , \2191 , \2192 ,
         \2193 , \2194 , \2195 , \2196 , \2197 , \2198 , \2199 , \2200 , \2201 , \2202 ,
         \2203 , \2204 , \2205 , \2206 , \2207 , \2208 , \2209 , \2210 , \2211 , \2212 ,
         \2213 , \2214 , \2215 , \2216 , \2217 , \2218 , \2219 , \2220 , \2221 , \2222 ,
         \2223 , \2224 , \2225 , \2226 , \2227 , \2228 , \2229 , \2230 , \2231 , \2232 ,
         \2233 , \2234 , \2235 , \2236 , \2237 , \2238 , \2239 , \2240 , \2241 , \2242 ,
         \2243 , \2244 , \2245 , \2246 , \2247 , \2248 , \2249 , \2250 , \2251 , \2252 ,
         \2253 , \2254 , \2255 , \2256 , \2257 , \2258 , \2259 , \2260 , \2261 , \2262 ,
         \2263 , \2264 , \2265 , \2266 , \2267 , \2268 , \2269 , \2270 , \2271 , \2272 ,
         \2273 , \2274 , \2275 , \2276 , \2277 , \2278 , \2279 , \2280 , \2281 , \2282 ,
         \2283 , \2284 , \2285 , \2286 , \2287 , \2288 , \2289 , \2290 , \2291 , \2292 ,
         \2293 , \2294 , \2295 , \2296 , \2297 , \2298 , \2299 , \2300 , \2301 , \2302 ,
         \2303 , \2304 , \2305 , \2306 , \2307 , \2308 , \2309 , \2310 , \2311 , \2312 ,
         \2313 , \2314 , \2315 , \2316 , \2317 , \2318 , \2319 , \2320 , \2321 , \2322 ,
         \2323 , \2324 , \2325 , \2326 , \2327 , \2328 , \2329 , \2330 , \2331 , \2332 ,
         \2333 , \2334 , \2335 , \2336 , \2337 , \2338 , \2339 , \2340 , \2341 , \2342 ,
         \2343 , \2344 , \2345 , \2346 , \2347 , \2348 , \2349 , \2350 , \2351 , \2352 ,
         \2353 , \2354 , \2355 , \2356 , \2357 , \2358 , \2359 , \2360 , \2361 , \2362 ,
         \2363 , \2364 , \2365 , \2366 , \2367 , \2368 , \2369 , \2370 , \2371 , \2372 ,
         \2373 , \2374 , \2375 , \2376 , \2377 , \2378 , \2379 , \2380 , \2381 , \2382 ,
         \2383 , \2384 , \2385 , \2386 , \2387 , \2388 , \2389 , \2390 , \2391 , \2392 ,
         \2393 , \2394 , \2395 , \2396 , \2397 , \2398 , \2399 , \2400 , \2401 , \2402 ,
         \2403 , \2404 , \2405 , \2406 , \2407 , \2408 , \2409 , \2410 , \2411 , \2412 ,
         \2413 , \2414 , \2415 , \2416 , \2417 , \2418 , \2419 , \2420 , \2421 , \2422 ,
         \2423 , \2424 , \2425 , \2426 , \2427 , \2428 , \2429 , \2430 , \2431 , \2432 ,
         \2433 , \2434 , \2435 , \2436 , \2437 , \2438 , \2439 , \2440 , \2441 , \2442 ,
         \2443 , \2444 , \2445 , \2446 , \2447 , \2448 , \2449 , \2450 , \2451 , \2452 ,
         \2453 , \2454 , \2455 , \2456 , \2457 , \2458 , \2459 , \2460 , \2461 , \2462 ,
         \2463 , \2464 , \2465 , \2466 , \2467 , \2468 , \2469 , \2470 , \2471 , \2472 ,
         \2473 , \2474 , \2475 , \2476 , \2477 , \2478 , \2479 , \2480 , \2481 , \2482 ,
         \2483 , \2484 , \2485 , \2486 , \2487 , \2488 , \2489 , \2490 , \2491 , \2492 ,
         \2493 , \2494 , \2495 , \2496 , \2497 , \2498 , \2499 , \2500 , \2501 , \2502 ,
         \2503 , \2504 , \2505 , \2506 , \2507 , \2508 , \2509 , \2510 , \2511 , \2512 ,
         \2513 , \2514 , \2515 , \2516 , \2517 , \2518 , \2519 , \2520 , \2521 , \2522 ,
         \2523 , \2524 , \2525 , \2526 , \2527 , \2528 , \2529 , \2530 , \2531 , \2532 ,
         \2533 , \2534 , \2535 , \2536 , \2537 , \2538 , \2539 , \2540 , \2541 , \2542 ,
         \2543 , \2544 , \2545 , \2546 , \2547 , \2548 , \2549 , \2550 , \2551 , \2552 ,
         \2553 , \2554 , \2555 , \2556 , \2557 , \2558 , \2559 , \2560 , \2561 , \2562 ,
         \2563 , \2564 , \2565 , \2566 , \2567 , \2568 , \2569 , \2570 , \2571 , \2572 ,
         \2573 , \2574 , \2575 , \2576 , \2577 , \2578 , \2579 , \2580 , \2581 , \2582 ,
         \2583 , \2584 , \2585 , \2586 , \2587 , \2588 , \2589 , \2590 , \2591 , \2592 ,
         \2593 , \2594 , \2595 , \2596 , \2597 , \2598 , \2599 , \2600 , \2601 , \2602 ,
         \2603 , \2604 , \2605 , \2606 , \2607 , \2608 , \2609 , \2610 , \2611 , \2612 ,
         \2613 , \2614 , \2615 , \2616 , \2617 , \2618 , \2619 , \2620 , \2621 , \2622 ,
         \2623 , \2624 , \2625 , \2626 , \2627 , \2628 , \2629 , \2630 , \2631 , \2632 ,
         \2633 , \2634 , \2635 , \2636 , \2637 , \2638 , \2639 , \2640 , \2641 , \2642 ,
         \2643 , \2644 , \2645 , \2646 , \2647 , \2648 , \2649 , \2650 , \2651 , \2652 ,
         \2653 , \2654 , \2655 , \2656 , \2657 , \2658 , \2659 , \2660 , \2661 , \2662 ,
         \2663 , \2664 , \2665 , \2666 , \2667 , \2668 , \2669 , \2670 , \2671 , \2672 ,
         \2673 , \2674 , \2675 , \2676 , \2677 , \2678 , \2679 , \2680 , \2681 , \2682 ,
         \2683 , \2684 , \2685 , \2686 , \2687 , \2688 , \2689 , \2690 , \2691 , \2692 ,
         \2693 , \2694 , \2695 , \2696 , \2697 , \2698 , \2699 , \2700 , \2701 , \2702 ,
         \2703 , \2704 , \2705 , \2706 , \2707 , \2708 , \2709 , \2710 , \2711 , \2712 ,
         \2713 , \2714 , \2715 , \2716 , \2717 , \2718 , \2719 , \2720 , \2721 , \2722 ,
         \2723 , \2724 , \2725 , \2726 , \2727 , \2728 , \2729 , \2730 , \2731 , \2732 ,
         \2733 , \2734 , \2735 , \2736 , \2737 , \2738 , \2739 , \2740 , \2741 , \2742 ,
         \2743 , \2744 , \2745 , \2746 , \2747 , \2748 , \2749 , \2750 , \2751 , \2752 ,
         \2753 , \2754 , \2755 , \2756 , \2757 , \2758 , \2759 , \2760 , \2761 , \2762 ,
         \2763 , \2764 , \2765 , \2766 , \2767 , \2768 , \2769 , \2770 , \2771 , \2772 ,
         \2773 , \2774 , \2775 , \2776 , \2777 , \2778 , \2779 , \2780 , \2781 , \2782 ,
         \2783 , \2784 , \2785 , \2786 , \2787 , \2788 , \2789 , \2790 , \2791 , \2792 ,
         \2793 , \2794 , \2795 , \2796 , \2797 , \2798 , \2799 , \2800 , \2801 , \2802 ,
         \2803 , \2804 , \2805 , \2806 , \2807 , \2808 , \2809 , \2810 , \2811 , \2812 ,
         \2813 , \2814 , \2815 , \2816 , \2817 , \2818 , \2819 , \2820 , \2821 , \2822 ,
         \2823 , \2824 , \2825 , \2826 , \2827 , \2828 , \2829 , \2830 , \2831 , \2832 ,
         \2833 , \2834 , \2835 , \2836 , \2837 , \2838 , \2839 , \2840 , \2841 , \2842 ,
         \2843 , \2844 , \2845 , \2846 , \2847 , \2848 , \2849 , \2850 , \2851 , \2852 ,
         \2853 , \2854 , \2855 , \2856 , \2857 , \2858 , \2859 , \2860 , \2861 , \2862 ,
         \2863 , \2864 , \2865 , \2866 , \2867 , \2868 , \2869 , \2870 , \2871 , \2872 ,
         \2873 , \2874 , \2875 , \2876 , \2877 , \2878 , \2879 , \2880 , \2881 , \2882 ,
         \2883 , \2884 , \2885 , \2886 , \2887 , \2888 , \2889 , \2890 , \2891 , \2892 ,
         \2893 , \2894 , \2895 , \2896 , \2897 , \2898 , \2899 , \2900 , \2901 , \2902 ,
         \2903 , \2904 , \2905 , \2906 , \2907 , \2908 , \2909 , \2910 , \2911 , \2912 ,
         \2913 , \2914 , \2915 , \2916 , \2917 , \2918 , \2919 , \2920 , \2921 , \2922 ,
         \2923 , \2924 , \2925 , \2926 , \2927 , \2928 , \2929 , \2930 , \2931 , \2932 ,
         \2933 , \2934 , \2935 , \2936 , \2937 , \2938 , \2939 , \2940 , \2941 , \2942 ,
         \2943 , \2944 , \2945 , \2946 , \2947 , \2948 , \2949 , \2950 , \2951 , \2952 ,
         \2953 , \2954 , \2955 , \2956 , \2957 , \2958 , \2959 , \2960 , \2961 , \2962 ,
         \2963 , \2964 , \2965 , \2966 , \2967 , \2968 , \2969 , \2970 , \2971 , \2972 ,
         \2973 , \2974 , \2975 , \2976 , \2977 , \2978 , \2979 , \2980 , \2981 , \2982 ,
         \2983 , \2984 , \2985 , \2986 , \2987 , \2988 , \2989 , \2990 , \2991 , \2992 ,
         \2993 , \2994 , \2995 , \2996 , \2997 , \2998 , \2999 , \3000 , \3001 , \3002 ,
         \3003 , \3004 , \3005 , \3006 , \3007 , \3008 , \3009 , \3010 , \3011 , \3012 ,
         \3013 , \3014 , \3015 , \3016 , \3017 , \3018 , \3019 , \3020 , \3021 , \3022 ,
         \3023 , \3024 , \3025 , \3026 , \3027 , \3028 , \3029 , \3030 , \3031 , \3032 ,
         \3033 , \3034 , \3035 , \3036 , \3037 , \3038 , \3039 , \3040 , \3041 , \3042 ,
         \3043 , \3044 , \3045 , \3046 , \3047 , \3048 , \3049 , \3050 , \3051 , \3052 ,
         \3053 , \3054 , \3055 , \3056 , \3057 , \3058 , \3059 , \3060 , \3061 , \3062 ,
         \3063 , \3064 , \3065 , \3066 , \3067 , \3068 , \3069 , \3070 , \3071 , \3072 ,
         \3073 , \3074 , \3075 , \3076 , \3077 , \3078 , \3079 , \3080 , \3081 , \3082 ,
         \3083 , \3084 , \3085 , \3086 , \3087 , \3088 , \3089 , \3090 , \3091 , \3092 ,
         \3093 , \3094 , \3095 , \3096 , \3097 , \3098 , \3099 , \3100 , \3101 , \3102 ,
         \3103 , \3104 , \3105 , \3106 , \3107 , \3108 , \3109 , \3110 , \3111 , \3112 ,
         \3113 , \3114 , \3115 , \3116 , \3117 , \3118 , \3119 , \3120 , \3121 , \3122 ,
         \3123 , \3124 , \3125 , \3126 , \3127 , \3128 , \3129 , \3130 , \3131 , \3132 ,
         \3133 , \3134 , \3135 , \3136 , \3137 , \3138 , \3139 , \3140 , \3141 , \3142 ,
         \3143 , \3144 , \3145 , \3146 , \3147 , \3148 , \3149 , \3150 , \3151 , \3152 ,
         \3153 , \3154 , \3155 , \3156 , \3157 , \3158 , \3159 , \3160 , \3161 , \3162 ,
         \3163 , \3164 , \3165 , \3166 , \3167 , \3168 , \3169 , \3170 , \3171 , \3172 ,
         \3173 , \3174 , \3175 , \3176 , \3177 , \3178 , \3179 , \3180 , \3181 , \3182 ,
         \3183 , \3184 , \3185 , \3186 , \3187 , \3188 , \3189 , \3190 , \3191 , \3192 ,
         \3193 , \3194 , \3195 , \3196 , \3197 , \3198 , \3199 , \3200 , \3201 , \3202 ,
         \3203 , \3204 , \3205 , \3206 , \3207 , \3208 , \3209 , \3210 , \3211 , \3212 ,
         \3213 , \3214 , \3215 , \3216 , \3217 , \3218 , \3219 , \3220 , \3221 , \3222 ,
         \3223 , \3224 , \3225 , \3226 , \3227 , \3228 , \3229 , \3230 , \3231 , \3232 ,
         \3233 , \3234 , \3235 , \3236 , \3237 , \3238 , \3239 , \3240 , \3241 , \3242 ,
         \3243 , \3244 , \3245 , \3246 , \3247 , \3248 , \3249 , \3250 , \3251 , \3252 ,
         \3253 , \3254 , \3255 , \3256 , \3257 , \3258 , \3259 , \3260 , \3261 , \3262 ,
         \3263 , \3264 , \3265 , \3266 , \3267 , \3268 , \3269 , \3270 , \3271 , \3272 ,
         \3273 , \3274 , \3275 , \3276 , \3277 , \3278 , \3279 , \3280 , \3281 , \3282 ,
         \3283 , \3284 , \3285 , \3286 , \3287 , \3288 , \3289 , \3290 , \3291 , \3292 ,
         \3293 , \3294 , \3295 , \3296 , \3297 , \3298 , \3299 , \3300 , \3301 , \3302 ,
         \3303 , \3304 , \3305 , \3306 , \3307 , \3308 , \3309 , \3310 , \3311 , \3312 ,
         \3313 , \3314 , \3315 , \3316 , \3317 , \3318 , \3319 , \3320 , \3321 , \3322 ,
         \3323 , \3324 , \3325 , \3326 , \3327 , \3328 , \3329 , \3330 , \3331 , \3332 ,
         \3333 , \3334 , \3335 , \3336 , \3337 , \3338 , \3339 , \3340 , \3341 , \3342 ,
         \3343 , \3344 , \3345 , \3346 , \3347 , \3348 , \3349 , \3350 , \3351 , \3352 ,
         \3353 , \3354 , \3355 , \3356 , \3357 , \3358 , \3359 , \3360 , \3361 , \3362 ,
         \3363 , \3364 , \3365 , \3366 , \3367 , \3368 , \3369 , \3370 , \3371 , \3372 ,
         \3373 , \3374 , \3375 , \3376 , \3377 , \3378 , \3379 , \3380 , \3381 , \3382 ,
         \3383 , \3384 , \3385 , \3386 , \3387 , \3388 , \3389 , \3390 , \3391 , \3392 ,
         \3393 , \3394 , \3395 , \3396 , \3397 , \3398 , \3399 , \3400 , \3401 , \3402 ,
         \3403 , \3404 , \3405 , \3406 , \3407 , \3408 , \3409 , \3410 , \3411 , \3412 ,
         \3413 , \3414 , \3415 , \3416 , \3417 , \3418 , \3419 , \3420 , \3421 , \3422 ,
         \3423 , \3424 , \3425 , \3426 , \3427 , \3428 , \3429 , \3430 , \3431 , \3432 ,
         \3433 , \3434 , \3435 , \3436 , \3437 , \3438 , \3439 , \3440 , \3441 , \3442 ,
         \3443 , \3444 , \3445 , \3446 , \3447 , \3448 , \3449 , \3450 , \3451 , \3452 ,
         \3453 , \3454 , \3455 , \3456 , \3457 , \3458 , \3459 , \3460 , \3461 , \3462 ,
         \3463 , \3464 , \3465 , \3466 , \3467 , \3468 , \3469 , \3470 , \3471 , \3472 ,
         \3473 , \3474 , \3475 , \3476 , \3477 , \3478 , \3479 , \3480 , \3481 , \3482 ,
         \3483 , \3484 , \3485 , \3486 , \3487 , \3488 , \3489 , \3490 , \3491 , \3492 ,
         \3493 , \3494 , \3495 , \3496 , \3497 , \3498 , \3499 , \3500 , \3501 , \3502 ,
         \3503 , \3504 , \3505 , \3506 , \3507 , \3508 , \3509 , \3510 , \3511 , \3512 ,
         \3513 , \3514 , \3515 , \3516 , \3517 , \3518 , \3519 , \3520 , \3521 , \3522 ,
         \3523 , \3524 , \3525 , \3526 , \3527 , \3528 , \3529 , \3530 , \3531 , \3532 ,
         \3533 , \3534 , \3535 , \3536 , \3537 , \3538 , \3539 , \3540 , \3541 , \3542 ,
         \3543 , \3544 , \3545 , \3546 , \3547 , \3548 , \3549 , \3550 , \3551 , \3552 ,
         \3553 , \3554 , \3555 , \3556 , \3557 , \3558 , \3559 , \3560 , \3561 , \3562 ,
         \3563 , \3564 , \3565 , \3566 , \3567 , \3568 , \3569 , \3570 , \3571 , \3572 ,
         \3573 , \3574 , \3575 , \3576 , \3577 , \3578 , \3579 , \3580 , \3581 , \3582 ,
         \3583 , \3584 , \3585 , \3586 , \3587 , \3588 , \3589 , \3590 , \3591 , \3592 ,
         \3593 , \3594 , \3595 , \3596 , \3597 , \3598 , \3599 , \3600 , \3601 , \3602 ,
         \3603 , \3604 , \3605 , \3606 , \3607 , \3608 , \3609 , \3610 , \3611 , \3612 ,
         \3613 , \3614 , \3615 , \3616 , \3617 , \3618 , \3619 , \3620 , \3621 , \3622 ,
         \3623 , \3624 , \3625 , \3626 , \3627 , \3628 , \3629 , \3630 , \3631 , \3632 ,
         \3633 , \3634 , \3635 , \3636 , \3637 , \3638 , \3639 , \3640 , \3641 , \3642 ,
         \3643 , \3644 , \3645 , \3646 , \3647 , \3648 , \3649 , \3650 , \3651 , \3652 ,
         \3653 , \3654 , \3655 , \3656 , \3657 , \3658 , \3659 , \3660 , \3661 , \3662 ,
         \3663 , \3664 , \3665 , \3666 , \3667 , \3668 , \3669 , \3670 , \3671 , \3672 ,
         \3673 , \3674 , \3675 , \3676 , \3677 , \3678 , \3679 , \3680 , \3681 , \3682 ,
         \3683 , \3684 , \3685 , \3686 , \3687 , \3688 , \3689 , \3690 , \3691 , \3692 ,
         \3693 , \3694 , \3695 , \3696 , \3697 , \3698 , \3699 , \3700 , \3701 , \3702 ,
         \3703 , \3704 , \3705 , \3706 , \3707 , \3708 , \3709 , \3710 , \3711 , \3712 ,
         \3713 , \3714 , \3715 , \3716 , \3717 , \3718 , \3719 , \3720 , \3721 , \3722 ,
         \3723 , \3724 , \3725 , \3726 , \3727 , \3728 , \3729 , \3730 , \3731 , \3732 ,
         \3733 , \3734 , \3735 , \3736 , \3737 , \3738 , \3739 , \3740 , \3741 , \3742 ,
         \3743 , \3744 , \3745 , \3746 , \3747 , \3748 , \3749 , \3750 , \3751 , \3752 ,
         \3753 , \3754 , \3755 , \3756 , \3757 , \3758 , \3759 , \3760 , \3761 , \3762 ,
         \3763 , \3764 , \3765 , \3766 , \3767 , \3768 , \3769 , \3770 , \3771 , \3772 ,
         \3773 , \3774 , \3775 , \3776 , \3777 , \3778 , \3779 , \3780 , \3781 , \3782 ,
         \3783 , \3784 , \3785 , \3786 , \3787 , \3788 , \3789 , \3790 , \3791 , \3792 ,
         \3793 , \3794 , \3795 , \3796 , \3797 , \3798 , \3799 , \3800 , \3801 , \3802 ,
         \3803 , \3804 , \3805 , \3806 , \3807 , \3808 , \3809 , \3810 , \3811 , \3812 ,
         \3813 , \3814 , \3815 , \3816 , \3817 , \3818 , \3819 , \3820 , \3821 , \3822 ,
         \3823 , \3824 , \3825 , \3826 , \3827 , \3828 , \3829 , \3830 , \3831 , \3832 ,
         \3833 , \3834 , \3835 , \3836 , \3837 , \3838 , \3839 , \3840 , \3841 , \3842 ,
         \3843 , \3844 , \3845 , \3846 , \3847 , \3848 , \3849 , \3850 , \3851 , \3852 ,
         \3853 , \3854 , \3855 , \3856 , \3857 , \3858 , \3859 , \3860 , \3861 , \3862 ,
         \3863 , \3864 , \3865 , \3866 , \3867 , \3868 , \3869 , \3870 , \3871 , \3872 ,
         \3873 , \3874 , \3875 , \3876 , \3877 , \3878 , \3879 , \3880 , \3881 , \3882 ,
         \3883 , \3884 , \3885 , \3886 , \3887 , \3888 , \3889 , \3890 , \3891 , \3892 ,
         \3893 , \3894 , \3895 , \3896 , \3897 , \3898 , \3899 , \3900 , \3901 , \3902 ,
         \3903 , \3904 , \3905 , \3906 , \3907 , \3908 , \3909 , \3910 , \3911 , \3912 ,
         \3913 , \3914 , \3915 , \3916 , \3917 , \3918 , \3919 , \3920 , \3921 , \3922 ,
         \3923 , \3924 , \3925 , \3926 , \3927 , \3928 , \3929 , \3930 , \3931 , \3932 ,
         \3933 , \3934 , \3935 , \3936 , \3937 , \3938 , \3939 , \3940 , \3941 , \3942 ,
         \3943 , \3944 , \3945 , \3946 , \3947 , \3948 , \3949 , \3950 , \3951 , \3952 ,
         \3953 , \3954 , \3955 , \3956 , \3957 , \3958 , \3959 , \3960 , \3961 , \3962 ,
         \3963 , \3964 , \3965 , \3966 , \3967 , \3968 , \3969 , \3970 , \3971 , \3972 ,
         \3973 , \3974 , \3975 , \3976 , \3977 , \3978 , \3979 , \3980 , \3981 , \3982 ,
         \3983 , \3984 , \3985 , \3986 , \3987 , \3988 , \3989 , \3990 , \3991 , \3992 ,
         \3993 , \3994 , \3995 , \3996 , \3997 , \3998 , \3999 , \4000 , \4001 , \4002 ,
         \4003 , \4004 , \4005 , \4006 , \4007 , \4008 , \4009 , \4010 , \4011 , \4012 ,
         \4013 , \4014 , \4015 , \4016 , \4017 , \4018 , \4019 , \4020 , \4021 , \4022 ,
         \4023 , \4024 , \4025 , \4026 , \4027 , \4028 , \4029 , \4030 , \4031 , \4032 ,
         \4033 , \4034 , \4035 , \4036 , \4037 , \4038 , \4039 , \4040 , \4041 , \4042 ,
         \4043 , \4044 , \4045 , \4046 , \4047 , \4048 , \4049 , \4050 , \4051 , \4052 ,
         \4053 , \4054 , \4055 , \4056 , \4057 , \4058 , \4059 , \4060 , \4061 , \4062 ,
         \4063 , \4064 , \4065 , \4066 , \4067 , \4068 , \4069 , \4070 , \4071 , \4072 ,
         \4073 , \4074 , \4075 , \4076 , \4077 , \4078 , \4079 , \4080 , \4081 , \4082 ,
         \4083 , \4084 , \4085 , \4086 , \4087 , \4088 , \4089 , \4090 , \4091 , \4092 ,
         \4093 , \4094 , \4095 , \4096 , \4097 , \4098 , \4099 , \4100 , \4101 , \4102 ,
         \4103 , \4104 , \4105 , \4106 , \4107 , \4108 , \4109 , \4110 , \4111 , \4112 ,
         \4113 , \4114 , \4115 , \4116 , \4117 , \4118 , \4119 , \4120 , \4121 , \4122 ,
         \4123 , \4124 , \4125 , \4126 , \4127 , \4128 , \4129 , \4130 , \4131 , \4132 ,
         \4133 , \4134 , \4135 , \4136 , \4137 , \4138 , \4139 , \4140 , \4141 , \4142 ,
         \4143 , \4144 , \4145 , \4146 , \4147 , \4148 , \4149 , \4150 , \4151 , \4152 ,
         \4153 , \4154 , \4155 , \4156 , \4157 , \4158 , \4159 , \4160 , \4161 , \4162 ,
         \4163 , \4164 , \4165 , \4166 , \4167 , \4168 , \4169 , \4170 , \4171 , \4172 ,
         \4173 , \4174 , \4175 , \4176 , \4177 , \4178 , \4179 , \4180 , \4181 , \4182 ,
         \4183 , \4184 , \4185 , \4186 , \4187 , \4188 , \4189 , \4190 , \4191 , \4192 ,
         \4193 , \4194 , \4195 , \4196 , \4197 , \4198 , \4199 , \4200 , \4201 , \4202 ,
         \4203 , \4204 , \4205 , \4206 , \4207 , \4208 , \4209 , \4210 , \4211 , \4212 ,
         \4213 , \4214 , \4215 , \4216 , \4217 , \4218 , \4219 , \4220 , \4221 , \4222 ,
         \4223 , \4224 , \4225 , \4226 , \4227 , \4228 , \4229 , \4230 , \4231 , \4232 ,
         \4233 , \4234 , \4235 , \4236 , \4237 , \4238 , \4239 , \4240 , \4241 , \4242 ,
         \4243 , \4244 , \4245 , \4246 , \4247 , \4248 , \4249 , \4250 , \4251 , \4252 ,
         \4253 , \4254 , \4255 , \4256 , \4257 , \4258 , \4259 , \4260 , \4261 , \4262 ,
         \4263 , \4264 , \4265 , \4266 , \4267 , \4268 , \4269 , \4270 , \4271 , \4272 ,
         \4273 , \4274 , \4275 , \4276 , \4277 , \4278 , \4279 , \4280 , \4281 , \4282 ,
         \4283 , \4284 , \4285 , \4286 , \4287 , \4288 , \4289 , \4290 , \4291 , \4292 ,
         \4293 , \4294 , \4295 , \4296 , \4297 , \4298 , \4299 , \4300 , \4301 , \4302 ,
         \4303 , \4304 , \4305 , \4306 , \4307 , \4308 , \4309 , \4310 , \4311 , \4312 ,
         \4313 , \4314 , \4315 , \4316 , \4317 , \4318 , \4319 , \4320 , \4321 , \4322 ,
         \4323 , \4324 , \4325 , \4326 , \4327 , \4328 , \4329 , \4330 , \4331 , \4332 ,
         \4333 , \4334 , \4335 , \4336 , \4337 , \4338 , \4339 , \4340 , \4341 , \4342 ,
         \4343 , \4344 , \4345 , \4346 , \4347 , \4348 , \4349 , \4350 , \4351 , \4352 ,
         \4353 , \4354 , \4355 , \4356 , \4357 , \4358 , \4359 , \4360 , \4361 , \4362 ,
         \4363 , \4364 , \4365 , \4366 , \4367 , \4368 , \4369 , \4370 , \4371 , \4372 ,
         \4373 , \4374 , \4375 , \4376 , \4377 , \4378 , \4379 , \4380 , \4381 , \4382 ,
         \4383 , \4384 , \4385 , \4386 , \4387 , \4388 , \4389 , \4390 , \4391 , \4392 ,
         \4393 , \4394 , \4395 , \4396 , \4397 , \4398 , \4399 , \4400 , \4401 , \4402 ,
         \4403 , \4404 , \4405 , \4406 , \4407 , \4408 , \4409 , \4410 , \4411 , \4412 ,
         \4413 , \4414 , \4415 , \4416 , \4417 , \4418 , \4419 , \4420 , \4421 , \4422 ,
         \4423 , \4424 , \4425 , \4426 , \4427 , \4428 , \4429 , \4430 , \4431 , \4432 ,
         \4433 , \4434 , \4435 , \4436 , \4437 , \4438 , \4439 , \4440 , \4441 , \4442 ,
         \4443 , \4444 , \4445 , \4446 , \4447 , \4448 , \4449 , \4450 , \4451 , \4452 ,
         \4453 , \4454 , \4455 , \4456 , \4457 , \4458 , \4459 , \4460 , \4461 , \4462 ,
         \4463 , \4464 , \4465 , \4466 , \4467 , \4468 , \4469 , \4470 , \4471 , \4472 ,
         \4473 , \4474 , \4475 , \4476 , \4477 , \4478 , \4479 , \4480 , \4481 , \4482 ,
         \4483 , \4484 , \4485 , \4486 , \4487 , \4488 , \4489 , \4490 , \4491 , \4492 ,
         \4493 , \4494 , \4495 , \4496 , \4497 , \4498 , \4499 , \4500 , \4501 , \4502 ,
         \4503 , \4504 , \4505 , \4506 , \4507 , \4508 , \4509 , \4510 , \4511 , \4512 ,
         \4513 , \4514 , \4515 , \4516 , \4517 , \4518 , \4519 , \4520 , \4521 , \4522 ,
         \4523 , \4524 , \4525 , \4526 , \4527 , \4528 , \4529 , \4530 , \4531 , \4532 ,
         \4533 , \4534 , \4535 , \4536 , \4537 , \4538 , \4539 , \4540 , \4541 , \4542 ,
         \4543 , \4544 , \4545 , \4546 , \4547 , \4548 , \4549 , \4550 , \4551 , \4552 ,
         \4553 , \4554 , \4555 , \4556 , \4557 , \4558 , \4559 , \4560 , \4561 , \4562 ,
         \4563 , \4564 , \4565 , \4566 , \4567 , \4568 , \4569 , \4570 , \4571 , \4572 ,
         \4573 , \4574 , \4575 , \4576 , \4577 , \4578 , \4579 , \4580 , \4581 , \4582 ,
         \4583 , \4584 , \4585 , \4586 , \4587 , \4588 , \4589 , \4590 , \4591 , \4592 ,
         \4593 , \4594 , \4595 , \4596 , \4597 , \4598 , \4599 , \4600 , \4601 , \4602 ,
         \4603 , \4604 , \4605 , \4606 , \4607 , \4608 , \4609 , \4610 , \4611 , \4612 ,
         \4613 , \4614 , \4615 , \4616 , \4617 , \4618 , \4619 , \4620 , \4621 , \4622 ,
         \4623 , \4624 , \4625 , \4626 , \4627 , \4628 , \4629 , \4630 , \4631 , \4632 ,
         \4633 , \4634 , \4635 , \4636 , \4637 , \4638 , \4639 , \4640 , \4641 , \4642 ,
         \4643 , \4644 , \4645 , \4646 , \4647 , \4648 , \4649 , \4650 , \4651 , \4652 ,
         \4653 , \4654 , \4655 , \4656 , \4657 , \4658 , \4659 , \4660 , \4661 , \4662 ,
         \4663 , \4664 , \4665 , \4666 , \4667 , \4668 , \4669 , \4670 , \4671 , \4672 ,
         \4673 , \4674 , \4675 , \4676 , \4677 , \4678 , \4679 , \4680 , \4681 , \4682 ,
         \4683 , \4684 , \4685 , \4686 , \4687 , \4688 , \4689 , \4690 , \4691 , \4692 ,
         \4693 , \4694 , \4695 , \4696 , \4697 , \4698 , \4699 , \4700 , \4701 , \4702 ,
         \4703 , \4704 , \4705 , \4706 , \4707 , \4708 , \4709 , \4710 , \4711 , \4712 ,
         \4713 , \4714 , \4715 , \4716 , \4717 , \4718 , \4719 , \4720 , \4721 , \4722 ,
         \4723 , \4724 , \4725 , \4726 , \4727 , \4728 , \4729 , \4730 , \4731 , \4732 ,
         \4733 , \4734 , \4735 , \4736 , \4737 , \4738 , \4739 , \4740 , \4741 , \4742 ,
         \4743 , \4744 , \4745 , \4746 , \4747 , \4748 , \4749 , \4750 , \4751 , \4752 ,
         \4753 , \4754 , \4755 , \4756 , \4757 , \4758 , \4759 , \4760 , \4761 , \4762 ,
         \4763 , \4764 , \4765 , \4766 , \4767 , \4768 , \4769 , \4770 , \4771 , \4772 ,
         \4773 , \4774 , \4775 , \4776 , \4777 , \4778 , \4779 , \4780 , \4781 , \4782 ,
         \4783 , \4784 , \4785 , \4786 , \4787 , \4788 , \4789 , \4790 , \4791 , \4792 ,
         \4793 , \4794 , \4795 , \4796 , \4797 , \4798 , \4799 , \4800 , \4801 , \4802 ,
         \4803 , \4804 , \4805 , \4806 , \4807 , \4808 , \4809 , \4810 , \4811 , \4812 ,
         \4813 , \4814 , \4815 , \4816 , \4817 , \4818 , \4819 , \4820 , \4821 , \4822 ,
         \4823 , \4824 , \4825 , \4826 , \4827 , \4828 , \4829 , \4830 , \4831 , \4832 ,
         \4833 , \4834 , \4835 , \4836 , \4837 , \4838 , \4839 , \4840 , \4841 , \4842 ,
         \4843 , \4844 , \4845 , \4846 , \4847 , \4848 , \4849 , \4850 , \4851 , \4852 ,
         \4853 , \4854 , \4855 , \4856 , \4857 , \4858 , \4859 , \4860 , \4861 , \4862 ,
         \4863 , \4864 , \4865 , \4866 , \4867 , \4868 , \4869 , \4870 , \4871 , \4872 ,
         \4873 , \4874 , \4875 , \4876 , \4877 , \4878 , \4879 , \4880 , \4881 , \4882 ,
         \4883 , \4884 , \4885 , \4886 , \4887 , \4888 , \4889 , \4890 , \4891 , \4892 ,
         \4893 , \4894 , \4895 , \4896 , \4897 , \4898 , \4899 , \4900 , \4901 , \4902 ,
         \4903 , \4904 , \4905 , \4906 , \4907 , \4908 , \4909 , \4910 , \4911 , \4912 ,
         \4913 , \4914 , \4915 , \4916 , \4917 , \4918 , \4919 , \4920 , \4921 , \4922 ,
         \4923 , \4924 , \4925 , \4926 , \4927 , \4928 , \4929 , \4930 , \4931 , \4932 ,
         \4933 , \4934 , \4935 , \4936 , \4937 , \4938 , \4939 , \4940 , \4941 , \4942 ,
         \4943 , \4944 , \4945 , \4946 , \4947 , \4948 , \4949 , \4950 , \4951 , \4952 ,
         \4953 , \4954 , \4955 , \4956 , \4957 , \4958 , \4959 , \4960 , \4961 , \4962 ,
         \4963 , \4964 , \4965 , \4966 , \4967 , \4968 , \4969 , \4970 , \4971 , \4972 ,
         \4973 , \4974 , \4975 , \4976 , \4977 , \4978 , \4979 , \4980 , \4981 , \4982 ,
         \4983 , \4984 , \4985 , \4986 , \4987 , \4988 , \4989 , \4990 , \4991 , \4992 ,
         \4993 , \4994 , \4995 , \4996 , \4997 , \4998 , \4999 , \5000 , \5001 , \5002 ,
         \5003 , \5004 , \5005 , \5006 , \5007 , \5008 , \5009 , \5010 , \5011 , \5012 ,
         \5013 , \5014 , \5015 , \5016 , \5017 , \5018 , \5019 , \5020 , \5021 , \5022 ,
         \5023 , \5024 , \5025 , \5026 , \5027 , \5028 , \5029 , \5030 , \5031 , \5032 ,
         \5033 , \5034 , \5035 , \5036 , \5037 , \5038 , \5039 , \5040 , \5041 , \5042 ,
         \5043 , \5044 , \5045 , \5046 , \5047 , \5048 , \5049 , \5050 , \5051 , \5052 ,
         \5053 , \5054 , \5055 , \5056 , \5057 , \5058 , \5059 , \5060 , \5061 , \5062 ,
         \5063 , \5064 , \5065 , \5066 , \5067 , \5068 , \5069 , \5070 , \5071 , \5072 ,
         \5073 , \5074 , \5075 , \5076 , \5077 , \5078 , \5079 , \5080 , \5081 , \5082 ,
         \5083 , \5084 , \5085 , \5086 , \5087 , \5088 , \5089 , \5090 , \5091 , \5092 ,
         \5093 , \5094 , \5095 , \5096 , \5097 , \5098 , \5099 , \5100 , \5101 , \5102 ,
         \5103 , \5104 , \5105 , \5106 , \5107 , \5108 , \5109 , \5110 , \5111 , \5112 ,
         \5113 , \5114 , \5115 , \5116 , \5117 , \5118 , \5119 , \5120 , \5121 , \5122 ,
         \5123 , \5124 , \5125 , \5126 , \5127 , \5128 , \5129 , \5130 , \5131 , \5132 ,
         \5133 , \5134 , \5135 , \5136 , \5137 , \5138 , \5139 , \5140 , \5141 , \5142 ,
         \5143 , \5144 , \5145 , \5146 , \5147 , \5148 , \5149 , \5150 , \5151 , \5152 ,
         \5153 , \5154 , \5155 , \5156 , \5157 , \5158 , \5159 , \5160 , \5161 , \5162 ,
         \5163 , \5164 , \5165 , \5166 , \5167 , \5168 , \5169 , \5170 , \5171 , \5172 ,
         \5173 , \5174 , \5175 , \5176 , \5177 , \5178 , \5179 , \5180 , \5181 , \5182 ,
         \5183 , \5184 , \5185 , \5186 , \5187 , \5188 , \5189 , \5190 , \5191 , \5192 ,
         \5193 , \5194 , \5195 , \5196 , \5197 , \5198 , \5199 , \5200 , \5201 , \5202 ,
         \5203 , \5204 , \5205 , \5206 , \5207 , \5208 , \5209 , \5210 , \5211 , \5212 ,
         \5213 , \5214 , \5215 , \5216 , \5217 , \5218 , \5219 , \5220 , \5221 , \5222 ,
         \5223 , \5224 , \5225 , \5226 , \5227 , \5228 , \5229 , \5230 , \5231 , \5232 ,
         \5233 , \5234 , \5235 , \5236 , \5237 , \5238 , \5239 , \5240 , \5241 , \5242 ,
         \5243 , \5244 , \5245 , \5246 , \5247 , \5248 , \5249 , \5250 , \5251 , \5252 ,
         \5253 , \5254 , \5255 , \5256 , \5257 , \5258 , \5259 , \5260 , \5261 , \5262 ,
         \5263 , \5264 , \5265 , \5266 , \5267 , \5268 , \5269 , \5270 , \5271 , \5272 ,
         \5273 , \5274 , \5275 , \5276 , \5277 , \5278 , \5279 , \5280 , \5281 , \5282 ,
         \5283 , \5284 , \5285 , \5286 , \5287 , \5288 , \5289 , \5290 , \5291 , \5292 ,
         \5293 , \5294 , \5295 , \5296 , \5297 , \5298 , \5299 , \5300 , \5301 , \5302 ,
         \5303 , \5304 , \5305 , \5306 , \5307 , \5308 , \5309 , \5310 , \5311 , \5312 ,
         \5313 , \5314 , \5315 , \5316 , \5317 , \5318 , \5319 , \5320 , \5321 , \5322 ,
         \5323 , \5324 , \5325 , \5326 , \5327 , \5328 , \5329 , \5330 , \5331 , \5332 ,
         \5333 , \5334 , \5335 , \5336 , \5337 , \5338 , \5339 , \5340 , \5341 , \5342 ,
         \5343 , \5344 , \5345 , \5346 , \5347 , \5348 , \5349 , \5350 , \5351 , \5352 ,
         \5353 , \5354 , \5355 , \5356 , \5357 , \5358 , \5359 , \5360 , \5361 , \5362 ,
         \5363 , \5364 , \5365 , \5366 , \5367 , \5368 , \5369 , \5370 , \5371 , \5372 ,
         \5373 , \5374 , \5375 , \5376 , \5377 , \5378 , \5379 , \5380 , \5381 , \5382 ,
         \5383 , \5384 , \5385 , \5386 , \5387 , \5388 , \5389 , \5390 , \5391 , \5392 ,
         \5393 , \5394 , \5395 , \5396 , \5397 , \5398 , \5399 , \5400 , \5401 , \5402 ,
         \5403 , \5404 , \5405 , \5406 , \5407 , \5408 , \5409 , \5410 , \5411 , \5412 ,
         \5413 , \5414 , \5415 , \5416 , \5417 , \5418 , \5419 , \5420 , \5421 , \5422 ,
         \5423 , \5424 , \5425 , \5426 , \5427 , \5428 , \5429 , \5430 , \5431 , \5432 ,
         \5433 , \5434 , \5435 , \5436 , \5437 , \5438 , \5439 , \5440 , \5441 , \5442 ,
         \5443 , \5444 , \5445 , \5446 , \5447 , \5448 , \5449 , \5450 , \5451 , \5452 ,
         \5453 , \5454 , \5455 , \5456 , \5457 , \5458 , \5459 , \5460 , \5461 , \5462 ,
         \5463 , \5464 , \5465 , \5466 , \5467 , \5468 , \5469 , \5470 , \5471 , \5472 ,
         \5473 , \5474 , \5475 , \5476 , \5477 , \5478 , \5479 , \5480 , \5481 , \5482 ,
         \5483 , \5484 , \5485 , \5486 , \5487 , \5488 , \5489 , \5490 , \5491 , \5492 ,
         \5493 , \5494 , \5495 , \5496 , \5497 , \5498 , \5499 , \5500 , \5501 , \5502 ,
         \5503 , \5504 , \5505 , \5506 , \5507 , \5508 , \5509 , \5510 , \5511 , \5512 ,
         \5513 , \5514 , \5515 , \5516 , \5517 , \5518 , \5519 , \5520 , \5521 , \5522 ,
         \5523 , \5524 , \5525 , \5526 , \5527 , \5528 , \5529 , \5530 , \5531 , \5532 ,
         \5533 , \5534 , \5535 , \5536 , \5537 , \5538 , \5539 , \5540 , \5541 , \5542 ,
         \5543 , \5544 , \5545 , \5546 , \5547 , \5548 , \5549 , \5550 , \5551 , \5552 ,
         \5553 , \5554 , \5555 , \5556 , \5557 , \5558 , \5559 , \5560 , \5561 , \5562 ,
         \5563 , \5564 , \5565 , \5566 , \5567 , \5568 , \5569 , \5570 , \5571 , \5572 ,
         \5573 , \5574 , \5575 , \5576 , \5577 , \5578 , \5579 , \5580 , \5581 , \5582 ,
         \5583 , \5584 , \5585 , \5586 , \5587 , \5588 , \5589 , \5590 , \5591 , \5592 ,
         \5593 , \5594 , \5595 , \5596 , \5597 , \5598 , \5599 , \5600 , \5601 , \5602 ,
         \5603 , \5604 , \5605 , \5606 , \5607 , \5608 , \5609 , \5610 , \5611 , \5612 ,
         \5613 , \5614 , \5615 , \5616 , \5617 , \5618 , \5619 , \5620 , \5621 , \5622 ,
         \5623 , \5624 , \5625 , \5626 , \5627 , \5628 , \5629 , \5630 , \5631 , \5632 ,
         \5633 , \5634 , \5635 , \5636 , \5637 , \5638 , \5639 , \5640 , \5641 , \5642 ,
         \5643 , \5644 , \5645 , \5646 , \5647 , \5648 , \5649 , \5650 , \5651 , \5652 ,
         \5653 , \5654 , \5655 , \5656 , \5657 , \5658 , \5659 , \5660 , \5661 , \5662 ,
         \5663 , \5664 , \5665 , \5666 , \5667 , \5668 , \5669 , \5670 , \5671 , \5672 ,
         \5673 , \5674 , \5675 , \5676 , \5677 , \5678 , \5679 , \5680 , \5681 , \5682 ,
         \5683 , \5684 , \5685 , \5686 , \5687 , \5688 , \5689 , \5690 , \5691 , \5692 ,
         \5693 , \5694 , \5695 , \5696 , \5697 , \5698 , \5699 , \5700 , \5701 , \5702 ,
         \5703 , \5704 , \5705 , \5706 , \5707 , \5708 , \5709 , \5710 , \5711 , \5712 ,
         \5713 , \5714 , \5715 , \5716 , \5717 , \5718 , \5719 , \5720 , \5721 , \5722 ,
         \5723 , \5724 , \5725 , \5726 , \5727 , \5728 , \5729 , \5730 , \5731 , \5732 ,
         \5733 , \5734 , \5735 , \5736 , \5737 , \5738 , \5739 , \5740 , \5741 , \5742 ,
         \5743 , \5744 , \5745 , \5746 , \5747 , \5748 , \5749 , \5750 , \5751 , \5752 ,
         \5753 , \5754 , \5755 , \5756 , \5757 , \5758 , \5759 , \5760 , \5761 , \5762 ,
         \5763 , \5764 , \5765 , \5766 , \5767 , \5768 , \5769 , \5770 , \5771 , \5772 ,
         \5773 , \5774 , \5775 , \5776 , \5777 , \5778 , \5779 , \5780 , \5781 , \5782 ,
         \5783 , \5784 , \5785 , \5786 , \5787 , \5788 , \5789 , \5790 , \5791 , \5792 ,
         \5793 , \5794 , \5795 , \5796 , \5797 , \5798 , \5799 , \5800 , \5801 , \5802 ,
         \5803 , \5804 , \5805 , \5806 , \5807 , \5808 , \5809 , \5810 , \5811 , \5812 ,
         \5813 , \5814 , \5815 , \5816 , \5817 , \5818 , \5819 , \5820 , \5821 , \5822 ,
         \5823 , \5824 , \5825 , \5826 , \5827 , \5828 , \5829 , \5830 , \5831 , \5832 ,
         \5833 , \5834 , \5835 , \5836 , \5837 , \5838 , \5839 , \5840 , \5841 , \5842 ,
         \5843 , \5844 , \5845 , \5846 , \5847 , \5848 , \5849 , \5850 , \5851 , \5852 ,
         \5853 , \5854 , \5855 , \5856 , \5857 , \5858 , \5859 , \5860 , \5861 , \5862 ,
         \5863 , \5864 , \5865 , \5866 , \5867 , \5868 , \5869 , \5870 , \5871 , \5872 ,
         \5873 , \5874 , \5875 , \5876 , \5877 , \5878 , \5879 , \5880 , \5881 , \5882 ,
         \5883 , \5884 , \5885 , \5886 , \5887 , \5888 , \5889 , \5890 , \5891 , \5892 ,
         \5893 , \5894 , \5895 , \5896 , \5897 , \5898 , \5899 , \5900 , \5901 , \5902 ,
         \5903 , \5904 , \5905 , \5906 , \5907 , \5908 , \5909 , \5910 , \5911 , \5912 ,
         \5913 , \5914 , \5915 , \5916 , \5917 , \5918 , \5919 , \5920 , \5921 , \5922 ,
         \5923 , \5924 , \5925 , \5926 , \5927 , \5928 , \5929 , \5930 , \5931 , \5932 ,
         \5933 , \5934 , \5935 , \5936 , \5937 , \5938 , \5939 , \5940 , \5941 , \5942 ,
         \5943 , \5944 , \5945 , \5946 , \5947 , \5948 , \5949 , \5950 , \5951 , \5952 ,
         \5953 , \5954 , \5955 , \5956 , \5957 , \5958 , \5959 , \5960 , \5961 , \5962 ,
         \5963 , \5964 , \5965 , \5966 , \5967 , \5968 , \5969 , \5970 , \5971 , \5972 ,
         \5973 , \5974 , \5975 , \5976 , \5977 , \5978 , \5979 , \5980 , \5981 , \5982 ,
         \5983 , \5984 , \5985 , \5986 , \5987 , \5988 , \5989 , \5990 , \5991 , \5992 ,
         \5993 , \5994 , \5995 , \5996 , \5997 , \5998 , \5999 , \6000 , \6001 , \6002 ,
         \6003 , \6004 , \6005 , \6006 , \6007 , \6008 , \6009 , \6010 , \6011 , \6012 ,
         \6013 , \6014 , \6015 , \6016 , \6017 , \6018 , \6019 , \6020 , \6021 , \6022 ,
         \6023 , \6024 , \6025 , \6026 , \6027 , \6028 , \6029 , \6030 , \6031 , \6032 ,
         \6033 , \6034 , \6035 , \6036 , \6037 , \6038 , \6039 , \6040 , \6041 , \6042 ,
         \6043 , \6044 , \6045 , \6046 , \6047 , \6048 , \6049 , \6050 , \6051 , \6052 ,
         \6053 , \6054 , \6055 , \6056 , \6057 , \6058 , \6059 , \6060 , \6061 , \6062 ,
         \6063 , \6064 , \6065 , \6066 , \6067 , \6068 , \6069 , \6070 , \6071 , \6072 ,
         \6073 , \6074 , \6075 , \6076 , \6077 , \6078 , \6079 , \6080 , \6081 , \6082 ,
         \6083 , \6084 , \6085 , \6086 , \6087 , \6088 , \6089 , \6090 , \6091 , \6092 ,
         \6093 , \6094 , \6095 , \6096 , \6097 , \6098 , \6099 , \6100 , \6101 , \6102 ,
         \6103 , \6104 , \6105 , \6106 , \6107 , \6108 , \6109 , \6110 , \6111 , \6112 ,
         \6113 , \6114 , \6115 , \6116 , \6117 , \6118 , \6119 , \6120 , \6121 , \6122 ,
         \6123 , \6124 , \6125 , \6126 , \6127 , \6128 , \6129 , \6130 , \6131 , \6132 ,
         \6133 , \6134 , \6135 , \6136 , \6137 , \6138 , \6139 , \6140 , \6141 , \6142 ,
         \6143 , \6144 , \6145 , \6146 , \6147 , \6148 , \6149 , \6150 , \6151 , \6152 ,
         \6153 , \6154 , \6155 , \6156 , \6157 , \6158 , \6159 , \6160 , \6161 , \6162 ,
         \6163 , \6164 , \6165 , \6166 , \6167 , \6168 , \6169 , \6170 , \6171 , \6172 ,
         \6173 , \6174 , \6175 , \6176 , \6177 , \6178 , \6179 , \6180 , \6181 , \6182 ,
         \6183 , \6184 , \6185 , \6186 , \6187 , \6188 , \6189 , \6190 , \6191 , \6192 ,
         \6193 , \6194 , \6195 , \6196 , \6197 , \6198 , \6199 , \6200 , \6201 , \6202 ,
         \6203 , \6204 , \6205 , \6206 , \6207 , \6208 , \6209 , \6210 , \6211 , \6212 ,
         \6213 , \6214 , \6215 , \6216 , \6217 , \6218 , \6219 , \6220 , \6221 , \6222 ,
         \6223 , \6224 , \6225 , \6226 , \6227 , \6228 , \6229 , \6230 , \6231 , \6232 ,
         \6233 , \6234 , \6235 , \6236 , \6237 , \6238 , \6239 , \6240 , \6241 , \6242 ,
         \6243 , \6244 , \6245 , \6246 , \6247 , \6248 , \6249 , \6250 , \6251 , \6252 ,
         \6253 , \6254 , \6255 , \6256 , \6257 , \6258 , \6259 , \6260 , \6261 , \6262 ,
         \6263 , \6264 , \6265 , \6266 , \6267 , \6268 , \6269 , \6270 , \6271 , \6272 ,
         \6273 , \6274 , \6275 , \6276 , \6277 , \6278 , \6279 , \6280 , \6281 , \6282 ,
         \6283 , \6284 , \6285 , \6286 , \6287 , \6288 , \6289 , \6290 , \6291 , \6292 ,
         \6293 , \6294 , \6295 , \6296 , \6297 , \6298 , \6299 , \6300 , \6301 , \6302 ,
         \6303 , \6304 , \6305 , \6306 , \6307 , \6308 , \6309 , \6310 , \6311 , \6312 ,
         \6313 , \6314 , \6315 , \6316 , \6317 , \6318 , \6319 , \6320 , \6321 , \6322 ,
         \6323 , \6324 , \6325 , \6326 , \6327 , \6328 , \6329 , \6330 , \6331 , \6332 ,
         \6333 , \6334 , \6335 , \6336 , \6337 , \6338 , \6339 , \6340 , \6341 , \6342 ,
         \6343 , \6344 , \6345 , \6346 , \6347 , \6348 , \6349 , \6350 , \6351 , \6352 ,
         \6353 , \6354 , \6355 , \6356 , \6357 , \6358 , \6359 , \6360 , \6361 , \6362 ,
         \6363 , \6364 , \6365 , \6366 , \6367 , \6368 , \6369 , \6370 , \6371 , \6372 ,
         \6373 , \6374 , \6375 , \6376 , \6377 , \6378 , \6379 , \6380 , \6381 , \6382 ,
         \6383 , \6384 , \6385 , \6386 , \6387 , \6388 , \6389 , \6390 , \6391 , \6392 ,
         \6393 , \6394 , \6395 , \6396 , \6397 , \6398 , \6399 , \6400 , \6401 , \6402 ,
         \6403 , \6404 , \6405 , \6406 , \6407 , \6408 , \6409 , \6410 , \6411 , \6412 ,
         \6413 , \6414 , \6415 , \6416 , \6417 , \6418 , \6419 , \6420 , \6421 , \6422 ,
         \6423 , \6424 , \6425 , \6426 , \6427 , \6428 , \6429 , \6430 , \6431 , \6432 ,
         \6433 , \6434 , \6435 , \6436 , \6437 , \6438 , \6439 , \6440 , \6441 , \6442 ,
         \6443 , \6444 , \6445 , \6446 , \6447 , \6448 , \6449 , \6450 , \6451 , \6452 ,
         \6453 , \6454 , \6455 , \6456 , \6457 , \6458 , \6459 , \6460 , \6461 , \6462 ,
         \6463 , \6464 , \6465 , \6466 , \6467 , \6468 , \6469 , \6470 , \6471 , \6472 ,
         \6473 , \6474 , \6475 , \6476 , \6477 , \6478 , \6479 , \6480 , \6481 , \6482 ,
         \6483 , \6484 , \6485 , \6486 , \6487 , \6488 , \6489 , \6490 , \6491 , \6492 ,
         \6493 , \6494 , \6495 , \6496 , \6497 , \6498 , \6499 , \6500 , \6501 , \6502 ,
         \6503 , \6504 , \6505 , \6506 , \6507 , \6508 , \6509 , \6510 , \6511 , \6512 ,
         \6513 , \6514 , \6515 , \6516 , \6517 , \6518 , \6519 , \6520 , \6521 , \6522 ,
         \6523 , \6524 , \6525 , \6526 , \6527 , \6528 , \6529 , \6530 , \6531 , \6532 ,
         \6533 , \6534 , \6535 , \6536 , \6537 , \6538 , \6539 , \6540 , \6541 , \6542 ,
         \6543 , \6544 , \6545 , \6546 , \6547 , \6548 , \6549 , \6550 , \6551 , \6552 ,
         \6553 , \6554 , \6555 , \6556 , \6557 , \6558 , \6559 , \6560 , \6561 , \6562 ,
         \6563 , \6564 , \6565 , \6566 , \6567 , \6568 , \6569 , \6570 , \6571 , \6572 ,
         \6573 , \6574 , \6575 , \6576 , \6577 , \6578 , \6579 , \6580 , \6581 , \6582 ,
         \6583 , \6584 , \6585 , \6586 , \6587 , \6588 , \6589 , \6590 , \6591 , \6592 ,
         \6593 , \6594 , \6595 , \6596 , \6597 , \6598 , \6599 , \6600 , \6601 , \6602 ,
         \6603 , \6604 , \6605 , \6606 , \6607 , \6608 , \6609 , \6610 , \6611 , \6612 ,
         \6613 , \6614 , \6615 , \6616 , \6617 , \6618 , \6619 , \6620 , \6621 , \6622 ,
         \6623 , \6624 , \6625 , \6626 , \6627 , \6628 , \6629 , \6630 , \6631 , \6632 ,
         \6633 , \6634 , \6635 , \6636 , \6637 , \6638 , \6639 , \6640 , \6641 , \6642 ,
         \6643 , \6644 , \6645 , \6646 , \6647 , \6648 , \6649 , \6650 , \6651 , \6652 ,
         \6653 , \6654 , \6655 , \6656 , \6657 , \6658 , \6659 , \6660 , \6661 , \6662 ,
         \6663 , \6664 , \6665 , \6666 , \6667 , \6668 , \6669 , \6670 , \6671 , \6672 ,
         \6673 , \6674 , \6675 , \6676 , \6677 , \6678 , \6679 , \6680 , \6681 , \6682 ,
         \6683 , \6684 , \6685 , \6686 , \6687 , \6688 , \6689 , \6690 , \6691 , \6692 ,
         \6693 , \6694 , \6695 , \6696 , \6697 , \6698 , \6699 , \6700 , \6701 , \6702 ,
         \6703 , \6704 , \6705 , \6706 , \6707 , \6708 , \6709 , \6710 , \6711 , \6712 ,
         \6713 , \6714 , \6715 , \6716 , \6717 , \6718 , \6719 , \6720 , \6721 , \6722 ,
         \6723 , \6724 , \6725 , \6726 , \6727 , \6728 , \6729 , \6730 , \6731 , \6732 ,
         \6733 , \6734 , \6735 , \6736 , \6737 , \6738 , \6739 , \6740 , \6741 , \6742 ,
         \6743 , \6744 , \6745 , \6746 , \6747 , \6748 , \6749 , \6750 , \6751 , \6752 ,
         \6753 , \6754 , \6755 , \6756 , \6757 , \6758 , \6759 , \6760 , \6761 , \6762 ,
         \6763 , \6764 , \6765 , \6766 , \6767 , \6768 , \6769 , \6770 , \6771 , \6772 ,
         \6773 , \6774 , \6775 , \6776 , \6777 , \6778 , \6779 , \6780 , \6781 , \6782 ,
         \6783 , \6784 , \6785 , \6786 , \6787 , \6788 , \6789 , \6790 , \6791 , \6792 ,
         \6793 , \6794 , \6795 , \6796 , \6797 , \6798 , \6799 , \6800 , \6801 , \6802 ,
         \6803 , \6804 , \6805 , \6806 , \6807 , \6808 , \6809 , \6810 , \6811 , \6812 ,
         \6813 , \6814 , \6815 , \6816 , \6817 , \6818 , \6819 , \6820 , \6821 , \6822 ,
         \6823 , \6824 , \6825 , \6826 , \6827 , \6828 , \6829 , \6830 , \6831 , \6832 ,
         \6833 , \6834 , \6835 , \6836 , \6837 , \6838 , \6839 , \6840 , \6841 , \6842 ,
         \6843 , \6844 , \6845 , \6846 , \6847 , \6848 , \6849 , \6850 , \6851 , \6852 ,
         \6853 , \6854 , \6855 , \6856 , \6857 , \6858 , \6859 , \6860 , \6861 , \6862 ,
         \6863 , \6864 , \6865 , \6866 , \6867 , \6868 , \6869 , \6870 , \6871 , \6872 ,
         \6873 , \6874 , \6875 , \6876 , \6877 , \6878 , \6879 , \6880 , \6881 , \6882 ,
         \6883 , \6884 , \6885 , \6886 , \6887 , \6888 , \6889 , \6890 , \6891 , \6892 ,
         \6893 , \6894 , \6895 , \6896 , \6897 , \6898 , \6899 , \6900 , \6901 , \6902 ,
         \6903 , \6904 , \6905 , \6906 , \6907 , \6908 , \6909 , \6910 , \6911 , \6912 ,
         \6913 , \6914 , \6915 , \6916 , \6917 , \6918 , \6919 , \6920 , \6921 , \6922 ,
         \6923 , \6924 , \6925 , \6926 , \6927 , \6928 , \6929 , \6930 , \6931 , \6932 ,
         \6933 , \6934 , \6935 , \6936 , \6937 , \6938 , \6939 , \6940 , \6941 , \6942 ,
         \6943 , \6944 , \6945 , \6946 , \6947 , \6948 , \6949 , \6950 , \6951 , \6952 ,
         \6953 , \6954 , \6955 , \6956 , \6957 , \6958 , \6959 , \6960 , \6961 , \6962 ,
         \6963 , \6964 , \6965 , \6966 , \6967 , \6968 , \6969 , \6970 , \6971 , \6972 ,
         \6973 , \6974 , \6975 , \6976 , \6977 , \6978 , \6979 , \6980 , \6981 , \6982 ,
         \6983 , \6984 , \6985 , \6986 , \6987 , \6988 , \6989 , \6990 , \6991 , \6992 ,
         \6993 , \6994 , \6995 , \6996 , \6997 , \6998 , \6999 , \7000 , \7001 , \7002 ,
         \7003 , \7004 , \7005 , \7006 , \7007 , \7008 , \7009 , \7010 , \7011 , \7012 ,
         \7013 , \7014 , \7015 , \7016 , \7017 , \7018 , \7019 , \7020 , \7021 , \7022 ,
         \7023 , \7024 , \7025 , \7026 , \7027 , \7028 , \7029 , \7030 , \7031 , \7032 ,
         \7033 , \7034 , \7035 , \7036 , \7037 , \7038 , \7039 , \7040 , \7041 , \7042 ,
         \7043 , \7044 , \7045 , \7046 , \7047 , \7048 , \7049 , \7050 , \7051 , \7052 ,
         \7053 , \7054 , \7055 , \7056 , \7057 , \7058 , \7059 , \7060 , \7061 , \7062 ,
         \7063 , \7064 , \7065 , \7066 , \7067 , \7068 , \7069 , \7070 , \7071 , \7072 ,
         \7073 , \7074 , \7075 , \7076 , \7077 , \7078 , \7079 , \7080 , \7081 , \7082 ,
         \7083 , \7084 , \7085 , \7086 , \7087 , \7088 , \7089 , \7090 , \7091 , \7092 ,
         \7093 , \7094 , \7095 , \7096 , \7097 , \7098 , \7099 , \7100 , \7101 , \7102 ,
         \7103 , \7104 , \7105 , \7106 , \7107 , \7108 , \7109 , \7110 , \7111 , \7112 ,
         \7113 , \7114 , \7115 , \7116 , \7117 , \7118 , \7119 , \7120 , \7121 , \7122 ,
         \7123 , \7124 , \7125 , \7126 , \7127 , \7128 , \7129 , \7130 , \7131 , \7132 ,
         \7133 , \7134 , \7135 , \7136 , \7137 , \7138 , \7139 , \7140 , \7141 , \7142 ,
         \7143 , \7144 , \7145 , \7146 , \7147 , \7148 , \7149 , \7150 , \7151 , \7152 ,
         \7153 , \7154 , \7155 , \7156 , \7157 , \7158 , \7159 , \7160 , \7161 , \7162 ,
         \7163 , \7164 , \7165 , \7166 , \7167 , \7168 , \7169 , \7170 , \7171 , \7172 ,
         \7173 , \7174 , \7175 , \7176 , \7177 , \7178 , \7179 , \7180 , \7181 , \7182 ,
         \7183 , \7184 , \7185 , \7186 , \7187 , \7188 , \7189 , \7190 , \7191 , \7192 ,
         \7193 , \7194 , \7195 , \7196 , \7197 , \7198 , \7199 , \7200 , \7201 , \7202 ,
         \7203 , \7204 , \7205 , \7206 , \7207 , \7208 , \7209 , \7210 , \7211 , \7212 ,
         \7213 , \7214 , \7215 , \7216 , \7217 , \7218 , \7219 , \7220 , \7221 , \7222 ,
         \7223 , \7224 , \7225 , \7226 , \7227 , \7228 , \7229 , \7230 , \7231 , \7232 ,
         \7233 , \7234 , \7235 , \7236 , \7237 , \7238 , \7239 , \7240 , \7241 , \7242 ,
         \7243 , \7244 , \7245 , \7246 , \7247 , \7248 , \7249 , \7250 , \7251 , \7252 ,
         \7253 , \7254 , \7255 , \7256 , \7257 , \7258 , \7259 , \7260 , \7261 , \7262 ,
         \7263 , \7264 , \7265 , \7266 , \7267 , \7268 , \7269 , \7270 , \7271 , \7272 ,
         \7273 , \7274 , \7275 , \7276 , \7277 , \7278 , \7279 , \7280 , \7281 , \7282 ,
         \7283 , \7284 , \7285 , \7286 , \7287 , \7288 , \7289 , \7290 , \7291 , \7292 ,
         \7293 , \7294 , \7295 , \7296 , \7297 , \7298 , \7299 , \7300 , \7301 , \7302 ,
         \7303 , \7304 , \7305 , \7306 , \7307 , \7308 , \7309 , \7310 , \7311 , \7312 ,
         \7313 , \7314 , \7315 , \7316 , \7317 , \7318 , \7319 , \7320 , \7321 , \7322 ,
         \7323 , \7324 , \7325 , \7326 , \7327 , \7328 , \7329 , \7330 , \7331 , \7332 ,
         \7333 , \7334 , \7335 , \7336 , \7337 , \7338 , \7339 , \7340 , \7341 , \7342 ,
         \7343 , \7344 , \7345 , \7346 , \7347 , \7348 , \7349 , \7350 , \7351 , \7352 ,
         \7353 , \7354 , \7355 , \7356 , \7357 , \7358 , \7359 , \7360 , \7361 , \7362 ,
         \7363 , \7364 , \7365 , \7366 , \7367 , \7368 , \7369 , \7370 , \7371 , \7372 ,
         \7373 , \7374 , \7375 , \7376 , \7377 , \7378 , \7379 , \7380 , \7381 , \7382 ,
         \7383 , \7384 , \7385 , \7386 , \7387 , \7388 , \7389 , \7390 , \7391 , \7392 ,
         \7393 , \7394 , \7395 , \7396 , \7397 , \7398 , \7399 , \7400 , \7401 , \7402 ,
         \7403 , \7404 , \7405 , \7406 , \7407 , \7408 , \7409 , \7410 , \7411 , \7412 ,
         \7413 , \7414 , \7415 , \7416 , \7417 , \7418 , \7419 , \7420 , \7421 , \7422 ,
         \7423 , \7424 , \7425 , \7426 , \7427 , \7428 , \7429 , \7430 , \7431 , \7432 ,
         \7433 , \7434 , \7435 , \7436 , \7437 , \7438 , \7439 , \7440 , \7441 , \7442 ,
         \7443 , \7444 , \7445 , \7446 , \7447 , \7448 , \7449 , \7450 , \7451 , \7452 ,
         \7453 , \7454 , \7455 , \7456 , \7457 , \7458 , \7459 , \7460 , \7461 , \7462 ,
         \7463 , \7464 , \7465 , \7466 , \7467 , \7468 , \7469 , \7470 , \7471 , \7472 ,
         \7473 , \7474 , \7475 , \7476 , \7477 , \7478 , \7479 , \7480 , \7481 , \7482 ,
         \7483 , \7484 , \7485 , \7486 , \7487 , \7488 , \7489 , \7490 , \7491 , \7492 ,
         \7493 , \7494 , \7495 , \7496 , \7497 , \7498 , \7499 , \7500 , \7501 , \7502 ,
         \7503 , \7504 , \7505 , \7506 , \7507 , \7508 , \7509 , \7510 , \7511 , \7512 ,
         \7513 , \7514 , \7515 , \7516 , \7517 , \7518 , \7519 , \7520 , \7521 , \7522 ,
         \7523 , \7524 , \7525 , \7526 , \7527 , \7528 , \7529 , \7530 , \7531 , \7532 ,
         \7533 , \7534 , \7535 , \7536 , \7537 , \7538 , \7539 , \7540 , \7541 , \7542 ,
         \7543 , \7544 , \7545 , \7546 , \7547 , \7548 , \7549 , \7550 , \7551 , \7552 ,
         \7553 , \7554 , \7555 , \7556 , \7557 , \7558 , \7559 , \7560 , \7561 , \7562 ,
         \7563 , \7564 , \7565 , \7566 , \7567 , \7568 , \7569 , \7570 , \7571 , \7572 ,
         \7573 , \7574 , \7575 , \7576 , \7577 , \7578 , \7579 , \7580 , \7581 , \7582 ,
         \7583 , \7584 , \7585 , \7586 , \7587 , \7588 , \7589 , \7590 , \7591 , \7592 ,
         \7593 , \7594 , \7595 , \7596 , \7597 , \7598 , \7599 , \7600 , \7601 , \7602 ,
         \7603 , \7604 , \7605 , \7606 , \7607 , \7608 , \7609 , \7610 , \7611 , \7612 ,
         \7613 , \7614 , \7615 , \7616 , \7617 , \7618 , \7619 , \7620 , \7621 , \7622 ,
         \7623 , \7624 , \7625 , \7626 , \7627 , \7628 , \7629 , \7630 , \7631 , \7632 ,
         \7633 , \7634 , \7635 , \7636 , \7637 , \7638 , \7639 , \7640 , \7641 , \7642 ,
         \7643 , \7644 , \7645 , \7646 , \7647 , \7648 , \7649 , \7650 , \7651 , \7652 ,
         \7653 , \7654 , \7655 , \7656 , \7657 , \7658 , \7659 , \7660 , \7661 , \7662 ,
         \7663 , \7664 , \7665 , \7666 , \7667 , \7668 , \7669 , \7670 , \7671 , \7672 ,
         \7673 , \7674 , \7675 , \7676 , \7677 , \7678 , \7679 , \7680 , \7681 , \7682 ,
         \7683 , \7684 , \7685 , \7686 , \7687 , \7688 , \7689 , \7690 , \7691 , \7692 ,
         \7693 , \7694 , \7695 , \7696 , \7697 , \7698 , \7699 , \7700 , \7701 , \7702 ,
         \7703 , \7704 , \7705 , \7706 , \7707 , \7708 , \7709 , \7710 , \7711 , \7712 ,
         \7713 , \7714 , \7715 , \7716 , \7717 , \7718 , \7719 , \7720 , \7721 , \7722 ,
         \7723 , \7724 , \7725 , \7726 , \7727 , \7728 , \7729 , \7730 , \7731 , \7732 ,
         \7733 , \7734 , \7735 , \7736 , \7737 , \7738 , \7739 , \7740 , \7741 , \7742 ,
         \7743 , \7744 , \7745 , \7746 , \7747 , \7748 , \7749 , \7750 , \7751 , \7752 ,
         \7753 , \7754 , \7755 , \7756 , \7757 , \7758 , \7759 , \7760 , \7761 , \7762 ,
         \7763 , \7764 , \7765 , \7766 , \7767 , \7768 , \7769 , \7770 , \7771 , \7772 ,
         \7773 , \7774 , \7775 , \7776 , \7777 , \7778 , \7779 , \7780 , \7781 , \7782 ,
         \7783 , \7784 , \7785 , \7786 , \7787 , \7788 , \7789 , \7790 , \7791 , \7792 ,
         \7793 , \7794 , \7795 , \7796 , \7797 , \7798 , \7799 , \7800 , \7801 , \7802 ,
         \7803 , \7804 , \7805 , \7806 , \7807 , \7808 , \7809 , \7810 , \7811 , \7812 ,
         \7813 , \7814 , \7815 , \7816 , \7817 , \7818 , \7819 , \7820 , \7821 , \7822 ,
         \7823 , \7824 , \7825 , \7826 , \7827 , \7828 , \7829 , \7830 , \7831 , \7832 ,
         \7833 , \7834 , \7835 , \7836 , \7837 , \7838 , \7839 , \7840 , \7841 , \7842 ,
         \7843 , \7844 , \7845 , \7846 , \7847 , \7848 , \7849 , \7850 , \7851 , \7852 ,
         \7853 , \7854 , \7855 , \7856 , \7857 , \7858 , \7859 , \7860 , \7861 , \7862 ,
         \7863 , \7864 , \7865 , \7866 , \7867 , \7868 , \7869 , \7870 , \7871 , \7872 ,
         \7873 , \7874 , \7875 , \7876 , \7877 , \7878 , \7879 , \7880 , \7881 , \7882 ,
         \7883 , \7884 , \7885 , \7886 , \7887 , \7888 , \7889 , \7890 , \7891 , \7892 ,
         \7893 , \7894 , \7895 , \7896 , \7897 , \7898 , \7899 , \7900 , \7901 , \7902 ,
         \7903 , \7904 , \7905 , \7906 , \7907 , \7908 , \7909 , \7910 , \7911 , \7912 ,
         \7913 , \7914 , \7915 , \7916 , \7917 , \7918 , \7919 , \7920 , \7921 , \7922 ,
         \7923 , \7924 , \7925 , \7926 , \7927 , \7928 , \7929 , \7930 , \7931 , \7932 ,
         \7933 , \7934 , \7935 , \7936 , \7937 , \7938 , \7939 , \7940 , \7941 , \7942 ,
         \7943 , \7944 , \7945 , \7946 , \7947 , \7948 , \7949 , \7950 , \7951 , \7952 ,
         \7953 , \7954 , \7955 , \7956 , \7957 , \7958 , \7959 , \7960 , \7961 , \7962 ,
         \7963 , \7964 , \7965 , \7966 , \7967 , \7968 , \7969 , \7970 , \7971 , \7972 ,
         \7973 , \7974 , \7975 , \7976 , \7977 , \7978 , \7979 , \7980 , \7981 , \7982 ,
         \7983 , \7984 , \7985 , \7986 , \7987 , \7988 , \7989 , \7990 , \7991 , \7992 ,
         \7993 , \7994 , \7995 , \7996 , \7997 , \7998 , \7999 , \8000 , \8001 , \8002 ,
         \8003 , \8004 , \8005 , \8006 , \8007 , \8008 , \8009 , \8010 , \8011 , \8012 ,
         \8013 , \8014 , \8015 , \8016 , \8017 , \8018 , \8019 , \8020 , \8021 , \8022 ,
         \8023 , \8024 , \8025 , \8026 , \8027 , \8028 , \8029 , \8030 , \8031 , \8032 ,
         \8033 , \8034 , \8035 , \8036 , \8037 , \8038 , \8039 , \8040 , \8041 , \8042 ,
         \8043 , \8044 , \8045 , \8046 , \8047 , \8048 , \8049 , \8050 , \8051 , \8052 ,
         \8053 , \8054 , \8055 , \8056 , \8057 , \8058 , \8059 , \8060 , \8061 , \8062 ,
         \8063 , \8064 , \8065 , \8066 , \8067 , \8068 , \8069 , \8070 , \8071 , \8072 ,
         \8073 , \8074 , \8075 , \8076 , \8077 , \8078 , \8079 , \8080 , \8081 , \8082 ,
         \8083 , \8084 , \8085 , \8086 , \8087 , \8088 , \8089 , \8090 , \8091 , \8092 ,
         \8093 , \8094 , \8095 , \8096 , \8097 , \8098 , \8099 , \8100 , \8101 , \8102 ,
         \8103 , \8104 , \8105 , \8106 , \8107 , \8108 , \8109 , \8110 , \8111 , \8112 ,
         \8113 , \8114 , \8115 , \8116 , \8117 , \8118 , \8119 , \8120 , \8121 , \8122 ,
         \8123 , \8124 , \8125 , \8126 , \8127 , \8128 , \8129 , \8130 , \8131 , \8132 ,
         \8133 , \8134 , \8135 , \8136 , \8137 , \8138 , \8139 , \8140 , \8141 , \8142 ,
         \8143 , \8144 , \8145 , \8146 , \8147 , \8148 , \8149 , \8150 , \8151 , \8152 ,
         \8153 , \8154 , \8155 , \8156 , \8157 , \8158 , \8159 , \8160 , \8161 , \8162 ,
         \8163 , \8164 , \8165 , \8166 , \8167 , \8168 , \8169 , \8170 , \8171 , \8172 ,
         \8173 , \8174 , \8175 , \8176 , \8177 , \8178 , \8179 , \8180 , \8181 , \8182 ,
         \8183 , \8184 , \8185 , \8186 , \8187 , \8188 , \8189 , \8190 , \8191 , \8192 ,
         \8193 , \8194 , \8195 , \8196 , \8197 , \8198 , \8199 , \8200 , \8201 , \8202 ,
         \8203 , \8204 , \8205 , \8206 , \8207 , \8208 , \8209 , \8210 , \8211 , \8212 ,
         \8213 , \8214 , \8215 , \8216 , \8217 , \8218 , \8219 , \8220 , \8221 , \8222 ,
         \8223 , \8224 , \8225 , \8226 , \8227 , \8228 , \8229 , \8230 , \8231 , \8232 ,
         \8233 , \8234 , \8235 , \8236 , \8237 , \8238 , \8239 , \8240 , \8241 , \8242 ,
         \8243 , \8244 , \8245 , \8246 , \8247 , \8248 , \8249 , \8250 , \8251 , \8252 ,
         \8253 , \8254 , \8255 , \8256 , \8257 , \8258 , \8259 , \8260 , \8261 , \8262 ,
         \8263 , \8264 , \8265 , \8266 , \8267 , \8268 , \8269 , \8270 , \8271 , \8272 ,
         \8273 , \8274 , \8275 , \8276 , \8277 , \8278 , \8279 , \8280 , \8281 , \8282 ,
         \8283 , \8284 , \8285 , \8286 , \8287 , \8288 , \8289 , \8290 , \8291 , \8292 ,
         \8293 , \8294 , \8295 , \8296 , \8297 , \8298 , \8299 , \8300 , \8301 , \8302 ,
         \8303 , \8304 , \8305 , \8306 , \8307 , \8308 , \8309 , \8310 , \8311 , \8312 ,
         \8313 , \8314 , \8315 , \8316 , \8317 , \8318 , \8319 , \8320 , \8321 , \8322 ,
         \8323 , \8324 , \8325 , \8326 , \8327 , \8328 , \8329 , \8330 , \8331 , \8332 ,
         \8333 , \8334 , \8335 , \8336 , \8337 , \8338 , \8339 , \8340 , \8341 , \8342 ,
         \8343 , \8344 , \8345 , \8346 , \8347 , \8348 , \8349 , \8350 , \8351 , \8352 ,
         \8353 , \8354 , \8355 , \8356 , \8357 , \8358 , \8359 , \8360 , \8361 , \8362 ,
         \8363 , \8364 , \8365 , \8366 , \8367 , \8368 , \8369 , \8370 , \8371 , \8372 ,
         \8373 , \8374 , \8375 , \8376 , \8377 , \8378 , \8379 , \8380 , \8381 , \8382 ,
         \8383 , \8384 , \8385 , \8386 , \8387 , \8388 , \8389 , \8390 , \8391 , \8392 ,
         \8393 , \8394 , \8395 , \8396 , \8397 , \8398 , \8399 , \8400 , \8401 , \8402 ,
         \8403 , \8404 , \8405 , \8406 , \8407 , \8408 , \8409 , \8410 , \8411 , \8412 ,
         \8413 , \8414 , \8415 , \8416 , \8417 , \8418 , \8419 , \8420 , \8421 , \8422 ,
         \8423 , \8424 , \8425 , \8426 , \8427 , \8428 , \8429 , \8430 , \8431 , \8432 ,
         \8433 , \8434 , \8435 , \8436 , \8437 , \8438 , \8439 , \8440 , \8441 , \8442 ,
         \8443 , \8444 , \8445 , \8446 , \8447 , \8448 , \8449 , \8450 , \8451 , \8452 ,
         \8453 , \8454 , \8455 , \8456 , \8457 , \8458 , \8459 , \8460 , \8461 , \8462 ,
         \8463 , \8464 , \8465 , \8466 , \8467 , \8468 , \8469 , \8470 , \8471 , \8472 ,
         \8473 , \8474 , \8475 , \8476 , \8477 , \8478 , \8479 , \8480 , \8481 , \8482 ,
         \8483 , \8484 , \8485 , \8486 , \8487 , \8488 , \8489 , \8490 , \8491 , \8492 ,
         \8493 , \8494 , \8495 , \8496 , \8497 , \8498 , \8499 , \8500 , \8501 , \8502 ,
         \8503 , \8504 , \8505 , \8506 , \8507 , \8508 , \8509 , \8510 , \8511 , \8512 ,
         \8513 , \8514 , \8515 , \8516 , \8517 , \8518 , \8519 , \8520 , \8521 , \8522 ,
         \8523 , \8524 , \8525 , \8526 , \8527 , \8528 , \8529 , \8530 , \8531 , \8532 ,
         \8533 , \8534 , \8535 , \8536 , \8537 , \8538 , \8539 , \8540 , \8541 , \8542 ,
         \8543 , \8544 , \8545 , \8546 , \8547 , \8548 , \8549 , \8550 , \8551 , \8552 ,
         \8553 , \8554 , \8555 , \8556 , \8557 , \8558 , \8559 , \8560 , \8561 , \8562 ,
         \8563 , \8564 , \8565 , \8566 , \8567 , \8568 , \8569 , \8570 , \8571 , \8572 ,
         \8573 , \8574 , \8575 , \8576 , \8577 , \8578 , \8579 , \8580 , \8581 , \8582 ,
         \8583 , \8584 , \8585 , \8586 , \8587 , \8588 , \8589 , \8590 , \8591 , \8592 ,
         \8593 , \8594 , \8595 , \8596 , \8597 , \8598 , \8599 , \8600 , \8601 , \8602 ,
         \8603 , \8604 , \8605 , \8606 , \8607 , \8608 , \8609 , \8610 , \8611 , \8612 ,
         \8613 , \8614 , \8615 , \8616 , \8617 , \8618 , \8619 , \8620 , \8621 , \8622 ,
         \8623 , \8624 , \8625 , \8626 , \8627 , \8628 , \8629 , \8630 , \8631 , \8632 ,
         \8633 , \8634 , \8635 , \8636 , \8637 , \8638 , \8639 , \8640 , \8641 , \8642 ,
         \8643 , \8644 , \8645 , \8646 , \8647 , \8648 , \8649 , \8650 , \8651 , \8652 ,
         \8653 , \8654 , \8655 , \8656 , \8657 , \8658 , \8659 , \8660 , \8661 , \8662 ,
         \8663 , \8664 , \8665 , \8666 , \8667 , \8668 , \8669 , \8670 , \8671 , \8672 ,
         \8673 , \8674 , \8675 , \8676 , \8677 , \8678 , \8679 , \8680 , \8681 , \8682 ,
         \8683 , \8684 , \8685 , \8686 , \8687 , \8688 , \8689 , \8690 , \8691 , \8692 ,
         \8693 , \8694 , \8695 , \8696 , \8697 , \8698 , \8699 , \8700 , \8701 , \8702 ,
         \8703 , \8704 , \8705 , \8706 , \8707 , \8708 , \8709 , \8710 , \8711 , \8712 ,
         \8713 , \8714 , \8715 , \8716 , \8717 , \8718 , \8719 , \8720 , \8721 , \8722 ,
         \8723 , \8724 , \8725 , \8726 , \8727 , \8728 , \8729 , \8730 , \8731 , \8732 ,
         \8733 , \8734 , \8735 , \8736 , \8737 , \8738 , \8739 , \8740 , \8741 , \8742 ,
         \8743 , \8744 , \8745 , \8746 , \8747 , \8748 , \8749 , \8750 , \8751 , \8752 ,
         \8753 , \8754 , \8755 , \8756 , \8757 , \8758 , \8759 , \8760 , \8761 , \8762 ,
         \8763 , \8764 , \8765 , \8766 , \8767 , \8768 , \8769 , \8770 , \8771 , \8772 ,
         \8773 , \8774 , \8775 , \8776 , \8777 , \8778 , \8779 , \8780 , \8781 , \8782 ,
         \8783 , \8784 , \8785 , \8786 , \8787 , \8788 , \8789 , \8790 , \8791 , \8792 ,
         \8793 , \8794 , \8795 , \8796 , \8797 , \8798 , \8799 , \8800 , \8801 , \8802 ,
         \8803 , \8804 , \8805 , \8806 , \8807 , \8808 , \8809 , \8810 , \8811 , \8812 ,
         \8813 , \8814 , \8815 , \8816 , \8817 , \8818 , \8819 , \8820 , \8821 , \8822 ,
         \8823 , \8824 , \8825 , \8826 , \8827 , \8828 , \8829 , \8830 , \8831 , \8832 ,
         \8833 , \8834 , \8835 , \8836 , \8837 , \8838 , \8839 , \8840 , \8841 , \8842 ,
         \8843 , \8844 , \8845 , \8846 , \8847 , \8848 , \8849 , \8850 , \8851 , \8852 ,
         \8853 , \8854 , \8855 , \8856 , \8857 , \8858 , \8859 , \8860 , \8861 , \8862 ,
         \8863 , \8864 , \8865 , \8866 , \8867 , \8868 , \8869 , \8870 , \8871 , \8872 ,
         \8873 , \8874 , \8875 , \8876 , \8877 , \8878 , \8879 , \8880 , \8881 , \8882 ,
         \8883 , \8884 , \8885 , \8886 , \8887 , \8888 , \8889 , \8890 , \8891 , \8892 ,
         \8893 , \8894 , \8895 , \8896 , \8897 , \8898 , \8899 , \8900 , \8901 , \8902 ,
         \8903 , \8904 , \8905 , \8906 , \8907 , \8908 , \8909 , \8910 , \8911 , \8912 ,
         \8913 , \8914 , \8915 , \8916 , \8917 , \8918 , \8919 , \8920 , \8921 , \8922 ,
         \8923 , \8924 , \8925 , \8926 , \8927 , \8928 , \8929 , \8930 , \8931 , \8932 ,
         \8933 , \8934 , \8935 , \8936 , \8937 , \8938 , \8939 , \8940 , \8941 , \8942 ,
         \8943 , \8944 , \8945 , \8946 , \8947 , \8948 , \8949 , \8950 , \8951 , \8952 ,
         \8953 , \8954 , \8955 , \8956 , \8957 , \8958 , \8959 , \8960 , \8961 , \8962 ,
         \8963 , \8964 , \8965 , \8966 , \8967 , \8968 , \8969 , \8970 , \8971 , \8972 ,
         \8973 , \8974 , \8975 , \8976 , \8977 , \8978 , \8979 , \8980 , \8981 , \8982 ,
         \8983 , \8984 , \8985 , \8986 , \8987 , \8988 , \8989 , \8990 , \8991 , \8992 ,
         \8993 , \8994 , \8995 , \8996 , \8997 , \8998 , \8999 , \9000 , \9001 , \9002 ,
         \9003 , \9004 , \9005 , \9006 , \9007 , \9008 , \9009 , \9010 , \9011 , \9012 ,
         \9013 , \9014 , \9015 , \9016 , \9017 , \9018 , \9019 , \9020 , \9021 , \9022 ,
         \9023 , \9024 , \9025 , \9026 , \9027 , \9028 , \9029 , \9030 , \9031 , \9032 ,
         \9033 , \9034 , \9035 , \9036 , \9037 , \9038 , \9039 , \9040 , \9041 , \9042 ,
         \9043 , \9044 , \9045 , \9046 , \9047 , \9048 , \9049 , \9050 , \9051 , \9052 ,
         \9053 , \9054 , \9055 , \9056 , \9057 , \9058 , \9059 , \9060 , \9061 , \9062 ,
         \9063 , \9064 , \9065 , \9066 , \9067 , \9068 , \9069 , \9070 , \9071 , \9072 ,
         \9073 , \9074 , \9075 , \9076 , \9077 , \9078 , \9079 , \9080 , \9081 , \9082 ,
         \9083 , \9084 , \9085 , \9086 , \9087 , \9088 , \9089 , \9090 , \9091 , \9092 ,
         \9093 , \9094 , \9095 , \9096 , \9097 , \9098 , \9099 , \9100 , \9101 , \9102 ,
         \9103 , \9104 , \9105 , \9106 , \9107 , \9108 , \9109 , \9110 , \9111 , \9112 ,
         \9113 , \9114 , \9115 , \9116 , \9117 , \9118 , \9119 , \9120 , \9121 , \9122 ,
         \9123 , \9124 , \9125 , \9126 , \9127 , \9128 , \9129 , \9130 , \9131 , \9132 ,
         \9133 , \9134 , \9135 , \9136 , \9137 , \9138 , \9139 , \9140 , \9141 , \9142 ,
         \9143 , \9144 , \9145 , \9146 , \9147 , \9148 , \9149 , \9150 , \9151 , \9152 ,
         \9153 , \9154 , \9155 , \9156 , \9157 , \9158 , \9159 , \9160 , \9161 , \9162 ,
         \9163 , \9164 , \9165 , \9166 , \9167 , \9168 , \9169 , \9170 , \9171 , \9172 ,
         \9173 , \9174 , \9175 , \9176 , \9177 , \9178 , \9179 , \9180 , \9181 , \9182 ,
         \9183 , \9184 , \9185 , \9186 , \9187 , \9188 , \9189 , \9190 , \9191 , \9192 ,
         \9193 , \9194 , \9195 , \9196 , \9197 , \9198 , \9199 , \9200 , \9201 , \9202 ,
         \9203 , \9204 , \9205 , \9206 , \9207 , \9208 , \9209 , \9210 , \9211 , \9212 ,
         \9213 , \9214 , \9215 , \9216 , \9217 , \9218 , \9219 , \9220 , \9221 , \9222 ,
         \9223 , \9224 , \9225 , \9226 , \9227 , \9228 , \9229 , \9230 , \9231 , \9232 ,
         \9233 , \9234 , \9235 , \9236 , \9237 , \9238 , \9239 , \9240 , \9241 , \9242 ,
         \9243 , \9244 , \9245 , \9246 , \9247 , \9248 , \9249 , \9250 , \9251 , \9252 ,
         \9253 , \9254 , \9255 , \9256 , \9257 , \9258 , \9259 , \9260 , \9261 , \9262 ,
         \9263 , \9264 , \9265 , \9266 , \9267 , \9268 , \9269 , \9270 , \9271 , \9272 ,
         \9273 , \9274 , \9275 , \9276 , \9277 , \9278 , \9279 , \9280 , \9281 , \9282 ,
         \9283 , \9284 , \9285 , \9286 , \9287 , \9288 , \9289 , \9290 , \9291 , \9292 ,
         \9293 , \9294 , \9295 , \9296 , \9297 , \9298 , \9299 , \9300 , \9301 , \9302 ,
         \9303 , \9304 , \9305 , \9306 , \9307 , \9308 , \9309 , \9310 , \9311 , \9312 ,
         \9313 , \9314 , \9315 , \9316 , \9317 , \9318 , \9319 , \9320 , \9321 , \9322 ,
         \9323 , \9324 , \9325 , \9326 , \9327 , \9328 , \9329 , \9330 , \9331 , \9332 ,
         \9333 , \9334 , \9335 , \9336 , \9337 , \9338 , \9339 , \9340 , \9341 , \9342 ,
         \9343 , \9344 , \9345 , \9346 , \9347 , \9348 , \9349 , \9350 , \9351 , \9352 ,
         \9353 , \9354 , \9355 , \9356 , \9357 , \9358 , \9359 , \9360 , \9361 , \9362 ,
         \9363 , \9364 , \9365 , \9366 , \9367 , \9368 , \9369 , \9370 , \9371 , \9372 ,
         \9373 , \9374 , \9375 , \9376 , \9377 , \9378 , \9379 , \9380 , \9381 , \9382 ,
         \9383 , \9384 , \9385 , \9386 , \9387 , \9388 , \9389 , \9390 , \9391 , \9392 ,
         \9393 , \9394 , \9395 , \9396 , \9397 , \9398 , \9399 , \9400 , \9401 , \9402 ,
         \9403 , \9404 , \9405 , \9406 , \9407 , \9408 , \9409 , \9410 , \9411 , \9412 ,
         \9413 , \9414 , \9415 , \9416 , \9417 , \9418 , \9419 , \9420 , \9421 , \9422 ,
         \9423 , \9424 , \9425 , \9426 , \9427 , \9428 , \9429 , \9430 , \9431 , \9432 ,
         \9433 , \9434 , \9435 , \9436 , \9437 , \9438 , \9439 , \9440 , \9441 , \9442 ,
         \9443 , \9444 , \9445 , \9446 , \9447 , \9448 , \9449 , \9450 , \9451 , \9452 ,
         \9453 , \9454 , \9455 , \9456 , \9457 , \9458 , \9459 , \9460 , \9461 , \9462 ,
         \9463 , \9464 , \9465 , \9466 , \9467 , \9468 , \9469 , \9470 , \9471 , \9472 ,
         \9473 , \9474 , \9475 , \9476 , \9477 , \9478 , \9479 , \9480 , \9481 , \9482 ,
         \9483 , \9484 , \9485 , \9486 , \9487 , \9488 , \9489 , \9490 , \9491 , \9492 ,
         \9493 , \9494 , \9495 , \9496 , \9497 , \9498 , \9499 , \9500 , \9501 , \9502 ,
         \9503 , \9504 , \9505 , \9506 , \9507 , \9508 , \9509 , \9510 , \9511 , \9512 ,
         \9513 , \9514 , \9515 , \9516 , \9517 , \9518 , \9519 , \9520 , \9521 , \9522 ,
         \9523 , \9524 , \9525 , \9526 , \9527 , \9528 , \9529 , \9530 , \9531 , \9532 ,
         \9533 , \9534 , \9535 , \9536 , \9537 , \9538 , \9539 , \9540 , \9541 , \9542 ,
         \9543 , \9544 , \9545 , \9546 , \9547 , \9548 , \9549 , \9550 , \9551 , \9552 ,
         \9553 , \9554 , \9555 , \9556 , \9557 , \9558 , \9559 , \9560 , \9561 , \9562 ,
         \9563 , \9564 , \9565 , \9566 , \9567 , \9568 , \9569 , \9570 , \9571 , \9572 ,
         \9573 , \9574 , \9575 , \9576 , \9577 , \9578 , \9579 , \9580 , \9581 , \9582 ,
         \9583 , \9584 , \9585 , \9586 , \9587 , \9588 , \9589 , \9590 , \9591 , \9592 ,
         \9593 , \9594 , \9595 , \9596 , \9597 , \9598 , \9599 , \9600 , \9601 , \9602 ,
         \9603 , \9604 , \9605 , \9606 , \9607 , \9608 , \9609 , \9610 , \9611 , \9612 ,
         \9613 , \9614 , \9615 , \9616 , \9617 , \9618 , \9619 , \9620 , \9621 , \9622 ,
         \9623 , \9624 , \9625 , \9626 , \9627 , \9628 , \9629 , \9630 , \9631 , \9632 ,
         \9633 , \9634 , \9635 , \9636 , \9637 , \9638 , \9639 , \9640 , \9641 , \9642 ,
         \9643 , \9644 , \9645 , \9646 , \9647 , \9648 , \9649 , \9650 , \9651 , \9652 ,
         \9653 , \9654 , \9655 , \9656 , \9657 , \9658 , \9659 , \9660 , \9661 , \9662 ,
         \9663 , \9664 , \9665 , \9666 , \9667 , \9668 , \9669 , \9670 , \9671 , \9672 ,
         \9673 , \9674 , \9675 , \9676 , \9677 , \9678 , \9679 , \9680 , \9681 , \9682 ,
         \9683 , \9684 , \9685 , \9686 , \9687 , \9688 , \9689 , \9690 , \9691 , \9692 ,
         \9693 , \9694 , \9695 , \9696 , \9697 , \9698 , \9699 , \9700 , \9701 , \9702 ,
         \9703 , \9704 , \9705 , \9706 , \9707 , \9708 , \9709 , \9710 , \9711 , \9712 ,
         \9713 , \9714 , \9715 , \9716 , \9717 , \9718 , \9719 , \9720 , \9721 , \9722 ,
         \9723 , \9724 , \9725 , \9726 , \9727 , \9728 , \9729 , \9730 , \9731 , \9732 ,
         \9733 , \9734 , \9735 , \9736 , \9737 , \9738 , \9739 , \9740 , \9741 , \9742 ,
         \9743 , \9744 , \9745 , \9746 , \9747 , \9748 , \9749 , \9750 , \9751 , \9752 ,
         \9753 , \9754 , \9755 , \9756 , \9757 , \9758 , \9759 , \9760 , \9761 , \9762 ,
         \9763 , \9764 , \9765 , \9766 , \9767 , \9768 , \9769 , \9770 , \9771 , \9772 ,
         \9773 , \9774 , \9775 , \9776 , \9777 , \9778 , \9779 , \9780 , \9781 , \9782 ,
         \9783 , \9784 , \9785 , \9786 , \9787 , \9788 , \9789 , \9790 , \9791 , \9792 ,
         \9793 , \9794 , \9795 , \9796 , \9797 , \9798 , \9799 , \9800 , \9801 , \9802 ,
         \9803 , \9804 , \9805 , \9806 , \9807 , \9808 , \9809 , \9810 , \9811 , \9812 ,
         \9813 , \9814 , \9815 , \9816 , \9817 , \9818 , \9819 , \9820 , \9821 , \9822 ,
         \9823 , \9824 , \9825 , \9826 , \9827 , \9828 , \9829 , \9830 , \9831 , \9832 ,
         \9833 , \9834 , \9835 , \9836 , \9837 , \9838 , \9839 , \9840 , \9841 , \9842 ,
         \9843 , \9844 , \9845 , \9846 , \9847 , \9848 , \9849 , \9850 , \9851 , \9852 ,
         \9853 , \9854 , \9855 , \9856 , \9857 , \9858 , \9859 , \9860 , \9861 , \9862 ,
         \9863 , \9864 , \9865 , \9866 , \9867 , \9868 , \9869 , \9870 , \9871 , \9872 ,
         \9873 , \9874 , \9875 , \9876 , \9877 , \9878 , \9879 , \9880 , \9881 , \9882 ,
         \9883 , \9884 , \9885 , \9886 , \9887 , \9888 , \9889 , \9890 , \9891 , \9892 ,
         \9893 , \9894 , \9895 , \9896 , \9897 , \9898 , \9899 , \9900 , \9901 , \9902 ,
         \9903 , \9904 , \9905 , \9906 , \9907 , \9908 , \9909 , \9910 , \9911 , \9912 ,
         \9913 , \9914 , \9915 , \9916 , \9917 , \9918 , \9919 , \9920 , \9921 , \9922 ,
         \9923 , \9924 , \9925 , \9926 , \9927 , \9928 , \9929 , \9930 , \9931 , \9932 ,
         \9933 , \9934 , \9935 , \9936 , \9937 , \9938 , \9939 , \9940 , \9941 , \9942 ,
         \9943 , \9944 , \9945 , \9946 , \9947 , \9948 , \9949 , \9950 , \9951 , \9952 ,
         \9953 , \9954 , \9955 , \9956 , \9957 , \9958 , \9959 , \9960 , \9961 , \9962 ,
         \9963 , \9964 , \9965 , \9966 , \9967 , \9968 , \9969 , \9970 , \9971 , \9972 ,
         \9973 , \9974 , \9975 , \9976 , \9977 , \9978 , \9979 , \9980 , \9981 , \9982 ,
         \9983 , \9984 , \9985 , \9986 , \9987 , \9988 , \9989 , \9990 , \9991 , \9992 ,
         \9993 , \9994 , \9995 , \9996 , \9997 , \9998 , \9999 , \10000 , \10001 , \10002 ,
         \10003 , \10004 , \10005 , \10006 , \10007 , \10008 , \10009 , \10010 , \10011 , \10012 ,
         \10013 , \10014 , \10015 , \10016 , \10017 , \10018 , \10019 , \10020 , \10021 , \10022 ,
         \10023 , \10024 , \10025 , \10026 , \10027 , \10028 , \10029 , \10030 , \10031 , \10032 ,
         \10033 , \10034 , \10035 , \10036 , \10037 , \10038 , \10039 , \10040 , \10041 , \10042 ,
         \10043 , \10044 , \10045 , \10046 , \10047 , \10048 , \10049 , \10050 , \10051 , \10052 ,
         \10053 , \10054 , \10055 , \10056 , \10057 , \10058 , \10059 , \10060 , \10061 , \10062 ,
         \10063 , \10064 , \10065 , \10066 , \10067 , \10068 , \10069 , \10070 , \10071 , \10072 ,
         \10073 , \10074 , \10075 , \10076 , \10077 , \10078 , \10079 , \10080 , \10081 , \10082 ,
         \10083 , \10084 , \10085 , \10086 , \10087 , \10088 , \10089 , \10090 , \10091 , \10092 ,
         \10093 , \10094 , \10095 , \10096 , \10097 , \10098 , \10099 , \10100 , \10101 , \10102 ,
         \10103 , \10104 , \10105 , \10106 , \10107 , \10108 , \10109 , \10110 , \10111 , \10112 ,
         \10113 , \10114 , \10115 , \10116 , \10117 , \10118 , \10119 , \10120 , \10121 , \10122 ,
         \10123 , \10124 , \10125 , \10126 , \10127 , \10128 , \10129 , \10130 , \10131 , \10132 ,
         \10133 , \10134 , \10135 , \10136 , \10137 , \10138 , \10139 , \10140 , \10141 , \10142 ,
         \10143 , \10144 , \10145 , \10146 , \10147 , \10148 , \10149 , \10150 , \10151 , \10152 ,
         \10153 , \10154 , \10155 , \10156 , \10157 , \10158 , \10159 , \10160 , \10161 , \10162 ,
         \10163 , \10164 , \10165 , \10166 , \10167 , \10168 , \10169 , \10170 , \10171 , \10172 ,
         \10173 , \10174 , \10175 , \10176 , \10177 , \10178 , \10179 , \10180 , \10181 , \10182 ,
         \10183 , \10184 , \10185 , \10186 , \10187 , \10188 , \10189 , \10190 , \10191 , \10192 ,
         \10193 , \10194 , \10195 , \10196 , \10197 , \10198 , \10199 , \10200 , \10201 , \10202 ,
         \10203 , \10204 , \10205 , \10206 , \10207 , \10208 , \10209 , \10210 , \10211 , \10212 ,
         \10213 , \10214 , \10215 , \10216 , \10217 , \10218 , \10219 , \10220 , \10221 , \10222 ,
         \10223 , \10224 , \10225 , \10226 , \10227 , \10228 , \10229 , \10230 , \10231 , \10232 ,
         \10233 , \10234 , \10235 , \10236 , \10237 , \10238 , \10239 , \10240 , \10241 , \10242 ,
         \10243 , \10244 , \10245 , \10246 , \10247 , \10248 , \10249 , \10250 , \10251 , \10252 ,
         \10253 , \10254 , \10255 , \10256 , \10257 , \10258 , \10259 , \10260 , \10261 , \10262 ,
         \10263 , \10264 , \10265 , \10266 , \10267 , \10268 , \10269 , \10270 , \10271 , \10272 ,
         \10273 , \10274 , \10275 , \10276 , \10277 , \10278 , \10279 , \10280 , \10281 , \10282 ,
         \10283 , \10284 , \10285 , \10286 , \10287 , \10288 , \10289 , \10290 , \10291 , \10292 ,
         \10293 , \10294 , \10295 , \10296 , \10297 , \10298 , \10299 , \10300 , \10301 , \10302 ,
         \10303 , \10304 , \10305 , \10306 , \10307 , \10308 , \10309 , \10310 , \10311 , \10312 ,
         \10313 , \10314 , \10315 , \10316 , \10317 , \10318 , \10319 , \10320 , \10321 , \10322 ,
         \10323 , \10324 , \10325 , \10326 , \10327 , \10328 , \10329 , \10330 , \10331 , \10332 ,
         \10333 , \10334 , \10335 , \10336 , \10337 , \10338 , \10339 , \10340 , \10341 , \10342 ,
         \10343 , \10344 , \10345 , \10346 , \10347 , \10348 , \10349 , \10350 , \10351 , \10352 ,
         \10353 , \10354 , \10355 , \10356 , \10357 , \10358 , \10359 , \10360 , \10361 , \10362 ,
         \10363 , \10364 , \10365 , \10366 , \10367 , \10368 , \10369 , \10370 , \10371 , \10372 ,
         \10373 , \10374 , \10375 , \10376 , \10377 , \10378 , \10379 , \10380 , \10381 , \10382 ,
         \10383 , \10384 , \10385 , \10386 , \10387 , \10388 , \10389 , \10390 , \10391 , \10392 ,
         \10393 , \10394 , \10395 , \10396 , \10397 , \10398 , \10399 , \10400 , \10401 , \10402 ,
         \10403 , \10404 , \10405 , \10406 , \10407 , \10408 , \10409 , \10410 , \10411 , \10412 ,
         \10413 , \10414 , \10415 , \10416 , \10417 , \10418 , \10419 , \10420 , \10421 , \10422 ,
         \10423 , \10424 , \10425 , \10426 , \10427 , \10428 , \10429 , \10430 , \10431 , \10432 ,
         \10433 , \10434 , \10435 , \10436 , \10437 , \10438 , \10439 , \10440 , \10441 , \10442 ,
         \10443 , \10444 , \10445 , \10446 , \10447 , \10448 , \10449 , \10450 , \10451 , \10452 ,
         \10453 , \10454 , \10455 , \10456 , \10457 , \10458 , \10459 , \10460 , \10461 , \10462 ,
         \10463 , \10464 , \10465 , \10466 , \10467 , \10468 , \10469 , \10470 , \10471 , \10472 ,
         \10473 , \10474 , \10475 , \10476 , \10477 , \10478 , \10479 , \10480 , \10481 , \10482 ,
         \10483 , \10484 , \10485 , \10486 , \10487 , \10488 , \10489 , \10490 , \10491 , \10492 ,
         \10493 , \10494 , \10495 , \10496 , \10497 , \10498 , \10499 , \10500 , \10501 , \10502 ,
         \10503 , \10504 , \10505 , \10506 , \10507 , \10508 , \10509 , \10510 , \10511 , \10512 ,
         \10513 , \10514 , \10515 , \10516 , \10517 , \10518 , \10519 , \10520 , \10521 , \10522 ,
         \10523 , \10524 , \10525 , \10526 , \10527 , \10528 , \10529 , \10530 , \10531 , \10532 ,
         \10533 , \10534 , \10535 , \10536 , \10537 , \10538 , \10539 , \10540 , \10541 , \10542 ,
         \10543 , \10544 , \10545 , \10546 , \10547 , \10548 , \10549 , \10550 , \10551 , \10552 ,
         \10553 , \10554 , \10555 , \10556 , \10557 , \10558 , \10559 , \10560 , \10561 , \10562 ,
         \10563 , \10564 , \10565 , \10566 , \10567 , \10568 , \10569 , \10570 , \10571 , \10572 ,
         \10573 , \10574 , \10575 , \10576 , \10577 , \10578 , \10579 , \10580 , \10581 , \10582 ,
         \10583 , \10584 , \10585 , \10586 , \10587 , \10588 , \10589 , \10590 , \10591 , \10592 ,
         \10593 , \10594 , \10595 , \10596 , \10597 , \10598 , \10599 , \10600 , \10601 , \10602 ,
         \10603 , \10604 , \10605 , \10606 , \10607 , \10608 , \10609 , \10610 , \10611 , \10612 ,
         \10613 , \10614 , \10615 , \10616 , \10617 , \10618 , \10619 , \10620 , \10621 , \10622 ,
         \10623 , \10624 , \10625 , \10626 , \10627 , \10628 , \10629 , \10630 , \10631 , \10632 ,
         \10633 , \10634 , \10635 , \10636 , \10637 , \10638 , \10639 , \10640 , \10641 , \10642 ,
         \10643 , \10644 , \10645 , \10646 , \10647 , \10648 , \10649 , \10650 , \10651 , \10652 ,
         \10653 , \10654 , \10655 , \10656 , \10657 , \10658 , \10659 , \10660 , \10661 , \10662 ,
         \10663 , \10664 , \10665 , \10666 , \10667 , \10668 , \10669 , \10670 , \10671 , \10672 ,
         \10673 , \10674 , \10675 , \10676 , \10677 , \10678 , \10679 , \10680 , \10681 , \10682 ,
         \10683 , \10684 , \10685 , \10686 , \10687 , \10688 , \10689 , \10690 , \10691 , \10692 ,
         \10693 , \10694 , \10695 , \10696 , \10697 , \10698 , \10699 , \10700 , \10701 , \10702 ,
         \10703 , \10704 , \10705 , \10706 , \10707 , \10708 , \10709 , \10710 , \10711 , \10712 ,
         \10713 , \10714 , \10715 , \10716 , \10717 , \10718 , \10719 , \10720 , \10721 , \10722 ,
         \10723 , \10724 , \10725 , \10726 , \10727 , \10728 , \10729 , \10730 , \10731 , \10732 ,
         \10733 , \10734 , \10735 , \10736 , \10737 , \10738 , \10739 , \10740 , \10741 , \10742 ,
         \10743 , \10744 , \10745 , \10746 , \10747 , \10748 , \10749 , \10750 , \10751 , \10752 ,
         \10753 , \10754 , \10755 , \10756 , \10757 , \10758 , \10759 , \10760 , \10761 , \10762 ,
         \10763 , \10764 , \10765 , \10766 , \10767 , \10768 , \10769 , \10770 , \10771 , \10772 ,
         \10773 , \10774 , \10775 , \10776 , \10777 , \10778 , \10779 , \10780 , \10781 , \10782 ,
         \10783 , \10784 , \10785 , \10786 , \10787 , \10788 , \10789 , \10790 , \10791 , \10792 ,
         \10793 , \10794 , \10795 , \10796 , \10797 , \10798 , \10799 , \10800 , \10801 , \10802 ,
         \10803 , \10804 , \10805 , \10806 , \10807 , \10808 , \10809 , \10810 , \10811 , \10812 ,
         \10813 , \10814 , \10815 , \10816 , \10817 , \10818 , \10819 , \10820 , \10821 , \10822 ,
         \10823 , \10824 , \10825 , \10826 , \10827 , \10828 , \10829 , \10830 , \10831 , \10832 ,
         \10833 , \10834 , \10835 , \10836 , \10837 , \10838 , \10839 , \10840 , \10841 , \10842 ,
         \10843 , \10844 , \10845 , \10846 , \10847 , \10848 , \10849 , \10850 , \10851 , \10852 ,
         \10853 , \10854 , \10855 , \10856 , \10857 , \10858 , \10859 , \10860 , \10861 , \10862 ,
         \10863 , \10864 , \10865 , \10866 , \10867 , \10868 , \10869 , \10870 , \10871 , \10872 ,
         \10873 , \10874 , \10875 , \10876 , \10877 , \10878 , \10879 , \10880 , \10881 , \10882 ,
         \10883 , \10884 , \10885 , \10886 , \10887 , \10888 , \10889 , \10890 , \10891 , \10892 ,
         \10893 , \10894 , \10895 , \10896 , \10897 , \10898 , \10899 , \10900 , \10901 , \10902 ,
         \10903 , \10904 , \10905 , \10906 , \10907 , \10908 , \10909 , \10910 , \10911 , \10912 ,
         \10913 , \10914 , \10915 , \10916 , \10917 , \10918 , \10919 , \10920 , \10921 , \10922 ,
         \10923 , \10924 , \10925 , \10926 , \10927 , \10928 , \10929 , \10930 , \10931 , \10932 ,
         \10933 , \10934 , \10935 , \10936 , \10937 , \10938 , \10939 , \10940 , \10941 , \10942 ,
         \10943 , \10944 , \10945 , \10946 , \10947 , \10948 , \10949 , \10950 , \10951 , \10952 ,
         \10953 , \10954 , \10955 , \10956 , \10957 , \10958 , \10959 , \10960 , \10961 , \10962 ,
         \10963 , \10964 , \10965 , \10966 , \10967 , \10968 , \10969 , \10970 , \10971 , \10972 ,
         \10973 , \10974 , \10975 , \10976 , \10977 , \10978 , \10979 , \10980 , \10981 , \10982 ,
         \10983 , \10984 , \10985 , \10986 , \10987 , \10988 , \10989 , \10990 , \10991 , \10992 ,
         \10993 , \10994 , \10995 , \10996 , \10997 , \10998 , \10999 , \11000 , \11001 , \11002 ,
         \11003 , \11004 , \11005 , \11006 , \11007 , \11008 , \11009 , \11010 , \11011 , \11012 ,
         \11013 , \11014 , \11015 , \11016 , \11017 , \11018 , \11019 , \11020 , \11021 , \11022 ,
         \11023 , \11024 , \11025 , \11026 , \11027 , \11028 , \11029 , \11030 , \11031 , \11032 ,
         \11033 , \11034 , \11035 , \11036 , \11037 , \11038 , \11039 , \11040 , \11041 , \11042 ,
         \11043 , \11044 , \11045 , \11046 , \11047 , \11048 , \11049 , \11050 , \11051 , \11052 ,
         \11053 , \11054 , \11055 , \11056 , \11057 , \11058 , \11059 , \11060 , \11061 , \11062 ,
         \11063 , \11064 , \11065 , \11066 , \11067 , \11068 , \11069 , \11070 , \11071 , \11072 ,
         \11073 , \11074 , \11075 , \11076 , \11077 , \11078 , \11079 , \11080 , \11081 , \11082 ,
         \11083 , \11084 , \11085 , \11086 , \11087 , \11088 , \11089 , \11090 , \11091 , \11092 ,
         \11093 , \11094 , \11095 , \11096 , \11097 , \11098 , \11099 , \11100 , \11101 , \11102 ,
         \11103 , \11104 , \11105 , \11106 , \11107 , \11108 , \11109 , \11110 , \11111 , \11112 ,
         \11113 , \11114 , \11115 , \11116 , \11117 , \11118 , \11119 , \11120 , \11121 , \11122 ,
         \11123 , \11124 , \11125 , \11126 , \11127 , \11128 , \11129 , \11130 , \11131 , \11132 ,
         \11133 , \11134 , \11135 , \11136 , \11137 , \11138 , \11139 , \11140 , \11141 , \11142 ,
         \11143 , \11144 , \11145 , \11146 , \11147 , \11148 , \11149 , \11150 , \11151 , \11152 ,
         \11153 , \11154 , \11155 , \11156 , \11157 , \11158 , \11159 , \11160 , \11161 , \11162 ,
         \11163 , \11164 , \11165 , \11166 , \11167 , \11168 , \11169 , \11170 , \11171 , \11172 ,
         \11173 , \11174 , \11175 , \11176 , \11177 , \11178 , \11179 , \11180 , \11181 , \11182 ,
         \11183 , \11184 , \11185 , \11186 , \11187 , \11188 , \11189 , \11190 , \11191 , \11192 ,
         \11193 , \11194 , \11195 , \11196 , \11197 , \11198 , \11199 , \11200 , \11201 , \11202 ,
         \11203 , \11204 , \11205 , \11206 , \11207 , \11208 , \11209 , \11210 , \11211 , \11212 ,
         \11213 , \11214 , \11215 , \11216 , \11217 , \11218 , \11219 , \11220 , \11221 , \11222 ,
         \11223 , \11224 , \11225 , \11226 , \11227 , \11228 , \11229 , \11230 , \11231 , \11232 ,
         \11233 , \11234 , \11235 , \11236 , \11237 , \11238 , \11239 , \11240 , \11241 , \11242 ,
         \11243 , \11244 , \11245 , \11246 , \11247 , \11248 , \11249 , \11250 , \11251 , \11252 ,
         \11253 , \11254 , \11255 , \11256 , \11257 , \11258 , \11259 , \11260 , \11261 , \11262 ,
         \11263 , \11264 , \11265 , \11266 , \11267 , \11268 , \11269 , \11270 , \11271 , \11272 ,
         \11273 , \11274 , \11275 , \11276 , \11277 , \11278 , \11279 , \11280 , \11281 , \11282 ,
         \11283 , \11284 , \11285 , \11286 , \11287 , \11288 , \11289 , \11290 , \11291 , \11292 ,
         \11293 , \11294 , \11295 , \11296 , \11297 , \11298 , \11299 , \11300 , \11301 , \11302 ,
         \11303 , \11304 , \11305 , \11306 , \11307 , \11308 , \11309 , \11310 , \11311 , \11312 ,
         \11313 , \11314 , \11315 , \11316 , \11317 , \11318 , \11319 , \11320 , \11321 , \11322 ,
         \11323 , \11324 , \11325 , \11326 , \11327 , \11328 , \11329 , \11330 , \11331 , \11332 ,
         \11333 , \11334 , \11335 , \11336 , \11337 , \11338 , \11339 , \11340 , \11341 , \11342 ,
         \11343 , \11344 , \11345 , \11346 , \11347 , \11348 , \11349 , \11350 , \11351 , \11352 ,
         \11353 , \11354 , \11355 , \11356 , \11357 , \11358 , \11359 , \11360 , \11361 , \11362 ,
         \11363 , \11364 , \11365 , \11366 , \11367 , \11368 , \11369 , \11370 , \11371 , \11372 ,
         \11373 , \11374 , \11375 , \11376 , \11377 , \11378 , \11379 , \11380 , \11381 , \11382 ,
         \11383 , \11384 , \11385 , \11386 , \11387 , \11388 , \11389 , \11390 , \11391 , \11392 ,
         \11393 , \11394 , \11395 , \11396 , \11397 , \11398 , \11399 , \11400 , \11401 , \11402 ,
         \11403 , \11404 , \11405 , \11406 , \11407 , \11408 , \11409 , \11410 , \11411 , \11412 ,
         \11413 , \11414 , \11415 , \11416 , \11417 , \11418 , \11419 , \11420 , \11421 , \11422 ,
         \11423 , \11424 , \11425 , \11426 , \11427 , \11428 , \11429 , \11430 , \11431 , \11432 ,
         \11433 , \11434 , \11435 , \11436 , \11437 , \11438 , \11439 , \11440 , \11441 , \11442 ,
         \11443 , \11444 , \11445 , \11446 , \11447 , \11448 , \11449 , \11450 , \11451 , \11452 ,
         \11453 , \11454 , \11455 , \11456 , \11457 , \11458 , \11459 , \11460 , \11461 , \11462 ,
         \11463 , \11464 , \11465 , \11466 , \11467 , \11468 , \11469 , \11470 , \11471 , \11472 ,
         \11473 , \11474 , \11475 , \11476 , \11477 , \11478 , \11479 , \11480 , \11481 , \11482 ,
         \11483 , \11484 , \11485 , \11486 , \11487 , \11488 , \11489 , \11490 , \11491 , \11492 ,
         \11493 , \11494 , \11495 , \11496 , \11497 , \11498 , \11499 , \11500 , \11501 , \11502 ,
         \11503 , \11504 , \11505 , \11506 , \11507 , \11508 , \11509 , \11510 , \11511 , \11512 ,
         \11513 , \11514 , \11515 , \11516 , \11517 , \11518 , \11519 , \11520 , \11521 , \11522 ,
         \11523 , \11524 , \11525 , \11526 , \11527 , \11528 , \11529 , \11530 , \11531 , \11532 ,
         \11533 , \11534 , \11535 , \11536 , \11537 , \11538 , \11539 , \11540 , \11541 , \11542 ,
         \11543 , \11544 , \11545 , \11546 , \11547 , \11548 , \11549 , \11550 , \11551 , \11552 ,
         \11553 , \11554 , \11555 , \11556 , \11557 , \11558 , \11559 , \11560 , \11561 , \11562 ,
         \11563 , \11564 , \11565 , \11566 , \11567 , \11568 , \11569 , \11570 , \11571 , \11572 ,
         \11573 , \11574 , \11575 , \11576 , \11577 , \11578 , \11579 , \11580 , \11581 , \11582 ,
         \11583 , \11584 , \11585 , \11586 , \11587 , \11588 , \11589 , \11590 , \11591 , \11592 ,
         \11593 , \11594 , \11595 , \11596 , \11597 , \11598 , \11599 , \11600 , \11601 , \11602 ,
         \11603 , \11604 , \11605 , \11606 , \11607 , \11608 , \11609 , \11610 , \11611 , \11612 ,
         \11613 , \11614 , \11615 , \11616 , \11617 , \11618 , \11619 , \11620 , \11621 , \11622 ,
         \11623 , \11624 , \11625 , \11626 , \11627 , \11628 , \11629 , \11630 , \11631 , \11632 ,
         \11633 , \11634 , \11635 , \11636 , \11637 , \11638 , \11639 , \11640 , \11641 , \11642 ,
         \11643 , \11644 , \11645 , \11646 , \11647 , \11648 , \11649 , \11650 , \11651 , \11652 ,
         \11653 , \11654 , \11655 , \11656 , \11657 , \11658 , \11659 , \11660 , \11661 , \11662 ,
         \11663 , \11664 , \11665 , \11666 , \11667 , \11668 , \11669 , \11670 , \11671 , \11672 ,
         \11673 , \11674 , \11675 , \11676 , \11677 , \11678 , \11679 , \11680 , \11681 , \11682 ,
         \11683 , \11684 , \11685 , \11686 , \11687 , \11688 , \11689 , \11690 , \11691 , \11692 ,
         \11693 , \11694 , \11695 , \11696 , \11697 , \11698 , \11699 , \11700 , \11701 , \11702 ,
         \11703 , \11704 , \11705 , \11706 , \11707 , \11708 , \11709 , \11710 , \11711 , \11712 ,
         \11713 , \11714 , \11715 , \11716 , \11717 , \11718 , \11719 , \11720 , \11721 , \11722 ,
         \11723 , \11724 , \11725 , \11726 , \11727 , \11728 , \11729 , \11730 , \11731 , \11732 ,
         \11733 , \11734 , \11735 , \11736 , \11737 , \11738 , \11739 , \11740 , \11741 , \11742 ,
         \11743 , \11744 , \11745 , \11746 , \11747 , \11748 , \11749 , \11750 , \11751 , \11752 ,
         \11753 , \11754 , \11755 , \11756 , \11757 , \11758 , \11759 , \11760 , \11761 , \11762 ,
         \11763 , \11764 , \11765 , \11766 , \11767 , \11768 , \11769 , \11770 , \11771 , \11772 ,
         \11773 , \11774 , \11775 , \11776 , \11777 , \11778 , \11779 , \11780 , \11781 , \11782 ,
         \11783 , \11784 , \11785 , \11786 , \11787 , \11788 , \11789 , \11790 , \11791 , \11792 ,
         \11793 , \11794 , \11795 , \11796 , \11797 , \11798 , \11799 , \11800 , \11801 , \11802 ,
         \11803 , \11804 , \11805 , \11806 , \11807 , \11808 , \11809 , \11810 , \11811 , \11812 ,
         \11813 , \11814 , \11815 , \11816 , \11817 , \11818 , \11819 , \11820 , \11821 , \11822 ,
         \11823 , \11824 , \11825 , \11826 , \11827 , \11828 , \11829 , \11830 , \11831 , \11832 ,
         \11833 , \11834 , \11835 , \11836 , \11837 , \11838 , \11839 , \11840 , \11841 , \11842 ,
         \11843 , \11844 , \11845 , \11846 , \11847 , \11848 , \11849 , \11850 , \11851 , \11852 ,
         \11853 , \11854 , \11855 , \11856 , \11857 , \11858 , \11859 , \11860 , \11861 , \11862 ,
         \11863 , \11864 , \11865 , \11866 , \11867 , \11868 , \11869 , \11870 , \11871 , \11872 ,
         \11873 , \11874 , \11875 , \11876 , \11877 , \11878 , \11879 , \11880 , \11881 , \11882 ,
         \11883 , \11884 , \11885 , \11886 , \11887 , \11888 , \11889 , \11890 , \11891 , \11892 ,
         \11893 , \11894 , \11895 , \11896 , \11897 , \11898 , \11899 , \11900 , \11901 , \11902 ,
         \11903 , \11904 , \11905 , \11906 , \11907 , \11908 , \11909 , \11910 , \11911 , \11912 ,
         \11913 , \11914 , \11915 , \11916 , \11917 , \11918 , \11919 , \11920 , \11921 , \11922 ,
         \11923 , \11924 , \11925 , \11926 , \11927 , \11928 , \11929 , \11930 , \11931 , \11932 ,
         \11933 , \11934 , \11935 , \11936 , \11937 , \11938 , \11939 , \11940 , \11941 , \11942 ,
         \11943 , \11944 , \11945 , \11946 , \11947 , \11948 , \11949 , \11950 , \11951 , \11952 ,
         \11953 , \11954 , \11955 , \11956 , \11957 , \11958 , \11959 , \11960 , \11961 , \11962 ,
         \11963 , \11964 , \11965 , \11966 , \11967 , \11968 , \11969 , \11970 , \11971 , \11972 ,
         \11973 , \11974 , \11975 , \11976 , \11977 , \11978 , \11979 , \11980 , \11981 , \11982 ,
         \11983 , \11984 , \11985 , \11986 , \11987 , \11988 , \11989 , \11990 , \11991 , \11992 ,
         \11993 , \11994 , \11995 , \11996 , \11997 , \11998 , \11999 , \12000 , \12001 , \12002 ,
         \12003 , \12004 , \12005 , \12006 , \12007 , \12008 , \12009 , \12010 , \12011 , \12012 ,
         \12013 , \12014 , \12015 , \12016 , \12017 , \12018 , \12019 , \12020 , \12021 , \12022 ,
         \12023 , \12024 , \12025 , \12026 , \12027 , \12028 , \12029 , \12030 , \12031 , \12032 ,
         \12033 , \12034 , \12035 , \12036 , \12037 , \12038 , \12039 , \12040 , \12041 , \12042 ,
         \12043 , \12044 , \12045 , \12046 , \12047 , \12048 , \12049 , \12050 , \12051 , \12052 ,
         \12053 , \12054 , \12055 , \12056 , \12057 , \12058 , \12059 , \12060 , \12061 , \12062 ,
         \12063 , \12064 , \12065 , \12066 , \12067 , \12068 , \12069 , \12070 , \12071 , \12072 ,
         \12073 , \12074 , \12075 , \12076 , \12077 , \12078 , \12079 , \12080 , \12081 , \12082 ,
         \12083 , \12084 , \12085 , \12086 , \12087 , \12088 , \12089 , \12090 , \12091 , \12092 ,
         \12093 , \12094 , \12095 , \12096 , \12097 , \12098 , \12099 , \12100 , \12101 , \12102 ,
         \12103 , \12104 , \12105 , \12106 , \12107 , \12108 , \12109 , \12110 , \12111 , \12112 ,
         \12113 , \12114 , \12115 , \12116 , \12117 , \12118 , \12119 , \12120 , \12121 , \12122 ,
         \12123 , \12124 , \12125 , \12126 , \12127 , \12128 , \12129 , \12130 , \12131 , \12132 ,
         \12133 , \12134 , \12135 , \12136 , \12137 , \12138 , \12139 , \12140 , \12141 , \12142 ,
         \12143 , \12144 , \12145 , \12146 , \12147 , \12148 , \12149 , \12150 , \12151 , \12152 ,
         \12153 , \12154 , \12155 , \12156 , \12157 , \12158 , \12159 , \12160 , \12161 , \12162 ,
         \12163 , \12164 , \12165 , \12166 , \12167 , \12168 , \12169 , \12170 , \12171 , \12172 ,
         \12173 , \12174 , \12175 , \12176 , \12177 , \12178 , \12179 , \12180 , \12181 , \12182 ,
         \12183 , \12184 , \12185 , \12186 , \12187 , \12188 , \12189 , \12190 , \12191 , \12192 ,
         \12193 , \12194 , \12195 , \12196 , \12197 , \12198 , \12199 , \12200 , \12201 , \12202 ,
         \12203 , \12204 , \12205 , \12206 , \12207 , \12208 , \12209 , \12210 , \12211 , \12212 ,
         \12213 , \12214 , \12215 , \12216 , \12217 , \12218 , \12219 , \12220 , \12221 , \12222 ,
         \12223 , \12224 , \12225 , \12226 , \12227 , \12228 , \12229 , \12230 , \12231 , \12232 ,
         \12233 , \12234 , \12235 , \12236 , \12237 , \12238 , \12239 , \12240 , \12241 , \12242 ,
         \12243 , \12244 , \12245 , \12246 , \12247 , \12248 , \12249 , \12250 , \12251 , \12252 ,
         \12253 , \12254 , \12255 , \12256 , \12257 , \12258 , \12259 , \12260 , \12261 , \12262 ,
         \12263 , \12264 , \12265 , \12266 , \12267 , \12268 , \12269 , \12270 , \12271 , \12272 ,
         \12273 , \12274 , \12275 , \12276 , \12277 , \12278 , \12279 , \12280 , \12281 , \12282 ,
         \12283 , \12284 , \12285 , \12286 , \12287 , \12288 , \12289 , \12290 , \12291 , \12292 ,
         \12293 , \12294 , \12295 , \12296 , \12297 , \12298 , \12299 , \12300 , \12301 , \12302 ,
         \12303 , \12304 , \12305 , \12306 , \12307 , \12308 , \12309 , \12310 , \12311 , \12312 ,
         \12313 , \12314 , \12315 , \12316 , \12317 , \12318 , \12319 , \12320 , \12321 , \12322 ,
         \12323 , \12324 , \12325 , \12326 , \12327 , \12328 , \12329 , \12330 , \12331 , \12332 ,
         \12333 , \12334 , \12335 , \12336 , \12337 , \12338 , \12339 , \12340 , \12341 , \12342 ,
         \12343 , \12344 , \12345 , \12346 , \12347 , \12348 , \12349 , \12350 , \12351 , \12352 ,
         \12353 , \12354 , \12355 , \12356 , \12357 , \12358 , \12359 , \12360 , \12361 , \12362 ,
         \12363 , \12364 , \12365 , \12366 , \12367 , \12368 , \12369 , \12370 , \12371 , \12372 ,
         \12373 , \12374 , \12375 , \12376 , \12377 , \12378 , \12379 , \12380 , \12381 , \12382 ,
         \12383 , \12384 , \12385 , \12386 , \12387 , \12388 , \12389 , \12390 , \12391 , \12392 ,
         \12393 , \12394 , \12395 , \12396 , \12397 , \12398 , \12399 , \12400 , \12401 , \12402 ,
         \12403 , \12404 , \12405 , \12406 , \12407 , \12408 , \12409 , \12410 , \12411 , \12412 ,
         \12413 , \12414 , \12415 , \12416 , \12417 , \12418 , \12419 , \12420 , \12421 , \12422 ,
         \12423 , \12424 , \12425 , \12426 , \12427 , \12428 , \12429 , \12430 , \12431 , \12432 ,
         \12433 , \12434 , \12435 , \12436 , \12437 , \12438 , \12439 , \12440 , \12441 , \12442 ,
         \12443 , \12444 , \12445 , \12446 , \12447 , \12448 , \12449 , \12450 , \12451 , \12452 ,
         \12453 , \12454 , \12455 , \12456 , \12457 , \12458 , \12459 , \12460 , \12461 , \12462 ,
         \12463 , \12464 , \12465 , \12466 , \12467 , \12468 , \12469 , \12470 , \12471 , \12472 ,
         \12473 , \12474 , \12475 , \12476 , \12477 , \12478 , \12479 , \12480 , \12481 , \12482 ,
         \12483 , \12484 , \12485 , \12486 , \12487 , \12488 , \12489 , \12490 , \12491 , \12492 ,
         \12493 , \12494 , \12495 , \12496 , \12497 , \12498 , \12499 , \12500 , \12501 , \12502 ,
         \12503 , \12504 , \12505 , \12506 , \12507 , \12508 , \12509 , \12510 , \12511 , \12512 ,
         \12513 , \12514 , \12515 , \12516 , \12517 , \12518 , \12519 , \12520 , \12521 , \12522 ,
         \12523 , \12524 , \12525 , \12526 , \12527 , \12528 , \12529 , \12530 , \12531 , \12532 ,
         \12533 , \12534 , \12535 , \12536 , \12537 , \12538 , \12539 , \12540 , \12541 , \12542 ,
         \12543 , \12544 , \12545 , \12546 , \12547 , \12548 , \12549 , \12550 , \12551 , \12552 ,
         \12553 , \12554 , \12555 , \12556 , \12557 , \12558 , \12559 , \12560 , \12561 , \12562 ,
         \12563 , \12564 , \12565 , \12566 , \12567 , \12568 , \12569 , \12570 , \12571 , \12572 ,
         \12573 , \12574 , \12575 , \12576 , \12577 , \12578 , \12579 , \12580 , \12581 , \12582 ,
         \12583 , \12584 , \12585 , \12586 , \12587 , \12588 , \12589 , \12590 , \12591 , \12592 ,
         \12593 , \12594 , \12595 , \12596 , \12597 , \12598 , \12599 , \12600 , \12601 , \12602 ,
         \12603 , \12604 , \12605 , \12606 , \12607 , \12608 , \12609 , \12610 , \12611 , \12612 ,
         \12613 , \12614 , \12615 , \12616 , \12617 , \12618 , \12619 , \12620 , \12621 , \12622 ,
         \12623 , \12624 , \12625 , \12626 , \12627 , \12628 , \12629 , \12630 , \12631 , \12632 ,
         \12633 , \12634 , \12635 , \12636 , \12637 , \12638 , \12639 , \12640 , \12641 , \12642 ,
         \12643 , \12644 , \12645 , \12646 , \12647 , \12648 , \12649 , \12650 , \12651 , \12652 ,
         \12653 , \12654 , \12655 , \12656 , \12657 , \12658 , \12659 , \12660 , \12661 , \12662 ,
         \12663 , \12664 , \12665 , \12666 , \12667 , \12668 , \12669 , \12670 , \12671 , \12672 ,
         \12673 , \12674 , \12675 , \12676 , \12677 , \12678 , \12679 , \12680 , \12681 , \12682 ,
         \12683 , \12684 , \12685 , \12686 , \12687 , \12688 , \12689 , \12690 , \12691 , \12692 ,
         \12693 , \12694 , \12695 , \12696 , \12697 , \12698 , \12699 , \12700 , \12701 , \12702 ,
         \12703 , \12704 , \12705 , \12706 , \12707 , \12708 , \12709 , \12710 , \12711 , \12712 ,
         \12713 , \12714 , \12715 , \12716 , \12717 , \12718 , \12719 , \12720 , \12721 , \12722 ,
         \12723 , \12724 , \12725 , \12726 , \12727 , \12728 , \12729 , \12730 , \12731 , \12732 ,
         \12733 , \12734 , \12735 , \12736 , \12737 , \12738 , \12739 , \12740 , \12741 , \12742 ,
         \12743 , \12744 , \12745 , \12746 , \12747 , \12748 , \12749 , \12750 , \12751 , \12752 ,
         \12753 , \12754 , \12755 , \12756 , \12757 , \12758 , \12759 , \12760 , \12761 , \12762 ,
         \12763 , \12764 , \12765 , \12766 , \12767 , \12768 , \12769 , \12770 , \12771 , \12772 ,
         \12773 , \12774 , \12775 , \12776 , \12777 , \12778 , \12779 , \12780 , \12781 , \12782 ,
         \12783 , \12784 , \12785 , \12786 , \12787 , \12788 , \12789 , \12790 , \12791 , \12792 ,
         \12793 , \12794 , \12795 , \12796 , \12797 , \12798 , \12799 , \12800 , \12801 , \12802 ,
         \12803 , \12804 , \12805 , \12806 , \12807 , \12808 , \12809 , \12810 , \12811 , \12812 ,
         \12813 , \12814 , \12815 , \12816 , \12817 , \12818 , \12819 , \12820 , \12821 , \12822 ,
         \12823 , \12824 , \12825 , \12826 , \12827 , \12828 , \12829 , \12830 , \12831 , \12832 ,
         \12833 , \12834 , \12835 , \12836 , \12837 , \12838 , \12839 , \12840 , \12841 , \12842 ,
         \12843 , \12844 , \12845 , \12846 , \12847 , \12848 , \12849 , \12850 , \12851 , \12852 ,
         \12853 , \12854 , \12855 , \12856 , \12857 , \12858 , \12859 , \12860 , \12861 , \12862 ,
         \12863 , \12864 , \12865 , \12866 , \12867 , \12868 , \12869 , \12870 , \12871 , \12872 ,
         \12873 , \12874 , \12875 , \12876 , \12877 , \12878 , \12879 , \12880 , \12881 , \12882 ,
         \12883 , \12884 , \12885 , \12886 , \12887 , \12888 , \12889 , \12890 , \12891 , \12892 ,
         \12893 , \12894 , \12895 , \12896 , \12897 , \12898 , \12899 , \12900 , \12901 , \12902 ,
         \12903 , \12904 , \12905 , \12906 , \12907 , \12908 , \12909 , \12910 , \12911 , \12912 ,
         \12913 , \12914 , \12915 , \12916 , \12917 , \12918 , \12919 , \12920 , \12921 , \12922 ,
         \12923 , \12924 , \12925 , \12926 , \12927 , \12928 , \12929 , \12930 , \12931 , \12932 ,
         \12933 , \12934 , \12935 , \12936 , \12937 , \12938 , \12939 , \12940 , \12941 , \12942 ,
         \12943 , \12944 , \12945 , \12946 , \12947 , \12948 , \12949 , \12950 , \12951 , \12952 ,
         \12953 , \12954 , \12955 , \12956 , \12957 , \12958 , \12959 , \12960 , \12961 , \12962 ,
         \12963 , \12964 , \12965 , \12966 , \12967 , \12968 , \12969 , \12970 , \12971 , \12972 ,
         \12973 , \12974 , \12975 , \12976 , \12977 , \12978 , \12979 , \12980 , \12981 , \12982 ,
         \12983 , \12984 , \12985 , \12986 , \12987 , \12988 , \12989 , \12990 , \12991 , \12992 ,
         \12993 , \12994 , \12995 , \12996 , \12997 , \12998 , \12999 , \13000 , \13001 , \13002 ,
         \13003 , \13004 , \13005 , \13006 , \13007 , \13008 , \13009 , \13010 , \13011 , \13012 ,
         \13013 , \13014 , \13015 , \13016 , \13017 , \13018 , \13019 , \13020 , \13021 , \13022 ,
         \13023 , \13024 , \13025 , \13026 , \13027 , \13028 , \13029 , \13030 , \13031 , \13032 ,
         \13033 , \13034 , \13035 , \13036 , \13037 , \13038 , \13039 , \13040 , \13041 , \13042 ,
         \13043 , \13044 , \13045 , \13046 , \13047 , \13048 , \13049 , \13050 , \13051 , \13052 ,
         \13053 , \13054 , \13055 , \13056 , \13057 , \13058 , \13059 , \13060 , \13061 , \13062 ,
         \13063 , \13064 , \13065 , \13066 , \13067 , \13068 , \13069 , \13070 , \13071 , \13072 ,
         \13073 , \13074 , \13075 , \13076 , \13077 , \13078 , \13079 , \13080 , \13081 , \13082 ,
         \13083 , \13084 , \13085 , \13086 , \13087 , \13088 , \13089 , \13090 , \13091 , \13092 ,
         \13093 , \13094 , \13095 , \13096 , \13097 , \13098 , \13099 , \13100 , \13101 , \13102 ,
         \13103 , \13104 , \13105 , \13106 , \13107 , \13108 , \13109 , \13110 , \13111 , \13112 ,
         \13113 , \13114 , \13115 , \13116 , \13117 , \13118 , \13119 , \13120 , \13121 , \13122 ,
         \13123 , \13124 , \13125 , \13126 , \13127 , \13128 , \13129 , \13130 , \13131 , \13132 ,
         \13133 , \13134 , \13135 , \13136 , \13137 , \13138 , \13139 , \13140 , \13141 , \13142 ,
         \13143 , \13144 , \13145 , \13146 , \13147 , \13148 , \13149 , \13150 , \13151 , \13152 ,
         \13153 , \13154 , \13155 , \13156 , \13157 , \13158 , \13159 , \13160 , \13161 , \13162 ,
         \13163 , \13164 , \13165 , \13166 , \13167 , \13168 , \13169 , \13170 , \13171 , \13172 ,
         \13173 , \13174 , \13175 , \13176 , \13177 , \13178 , \13179 , \13180 , \13181 , \13182 ,
         \13183 , \13184 , \13185 , \13186 , \13187 , \13188 , \13189 , \13190 , \13191 , \13192 ,
         \13193 , \13194 , \13195 , \13196 , \13197 , \13198 , \13199 , \13200 , \13201 , \13202 ,
         \13203 , \13204 , \13205 , \13206 , \13207 , \13208 , \13209 , \13210 , \13211 , \13212 ,
         \13213 , \13214 , \13215 , \13216 , \13217 , \13218 , \13219 , \13220 , \13221 , \13222 ,
         \13223 , \13224 , \13225 , \13226 , \13227 , \13228 , \13229 , \13230 , \13231 , \13232 ,
         \13233 , \13234 , \13235 , \13236 , \13237 , \13238 , \13239 , \13240 , \13241 , \13242 ,
         \13243 , \13244 , \13245 , \13246 , \13247 , \13248 , \13249 , \13250 , \13251 , \13252 ,
         \13253 , \13254 , \13255 , \13256 , \13257 , \13258 , \13259 , \13260 , \13261 , \13262 ,
         \13263 , \13264 , \13265 , \13266 , \13267 , \13268 , \13269 , \13270 , \13271 , \13272 ,
         \13273 , \13274 , \13275 , \13276 , \13277 , \13278 , \13279 , \13280 , \13281 , \13282 ,
         \13283 , \13284 , \13285 , \13286 , \13287 , \13288 , \13289 , \13290 , \13291 , \13292 ,
         \13293 , \13294 , \13295 , \13296 , \13297 , \13298 , \13299 , \13300 , \13301 , \13302 ,
         \13303 , \13304 , \13305 , \13306 , \13307 , \13308 , \13309 , \13310 , \13311 , \13312 ,
         \13313 , \13314 , \13315 , \13316 , \13317 , \13318 , \13319 , \13320 , \13321 , \13322 ,
         \13323 , \13324 , \13325 , \13326 , \13327 , \13328 , \13329 , \13330 , \13331 , \13332 ,
         \13333 , \13334 , \13335 , \13336 , \13337 , \13338 , \13339 , \13340 , \13341 , \13342 ,
         \13343 , \13344 , \13345 , \13346 , \13347 , \13348 , \13349 , \13350 , \13351 , \13352 ,
         \13353 , \13354 , \13355 , \13356 , \13357 , \13358 , \13359 , \13360 , \13361 , \13362 ,
         \13363 , \13364 , \13365 , \13366 , \13367 , \13368 , \13369 , \13370 , \13371 , \13372 ,
         \13373 , \13374 , \13375 , \13376 , \13377 , \13378 , \13379 , \13380 , \13381 , \13382 ,
         \13383 , \13384 , \13385 , \13386 , \13387 , \13388 , \13389 , \13390 , \13391 , \13392 ,
         \13393 , \13394 , \13395 , \13396 , \13397 , \13398 , \13399 , \13400 , \13401 , \13402 ,
         \13403 , \13404 , \13405 , \13406 , \13407 , \13408 , \13409 , \13410 , \13411 , \13412 ,
         \13413 , \13414 , \13415 , \13416 , \13417 , \13418 , \13419 , \13420 , \13421 , \13422 ,
         \13423 , \13424 , \13425 , \13426 , \13427 , \13428 , \13429 , \13430 , \13431 , \13432 ,
         \13433 , \13434 , \13435 , \13436 , \13437 , \13438 , \13439 , \13440 , \13441 , \13442 ,
         \13443 , \13444 , \13445 , \13446 , \13447 , \13448 , \13449 , \13450 , \13451 , \13452 ,
         \13453 , \13454 , \13455 , \13456 , \13457 , \13458 , \13459 , \13460 , \13461 , \13462 ,
         \13463 , \13464 , \13465 , \13466 , \13467 , \13468 , \13469 , \13470 , \13471 , \13472 ,
         \13473 , \13474 , \13475 , \13476 , \13477 , \13478 , \13479 , \13480 , \13481 , \13482 ,
         \13483 , \13484 , \13485 , \13486 , \13487 , \13488 , \13489 , \13490 , \13491 , \13492 ,
         \13493 , \13494 , \13495 , \13496 , \13497 , \13498 , \13499 , \13500 , \13501 , \13502 ,
         \13503 , \13504 , \13505 , \13506 , \13507 , \13508 , \13509 , \13510 , \13511 , \13512 ,
         \13513 , \13514 , \13515 , \13516 , \13517 , \13518 , \13519 , \13520 , \13521 , \13522 ,
         \13523 , \13524 , \13525 , \13526 , \13527 , \13528 , \13529 , \13530 , \13531 , \13532 ,
         \13533 , \13534 , \13535 , \13536 , \13537 , \13538 , \13539 , \13540 , \13541 , \13542 ,
         \13543 , \13544 , \13545 , \13546 , \13547 , \13548 , \13549 , \13550 , \13551 , \13552 ,
         \13553 , \13554 , \13555 , \13556 , \13557 , \13558 , \13559 , \13560 , \13561 , \13562 ,
         \13563 , \13564 , \13565 , \13566 , \13567 , \13568 , \13569 , \13570 , \13571 , \13572 ,
         \13573 , \13574 , \13575 , \13576 , \13577 , \13578 , \13579 , \13580 , \13581 , \13582 ,
         \13583 , \13584 , \13585 , \13586 , \13587 , \13588 , \13589 , \13590 , \13591 , \13592 ,
         \13593 , \13594 , \13595 , \13596 , \13597 , \13598 , \13599 , \13600 , \13601 , \13602 ,
         \13603 , \13604 , \13605 , \13606 , \13607 , \13608 , \13609 , \13610 , \13611 , \13612 ,
         \13613 , \13614 , \13615 , \13616 , \13617 , \13618 , \13619 , \13620 , \13621 , \13622 ,
         \13623 , \13624 , \13625 , \13626 , \13627 , \13628 , \13629 , \13630 , \13631 , \13632 ,
         \13633 , \13634 , \13635 , \13636 , \13637 , \13638 , \13639 , \13640 , \13641 , \13642 ,
         \13643 , \13644 , \13645 , \13646 , \13647 , \13648 , \13649 , \13650 , \13651 , \13652 ,
         \13653 , \13654 , \13655 , \13656 , \13657 , \13658 , \13659 , \13660 , \13661 , \13662 ,
         \13663 , \13664 , \13665 , \13666 , \13667 , \13668 , \13669 , \13670 , \13671 , \13672 ,
         \13673 , \13674 , \13675 , \13676 , \13677 , \13678 , \13679 , \13680 , \13681 , \13682 ,
         \13683 , \13684 , \13685 , \13686 , \13687 , \13688 , \13689 , \13690 , \13691 , \13692 ,
         \13693 , \13694 , \13695 , \13696 , \13697 , \13698 , \13699 , \13700 , \13701 , \13702 ,
         \13703 , \13704 , \13705 , \13706 , \13707 , \13708 , \13709 , \13710 , \13711 , \13712 ,
         \13713 , \13714 , \13715 , \13716 , \13717 , \13718 , \13719 , \13720 , \13721 , \13722 ,
         \13723 , \13724 , \13725 , \13726 , \13727 , \13728 , \13729 , \13730 , \13731 , \13732 ,
         \13733 , \13734 , \13735 , \13736 , \13737 , \13738 , \13739 , \13740 , \13741 , \13742 ,
         \13743 , \13744 , \13745 , \13746 , \13747 , \13748 , \13749 , \13750 , \13751 , \13752 ,
         \13753 , \13754 , \13755 , \13756 , \13757 , \13758 , \13759 , \13760 , \13761 , \13762 ,
         \13763 , \13764 , \13765 , \13766 , \13767 , \13768 , \13769 , \13770 , \13771 , \13772 ,
         \13773 , \13774 , \13775 , \13776 , \13777 , \13778 , \13779 , \13780 , \13781 , \13782 ,
         \13783 , \13784 , \13785 , \13786 , \13787 , \13788 , \13789 , \13790 , \13791 , \13792 ,
         \13793 , \13794 , \13795 , \13796 , \13797 , \13798 , \13799 , \13800 , \13801 , \13802 ,
         \13803 , \13804 , \13805 , \13806 , \13807 , \13808 , \13809 , \13810 , \13811 , \13812 ,
         \13813 , \13814 , \13815 , \13816 , \13817 , \13818 , \13819 , \13820 , \13821 , \13822 ,
         \13823 , \13824 , \13825 , \13826 , \13827 , \13828 , \13829 , \13830 , \13831 , \13832 ,
         \13833 , \13834 , \13835 , \13836 , \13837 , \13838 , \13839 , \13840 , \13841 , \13842 ,
         \13843 , \13844 , \13845 , \13846 , \13847 , \13848 , \13849 , \13850 , \13851 , \13852 ,
         \13853 , \13854 , \13855 , \13856 , \13857 , \13858 , \13859 , \13860 , \13861 , \13862 ,
         \13863 , \13864 , \13865 , \13866 , \13867 , \13868 , \13869 , \13870 , \13871 , \13872 ,
         \13873 , \13874 , \13875 , \13876 , \13877 , \13878 , \13879 , \13880 , \13881 , \13882 ,
         \13883 , \13884 , \13885 , \13886 , \13887 , \13888 , \13889 , \13890 , \13891 , \13892 ,
         \13893 , \13894 , \13895 , \13896 , \13897 , \13898 , \13899 , \13900 , \13901 , \13902 ,
         \13903 , \13904 , \13905 , \13906 , \13907 , \13908 , \13909 , \13910 , \13911 , \13912 ,
         \13913 , \13914 , \13915 , \13916 , \13917 , \13918 , \13919 , \13920 , \13921 , \13922 ,
         \13923 , \13924 , \13925 , \13926 , \13927 , \13928 , \13929 , \13930 , \13931 , \13932 ,
         \13933 , \13934 , \13935 , \13936 , \13937 , \13938 , \13939 , \13940 , \13941 , \13942 ,
         \13943 , \13944 , \13945 , \13946 , \13947 , \13948 , \13949 , \13950 , \13951 , \13952 ,
         \13953 , \13954 , \13955 , \13956 , \13957 , \13958 , \13959 , \13960 , \13961 , \13962 ,
         \13963 , \13964 , \13965 , \13966 , \13967 , \13968 , \13969 , \13970 , \13971 , \13972 ,
         \13973 , \13974 , \13975 , \13976 , \13977 , \13978 , \13979 , \13980 , \13981 , \13982 ,
         \13983 , \13984 , \13985 , \13986 , \13987 , \13988 , \13989 , \13990 , \13991 , \13992 ,
         \13993 , \13994 , \13995 , \13996 , \13997 , \13998 , \13999 , \14000 , \14001 , \14002 ,
         \14003 , \14004 , \14005 , \14006 , \14007 , \14008 , \14009 , \14010 , \14011 , \14012 ,
         \14013 , \14014 , \14015 , \14016 , \14017 , \14018 , \14019 , \14020 , \14021 , \14022 ,
         \14023 , \14024 , \14025 , \14026 , \14027 , \14028 , \14029 , \14030 , \14031 , \14032 ,
         \14033 , \14034 , \14035 , \14036 , \14037 , \14038 , \14039 , \14040 , \14041 , \14042 ,
         \14043 , \14044 , \14045 , \14046 , \14047 , \14048 , \14049 , \14050 , \14051 , \14052 ,
         \14053 , \14054 , \14055 , \14056 , \14057 , \14058 , \14059 , \14060 , \14061 , \14062 ,
         \14063 , \14064 , \14065 , \14066 , \14067 , \14068 , \14069 , \14070 , \14071 , \14072 ,
         \14073 , \14074 , \14075 , \14076 , \14077 , \14078 , \14079 , \14080 , \14081 , \14082 ,
         \14083 , \14084 , \14085 , \14086 , \14087 , \14088 , \14089 , \14090 , \14091 , \14092 ,
         \14093 , \14094 , \14095 , \14096 , \14097 , \14098 , \14099 , \14100 , \14101 , \14102 ,
         \14103 , \14104 , \14105 , \14106 , \14107 , \14108 , \14109 , \14110 , \14111 , \14112 ,
         \14113 , \14114 , \14115 , \14116 , \14117 , \14118 , \14119 , \14120 , \14121 , \14122 ,
         \14123 , \14124 , \14125 , \14126 , \14127 , \14128 , \14129 , \14130 , \14131 , \14132 ,
         \14133 , \14134 , \14135 , \14136 , \14137 , \14138 , \14139 , \14140 , \14141 , \14142 ,
         \14143 , \14144 , \14145 , \14146 , \14147 , \14148 , \14149 , \14150 , \14151 , \14152 ,
         \14153 , \14154 , \14155 , \14156 , \14157 , \14158 , \14159 , \14160 , \14161 , \14162 ,
         \14163 , \14164 , \14165 , \14166 , \14167 , \14168 , \14169 , \14170 , \14171 , \14172 ,
         \14173 , \14174 , \14175 , \14176 , \14177 , \14178 , \14179 , \14180 , \14181 , \14182 ,
         \14183 , \14184 , \14185 , \14186 , \14187 , \14188 , \14189 , \14190 , \14191 , \14192 ,
         \14193 , \14194 , \14195 , \14196 , \14197 , \14198 , \14199 , \14200 , \14201 , \14202 ,
         \14203 , \14204 , \14205 , \14206 , \14207 , \14208 , \14209 , \14210 , \14211 , \14212 ,
         \14213 , \14214 , \14215 , \14216 , \14217 , \14218 , \14219 , \14220 , \14221 , \14222 ,
         \14223 , \14224 , \14225 , \14226 , \14227 , \14228 , \14229 , \14230 , \14231 , \14232 ,
         \14233 , \14234 , \14235 , \14236 , \14237 , \14238 , \14239 , \14240 , \14241 , \14242 ,
         \14243 , \14244 , \14245 , \14246 , \14247 , \14248 , \14249 , \14250 , \14251 , \14252 ,
         \14253 , \14254 , \14255 , \14256 , \14257 , \14258 , \14259 , \14260 , \14261 , \14262 ,
         \14263 , \14264 , \14265 , \14266 , \14267 , \14268 , \14269 , \14270 , \14271 , \14272 ,
         \14273 , \14274 , \14275 , \14276 , \14277 , \14278 , \14279 , \14280 , \14281 , \14282 ,
         \14283 , \14284 , \14285 , \14286 , \14287 , \14288 , \14289 , \14290 , \14291 , \14292 ,
         \14293 , \14294 , \14295 , \14296 , \14297 , \14298 , \14299 , \14300 , \14301 , \14302 ,
         \14303 , \14304 , \14305 , \14306 , \14307 , \14308 , \14309 , \14310 , \14311 , \14312 ,
         \14313 , \14314 , \14315 , \14316 , \14317 , \14318 , \14319 , \14320 , \14321 , \14322 ,
         \14323 , \14324 , \14325 , \14326 , \14327 , \14328 , \14329 , \14330 , \14331 , \14332 ,
         \14333 , \14334 , \14335 , \14336 , \14337 , \14338 , \14339 , \14340 , \14341 , \14342 ,
         \14343 , \14344 , \14345 , \14346 , \14347 , \14348 , \14349 , \14350 , \14351 , \14352 ,
         \14353 , \14354 , \14355 , \14356 , \14357 , \14358 , \14359 , \14360 , \14361 , \14362 ,
         \14363 , \14364 , \14365 , \14366 , \14367 , \14368 , \14369 , \14370 , \14371 , \14372 ,
         \14373 , \14374 , \14375 , \14376 , \14377 , \14378 , \14379 , \14380 , \14381 , \14382 ,
         \14383 , \14384 , \14385 , \14386 , \14387 , \14388 , \14389 , \14390 , \14391 , \14392 ,
         \14393 , \14394 , \14395 , \14396 , \14397 , \14398 , \14399 , \14400 , \14401 , \14402 ,
         \14403 , \14404 , \14405 , \14406 , \14407 , \14408 , \14409 , \14410 , \14411 , \14412 ,
         \14413 , \14414 , \14415 , \14416 , \14417 , \14418 , \14419 , \14420 , \14421 , \14422 ,
         \14423 , \14424 , \14425 , \14426 , \14427 , \14428 , \14429 , \14430 , \14431 , \14432 ,
         \14433 , \14434 , \14435 , \14436 , \14437 , \14438 , \14439 , \14440 , \14441 , \14442 ,
         \14443 , \14444 , \14445 , \14446 , \14447 , \14448 , \14449 , \14450 , \14451 , \14452 ,
         \14453 , \14454 , \14455 , \14456 , \14457 , \14458 , \14459 , \14460 , \14461 , \14462 ,
         \14463 , \14464 , \14465 , \14466 , \14467 , \14468 , \14469 , \14470 , \14471 , \14472 ,
         \14473 , \14474 , \14475 , \14476 , \14477 , \14478 , \14479 , \14480 , \14481 , \14482 ,
         \14483 , \14484 , \14485 , \14486 , \14487 , \14488 , \14489 , \14490 , \14491 , \14492 ,
         \14493 , \14494 , \14495 , \14496 , \14497 , \14498 , \14499 , \14500 , \14501 , \14502 ,
         \14503 , \14504 , \14505 , \14506 , \14507 , \14508 , \14509 , \14510 , \14511 , \14512 ,
         \14513 , \14514 , \14515 , \14516 , \14517 , \14518 , \14519 , \14520 , \14521 , \14522 ,
         \14523 , \14524 , \14525 , \14526 , \14527 , \14528 , \14529 , \14530 , \14531 , \14532 ,
         \14533 , \14534 , \14535 , \14536 , \14537 , \14538 , \14539 , \14540 , \14541 , \14542 ,
         \14543 , \14544 , \14545 , \14546 , \14547 , \14548 , \14549 , \14550 , \14551 , \14552 ,
         \14553 , \14554 , \14555 , \14556 , \14557 , \14558 , \14559 , \14560 , \14561 , \14562 ,
         \14563 , \14564 , \14565 , \14566 , \14567 , \14568 , \14569 , \14570 , \14571 , \14572 ,
         \14573 , \14574 , \14575 , \14576 , \14577 , \14578 , \14579 , \14580 , \14581 , \14582 ,
         \14583 , \14584 , \14585 , \14586 , \14587 , \14588 , \14589 , \14590 , \14591 , \14592 ,
         \14593 , \14594 , \14595 , \14596 , \14597 , \14598 , \14599 , \14600 , \14601 , \14602 ,
         \14603 , \14604 , \14605 , \14606 , \14607 , \14608 , \14609 , \14610 , \14611 , \14612 ,
         \14613 , \14614 , \14615 , \14616 , \14617 , \14618 , \14619 , \14620 , \14621 , \14622 ,
         \14623 , \14624 , \14625 , \14626 , \14627 , \14628 , \14629 , \14630 , \14631 , \14632 ,
         \14633 , \14634 , \14635 , \14636 , \14637 , \14638 , \14639 , \14640 , \14641 , \14642 ,
         \14643 , \14644 , \14645 , \14646 , \14647 , \14648 , \14649 , \14650 , \14651 , \14652 ,
         \14653 , \14654 , \14655 , \14656 , \14657 , \14658 , \14659 , \14660 , \14661 , \14662 ,
         \14663 , \14664 , \14665 , \14666 , \14667 , \14668 , \14669 , \14670 , \14671 , \14672 ,
         \14673 , \14674 , \14675 , \14676 , \14677 , \14678 , \14679 , \14680 , \14681 , \14682 ,
         \14683 , \14684 , \14685 , \14686 , \14687 , \14688 , \14689 , \14690 , \14691 , \14692 ,
         \14693 , \14694 , \14695 , \14696 , \14697 , \14698 , \14699 , \14700 , \14701 , \14702 ,
         \14703 , \14704 , \14705 , \14706 , \14707 , \14708 , \14709 , \14710 , \14711 , \14712 ,
         \14713 , \14714 , \14715 , \14716 , \14717 , \14718 , \14719 , \14720 , \14721 , \14722 ,
         \14723 , \14724 , \14725 , \14726 , \14727 , \14728 , \14729 , \14730 , \14731 , \14732 ,
         \14733 , \14734 , \14735 , \14736 , \14737 , \14738 , \14739 , \14740 , \14741 , \14742 ,
         \14743 , \14744 , \14745 , \14746 , \14747 , \14748 , \14749 , \14750 , \14751 , \14752 ,
         \14753 , \14754 , \14755 , \14756 , \14757 , \14758 , \14759 , \14760 , \14761 , \14762 ,
         \14763 , \14764 , \14765 , \14766 , \14767 , \14768 , \14769 , \14770 , \14771 , \14772 ,
         \14773 , \14774 , \14775 , \14776 , \14777 , \14778 , \14779 , \14780 , \14781 , \14782 ,
         \14783 , \14784 , \14785 , \14786 , \14787 , \14788 , \14789 , \14790 , \14791 , \14792 ,
         \14793 , \14794 , \14795 , \14796 , \14797 , \14798 , \14799 , \14800 , \14801 , \14802 ,
         \14803 , \14804 , \14805 , \14806 , \14807 , \14808 , \14809 , \14810 , \14811 , \14812 ,
         \14813 , \14814 , \14815 , \14816 , \14817 , \14818 , \14819 , \14820 , \14821 , \14822 ,
         \14823 , \14824 , \14825 , \14826 , \14827 , \14828 , \14829 , \14830 , \14831 , \14832 ,
         \14833 , \14834 , \14835 , \14836 , \14837 , \14838 , \14839 , \14840 , \14841 , \14842 ,
         \14843 , \14844 , \14845 , \14846 , \14847 , \14848 , \14849 , \14850 , \14851 , \14852 ,
         \14853 , \14854 , \14855 , \14856 , \14857 , \14858 , \14859 , \14860 , \14861 , \14862 ,
         \14863 , \14864 , \14865 , \14866 , \14867 , \14868 , \14869 , \14870 , \14871 , \14872 ,
         \14873 , \14874 , \14875 , \14876 , \14877 , \14878 , \14879 , \14880 , \14881 , \14882 ,
         \14883 , \14884 , \14885 , \14886 , \14887 , \14888 , \14889 , \14890 , \14891 , \14892 ,
         \14893 , \14894 , \14895 , \14896 , \14897 , \14898 , \14899 , \14900 , \14901 , \14902 ,
         \14903 , \14904 , \14905 , \14906 , \14907 , \14908 , \14909 , \14910 , \14911 , \14912 ,
         \14913 , \14914 , \14915 , \14916 , \14917 , \14918 , \14919 , \14920 , \14921 , \14922 ,
         \14923 , \14924 , \14925 , \14926 , \14927 , \14928 , \14929 , \14930 , \14931 , \14932 ,
         \14933 , \14934 , \14935 , \14936 , \14937 , \14938 , \14939 , \14940 , \14941 , \14942 ,
         \14943 , \14944 , \14945 , \14946 , \14947 , \14948 , \14949 , \14950 , \14951 , \14952 ,
         \14953 , \14954 , \14955 , \14956 , \14957 , \14958 , \14959 , \14960 , \14961 , \14962 ,
         \14963 , \14964 , \14965 , \14966 , \14967 , \14968 , \14969 , \14970 , \14971 , \14972 ,
         \14973 , \14974 , \14975 , \14976 , \14977 , \14978 , \14979 , \14980 , \14981 , \14982 ,
         \14983 , \14984 , \14985 , \14986 , \14987 , \14988 , \14989 , \14990 , \14991 , \14992 ,
         \14993 , \14994 , \14995 , \14996 , \14997 , \14998 , \14999 , \15000 , \15001 , \15002 ,
         \15003 , \15004 , \15005 , \15006 , \15007 , \15008 , \15009 , \15010 , \15011 , \15012 ,
         \15013 , \15014 , \15015 , \15016 , \15017 , \15018 , \15019 , \15020 , \15021 , \15022 ,
         \15023 , \15024 , \15025 , \15026 , \15027 , \15028 , \15029 , \15030 , \15031 , \15032 ,
         \15033 , \15034 , \15035 , \15036 , \15037 , \15038 , \15039 , \15040 , \15041 , \15042 ,
         \15043 , \15044 , \15045 , \15046 , \15047 , \15048 , \15049 , \15050 , \15051 , \15052 ,
         \15053 , \15054 , \15055 , \15056 , \15057 , \15058 , \15059 , \15060 , \15061 , \15062 ,
         \15063 , \15064 , \15065 , \15066 , \15067 , \15068 , \15069 , \15070 , \15071 , \15072 ,
         \15073 , \15074 , \15075 , \15076 , \15077 , \15078 , \15079 , \15080 , \15081 , \15082 ,
         \15083 , \15084 , \15085 , \15086 , \15087 , \15088 , \15089 , \15090 , \15091 , \15092 ,
         \15093 , \15094 , \15095 , \15096 , \15097 , \15098 , \15099 , \15100 , \15101 , \15102 ,
         \15103 , \15104 , \15105 , \15106 , \15107 , \15108 , \15109 , \15110 , \15111 , \15112 ,
         \15113 , \15114 , \15115 , \15116 , \15117 , \15118 , \15119 , \15120 , \15121 , \15122 ,
         \15123 , \15124 , \15125 , \15126 , \15127 , \15128 , \15129 , \15130 , \15131 , \15132 ,
         \15133 , \15134 , \15135 , \15136 , \15137 , \15138 , \15139 , \15140 , \15141 , \15142 ,
         \15143 , \15144 , \15145 , \15146 , \15147 , \15148 , \15149 , \15150 , \15151 , \15152 ,
         \15153 , \15154 , \15155 , \15156 , \15157 , \15158 , \15159 , \15160 , \15161 , \15162 ,
         \15163 , \15164 , \15165 , \15166 , \15167 , \15168 , \15169 , \15170 , \15171 , \15172 ,
         \15173 , \15174 , \15175 , \15176 , \15177 , \15178 , \15179 , \15180 , \15181 , \15182 ,
         \15183 , \15184 , \15185 , \15186 , \15187 , \15188 , \15189 , \15190 , \15191 , \15192 ,
         \15193 , \15194 , \15195 , \15196 , \15197 , \15198 , \15199 , \15200 , \15201 , \15202 ,
         \15203 , \15204 , \15205 , \15206 , \15207 , \15208 , \15209 , \15210 , \15211 , \15212 ,
         \15213 , \15214 , \15215 , \15216 , \15217 , \15218 , \15219 , \15220 , \15221 , \15222 ,
         \15223 , \15224 , \15225 , \15226 , \15227 , \15228 , \15229 , \15230 , \15231 , \15232 ,
         \15233 , \15234 , \15235 , \15236 , \15237 , \15238 , \15239 , \15240 , \15241 , \15242 ,
         \15243 , \15244 , \15245 , \15246 , \15247 , \15248 , \15249 , \15250 , \15251 , \15252 ,
         \15253 , \15254 , \15255 , \15256 , \15257 , \15258 , \15259 , \15260 , \15261 , \15262 ,
         \15263 , \15264 , \15265 , \15266 , \15267 , \15268 , \15269 , \15270 , \15271 , \15272 ,
         \15273 , \15274 , \15275 , \15276 , \15277 , \15278 , \15279 , \15280 , \15281 , \15282 ,
         \15283 , \15284 , \15285 , \15286 , \15287 , \15288 , \15289 , \15290 , \15291 , \15292 ,
         \15293 , \15294 , \15295 , \15296 , \15297 , \15298 , \15299 , \15300 , \15301 , \15302 ,
         \15303 , \15304 , \15305 , \15306 , \15307 , \15308 , \15309 , \15310 , \15311 , \15312 ,
         \15313 , \15314 , \15315 , \15316 , \15317 , \15318 , \15319 , \15320 , \15321 , \15322 ,
         \15323 , \15324 , \15325 , \15326 , \15327 , \15328 , \15329 , \15330 , \15331 , \15332 ,
         \15333 , \15334 , \15335 , \15336 , \15337 , \15338 , \15339 , \15340 , \15341 , \15342 ,
         \15343 , \15344 , \15345 , \15346 , \15347 , \15348 , \15349 , \15350 , \15351 , \15352 ,
         \15353 , \15354 , \15355 , \15356 , \15357 , \15358 , \15359 , \15360 , \15361 , \15362 ,
         \15363 , \15364 , \15365 , \15366 , \15367 , \15368 , \15369 , \15370 , \15371 , \15372 ,
         \15373 , \15374 , \15375 , \15376 , \15377 , \15378 , \15379 , \15380 , \15381 , \15382 ,
         \15383 , \15384 , \15385 , \15386 , \15387 , \15388 , \15389 , \15390 , \15391 , \15392 ,
         \15393 , \15394 , \15395 , \15396 , \15397 , \15398 , \15399 , \15400 , \15401 , \15402 ,
         \15403 , \15404 , \15405 , \15406 , \15407 , \15408 , \15409 , \15410 , \15411 , \15412 ,
         \15413 , \15414 , \15415 , \15416 , \15417 , \15418 , \15419 , \15420 , \15421 , \15422 ,
         \15423 , \15424 , \15425 , \15426 , \15427 , \15428 , \15429 , \15430 , \15431 , \15432 ,
         \15433 , \15434 , \15435 , \15436 , \15437 , \15438 , \15439 , \15440 , \15441 , \15442 ,
         \15443 , \15444 , \15445 , \15446 , \15447 , \15448 , \15449 , \15450 , \15451 , \15452 ,
         \15453 , \15454 , \15455 , \15456 , \15457 , \15458 , \15459 , \15460 , \15461 , \15462 ,
         \15463 , \15464 , \15465 , \15466 , \15467 , \15468 , \15469 , \15470 , \15471 , \15472 ,
         \15473 , \15474 , \15475 , \15476 , \15477 , \15478 , \15479 , \15480 , \15481 , \15482 ,
         \15483 , \15484 , \15485 , \15486 , \15487 , \15488 , \15489 , \15490 , \15491 , \15492 ,
         \15493 , \15494 , \15495 , \15496 , \15497 , \15498 , \15499 , \15500 , \15501 , \15502 ,
         \15503 , \15504 , \15505 , \15506 , \15507 , \15508 , \15509 , \15510 , \15511 , \15512 ,
         \15513 , \15514 , \15515 , \15516 , \15517 , \15518 , \15519 , \15520 , \15521 , \15522 ,
         \15523 , \15524 , \15525 , \15526 , \15527 , \15528 , \15529 , \15530 , \15531 , \15532 ,
         \15533 , \15534 , \15535 , \15536 , \15537 , \15538 , \15539 , \15540 , \15541 , \15542 ,
         \15543 , \15544 , \15545 , \15546 , \15547 , \15548 , \15549 , \15550 , \15551 , \15552 ,
         \15553 , \15554 , \15555 , \15556 , \15557 , \15558 , \15559 , \15560 , \15561 , \15562 ,
         \15563 , \15564 , \15565 , \15566 , \15567 , \15568 , \15569 , \15570 , \15571 , \15572 ,
         \15573 , \15574 , \15575 , \15576 , \15577 , \15578 , \15579 , \15580 , \15581 , \15582 ,
         \15583 , \15584 , \15585 , \15586 , \15587 , \15588 , \15589 , \15590 , \15591 , \15592 ,
         \15593 , \15594 , \15595 , \15596 , \15597 , \15598 , \15599 , \15600 , \15601 , \15602 ,
         \15603 , \15604 , \15605 , \15606 , \15607 , \15608 , \15609 , \15610 , \15611 , \15612 ,
         \15613 , \15614 , \15615 , \15616 , \15617 , \15618 , \15619 , \15620 , \15621 , \15622 ,
         \15623 , \15624 , \15625 , \15626 , \15627 , \15628 , \15629 , \15630 , \15631 , \15632 ,
         \15633 , \15634 , \15635 , \15636 , \15637 , \15638 , \15639 , \15640 , \15641 , \15642 ,
         \15643 , \15644 , \15645 , \15646 , \15647 , \15648 , \15649 , \15650 , \15651 , \15652 ,
         \15653 , \15654 , \15655 , \15656 , \15657 , \15658 , \15659 , \15660 , \15661 , \15662 ,
         \15663 , \15664 , \15665 , \15666 , \15667 , \15668 , \15669 , \15670 , \15671 , \15672 ,
         \15673 , \15674 , \15675 , \15676 , \15677 , \15678 , \15679 , \15680 , \15681 , \15682 ,
         \15683 , \15684 , \15685 , \15686 , \15687 , \15688 , \15689 , \15690 , \15691 , \15692 ,
         \15693 , \15694 , \15695 , \15696 , \15697 , \15698 , \15699 , \15700 , \15701 , \15702 ,
         \15703 , \15704 , \15705 , \15706 , \15707 , \15708 , \15709 , \15710 , \15711 , \15712 ,
         \15713 , \15714 , \15715 , \15716 , \15717 , \15718 , \15719 , \15720 , \15721 , \15722 ,
         \15723 , \15724 , \15725 , \15726 , \15727 , \15728 , \15729 , \15730 , \15731 , \15732 ,
         \15733 , \15734 , \15735 , \15736 , \15737 , \15738 , \15739 , \15740 , \15741 , \15742 ,
         \15743 , \15744 , \15745 , \15746 , \15747 , \15748 , \15749 , \15750 , \15751 , \15752 ,
         \15753 , \15754 , \15755 , \15756 , \15757 , \15758 , \15759 , \15760 , \15761 , \15762 ,
         \15763 , \15764 , \15765 , \15766 , \15767 , \15768 , \15769 , \15770 , \15771 , \15772 ,
         \15773 , \15774 , \15775 , \15776 , \15777 , \15778 , \15779 , \15780 , \15781 , \15782 ,
         \15783 , \15784 , \15785 , \15786 , \15787 , \15788 , \15789 , \15790 , \15791 , \15792 ,
         \15793 , \15794 , \15795 , \15796 , \15797 , \15798 , \15799 , \15800 , \15801 , \15802 ,
         \15803 , \15804 , \15805 , \15806 , \15807 , \15808 , \15809 , \15810 , \15811 , \15812 ,
         \15813 , \15814 , \15815 , \15816 , \15817 , \15818 , \15819 , \15820 , \15821 , \15822 ,
         \15823 , \15824 , \15825 , \15826 , \15827 , \15828 , \15829 , \15830 , \15831 , \15832 ,
         \15833 , \15834 , \15835 , \15836 , \15837 , \15838 , \15839 , \15840 , \15841 , \15842 ,
         \15843 , \15844 , \15845 , \15846 , \15847 , \15848 , \15849 , \15850 , \15851 , \15852 ,
         \15853 , \15854 , \15855 , \15856 , \15857 , \15858 , \15859 , \15860 , \15861 , \15862 ,
         \15863 , \15864 , \15865 , \15866 , \15867 , \15868 , \15869 , \15870 , \15871 , \15872 ,
         \15873 , \15874 , \15875 , \15876 , \15877 , \15878 , \15879 , \15880 , \15881 , \15882 ,
         \15883 , \15884 , \15885 , \15886 , \15887 , \15888 , \15889 , \15890 , \15891 , \15892 ,
         \15893 , \15894 , \15895 , \15896 , \15897 , \15898 , \15899 , \15900 , \15901 , \15902 ,
         \15903 , \15904 , \15905 , \15906 , \15907 , \15908 , \15909 , \15910 , \15911 , \15912 ,
         \15913 , \15914 , \15915 , \15916 , \15917 , \15918 , \15919 , \15920 , \15921 , \15922 ,
         \15923 , \15924 , \15925 , \15926 , \15927 , \15928 , \15929 , \15930 , \15931 , \15932 ,
         \15933 , \15934 , \15935 , \15936 , \15937 , \15938 , \15939 , \15940 , \15941 , \15942 ,
         \15943 , \15944 , \15945 , \15946 , \15947 , \15948 , \15949 , \15950 , \15951 , \15952 ,
         \15953 , \15954 , \15955 , \15956 , \15957 , \15958 , \15959 , \15960 , \15961 , \15962 ,
         \15963 , \15964 , \15965 , \15966 , \15967 , \15968 , \15969 , \15970 , \15971 , \15972 ,
         \15973 , \15974 , \15975 , \15976 , \15977 , \15978 , \15979 , \15980 , \15981 , \15982 ,
         \15983 , \15984 , \15985 , \15986 , \15987 , \15988 , \15989 , \15990 , \15991 , \15992 ,
         \15993 , \15994 , \15995 , \15996 , \15997 , \15998 , \15999 , \16000 , \16001 , \16002 ,
         \16003 , \16004 , \16005 , \16006 , \16007 , \16008 , \16009 , \16010 , \16011 , \16012 ,
         \16013 , \16014 , \16015 , \16016 , \16017 , \16018 , \16019 , \16020 , \16021 , \16022 ,
         \16023 , \16024 , \16025 , \16026 , \16027 , \16028 , \16029 , \16030 , \16031 , \16032 ,
         \16033 , \16034 , \16035 , \16036 , \16037 , \16038 , \16039 , \16040 , \16041 , \16042 ,
         \16043 , \16044 , \16045 , \16046 , \16047 , \16048 , \16049 , \16050 , \16051 , \16052 ,
         \16053 , \16054 , \16055 , \16056 , \16057 , \16058 , \16059 , \16060 , \16061 , \16062 ,
         \16063 , \16064 , \16065 , \16066 , \16067 , \16068 , \16069 , \16070 , \16071 , \16072 ,
         \16073 , \16074 , \16075 , \16076 , \16077 , \16078 , \16079 , \16080 , \16081 , \16082 ,
         \16083 , \16084 , \16085 , \16086 , \16087 , \16088 , \16089 , \16090 , \16091 , \16092 ,
         \16093 , \16094 , \16095 , \16096 , \16097 , \16098 , \16099 , \16100 , \16101 , \16102 ,
         \16103 , \16104 , \16105 , \16106 , \16107 , \16108 , \16109 , \16110 , \16111 , \16112 ,
         \16113 , \16114 , \16115 , \16116 , \16117 , \16118 , \16119 , \16120 , \16121 , \16122 ,
         \16123 , \16124 , \16125 , \16126 , \16127 , \16128 , \16129 , \16130 , \16131 , \16132 ,
         \16133 , \16134 , \16135 , \16136 , \16137 , \16138 , \16139 , \16140 , \16141 , \16142 ,
         \16143 , \16144 , \16145 , \16146 , \16147 , \16148 , \16149 , \16150 , \16151 , \16152 ,
         \16153 , \16154 , \16155 , \16156 , \16157 , \16158 , \16159 , \16160 , \16161 , \16162 ,
         \16163 , \16164 , \16165 , \16166 , \16167 , \16168 , \16169 , \16170 , \16171 , \16172 ,
         \16173 , \16174 , \16175 , \16176 , \16177 , \16178 , \16179 , \16180 , \16181 , \16182 ,
         \16183 , \16184 , \16185 , \16186 , \16187 , \16188 , \16189 , \16190 , \16191 , \16192 ,
         \16193 , \16194 , \16195 , \16196 , \16197 , \16198 , \16199 , \16200 , \16201 , \16202 ,
         \16203 , \16204 , \16205 , \16206 , \16207 , \16208 , \16209 , \16210 , \16211 , \16212 ,
         \16213 , \16214 , \16215 , \16216 , \16217 , \16218 , \16219 , \16220 , \16221 , \16222 ,
         \16223 , \16224 , \16225 , \16226 , \16227 , \16228 , \16229 , \16230 , \16231 , \16232 ,
         \16233 , \16234 , \16235 , \16236 , \16237 , \16238 , \16239 , \16240 , \16241 , \16242 ,
         \16243 , \16244 , \16245 , \16246 , \16247 , \16248 , \16249 , \16250 , \16251 , \16252 ,
         \16253 , \16254 , \16255 , \16256 , \16257 , \16258 , \16259 , \16260 , \16261 , \16262 ,
         \16263 , \16264 , \16265 , \16266 , \16267 , \16268 , \16269 , \16270 , \16271 , \16272 ,
         \16273 , \16274 , \16275 , \16276 , \16277 , \16278 , \16279 , \16280 , \16281 , \16282 ,
         \16283 , \16284 , \16285 , \16286 , \16287 , \16288 , \16289 , \16290 , \16291 , \16292 ,
         \16293 , \16294 , \16295 , \16296 , \16297 , \16298 , \16299 , \16300 , \16301 , \16302 ,
         \16303 , \16304 , \16305 , \16306 , \16307 , \16308 , \16309 , \16310 , \16311 , \16312 ,
         \16313 , \16314 , \16315 , \16316 , \16317 , \16318 , \16319 , \16320 , \16321 , \16322 ,
         \16323 , \16324 , \16325 , \16326 , \16327 , \16328 , \16329 , \16330 , \16331 , \16332 ,
         \16333 , \16334 , \16335 , \16336 , \16337 , \16338 , \16339 , \16340 , \16341 , \16342 ,
         \16343 , \16344 , \16345 , \16346 , \16347 , \16348 , \16349 , \16350 , \16351 , \16352 ,
         \16353 , \16354 , \16355 , \16356 , \16357 , \16358 , \16359 , \16360 , \16361 , \16362 ,
         \16363 , \16364 , \16365 , \16366 , \16367 , \16368 , \16369 , \16370 , \16371 , \16372 ,
         \16373 , \16374 , \16375 , \16376 , \16377 , \16378 , \16379 , \16380 , \16381 , \16382 ,
         \16383 , \16384 , \16385 , \16386 , \16387 , \16388 , \16389 , \16390 , \16391 , \16392 ,
         \16393 , \16394 , \16395 , \16396 , \16397 , \16398 , \16399 , \16400 , \16401 , \16402 ,
         \16403 , \16404 , \16405 , \16406 , \16407 , \16408 , \16409 , \16410 , \16411 , \16412 ,
         \16413 , \16414 , \16415 , \16416 , \16417 , \16418 , \16419 , \16420 , \16421 , \16422 ,
         \16423 , \16424 , \16425 , \16426 , \16427 , \16428 , \16429 , \16430 , \16431 , \16432 ,
         \16433 , \16434 , \16435 , \16436 , \16437 , \16438 , \16439 , \16440 , \16441 , \16442 ,
         \16443 , \16444 , \16445 , \16446 , \16447 , \16448 , \16449 , \16450 , \16451 , \16452 ,
         \16453 , \16454 , \16455 , \16456 , \16457 , \16458 , \16459 , \16460 , \16461 , \16462 ,
         \16463 , \16464 , \16465 , \16466 , \16467 , \16468 , \16469 , \16470 , \16471 , \16472 ,
         \16473 , \16474 , \16475 , \16476 , \16477 , \16478 , \16479 , \16480 , \16481 , \16482 ,
         \16483 , \16484 , \16485 , \16486 , \16487 , \16488 , \16489 , \16490 , \16491 , \16492 ,
         \16493 , \16494 , \16495 , \16496 , \16497 , \16498 , \16499 , \16500 , \16501 , \16502 ,
         \16503 , \16504 , \16505 , \16506 , \16507 , \16508 , \16509 , \16510 , \16511 , \16512 ,
         \16513 , \16514 , \16515 , \16516 , \16517 , \16518 , \16519 , \16520 , \16521 , \16522 ,
         \16523 , \16524 , \16525 , \16526 , \16527 , \16528 , \16529 , \16530 , \16531 , \16532 ,
         \16533 , \16534 , \16535 , \16536 , \16537 , \16538 , \16539 , \16540 , \16541 , \16542 ,
         \16543 , \16544 , \16545 , \16546 , \16547 , \16548 , \16549 , \16550 , \16551 , \16552 ,
         \16553 , \16554 , \16555 , \16556 , \16557 , \16558 , \16559 , \16560 , \16561 , \16562 ,
         \16563 , \16564 , \16565 , \16566 , \16567 , \16568 , \16569 , \16570 , \16571 , \16572 ,
         \16573 , \16574 , \16575 , \16576 , \16577 , \16578 , \16579 , \16580 , \16581 , \16582 ,
         \16583 , \16584 , \16585 , \16586 , \16587 , \16588 , \16589 , \16590 , \16591 , \16592 ,
         \16593 , \16594 , \16595 , \16596 , \16597 , \16598 , \16599 , \16600 , \16601 , \16602 ,
         \16603 , \16604 , \16605 , \16606 , \16607 , \16608 , \16609 , \16610 , \16611 , \16612 ,
         \16613 , \16614 , \16615 , \16616 , \16617 , \16618 , \16619 , \16620 , \16621 , \16622 ,
         \16623 , \16624 , \16625 , \16626 , \16627 , \16628 , \16629 , \16630 , \16631 , \16632 ,
         \16633 , \16634 , \16635 , \16636 , \16637 , \16638 , \16639 , \16640 , \16641 , \16642 ,
         \16643 , \16644 , \16645 , \16646 , \16647 , \16648 , \16649 , \16650 , \16651 , \16652 ,
         \16653 , \16654 , \16655 , \16656 , \16657 , \16658 , \16659 , \16660 , \16661 , \16662 ,
         \16663 , \16664 , \16665 , \16666 , \16667 , \16668 , \16669 , \16670 , \16671 , \16672 ,
         \16673 , \16674 , \16675 , \16676 , \16677 , \16678 , \16679 , \16680 , \16681 , \16682 ,
         \16683 , \16684 , \16685 , \16686 , \16687 , \16688 , \16689 , \16690 , \16691 , \16692 ,
         \16693 , \16694 , \16695 , \16696 , \16697 , \16698 , \16699 , \16700 , \16701 , \16702 ,
         \16703 , \16704 , \16705 , \16706 , \16707 , \16708 , \16709 , \16710 , \16711 , \16712 ,
         \16713 , \16714 , \16715 , \16716 , \16717 , \16718 , \16719 , \16720 , \16721 , \16722 ,
         \16723 , \16724 , \16725 , \16726 , \16727 , \16728 , \16729 , \16730 , \16731 , \16732 ,
         \16733 , \16734 , \16735 , \16736 , \16737 , \16738 , \16739 , \16740 , \16741 , \16742 ,
         \16743 , \16744 , \16745 , \16746 , \16747 , \16748 , \16749 , \16750 , \16751 , \16752 ,
         \16753 , \16754 , \16755 , \16756 , \16757 , \16758 , \16759 , \16760 , \16761 , \16762 ,
         \16763 , \16764 , \16765 , \16766 , \16767 , \16768 , \16769 , \16770 , \16771 , \16772 ,
         \16773 , \16774 , \16775 , \16776 , \16777 , \16778 , \16779 , \16780 , \16781 , \16782 ,
         \16783 , \16784 , \16785 , \16786 , \16787 , \16788 , \16789 , \16790 , \16791 , \16792 ,
         \16793 , \16794 , \16795 , \16796 , \16797 , \16798 , \16799 , \16800 , \16801 , \16802 ,
         \16803 , \16804 , \16805 , \16806 , \16807 , \16808 , \16809 , \16810 , \16811 , \16812 ,
         \16813 , \16814 , \16815 , \16816 , \16817 , \16818 , \16819 , \16820 , \16821 , \16822 ,
         \16823 , \16824 , \16825 , \16826 , \16827 , \16828 , \16829 , \16830 , \16831 , \16832 ,
         \16833 , \16834 , \16835 , \16836 , \16837 , \16838 , \16839 , \16840 , \16841 , \16842 ,
         \16843 , \16844 , \16845 , \16846 , \16847 , \16848 , \16849 , \16850 , \16851 , \16852 ,
         \16853 , \16854 , \16855 , \16856 , \16857 , \16858 , \16859 , \16860 , \16861 , \16862 ,
         \16863 , \16864 , \16865 , \16866 , \16867 , \16868 , \16869 , \16870 , \16871 , \16872 ,
         \16873 , \16874 , \16875 , \16876 , \16877 , \16878 , \16879 , \16880 , \16881 , \16882 ,
         \16883 , \16884 , \16885 , \16886 , \16887 , \16888 , \16889 , \16890 , \16891 , \16892 ,
         \16893 , \16894 , \16895 , \16896 , \16897 , \16898 , \16899 , \16900 , \16901 , \16902 ,
         \16903 , \16904 , \16905 , \16906 , \16907 , \16908 , \16909 , \16910 , \16911 , \16912 ,
         \16913 , \16914 , \16915 , \16916 , \16917 , \16918 , \16919 , \16920 , \16921 , \16922 ,
         \16923 , \16924 , \16925 , \16926 , \16927 , \16928 , \16929 , \16930 , \16931 , \16932 ,
         \16933 , \16934 , \16935 , \16936 , \16937 , \16938 , \16939 , \16940 , \16941 , \16942 ,
         \16943 , \16944 , \16945 , \16946 , \16947 , \16948 , \16949 , \16950 , \16951 , \16952 ,
         \16953 , \16954 , \16955 , \16956 , \16957 , \16958 , \16959 , \16960 , \16961 , \16962 ,
         \16963 , \16964 , \16965 , \16966 , \16967 , \16968 , \16969 , \16970 , \16971 , \16972 ,
         \16973 , \16974 , \16975 , \16976 , \16977 , \16978 , \16979 , \16980 , \16981 , \16982 ,
         \16983 , \16984 , \16985 , \16986 , \16987 , \16988 , \16989 , \16990 , \16991 , \16992 ,
         \16993 , \16994 , \16995 , \16996 , \16997 , \16998 , \16999 , \17000 , \17001 , \17002 ,
         \17003 , \17004 , \17005 , \17006 , \17007 , \17008 , \17009 , \17010 , \17011 , \17012 ,
         \17013 , \17014 , \17015 , \17016 , \17017 , \17018 , \17019 , \17020 , \17021 , \17022 ,
         \17023 , \17024 , \17025 , \17026 , \17027 , \17028 , \17029 , \17030 , \17031 , \17032 ,
         \17033 , \17034 , \17035 , \17036 , \17037 , \17038 , \17039 , \17040 , \17041 , \17042 ,
         \17043 , \17044 , \17045 , \17046 , \17047 , \17048 , \17049 , \17050 , \17051 , \17052 ,
         \17053 , \17054 , \17055 , \17056 , \17057 , \17058 , \17059 , \17060 , \17061 , \17062 ,
         \17063 , \17064 , \17065 , \17066 , \17067 , \17068 , \17069 , \17070 , \17071 , \17072 ,
         \17073 , \17074 , \17075 , \17076 , \17077 , \17078 , \17079 , \17080 , \17081 , \17082 ,
         \17083 , \17084 , \17085 , \17086 , \17087 , \17088 , \17089 , \17090 , \17091 , \17092 ,
         \17093 , \17094 , \17095 , \17096 , \17097 , \17098 , \17099 , \17100 , \17101 , \17102 ,
         \17103 , \17104 , \17105 , \17106 , \17107 , \17108 , \17109 , \17110 , \17111 , \17112 ,
         \17113 , \17114 , \17115 , \17116 , \17117 , \17118 , \17119 , \17120 , \17121 , \17122 ,
         \17123 , \17124 , \17125 , \17126 , \17127 , \17128 , \17129 , \17130 , \17131 , \17132 ,
         \17133 , \17134 , \17135 , \17136 , \17137 , \17138 , \17139 , \17140 , \17141 , \17142 ,
         \17143 , \17144 , \17145 , \17146 , \17147 , \17148 , \17149 , \17150 , \17151 , \17152 ,
         \17153 , \17154 , \17155 , \17156 , \17157 , \17158 , \17159 , \17160 , \17161 , \17162 ,
         \17163 , \17164 , \17165 , \17166 , \17167 , \17168 , \17169 , \17170 , \17171 , \17172 ,
         \17173 , \17174 , \17175 , \17176 , \17177 , \17178 , \17179 , \17180 , \17181 , \17182 ,
         \17183 , \17184 , \17185 , \17186 , \17187 , \17188 , \17189 , \17190 , \17191 , \17192 ,
         \17193 , \17194 , \17195 , \17196 , \17197 , \17198 , \17199 , \17200 , \17201 , \17202 ,
         \17203 , \17204 , \17205 , \17206 , \17207 , \17208 , \17209 , \17210 , \17211 , \17212 ,
         \17213 , \17214 , \17215 , \17216 , \17217 , \17218 , \17219 , \17220 , \17221 , \17222 ,
         \17223 , \17224 , \17225 , \17226 , \17227 , \17228 , \17229 , \17230 , \17231 , \17232 ,
         \17233 , \17234 , \17235 , \17236 , \17237 , \17238 , \17239 , \17240 , \17241 , \17242 ,
         \17243 , \17244 , \17245 , \17246 , \17247 , \17248 , \17249 , \17250 , \17251 , \17252 ,
         \17253 , \17254 , \17255 , \17256 , \17257 , \17258 , \17259 , \17260 , \17261 , \17262 ,
         \17263 , \17264 , \17265 , \17266 , \17267 , \17268 , \17269 , \17270 , \17271 , \17272 ,
         \17273 , \17274 , \17275 , \17276 , \17277 , \17278 , \17279 , \17280 , \17281 , \17282 ,
         \17283 , \17284 , \17285 , \17286 , \17287 , \17288 , \17289 , \17290 , \17291 , \17292 ,
         \17293 , \17294 , \17295 , \17296 , \17297 , \17298 , \17299 , \17300 , \17301 , \17302 ,
         \17303 , \17304 , \17305 , \17306 , \17307 , \17308 , \17309 , \17310 , \17311 , \17312 ,
         \17313 , \17314 , \17315 , \17316 , \17317 , \17318 , \17319 , \17320 , \17321 , \17322 ,
         \17323 , \17324 , \17325 , \17326 , \17327 , \17328 , \17329 , \17330 , \17331 , \17332 ,
         \17333 , \17334 , \17335 , \17336 , \17337 , \17338 , \17339 , \17340 , \17341 , \17342 ,
         \17343 , \17344 , \17345 , \17346 , \17347 , \17348 , \17349 , \17350 , \17351 , \17352 ,
         \17353 , \17354 , \17355 , \17356 , \17357 , \17358 , \17359 , \17360 , \17361 , \17362 ,
         \17363 , \17364 , \17365 , \17366 , \17367 , \17368 , \17369 , \17370 , \17371 , \17372 ,
         \17373 , \17374 , \17375 , \17376 , \17377 , \17378 , \17379 , \17380 , \17381 , \17382 ,
         \17383 , \17384 , \17385 , \17386 , \17387 , \17388 , \17389 , \17390 , \17391 , \17392 ,
         \17393 , \17394 , \17395 , \17396 , \17397 , \17398 , \17399 , \17400 , \17401 , \17402 ,
         \17403 , \17404 , \17405 , \17406 , \17407 , \17408 , \17409 , \17410 , \17411 , \17412 ,
         \17413 , \17414 , \17415 , \17416 , \17417 , \17418 , \17419 , \17420 , \17421 , \17422 ,
         \17423 , \17424 , \17425 , \17426 , \17427 , \17428 , \17429 , \17430 , \17431 , \17432 ,
         \17433 , \17434 , \17435 , \17436 , \17437 , \17438 , \17439 , \17440 , \17441 , \17442 ,
         \17443 , \17444 , \17445 , \17446 , \17447 , \17448 , \17449 , \17450 , \17451 , \17452 ,
         \17453 , \17454 , \17455 , \17456 , \17457 , \17458 , \17459 , \17460 , \17461 , \17462 ,
         \17463 , \17464 , \17465 , \17466 , \17467 , \17468 , \17469 , \17470 , \17471 , \17472 ,
         \17473 , \17474 , \17475 , \17476 , \17477 , \17478 , \17479 , \17480 , \17481 , \17482 ,
         \17483 , \17484 , \17485 , \17486 , \17487 , \17488 , \17489 , \17490 , \17491 , \17492 ,
         \17493 , \17494 , \17495 , \17496 , \17497 , \17498 , \17499 , \17500 , \17501 , \17502 ,
         \17503 , \17504 , \17505 , \17506 , \17507 , \17508 , \17509 , \17510 , \17511 , \17512 ,
         \17513 , \17514 , \17515 , \17516 , \17517 , \17518 , \17519 , \17520 , \17521 , \17522 ,
         \17523 , \17524 , \17525 , \17526 , \17527 , \17528 , \17529 , \17530 , \17531 , \17532 ,
         \17533 , \17534 , \17535 , \17536 , \17537 , \17538 , \17539 , \17540 , \17541 , \17542 ,
         \17543 , \17544 , \17545 , \17546 , \17547 , \17548 , \17549 , \17550 , \17551 , \17552 ,
         \17553 , \17554 , \17555 , \17556 , \17557 , \17558 , \17559 , \17560 , \17561 , \17562 ,
         \17563 , \17564 , \17565 , \17566 , \17567 , \17568 , \17569 , \17570 , \17571 , \17572 ,
         \17573 , \17574 , \17575 , \17576 , \17577 , \17578 , \17579 , \17580 , \17581 , \17582 ,
         \17583 , \17584 , \17585 , \17586 , \17587 , \17588 , \17589 , \17590 , \17591 , \17592 ,
         \17593 , \17594 , \17595 , \17596 , \17597 , \17598 , \17599 , \17600 , \17601 , \17602 ,
         \17603 , \17604 , \17605 , \17606 , \17607 , \17608 , \17609 , \17610 , \17611 , \17612 ,
         \17613 , \17614 , \17615 , \17616 , \17617 , \17618 , \17619 , \17620 , \17621 , \17622 ,
         \17623 , \17624 , \17625 , \17626 , \17627 , \17628 , \17629 , \17630 , \17631 , \17632 ,
         \17633 , \17634 , \17635 , \17636 , \17637 , \17638 , \17639 , \17640 , \17641 , \17642 ,
         \17643 , \17644 , \17645 , \17646 , \17647 , \17648 , \17649 , \17650 , \17651 , \17652 ,
         \17653 , \17654 , \17655 , \17656 , \17657 , \17658 , \17659 , \17660 , \17661 , \17662 ,
         \17663 , \17664 , \17665 , \17666 , \17667 , \17668 , \17669 , \17670 , \17671 , \17672 ,
         \17673 , \17674 , \17675 , \17676 , \17677 , \17678 , \17679 , \17680 , \17681 , \17682 ,
         \17683 , \17684 , \17685 , \17686 , \17687 , \17688 , \17689 , \17690 , \17691 , \17692 ,
         \17693 , \17694 , \17695 , \17696 , \17697 , \17698 , \17699 , \17700 , \17701 , \17702 ,
         \17703 , \17704 , \17705 , \17706 , \17707 , \17708 , \17709 , \17710 , \17711 , \17712 ,
         \17713 , \17714 , \17715 , \17716 , \17717 , \17718 , \17719 , \17720 , \17721 , \17722 ,
         \17723 , \17724 , \17725 , \17726 , \17727 , \17728 , \17729 , \17730 , \17731 , \17732 ,
         \17733 , \17734 , \17735 , \17736 , \17737 , \17738 , \17739 , \17740 , \17741 , \17742 ,
         \17743 , \17744 , \17745 , \17746 , \17747 , \17748 , \17749 , \17750 , \17751 , \17752 ,
         \17753 , \17754 , \17755 , \17756 , \17757 , \17758 , \17759 , \17760 , \17761 , \17762 ,
         \17763 , \17764 , \17765 , \17766 , \17767 , \17768 , \17769 , \17770 , \17771 , \17772 ,
         \17773 , \17774 , \17775 , \17776 , \17777 , \17778 , \17779 , \17780 , \17781 , \17782 ,
         \17783 , \17784 , \17785 , \17786 , \17787 , \17788 , \17789 , \17790 , \17791 , \17792 ,
         \17793 , \17794 , \17795 , \17796 , \17797 , \17798 , \17799 , \17800 , \17801 , \17802 ,
         \17803 , \17804 , \17805 , \17806 , \17807 , \17808 , \17809 , \17810 , \17811 , \17812 ,
         \17813 , \17814 , \17815 , \17816 , \17817 , \17818 , \17819 , \17820 , \17821 , \17822 ,
         \17823 , \17824 , \17825 , \17826 , \17827 , \17828 , \17829 , \17830 , \17831 , \17832 ,
         \17833 , \17834 , \17835 , \17836 , \17837 , \17838 , \17839 , \17840 , \17841 , \17842 ,
         \17843 , \17844 , \17845 , \17846 , \17847 , \17848 , \17849 , \17850 , \17851 , \17852 ,
         \17853 , \17854 , \17855 , \17856 , \17857 , \17858 , \17859 , \17860 , \17861 , \17862 ,
         \17863 , \17864 , \17865 , \17866 , \17867 , \17868 , \17869 , \17870 , \17871 , \17872 ,
         \17873 , \17874 , \17875 , \17876 , \17877 , \17878 , \17879 , \17880 , \17881 , \17882 ,
         \17883 , \17884 , \17885 , \17886 , \17887 , \17888 , \17889 , \17890 , \17891 , \17892 ,
         \17893 , \17894 , \17895 , \17896 , \17897 , \17898 , \17899 , \17900 , \17901 , \17902 ,
         \17903 , \17904 , \17905 , \17906 , \17907 , \17908 , \17909 , \17910 , \17911 , \17912 ,
         \17913 , \17914 , \17915 , \17916 , \17917 , \17918 , \17919 , \17920 , \17921 , \17922 ,
         \17923 , \17924 , \17925 , \17926 , \17927 , \17928 , \17929 , \17930 , \17931 , \17932 ,
         \17933 , \17934 , \17935 , \17936 , \17937 , \17938 , \17939 , \17940 , \17941 , \17942 ,
         \17943 , \17944 , \17945 , \17946 , \17947 , \17948 , \17949 , \17950 , \17951 , \17952 ,
         \17953 , \17954 , \17955 , \17956 , \17957 , \17958 , \17959 , \17960 , \17961 , \17962 ,
         \17963 , \17964 , \17965 , \17966 , \17967 , \17968 , \17969 , \17970 , \17971 , \17972 ,
         \17973 , \17974 , \17975 , \17976 , \17977 , \17978 , \17979 , \17980 , \17981 , \17982 ,
         \17983 , \17984 , \17985 , \17986 , \17987 , \17988 , \17989 , \17990 , \17991 , \17992 ,
         \17993 , \17994 , \17995 , \17996 , \17997 , \17998 , \17999 , \18000 , \18001 , \18002 ,
         \18003 , \18004 , \18005 , \18006 , \18007 , \18008 , \18009 , \18010 , \18011 , \18012 ,
         \18013 , \18014 , \18015 , \18016 , \18017 , \18018 , \18019 , \18020 , \18021 , \18022 ,
         \18023 , \18024 , \18025 , \18026 , \18027 , \18028 , \18029 , \18030 , \18031 , \18032 ,
         \18033 , \18034 , \18035 , \18036 , \18037 , \18038 , \18039 , \18040 , \18041 , \18042 ,
         \18043 , \18044 , \18045 , \18046 , \18047 , \18048 , \18049 , \18050 , \18051 , \18052 ,
         \18053 , \18054 , \18055 , \18056 , \18057 , \18058 , \18059 , \18060 , \18061 , \18062 ,
         \18063 , \18064 , \18065 , \18066 , \18067 , \18068 , \18069 , \18070 , \18071 , \18072 ,
         \18073 , \18074 , \18075 , \18076 , \18077 , \18078 , \18079 , \18080 , \18081 , \18082 ,
         \18083 , \18084 , \18085 , \18086 , \18087 , \18088 , \18089 , \18090 , \18091 , \18092 ,
         \18093 , \18094 , \18095 , \18096 , \18097 , \18098 , \18099 , \18100 , \18101 , \18102 ,
         \18103 , \18104 , \18105 , \18106 , \18107 , \18108 , \18109 , \18110 , \18111 , \18112 ,
         \18113 , \18114 , \18115 , \18116 , \18117 , \18118 , \18119 , \18120 , \18121 , \18122 ,
         \18123 , \18124 , \18125 , \18126 , \18127 , \18128 , \18129 , \18130 , \18131 , \18132 ,
         \18133 , \18134 , \18135 , \18136 , \18137 , \18138 , \18139 , \18140 , \18141 , \18142 ,
         \18143 , \18144 , \18145 , \18146 , \18147 , \18148 , \18149 , \18150 , \18151 , \18152 ,
         \18153 , \18154 , \18155 , \18156 , \18157 , \18158 , \18159 , \18160 , \18161 , \18162 ,
         \18163 , \18164 , \18165 , \18166 , \18167 , \18168 , \18169 , \18170 , \18171 , \18172 ,
         \18173 , \18174 , \18175 , \18176 , \18177 , \18178 , \18179 , \18180 , \18181 , \18182 ,
         \18183 , \18184 , \18185 , \18186 , \18187 , \18188 , \18189 , \18190 , \18191 , \18192 ,
         \18193 , \18194 , \18195 , \18196 , \18197 , \18198 , \18199 , \18200 , \18201 , \18202 ,
         \18203 , \18204 , \18205 , \18206 , \18207 , \18208 , \18209 , \18210 , \18211 , \18212 ,
         \18213 , \18214 , \18215 , \18216 , \18217 , \18218 , \18219 , \18220 , \18221 , \18222 ,
         \18223 , \18224 , \18225 , \18226 , \18227 , \18228 , \18229 , \18230 , \18231 , \18232 ,
         \18233 , \18234 , \18235 , \18236 , \18237 , \18238 , \18239 , \18240 , \18241 , \18242 ,
         \18243 , \18244 , \18245 , \18246 , \18247 , \18248 , \18249 , \18250 , \18251 , \18252 ,
         \18253 , \18254 , \18255 , \18256 , \18257 , \18258 , \18259 , \18260 , \18261 , \18262 ,
         \18263 , \18264 , \18265 , \18266 , \18267 , \18268 , \18269 , \18270 , \18271 , \18272 ,
         \18273 , \18274 , \18275 , \18276 , \18277 , \18278 , \18279 , \18280 , \18281 , \18282 ,
         \18283 , \18284 , \18285 , \18286 , \18287 , \18288 , \18289 , \18290 , \18291 , \18292 ,
         \18293 , \18294 , \18295 , \18296 , \18297 , \18298 , \18299 , \18300 , \18301 , \18302 ,
         \18303 , \18304 , \18305 , \18306 , \18307 , \18308 , \18309 , \18310 , \18311 , \18312 ,
         \18313 , \18314 , \18315 , \18316 , \18317 , \18318 , \18319 , \18320 , \18321 , \18322 ,
         \18323 , \18324 , \18325 , \18326 , \18327 , \18328 , \18329 , \18330 , \18331 , \18332 ,
         \18333 , \18334 , \18335 , \18336 , \18337 , \18338 , \18339 , \18340 , \18341 , \18342 ,
         \18343 , \18344 , \18345 , \18346 , \18347 , \18348 , \18349 , \18350 , \18351 , \18352 ,
         \18353 , \18354 , \18355 , \18356 , \18357 , \18358 , \18359 , \18360 , \18361 , \18362 ,
         \18363 , \18364 , \18365 , \18366 , \18367 , \18368 , \18369 , \18370 , \18371 , \18372 ,
         \18373 , \18374 , \18375 , \18376 , \18377 , \18378 , \18379 , \18380 , \18381 , \18382 ,
         \18383 , \18384 , \18385 , \18386 , \18387 , \18388 , \18389 , \18390 , \18391 , \18392 ,
         \18393 , \18394 , \18395 , \18396 , \18397 , \18398 , \18399 , \18400 , \18401 , \18402 ,
         \18403 , \18404 , \18405 , \18406 , \18407 , \18408 , \18409 , \18410 , \18411 , \18412 ,
         \18413 , \18414 , \18415 , \18416 , \18417 , \18418 , \18419 , \18420 , \18421 , \18422 ,
         \18423 , \18424 , \18425 , \18426 , \18427 , \18428 , \18429 , \18430 , \18431 , \18432 ,
         \18433 , \18434 , \18435 , \18436 , \18437 , \18438 , \18439 , \18440 , \18441 , \18442 ,
         \18443 , \18444 , \18445 , \18446 , \18447 , \18448 , \18449 , \18450 , \18451 , \18452 ,
         \18453 , \18454 , \18455 , \18456 , \18457 , \18458 , \18459 , \18460 , \18461 , \18462 ,
         \18463 , \18464 , \18465 , \18466 , \18467 , \18468 , \18469 , \18470 , \18471 , \18472 ,
         \18473 , \18474 , \18475 , \18476 , \18477 , \18478 , \18479 , \18480 , \18481 , \18482 ,
         \18483 , \18484 , \18485 , \18486 , \18487 , \18488 , \18489 , \18490 , \18491 , \18492 ,
         \18493 , \18494 , \18495 , \18496 , \18497 , \18498 , \18499 , \18500 , \18501 , \18502 ,
         \18503 , \18504 , \18505 , \18506 , \18507 , \18508 , \18509 , \18510 , \18511 , \18512 ,
         \18513 , \18514 , \18515 , \18516 , \18517 , \18518 , \18519 , \18520 , \18521 , \18522 ,
         \18523 , \18524 , \18525 , \18526 , \18527 , \18528 , \18529 , \18530 , \18531 , \18532 ,
         \18533 , \18534 , \18535 , \18536 , \18537 , \18538 , \18539 , \18540 , \18541 , \18542 ,
         \18543 , \18544 , \18545 , \18546 , \18547 , \18548 , \18549 , \18550 , \18551 , \18552 ,
         \18553 , \18554 , \18555 , \18556 , \18557 , \18558 , \18559 , \18560 , \18561 , \18562 ,
         \18563 , \18564 , \18565 , \18566 , \18567 , \18568 , \18569 , \18570 , \18571 , \18572 ,
         \18573 , \18574 , \18575 , \18576 , \18577 , \18578 , \18579 , \18580 , \18581 , \18582 ,
         \18583 , \18584 , \18585 , \18586 , \18587 , \18588 , \18589 , \18590 , \18591 , \18592 ,
         \18593 , \18594 , \18595 , \18596 , \18597 , \18598 , \18599 , \18600 , \18601 , \18602 ,
         \18603 , \18604 , \18605 , \18606 , \18607 , \18608 , \18609 , \18610 , \18611 , \18612 ,
         \18613 , \18614 , \18615 , \18616 , \18617 , \18618 , \18619 , \18620 , \18621 , \18622 ,
         \18623 , \18624 , \18625 , \18626 , \18627 , \18628 , \18629 , \18630 , \18631 , \18632 ,
         \18633 , \18634 , \18635 , \18636 , \18637 , \18638 , \18639 , \18640 , \18641 , \18642 ,
         \18643 , \18644 , \18645 , \18646 , \18647 , \18648 , \18649 , \18650 , \18651 , \18652 ,
         \18653 , \18654 , \18655 , \18656 , \18657 , \18658 , \18659 , \18660 , \18661 , \18662 ,
         \18663 , \18664 , \18665 , \18666 , \18667 , \18668 , \18669 , \18670 , \18671 , \18672 ,
         \18673 , \18674 , \18675 , \18676 , \18677 , \18678 , \18679 , \18680 , \18681 , \18682 ,
         \18683 , \18684 , \18685 , \18686 , \18687 , \18688 , \18689 , \18690 , \18691 , \18692 ,
         \18693 , \18694 , \18695 , \18696 , \18697 , \18698 , \18699 , \18700 , \18701 , \18702 ,
         \18703 , \18704 , \18705 , \18706 , \18707 , \18708 , \18709 , \18710 , \18711 , \18712 ,
         \18713 , \18714 , \18715 , \18716 , \18717 , \18718 , \18719 , \18720 , \18721 , \18722 ,
         \18723 , \18724 , \18725 , \18726 , \18727 , \18728 , \18729 , \18730 , \18731 , \18732 ,
         \18733 , \18734 , \18735 , \18736 , \18737 , \18738 , \18739 , \18740 , \18741 , \18742 ,
         \18743 , \18744 , \18745 , \18746 , \18747 , \18748 , \18749 , \18750 , \18751 , \18752 ,
         \18753 , \18754 , \18755 , \18756 , \18757 , \18758 , \18759 , \18760 , \18761 , \18762 ,
         \18763 , \18764 , \18765 , \18766 , \18767 , \18768 , \18769 , \18770 , \18771 , \18772 ,
         \18773 , \18774 , \18775 , \18776 , \18777 , \18778 , \18779 , \18780 , \18781 , \18782 ,
         \18783 , \18784 , \18785 , \18786 , \18787 , \18788 , \18789 , \18790 , \18791 , \18792 ,
         \18793 , \18794 , \18795 , \18796 , \18797 , \18798 , \18799 , \18800 , \18801 , \18802 ,
         \18803 , \18804 , \18805 , \18806 , \18807 , \18808 , \18809 , \18810 , \18811 , \18812 ,
         \18813 , \18814 , \18815 , \18816 , \18817 , \18818 , \18819 , \18820 , \18821 , \18822 ,
         \18823 , \18824 , \18825 , \18826 , \18827 , \18828 , \18829 , \18830 , \18831 , \18832 ,
         \18833 , \18834 , \18835 , \18836 , \18837 , \18838 , \18839 , \18840 , \18841 , \18842 ,
         \18843 , \18844 , \18845 , \18846 , \18847 , \18848 , \18849 , \18850 , \18851 , \18852 ,
         \18853 , \18854 , \18855 , \18856 , \18857 , \18858 , \18859 , \18860 , \18861 , \18862 ,
         \18863 , \18864 , \18865 , \18866 , \18867 , \18868 , \18869 , \18870 , \18871 , \18872 ,
         \18873 , \18874 , \18875 , \18876 , \18877 , \18878 , \18879 , \18880 , \18881 , \18882 ,
         \18883 , \18884 , \18885 , \18886 , \18887 , \18888 , \18889 , \18890 , \18891 , \18892 ,
         \18893 , \18894 , \18895 , \18896 , \18897 , \18898 , \18899 , \18900 , \18901 , \18902 ,
         \18903 , \18904 , \18905 , \18906 , \18907 , \18908 , \18909 , \18910 , \18911 , \18912 ,
         \18913 , \18914 , \18915 , \18916 , \18917 , \18918 , \18919 , \18920 , \18921 , \18922 ,
         \18923 , \18924 , \18925 , \18926 , \18927 , \18928 , \18929 , \18930 , \18931 , \18932 ,
         \18933 , \18934 , \18935 , \18936 , \18937 , \18938 , \18939 , \18940 , \18941 , \18942 ,
         \18943 , \18944 , \18945 , \18946 , \18947 , \18948 , \18949 , \18950 , \18951 , \18952 ,
         \18953 , \18954 , \18955 , \18956 , \18957 , \18958 , \18959 , \18960 , \18961 , \18962 ,
         \18963 , \18964 , \18965 , \18966 , \18967 , \18968 , \18969 , \18970 , \18971 , \18972 ,
         \18973 , \18974 , \18975 , \18976 , \18977 , \18978 , \18979 , \18980 , \18981 , \18982 ,
         \18983 , \18984 , \18985 , \18986 , \18987 , \18988 , \18989 , \18990 , \18991 , \18992 ,
         \18993 , \18994 , \18995 , \18996 , \18997 , \18998 , \18999 , \19000 , \19001 , \19002 ,
         \19003 , \19004 , \19005 , \19006 , \19007 , \19008 , \19009 , \19010 , \19011 , \19012 ,
         \19013 , \19014 , \19015 , \19016 , \19017 , \19018 , \19019 , \19020 , \19021 , \19022 ,
         \19023 , \19024 , \19025 , \19026 , \19027 , \19028 , \19029 , \19030 , \19031 , \19032 ,
         \19033 , \19034 , \19035 , \19036 , \19037 , \19038 , \19039 , \19040 , \19041 , \19042 ,
         \19043 , \19044 , \19045 , \19046 , \19047 , \19048 , \19049 , \19050 , \19051 , \19052 ,
         \19053 , \19054 , \19055 , \19056 , \19057 , \19058 , \19059 , \19060 , \19061 , \19062 ,
         \19063 , \19064 , \19065 , \19066 , \19067 , \19068 , \19069 , \19070 , \19071 , \19072 ,
         \19073 , \19074 , \19075 , \19076 , \19077 , \19078 , \19079 , \19080 , \19081 , \19082 ,
         \19083 , \19084 , \19085 , \19086 , \19087 , \19088 , \19089 , \19090 , \19091 , \19092 ,
         \19093 , \19094 , \19095 , \19096 , \19097 , \19098 , \19099 , \19100 , \19101 , \19102 ,
         \19103 , \19104 , \19105 , \19106 , \19107 , \19108 , \19109 , \19110 , \19111 , \19112 ,
         \19113 , \19114 , \19115 , \19116 , \19117 , \19118 , \19119 , \19120 , \19121 , \19122 ,
         \19123 , \19124 , \19125 , \19126 , \19127 , \19128 , \19129 , \19130 , \19131 , \19132 ,
         \19133 , \19134 , \19135 , \19136 , \19137 , \19138 , \19139 , \19140 , \19141 , \19142 ,
         \19143 , \19144 , \19145 , \19146 , \19147 , \19148 , \19149 , \19150 , \19151 , \19152 ,
         \19153 , \19154 , \19155 , \19156 , \19157 , \19158 , \19159 , \19160 , \19161 , \19162 ,
         \19163 , \19164 , \19165 , \19166 , \19167 , \19168 , \19169 , \19170 , \19171 , \19172 ,
         \19173 , \19174 , \19175 , \19176 , \19177 , \19178 , \19179 , \19180 , \19181 , \19182 ,
         \19183 , \19184 , \19185 , \19186 , \19187 , \19188 , \19189 , \19190 , \19191 , \19192 ,
         \19193 , \19194 , \19195 , \19196 , \19197 , \19198 , \19199 , \19200 , \19201 , \19202 ,
         \19203 , \19204 , \19205 , \19206 , \19207 , \19208 , \19209 , \19210 , \19211 , \19212 ,
         \19213 , \19214 , \19215 , \19216 , \19217 , \19218 , \19219 , \19220 , \19221 , \19222 ,
         \19223 , \19224 , \19225 , \19226 , \19227 , \19228 , \19229 , \19230 , \19231 , \19232 ,
         \19233 , \19234 , \19235 , \19236 , \19237 , \19238 , \19239 , \19240 , \19241 , \19242 ,
         \19243 , \19244 , \19245 , \19246 , \19247 , \19248 , \19249 , \19250 , \19251 , \19252 ,
         \19253 , \19254 , \19255 , \19256 , \19257 , \19258 , \19259 , \19260 , \19261 , \19262 ,
         \19263 , \19264 , \19265 , \19266 , \19267 , \19268 , \19269 , \19270 , \19271 , \19272 ,
         \19273 , \19274 , \19275 , \19276 , \19277 , \19278 , \19279 , \19280 , \19281 , \19282 ,
         \19283 , \19284 , \19285 , \19286 , \19287 , \19288 , \19289 , \19290 , \19291 , \19292 ,
         \19293 , \19294 , \19295 , \19296 , \19297 , \19298 , \19299 , \19300 , \19301 , \19302 ,
         \19303 , \19304 , \19305 , \19306 , \19307 , \19308 , \19309 , \19310 , \19311 , \19312 ,
         \19313 , \19314 , \19315 , \19316 , \19317 , \19318 , \19319 , \19320 , \19321 , \19322 ,
         \19323 , \19324 , \19325 , \19326 , \19327 , \19328 , \19329 , \19330 , \19331 , \19332 ,
         \19333 , \19334 , \19335 , \19336 , \19337 , \19338 , \19339 , \19340 , \19341 , \19342 ,
         \19343 , \19344 , \19345 , \19346 , \19347 , \19348 , \19349 , \19350 , \19351 , \19352 ,
         \19353 , \19354 , \19355 , \19356 , \19357 , \19358 , \19359 , \19360 , \19361 , \19362 ,
         \19363 , \19364 , \19365 , \19366 , \19367 , \19368 , \19369 , \19370 , \19371 , \19372 ,
         \19373 , \19374 , \19375 , \19376 , \19377 , \19378 , \19379 , \19380 , \19381 , \19382 ,
         \19383 , \19384 , \19385 , \19386 , \19387 , \19388 , \19389 , \19390 , \19391 , \19392 ,
         \19393 , \19394 , \19395 , \19396 , \19397 , \19398 , \19399 , \19400 , \19401 , \19402 ,
         \19403 , \19404 , \19405 , \19406 , \19407 , \19408 , \19409 , \19410 , \19411 , \19412 ,
         \19413 , \19414 , \19415 , \19416 , \19417 , \19418 , \19419 , \19420 , \19421 , \19422 ,
         \19423 , \19424 , \19425 , \19426 , \19427 , \19428 , \19429 , \19430 , \19431 , \19432 ,
         \19433 , \19434 , \19435 , \19436 , \19437 , \19438 , \19439 , \19440 , \19441 , \19442 ,
         \19443 , \19444 , \19445 , \19446 , \19447 , \19448 , \19449 , \19450 , \19451 , \19452 ,
         \19453 , \19454 , \19455 , \19456 , \19457 , \19458 , \19459 , \19460 , \19461 , \19462 ,
         \19463 , \19464 , \19465 , \19466 , \19467 , \19468 , \19469 , \19470 , \19471 , \19472 ,
         \19473 , \19474 , \19475 , \19476 , \19477 , \19478 , \19479 , \19480 , \19481 , \19482 ,
         \19483 , \19484 , \19485 , \19486 , \19487 , \19488 , \19489 , \19490 , \19491 , \19492 ,
         \19493 , \19494 , \19495 , \19496 , \19497 , \19498 , \19499 , \19500 , \19501 , \19502 ,
         \19503 , \19504 , \19505 , \19506 , \19507 , \19508 , \19509 , \19510 , \19511 , \19512 ,
         \19513 , \19514 , \19515 , \19516 , \19517 , \19518 , \19519 , \19520 , \19521 , \19522 ,
         \19523 , \19524 , \19525 , \19526 , \19527 , \19528 , \19529 , \19530 , \19531 , \19532 ,
         \19533 , \19534 , \19535 , \19536 , \19537 , \19538 , \19539 , \19540 , \19541 , \19542 ,
         \19543 , \19544 , \19545 , \19546 , \19547 , \19548 , \19549 , \19550 , \19551 , \19552 ,
         \19553 , \19554 , \19555 , \19556 , \19557 , \19558 , \19559 , \19560 , \19561 , \19562 ,
         \19563 , \19564 , \19565 , \19566 , \19567 , \19568 , \19569 , \19570 , \19571 , \19572 ,
         \19573 , \19574 , \19575 , \19576 , \19577 , \19578 , \19579 , \19580 , \19581 , \19582 ,
         \19583 , \19584 , \19585 , \19586 , \19587 , \19588 , \19589 , \19590 , \19591 , \19592 ,
         \19593 , \19594 , \19595 , \19596 , \19597 , \19598 , \19599 , \19600 , \19601 , \19602 ,
         \19603 , \19604 , \19605 , \19606 , \19607 , \19608 , \19609 , \19610 , \19611 , \19612 ,
         \19613 , \19614 , \19615 , \19616 , \19617 , \19618 , \19619 , \19620 , \19621 , \19622 ,
         \19623 , \19624 , \19625 , \19626 , \19627 , \19628 , \19629 , \19630 , \19631 , \19632 ,
         \19633 , \19634 , \19635 , \19636 , \19637 , \19638 , \19639 , \19640 , \19641 , \19642 ,
         \19643 , \19644 , \19645 , \19646 , \19647 , \19648 , \19649 , \19650 , \19651 , \19652 ,
         \19653 , \19654 , \19655 , \19656 , \19657 , \19658 , \19659 , \19660 , \19661 , \19662 ,
         \19663 , \19664 , \19665 , \19666 , \19667 , \19668 , \19669 , \19670 , \19671 , \19672 ,
         \19673 , \19674 , \19675 , \19676 , \19677 , \19678 , \19679 , \19680 , \19681 , \19682 ,
         \19683 , \19684 , \19685 , \19686 , \19687 , \19688 , \19689 , \19690 , \19691 , \19692 ,
         \19693 , \19694 , \19695 , \19696 , \19697 , \19698 , \19699 , \19700 , \19701 , \19702 ,
         \19703 , \19704 , \19705 , \19706 , \19707 , \19708 , \19709 , \19710 , \19711 , \19712 ,
         \19713 , \19714 , \19715 , \19716 , \19717 , \19718 , \19719 , \19720 , \19721 , \19722 ,
         \19723 , \19724 , \19725 , \19726 , \19727 , \19728 , \19729 , \19730 , \19731 , \19732 ,
         \19733 , \19734 , \19735 , \19736 , \19737 , \19738 , \19739 , \19740 , \19741 , \19742 ,
         \19743 , \19744 , \19745 , \19746 , \19747 , \19748 , \19749 , \19750 , \19751 , \19752 ,
         \19753 , \19754 , \19755 , \19756 , \19757 , \19758 , \19759 , \19760 , \19761 , \19762 ,
         \19763 , \19764 , \19765 , \19766 , \19767 , \19768 , \19769 , \19770 , \19771 , \19772 ,
         \19773 , \19774 , \19775 , \19776 , \19777 , \19778 , \19779 , \19780 , \19781 , \19782 ,
         \19783 , \19784 , \19785 , \19786 , \19787 , \19788 , \19789 , \19790 , \19791 , \19792 ,
         \19793 , \19794 , \19795 , \19796 , \19797 , \19798 , \19799 , \19800 , \19801 , \19802 ,
         \19803 , \19804 , \19805 , \19806 , \19807 , \19808 , \19809 , \19810 , \19811 , \19812 ,
         \19813 , \19814 , \19815 , \19816 , \19817 , \19818 , \19819 , \19820 , \19821 , \19822 ,
         \19823 , \19824 , \19825 , \19826 , \19827 , \19828 , \19829 , \19830 , \19831 , \19832 ,
         \19833 , \19834 , \19835 , \19836 , \19837 , \19838 , \19839 , \19840 , \19841 , \19842 ,
         \19843 , \19844 , \19845 , \19846 , \19847 , \19848 , \19849 , \19850 , \19851 , \19852 ,
         \19853 , \19854 , \19855 , \19856 , \19857 , \19858 , \19859 , \19860 , \19861 , \19862 ,
         \19863 , \19864 , \19865 , \19866 , \19867 , \19868 , \19869 , \19870 , \19871 , \19872 ,
         \19873 , \19874 , \19875 , \19876 , \19877 , \19878 , \19879 , \19880 , \19881 , \19882 ,
         \19883 , \19884 , \19885 , \19886 , \19887 , \19888 , \19889 , \19890 , \19891 , \19892 ,
         \19893 , \19894 , \19895 , \19896 , \19897 , \19898 , \19899 , \19900 , \19901 , \19902 ,
         \19903 , \19904 , \19905 , \19906 , \19907 , \19908 , \19909 , \19910 , \19911 , \19912 ,
         \19913 , \19914 , \19915 , \19916 , \19917 , \19918 , \19919 , \19920 , \19921 , \19922 ,
         \19923 , \19924 , \19925 , \19926 , \19927 , \19928 , \19929 , \19930 , \19931 , \19932 ,
         \19933 , \19934 , \19935 , \19936 , \19937 , \19938 , \19939 , \19940 , \19941 , \19942 ,
         \19943 , \19944 , \19945 , \19946 , \19947 , \19948 , \19949 , \19950 , \19951 , \19952 ,
         \19953 , \19954 , \19955 , \19956 , \19957 , \19958 , \19959 , \19960 , \19961 , \19962 ,
         \19963 , \19964 , \19965 , \19966 , \19967 , \19968 , \19969 , \19970 , \19971 , \19972 ,
         \19973 , \19974 , \19975 , \19976 , \19977 , \19978 , \19979 , \19980 , \19981 , \19982 ,
         \19983 , \19984 , \19985 , \19986 , \19987 , \19988 , \19989 , \19990 , \19991 , \19992 ,
         \19993 , \19994 , \19995 , \19996 , \19997 , \19998 , \19999 , \20000 , \20001 , \20002 ,
         \20003 , \20004 , \20005 , \20006 , \20007 , \20008 , \20009 , \20010 , \20011 , \20012 ,
         \20013 , \20014 , \20015 , \20016 , \20017 , \20018 , \20019 , \20020 , \20021 , \20022 ,
         \20023 , \20024 , \20025 , \20026 , \20027 , \20028 , \20029 , \20030 , \20031 , \20032 ,
         \20033 , \20034 , \20035 , \20036 , \20037 , \20038 , \20039 , \20040 , \20041 , \20042 ,
         \20043 , \20044 , \20045 , \20046 , \20047 , \20048 , \20049 , \20050 , \20051 , \20052 ,
         \20053 , \20054 , \20055 , \20056 , \20057 , \20058 , \20059 , \20060 , \20061 , \20062 ,
         \20063 , \20064 , \20065 , \20066 , \20067 , \20068 , \20069 , \20070 , \20071 , \20072 ,
         \20073 , \20074 , \20075 , \20076 , \20077 , \20078 , \20079 , \20080 , \20081 , \20082 ,
         \20083 , \20084 , \20085 , \20086 , \20087 , \20088 , \20089 , \20090 , \20091 , \20092 ,
         \20093 , \20094 , \20095 , \20096 , \20097 , \20098 , \20099 , \20100 , \20101 , \20102 ,
         \20103 , \20104 , \20105 , \20106 , \20107 , \20108 , \20109 , \20110 , \20111 , \20112 ,
         \20113 , \20114 , \20115 , \20116 , \20117 , \20118 , \20119 , \20120 , \20121 , \20122 ,
         \20123 , \20124 , \20125 , \20126 , \20127 , \20128 , \20129 , \20130 , \20131 , \20132 ,
         \20133 , \20134 , \20135 , \20136 , \20137 , \20138 , \20139 , \20140 , \20141 , \20142 ,
         \20143 , \20144 , \20145 , \20146 , \20147 , \20148 , \20149 , \20150 , \20151 , \20152 ,
         \20153 , \20154 , \20155 , \20156 , \20157 , \20158 , \20159 , \20160 , \20161 , \20162 ,
         \20163 , \20164 , \20165 , \20166 , \20167 , \20168 , \20169 , \20170 , \20171 , \20172 ,
         \20173 , \20174 , \20175 , \20176 , \20177 , \20178 , \20179 , \20180 , \20181 , \20182 ,
         \20183 , \20184 , \20185 , \20186 , \20187 , \20188 , \20189 , \20190 , \20191 , \20192 ,
         \20193 , \20194 , \20195 , \20196 , \20197 , \20198 , \20199 , \20200 , \20201 , \20202 ,
         \20203 , \20204 , \20205 , \20206 , \20207 , \20208 , \20209 , \20210 , \20211 , \20212 ,
         \20213 , \20214 , \20215 , \20216 , \20217 , \20218 , \20219 , \20220 , \20221 , \20222 ,
         \20223 , \20224 , \20225 , \20226 , \20227 , \20228 , \20229 , \20230 , \20231 , \20232 ,
         \20233 , \20234 , \20235 , \20236 , \20237 , \20238 , \20239 , \20240 , \20241 , \20242 ,
         \20243 , \20244 , \20245 , \20246 , \20247 , \20248 , \20249 , \20250 , \20251 , \20252 ,
         \20253 , \20254 , \20255 , \20256 , \20257 , \20258 , \20259 , \20260 , \20261 , \20262 ,
         \20263 , \20264 , \20265 , \20266 , \20267 , \20268 , \20269 , \20270 , \20271 , \20272 ,
         \20273 , \20274 , \20275 , \20276 , \20277 , \20278 , \20279 , \20280 , \20281 , \20282 ,
         \20283 , \20284 , \20285 , \20286 , \20287 , \20288 , \20289 , \20290 , \20291 , \20292 ,
         \20293 , \20294 , \20295 , \20296 , \20297 , \20298 , \20299 , \20300 , \20301 , \20302 ,
         \20303 , \20304 , \20305 , \20306 , \20307 , \20308 , \20309 , \20310 , \20311 , \20312 ,
         \20313 , \20314 , \20315 , \20316 , \20317 , \20318 , \20319 , \20320 , \20321 , \20322 ,
         \20323 , \20324 , \20325 , \20326 , \20327 , \20328 , \20329 , \20330 , \20331 , \20332 ,
         \20333 , \20334 , \20335 , \20336 , \20337 , \20338 , \20339 , \20340 , \20341 , \20342 ,
         \20343 , \20344 , \20345 , \20346 , \20347 , \20348 , \20349 , \20350 , \20351 , \20352 ,
         \20353 , \20354 , \20355 , \20356 , \20357 , \20358 , \20359 , \20360 , \20361 , \20362 ,
         \20363 , \20364 , \20365 , \20366 , \20367 , \20368 , \20369 , \20370 , \20371 , \20372 ,
         \20373 , \20374 , \20375 , \20376 , \20377 , \20378 , \20379 , \20380 , \20381 , \20382 ,
         \20383 , \20384 , \20385 , \20386 , \20387 , \20388 , \20389 , \20390 , \20391 , \20392 ,
         \20393 , \20394 , \20395 , \20396 , \20397 , \20398 , \20399 , \20400 , \20401 , \20402 ,
         \20403 , \20404 , \20405 , \20406 , \20407 , \20408 , \20409 , \20410 , \20411 , \20412 ,
         \20413 , \20414 , \20415 , \20416 , \20417 , \20418 , \20419 , \20420 , \20421 , \20422 ,
         \20423 , \20424 , \20425 , \20426 , \20427 , \20428 , \20429 , \20430 , \20431 , \20432 ,
         \20433 , \20434 , \20435 , \20436 , \20437 , \20438 , \20439 , \20440 , \20441 , \20442 ,
         \20443 , \20444 , \20445 , \20446 , \20447 , \20448 , \20449 , \20450 , \20451 , \20452 ,
         \20453 , \20454 , \20455 , \20456 , \20457 , \20458 , \20459 , \20460 , \20461 , \20462 ,
         \20463 , \20464 , \20465 , \20466 , \20467 , \20468 , \20469 , \20470 , \20471 , \20472 ,
         \20473 , \20474 , \20475 , \20476 , \20477 , \20478 , \20479 , \20480 , \20481 , \20482 ,
         \20483 , \20484 , \20485 , \20486 , \20487 , \20488 , \20489 , \20490 , \20491 , \20492 ,
         \20493 , \20494 , \20495 , \20496 , \20497 , \20498 , \20499 , \20500 , \20501 , \20502 ,
         \20503 , \20504 , \20505 , \20506 , \20507 , \20508 , \20509 , \20510 , \20511 , \20512 ,
         \20513 , \20514 , \20515 , \20516 , \20517 , \20518 , \20519 , \20520 , \20521 , \20522 ,
         \20523 , \20524 , \20525 , \20526 , \20527 , \20528 , \20529 , \20530 , \20531 , \20532 ,
         \20533 , \20534 , \20535 , \20536 , \20537 , \20538 , \20539 , \20540 , \20541 , \20542 ,
         \20543 , \20544 , \20545 , \20546 , \20547 , \20548 , \20549 , \20550 , \20551 , \20552 ,
         \20553 , \20554 , \20555 , \20556 , \20557 , \20558 , \20559 , \20560 , \20561 , \20562 ,
         \20563 , \20564 , \20565 , \20566 , \20567 , \20568 , \20569 , \20570 , \20571 , \20572 ,
         \20573 , \20574 , \20575 , \20576 , \20577 , \20578 , \20579 , \20580 , \20581 , \20582 ,
         \20583 , \20584 , \20585 , \20586 , \20587 , \20588 , \20589 , \20590 , \20591 , \20592 ,
         \20593 , \20594 , \20595 , \20596 , \20597 , \20598 , \20599 , \20600 , \20601 , \20602 ,
         \20603 , \20604 , \20605 , \20606 , \20607 , \20608 , \20609 , \20610 , \20611 , \20612 ,
         \20613 , \20614 , \20615 , \20616 , \20617 , \20618 , \20619 , \20620 , \20621 , \20622 ,
         \20623 , \20624 , \20625 , \20626 , \20627 , \20628 , \20629 , \20630 , \20631 , \20632 ,
         \20633 , \20634 , \20635 , \20636 , \20637 , \20638 , \20639 , \20640 , \20641 , \20642 ,
         \20643 , \20644 , \20645 , \20646 , \20647 , \20648 , \20649 , \20650 , \20651 , \20652 ,
         \20653 , \20654 , \20655 , \20656 , \20657 , \20658 , \20659 , \20660 , \20661 , \20662 ,
         \20663 , \20664 , \20665 , \20666 , \20667 , \20668 , \20669 , \20670 , \20671 , \20672 ,
         \20673 , \20674 , \20675 , \20676 , \20677 , \20678 , \20679 , \20680 , \20681 , \20682 ,
         \20683 , \20684 , \20685 , \20686 , \20687 , \20688 , \20689 , \20690 , \20691 , \20692 ,
         \20693 , \20694 , \20695 , \20696 , \20697 , \20698 , \20699 , \20700 , \20701 , \20702 ,
         \20703 , \20704 , \20705 , \20706 , \20707 , \20708 , \20709 , \20710 , \20711 , \20712 ,
         \20713 , \20714 , \20715 , \20716 , \20717 , \20718 , \20719 , \20720 , \20721 , \20722 ,
         \20723 , \20724 , \20725 , \20726 , \20727 , \20728 , \20729 , \20730 , \20731 , \20732 ,
         \20733 , \20734 , \20735 , \20736 , \20737 , \20738 , \20739 , \20740 , \20741 , \20742 ,
         \20743 , \20744 , \20745 , \20746 , \20747 , \20748 , \20749 , \20750 , \20751 , \20752 ,
         \20753 , \20754 , \20755 , \20756 , \20757 , \20758 , \20759 , \20760 , \20761 , \20762 ,
         \20763 , \20764 , \20765 , \20766 , \20767 , \20768 , \20769 , \20770 , \20771 , \20772 ,
         \20773 , \20774 , \20775 , \20776 , \20777 , \20778 , \20779 , \20780 , \20781 , \20782 ,
         \20783 , \20784 , \20785 , \20786 , \20787 , \20788 , \20789 , \20790 , \20791 , \20792 ,
         \20793 , \20794 , \20795 , \20796 , \20797 , \20798 , \20799 , \20800 , \20801 , \20802 ,
         \20803 , \20804 , \20805 , \20806 , \20807 , \20808 , \20809 , \20810 , \20811 , \20812 ,
         \20813 , \20814 , \20815 , \20816 , \20817 , \20818 , \20819 , \20820 , \20821 , \20822 ,
         \20823 , \20824 , \20825 , \20826 , \20827 , \20828 , \20829 , \20830 , \20831 , \20832 ,
         \20833 , \20834 , \20835 , \20836 , \20837 , \20838 , \20839 , \20840 , \20841 , \20842 ,
         \20843 , \20844 , \20845 , \20846 , \20847 , \20848 , \20849 , \20850 , \20851 , \20852 ,
         \20853 , \20854 , \20855 , \20856 , \20857 , \20858 , \20859 , \20860 , \20861 , \20862 ,
         \20863 , \20864 , \20865 , \20866 , \20867 , \20868 , \20869 , \20870 , \20871 , \20872 ,
         \20873 , \20874 , \20875 , \20876 , \20877 , \20878 , \20879 , \20880 , \20881 , \20882 ,
         \20883 , \20884 , \20885 , \20886 , \20887 , \20888 , \20889 , \20890 , \20891 , \20892 ,
         \20893 , \20894 , \20895 , \20896 , \20897 , \20898 , \20899 , \20900 , \20901 , \20902 ,
         \20903 , \20904 , \20905 , \20906 , \20907 , \20908 , \20909 , \20910 , \20911 , \20912 ,
         \20913 , \20914 , \20915 , \20916 , \20917 , \20918 , \20919 , \20920 , \20921 , \20922 ,
         \20923 , \20924 , \20925 , \20926 , \20927 , \20928 , \20929 , \20930 , \20931 , \20932 ,
         \20933 , \20934 , \20935 , \20936 , \20937 , \20938 , \20939 , \20940 , \20941 , \20942 ,
         \20943 , \20944 , \20945 , \20946 , \20947 , \20948 , \20949 , \20950 , \20951 , \20952 ,
         \20953 , \20954 , \20955 , \20956 , \20957 , \20958 , \20959 , \20960 , \20961 , \20962 ,
         \20963 , \20964 , \20965 , \20966 , \20967 , \20968 , \20969 , \20970 , \20971 , \20972 ,
         \20973 , \20974 , \20975 , \20976 , \20977 , \20978 , \20979 , \20980 , \20981 , \20982 ,
         \20983 , \20984 , \20985 , \20986 , \20987 , \20988 , \20989 , \20990 , \20991 , \20992 ,
         \20993 , \20994 , \20995 , \20996 , \20997 , \20998 , \20999 , \21000 , \21001 , \21002 ,
         \21003 , \21004 , \21005 , \21006 , \21007 , \21008 , \21009 , \21010 , \21011 , \21012 ,
         \21013 , \21014 , \21015 , \21016 , \21017 , \21018 , \21019 , \21020 , \21021 , \21022 ,
         \21023 , \21024 , \21025 , \21026 , \21027 , \21028 , \21029 , \21030 , \21031 , \21032 ,
         \21033 , \21034 , \21035 , \21036 , \21037 , \21038 , \21039 , \21040 , \21041 , \21042 ,
         \21043 , \21044 , \21045 , \21046 , \21047 , \21048 , \21049 , \21050 , \21051 , \21052 ,
         \21053 , \21054 , \21055 , \21056 , \21057 , \21058 , \21059 , \21060 , \21061 , \21062 ,
         \21063 , \21064 , \21065 , \21066 , \21067 , \21068 , \21069 , \21070 , \21071 , \21072 ,
         \21073 , \21074 , \21075 , \21076 , \21077 , \21078 , \21079 , \21080 , \21081 , \21082 ,
         \21083 , \21084 , \21085 , \21086 , \21087 , \21088 , \21089 , \21090 , \21091 , \21092 ,
         \21093 , \21094 , \21095 , \21096 , \21097 , \21098 , \21099 , \21100 , \21101 , \21102 ,
         \21103 , \21104 , \21105 , \21106 , \21107 , \21108 , \21109 , \21110 , \21111 , \21112 ,
         \21113 , \21114 , \21115 , \21116 , \21117 , \21118 , \21119 , \21120 , \21121 , \21122 ,
         \21123 , \21124 , \21125 , \21126 , \21127 , \21128 , \21129 , \21130 , \21131 , \21132 ,
         \21133 , \21134 , \21135 , \21136 , \21137 , \21138 , \21139 , \21140 , \21141 , \21142 ,
         \21143 , \21144 , \21145 , \21146 , \21147 , \21148 , \21149 , \21150 , \21151 , \21152 ,
         \21153 , \21154 , \21155 , \21156 , \21157 , \21158 , \21159 , \21160 , \21161 , \21162 ,
         \21163 , \21164 , \21165 , \21166 , \21167 , \21168 , \21169 , \21170 , \21171 , \21172 ,
         \21173 , \21174 , \21175 , \21176 , \21177 , \21178 , \21179 , \21180 , \21181 , \21182 ,
         \21183 , \21184 , \21185 , \21186 , \21187 , \21188 , \21189 , \21190 , \21191 , \21192 ,
         \21193 , \21194 , \21195 , \21196 , \21197 , \21198 , \21199 , \21200 , \21201 , \21202 ,
         \21203 , \21204 , \21205 , \21206 , \21207 , \21208 , \21209 , \21210 , \21211 , \21212 ,
         \21213 , \21214 , \21215 , \21216 , \21217 , \21218 , \21219 , \21220 , \21221 , \21222 ,
         \21223 , \21224 , \21225 , \21226 , \21227 , \21228 , \21229 , \21230 , \21231 , \21232 ,
         \21233 , \21234 , \21235 , \21236 , \21237 , \21238 , \21239 , \21240 , \21241 , \21242 ,
         \21243 , \21244 , \21245 , \21246 , \21247 , \21248 , \21249 , \21250 , \21251 , \21252 ,
         \21253 , \21254 , \21255 , \21256 , \21257 , \21258 , \21259 , \21260 , \21261 , \21262 ,
         \21263 , \21264 , \21265 , \21266 , \21267 , \21268 , \21269 , \21270 , \21271 , \21272 ,
         \21273 , \21274 , \21275 , \21276 , \21277 , \21278 , \21279 , \21280 , \21281 , \21282 ,
         \21283 , \21284 , \21285 , \21286 , \21287 , \21288 , \21289 , \21290 , \21291 , \21292 ,
         \21293 , \21294 , \21295 , \21296 , \21297 , \21298 , \21299 , \21300 , \21301 , \21302 ,
         \21303 , \21304 , \21305 , \21306 , \21307 , \21308 , \21309 , \21310 , \21311 , \21312 ,
         \21313 , \21314 , \21315 , \21316 , \21317 , \21318 , \21319 , \21320 , \21321 , \21322 ,
         \21323 , \21324 , \21325 , \21326 , \21327 , \21328 , \21329 , \21330 , \21331 , \21332 ,
         \21333 , \21334 , \21335 , \21336 , \21337 , \21338 , \21339 , \21340 , \21341 , \21342 ,
         \21343 , \21344 , \21345 , \21346 , \21347 , \21348 , \21349 , \21350 , \21351 , \21352 ,
         \21353 , \21354 , \21355 , \21356 , \21357 , \21358 , \21359 , \21360 , \21361 , \21362 ,
         \21363 , \21364 , \21365 , \21366 , \21367 , \21368 , \21369 , \21370 , \21371 , \21372 ,
         \21373 , \21374 , \21375 , \21376 , \21377 , \21378 , \21379 , \21380 , \21381 , \21382 ,
         \21383 , \21384 , \21385 , \21386 , \21387 , \21388 , \21389 , \21390 , \21391 , \21392 ,
         \21393 , \21394 , \21395 , \21396 , \21397 , \21398 , \21399 , \21400 , \21401 , \21402 ,
         \21403 , \21404 , \21405 , \21406 , \21407 , \21408 , \21409 , \21410 , \21411 , \21412 ,
         \21413 , \21414 , \21415 , \21416 , \21417 , \21418 , \21419 , \21420 , \21421 , \21422 ,
         \21423 , \21424 , \21425 , \21426 , \21427 , \21428 , \21429 , \21430 , \21431 , \21432 ,
         \21433 , \21434 , \21435 , \21436 , \21437 , \21438 , \21439 , \21440 , \21441 , \21442 ,
         \21443 , \21444 , \21445 , \21446 , \21447 , \21448 , \21449 , \21450 , \21451 , \21452 ,
         \21453 , \21454 , \21455 , \21456 , \21457 , \21458 , \21459 , \21460 , \21461 , \21462 ,
         \21463 , \21464 , \21465 , \21466 , \21467 , \21468 , \21469 , \21470 , \21471 , \21472 ,
         \21473 , \21474 , \21475 , \21476 , \21477 , \21478 , \21479 , \21480 , \21481 , \21482 ,
         \21483 , \21484 , \21485 , \21486 , \21487 , \21488 , \21489 , \21490 , \21491 , \21492 ,
         \21493 , \21494 , \21495 , \21496 , \21497 , \21498 , \21499 , \21500 , \21501 , \21502 ,
         \21503 , \21504 , \21505 , \21506 , \21507 , \21508 , \21509 , \21510 , \21511 , \21512 ,
         \21513 , \21514 , \21515 , \21516 , \21517 , \21518 , \21519 , \21520 , \21521 , \21522 ,
         \21523 , \21524 , \21525 , \21526 , \21527 , \21528 , \21529 , \21530 , \21531 , \21532 ,
         \21533 , \21534 , \21535 , \21536 , \21537 , \21538 , \21539 , \21540 , \21541 , \21542 ,
         \21543 , \21544 , \21545 , \21546 , \21547 , \21548 , \21549 , \21550 , \21551 , \21552 ,
         \21553 , \21554 , \21555 , \21556 , \21557 , \21558 , \21559 , \21560 , \21561 , \21562 ,
         \21563 , \21564 , \21565 , \21566 , \21567 , \21568 , \21569 , \21570 , \21571 , \21572 ,
         \21573 , \21574 , \21575 , \21576 , \21577 , \21578 , \21579 , \21580 , \21581 , \21582 ,
         \21583 , \21584 , \21585 , \21586 , \21587 , \21588 , \21589 , \21590 , \21591 , \21592 ,
         \21593 , \21594 , \21595 , \21596 , \21597 , \21598 , \21599 , \21600 , \21601 , \21602 ,
         \21603 , \21604 , \21605 , \21606 , \21607 , \21608 , \21609 , \21610 , \21611 , \21612 ,
         \21613 , \21614 , \21615 , \21616 , \21617 , \21618 , \21619 , \21620 , \21621 , \21622 ,
         \21623 , \21624 , \21625 , \21626 , \21627 , \21628 , \21629 , \21630 , \21631 , \21632 ,
         \21633 , \21634 , \21635 , \21636 , \21637 , \21638 , \21639 , \21640 , \21641 , \21642 ,
         \21643 , \21644 , \21645 , \21646 , \21647 , \21648 , \21649 , \21650 , \21651 , \21652 ,
         \21653 , \21654 , \21655 , \21656 , \21657 , \21658 , \21659 , \21660 , \21661 , \21662 ,
         \21663 , \21664 , \21665 , \21666 , \21667 , \21668 , \21669 , \21670 , \21671 , \21672 ,
         \21673 , \21674 , \21675 , \21676 , \21677 , \21678 , \21679 , \21680 , \21681 , \21682 ,
         \21683 , \21684 , \21685 , \21686 , \21687 , \21688 , \21689 , \21690 , \21691 , \21692 ,
         \21693 , \21694 , \21695 , \21696 , \21697 , \21698 , \21699 , \21700 , \21701 , \21702 ,
         \21703 , \21704 , \21705 , \21706 , \21707 , \21708 , \21709 , \21710 , \21711 , \21712 ,
         \21713 , \21714 , \21715 , \21716 , \21717 , \21718 , \21719 , \21720 , \21721 , \21722 ,
         \21723 , \21724 , \21725 , \21726 , \21727 , \21728 , \21729 , \21730 , \21731 , \21732 ,
         \21733 , \21734 , \21735 , \21736 , \21737 , \21738 , \21739 , \21740 , \21741 , \21742 ,
         \21743 , \21744 , \21745 , \21746 , \21747 , \21748 , \21749 , \21750 , \21751 , \21752 ,
         \21753 , \21754 , \21755 , \21756 , \21757 , \21758 , \21759 , \21760 , \21761 , \21762 ,
         \21763 , \21764 , \21765 , \21766 , \21767 , \21768 , \21769 , \21770 , \21771 , \21772 ,
         \21773 , \21774 , \21775 , \21776 , \21777 , \21778 , \21779 , \21780 , \21781 , \21782 ,
         \21783 , \21784 , \21785 , \21786 , \21787 , \21788 , \21789 , \21790 , \21791 , \21792 ,
         \21793 , \21794 , \21795 , \21796 , \21797 , \21798 , \21799 , \21800 , \21801 , \21802 ,
         \21803 , \21804 , \21805 , \21806 , \21807 , \21808 , \21809 , \21810 , \21811 , \21812 ,
         \21813 , \21814 , \21815 , \21816 , \21817 , \21818 , \21819 , \21820 , \21821 , \21822 ,
         \21823 , \21824 , \21825 , \21826 , \21827 , \21828 , \21829 , \21830 , \21831 , \21832 ,
         \21833 , \21834 , \21835 , \21836 , \21837 , \21838 , \21839 , \21840 , \21841 , \21842 ,
         \21843 , \21844 , \21845 , \21846 , \21847 , \21848 , \21849 , \21850 , \21851 , \21852 ,
         \21853 , \21854 , \21855 , \21856 , \21857 , \21858 , \21859 , \21860 , \21861 , \21862 ,
         \21863 , \21864 , \21865 , \21866 , \21867 , \21868 , \21869 , \21870 , \21871 , \21872 ,
         \21873 , \21874 , \21875 , \21876 , \21877 , \21878 , \21879 , \21880 , \21881 , \21882 ,
         \21883 , \21884 , \21885 , \21886 , \21887 , \21888 , \21889 , \21890 , \21891 , \21892 ,
         \21893 , \21894 , \21895 , \21896 , \21897 , \21898 , \21899 , \21900 , \21901 , \21902 ,
         \21903 , \21904 , \21905 , \21906 , \21907 , \21908 , \21909 , \21910 , \21911 , \21912 ,
         \21913 , \21914 , \21915 , \21916 , \21917 , \21918 , \21919 , \21920 , \21921 , \21922 ,
         \21923 , \21924 , \21925 , \21926 , \21927 , \21928 , \21929 , \21930 , \21931 , \21932 ,
         \21933 , \21934 , \21935 , \21936 , \21937 , \21938 , \21939 , \21940 , \21941 , \21942 ,
         \21943 , \21944 , \21945 , \21946 , \21947 , \21948 , \21949 , \21950 , \21951 , \21952 ,
         \21953 , \21954 , \21955 , \21956 , \21957 , \21958 , \21959 , \21960 , \21961 , \21962 ,
         \21963 , \21964 , \21965 , \21966 , \21967 , \21968 , \21969 , \21970 , \21971 , \21972 ,
         \21973 , \21974 , \21975 , \21976 , \21977 , \21978 , \21979 , \21980 , \21981 , \21982 ,
         \21983 , \21984 , \21985 , \21986 , \21987 , \21988 , \21989 , \21990 , \21991 , \21992 ,
         \21993 , \21994 , \21995 , \21996 , \21997 , \21998 , \21999 , \22000 , \22001 , \22002 ,
         \22003 , \22004 , \22005 , \22006 , \22007 , \22008 , \22009 , \22010 , \22011 , \22012 ,
         \22013 , \22014 , \22015 , \22016 , \22017 , \22018 , \22019 , \22020 , \22021 , \22022 ,
         \22023 , \22024 , \22025 , \22026 , \22027 , \22028 , \22029 , \22030 , \22031 , \22032 ,
         \22033 , \22034 , \22035 , \22036 , \22037 , \22038 , \22039 , \22040 , \22041 , \22042 ,
         \22043 , \22044 , \22045 , \22046 , \22047 , \22048 , \22049 , \22050 , \22051 , \22052 ,
         \22053 , \22054 , \22055 , \22056 , \22057 , \22058 , \22059 , \22060 , \22061 , \22062 ,
         \22063 , \22064 , \22065 , \22066 , \22067 , \22068 , \22069 , \22070 , \22071 , \22072 ,
         \22073 , \22074 , \22075 , \22076 , \22077 , \22078 , \22079 , \22080 , \22081 , \22082 ,
         \22083 , \22084 , \22085 , \22086 , \22087 , \22088 , \22089 , \22090 , \22091 , \22092 ,
         \22093 , \22094 , \22095 , \22096 , \22097 , \22098 , \22099 , \22100 , \22101 , \22102 ,
         \22103 , \22104 , \22105 , \22106 , \22107 , \22108 , \22109 , \22110 , \22111 , \22112 ,
         \22113 , \22114 , \22115 , \22116 , \22117 , \22118 , \22119 , \22120 , \22121 , \22122 ,
         \22123 , \22124 , \22125 , \22126 , \22127 , \22128 , \22129 , \22130 , \22131 , \22132 ,
         \22133 , \22134 , \22135 , \22136 , \22137 , \22138 , \22139 , \22140 , \22141 , \22142 ,
         \22143 , \22144 , \22145 , \22146 , \22147 , \22148 , \22149 , \22150 , \22151 , \22152 ,
         \22153 , \22154 , \22155 , \22156 , \22157 , \22158 , \22159 , \22160 , \22161 , \22162 ,
         \22163 , \22164 , \22165 , \22166 , \22167 , \22168 , \22169 , \22170 , \22171 , \22172 ,
         \22173 , \22174 , \22175 , \22176 , \22177 , \22178 , \22179 , \22180 , \22181 , \22182 ,
         \22183 , \22184 , \22185 , \22186 , \22187 , \22188 , \22189 , \22190 , \22191 , \22192 ,
         \22193 , \22194 , \22195 , \22196 , \22197 , \22198 , \22199 , \22200 , \22201 , \22202 ,
         \22203 , \22204 , \22205 , \22206 , \22207 , \22208 , \22209 , \22210 , \22211 , \22212 ,
         \22213 , \22214 , \22215 , \22216 , \22217 , \22218 , \22219 , \22220 , \22221 , \22222 ,
         \22223 , \22224 , \22225 , \22226 , \22227 , \22228 , \22229 , \22230 , \22231 , \22232 ,
         \22233 , \22234 , \22235 , \22236 , \22237 , \22238 , \22239 , \22240 , \22241 , \22242 ,
         \22243 , \22244 , \22245 , \22246 , \22247 , \22248 , \22249 , \22250 , \22251 , \22252 ,
         \22253 , \22254 , \22255 , \22256 , \22257 , \22258 , \22259 , \22260 , \22261 , \22262 ,
         \22263 , \22264 , \22265 , \22266 , \22267 , \22268 , \22269 , \22270 , \22271 , \22272 ,
         \22273 , \22274 , \22275 , \22276 , \22277 , \22278 , \22279 , \22280 , \22281 , \22282 ,
         \22283 , \22284 , \22285 , \22286 , \22287 , \22288 , \22289 , \22290 , \22291 , \22292 ,
         \22293 , \22294 , \22295 , \22296 , \22297 , \22298 , \22299 , \22300 , \22301 , \22302 ,
         \22303 , \22304 , \22305 , \22306 , \22307 , \22308 , \22309 , \22310 , \22311 , \22312 ,
         \22313 , \22314 , \22315 , \22316 , \22317 , \22318 , \22319 , \22320 , \22321 , \22322 ,
         \22323 , \22324 , \22325 , \22326 , \22327 , \22328 , \22329 , \22330 , \22331 , \22332 ,
         \22333 , \22334 , \22335 , \22336 , \22337 , \22338 , \22339 , \22340 , \22341 , \22342 ,
         \22343 , \22344 , \22345 , \22346 , \22347 , \22348 , \22349 , \22350 , \22351 , \22352 ,
         \22353 , \22354 , \22355 , \22356 , \22357 , \22358 , \22359 , \22360 , \22361 , \22362 ,
         \22363 , \22364 , \22365 , \22366 , \22367 , \22368 , \22369 , \22370 , \22371 , \22372 ,
         \22373 , \22374 , \22375 , \22376 , \22377 , \22378 , \22379 , \22380 , \22381 , \22382 ,
         \22383 , \22384 , \22385 , \22386 , \22387 , \22388 , \22389 , \22390 , \22391 , \22392 ,
         \22393 , \22394 , \22395 , \22396 , \22397 , \22398 , \22399 , \22400 , \22401 , \22402 ,
         \22403 , \22404 , \22405 , \22406 , \22407 , \22408 , \22409 , \22410 , \22411 , \22412 ,
         \22413 , \22414 , \22415 , \22416 , \22417 , \22418 , \22419 , \22420 , \22421 , \22422 ,
         \22423 , \22424 , \22425 , \22426 , \22427 , \22428 , \22429 , \22430 , \22431 , \22432 ,
         \22433 , \22434 , \22435 , \22436 , \22437 , \22438 , \22439 , \22440 , \22441 , \22442 ,
         \22443 , \22444 , \22445 , \22446 , \22447 , \22448 , \22449 , \22450 , \22451 , \22452 ,
         \22453 , \22454 , \22455 , \22456 , \22457 , \22458 , \22459 , \22460 , \22461 , \22462 ,
         \22463 , \22464 , \22465 , \22466 , \22467 , \22468 , \22469 , \22470 , \22471 , \22472 ,
         \22473 , \22474 , \22475 , \22476 , \22477 , \22478 , \22479 , \22480 , \22481 , \22482 ,
         \22483 , \22484 , \22485 , \22486 , \22487 , \22488 , \22489 , \22490 , \22491 , \22492 ,
         \22493 , \22494 , \22495 , \22496 , \22497 , \22498 , \22499 , \22500 , \22501 , \22502 ,
         \22503 , \22504 , \22505 , \22506 , \22507 , \22508 , \22509 , \22510 , \22511 , \22512 ,
         \22513 , \22514 , \22515 , \22516 , \22517 , \22518 , \22519 , \22520 , \22521 , \22522 ,
         \22523 , \22524 , \22525 , \22526 , \22527 , \22528 , \22529 , \22530 , \22531 , \22532 ,
         \22533 , \22534 , \22535 , \22536 , \22537 , \22538 , \22539 , \22540 , \22541 , \22542 ,
         \22543 , \22544 , \22545 , \22546 , \22547 , \22548 , \22549 , \22550 , \22551 , \22552 ,
         \22553 , \22554 , \22555 , \22556 , \22557 , \22558 , \22559 , \22560 , \22561 , \22562 ,
         \22563 , \22564 , \22565 , \22566 , \22567 , \22568 , \22569 , \22570 , \22571 , \22572 ,
         \22573 , \22574 , \22575 , \22576 , \22577 , \22578 , \22579 , \22580 , \22581 , \22582 ,
         \22583 , \22584 , \22585 , \22586 , \22587 , \22588 , \22589 , \22590 , \22591 , \22592 ,
         \22593 , \22594 , \22595 , \22596 , \22597 , \22598 , \22599 , \22600 , \22601 , \22602 ,
         \22603 , \22604 , \22605 , \22606 , \22607 , \22608 , \22609 , \22610 , \22611 , \22612 ,
         \22613 , \22614 , \22615 , \22616 , \22617 , \22618 , \22619 , \22620 , \22621 , \22622 ,
         \22623 , \22624 , \22625 , \22626 , \22627 , \22628 , \22629 , \22630 , \22631 , \22632 ,
         \22633 , \22634 , \22635 , \22636 , \22637 , \22638 , \22639 , \22640 , \22641 , \22642 ,
         \22643 , \22644 , \22645 , \22646 , \22647 , \22648 , \22649 , \22650 , \22651 , \22652 ,
         \22653 , \22654 , \22655 , \22656 , \22657 , \22658 , \22659 , \22660 , \22661 , \22662 ,
         \22663 , \22664 , \22665 , \22666 , \22667 , \22668 , \22669 , \22670 , \22671 , \22672 ,
         \22673 , \22674 , \22675 , \22676 , \22677 , \22678 , \22679 , \22680 , \22681 , \22682 ,
         \22683 , \22684 , \22685 , \22686 , \22687 , \22688 , \22689 , \22690 , \22691 , \22692 ,
         \22693 , \22694 , \22695 , \22696 , \22697 , \22698 , \22699 , \22700 , \22701 , \22702 ,
         \22703 , \22704 , \22705 , \22706 , \22707 , \22708 , \22709 , \22710 , \22711 , \22712 ,
         \22713 , \22714 , \22715 , \22716 , \22717 , \22718 , \22719 , \22720 , \22721 , \22722 ,
         \22723 , \22724 , \22725 , \22726 , \22727 , \22728 , \22729 , \22730 , \22731 , \22732 ,
         \22733 , \22734 , \22735 , \22736 , \22737 , \22738 , \22739 , \22740 , \22741 , \22742 ,
         \22743 , \22744 , \22745 , \22746 , \22747 , \22748 , \22749 , \22750 , \22751 , \22752 ,
         \22753 , \22754 , \22755 , \22756 , \22757 , \22758 , \22759 , \22760 , \22761 , \22762 ,
         \22763 , \22764 , \22765 , \22766 , \22767 , \22768 , \22769 , \22770 , \22771 , \22772 ,
         \22773 , \22774 , \22775 , \22776 , \22777 , \22778 , \22779 , \22780 , \22781 , \22782 ,
         \22783 , \22784 , \22785 , \22786 , \22787 , \22788 , \22789 , \22790 , \22791 , \22792 ,
         \22793 , \22794 , \22795 , \22796 , \22797 , \22798 , \22799 , \22800 , \22801 , \22802 ,
         \22803 , \22804 , \22805 , \22806 , \22807 , \22808 , \22809 , \22810 , \22811 , \22812 ,
         \22813 , \22814 , \22815 , \22816 , \22817 , \22818 , \22819 , \22820 , \22821 , \22822 ,
         \22823 , \22824 , \22825 , \22826 , \22827 , \22828 , \22829 , \22830 , \22831 , \22832 ,
         \22833 , \22834 , \22835 , \22836 , \22837 , \22838 , \22839 , \22840 , \22841 , \22842 ,
         \22843 , \22844 , \22845 , \22846 , \22847 , \22848 , \22849 , \22850 , \22851 , \22852 ,
         \22853 , \22854 , \22855 , \22856 , \22857 , \22858 , \22859 , \22860 , \22861 , \22862 ,
         \22863 , \22864 , \22865 , \22866 , \22867 , \22868 , \22869 , \22870 , \22871 , \22872 ,
         \22873 , \22874 , \22875 , \22876 , \22877 , \22878 , \22879 , \22880 , \22881 , \22882 ,
         \22883 , \22884 , \22885 , \22886 , \22887 , \22888 , \22889 , \22890 , \22891 , \22892 ,
         \22893 , \22894 , \22895 , \22896 , \22897 , \22898 , \22899 , \22900 , \22901 , \22902 ,
         \22903 , \22904 , \22905 , \22906 , \22907 , \22908 , \22909 , \22910 , \22911 , \22912 ,
         \22913 , \22914 , \22915 , \22916 , \22917 , \22918 , \22919 , \22920 , \22921 , \22922 ,
         \22923 , \22924 , \22925 , \22926 , \22927 , \22928 , \22929 , \22930 , \22931 , \22932 ,
         \22933 , \22934 , \22935 , \22936 , \22937 , \22938 , \22939 , \22940 , \22941 , \22942 ,
         \22943 , \22944 , \22945 , \22946 , \22947 , \22948 , \22949 , \22950 , \22951 , \22952 ,
         \22953 , \22954 , \22955 , \22956 , \22957 , \22958 , \22959 , \22960 , \22961 , \22962 ,
         \22963 , \22964 , \22965 , \22966 , \22967 , \22968 , \22969 , \22970 , \22971 , \22972 ,
         \22973 , \22974 , \22975 , \22976 , \22977 , \22978 , \22979 , \22980 , \22981 , \22982 ,
         \22983 , \22984 , \22985 , \22986 , \22987 , \22988 , \22989 , \22990 , \22991 , \22992 ,
         \22993 , \22994 , \22995 , \22996 , \22997 , \22998 , \22999 , \23000 , \23001 , \23002 ,
         \23003 , \23004 , \23005 , \23006 , \23007 , \23008 , \23009 , \23010 , \23011 , \23012 ,
         \23013 , \23014 , \23015 , \23016 , \23017 , \23018 , \23019 , \23020 , \23021 , \23022 ,
         \23023 , \23024 , \23025 , \23026 , \23027 , \23028 , \23029 , \23030 , \23031 , \23032 ,
         \23033 , \23034 , \23035 , \23036 , \23037 , \23038 , \23039 , \23040 , \23041 , \23042 ,
         \23043 , \23044 , \23045 , \23046 , \23047 , \23048 , \23049 , \23050 , \23051 , \23052 ,
         \23053 , \23054 , \23055 , \23056 , \23057 , \23058 , \23059 , \23060 , \23061 , \23062 ,
         \23063 , \23064 , \23065 , \23066 , \23067 , \23068 , \23069 , \23070 , \23071 , \23072 ,
         \23073 , \23074 , \23075 , \23076 , \23077 , \23078 , \23079 , \23080 , \23081 , \23082 ,
         \23083 , \23084 , \23085 , \23086 , \23087 , \23088 , \23089 , \23090 , \23091 , \23092 ,
         \23093 , \23094 , \23095 , \23096 , \23097 , \23098 , \23099 , \23100 , \23101 , \23102 ,
         \23103 , \23104 , \23105 , \23106 , \23107 , \23108 , \23109 , \23110 , \23111 , \23112 ,
         \23113 , \23114 , \23115 , \23116 , \23117 , \23118 , \23119 , \23120 , \23121 , \23122 ,
         \23123 , \23124 , \23125 , \23126 , \23127 , \23128 , \23129 , \23130 , \23131 , \23132 ,
         \23133 , \23134 , \23135 , \23136 , \23137 , \23138 , \23139 , \23140 , \23141 , \23142 ,
         \23143 , \23144 , \23145 , \23146 , \23147 , \23148 , \23149 , \23150 , \23151 , \23152 ,
         \23153 , \23154 , \23155 , \23156 , \23157 , \23158 , \23159 , \23160 , \23161 , \23162 ,
         \23163 , \23164 , \23165 , \23166 , \23167 , \23168 , \23169 , \23170 , \23171 , \23172 ,
         \23173 , \23174 , \23175 , \23176 , \23177 , \23178 , \23179 , \23180 , \23181 , \23182 ,
         \23183 , \23184 , \23185 , \23186 , \23187 , \23188 , \23189 , \23190 , \23191 , \23192 ,
         \23193 , \23194 , \23195 , \23196 , \23197 , \23198 , \23199 , \23200 , \23201 , \23202 ,
         \23203 , \23204 , \23205 , \23206 , \23207 , \23208 , \23209 , \23210 , \23211 , \23212 ,
         \23213 , \23214 , \23215 , \23216 , \23217 , \23218 , \23219 , \23220 , \23221 , \23222 ,
         \23223 , \23224 , \23225 , \23226 , \23227 , \23228 , \23229 , \23230 , \23231 , \23232 ,
         \23233 , \23234 , \23235 , \23236 , \23237 , \23238 , \23239 , \23240 , \23241 , \23242 ,
         \23243 , \23244 , \23245 , \23246 , \23247 , \23248 , \23249 , \23250 , \23251 , \23252 ,
         \23253 , \23254 , \23255 , \23256 , \23257 , \23258 , \23259 , \23260 , \23261 , \23262 ,
         \23263 , \23264 , \23265 , \23266 , \23267 , \23268 , \23269 , \23270 , \23271 , \23272 ,
         \23273 , \23274 , \23275 , \23276 , \23277 , \23278 , \23279 , \23280 , \23281 , \23282 ,
         \23283 , \23284 , \23285 , \23286 , \23287 , \23288 , \23289 , \23290 , \23291 , \23292 ,
         \23293 , \23294 , \23295 , \23296 , \23297 , \23298 , \23299 , \23300 , \23301 , \23302 ,
         \23303 , \23304 , \23305 , \23306 , \23307 , \23308 , \23309 , \23310 , \23311 , \23312 ,
         \23313 , \23314 , \23315 , \23316 , \23317 , \23318 , \23319 , \23320 , \23321 , \23322 ,
         \23323 , \23324 , \23325 , \23326 , \23327 , \23328 , \23329 , \23330 , \23331 , \23332 ,
         \23333 , \23334 , \23335 , \23336 , \23337 , \23338 , \23339 , \23340 , \23341 , \23342 ,
         \23343 , \23344 , \23345 , \23346 , \23347 , \23348 , \23349 , \23350 , \23351 , \23352 ,
         \23353 , \23354 , \23355 , \23356 , \23357 , \23358 , \23359 , \23360 , \23361 , \23362 ,
         \23363 , \23364 , \23365 , \23366 , \23367 , \23368 , \23369 , \23370 , \23371 , \23372 ,
         \23373 , \23374 , \23375 , \23376 , \23377 , \23378 , \23379 , \23380 , \23381 , \23382 ,
         \23383 , \23384 , \23385 , \23386 , \23387 , \23388 , \23389 , \23390 , \23391 , \23392 ,
         \23393 , \23394 , \23395 , \23396 , \23397 , \23398 , \23399 , \23400 , \23401 , \23402 ,
         \23403 , \23404 , \23405 , \23406 , \23407 , \23408 , \23409 , \23410 , \23411 , \23412 ,
         \23413 , \23414 , \23415 , \23416 , \23417 , \23418 , \23419 , \23420 , \23421 , \23422 ,
         \23423 , \23424 , \23425 , \23426 , \23427 , \23428 , \23429 , \23430 , \23431 , \23432 ,
         \23433 , \23434 , \23435 , \23436 , \23437 , \23438 , \23439 , \23440 , \23441 , \23442 ,
         \23443 , \23444 , \23445 , \23446 , \23447 , \23448 , \23449 , \23450 , \23451 , \23452 ,
         \23453 , \23454 , \23455 , \23456 , \23457 , \23458 , \23459 , \23460 , \23461 , \23462 ,
         \23463 , \23464 , \23465 , \23466 , \23467 , \23468 , \23469 , \23470 , \23471 , \23472 ,
         \23473 , \23474 , \23475 , \23476 , \23477 , \23478 , \23479 , \23480 , \23481 , \23482 ,
         \23483 , \23484 , \23485 , \23486 , \23487 , \23488 , \23489 , \23490 , \23491 , \23492 ,
         \23493 , \23494 , \23495 , \23496 , \23497 , \23498 , \23499 , \23500 , \23501 , \23502 ,
         \23503 , \23504 , \23505 , \23506 , \23507 , \23508 , \23509 , \23510 , \23511 , \23512 ,
         \23513 , \23514 , \23515 , \23516 , \23517 , \23518 , \23519 , \23520 , \23521 , \23522 ,
         \23523 , \23524 , \23525 , \23526 , \23527 , \23528 , \23529 , \23530 , \23531 , \23532 ,
         \23533 , \23534 , \23535 , \23536 , \23537 , \23538 , \23539 , \23540 , \23541 , \23542 ,
         \23543 , \23544 , \23545 , \23546 , \23547 , \23548 , \23549 , \23550 , \23551 , \23552 ,
         \23553 , \23554 , \23555 , \23556 , \23557 , \23558 , \23559 , \23560 , \23561 , \23562 ,
         \23563 , \23564 , \23565 , \23566 , \23567 , \23568 , \23569 , \23570 , \23571 , \23572 ,
         \23573 , \23574 , \23575 , \23576 , \23577 , \23578 , \23579 , \23580 , \23581 , \23582 ,
         \23583 , \23584 , \23585 , \23586 , \23587 , \23588 , \23589 , \23590 , \23591 , \23592 ,
         \23593 , \23594 , \23595 , \23596 , \23597 , \23598 , \23599 , \23600 , \23601 , \23602 ,
         \23603 , \23604 , \23605 , \23606 , \23607 , \23608 , \23609 , \23610 , \23611 , \23612 ,
         \23613 , \23614 , \23615 , \23616 , \23617 , \23618 , \23619 , \23620 , \23621 , \23622 ,
         \23623 , \23624 , \23625 , \23626 , \23627 , \23628 , \23629 , \23630 , \23631 , \23632 ,
         \23633 , \23634 , \23635 , \23636 , \23637 , \23638 , \23639 , \23640 , \23641 , \23642 ,
         \23643 , \23644 , \23645 , \23646 , \23647 , \23648 , \23649 , \23650 , \23651 , \23652 ,
         \23653 , \23654 , \23655 , \23656 , \23657 , \23658 , \23659 , \23660 , \23661 , \23662 ,
         \23663 , \23664 , \23665 , \23666 , \23667 , \23668 , \23669 , \23670 , \23671 , \23672 ,
         \23673 , \23674 , \23675 , \23676 , \23677 , \23678 , \23679 , \23680 , \23681 , \23682 ,
         \23683 , \23684 , \23685 , \23686 , \23687 , \23688 , \23689 , \23690 , \23691 , \23692 ,
         \23693 , \23694 , \23695 , \23696 , \23697 , \23698 , \23699 , \23700 , \23701 , \23702 ,
         \23703 , \23704 , \23705 , \23706 , \23707 , \23708 , \23709 , \23710 , \23711 , \23712 ,
         \23713 , \23714 , \23715 , \23716 , \23717 , \23718 , \23719 , \23720 , \23721 , \23722 ,
         \23723 , \23724 , \23725 , \23726 , \23727 , \23728 , \23729 , \23730 , \23731 , \23732 ,
         \23733 , \23734 , \23735 , \23736 , \23737 , \23738 , \23739 , \23740 , \23741 , \23742 ,
         \23743 , \23744 , \23745 , \23746 , \23747 , \23748 , \23749 , \23750 , \23751 , \23752 ,
         \23753 , \23754 , \23755 , \23756 , \23757 , \23758 , \23759 , \23760 , \23761 , \23762 ,
         \23763 , \23764 , \23765 , \23766 , \23767 , \23768 , \23769 , \23770 , \23771 , \23772 ,
         \23773 , \23774 , \23775 , \23776 , \23777 , \23778 , \23779 , \23780 , \23781 , \23782 ,
         \23783 , \23784 , \23785 , \23786 , \23787 , \23788 , \23789 , \23790 , \23791 , \23792 ,
         \23793 , \23794 , \23795 , \23796 , \23797 , \23798 , \23799 , \23800 , \23801 , \23802 ,
         \23803 , \23804 , \23805 , \23806 , \23807 , \23808 , \23809 , \23810 , \23811 , \23812 ,
         \23813 , \23814 , \23815 , \23816 , \23817 , \23818 , \23819 , \23820 , \23821 , \23822 ,
         \23823 , \23824 , \23825 , \23826 , \23827 , \23828 , \23829 , \23830 , \23831 , \23832 ,
         \23833 , \23834 , \23835 , \23836 , \23837 , \23838 , \23839 , \23840 , \23841 , \23842 ,
         \23843 , \23844 , \23845 , \23846 , \23847 , \23848 , \23849 , \23850 , \23851 , \23852 ,
         \23853 , \23854 , \23855 , \23856 , \23857 , \23858 , \23859 , \23860 , \23861 , \23862 ,
         \23863 , \23864 , \23865 , \23866 , \23867 , \23868 , \23869 , \23870 , \23871 , \23872 ,
         \23873 , \23874 , \23875 , \23876 , \23877 , \23878 , \23879 , \23880 , \23881 , \23882 ,
         \23883 , \23884 , \23885 , \23886 , \23887 , \23888 , \23889 , \23890 , \23891 , \23892 ,
         \23893 , \23894 , \23895 , \23896 , \23897 , \23898 , \23899 , \23900 , \23901 , \23902 ,
         \23903 , \23904 , \23905 , \23906 , \23907 , \23908 , \23909 , \23910 , \23911 , \23912 ,
         \23913 , \23914 , \23915 , \23916 , \23917 , \23918 , \23919 , \23920 , \23921 , \23922 ,
         \23923 , \23924 , \23925 , \23926 , \23927 , \23928 , \23929 , \23930 , \23931 , \23932 ,
         \23933 , \23934 , \23935 , \23936 , \23937 , \23938 , \23939 , \23940 , \23941 , \23942 ,
         \23943 , \23944 , \23945 , \23946 , \23947 , \23948 , \23949 , \23950 , \23951 , \23952 ,
         \23953 , \23954 , \23955 , \23956 , \23957 , \23958 , \23959 , \23960 , \23961 , \23962 ,
         \23963 , \23964 , \23965 , \23966 , \23967 , \23968 , \23969 , \23970 , \23971 , \23972 ,
         \23973 , \23974 , \23975 , \23976 , \23977 , \23978 , \23979 , \23980 , \23981 , \23982 ,
         \23983 , \23984 , \23985 , \23986 , \23987 , \23988 , \23989 , \23990 , \23991 , \23992 ,
         \23993 , \23994 , \23995 , \23996 , \23997 , \23998 , \23999 , \24000 , \24001 , \24002 ,
         \24003 , \24004 , \24005 , \24006 , \24007 , \24008 , \24009 , \24010 , \24011 , \24012 ,
         \24013 , \24014 , \24015 , \24016 , \24017 , \24018 , \24019 , \24020 , \24021 , \24022 ,
         \24023 , \24024 , \24025 , \24026 , \24027 , \24028 , \24029 , \24030 , \24031 , \24032 ,
         \24033 , \24034 , \24035 , \24036 , \24037 , \24038 , \24039 , \24040 , \24041 , \24042 ,
         \24043 , \24044 , \24045 , \24046 , \24047 , \24048 , \24049 , \24050 , \24051 , \24052 ,
         \24053 , \24054 , \24055 , \24056 , \24057 , \24058 , \24059 , \24060 , \24061 , \24062 ,
         \24063 , \24064 , \24065 , \24066 , \24067 , \24068 , \24069 , \24070 , \24071 , \24072 ,
         \24073 , \24074 , \24075 , \24076 , \24077 , \24078 , \24079 , \24080 , \24081 , \24082 ,
         \24083 , \24084 , \24085 , \24086 , \24087 , \24088 , \24089 , \24090 , \24091 , \24092 ,
         \24093 , \24094 , \24095 , \24096 , \24097 , \24098 , \24099 , \24100 , \24101 , \24102 ,
         \24103 , \24104 , \24105 , \24106 , \24107 , \24108 , \24109 , \24110 , \24111 , \24112 ,
         \24113 , \24114 , \24115 , \24116 , \24117 , \24118 , \24119 , \24120 , \24121 , \24122 ,
         \24123 , \24124 , \24125 , \24126 , \24127 , \24128 , \24129 , \24130 , \24131 , \24132 ,
         \24133 , \24134 , \24135 , \24136 , \24137 , \24138 , \24139 , \24140 , \24141 , \24142 ,
         \24143 , \24144 , \24145 , \24146 , \24147 , \24148 , \24149 , \24150 , \24151 , \24152 ,
         \24153 , \24154 , \24155 , \24156 , \24157 , \24158 , \24159 , \24160 , \24161 , \24162 ,
         \24163 , \24164 , \24165 , \24166 , \24167 , \24168 , \24169 , \24170 , \24171 , \24172 ,
         \24173 , \24174 , \24175 , \24176 , \24177 , \24178 , \24179 , \24180 , \24181 , \24182 ,
         \24183 , \24184 , \24185 , \24186 , \24187 , \24188 , \24189 , \24190 , \24191 , \24192 ,
         \24193 , \24194 , \24195 , \24196 , \24197 , \24198 , \24199 , \24200 , \24201 , \24202 ,
         \24203 , \24204 , \24205 , \24206 , \24207 , \24208 , \24209 , \24210 , \24211 , \24212 ,
         \24213 , \24214 , \24215 , \24216 , \24217 , \24218 , \24219 , \24220 , \24221 , \24222 ,
         \24223 , \24224 , \24225 , \24226 , \24227 , \24228 , \24229 , \24230 , \24231 , \24232 ,
         \24233 , \24234 , \24235 , \24236 , \24237 , \24238 , \24239 , \24240 , \24241 , \24242 ,
         \24243 , \24244 , \24245 , \24246 , \24247 , \24248 , \24249 , \24250 , \24251 , \24252 ,
         \24253 , \24254 , \24255 , \24256 , \24257 , \24258 , \24259 , \24260 , \24261 , \24262 ,
         \24263 , \24264 , \24265 , \24266 , \24267 , \24268 , \24269 , \24270 , \24271 , \24272 ,
         \24273 , \24274 , \24275 , \24276 , \24277 , \24278 , \24279 , \24280 , \24281 , \24282 ,
         \24283 , \24284 , \24285 , \24286 , \24287 , \24288 , \24289 , \24290 , \24291 , \24292 ,
         \24293 , \24294 , \24295 , \24296 , \24297 , \24298 , \24299 , \24300 , \24301 , \24302 ,
         \24303 , \24304 , \24305 , \24306 , \24307 , \24308 , \24309 , \24310 , \24311 , \24312 ,
         \24313 , \24314 , \24315 , \24316 , \24317 , \24318 , \24319 , \24320 , \24321 , \24322 ,
         \24323 , \24324 , \24325 , \24326 , \24327 , \24328 , \24329 , \24330 , \24331 , \24332 ,
         \24333 , \24334 , \24335 , \24336 , \24337 , \24338 , \24339 , \24340 , \24341 , \24342 ,
         \24343 , \24344 , \24345 , \24346 , \24347 , \24348 , \24349 , \24350 , \24351 , \24352 ,
         \24353 , \24354 , \24355 , \24356 , \24357 , \24358 , \24359 , \24360 , \24361 , \24362 ,
         \24363 , \24364 , \24365 , \24366 , \24367 , \24368 , \24369 , \24370 , \24371 , \24372 ,
         \24373 , \24374 , \24375 , \24376 , \24377 , \24378 , \24379 , \24380 , \24381 , \24382 ,
         \24383 , \24384 , \24385 , \24386 , \24387 , \24388 , \24389 , \24390 , \24391 , \24392 ,
         \24393 , \24394 , \24395 , \24396 , \24397 , \24398 , \24399 , \24400 , \24401 , \24402 ,
         \24403 , \24404 , \24405 , \24406 , \24407 , \24408 , \24409 , \24410 , \24411 , \24412 ,
         \24413 , \24414 , \24415 , \24416 , \24417 , \24418 , \24419 , \24420 , \24421 , \24422 ,
         \24423 , \24424 , \24425 , \24426 , \24427 , \24428 , \24429 , \24430 , \24431 , \24432 ,
         \24433 , \24434 , \24435 , \24436 , \24437 , \24438 , \24439 , \24440 , \24441 , \24442 ,
         \24443 , \24444 , \24445 , \24446 , \24447 , \24448 , \24449 , \24450 , \24451 , \24452 ,
         \24453 , \24454 , \24455 , \24456 , \24457 , \24458 , \24459 , \24460 , \24461 , \24462 ,
         \24463 , \24464 , \24465 , \24466 , \24467 , \24468 , \24469 , \24470 , \24471 , \24472 ,
         \24473 , \24474 , \24475 , \24476 , \24477 , \24478 , \24479 , \24480 , \24481 , \24482 ,
         \24483 , \24484 , \24485 , \24486 , \24487 , \24488 , \24489 , \24490 , \24491 , \24492 ,
         \24493 , \24494 , \24495 , \24496 , \24497 , \24498 , \24499 , \24500 , \24501 , \24502 ,
         \24503 , \24504 , \24505 , \24506 , \24507 , \24508 , \24509 , \24510 , \24511 , \24512 ,
         \24513 , \24514 , \24515 , \24516 , \24517 , \24518 , \24519 , \24520 , \24521 , \24522 ,
         \24523 , \24524 , \24525 , \24526 , \24527 , \24528 , \24529 , \24530 , \24531 , \24532 ,
         \24533 , \24534 , \24535 , \24536 , \24537 , \24538 , \24539 , \24540 , \24541 , \24542 ,
         \24543 , \24544 , \24545 , \24546 , \24547 , \24548 , \24549 , \24550 , \24551 , \24552 ,
         \24553 , \24554 , \24555 , \24556 , \24557 , \24558 , \24559 , \24560 , \24561 , \24562 ,
         \24563 , \24564 , \24565 , \24566 , \24567 , \24568 , \24569 , \24570 , \24571 , \24572 ,
         \24573 , \24574 , \24575 , \24576 , \24577 , \24578 , \24579 , \24580 , \24581 , \24582 ,
         \24583 , \24584 , \24585 , \24586 , \24587 , \24588 , \24589 , \24590 , \24591 , \24592 ,
         \24593 , \24594 , \24595 , \24596 , \24597 , \24598 , \24599 , \24600 , \24601 , \24602 ,
         \24603 , \24604 , \24605 , \24606 , \24607 , \24608 , \24609 , \24610 , \24611 , \24612 ,
         \24613 , \24614 , \24615 , \24616 , \24617 , \24618 , \24619 , \24620 , \24621 , \24622 ,
         \24623 , \24624 , \24625 , \24626 , \24627 , \24628 , \24629 , \24630 , \24631 , \24632 ,
         \24633 , \24634 , \24635 , \24636 , \24637 , \24638 , \24639 , \24640 , \24641 , \24642 ,
         \24643 , \24644 , \24645 , \24646 , \24647 , \24648 , \24649 , \24650 , \24651 , \24652 ,
         \24653 , \24654 , \24655 , \24656 , \24657 , \24658 , \24659 , \24660 , \24661 , \24662 ,
         \24663 , \24664 , \24665 , \24666 , \24667 , \24668 , \24669 , \24670 , \24671 , \24672 ,
         \24673 , \24674 , \24675 , \24676 , \24677 , \24678 , \24679 , \24680 , \24681 , \24682 ,
         \24683 , \24684 , \24685 , \24686 , \24687 , \24688 , \24689 , \24690 , \24691 , \24692 ,
         \24693 , \24694 , \24695 , \24696 , \24697 , \24698 , \24699 , \24700 , \24701 , \24702 ,
         \24703 , \24704 , \24705 , \24706 , \24707 , \24708 , \24709 , \24710 , \24711 , \24712 ,
         \24713 , \24714 , \24715 , \24716 , \24717 , \24718 , \24719 , \24720 , \24721 , \24722 ,
         \24723 , \24724 , \24725 , \24726 , \24727 , \24728 , \24729 , \24730 , \24731 , \24732 ,
         \24733 , \24734 , \24735 , \24736 , \24737 , \24738 , \24739 , \24740 , \24741 , \24742 ,
         \24743 , \24744 , \24745 , \24746 , \24747 , \24748 , \24749 , \24750 , \24751 , \24752 ,
         \24753 , \24754 , \24755 , \24756 , \24757 , \24758 , \24759 , \24760 , \24761 , \24762 ,
         \24763 , \24764 , \24765 , \24766 , \24767 , \24768 , \24769 , \24770 , \24771 , \24772 ,
         \24773 , \24774 , \24775 , \24776 , \24777 , \24778 , \24779 , \24780 , \24781 , \24782 ,
         \24783 , \24784 , \24785 , \24786 , \24787 , \24788 , \24789 , \24790 , \24791 , \24792 ,
         \24793 , \24794 , \24795 , \24796 , \24797 , \24798 , \24799 , \24800 , \24801 , \24802 ,
         \24803 , \24804 , \24805 , \24806 , \24807 , \24808 , \24809 , \24810 , \24811 , \24812 ,
         \24813 , \24814 , \24815 , \24816 , \24817 , \24818 , \24819 , \24820 , \24821 , \24822 ,
         \24823 , \24824 , \24825 , \24826 , \24827 , \24828 , \24829 , \24830 , \24831 , \24832 ,
         \24833 , \24834 , \24835 , \24836 , \24837 , \24838 , \24839 , \24840 , \24841 , \24842 ,
         \24843 , \24844 , \24845 , \24846 , \24847 , \24848 , \24849 , \24850 , \24851 , \24852 ,
         \24853 , \24854 , \24855 , \24856 , \24857 , \24858 , \24859 , \24860 , \24861 , \24862 ,
         \24863 , \24864 , \24865 , \24866 , \24867 , \24868 , \24869 , \24870 , \24871 , \24872 ,
         \24873 , \24874 , \24875 , \24876 , \24877 , \24878 , \24879 , \24880 , \24881 , \24882 ,
         \24883 , \24884 , \24885 , \24886 , \24887 , \24888 , \24889 , \24890 , \24891 , \24892 ,
         \24893 , \24894 , \24895 , \24896 , \24897 , \24898 , \24899 , \24900 , \24901 , \24902 ,
         \24903 , \24904 , \24905 , \24906 , \24907 , \24908 , \24909 , \24910 , \24911 , \24912 ,
         \24913 , \24914 , \24915 , \24916 , \24917 , \24918 , \24919 , \24920 , \24921 , \24922 ,
         \24923 , \24924 , \24925 , \24926 , \24927 , \24928 , \24929 , \24930 , \24931 , \24932 ,
         \24933 , \24934 , \24935 , \24936 , \24937 , \24938 , \24939 , \24940 , \24941 , \24942 ,
         \24943 , \24944 , \24945 , \24946 , \24947 , \24948 , \24949 , \24950 , \24951 , \24952 ,
         \24953 , \24954 , \24955 , \24956 , \24957 , \24958 , \24959 , \24960 , \24961 , \24962 ,
         \24963 , \24964 , \24965 , \24966 , \24967 , \24968 , \24969 , \24970 , \24971 , \24972 ,
         \24973 , \24974 , \24975 , \24976 , \24977 , \24978 , \24979 , \24980 , \24981 , \24982 ,
         \24983 , \24984 , \24985 , \24986 , \24987 , \24988 , \24989 , \24990 , \24991 , \24992 ,
         \24993 , \24994 , \24995 , \24996 , \24997 , \24998 , \24999 , \25000 , \25001 , \25002 ,
         \25003 , \25004 , \25005 , \25006 , \25007 , \25008 , \25009 , \25010 , \25011 , \25012 ,
         \25013 , \25014 , \25015 , \25016 , \25017 , \25018 , \25019 , \25020 , \25021 , \25022 ,
         \25023 , \25024 , \25025 , \25026 , \25027 , \25028 , \25029 , \25030 , \25031 , \25032 ,
         \25033 , \25034 , \25035 , \25036 , \25037 , \25038 , \25039 , \25040 , \25041 , \25042 ,
         \25043 , \25044 , \25045 , \25046 , \25047 , \25048 , \25049 , \25050 , \25051 , \25052 ,
         \25053 , \25054 , \25055 , \25056 , \25057 , \25058 , \25059 , \25060 , \25061 , \25062 ,
         \25063 , \25064 , \25065 , \25066 , \25067 , \25068 , \25069 , \25070 , \25071 , \25072 ,
         \25073 , \25074 , \25075 , \25076 , \25077 , \25078 , \25079 , \25080 , \25081 , \25082 ,
         \25083 , \25084 , \25085 , \25086 , \25087 , \25088 , \25089 , \25090 , \25091 , \25092 ,
         \25093 , \25094 , \25095 , \25096 , \25097 , \25098 , \25099 , \25100 , \25101 , \25102 ,
         \25103 , \25104 , \25105 , \25106 , \25107 , \25108 , \25109 , \25110 , \25111 , \25112 ,
         \25113 , \25114 , \25115 , \25116 , \25117 , \25118 , \25119 , \25120 , \25121 , \25122 ,
         \25123 , \25124 , \25125 , \25126 , \25127 , \25128 , \25129 , \25130 , \25131 , \25132 ,
         \25133 , \25134 , \25135 , \25136 , \25137 , \25138 , \25139 , \25140 , \25141 , \25142 ,
         \25143 , \25144 , \25145 , \25146 , \25147 , \25148 , \25149 , \25150 , \25151 , \25152 ,
         \25153 , \25154 , \25155 , \25156 , \25157 , \25158 , \25159 , \25160 , \25161 , \25162 ,
         \25163 , \25164 , \25165 , \25166 , \25167 , \25168 , \25169 , \25170 , \25171 , \25172 ,
         \25173 , \25174 , \25175 , \25176 , \25177 , \25178 , \25179 , \25180 , \25181 , \25182 ,
         \25183 , \25184 , \25185 , \25186 , \25187 , \25188 , \25189 , \25190 , \25191 , \25192 ,
         \25193 , \25194 , \25195 , \25196 , \25197 , \25198 , \25199 , \25200 , \25201 , \25202 ,
         \25203 , \25204 , \25205 , \25206 , \25207 , \25208 , \25209 , \25210 , \25211 , \25212 ,
         \25213 , \25214 , \25215 , \25216 , \25217 , \25218 , \25219 , \25220 , \25221 , \25222 ,
         \25223 , \25224 , \25225 , \25226 , \25227 , \25228 , \25229 , \25230 , \25231 , \25232 ,
         \25233 , \25234 , \25235 , \25236 , \25237 , \25238 , \25239 , \25240 , \25241 , \25242 ,
         \25243 , \25244 , \25245 , \25246 , \25247 , \25248 , \25249 , \25250 , \25251 , \25252 ,
         \25253 , \25254 , \25255 , \25256 , \25257 , \25258 , \25259 , \25260 , \25261 , \25262 ,
         \25263 , \25264 , \25265 , \25266 , \25267 , \25268 , \25269 , \25270 , \25271 , \25272 ,
         \25273 , \25274 , \25275 , \25276 , \25277 , \25278 , \25279 , \25280 , \25281 , \25282 ,
         \25283 , \25284 , \25285 , \25286 , \25287 , \25288 , \25289 , \25290 , \25291 , \25292 ,
         \25293 , \25294 , \25295 , \25296 , \25297 , \25298 , \25299 , \25300 , \25301 , \25302 ,
         \25303 , \25304 , \25305 , \25306 , \25307 , \25308 , \25309 , \25310 , \25311 , \25312 ,
         \25313 , \25314 , \25315 , \25316 , \25317 , \25318 , \25319 , \25320 , \25321 , \25322 ,
         \25323 , \25324 , \25325 , \25326 , \25327 , \25328 , \25329 , \25330 , \25331 , \25332 ,
         \25333 , \25334 , \25335 , \25336 , \25337 , \25338 , \25339 , \25340 , \25341 , \25342 ,
         \25343 , \25344 , \25345 , \25346 , \25347 , \25348 , \25349 , \25350 , \25351 , \25352 ,
         \25353 , \25354 , \25355 , \25356 , \25357 , \25358 , \25359 , \25360 , \25361 , \25362 ,
         \25363 , \25364 , \25365 , \25366 , \25367 , \25368 , \25369 , \25370 , \25371 , \25372 ,
         \25373 , \25374 , \25375 , \25376 , \25377 , \25378 , \25379 , \25380 , \25381 , \25382 ,
         \25383 , \25384 , \25385 , \25386 , \25387 , \25388 , \25389 , \25390 , \25391 , \25392 ,
         \25393 , \25394 , \25395 , \25396 , \25397 , \25398 , \25399 , \25400 , \25401 , \25402 ,
         \25403 , \25404 , \25405 , \25406 , \25407 , \25408 , \25409 , \25410 , \25411 , \25412 ,
         \25413 , \25414 , \25415 , \25416 , \25417 , \25418 , \25419 , \25420 , \25421 , \25422 ,
         \25423 , \25424 , \25425 , \25426 , \25427 , \25428 , \25429 , \25430 , \25431 , \25432 ,
         \25433 , \25434 , \25435 , \25436 , \25437 , \25438 , \25439 , \25440 , \25441 , \25442 ,
         \25443 , \25444 , \25445 , \25446 , \25447 , \25448 , \25449 , \25450 , \25451 , \25452 ,
         \25453 , \25454 , \25455 , \25456 , \25457 , \25458 , \25459 , \25460 , \25461 , \25462 ,
         \25463 , \25464 , \25465 , \25466 , \25467 , \25468 , \25469 , \25470 , \25471 , \25472 ,
         \25473 , \25474 , \25475 , \25476 , \25477 , \25478 , \25479 , \25480 , \25481 , \25482 ,
         \25483 , \25484 , \25485 , \25486 , \25487 , \25488 , \25489 , \25490 , \25491 , \25492 ,
         \25493 , \25494 , \25495 , \25496 , \25497 , \25498 , \25499 , \25500 , \25501 , \25502 ,
         \25503 , \25504 , \25505 , \25506 , \25507 , \25508 , \25509 , \25510 , \25511 , \25512 ,
         \25513 , \25514 , \25515 , \25516 , \25517 , \25518 , \25519 , \25520 , \25521 , \25522 ,
         \25523 , \25524 , \25525 , \25526 , \25527 , \25528 , \25529 , \25530 , \25531 , \25532 ,
         \25533 , \25534 , \25535 , \25536 , \25537 , \25538 , \25539 , \25540 , \25541 , \25542 ,
         \25543 , \25544 , \25545 , \25546 , \25547 , \25548 , \25549 , \25550 , \25551 , \25552 ,
         \25553 , \25554 , \25555 , \25556 , \25557 , \25558 , \25559 , \25560 , \25561 , \25562 ,
         \25563 , \25564 , \25565 , \25566 , \25567 , \25568 , \25569 , \25570 , \25571 , \25572 ,
         \25573 , \25574 , \25575 , \25576 , \25577 , \25578 , \25579 , \25580 , \25581 , \25582 ,
         \25583 , \25584 , \25585 , \25586 , \25587 , \25588 , \25589 , \25590 , \25591 , \25592 ,
         \25593 , \25594 , \25595 , \25596 , \25597 , \25598 , \25599 , \25600 , \25601 , \25602 ,
         \25603 , \25604 , \25605 , \25606 , \25607 , \25608 , \25609 , \25610 , \25611 , \25612 ,
         \25613 , \25614 , \25615 , \25616 , \25617 , \25618 , \25619 , \25620 , \25621 , \25622 ,
         \25623 , \25624 , \25625 , \25626 , \25627 , \25628 , \25629 , \25630 , \25631 , \25632 ,
         \25633 , \25634 , \25635 , \25636 , \25637 , \25638 , \25639 , \25640 , \25641 , \25642 ,
         \25643 , \25644 , \25645 , \25646 , \25647 , \25648 , \25649 , \25650 , \25651 , \25652 ,
         \25653 , \25654 , \25655 , \25656 , \25657 , \25658 , \25659 , \25660 , \25661 , \25662 ,
         \25663 , \25664 , \25665 , \25666 , \25667 , \25668 , \25669 , \25670 , \25671 , \25672 ,
         \25673 , \25674 , \25675 , \25676 , \25677 , \25678 , \25679 , \25680 , \25681 , \25682 ,
         \25683 , \25684 , \25685 , \25686 , \25687 , \25688 , \25689 , \25690 , \25691 , \25692 ,
         \25693 , \25694 , \25695 , \25696 , \25697 , \25698 , \25699 , \25700 , \25701 , \25702 ,
         \25703 , \25704 , \25705 , \25706 , \25707 , \25708 , \25709 , \25710 , \25711 , \25712 ,
         \25713 , \25714 , \25715 , \25716 , \25717 , \25718 , \25719 , \25720 , \25721 , \25722 ,
         \25723 , \25724 , \25725 , \25726 , \25727 , \25728 , \25729 , \25730 , \25731 , \25732 ,
         \25733 , \25734 , \25735 , \25736 , \25737 , \25738 , \25739 , \25740 , \25741 , \25742 ,
         \25743 , \25744 , \25745 , \25746 , \25747 , \25748 , \25749 , \25750 , \25751 , \25752 ,
         \25753 , \25754 , \25755 , \25756 , \25757 , \25758 , \25759 , \25760 , \25761 , \25762 ,
         \25763 , \25764 , \25765 , \25766 , \25767 , \25768 , \25769 , \25770 , \25771 , \25772 ,
         \25773 , \25774 , \25775 , \25776 , \25777 , \25778 , \25779 , \25780 , \25781 , \25782 ,
         \25783 , \25784 , \25785 , \25786 , \25787 , \25788 , \25789 , \25790 , \25791 , \25792 ,
         \25793 , \25794 , \25795 , \25796 , \25797 , \25798 , \25799 , \25800 , \25801 , \25802 ,
         \25803 , \25804 , \25805 , \25806 , \25807 , \25808 , \25809 , \25810 , \25811 , \25812 ,
         \25813 , \25814 , \25815 , \25816 , \25817 , \25818 , \25819 , \25820 , \25821 , \25822 ,
         \25823 , \25824 , \25825 , \25826 , \25827 , \25828 , \25829 , \25830 , \25831 , \25832 ,
         \25833 , \25834 , \25835 , \25836 , \25837 , \25838 , \25839 , \25840 , \25841 , \25842 ,
         \25843 , \25844 , \25845 , \25846 , \25847 , \25848 , \25849 , \25850 , \25851 , \25852 ,
         \25853 , \25854 , \25855 , \25856 , \25857 , \25858 , \25859 , \25860 , \25861 , \25862 ,
         \25863 , \25864 , \25865 , \25866 , \25867 , \25868 , \25869 , \25870 , \25871 , \25872 ,
         \25873 , \25874 , \25875 , \25876 , \25877 , \25878 , \25879 , \25880 , \25881 , \25882 ,
         \25883 , \25884 , \25885 , \25886 , \25887 , \25888 , \25889 , \25890 , \25891 , \25892 ,
         \25893 , \25894 , \25895 , \25896 , \25897 , \25898 , \25899 , \25900 , \25901 , \25902 ,
         \25903 , \25904 , \25905 , \25906 , \25907 , \25908 , \25909 , \25910 , \25911 , \25912 ,
         \25913 , \25914 , \25915 , \25916 , \25917 , \25918 , \25919 , \25920 , \25921 , \25922 ,
         \25923 , \25924 , \25925 , \25926 , \25927 , \25928 , \25929 , \25930 , \25931 , \25932 ,
         \25933 , \25934 , \25935 , \25936 , \25937 , \25938 , \25939 , \25940 , \25941 , \25942 ,
         \25943 , \25944 , \25945 , \25946 , \25947 , \25948 , \25949 , \25950 , \25951 , \25952 ,
         \25953 , \25954 , \25955 , \25956 , \25957 , \25958 , \25959 , \25960 , \25961 , \25962 ,
         \25963 , \25964 , \25965 , \25966 , \25967 , \25968 , \25969 , \25970 , \25971 , \25972 ,
         \25973 , \25974 , \25975 , \25976 , \25977 , \25978 , \25979 , \25980 , \25981 , \25982 ,
         \25983 , \25984 , \25985 , \25986 , \25987 , \25988 , \25989 , \25990 , \25991 , \25992 ,
         \25993 , \25994 , \25995 , \25996 , \25997 , \25998 , \25999 , \26000 , \26001 , \26002 ,
         \26003 , \26004 , \26005 , \26006 , \26007 , \26008 , \26009 , \26010 , \26011 , \26012 ,
         \26013 , \26014 , \26015 , \26016 , \26017 , \26018 , \26019 , \26020 , \26021 , \26022 ,
         \26023 , \26024 , \26025 , \26026 , \26027 , \26028 , \26029 , \26030 , \26031 , \26032 ,
         \26033 , \26034 , \26035 , \26036 , \26037 , \26038 , \26039 , \26040 , \26041 , \26042 ,
         \26043 , \26044 , \26045 , \26046 , \26047 , \26048 , \26049 , \26050 , \26051 , \26052 ,
         \26053 , \26054 , \26055 , \26056 , \26057 , \26058 , \26059 , \26060 , \26061 , \26062 ,
         \26063 , \26064 , \26065 , \26066 , \26067 , \26068 , \26069 , \26070 , \26071 , \26072 ,
         \26073 , \26074 , \26075 , \26076 , \26077 , \26078 , \26079 , \26080 , \26081 , \26082 ,
         \26083 , \26084 , \26085 , \26086 , \26087 , \26088 , \26089 , \26090 , \26091 , \26092 ,
         \26093 , \26094 , \26095 , \26096 , \26097 , \26098 , \26099 , \26100 , \26101 , \26102 ,
         \26103 , \26104 , \26105 , \26106 , \26107 , \26108 , \26109 , \26110 , \26111 , \26112 ,
         \26113 , \26114 , \26115 , \26116 , \26117 , \26118 , \26119 , \26120 , \26121 , \26122 ,
         \26123 , \26124 , \26125 , \26126 , \26127 , \26128 , \26129 , \26130 , \26131 , \26132 ,
         \26133 , \26134 , \26135 , \26136 , \26137 , \26138 , \26139 , \26140 , \26141 , \26142 ,
         \26143 , \26144 , \26145 , \26146 , \26147 , \26148 , \26149 , \26150 , \26151 , \26152 ,
         \26153 , \26154 , \26155 , \26156 , \26157 , \26158 , \26159 , \26160 , \26161 , \26162 ,
         \26163 , \26164 , \26165 , \26166 , \26167 , \26168 , \26169 , \26170 , \26171 , \26172 ,
         \26173 , \26174 , \26175 , \26176 , \26177 , \26178 , \26179 , \26180 , \26181 , \26182 ,
         \26183 , \26184 , \26185 , \26186 , \26187 , \26188 , \26189 , \26190 , \26191 , \26192 ,
         \26193 , \26194 , \26195 , \26196 , \26197 , \26198 , \26199 , \26200 , \26201 , \26202 ,
         \26203 , \26204 , \26205 , \26206 , \26207 , \26208 , \26209 , \26210 , \26211 , \26212 ,
         \26213 , \26214 , \26215 , \26216 , \26217 , \26218 , \26219 , \26220 , \26221 , \26222 ,
         \26223 , \26224 , \26225 , \26226 , \26227 , \26228 , \26229 , \26230 , \26231 , \26232 ,
         \26233 , \26234 , \26235 , \26236 , \26237 , \26238 , \26239 , \26240 , \26241 , \26242 ,
         \26243 , \26244 , \26245 , \26246 , \26247 , \26248 , \26249 , \26250 , \26251 , \26252 ,
         \26253 , \26254 , \26255 , \26256 , \26257 , \26258 , \26259 , \26260 , \26261 , \26262 ,
         \26263 , \26264 , \26265 , \26266 , \26267 , \26268 , \26269 , \26270 , \26271 , \26272 ,
         \26273 , \26274 , \26275 , \26276 , \26277 , \26278 , \26279 , \26280 , \26281 , \26282 ,
         \26283 , \26284 , \26285 , \26286 , \26287 , \26288 , \26289 , \26290 , \26291 , \26292 ,
         \26293 , \26294 , \26295 , \26296 , \26297 , \26298 , \26299 , \26300 , \26301 , \26302 ,
         \26303 , \26304 , \26305 , \26306 , \26307 , \26308 , \26309 , \26310 , \26311 , \26312 ,
         \26313 , \26314 , \26315 , \26316 , \26317 , \26318 , \26319 , \26320 , \26321 , \26322 ,
         \26323 , \26324 , \26325 , \26326 , \26327 , \26328 , \26329 , \26330 , \26331 , \26332 ,
         \26333 , \26334 , \26335 , \26336 , \26337 , \26338 , \26339 , \26340 , \26341 , \26342 ,
         \26343 , \26344 , \26345 , \26346 , \26347 , \26348 , \26349 , \26350 , \26351 , \26352 ,
         \26353 , \26354 , \26355 , \26356 , \26357 , \26358 , \26359 , \26360 , \26361 , \26362 ,
         \26363 , \26364 , \26365 , \26366 , \26367 , \26368 , \26369 , \26370 , \26371 , \26372 ,
         \26373 , \26374 , \26375 , \26376 , \26377 , \26378 , \26379 , \26380 , \26381 , \26382 ,
         \26383 , \26384 , \26385 , \26386 , \26387 , \26388 , \26389 , \26390 , \26391 , \26392 ,
         \26393 , \26394 , \26395 , \26396 , \26397 , \26398 , \26399 , \26400 , \26401 , \26402 ,
         \26403 , \26404 , \26405 , \26406 , \26407 , \26408 , \26409 , \26410 , \26411 , \26412 ,
         \26413 , \26414 , \26415 , \26416 , \26417 , \26418 , \26419 , \26420 , \26421 , \26422 ,
         \26423 , \26424 , \26425 , \26426 , \26427 , \26428 , \26429 , \26430 , \26431 , \26432 ,
         \26433 , \26434 , \26435 , \26436 , \26437 , \26438 , \26439 , \26440 , \26441 , \26442 ,
         \26443 , \26444 , \26445 , \26446 , \26447 , \26448 , \26449 , \26450 , \26451 , \26452 ,
         \26453 , \26454 , \26455 , \26456 , \26457 , \26458 , \26459 , \26460 , \26461 , \26462 ,
         \26463 , \26464 , \26465 , \26466 , \26467 , \26468 , \26469 , \26470 , \26471 , \26472 ,
         \26473 , \26474 , \26475 , \26476 , \26477 , \26478 , \26479 , \26480 , \26481 , \26482 ,
         \26483 , \26484 , \26485 , \26486 , \26487 , \26488 , \26489 , \26490 , \26491 , \26492 ,
         \26493 , \26494 , \26495 , \26496 , \26497 , \26498 , \26499 , \26500 , \26501 , \26502 ,
         \26503 , \26504 , \26505 , \26506 , \26507 , \26508 , \26509 , \26510 , \26511 , \26512 ,
         \26513 , \26514 , \26515 , \26516 , \26517 , \26518 , \26519 , \26520 , \26521 , \26522 ,
         \26523 , \26524 , \26525 , \26526 , \26527 , \26528 , \26529 , \26530 , \26531 , \26532 ,
         \26533 , \26534 , \26535 , \26536 , \26537 , \26538 , \26539 , \26540 , \26541 , \26542 ,
         \26543 , \26544 , \26545 , \26546 , \26547 , \26548 , \26549 , \26550 , \26551 , \26552 ,
         \26553 , \26554 , \26555 , \26556 , \26557 , \26558 , \26559 , \26560 , \26561 , \26562 ,
         \26563 , \26564 , \26565 , \26566 , \26567 , \26568 , \26569 , \26570 , \26571 , \26572 ,
         \26573 , \26574 , \26575 , \26576 , \26577 , \26578 , \26579 , \26580 , \26581 , \26582 ,
         \26583 , \26584 , \26585 , \26586 , \26587 , \26588 , \26589 , \26590 , \26591 , \26592 ,
         \26593 , \26594 , \26595 , \26596 , \26597 , \26598 , \26599 , \26600 , \26601 , \26602 ,
         \26603 , \26604 , \26605 , \26606 , \26607 , \26608 , \26609 , \26610 , \26611 , \26612 ,
         \26613 , \26614 , \26615 , \26616 , \26617 , \26618 , \26619 , \26620 , \26621 , \26622 ,
         \26623 , \26624 , \26625 , \26626 , \26627 , \26628 , \26629 , \26630 , \26631 , \26632 ,
         \26633 , \26634 , \26635 , \26636 , \26637 , \26638 , \26639 , \26640 , \26641 , \26642 ,
         \26643 , \26644 , \26645 , \26646 , \26647 , \26648 , \26649 , \26650 , \26651 , \26652 ,
         \26653 , \26654 , \26655 , \26656 , \26657 , \26658 , \26659 , \26660 , \26661 , \26662 ,
         \26663 , \26664 , \26665 , \26666 , \26667 , \26668 , \26669 , \26670 , \26671 , \26672 ,
         \26673 , \26674 , \26675 , \26676 , \26677 , \26678 , \26679 , \26680 , \26681 , \26682 ,
         \26683 , \26684 , \26685 , \26686 , \26687 , \26688 , \26689 , \26690 , \26691 , \26692 ,
         \26693 , \26694 , \26695 , \26696 , \26697 , \26698 , \26699 , \26700 , \26701 , \26702 ,
         \26703 , \26704 , \26705 , \26706 , \26707 , \26708 , \26709 , \26710 , \26711 , \26712 ,
         \26713 , \26714 , \26715 , \26716 , \26717 , \26718 , \26719 , \26720 , \26721 , \26722 ,
         \26723 , \26724 , \26725 , \26726 , \26727 , \26728 , \26729 , \26730 , \26731 , \26732 ,
         \26733 , \26734 , \26735 , \26736 , \26737 , \26738 , \26739 , \26740 , \26741 , \26742 ,
         \26743 , \26744 , \26745 , \26746 , \26747 , \26748 , \26749 , \26750 , \26751 , \26752 ,
         \26753 , \26754 , \26755 , \26756 , \26757 , \26758 , \26759 , \26760 , \26761 , \26762 ,
         \26763 , \26764 , \26765 , \26766 , \26767 , \26768 , \26769 , \26770 , \26771 , \26772 ,
         \26773 , \26774 , \26775 , \26776 , \26777 , \26778 , \26779 , \26780 , \26781 , \26782 ,
         \26783 , \26784 , \26785 , \26786 , \26787 , \26788 , \26789 , \26790 , \26791 , \26792 ,
         \26793 , \26794 , \26795 , \26796 , \26797 , \26798 , \26799 , \26800 , \26801 , \26802 ,
         \26803 , \26804 , \26805 , \26806 , \26807 , \26808 , \26809 , \26810 , \26811 , \26812 ,
         \26813 , \26814 , \26815 , \26816 , \26817 , \26818 , \26819 , \26820 , \26821 , \26822 ,
         \26823 , \26824 , \26825 , \26826 , \26827 , \26828 , \26829 , \26830 , \26831 , \26832 ,
         \26833 , \26834 , \26835 , \26836 , \26837 , \26838 , \26839 , \26840 , \26841 , \26842 ,
         \26843 , \26844 , \26845 , \26846 , \26847 , \26848 , \26849 , \26850 , \26851 , \26852 ,
         \26853 , \26854 , \26855 , \26856 , \26857 , \26858 , \26859 , \26860 , \26861 , \26862 ,
         \26863 , \26864 , \26865 , \26866 , \26867 , \26868 , \26869 , \26870 , \26871 , \26872 ,
         \26873 , \26874 , \26875 , \26876 , \26877 , \26878 , \26879 , \26880 , \26881 , \26882 ,
         \26883 , \26884 , \26885 , \26886 , \26887 , \26888 , \26889 , \26890 , \26891 , \26892 ,
         \26893 , \26894 , \26895 , \26896 , \26897 , \26898 , \26899 , \26900 , \26901 , \26902 ,
         \26903 , \26904 , \26905 , \26906 , \26907 , \26908 , \26909 , \26910 , \26911 , \26912 ,
         \26913 , \26914 , \26915 , \26916 , \26917 , \26918 , \26919 , \26920 , \26921 , \26922 ,
         \26923 , \26924 , \26925 , \26926 , \26927 , \26928 , \26929 , \26930 , \26931 , \26932 ,
         \26933 , \26934 , \26935 , \26936 , \26937 , \26938 , \26939 , \26940 , \26941 , \26942 ,
         \26943 , \26944 , \26945 , \26946 , \26947 , \26948 , \26949 , \26950 , \26951 , \26952 ,
         \26953 , \26954 , \26955 , \26956 , \26957 , \26958 , \26959 , \26960 , \26961 , \26962 ,
         \26963 , \26964 , \26965 , \26966 , \26967 , \26968 , \26969 , \26970 , \26971 , \26972 ,
         \26973 , \26974 , \26975 , \26976 , \26977 , \26978 , \26979 , \26980 , \26981 , \26982 ,
         \26983 , \26984 , \26985 , \26986 , \26987 , \26988 , \26989 , \26990 , \26991 , \26992 ,
         \26993 , \26994 , \26995 , \26996 , \26997 , \26998 , \26999 , \27000 , \27001 , \27002 ,
         \27003 , \27004 , \27005 , \27006 , \27007 , \27008 , \27009 , \27010 , \27011 , \27012 ,
         \27013 , \27014 , \27015 , \27016 , \27017 , \27018 , \27019 , \27020 , \27021 , \27022 ,
         \27023 , \27024 , \27025 , \27026 , \27027 , \27028 , \27029 , \27030 , \27031 , \27032 ,
         \27033 , \27034 , \27035 , \27036 , \27037 , \27038 , \27039 , \27040 , \27041 , \27042 ,
         \27043 , \27044 , \27045 , \27046 , \27047 , \27048 , \27049 , \27050 , \27051 , \27052 ,
         \27053 , \27054 , \27055 , \27056 , \27057 , \27058 , \27059 , \27060 , \27061 , \27062 ,
         \27063 , \27064 , \27065 , \27066 , \27067 , \27068 , \27069 , \27070 , \27071 , \27072 ,
         \27073 , \27074 , \27075 , \27076 , \27077 , \27078 , \27079 , \27080 , \27081 , \27082 ,
         \27083 , \27084 , \27085 , \27086 , \27087 , \27088 , \27089 , \27090 , \27091 , \27092 ,
         \27093 , \27094 , \27095 , \27096 , \27097 , \27098 , \27099 , \27100 , \27101 , \27102 ,
         \27103 , \27104 , \27105 , \27106 , \27107 , \27108 , \27109 , \27110 , \27111 , \27112 ,
         \27113 , \27114 , \27115 , \27116 , \27117 , \27118 , \27119 , \27120 , \27121 , \27122 ,
         \27123 , \27124 , \27125 , \27126 , \27127 , \27128 , \27129 , \27130 , \27131 , \27132 ,
         \27133 , \27134 , \27135 , \27136 , \27137 , \27138 , \27139 , \27140 , \27141 , \27142 ,
         \27143 , \27144 , \27145 , \27146 , \27147 , \27148 , \27149 , \27150 , \27151 , \27152 ,
         \27153 , \27154 , \27155 , \27156 , \27157 , \27158 , \27159 , \27160 , \27161 , \27162 ,
         \27163 , \27164 , \27165 , \27166 , \27167 , \27168 , \27169 , \27170 , \27171 , \27172 ,
         \27173 , \27174 , \27175 , \27176 , \27177 , \27178 , \27179 , \27180 , \27181 , \27182 ,
         \27183 , \27184 , \27185 , \27186 , \27187 , \27188 , \27189 , \27190 , \27191 , \27192 ,
         \27193 , \27194 , \27195 , \27196 , \27197 , \27198 , \27199 , \27200 , \27201 , \27202 ,
         \27203 , \27204 , \27205 , \27206 , \27207 , \27208 , \27209 , \27210 , \27211 , \27212 ,
         \27213 , \27214 , \27215 , \27216 , \27217 , \27218 , \27219 , \27220 , \27221 , \27222 ,
         \27223 , \27224 , \27225 , \27226 , \27227 , \27228 , \27229 , \27230 , \27231 , \27232 ,
         \27233 , \27234 , \27235 , \27236 , \27237 , \27238 , \27239 , \27240 , \27241 , \27242 ,
         \27243 , \27244 , \27245 , \27246 , \27247 , \27248 , \27249 , \27250 , \27251 , \27252 ,
         \27253 , \27254 , \27255 , \27256 , \27257 , \27258 , \27259 , \27260 , \27261 , \27262 ,
         \27263 , \27264 , \27265 , \27266 , \27267 , \27268 , \27269 , \27270 , \27271 , \27272 ,
         \27273 , \27274 , \27275 , \27276 , \27277 , \27278 , \27279 , \27280 , \27281 , \27282 ,
         \27283 , \27284 , \27285 , \27286 , \27287 , \27288 , \27289 , \27290 , \27291 , \27292 ,
         \27293 , \27294 , \27295 , \27296 , \27297 , \27298 , \27299 , \27300 , \27301 , \27302 ,
         \27303 , \27304 , \27305 , \27306 , \27307 , \27308 , \27309 , \27310 , \27311 , \27312 ,
         \27313 , \27314 , \27315 , \27316 , \27317 , \27318 , \27319 , \27320 , \27321 , \27322 ,
         \27323 , \27324 , \27325 , \27326 , \27327 , \27328 , \27329 , \27330 , \27331 , \27332 ,
         \27333 , \27334 , \27335 , \27336 , \27337 , \27338 , \27339 , \27340 , \27341 , \27342 ,
         \27343 , \27344 , \27345 , \27346 , \27347 , \27348 , \27349 , \27350 , \27351 , \27352 ,
         \27353 , \27354 , \27355 , \27356 , \27357 , \27358 , \27359 , \27360 , \27361 , \27362 ,
         \27363 , \27364 , \27365 , \27366 , \27367 , \27368 , \27369 , \27370 , \27371 , \27372 ,
         \27373 , \27374 , \27375 , \27376 , \27377 , \27378 , \27379 , \27380 , \27381 , \27382 ,
         \27383 , \27384 , \27385 , \27386 , \27387 , \27388 , \27389 , \27390 , \27391 , \27392 ,
         \27393 , \27394 , \27395 , \27396 , \27397 , \27398 , \27399 , \27400 , \27401 , \27402 ,
         \27403 , \27404 , \27405 , \27406 , \27407 , \27408 , \27409 , \27410 , \27411 , \27412 ,
         \27413 , \27414 , \27415 , \27416 , \27417 , \27418 , \27419 , \27420 , \27421 , \27422 ,
         \27423 , \27424 , \27425 , \27426 , \27427 , \27428 , \27429 , \27430 , \27431 , \27432 ,
         \27433 , \27434 , \27435 , \27436 , \27437 , \27438 , \27439 , \27440 , \27441 , \27442 ,
         \27443 , \27444 , \27445 , \27446 , \27447 , \27448 , \27449 , \27450 , \27451 , \27452 ,
         \27453 , \27454 , \27455 , \27456 , \27457 , \27458 , \27459 , \27460 , \27461 , \27462 ,
         \27463 , \27464 , \27465 , \27466 , \27467 , \27468 , \27469 , \27470 , \27471 , \27472 ,
         \27473 , \27474 , \27475 , \27476 , \27477 , \27478 , \27479 , \27480 , \27481 , \27482 ,
         \27483 , \27484 , \27485 , \27486 , \27487 , \27488 , \27489 , \27490 , \27491 , \27492 ,
         \27493 , \27494 , \27495 , \27496 , \27497 , \27498 , \27499 , \27500 , \27501 , \27502 ,
         \27503 , \27504 , \27505 , \27506 , \27507 , \27508 , \27509 , \27510 , \27511 , \27512 ,
         \27513 , \27514 , \27515 , \27516 , \27517 , \27518 , \27519 , \27520 , \27521 , \27522 ,
         \27523 , \27524 , \27525 , \27526 , \27527 , \27528 , \27529 , \27530 , \27531 , \27532 ,
         \27533 , \27534 , \27535 , \27536 , \27537 , \27538 , \27539 , \27540 , \27541 , \27542 ,
         \27543 , \27544 , \27545 , \27546 , \27547 , \27548 , \27549 , \27550 , \27551 , \27552 ,
         \27553 , \27554 , \27555 , \27556 , \27557 , \27558 , \27559 , \27560 , \27561 , \27562 ,
         \27563 , \27564 , \27565 , \27566 , \27567 , \27568 , \27569 , \27570 , \27571 , \27572 ,
         \27573 , \27574 , \27575 , \27576 , \27577 , \27578 , \27579 , \27580 , \27581 , \27582 ,
         \27583 , \27584 , \27585 , \27586 , \27587 , \27588 , \27589 , \27590 , \27591 , \27592 ,
         \27593 , \27594 , \27595 , \27596 , \27597 , \27598 , \27599 , \27600 , \27601 , \27602 ,
         \27603 , \27604 , \27605 , \27606 , \27607 , \27608 , \27609 , \27610 , \27611 , \27612 ,
         \27613 , \27614 , \27615 , \27616 , \27617 , \27618 , \27619 , \27620 , \27621 , \27622 ,
         \27623 , \27624 , \27625 , \27626 , \27627 , \27628 , \27629 , \27630 , \27631 , \27632 ,
         \27633 , \27634 , \27635 , \27636 , \27637 , \27638 , \27639 , \27640 , \27641 , \27642 ,
         \27643 , \27644 , \27645 , \27646 , \27647 , \27648 , \27649 , \27650 , \27651 , \27652 ,
         \27653 , \27654 , \27655 , \27656 , \27657 , \27658 , \27659 , \27660 , \27661 , \27662 ,
         \27663 , \27664 , \27665 , \27666 , \27667 , \27668 , \27669 , \27670 , \27671 , \27672 ,
         \27673 , \27674 , \27675 , \27676 , \27677 , \27678 , \27679 , \27680 , \27681 , \27682 ,
         \27683 , \27684 , \27685 , \27686 , \27687 , \27688 , \27689 , \27690 , \27691 , \27692 ,
         \27693 , \27694 , \27695 , \27696 , \27697 , \27698 , \27699 , \27700 , \27701 , \27702 ,
         \27703 , \27704 , \27705 , \27706 , \27707 , \27708 , \27709 , \27710 , \27711 , \27712 ,
         \27713 , \27714 , \27715 , \27716 , \27717 , \27718 , \27719 , \27720 , \27721 , \27722 ,
         \27723 , \27724 , \27725 , \27726 , \27727 , \27728 , \27729 , \27730 , \27731 , \27732 ,
         \27733 , \27734 , \27735 , \27736 , \27737 , \27738 , \27739 , \27740 , \27741 , \27742 ,
         \27743 , \27744 , \27745 , \27746 , \27747 , \27748 , \27749 , \27750 , \27751 , \27752 ,
         \27753 , \27754 , \27755 , \27756 , \27757 , \27758 , \27759 , \27760 , \27761 , \27762 ,
         \27763 , \27764 , \27765 , \27766 , \27767 , \27768 , \27769 , \27770 , \27771 , \27772 ,
         \27773 , \27774 , \27775 , \27776 , \27777 , \27778 , \27779 , \27780 , \27781 , \27782 ,
         \27783 , \27784 , \27785 , \27786 , \27787 , \27788 , \27789 , \27790 , \27791 , \27792 ,
         \27793 , \27794 , \27795 , \27796 , \27797 , \27798 , \27799 , \27800 , \27801 , \27802 ,
         \27803 , \27804 , \27805 , \27806 , \27807 , \27808 , \27809 , \27810 , \27811 , \27812 ,
         \27813 , \27814 , \27815 , \27816 , \27817 , \27818 , \27819 , \27820 , \27821 , \27822 ,
         \27823 , \27824 , \27825 , \27826 , \27827 , \27828 , \27829 , \27830 , \27831 , \27832 ,
         \27833 , \27834 , \27835 , \27836 , \27837 , \27838 , \27839 , \27840 , \27841 , \27842 ,
         \27843 , \27844 , \27845 , \27846 , \27847 , \27848 , \27849 , \27850 , \27851 , \27852 ,
         \27853 , \27854 , \27855 , \27856 , \27857 , \27858 , \27859 , \27860 , \27861 , \27862 ,
         \27863 , \27864 , \27865 , \27866 , \27867 , \27868 , \27869 , \27870 , \27871 , \27872 ,
         \27873 , \27874 , \27875 , \27876 , \27877 , \27878 , \27879 , \27880 , \27881 , \27882 ,
         \27883 , \27884 , \27885 , \27886 , \27887 , \27888 , \27889 , \27890 , \27891 , \27892 ,
         \27893 , \27894 , \27895 , \27896 , \27897 , \27898 , \27899 , \27900 , \27901 , \27902 ,
         \27903 , \27904 , \27905 , \27906 , \27907 , \27908 , \27909 , \27910 , \27911 , \27912 ,
         \27913 , \27914 , \27915 , \27916 , \27917 , \27918 , \27919 , \27920 , \27921 , \27922 ,
         \27923 , \27924 , \27925 , \27926 , \27927 , \27928 , \27929 , \27930 , \27931 , \27932 ,
         \27933 , \27934 , \27935 , \27936 , \27937 , \27938 , \27939 , \27940 , \27941 , \27942 ,
         \27943 , \27944 , \27945 , \27946 , \27947 , \27948 , \27949 , \27950 , \27951 , \27952 ,
         \27953 , \27954 , \27955 , \27956 , \27957 , \27958 , \27959 , \27960 , \27961 , \27962 ,
         \27963 , \27964 , \27965 , \27966 , \27967 , \27968 , \27969 , \27970 , \27971 , \27972 ,
         \27973 , \27974 , \27975 , \27976 , \27977 , \27978 , \27979 , \27980 , \27981 , \27982 ,
         \27983 , \27984 , \27985 , \27986 , \27987 , \27988 , \27989 , \27990 , \27991 , \27992 ,
         \27993 , \27994 , \27995 , \27996 , \27997 , \27998 , \27999 , \28000 , \28001 , \28002 ,
         \28003 , \28004 , \28005 , \28006 , \28007 , \28008 , \28009 , \28010 , \28011 , \28012 ,
         \28013 , \28014 , \28015 , \28016 , \28017 , \28018 , \28019 , \28020 , \28021 , \28022 ,
         \28023 , \28024 , \28025 , \28026 , \28027 , \28028 , \28029 , \28030 , \28031 , \28032 ,
         \28033 , \28034 , \28035 , \28036 , \28037 , \28038 , \28039 , \28040 , \28041 , \28042 ,
         \28043 , \28044 , \28045 , \28046 , \28047 , \28048 , \28049 , \28050 , \28051 , \28052 ,
         \28053 , \28054 , \28055 , \28056 , \28057 , \28058 , \28059 , \28060 , \28061 , \28062 ,
         \28063 , \28064 , \28065 , \28066 , \28067 , \28068 , \28069 , \28070 , \28071 , \28072 ,
         \28073 , \28074 , \28075 , \28076 , \28077 , \28078 , \28079 , \28080 , \28081 , \28082 ,
         \28083 , \28084 , \28085 , \28086 , \28087 , \28088 , \28089 , \28090 , \28091 , \28092 ,
         \28093 , \28094 , \28095 , \28096 , \28097 , \28098 , \28099 , \28100 , \28101 , \28102 ,
         \28103 , \28104 , \28105 , \28106 , \28107 , \28108 , \28109 , \28110 , \28111 , \28112 ,
         \28113 , \28114 , \28115 , \28116 , \28117 , \28118 , \28119 , \28120 , \28121 , \28122 ,
         \28123 , \28124 , \28125 , \28126 , \28127 , \28128 , \28129 , \28130 , \28131 , \28132 ,
         \28133 , \28134 , \28135 , \28136 , \28137 , \28138 , \28139 , \28140 , \28141 , \28142 ,
         \28143 , \28144 , \28145 , \28146 , \28147 , \28148 , \28149 , \28150 , \28151 , \28152 ,
         \28153 , \28154 , \28155 , \28156 , \28157 , \28158 , \28159 , \28160 , \28161 , \28162 ,
         \28163 , \28164 , \28165 , \28166 , \28167 , \28168 , \28169 , \28170 , \28171 , \28172 ,
         \28173 , \28174 , \28175 , \28176 , \28177 , \28178 , \28179 , \28180 , \28181 , \28182 ,
         \28183 , \28184 , \28185 , \28186 , \28187 , \28188 , \28189 , \28190 , \28191 , \28192 ,
         \28193 , \28194 , \28195 , \28196 , \28197 , \28198 , \28199 , \28200 , \28201 , \28202 ,
         \28203 , \28204 , \28205 , \28206 , \28207 , \28208 , \28209 , \28210 , \28211 , \28212 ,
         \28213 , \28214 , \28215 , \28216 , \28217 , \28218 , \28219 , \28220 , \28221 , \28222 ,
         \28223 , \28224 , \28225 , \28226 , \28227 , \28228 , \28229 , \28230 , \28231 , \28232 ,
         \28233 , \28234 , \28235 , \28236 , \28237 , \28238 , \28239 , \28240 , \28241 , \28242 ,
         \28243 , \28244 , \28245 , \28246 , \28247 , \28248 , \28249 , \28250 , \28251 , \28252 ,
         \28253 , \28254 , \28255 , \28256 , \28257 , \28258 , \28259 , \28260 , \28261 , \28262 ,
         \28263 , \28264 , \28265 , \28266 , \28267 , \28268 , \28269 , \28270 , \28271 , \28272 ,
         \28273 , \28274 , \28275 , \28276 , \28277 , \28278 , \28279 , \28280 , \28281 , \28282 ,
         \28283 , \28284 , \28285 , \28286 , \28287 , \28288 , \28289 , \28290 , \28291 , \28292 ,
         \28293 , \28294 , \28295 , \28296 , \28297 , \28298 , \28299 , \28300 , \28301 , \28302 ,
         \28303 , \28304 , \28305 , \28306 , \28307 , \28308 , \28309 , \28310 , \28311 , \28312 ,
         \28313 , \28314 , \28315 , \28316 , \28317 , \28318 , \28319 , \28320 , \28321 , \28322 ,
         \28323 , \28324 , \28325 , \28326 , \28327 , \28328 , \28329 , \28330 , \28331 , \28332 ,
         \28333 , \28334 , \28335 , \28336 , \28337 , \28338 , \28339 , \28340 , \28341 , \28342 ,
         \28343 , \28344 , \28345 , \28346 , \28347 , \28348 , \28349 , \28350 , \28351 , \28352 ,
         \28353 , \28354 , \28355 , \28356 , \28357 , \28358 , \28359 , \28360 , \28361 , \28362 ,
         \28363 , \28364 , \28365 , \28366 , \28367 , \28368 , \28369 , \28370 , \28371 , \28372 ,
         \28373 , \28374 , \28375 , \28376 , \28377 , \28378 , \28379 , \28380 , \28381 , \28382 ,
         \28383 , \28384 , \28385 , \28386 , \28387 , \28388 , \28389 , \28390 , \28391 , \28392 ,
         \28393 , \28394 , \28395 , \28396 , \28397 , \28398 , \28399 , \28400 , \28401 , \28402 ,
         \28403 , \28404 , \28405 , \28406 , \28407 , \28408 , \28409 , \28410 , \28411 , \28412 ,
         \28413 , \28414 , \28415 , \28416 , \28417 , \28418 , \28419 , \28420 , \28421 , \28422 ,
         \28423 , \28424 , \28425 , \28426 , \28427 , \28428 , \28429 , \28430 , \28431 , \28432 ,
         \28433 , \28434 , \28435 , \28436 , \28437 , \28438 , \28439 , \28440 , \28441 , \28442 ,
         \28443 , \28444 , \28445 , \28446 , \28447 , \28448 , \28449 , \28450 , \28451 , \28452 ,
         \28453 , \28454 , \28455 , \28456 , \28457 , \28458 , \28459 , \28460 , \28461 , \28462 ,
         \28463 , \28464 , \28465 , \28466 , \28467 , \28468 , \28469 , \28470 , \28471 , \28472 ,
         \28473 , \28474 , \28475 , \28476 , \28477 , \28478 , \28479 , \28480 , \28481 , \28482 ,
         \28483 , \28484 , \28485 , \28486 , \28487 , \28488 , \28489 , \28490 , \28491 , \28492 ,
         \28493 , \28494 , \28495 , \28496 , \28497 , \28498 , \28499 , \28500 , \28501 , \28502 ,
         \28503 , \28504 , \28505 , \28506 , \28507 , \28508 , \28509 , \28510 , \28511 , \28512 ,
         \28513 , \28514 , \28515 , \28516 , \28517 , \28518 , \28519 , \28520 , \28521 , \28522 ,
         \28523 , \28524 , \28525 , \28526 , \28527 , \28528 , \28529 , \28530 , \28531 , \28532 ,
         \28533 , \28534 , \28535 , \28536 , \28537 , \28538 , \28539 , \28540 , \28541 , \28542 ,
         \28543 , \28544 , \28545 , \28546 , \28547 , \28548 , \28549 , \28550 , \28551 , \28552 ,
         \28553 , \28554 , \28555 , \28556 , \28557 , \28558 , \28559 , \28560 , \28561 , \28562 ,
         \28563 , \28564 , \28565 , \28566 , \28567 , \28568 , \28569 , \28570 , \28571 , \28572 ,
         \28573 , \28574 , \28575 , \28576 , \28577 , \28578 , \28579 , \28580 , \28581 , \28582 ,
         \28583 , \28584 , \28585 , \28586 , \28587 , \28588 , \28589 , \28590 , \28591 , \28592 ,
         \28593 , \28594 , \28595 , \28596 , \28597 , \28598 , \28599 , \28600 , \28601 , \28602 ,
         \28603 , \28604 , \28605 , \28606 , \28607 , \28608 , \28609 , \28610 , \28611 , \28612 ,
         \28613 , \28614 , \28615 , \28616 , \28617 , \28618 , \28619 , \28620 , \28621 , \28622 ,
         \28623 , \28624 , \28625 , \28626 , \28627 , \28628 , \28629 , \28630 , \28631 , \28632 ,
         \28633 , \28634 , \28635 , \28636 , \28637 , \28638 , \28639 , \28640 , \28641 , \28642 ,
         \28643 , \28644 , \28645 , \28646 , \28647 , \28648 , \28649 , \28650 , \28651 , \28652 ,
         \28653 , \28654 , \28655 , \28656 , \28657 , \28658 , \28659 , \28660 , \28661 , \28662 ,
         \28663 , \28664 , \28665 , \28666 , \28667 , \28668 , \28669 , \28670 , \28671 , \28672 ,
         \28673 , \28674 , \28675 , \28676 , \28677 , \28678 , \28679 , \28680 , \28681 , \28682 ,
         \28683 , \28684 , \28685 , \28686 , \28687 , \28688 , \28689 , \28690 , \28691 , \28692 ,
         \28693 , \28694 , \28695 , \28696 , \28697 , \28698 , \28699 , \28700 , \28701 , \28702 ,
         \28703 , \28704 , \28705 , \28706 , \28707 , \28708 , \28709 , \28710 , \28711 , \28712 ,
         \28713 , \28714 , \28715 , \28716 , \28717 , \28718 , \28719 , \28720 , \28721 , \28722 ,
         \28723 , \28724 , \28725 , \28726 , \28727 , \28728 , \28729 , \28730 , \28731 , \28732 ,
         \28733 , \28734 , \28735 , \28736 , \28737 , \28738 , \28739 , \28740 , \28741 , \28742 ,
         \28743 , \28744 , \28745 , \28746 , \28747 , \28748 , \28749 , \28750 , \28751 , \28752 ,
         \28753 , \28754 , \28755 , \28756 , \28757 , \28758 , \28759 , \28760 , \28761 , \28762 ,
         \28763 , \28764 , \28765 , \28766 , \28767 , \28768 , \28769 , \28770 , \28771 , \28772 ,
         \28773 , \28774 , \28775 , \28776 , \28777 , \28778 , \28779 , \28780 , \28781 , \28782 ,
         \28783 , \28784 , \28785 , \28786 , \28787 , \28788 , \28789 , \28790 , \28791 , \28792 ,
         \28793 , \28794 , \28795 , \28796 , \28797 , \28798 , \28799 , \28800 , \28801 , \28802 ,
         \28803 , \28804 , \28805 , \28806 , \28807 , \28808 , \28809 , \28810 , \28811 , \28812 ,
         \28813 , \28814 , \28815 , \28816 , \28817 , \28818 , \28819 , \28820 , \28821 , \28822 ,
         \28823 , \28824 , \28825 , \28826 , \28827 , \28828 , \28829 , \28830 , \28831 , \28832 ,
         \28833 , \28834 , \28835 , \28836 , \28837 , \28838 , \28839 , \28840 , \28841 , \28842 ,
         \28843 , \28844 , \28845 , \28846 , \28847 , \28848 , \28849 , \28850 , \28851 , \28852 ,
         \28853 , \28854 , \28855 , \28856 , \28857 , \28858 , \28859 , \28860 , \28861 , \28862 ,
         \28863 , \28864 , \28865 , \28866 , \28867 , \28868 , \28869 , \28870 , \28871 , \28872 ,
         \28873 , \28874 , \28875 , \28876 , \28877 , \28878 , \28879 , \28880 , \28881 , \28882 ,
         \28883 , \28884 , \28885 , \28886 , \28887 , \28888 , \28889 , \28890 , \28891 , \28892 ,
         \28893 , \28894 , \28895 , \28896 , \28897 , \28898 , \28899 , \28900 , \28901 , \28902 ,
         \28903 , \28904 , \28905 , \28906 , \28907 , \28908 , \28909 , \28910 , \28911 , \28912 ,
         \28913 , \28914 , \28915 , \28916 , \28917 , \28918 , \28919 , \28920 , \28921 , \28922 ,
         \28923 , \28924 , \28925 , \28926 , \28927 , \28928 , \28929 , \28930 , \28931 , \28932 ,
         \28933 , \28934 , \28935 , \28936 , \28937 , \28938 , \28939 , \28940 , \28941 , \28942 ,
         \28943 , \28944 , \28945 , \28946 , \28947 , \28948 , \28949 , \28950 , \28951 , \28952 ,
         \28953 , \28954 , \28955 , \28956 , \28957 , \28958 , \28959 , \28960 , \28961 , \28962 ,
         \28963 , \28964 , \28965 , \28966 , \28967 , \28968 , \28969 , \28970 , \28971 , \28972 ,
         \28973 , \28974 , \28975 , \28976 , \28977 , \28978 , \28979 , \28980 , \28981 , \28982 ,
         \28983 , \28984 , \28985 , \28986 , \28987 , \28988 , \28989 , \28990 , \28991 , \28992 ,
         \28993 , \28994 , \28995 , \28996 , \28997 , \28998 , \28999 , \29000 , \29001 , \29002 ,
         \29003 , \29004 , \29005 , \29006 , \29007 , \29008 , \29009 , \29010 , \29011 , \29012 ,
         \29013 , \29014 , \29015 , \29016 , \29017 , \29018 , \29019 , \29020 , \29021 , \29022 ,
         \29023 , \29024 , \29025 , \29026 , \29027 , \29028 , \29029 , \29030 , \29031 , \29032 ,
         \29033 , \29034 , \29035 , \29036 , \29037 , \29038 , \29039 , \29040 , \29041 , \29042 ,
         \29043 , \29044 , \29045 , \29046 , \29047 , \29048 , \29049 , \29050 , \29051 , \29052 ,
         \29053 , \29054 , \29055 , \29056 , \29057 , \29058 , \29059 , \29060 , \29061 , \29062 ,
         \29063 , \29064 , \29065 , \29066 , \29067 , \29068 , \29069 , \29070 , \29071 , \29072 ,
         \29073 , \29074 , \29075 , \29076 , \29077 , \29078 , \29079 , \29080 , \29081 , \29082 ,
         \29083 , \29084 , \29085 , \29086 , \29087 , \29088 , \29089 , \29090 , \29091 , \29092 ,
         \29093 , \29094 , \29095 , \29096 , \29097 , \29098 , \29099 , \29100 , \29101 , \29102 ,
         \29103 , \29104 , \29105 , \29106 , \29107 , \29108 , \29109 , \29110 , \29111 , \29112 ,
         \29113 , \29114 , \29115 , \29116 , \29117 , \29118 , \29119 , \29120 , \29121 , \29122 ,
         \29123 , \29124 , \29125 , \29126 , \29127 , \29128 , \29129 , \29130 , \29131 , \29132 ,
         \29133 , \29134 , \29135 , \29136 , \29137 , \29138 , \29139 , \29140 , \29141 , \29142 ,
         \29143 , \29144 , \29145 , \29146 , \29147 , \29148 , \29149 , \29150 , \29151 , \29152 ,
         \29153 , \29154 , \29155 , \29156 , \29157 , \29158 , \29159 , \29160 , \29161 , \29162 ,
         \29163 , \29164 , \29165 , \29166 , \29167 , \29168 , \29169 , \29170 , \29171 , \29172 ,
         \29173 , \29174 , \29175 , \29176 , \29177 , \29178 , \29179 , \29180 , \29181 , \29182 ,
         \29183 , \29184 , \29185 , \29186 , \29187 , \29188 , \29189 , \29190 , \29191 , \29192 ,
         \29193 , \29194 , \29195 , \29196 , \29197 , \29198 , \29199 , \29200 , \29201 , \29202 ,
         \29203 , \29204 , \29205 , \29206 , \29207 , \29208 , \29209 , \29210 , \29211 , \29212 ,
         \29213 , \29214 , \29215 , \29216 , \29217 , \29218 , \29219 , \29220 , \29221 , \29222 ,
         \29223 , \29224 , \29225 , \29226 , \29227 , \29228 , \29229 , \29230 , \29231 , \29232 ,
         \29233 , \29234 , \29235 , \29236 , \29237 , \29238 , \29239 , \29240 , \29241 , \29242 ,
         \29243 , \29244 , \29245 , \29246 , \29247 , \29248 , \29249 , \29250 , \29251 , \29252 ,
         \29253 , \29254 , \29255 , \29256 , \29257 , \29258 , \29259 , \29260 , \29261 , \29262 ,
         \29263 , \29264 , \29265 , \29266 , \29267 , \29268 , \29269 , \29270 , \29271 , \29272 ,
         \29273 , \29274 , \29275 , \29276 , \29277 , \29278 , \29279 , \29280 , \29281 , \29282 ,
         \29283 , \29284 , \29285 , \29286 , \29287 , \29288 , \29289 , \29290 , \29291 , \29292 ,
         \29293 , \29294 , \29295 , \29296 , \29297 , \29298 , \29299 , \29300 , \29301 , \29302 ,
         \29303 , \29304 , \29305 , \29306 , \29307 , \29308 , \29309 , \29310 , \29311 , \29312 ,
         \29313 , \29314 , \29315 , \29316 , \29317 , \29318 , \29319 , \29320 , \29321 , \29322 ,
         \29323 , \29324 , \29325 , \29326 , \29327 , \29328 , \29329 , \29330 , \29331 , \29332 ,
         \29333 , \29334 , \29335 , \29336 , \29337 , \29338 , \29339 , \29340 , \29341 , \29342 ,
         \29343 , \29344 , \29345 , \29346 , \29347 , \29348 , \29349 , \29350 , \29351 , \29352 ,
         \29353 , \29354 , \29355 , \29356 , \29357 , \29358 , \29359 , \29360 , \29361 , \29362 ,
         \29363 , \29364 , \29365 , \29366 , \29367 , \29368 , \29369 , \29370 , \29371 , \29372 ,
         \29373 , \29374 , \29375 , \29376 , \29377 , \29378 , \29379 , \29380 , \29381 , \29382 ,
         \29383 , \29384 , \29385 , \29386 , \29387 , \29388 , \29389 , \29390 , \29391 , \29392 ,
         \29393 , \29394 , \29395 , \29396 , \29397 , \29398 , \29399 , \29400 , \29401 , \29402 ,
         \29403 , \29404 , \29405 , \29406 , \29407 , \29408 , \29409 , \29410 , \29411 , \29412 ,
         \29413 , \29414 , \29415 , \29416 , \29417 , \29418 , \29419 , \29420 , \29421 , \29422 ,
         \29423 , \29424 , \29425 , \29426 , \29427 , \29428 , \29429 , \29430 , \29431 , \29432 ,
         \29433 , \29434 , \29435 , \29436 , \29437 , \29438 , \29439 , \29440 , \29441 , \29442 ,
         \29443 , \29444 , \29445 , \29446 , \29447 , \29448 , \29449 , \29450 , \29451 , \29452 ,
         \29453 , \29454 , \29455 , \29456 , \29457 , \29458 , \29459 , \29460 , \29461 , \29462 ,
         \29463 , \29464 , \29465 , \29466 , \29467 , \29468 , \29469 , \29470 , \29471 , \29472 ,
         \29473 , \29474 , \29475 , \29476 , \29477 , \29478 , \29479 , \29480 , \29481 , \29482 ,
         \29483 , \29484 , \29485 , \29486 , \29487 , \29488 , \29489 , \29490 , \29491 , \29492 ,
         \29493 , \29494 , \29495 , \29496 , \29497 , \29498 , \29499 , \29500 , \29501 , \29502 ,
         \29503 , \29504 , \29505 , \29506 , \29507 , \29508 , \29509 , \29510 , \29511 , \29512 ,
         \29513 , \29514 , \29515 , \29516 , \29517 , \29518 , \29519 , \29520 , \29521 , \29522 ,
         \29523 , \29524 , \29525 , \29526 , \29527 , \29528 , \29529 , \29530 , \29531 , \29532 ,
         \29533 , \29534 , \29535 , \29536 , \29537 , \29538 , \29539 , \29540 , \29541 , \29542 ,
         \29543 , \29544 , \29545 , \29546 , \29547 , \29548 , \29549 , \29550 , \29551 , \29552 ,
         \29553 , \29554 , \29555 , \29556 , \29557 , \29558 , \29559 , \29560 , \29561 , \29562 ,
         \29563 , \29564 , \29565 , \29566 , \29567 , \29568 , \29569 , \29570 , \29571 , \29572 ,
         \29573 , \29574 , \29575 , \29576 , \29577 , \29578 , \29579 , \29580 , \29581 , \29582 ,
         \29583 , \29584 , \29585 , \29586 , \29587 , \29588 , \29589 , \29590 , \29591 , \29592 ,
         \29593 , \29594 , \29595 , \29596 , \29597 , \29598 , \29599 , \29600 , \29601 , \29602 ,
         \29603 , \29604 , \29605 , \29606 , \29607 , \29608 , \29609 , \29610 , \29611 , \29612 ,
         \29613 , \29614 , \29615 , \29616 , \29617 , \29618 , \29619 , \29620 , \29621 , \29622 ,
         \29623 , \29624 , \29625 , \29626 , \29627 , \29628 , \29629 , \29630 , \29631 , \29632 ,
         \29633 , \29634 , \29635 , \29636 , \29637 , \29638 , \29639 , \29640 , \29641 , \29642 ,
         \29643 , \29644 , \29645 , \29646 , \29647 , \29648 , \29649 , \29650 , \29651 , \29652 ,
         \29653 , \29654 , \29655 , \29656 , \29657 , \29658 , \29659 , \29660 , \29661 , \29662 ,
         \29663 , \29664 , \29665 , \29666 , \29667 , \29668 , \29669 , \29670 , \29671 , \29672 ,
         \29673 , \29674 , \29675 , \29676 , \29677 , \29678 , \29679 , \29680 , \29681 , \29682 ,
         \29683 , \29684 , \29685 , \29686 , \29687 , \29688 , \29689 , \29690 , \29691 , \29692 ,
         \29693 , \29694 , \29695 , \29696 , \29697 , \29698 , \29699 , \29700 , \29701 , \29702 ,
         \29703 , \29704 , \29705 , \29706 , \29707 , \29708 , \29709 , \29710 , \29711 , \29712 ,
         \29713 , \29714 , \29715 , \29716 , \29717 , \29718 , \29719 , \29720 , \29721 , \29722 ,
         \29723 , \29724 , \29725 , \29726 , \29727 , \29728 , \29729 , \29730 , \29731 , \29732 ,
         \29733 , \29734 , \29735 , \29736 , \29737 , \29738 , \29739 , \29740 , \29741 , \29742 ,
         \29743 , \29744 , \29745 , \29746 , \29747 , \29748 , \29749 , \29750 , \29751 , \29752 ,
         \29753 , \29754 , \29755 , \29756 , \29757 , \29758 , \29759 , \29760 , \29761 , \29762 ,
         \29763 , \29764 , \29765 , \29766 , \29767 , \29768 , \29769 , \29770 , \29771 , \29772 ,
         \29773 , \29774 , \29775 , \29776 , \29777 , \29778 , \29779 , \29780 , \29781 , \29782 ,
         \29783 , \29784 , \29785 , \29786 , \29787 , \29788 , \29789 , \29790 , \29791 , \29792 ,
         \29793 , \29794 , \29795 , \29796 , \29797 , \29798 , \29799 , \29800 , \29801 , \29802 ,
         \29803 , \29804 , \29805 , \29806 , \29807 , \29808 , \29809 , \29810 , \29811 , \29812 ,
         \29813 , \29814 , \29815 , \29816 , \29817 , \29818 , \29819 , \29820 , \29821 , \29822 ,
         \29823 , \29824 , \29825 , \29826 , \29827 , \29828 , \29829 , \29830 , \29831 , \29832 ,
         \29833 , \29834 , \29835 , \29836 , \29837 , \29838 , \29839 , \29840 , \29841 , \29842 ,
         \29843 , \29844 , \29845 , \29846 , \29847 , \29848 , \29849 , \29850 , \29851 , \29852 ,
         \29853 , \29854 , \29855 , \29856 , \29857 , \29858 , \29859 , \29860 , \29861 , \29862 ,
         \29863 , \29864 , \29865 , \29866 , \29867 , \29868 , \29869 , \29870 , \29871 , \29872 ,
         \29873 , \29874 , \29875 , \29876 , \29877 , \29878 , \29879 , \29880 , \29881 , \29882 ,
         \29883 , \29884 , \29885 , \29886 , \29887 , \29888 , \29889 , \29890 , \29891 , \29892 ,
         \29893 , \29894 , \29895 , \29896 , \29897 , \29898 , \29899 , \29900 , \29901 , \29902 ,
         \29903 , \29904 , \29905 , \29906 , \29907 , \29908 , \29909 , \29910 , \29911 , \29912 ,
         \29913 , \29914 , \29915 , \29916 , \29917 , \29918 , \29919 , \29920 , \29921 , \29922 ,
         \29923 , \29924 , \29925 , \29926 , \29927 , \29928 , \29929 , \29930 , \29931 , \29932 ,
         \29933 , \29934 , \29935 , \29936 , \29937 , \29938 , \29939 , \29940 , \29941 , \29942 ,
         \29943 , \29944 , \29945 , \29946 , \29947 , \29948 , \29949 , \29950 , \29951 , \29952 ,
         \29953 , \29954 , \29955 , \29956 , \29957 , \29958 , \29959 , \29960 , \29961 , \29962 ,
         \29963 , \29964 , \29965 , \29966 , \29967 , \29968 , \29969 , \29970 , \29971 , \29972 ,
         \29973 , \29974 , \29975 , \29976 , \29977 , \29978 , \29979 , \29980 , \29981 , \29982 ,
         \29983 , \29984 , \29985 , \29986 , \29987 , \29988 , \29989 , \29990 , \29991 , \29992 ,
         \29993 , \29994 , \29995 , \29996 , \29997 , \29998 , \29999 , \30000 , \30001 , \30002 ,
         \30003 , \30004 , \30005 , \30006 , \30007 , \30008 , \30009 , \30010 , \30011 , \30012 ,
         \30013 , \30014 , \30015 , \30016 , \30017 , \30018 , \30019 , \30020 , \30021 , \30022 ,
         \30023 , \30024 , \30025 , \30026 , \30027 , \30028 , \30029 , \30030 , \30031 , \30032 ,
         \30033 , \30034 , \30035 , \30036 , \30037 , \30038 , \30039 , \30040 , \30041 , \30042 ,
         \30043 , \30044 , \30045 , \30046 , \30047 , \30048 , \30049 , \30050 , \30051 , \30052 ,
         \30053 , \30054 , \30055 , \30056 , \30057 , \30058 , \30059 , \30060 , \30061 , \30062 ,
         \30063 , \30064 , \30065 , \30066 , \30067 , \30068 , \30069 , \30070 , \30071 , \30072 ,
         \30073 , \30074 , \30075 , \30076 , \30077 , \30078 , \30079 , \30080 , \30081 , \30082 ,
         \30083 , \30084 , \30085 , \30086 , \30087 , \30088 , \30089 , \30090 , \30091 , \30092 ,
         \30093 , \30094 , \30095 , \30096 , \30097 , \30098 , \30099 , \30100 , \30101 , \30102 ,
         \30103 , \30104 , \30105 , \30106 , \30107 , \30108 , \30109 , \30110 , \30111 , \30112 ,
         \30113 , \30114 , \30115 , \30116 , \30117 , \30118 , \30119 , \30120 , \30121 , \30122 ,
         \30123 , \30124 , \30125 , \30126 , \30127 , \30128 , \30129 , \30130 , \30131 , \30132 ,
         \30133 , \30134 , \30135 , \30136 , \30137 , \30138 , \30139 , \30140 , \30141 , \30142 ,
         \30143 , \30144 , \30145 , \30146 , \30147 , \30148 , \30149 , \30150 , \30151 , \30152 ,
         \30153 , \30154 , \30155 , \30156 , \30157 , \30158 , \30159 , \30160 , \30161 , \30162 ,
         \30163 , \30164 , \30165 , \30166 , \30167 , \30168 , \30169 , \30170 , \30171 , \30172 ,
         \30173 , \30174 , \30175 , \30176 , \30177 , \30178 , \30179 , \30180 , \30181 , \30182 ,
         \30183 , \30184 , \30185 , \30186 , \30187 , \30188 , \30189 , \30190 , \30191 , \30192 ,
         \30193 , \30194 , \30195 , \30196 , \30197 , \30198 , \30199 , \30200 , \30201 , \30202 ,
         \30203 , \30204 , \30205 , \30206 , \30207 , \30208 , \30209 , \30210 , \30211 , \30212 ,
         \30213 , \30214 , \30215 , \30216 , \30217 , \30218 , \30219 , \30220 , \30221 , \30222 ,
         \30223 , \30224 , \30225 , \30226 , \30227 , \30228 , \30229 , \30230 , \30231 , \30232 ,
         \30233 , \30234 , \30235 , \30236 , \30237 , \30238 , \30239 , \30240 , \30241 , \30242 ,
         \30243 , \30244 , \30245 , \30246 , \30247 , \30248 , \30249 , \30250 , \30251 , \30252 ,
         \30253 , \30254 , \30255 , \30256 , \30257 , \30258 , \30259 , \30260 , \30261 , \30262 ,
         \30263 , \30264 , \30265 , \30266 , \30267 , \30268 , \30269 , \30270 , \30271 , \30272 ,
         \30273 , \30274 , \30275 , \30276 , \30277 , \30278 , \30279 , \30280 , \30281 , \30282 ,
         \30283 , \30284 , \30285 , \30286 , \30287 , \30288 , \30289 , \30290 , \30291 , \30292 ,
         \30293 , \30294 , \30295 , \30296 , \30297 , \30298 , \30299 , \30300 , \30301 , \30302 ,
         \30303 , \30304 , \30305 , \30306 , \30307 , \30308 , \30309 , \30310 , \30311 , \30312 ,
         \30313 , \30314 , \30315 , \30316 , \30317 , \30318 , \30319 , \30320 , \30321 , \30322 ,
         \30323 , \30324 , \30325 , \30326 , \30327 , \30328 , \30329 , \30330 , \30331 , \30332 ,
         \30333 , \30334 , \30335 , \30336 , \30337 , \30338 , \30339 , \30340 , \30341 , \30342 ,
         \30343 , \30344 , \30345 , \30346 , \30347 , \30348 , \30349 , \30350 , \30351 , \30352 ,
         \30353 , \30354 , \30355 , \30356 , \30357 , \30358 , \30359 , \30360 , \30361 , \30362 ,
         \30363 , \30364 , \30365 , \30366 , \30367 , \30368 , \30369 , \30370 , \30371 , \30372 ,
         \30373 , \30374 , \30375 , \30376 , \30377 , \30378 , \30379 , \30380 , \30381 , \30382 ,
         \30383 , \30384 , \30385 , \30386 , \30387 , \30388 , \30389 , \30390 , \30391 , \30392 ,
         \30393 , \30394 , \30395 , \30396 , \30397 , \30398 , \30399 , \30400 , \30401 , \30402 ,
         \30403 , \30404 , \30405 , \30406 , \30407 , \30408 , \30409 , \30410 , \30411 , \30412 ,
         \30413 , \30414 , \30415 , \30416 , \30417 , \30418 , \30419 , \30420 , \30421 , \30422 ,
         \30423 , \30424 , \30425 , \30426 , \30427 , \30428 , \30429 , \30430 , \30431 , \30432 ,
         \30433 , \30434 , \30435 , \30436 , \30437 , \30438 , \30439 , \30440 , \30441 , \30442 ,
         \30443 , \30444 , \30445 , \30446 , \30447 , \30448 , \30449 , \30450 , \30451 , \30452 ,
         \30453 , \30454 , \30455 , \30456 , \30457 , \30458 , \30459 , \30460 , \30461 , \30462 ,
         \30463 , \30464 , \30465 , \30466 , \30467 , \30468 , \30469 , \30470 , \30471 , \30472 ,
         \30473 , \30474 , \30475 , \30476 , \30477 , \30478 , \30479 , \30480 , \30481 , \30482 ,
         \30483 , \30484 , \30485 , \30486 , \30487 , \30488 , \30489 , \30490 , \30491 , \30492 ,
         \30493 , \30494 , \30495 , \30496 , \30497 , \30498 , \30499 , \30500 , \30501 , \30502 ,
         \30503 , \30504 , \30505 , \30506 , \30507 , \30508 , \30509 , \30510 , \30511 , \30512 ,
         \30513 , \30514 , \30515 , \30516 , \30517 , \30518 , \30519 , \30520 , \30521 , \30522 ,
         \30523 , \30524 , \30525 , \30526 , \30527 , \30528 , \30529 , \30530 , \30531 , \30532 ,
         \30533 , \30534 , \30535 , \30536 , \30537 , \30538 , \30539 , \30540 , \30541 , \30542 ,
         \30543 , \30544 , \30545 , \30546 , \30547 , \30548 , \30549 , \30550 , \30551 , \30552 ,
         \30553 , \30554 , \30555 , \30556 , \30557 , \30558 , \30559 , \30560 , \30561 , \30562 ,
         \30563 , \30564 , \30565 , \30566 , \30567 , \30568 , \30569 , \30570 , \30571 , \30572 ,
         \30573 , \30574 , \30575 , \30576 , \30577 , \30578 , \30579 , \30580 , \30581 , \30582 ,
         \30583 , \30584 , \30585 , \30586 , \30587 , \30588 , \30589 , \30590 , \30591 , \30592 ,
         \30593 , \30594 , \30595 , \30596 , \30597 , \30598 , \30599 , \30600 , \30601 , \30602 ,
         \30603 , \30604 , \30605 , \30606 , \30607 , \30608 , \30609 , \30610 , \30611 , \30612 ,
         \30613 , \30614 , \30615 , \30616 , \30617 , \30618 , \30619 , \30620 , \30621 , \30622 ,
         \30623 , \30624 , \30625 , \30626 , \30627 , \30628 , \30629 , \30630 , \30631 , \30632 ,
         \30633 , \30634 , \30635 , \30636 , \30637 , \30638 , \30639 , \30640 , \30641 , \30642 ,
         \30643 , \30644 , \30645 , \30646 , \30647 , \30648 , \30649 , \30650 , \30651 , \30652 ,
         \30653 , \30654 , \30655 , \30656 , \30657 , \30658 , \30659 , \30660 , \30661 , \30662 ,
         \30663 , \30664 , \30665 , \30666 , \30667 , \30668 , \30669 , \30670 , \30671 , \30672 ,
         \30673 , \30674 , \30675 , \30676 , \30677 , \30678 , \30679 , \30680 , \30681 , \30682 ,
         \30683 , \30684 , \30685 , \30686 , \30687 , \30688 , \30689 , \30690 , \30691 , \30692 ,
         \30693 , \30694 , \30695 , \30696 , \30697 , \30698 , \30699 , \30700 , \30701 , \30702 ,
         \30703 , \30704 , \30705 , \30706 , \30707 , \30708 , \30709 , \30710 , \30711 , \30712 ,
         \30713 , \30714 , \30715 , \30716 , \30717 , \30718 , \30719 , \30720 , \30721 , \30722 ,
         \30723 , \30724 , \30725 , \30726 , \30727 , \30728 , \30729 , \30730 , \30731 , \30732 ,
         \30733 , \30734 , \30735 , \30736 , \30737 , \30738 , \30739 , \30740 , \30741 , \30742 ,
         \30743 , \30744 , \30745 , \30746 , \30747 , \30748 , \30749 , \30750 , \30751 , \30752 ,
         \30753 , \30754 , \30755 , \30756 , \30757 , \30758 , \30759 , \30760 , \30761 , \30762 ,
         \30763 , \30764 , \30765 , \30766 , \30767 , \30768 , \30769 , \30770 , \30771 , \30772 ,
         \30773 , \30774 , \30775 , \30776 , \30777 , \30778 , \30779 , \30780 , \30781 , \30782 ,
         \30783 , \30784 , \30785 , \30786 , \30787 , \30788 , \30789 , \30790 , \30791 , \30792 ,
         \30793 , \30794 , \30795 , \30796 , \30797 , \30798 , \30799 , \30800 , \30801 , \30802 ,
         \30803 , \30804 , \30805 , \30806 , \30807 , \30808 , \30809 , \30810 , \30811 , \30812 ,
         \30813 , \30814 , \30815 , \30816 , \30817 , \30818 , \30819 , \30820 , \30821 , \30822 ,
         \30823 , \30824 , \30825 , \30826 , \30827 , \30828 , \30829 , \30830 , \30831 , \30832 ,
         \30833 , \30834 , \30835 , \30836 , \30837 , \30838 , \30839 , \30840 , \30841 , \30842 ,
         \30843 , \30844 , \30845 , \30846 , \30847 , \30848 , \30849 , \30850 , \30851 , \30852 ,
         \30853 , \30854 , \30855 , \30856 , \30857 , \30858 , \30859 , \30860 , \30861 , \30862 ,
         \30863 , \30864 , \30865 , \30866 , \30867 , \30868 , \30869 , \30870 , \30871 , \30872 ,
         \30873 , \30874 , \30875 , \30876 , \30877 , \30878 , \30879 , \30880 , \30881 , \30882 ,
         \30883 , \30884 , \30885 , \30886 , \30887 , \30888 , \30889 , \30890 , \30891 , \30892 ,
         \30893 , \30894 , \30895 , \30896 , \30897 , \30898 , \30899 , \30900 , \30901 , \30902 ,
         \30903 , \30904 , \30905 , \30906 , \30907 , \30908 , \30909 , \30910 , \30911 , \30912 ,
         \30913 , \30914 , \30915 , \30916 , \30917 , \30918 , \30919 , \30920 , \30921 , \30922 ,
         \30923 , \30924 , \30925 , \30926 , \30927 , \30928 , \30929 , \30930 , \30931 , \30932 ,
         \30933 , \30934 , \30935 , \30936 , \30937 , \30938 , \30939 , \30940 , \30941 , \30942 ,
         \30943 , \30944 , \30945 , \30946 , \30947 , \30948 , \30949 , \30950 , \30951 , \30952 ,
         \30953 , \30954 , \30955 , \30956 , \30957 , \30958 , \30959 , \30960 , \30961 , \30962 ,
         \30963 , \30964 , \30965 , \30966 , \30967 , \30968 , \30969 , \30970 , \30971 , \30972 ,
         \30973 , \30974 , \30975 , \30976 , \30977 , \30978 , \30979 , \30980 , \30981 , \30982 ,
         \30983 , \30984 , \30985 , \30986 , \30987 , \30988 , \30989 , \30990 , \30991 , \30992 ,
         \30993 , \30994 , \30995 , \30996 , \30997 , \30998 , \30999 , \31000 , \31001 , \31002 ,
         \31003 , \31004 , \31005 , \31006 , \31007 , \31008 , \31009 , \31010 , \31011 , \31012 ,
         \31013 , \31014 , \31015 , \31016 , \31017 , \31018 , \31019 , \31020 , \31021 , \31022 ,
         \31023 , \31024 , \31025 , \31026 , \31027 , \31028 , \31029 , \31030 , \31031 , \31032 ,
         \31033 , \31034 , \31035 , \31036 , \31037 , \31038 , \31039 , \31040 , \31041 , \31042 ,
         \31043 , \31044 , \31045 , \31046 , \31047 , \31048 , \31049 , \31050 , \31051 , \31052 ,
         \31053 , \31054 , \31055 , \31056 , \31057 , \31058 , \31059 , \31060 , \31061 , \31062 ,
         \31063 , \31064 , \31065 , \31066 , \31067 , \31068 , \31069 , \31070 , \31071 , \31072 ,
         \31073 , \31074 , \31075 , \31076 , \31077 , \31078 , \31079 , \31080 , \31081 , \31082 ,
         \31083 , \31084 , \31085 , \31086 , \31087 , \31088 , \31089 , \31090 , \31091 , \31092 ,
         \31093 , \31094 , \31095 , \31096 , \31097 , \31098 , \31099 , \31100 , \31101 , \31102 ,
         \31103 , \31104 , \31105 , \31106 , \31107 , \31108 , \31109 , \31110 , \31111 , \31112 ,
         \31113 , \31114 , \31115 , \31116 , \31117 , \31118 , \31119 , \31120 , \31121 , \31122 ,
         \31123 , \31124 , \31125 , \31126 , \31127 , \31128 , \31129 , \31130 , \31131 , \31132 ,
         \31133 , \31134 , \31135 , \31136 , \31137 , \31138 , \31139 , \31140 , \31141 , \31142 ,
         \31143 , \31144 , \31145 , \31146 , \31147 , \31148 , \31149 , \31150 , \31151 , \31152 ,
         \31153 , \31154 , \31155 , \31156 , \31157 , \31158 , \31159 , \31160 , \31161 , \31162 ,
         \31163 , \31164 , \31165 , \31166 , \31167 , \31168 , \31169 , \31170 , \31171 , \31172 ,
         \31173 , \31174 , \31175 , \31176 , \31177 , \31178 , \31179 , \31180 , \31181 , \31182 ,
         \31183 , \31184 , \31185 , \31186 , \31187 , \31188 , \31189 , \31190 , \31191 , \31192 ,
         \31193 , \31194 , \31195 , \31196 , \31197 , \31198 , \31199 , \31200 , \31201 , \31202 ,
         \31203 , \31204 , \31205 , \31206 , \31207 , \31208 , \31209 , \31210 , \31211 , \31212 ,
         \31213 , \31214 , \31215 , \31216 , \31217 , \31218 , \31219 , \31220 , \31221 , \31222 ,
         \31223 , \31224 , \31225 , \31226 , \31227 , \31228 , \31229 , \31230 , \31231 , \31232 ,
         \31233 , \31234 , \31235 , \31236 , \31237 , \31238 , \31239 , \31240 , \31241 , \31242 ,
         \31243 , \31244 , \31245 , \31246 , \31247 , \31248 , \31249 , \31250 , \31251 , \31252 ,
         \31253 , \31254 , \31255 , \31256 , \31257 , \31258 , \31259 , \31260 , \31261 , \31262 ,
         \31263 , \31264 , \31265 , \31266 , \31267 , \31268 , \31269 , \31270 , \31271 , \31272 ,
         \31273 , \31274 , \31275 , \31276 , \31277 , \31278 , \31279 , \31280 , \31281 , \31282 ,
         \31283 , \31284 , \31285 , \31286 , \31287 , \31288 , \31289 , \31290 , \31291 , \31292 ,
         \31293 , \31294 , \31295 , \31296 , \31297 , \31298 , \31299 , \31300 , \31301 , \31302 ,
         \31303 , \31304 , \31305 , \31306 , \31307 , \31308 , \31309 , \31310 , \31311 , \31312 ,
         \31313 , \31314 , \31315 , \31316 , \31317 , \31318 , \31319 , \31320 , \31321 , \31322 ,
         \31323 , \31324 , \31325 , \31326 , \31327 , \31328 , \31329 , \31330 , \31331 , \31332 ,
         \31333 , \31334 , \31335 , \31336 , \31337 , \31338 , \31339 , \31340 , \31341 , \31342 ,
         \31343 , \31344 , \31345 , \31346 , \31347 , \31348 , \31349 , \31350 , \31351 , \31352 ,
         \31353 , \31354 , \31355 , \31356 , \31357 , \31358 , \31359 , \31360 , \31361 , \31362 ,
         \31363 , \31364 , \31365 , \31366 , \31367 , \31368 , \31369 , \31370 , \31371 , \31372 ,
         \31373 , \31374 , \31375 , \31376 , \31377 , \31378 , \31379 , \31380 , \31381 , \31382 ,
         \31383 , \31384 , \31385 , \31386 , \31387 , \31388 , \31389 , \31390 , \31391 , \31392 ,
         \31393 , \31394 , \31395 , \31396 , \31397 , \31398 , \31399 , \31400 , \31401 , \31402 ,
         \31403 , \31404 , \31405 , \31406 , \31407 , \31408 , \31409 , \31410 , \31411 , \31412 ,
         \31413 , \31414 , \31415 , \31416 , \31417 , \31418 , \31419 , \31420 , \31421 , \31422 ,
         \31423 , \31424 , \31425 , \31426 , \31427 , \31428 , \31429 , \31430 , \31431 , \31432 ,
         \31433 , \31434 , \31435 , \31436 , \31437 , \31438 , \31439 , \31440 , \31441 , \31442 ,
         \31443 , \31444 , \31445 , \31446 , \31447 , \31448 , \31449 , \31450 , \31451 , \31452 ,
         \31453 , \31454 , \31455 , \31456 , \31457 , \31458 , \31459 , \31460 , \31461 , \31462 ,
         \31463 , \31464 , \31465 , \31466 , \31467 , \31468 , \31469 , \31470 , \31471 , \31472 ,
         \31473 , \31474 , \31475 , \31476 , \31477 , \31478 , \31479 , \31480 , \31481 , \31482 ,
         \31483 , \31484 , \31485 , \31486 , \31487 , \31488 , \31489 , \31490 , \31491 , \31492 ,
         \31493 , \31494 , \31495 , \31496 , \31497 , \31498 , \31499 , \31500 , \31501 , \31502 ,
         \31503 , \31504 , \31505 , \31506 , \31507 , \31508 , \31509 , \31510 , \31511 , \31512 ,
         \31513 , \31514 , \31515 , \31516 , \31517 , \31518 , \31519 , \31520 , \31521 , \31522 ,
         \31523 , \31524 , \31525 , \31526 , \31527 , \31528 , \31529 , \31530 , \31531 , \31532 ,
         \31533 , \31534 , \31535 , \31536 , \31537 , \31538 , \31539 , \31540 , \31541 , \31542 ,
         \31543 , \31544 , \31545 , \31546 , \31547 , \31548 , \31549 , \31550 , \31551 , \31552 ,
         \31553 , \31554 , \31555 , \31556 , \31557 , \31558 , \31559 , \31560 , \31561 , \31562 ,
         \31563 , \31564 , \31565 , \31566 , \31567 , \31568 , \31569 , \31570 , \31571 , \31572 ,
         \31573 , \31574 , \31575 , \31576 , \31577 , \31578 , \31579 , \31580 , \31581 , \31582 ,
         \31583 , \31584 , \31585 , \31586 , \31587 , \31588 , \31589 , \31590 , \31591 , \31592 ,
         \31593 , \31594 , \31595 , \31596 , \31597 , \31598 , \31599 , \31600 , \31601 , \31602 ,
         \31603 , \31604 , \31605 , \31606 , \31607 , \31608 , \31609 , \31610 , \31611 , \31612 ,
         \31613 , \31614 , \31615 , \31616 , \31617 , \31618 , \31619 , \31620 , \31621 , \31622 ,
         \31623 , \31624 , \31625 , \31626 , \31627 , \31628 , \31629 , \31630 , \31631 , \31632 ,
         \31633 , \31634 , \31635 , \31636 , \31637 , \31638 , \31639 , \31640 , \31641 , \31642 ,
         \31643 , \31644 , \31645 , \31646 , \31647 , \31648 , \31649 , \31650 , \31651 , \31652 ,
         \31653 , \31654 , \31655 , \31656 , \31657 , \31658 , \31659 , \31660 , \31661 , \31662 ,
         \31663 , \31664 , \31665 , \31666 , \31667 , \31668 , \31669 , \31670 , \31671 , \31672 ,
         \31673 , \31674 , \31675 , \31676 , \31677 , \31678 , \31679 , \31680 , \31681 , \31682 ,
         \31683 , \31684 , \31685 , \31686 , \31687 , \31688 , \31689 , \31690 , \31691 , \31692 ,
         \31693 , \31694 , \31695 , \31696 , \31697 , \31698 , \31699 , \31700 , \31701 , \31702 ,
         \31703 , \31704 , \31705 , \31706 , \31707 , \31708 , \31709 , \31710 , \31711 , \31712 ,
         \31713 , \31714 , \31715 , \31716 , \31717 , \31718 , \31719 , \31720 , \31721 , \31722 ,
         \31723 , \31724 , \31725 , \31726 , \31727 , \31728 , \31729 , \31730 , \31731 , \31732 ,
         \31733 , \31734 , \31735 , \31736 , \31737 , \31738 , \31739 , \31740 , \31741 , \31742 ,
         \31743 , \31744 , \31745 , \31746 , \31747 , \31748 , \31749 , \31750 , \31751 , \31752 ,
         \31753 , \31754 , \31755 , \31756 , \31757 , \31758 , \31759 , \31760 , \31761 , \31762 ,
         \31763 , \31764 , \31765 , \31766 , \31767 , \31768 , \31769 , \31770 , \31771 , \31772 ,
         \31773 , \31774 , \31775 , \31776 , \31777 , \31778 , \31779 , \31780 , \31781 , \31782 ,
         \31783 , \31784 , \31785 , \31786 , \31787 , \31788 , \31789 , \31790 , \31791 , \31792 ,
         \31793 , \31794 , \31795 , \31796 , \31797 , \31798 , \31799 , \31800 , \31801 , \31802 ,
         \31803 , \31804 , \31805 , \31806 , \31807 , \31808 , \31809 , \31810 , \31811 , \31812 ,
         \31813 , \31814 , \31815 , \31816 , \31817 , \31818 , \31819 , \31820 , \31821 , \31822 ,
         \31823 , \31824 , \31825 , \31826 , \31827 , \31828 , \31829 , \31830 , \31831 , \31832 ,
         \31833 , \31834 , \31835 , \31836 , \31837 , \31838 , \31839 , \31840 , \31841 , \31842 ,
         \31843 , \31844 , \31845 , \31846 , \31847 , \31848 , \31849 , \31850 , \31851 , \31852 ,
         \31853 , \31854 , \31855 , \31856 , \31857 , \31858 , \31859 , \31860 , \31861 , \31862 ,
         \31863 , \31864 , \31865 , \31866 , \31867 , \31868 , \31869 , \31870 , \31871 , \31872 ,
         \31873 , \31874 , \31875 , \31876 , \31877 , \31878 , \31879 , \31880 , \31881 , \31882 ,
         \31883 , \31884 , \31885 , \31886 , \31887 , \31888 , \31889 , \31890 , \31891 , \31892 ,
         \31893 , \31894 , \31895 , \31896 , \31897 , \31898 , \31899 , \31900 , \31901 , \31902 ,
         \31903 , \31904 , \31905 , \31906 , \31907 , \31908 , \31909 , \31910 , \31911 , \31912 ,
         \31913 , \31914 , \31915 , \31916 , \31917 , \31918 , \31919 , \31920 , \31921 , \31922 ,
         \31923 , \31924 , \31925 , \31926 , \31927 , \31928 , \31929 , \31930 , \31931 , \31932 ,
         \31933 , \31934 , \31935 , \31936 , \31937 , \31938 , \31939 , \31940 , \31941 , \31942 ,
         \31943 , \31944 , \31945 , \31946 , \31947 , \31948 , \31949 , \31950 , \31951 , \31952 ,
         \31953 , \31954 , \31955 , \31956 , \31957 , \31958 , \31959 , \31960 , \31961 , \31962 ,
         \31963 , \31964 , \31965 , \31966 , \31967 , \31968 , \31969 , \31970 , \31971 , \31972 ,
         \31973 , \31974 , \31975 , \31976 , \31977 , \31978 , \31979 , \31980 , \31981 , \31982 ,
         \31983 , \31984 , \31985 , \31986 , \31987 , \31988 , \31989 , \31990 , \31991 , \31992 ,
         \31993 , \31994 , \31995 , \31996 , \31997 , \31998 , \31999 , \32000 , \32001 , \32002 ,
         \32003 , \32004 , \32005 , \32006 , \32007 , \32008 , \32009 , \32010 , \32011 , \32012 ,
         \32013 , \32014 , \32015 , \32016 , \32017 , \32018 , \32019 , \32020 , \32021 , \32022 ,
         \32023 , \32024 , \32025 , \32026 , \32027 , \32028 , \32029 , \32030 , \32031 , \32032 ,
         \32033 , \32034 , \32035 , \32036 , \32037 , \32038 , \32039 , \32040 , \32041 , \32042 ,
         \32043 , \32044 , \32045 , \32046 , \32047 , \32048 , \32049 , \32050 , \32051 , \32052 ,
         \32053 , \32054 , \32055 , \32056 , \32057 , \32058 , \32059 , \32060 , \32061 , \32062 ,
         \32063 , \32064 , \32065 , \32066 , \32067 , \32068 , \32069 , \32070 , \32071 , \32072 ,
         \32073 , \32074 , \32075 , \32076 , \32077 , \32078 , \32079 , \32080 , \32081 , \32082 ,
         \32083 , \32084 , \32085 , \32086 , \32087 , \32088 , \32089 , \32090 , \32091 , \32092 ,
         \32093 , \32094 , \32095 , \32096 , \32097 , \32098 , \32099 , \32100 , \32101 , \32102 ,
         \32103 , \32104 , \32105 , \32106 , \32107 , \32108 , \32109 , \32110 , \32111 , \32112 ,
         \32113 , \32114 , \32115 , \32116 , \32117 , \32118 , \32119 , \32120 , \32121 , \32122 ,
         \32123 , \32124 , \32125 , \32126 , \32127 , \32128 , \32129 , \32130 , \32131 , \32132 ,
         \32133 , \32134 , \32135 , \32136 , \32137 , \32138 , \32139 , \32140 , \32141 , \32142 ,
         \32143 , \32144 , \32145 , \32146 , \32147 , \32148 , \32149 , \32150 , \32151 , \32152 ,
         \32153 , \32154 , \32155 , \32156 , \32157 , \32158 , \32159 , \32160 , \32161 , \32162 ,
         \32163 , \32164 , \32165 , \32166 , \32167 , \32168 , \32169 , \32170 , \32171 , \32172 ,
         \32173 , \32174 , \32175 , \32176 , \32177 , \32178 , \32179 , \32180 , \32181 , \32182 ,
         \32183 , \32184 , \32185 , \32186 , \32187 , \32188 , \32189 , \32190 , \32191 , \32192 ,
         \32193 , \32194 , \32195 , \32196 , \32197 , \32198 , \32199 , \32200 , \32201 , \32202 ,
         \32203 , \32204 , \32205 , \32206 , \32207 , \32208 , \32209 , \32210 , \32211 , \32212 ,
         \32213 , \32214 , \32215 , \32216 , \32217 , \32218 , \32219 , \32220 , \32221 , \32222 ,
         \32223 , \32224 , \32225 , \32226 , \32227 , \32228 , \32229 , \32230 , \32231 , \32232 ,
         \32233 , \32234 , \32235 , \32236 , \32237 , \32238 , \32239 , \32240 , \32241 , \32242 ,
         \32243 , \32244 , \32245 , \32246 , \32247 , \32248 , \32249 , \32250 , \32251 , \32252 ,
         \32253 , \32254 , \32255 , \32256 , \32257 , \32258 , \32259 , \32260 , \32261 , \32262 ,
         \32263 , \32264 , \32265 , \32266 , \32267 , \32268 , \32269 , \32270 , \32271 , \32272 ,
         \32273 , \32274 , \32275 , \32276 , \32277 , \32278 , \32279 , \32280 , \32281 , \32282 ,
         \32283 , \32284 , \32285 , \32286 , \32287 , \32288 , \32289 , \32290 , \32291 , \32292 ,
         \32293 , \32294 , \32295 , \32296 , \32297 , \32298 , \32299 , \32300 , \32301 , \32302 ,
         \32303 , \32304 , \32305 , \32306 , \32307 , \32308 , \32309 , \32310 , \32311 , \32312 ,
         \32313 , \32314 , \32315 , \32316 , \32317 , \32318 , \32319 , \32320 , \32321 , \32322 ,
         \32323 , \32324 , \32325 , \32326 , \32327 , \32328 , \32329 , \32330 , \32331 , \32332 ,
         \32333 , \32334 , \32335 , \32336 , \32337 , \32338 , \32339 , \32340 , \32341 , \32342 ,
         \32343 , \32344 , \32345 , \32346 , \32347 , \32348 , \32349 , \32350 , \32351 , \32352 ,
         \32353 , \32354 , \32355 , \32356 , \32357 , \32358 , \32359 , \32360 , \32361 , \32362 ,
         \32363 , \32364 , \32365 , \32366 , \32367 , \32368 , \32369 , \32370 , \32371 , \32372 ,
         \32373 , \32374 , \32375 , \32376 , \32377 , \32378 , \32379 , \32380 , \32381 , \32382 ,
         \32383 , \32384 , \32385 , \32386 , \32387 , \32388 , \32389 , \32390 , \32391 , \32392 ,
         \32393 , \32394 , \32395 , \32396 , \32397 , \32398 , \32399 , \32400 , \32401 , \32402 ,
         \32403 , \32404 , \32405 , \32406 , \32407 , \32408 , \32409 , \32410 , \32411 , \32412 ,
         \32413 , \32414 , \32415 , \32416 , \32417 , \32418 , \32419 , \32420 , \32421 , \32422 ,
         \32423 , \32424 , \32425 , \32426 , \32427 , \32428 , \32429 , \32430 , \32431 , \32432 ,
         \32433 , \32434 , \32435 , \32436 , \32437 , \32438 , \32439 , \32440 , \32441 , \32442 ,
         \32443 , \32444 , \32445 , \32446 , \32447 , \32448 , \32449 , \32450 , \32451 , \32452 ,
         \32453 , \32454 , \32455 , \32456 , \32457 , \32458 , \32459 , \32460 , \32461 , \32462 ,
         \32463 , \32464 , \32465 , \32466 , \32467 , \32468 , \32469 , \32470 , \32471 , \32472 ,
         \32473 , \32474 , \32475 , \32476 , \32477 , \32478 , \32479 , \32480 , \32481 , \32482 ,
         \32483 , \32484 , \32485 , \32486 , \32487 , \32488 , \32489 , \32490 , \32491 , \32492 ,
         \32493 , \32494 , \32495 , \32496 , \32497 , \32498 , \32499 , \32500 , \32501 , \32502 ,
         \32503 , \32504 , \32505 , \32506 , \32507 , \32508 , \32509 , \32510 , \32511 , \32512 ,
         \32513 , \32514 , \32515 , \32516 , \32517 , \32518 , \32519 , \32520 , \32521 , \32522 ,
         \32523 , \32524 , \32525 , \32526 , \32527 , \32528 , \32529 , \32530 , \32531 , \32532 ,
         \32533 , \32534 , \32535 , \32536 , \32537 , \32538 , \32539 , \32540 , \32541 , \32542 ,
         \32543 , \32544 , \32545 , \32546 , \32547 , \32548 , \32549 , \32550 , \32551 , \32552 ,
         \32553 , \32554 , \32555 , \32556 , \32557 , \32558 , \32559 , \32560 , \32561 , \32562 ,
         \32563 , \32564 , \32565 , \32566 , \32567 , \32568 , \32569 , \32570 , \32571 , \32572 ,
         \32573 , \32574 , \32575 , \32576 , \32577 , \32578 , \32579 , \32580 , \32581 , \32582 ,
         \32583 , \32584 , \32585 , \32586 , \32587 , \32588 , \32589 , \32590 , \32591 , \32592 ,
         \32593 , \32594 , \32595 , \32596 , \32597 , \32598 , \32599 , \32600 , \32601 , \32602 ,
         \32603 , \32604 , \32605 , \32606 , \32607 , \32608 , \32609 , \32610 , \32611 , \32612 ,
         \32613 , \32614 , \32615 , \32616 , \32617 , \32618 , \32619 , \32620 , \32621 , \32622 ,
         \32623 , \32624 , \32625 , \32626 , \32627 , \32628 , \32629 , \32630 , \32631 , \32632 ,
         \32633 , \32634 , \32635 , \32636 , \32637 , \32638 , \32639 , \32640 , \32641 , \32642 ,
         \32643 , \32644 , \32645 , \32646 , \32647 , \32648 , \32649 , \32650 , \32651 , \32652 ,
         \32653 , \32654 , \32655 , \32656 , \32657 , \32658 , \32659 , \32660 , \32661 , \32662 ,
         \32663 , \32664 , \32665 , \32666 , \32667 , \32668 , \32669 , \32670 , \32671 , \32672 ,
         \32673 , \32674 , \32675 , \32676 , \32677 , \32678 , \32679 , \32680 , \32681 , \32682 ,
         \32683 , \32684 , \32685 , \32686 , \32687 , \32688 , \32689 , \32690 , \32691 , \32692 ,
         \32693 , \32694 , \32695 , \32696 , \32697 , \32698 , \32699 , \32700 , \32701 , \32702 ,
         \32703 , \32704 , \32705 , \32706 , \32707 , \32708 , \32709 , \32710 , \32711 , \32712 ,
         \32713 , \32714 , \32715 , \32716 , \32717 , \32718 , \32719 , \32720 , \32721 , \32722 ,
         \32723 , \32724 , \32725 , \32726 , \32727 , \32728 , \32729 , \32730 , \32731 , \32732 ,
         \32733 , \32734 , \32735 , \32736 , \32737 , \32738 , \32739 , \32740 , \32741 , \32742 ,
         \32743 , \32744 , \32745 , \32746 , \32747 , \32748 , \32749 , \32750 , \32751 , \32752 ,
         \32753 , \32754 , \32755 , \32756 , \32757 , \32758 , \32759 , \32760 , \32761 , \32762 ,
         \32763 , \32764 , \32765 , \32766 , \32767 , \32768 , \32769 , \32770 , \32771 , \32772 ,
         \32773 , \32774 , \32775 , \32776 , \32777 , \32778 , \32779 , \32780 , \32781 , \32782 ,
         \32783 , \32784 , \32785 , \32786 , \32787 , \32788 , \32789 , \32790 , \32791 , \32792 ,
         \32793 , \32794 , \32795 , \32796 , \32797 , \32798 , \32799 , \32800 , \32801 , \32802 ,
         \32803 , \32804 , \32805 , \32806 , \32807 , \32808 , \32809 , \32810 , \32811 , \32812 ,
         \32813 , \32814 , \32815 , \32816 , \32817 , \32818 , \32819 , \32820 , \32821 , \32822 ,
         \32823 , \32824 , \32825 , \32826 , \32827 , \32828 , \32829 , \32830 , \32831 , \32832 ,
         \32833 , \32834 , \32835 , \32836 , \32837 , \32838 , \32839 , \32840 , \32841 , \32842 ,
         \32843 , \32844 , \32845 , \32846 , \32847 , \32848 , \32849 , \32850 , \32851 , \32852 ,
         \32853 , \32854 , \32855 , \32856 , \32857 , \32858 , \32859 , \32860 , \32861 , \32862 ,
         \32863 , \32864 , \32865 , \32866 , \32867 , \32868 , \32869 , \32870 , \32871 , \32872 ,
         \32873 , \32874 , \32875 , \32876 , \32877 , \32878 , \32879 , \32880 , \32881 , \32882 ,
         \32883 , \32884 , \32885 , \32886 , \32887 , \32888 , \32889 , \32890 , \32891 , \32892 ,
         \32893 , \32894 , \32895 , \32896 , \32897 , \32898 , \32899 , \32900 , \32901 , \32902 ,
         \32903 , \32904 , \32905 , \32906 , \32907 , \32908 , \32909 , \32910 , \32911 , \32912 ,
         \32913 , \32914 , \32915 , \32916 , \32917 , \32918 , \32919 , \32920 , \32921 , \32922 ,
         \32923 , \32924 , \32925 , \32926 , \32927 , \32928 , \32929 , \32930 , \32931 , \32932 ,
         \32933 , \32934 , \32935 , \32936 , \32937 , \32938 , \32939 , \32940 , \32941 , \32942 ,
         \32943 , \32944 , \32945 , \32946 , \32947 , \32948 , \32949 , \32950 , \32951 , \32952 ,
         \32953 , \32954 , \32955 , \32956 , \32957 , \32958 , \32959 , \32960 , \32961 , \32962 ,
         \32963 , \32964 , \32965 , \32966 , \32967 , \32968 , \32969 , \32970 , \32971 , \32972 ,
         \32973 , \32974 , \32975 , \32976 , \32977 , \32978 , \32979 , \32980 , \32981 , \32982 ,
         \32983 , \32984 , \32985 , \32986 , \32987 , \32988 , \32989 , \32990 , \32991 , \32992 ,
         \32993 , \32994 , \32995 , \32996 , \32997 , \32998 , \32999 , \33000 , \33001 , \33002 ,
         \33003 , \33004 , \33005 , \33006 , \33007 , \33008 , \33009 , \33010 , \33011 , \33012 ,
         \33013 , \33014 , \33015 , \33016 , \33017 , \33018 , \33019 , \33020 , \33021 , \33022 ,
         \33023 , \33024 , \33025 , \33026 , \33027 , \33028 , \33029 , \33030 , \33031 , \33032 ,
         \33033 , \33034 , \33035 , \33036 , \33037 , \33038 , \33039 , \33040 , \33041 , \33042 ,
         \33043 , \33044 , \33045 , \33046 , \33047 , \33048 , \33049 , \33050 , \33051 , \33052 ,
         \33053 , \33054 , \33055 , \33056 , \33057 , \33058 , \33059 , \33060 , \33061 , \33062 ,
         \33063 , \33064 , \33065 , \33066 , \33067 , \33068 , \33069 , \33070 , \33071 , \33072 ,
         \33073 , \33074 , \33075 , \33076 , \33077 , \33078 , \33079 , \33080 , \33081 , \33082 ,
         \33083 , \33084 , \33085 , \33086 , \33087 , \33088 , \33089 , \33090 , \33091 , \33092 ,
         \33093 , \33094 , \33095 , \33096 , \33097 , \33098 , \33099 , \33100 , \33101 , \33102 ,
         \33103 , \33104 , \33105 , \33106 , \33107 , \33108 , \33109 , \33110 , \33111 , \33112 ,
         \33113 , \33114 , \33115 , \33116 , \33117 , \33118 , \33119 , \33120 , \33121 , \33122 ,
         \33123 , \33124 , \33125 , \33126 , \33127 , \33128 , \33129 , \33130 , \33131 , \33132 ,
         \33133 , \33134 , \33135 , \33136 , \33137 , \33138 , \33139 , \33140 , \33141 , \33142 ,
         \33143 , \33144 , \33145 , \33146 , \33147 , \33148 , \33149 , \33150 , \33151 , \33152 ,
         \33153 , \33154 , \33155 , \33156 , \33157 , \33158 , \33159 , \33160 , \33161 , \33162 ,
         \33163 , \33164 , \33165 , \33166 , \33167 , \33168 , \33169 , \33170 , \33171 , \33172 ,
         \33173 , \33174 , \33175 , \33176 , \33177 , \33178 , \33179 , \33180 , \33181 , \33182 ,
         \33183 , \33184 , \33185 , \33186 , \33187 , \33188 , \33189 , \33190 , \33191 , \33192 ,
         \33193 , \33194 , \33195 , \33196 , \33197 , \33198 , \33199 , \33200 , \33201 , \33202 ,
         \33203 , \33204 , \33205 , \33206 , \33207 , \33208 , \33209 , \33210 , \33211 , \33212 ,
         \33213 , \33214 , \33215 , \33216 , \33217 , \33218 , \33219 , \33220 , \33221 , \33222 ,
         \33223 , \33224 , \33225 , \33226 , \33227 , \33228 , \33229 , \33230 , \33231 , \33232 ,
         \33233 , \33234 , \33235 , \33236 , \33237 , \33238 , \33239 , \33240 , \33241 , \33242 ,
         \33243 , \33244 , \33245 , \33246 , \33247 , \33248 , \33249 , \33250 , \33251 , \33252 ,
         \33253 , \33254 , \33255 , \33256 , \33257 , \33258 , \33259 , \33260 , \33261 , \33262 ,
         \33263 , \33264 , \33265 , \33266 , \33267 , \33268 , \33269 , \33270 , \33271 , \33272 ,
         \33273 , \33274 , \33275 , \33276 , \33277 , \33278 , \33279 , \33280 , \33281 , \33282 ,
         \33283 , \33284 , \33285 , \33286 , \33287 , \33288 , \33289 , \33290 , \33291 , \33292 ,
         \33293 , \33294 , \33295 , \33296 , \33297 , \33298 , \33299 , \33300 , \33301 , \33302 ,
         \33303 , \33304 , \33305 , \33306 , \33307 , \33308 , \33309 , \33310 , \33311 , \33312 ,
         \33313 , \33314 , \33315 , \33316 , \33317 , \33318 , \33319 , \33320 , \33321 , \33322 ,
         \33323 , \33324 , \33325 , \33326 , \33327 , \33328 , \33329 , \33330 , \33331 , \33332 ,
         \33333 , \33334 , \33335 , \33336 , \33337 , \33338 , \33339 , \33340 , \33341 , \33342 ,
         \33343 , \33344 , \33345 , \33346 , \33347 , \33348 , \33349 , \33350 , \33351 , \33352 ,
         \33353 , \33354 , \33355 , \33356 , \33357 , \33358 , \33359 , \33360 , \33361 , \33362 ,
         \33363 , \33364 , \33365 , \33366 , \33367 , \33368 , \33369 , \33370 , \33371 , \33372 ,
         \33373 , \33374 , \33375 , \33376 , \33377 , \33378 , \33379 , \33380 , \33381 , \33382 ,
         \33383 , \33384 , \33385 , \33386 , \33387 , \33388 , \33389 , \33390 , \33391 , \33392 ,
         \33393 , \33394 , \33395 , \33396 , \33397 , \33398 , \33399 , \33400 , \33401 , \33402 ,
         \33403 , \33404 , \33405 , \33406 , \33407 , \33408 , \33409 , \33410 , \33411 , \33412 ,
         \33413 , \33414 , \33415 , \33416 , \33417 , \33418 , \33419 , \33420 , \33421 , \33422 ,
         \33423 , \33424 , \33425 , \33426 , \33427 , \33428 , \33429 , \33430 , \33431 , \33432 ,
         \33433 , \33434 , \33435 , \33436 , \33437 , \33438 , \33439 , \33440 , \33441 , \33442 ,
         \33443 , \33444 , \33445 , \33446 , \33447 , \33448 , \33449 , \33450 , \33451 , \33452 ,
         \33453 , \33454 , \33455 , \33456 , \33457 , \33458 , \33459 , \33460 , \33461 , \33462 ,
         \33463 , \33464 , \33465 , \33466 , \33467 , \33468 , \33469 , \33470 , \33471 , \33472 ,
         \33473 , \33474 , \33475 , \33476 , \33477 , \33478 , \33479 , \33480 , \33481 , \33482 ,
         \33483 , \33484 , \33485 , \33486 , \33487 , \33488 , \33489 , \33490 , \33491 , \33492 ,
         \33493 , \33494 , \33495 , \33496 , \33497 , \33498 , \33499 , \33500 , \33501 , \33502 ,
         \33503 , \33504 , \33505 , \33506 , \33507 , \33508 , \33509 , \33510 , \33511 , \33512 ,
         \33513 , \33514 , \33515 , \33516 , \33517 , \33518 , \33519 , \33520 , \33521 , \33522 ,
         \33523 , \33524 , \33525 , \33526 , \33527 , \33528 , \33529 , \33530 , \33531 , \33532 ,
         \33533 , \33534 , \33535 , \33536 , \33537 , \33538 , \33539 , \33540 , \33541 , \33542 ,
         \33543 , \33544 , \33545 , \33546 , \33547 , \33548 , \33549 , \33550 , \33551 , \33552 ,
         \33553 , \33554 , \33555 , \33556 , \33557 , \33558 , \33559 , \33560 , \33561 , \33562 ,
         \33563 , \33564 , \33565 , \33566 , \33567 , \33568 , \33569 , \33570 , \33571 , \33572 ,
         \33573 , \33574 , \33575 , \33576 , \33577 , \33578 , \33579 , \33580 , \33581 , \33582 ,
         \33583 , \33584 , \33585 , \33586 , \33587 , \33588 , \33589 , \33590 , \33591 , \33592 ,
         \33593 , \33594 , \33595 , \33596 , \33597 , \33598 , \33599 , \33600 , \33601 , \33602 ,
         \33603 , \33604 , \33605 , \33606 , \33607 , \33608 , \33609 , \33610 , \33611 , \33612 ,
         \33613 , \33614 , \33615 , \33616 , \33617 , \33618 , \33619 , \33620 , \33621 , \33622 ,
         \33623 , \33624 , \33625 , \33626 , \33627 , \33628 , \33629 , \33630 , \33631 , \33632 ,
         \33633 , \33634 , \33635 , \33636 , \33637 , \33638 , \33639 , \33640 , \33641 , \33642 ,
         \33643 , \33644 , \33645 , \33646 , \33647 , \33648 , \33649 , \33650 , \33651 , \33652 ,
         \33653 , \33654 , \33655 , \33656 , \33657 , \33658 , \33659 , \33660 , \33661 , \33662 ,
         \33663 , \33664 , \33665 , \33666 , \33667 , \33668 , \33669 , \33670 , \33671 , \33672 ,
         \33673 , \33674 , \33675 , \33676 , \33677 , \33678 , \33679 , \33680 , \33681 , \33682 ,
         \33683 , \33684 , \33685 , \33686 , \33687 , \33688 , \33689 , \33690 , \33691 , \33692 ,
         \33693 , \33694 , \33695 , \33696 , \33697 , \33698 , \33699 , \33700 , \33701 , \33702 ,
         \33703 , \33704 , \33705 , \33706 , \33707 , \33708 , \33709 , \33710 , \33711 , \33712 ,
         \33713 , \33714 , \33715 , \33716 , \33717 , \33718 , \33719 , \33720 , \33721 , \33722 ,
         \33723 , \33724 , \33725 , \33726 , \33727 , \33728 , \33729 , \33730 , \33731 , \33732 ,
         \33733 , \33734 , \33735 , \33736 , \33737 , \33738 , \33739 , \33740 , \33741 , \33742 ,
         \33743 , \33744 , \33745 , \33746 , \33747 , \33748 , \33749 , \33750 , \33751 , \33752 ,
         \33753 , \33754 , \33755 , \33756 , \33757 , \33758 , \33759 , \33760 , \33761 , \33762 ,
         \33763 , \33764 , \33765 , \33766 , \33767 , \33768 , \33769 , \33770 , \33771 , \33772 ,
         \33773 , \33774 , \33775 , \33776 , \33777 , \33778 , \33779 , \33780 , \33781 , \33782 ,
         \33783 , \33784 , \33785 , \33786 , \33787 , \33788 , \33789 , \33790 , \33791 , \33792 ,
         \33793 , \33794 , \33795 , \33796 , \33797 , \33798 , \33799 , \33800 , \33801 , \33802 ,
         \33803 , \33804 , \33805 , \33806 , \33807 , \33808 , \33809 , \33810 , \33811 , \33812 ,
         \33813 , \33814 , \33815 , \33816 , \33817 , \33818 , \33819 , \33820 , \33821 , \33822 ,
         \33823 , \33824 , \33825 , \33826 , \33827 , \33828 , \33829 , \33830 , \33831 , \33832 ,
         \33833 , \33834 , \33835 , \33836 , \33837 , \33838 , \33839 , \33840 , \33841 , \33842 ,
         \33843 , \33844 , \33845 , \33846 , \33847 , \33848 , \33849 , \33850 , \33851 , \33852 ,
         \33853 , \33854 , \33855 , \33856 , \33857 , \33858 , \33859 , \33860 , \33861 , \33862 ,
         \33863 , \33864 , \33865 , \33866 , \33867 , \33868 , \33869 , \33870 , \33871 , \33872 ,
         \33873 , \33874 , \33875 , \33876 , \33877 , \33878 , \33879 , \33880 , \33881 , \33882 ,
         \33883 , \33884 , \33885 , \33886 , \33887 , \33888 , \33889 , \33890 , \33891 , \33892 ,
         \33893 , \33894 , \33895 , \33896 , \33897 , \33898 , \33899 , \33900 , \33901 , \33902 ,
         \33903 , \33904 , \33905 , \33906 , \33907 , \33908 , \33909 , \33910 , \33911 , \33912 ,
         \33913 , \33914 , \33915 , \33916 , \33917 , \33918 , \33919 , \33920 , \33921 , \33922 ,
         \33923 , \33924 , \33925 , \33926 , \33927 , \33928 , \33929 , \33930 , \33931 , \33932 ,
         \33933 , \33934 , \33935 , \33936 , \33937 , \33938 , \33939 , \33940 , \33941 , \33942 ,
         \33943 , \33944 , \33945 , \33946 , \33947 , \33948 , \33949 , \33950 , \33951 , \33952 ,
         \33953 , \33954 , \33955 , \33956 , \33957 , \33958 , \33959 , \33960 , \33961 , \33962 ,
         \33963 , \33964 , \33965 , \33966 , \33967 , \33968 , \33969 , \33970 , \33971 , \33972 ,
         \33973 , \33974 , \33975 , \33976 , \33977 , \33978 , \33979 , \33980 , \33981 , \33982 ,
         \33983 , \33984 , \33985 , \33986 , \33987 , \33988 , \33989 , \33990 , \33991 , \33992 ,
         \33993 , \33994 , \33995 , \33996 , \33997 , \33998 , \33999 , \34000 , \34001 , \34002 ,
         \34003 , \34004 , \34005 , \34006 , \34007 , \34008 , \34009 , \34010 , \34011 , \34012 ,
         \34013 , \34014 , \34015 , \34016 , \34017 , \34018 , \34019 , \34020 , \34021 , \34022 ,
         \34023 , \34024 , \34025 , \34026 , \34027 , \34028 , \34029 , \34030 , \34031 , \34032 ,
         \34033 , \34034 , \34035 , \34036 , \34037 , \34038 , \34039 , \34040 , \34041 , \34042 ,
         \34043 , \34044 , \34045 , \34046 , \34047 , \34048 , \34049 , \34050 , \34051 , \34052 ,
         \34053 , \34054 , \34055 , \34056 , \34057 , \34058 , \34059 , \34060 , \34061 , \34062 ,
         \34063 , \34064 , \34065 , \34066 , \34067 , \34068 , \34069 , \34070 , \34071 , \34072 ,
         \34073 , \34074 , \34075 , \34076 , \34077 , \34078 , \34079 , \34080 , \34081 , \34082 ,
         \34083 , \34084 , \34085 , \34086 , \34087 , \34088 , \34089 , \34090 , \34091 , \34092 ,
         \34093 , \34094 , \34095 , \34096 , \34097 , \34098 , \34099 , \34100 , \34101 , \34102 ,
         \34103 , \34104 , \34105 , \34106 , \34107 , \34108 , \34109 , \34110 , \34111 , \34112 ,
         \34113 , \34114 , \34115 , \34116 , \34117 , \34118 , \34119 , \34120 , \34121 , \34122 ,
         \34123 , \34124 , \34125 , \34126 , \34127 , \34128 , \34129 , \34130 , \34131 , \34132 ,
         \34133 , \34134 , \34135 , \34136 , \34137 , \34138 , \34139 , \34140 , \34141 , \34142 ,
         \34143 , \34144 , \34145 , \34146 , \34147 , \34148 , \34149 , \34150 , \34151 , \34152 ,
         \34153 , \34154 , \34155 , \34156 , \34157 , \34158 , \34159 , \34160 , \34161 , \34162 ,
         \34163 , \34164 , \34165 , \34166 , \34167 , \34168 , \34169 , \34170 , \34171 , \34172 ,
         \34173 , \34174 , \34175 , \34176 , \34177 , \34178 , \34179 , \34180 , \34181 , \34182 ,
         \34183 , \34184 , \34185 , \34186 , \34187 , \34188 , \34189 , \34190 , \34191 , \34192 ,
         \34193 , \34194 , \34195 , \34196 , \34197 , \34198 , \34199 , \34200 , \34201 , \34202 ,
         \34203 , \34204 , \34205 , \34206 , \34207 , \34208 , \34209 , \34210 , \34211 , \34212 ,
         \34213 , \34214 , \34215 , \34216 , \34217 , \34218 , \34219 , \34220 , \34221 , \34222 ,
         \34223 , \34224 , \34225 , \34226 , \34227 , \34228 , \34229 , \34230 , \34231 , \34232 ,
         \34233 , \34234 , \34235 , \34236 , \34237 , \34238 , \34239 , \34240 , \34241 , \34242 ,
         \34243 , \34244 , \34245 , \34246 , \34247 , \34248 , \34249 , \34250 , \34251 , \34252 ,
         \34253 , \34254 , \34255 , \34256 , \34257 , \34258 , \34259 , \34260 , \34261 , \34262 ,
         \34263 , \34264 , \34265 , \34266 , \34267 , \34268 , \34269 , \34270 , \34271 , \34272 ,
         \34273 , \34274 , \34275 , \34276 , \34277 , \34278 , \34279 , \34280 , \34281 , \34282 ,
         \34283 , \34284 , \34285 , \34286 , \34287 , \34288 , \34289 , \34290 , \34291 , \34292 ,
         \34293 , \34294 , \34295 , \34296 , \34297 , \34298 , \34299 , \34300 , \34301 , \34302 ,
         \34303 , \34304 , \34305 , \34306 , \34307 , \34308 , \34309 , \34310 , \34311 , \34312 ,
         \34313 , \34314 , \34315 , \34316 , \34317 , \34318 , \34319 , \34320 , \34321 , \34322 ,
         \34323 , \34324 , \34325 , \34326 , \34327 , \34328 , \34329 , \34330 , \34331 , \34332 ,
         \34333 , \34334 , \34335 , \34336 , \34337 , \34338 , \34339 , \34340 , \34341 , \34342 ,
         \34343 , \34344 , \34345 , \34346 , \34347 , \34348 , \34349 , \34350 , \34351 , \34352 ,
         \34353 , \34354 , \34355 , \34356 , \34357 , \34358 , \34359 , \34360 , \34361 , \34362 ,
         \34363 , \34364 , \34365 , \34366 , \34367 , \34368 , \34369 , \34370 , \34371 , \34372 ,
         \34373 , \34374 , \34375 , \34376 , \34377 , \34378 , \34379 , \34380 , \34381 , \34382 ,
         \34383 , \34384 , \34385 , \34386 , \34387 , \34388 , \34389 , \34390 , \34391 , \34392 ,
         \34393 , \34394 , \34395 , \34396 , \34397 , \34398 , \34399 , \34400 , \34401 , \34402 ,
         \34403 , \34404 , \34405 , \34406 , \34407 , \34408 , \34409 , \34410 , \34411 , \34412 ,
         \34413 , \34414 , \34415 , \34416 , \34417 , \34418 , \34419 , \34420 , \34421 , \34422 ,
         \34423 , \34424 , \34425 , \34426 , \34427 , \34428 , \34429 , \34430 , \34431 , \34432 ,
         \34433 , \34434 , \34435 , \34436 , \34437 , \34438 , \34439 , \34440 , \34441 , \34442 ,
         \34443 , \34444 , \34445 , \34446 , \34447 , \34448 , \34449 , \34450 , \34451 , \34452 ,
         \34453 , \34454 , \34455 , \34456 , \34457 , \34458 , \34459 , \34460 , \34461 , \34462 ,
         \34463 , \34464 , \34465 , \34466 , \34467 , \34468 , \34469 , \34470 , \34471 , \34472 ,
         \34473 , \34474 , \34475 , \34476 , \34477 , \34478 , \34479 , \34480 , \34481 , \34482 ,
         \34483 , \34484 , \34485 , \34486 , \34487 , \34488 , \34489 , \34490 , \34491 , \34492 ,
         \34493 , \34494 , \34495 , \34496 , \34497 , \34498 , \34499 , \34500 , \34501 , \34502 ,
         \34503 , \34504 , \34505 , \34506 , \34507 , \34508 , \34509 , \34510 , \34511 , \34512 ,
         \34513 , \34514 , \34515 , \34516 , \34517 , \34518 , \34519 , \34520 , \34521 , \34522 ,
         \34523 , \34524 , \34525 , \34526 , \34527 , \34528 , \34529 , \34530 , \34531 , \34532 ,
         \34533 , \34534 , \34535 , \34536 , \34537 , \34538 , \34539 , \34540 , \34541 , \34542 ,
         \34543 , \34544 , \34545 , \34546 , \34547 , \34548 , \34549 , \34550 , \34551 , \34552 ,
         \34553 , \34554 , \34555 , \34556 , \34557 , \34558 , \34559 , \34560 , \34561 , \34562 ,
         \34563 , \34564 , \34565 , \34566 , \34567 , \34568 , \34569 , \34570 , \34571 , \34572 ,
         \34573 , \34574 , \34575 , \34576 , \34577 , \34578 , \34579 , \34580 , \34581 , \34582 ,
         \34583 , \34584 , \34585 , \34586 , \34587 , \34588 , \34589 , \34590 , \34591 , \34592 ,
         \34593 , \34594 , \34595 , \34596 , \34597 , \34598 , \34599 , \34600 , \34601 , \34602 ,
         \34603 , \34604 , \34605 , \34606 , \34607 , \34608 , \34609 , \34610 , \34611 , \34612 ,
         \34613 , \34614 , \34615 , \34616 , \34617 , \34618 , \34619 , \34620 , \34621 , \34622 ,
         \34623 , \34624 , \34625 , \34626 , \34627 , \34628 , \34629 , \34630 , \34631 , \34632 ,
         \34633 , \34634 , \34635 , \34636 , \34637 , \34638 , \34639 , \34640 , \34641 , \34642 ,
         \34643 , \34644 , \34645 , \34646 , \34647 , \34648 , \34649 , \34650 , \34651 , \34652 ,
         \34653 , \34654 , \34655 , \34656 , \34657 , \34658 , \34659 , \34660 , \34661 , \34662 ,
         \34663 , \34664 , \34665 , \34666 , \34667 , \34668 , \34669 , \34670 , \34671 , \34672 ,
         \34673 , \34674 , \34675 , \34676 , \34677 , \34678 , \34679 , \34680 , \34681 , \34682 ,
         \34683 , \34684 , \34685 , \34686 , \34687 , \34688 , \34689 , \34690 , \34691 , \34692 ,
         \34693 , \34694 , \34695 , \34696 , \34697 , \34698 , \34699 , \34700 , \34701 , \34702 ,
         \34703 , \34704 , \34705 , \34706 , \34707 , \34708 , \34709 , \34710 , \34711 , \34712 ,
         \34713 , \34714 , \34715 , \34716 , \34717 , \34718 , \34719 , \34720 , \34721 , \34722 ,
         \34723 , \34724 , \34725 , \34726 , \34727 , \34728 , \34729 , \34730 , \34731 , \34732 ,
         \34733 , \34734 , \34735 , \34736 , \34737 , \34738 , \34739 , \34740 , \34741 , \34742 ,
         \34743 , \34744 , \34745 , \34746 , \34747 , \34748 , \34749 , \34750 , \34751 , \34752 ,
         \34753 , \34754 , \34755 , \34756 , \34757 , \34758 , \34759 , \34760 , \34761 , \34762 ,
         \34763 , \34764 , \34765 , \34766 , \34767 , \34768 , \34769 , \34770 , \34771 , \34772 ,
         \34773 , \34774 , \34775 , \34776 , \34777 , \34778 , \34779 , \34780 , \34781 , \34782 ,
         \34783 , \34784 , \34785 , \34786 , \34787 , \34788 , \34789 , \34790 , \34791 , \34792 ,
         \34793 , \34794 , \34795 , \34796 , \34797 , \34798 , \34799 , \34800 , \34801 , \34802 ,
         \34803 , \34804 , \34805 , \34806 , \34807 , \34808 , \34809 , \34810 , \34811 , \34812 ,
         \34813 , \34814 , \34815 , \34816 , \34817 , \34818 , \34819 , \34820 , \34821 , \34822 ,
         \34823 , \34824 , \34825 , \34826 , \34827 , \34828 , \34829 , \34830 , \34831 , \34832 ,
         \34833 , \34834 , \34835 , \34836 , \34837 , \34838 , \34839 , \34840 , \34841 , \34842 ,
         \34843 , \34844 , \34845 , \34846 , \34847 , \34848 , \34849 , \34850 , \34851 , \34852 ,
         \34853 , \34854 , \34855 , \34856 , \34857 , \34858 , \34859 , \34860 , \34861 , \34862 ,
         \34863 , \34864 , \34865 , \34866 , \34867 , \34868 , \34869 , \34870 , \34871 , \34872 ,
         \34873 , \34874 , \34875 , \34876 , \34877 , \34878 , \34879 , \34880 , \34881 , \34882 ,
         \34883 , \34884 , \34885 , \34886 , \34887 , \34888 , \34889 , \34890 , \34891 , \34892 ,
         \34893 , \34894 , \34895 , \34896 , \34897 , \34898 , \34899 , \34900 , \34901 , \34902 ,
         \34903 , \34904 , \34905 , \34906 , \34907 , \34908 , \34909 , \34910 , \34911 , \34912 ,
         \34913 , \34914 , \34915 , \34916 , \34917 , \34918 , \34919 , \34920 , \34921 , \34922 ,
         \34923 , \34924 , \34925 , \34926 , \34927 , \34928 , \34929 , \34930 , \34931 , \34932 ,
         \34933 , \34934 , \34935 , \34936 , \34937 , \34938 , \34939 , \34940 , \34941 , \34942 ,
         \34943 , \34944 , \34945 , \34946 , \34947 , \34948 , \34949 , \34950 , \34951 , \34952 ,
         \34953 , \34954 , \34955 , \34956 , \34957 , \34958 , \34959 , \34960 , \34961 , \34962 ,
         \34963 , \34964 , \34965 , \34966 , \34967 , \34968 , \34969 , \34970 , \34971 , \34972 ,
         \34973 , \34974 , \34975 , \34976 , \34977 , \34978 , \34979 , \34980 , \34981 , \34982 ,
         \34983 , \34984 , \34985 , \34986 , \34987 , \34988 , \34989 , \34990 , \34991 , \34992 ,
         \34993 , \34994 , \34995 , \34996 , \34997 , \34998 , \34999 , \35000 , \35001 , \35002 ,
         \35003 , \35004 , \35005 , \35006 , \35007 , \35008 , \35009 , \35010 , \35011 , \35012 ,
         \35013 , \35014 , \35015 , \35016 , \35017 , \35018 , \35019 , \35020 , \35021 , \35022 ,
         \35023 , \35024 , \35025 , \35026 , \35027 , \35028 , \35029 , \35030 , \35031 , \35032 ,
         \35033 , \35034 , \35035 , \35036 , \35037 , \35038 , \35039 , \35040 , \35041 , \35042 ,
         \35043 , \35044 , \35045 , \35046 , \35047 , \35048 , \35049 , \35050 , \35051 , \35052 ,
         \35053 , \35054 , \35055 , \35056 , \35057 , \35058 , \35059 , \35060 , \35061 , \35062 ,
         \35063 , \35064 , \35065 , \35066 , \35067 , \35068 , \35069 , \35070 , \35071 , \35072 ,
         \35073 , \35074 , \35075 , \35076 , \35077 , \35078 , \35079 , \35080 , \35081 , \35082 ,
         \35083 , \35084 , \35085 , \35086 , \35087 , \35088 , \35089 , \35090 , \35091 , \35092 ,
         \35093 , \35094 , \35095 , \35096 , \35097 , \35098 , \35099 , \35100 , \35101 , \35102 ,
         \35103 , \35104 , \35105 , \35106 , \35107 , \35108 , \35109 , \35110 , \35111 , \35112 ,
         \35113 , \35114 , \35115 , \35116 , \35117 , \35118 , \35119 , \35120 , \35121 , \35122 ,
         \35123 , \35124 , \35125 , \35126 , \35127 , \35128 , \35129 , \35130 , \35131 , \35132 ,
         \35133 , \35134 , \35135 , \35136 , \35137 , \35138 , \35139 , \35140 , \35141 , \35142 ,
         \35143 , \35144 , \35145 , \35146 , \35147 , \35148 , \35149 , \35150 , \35151 , \35152 ,
         \35153 , \35154 , \35155 , \35156 , \35157 , \35158 , \35159 , \35160 , \35161 , \35162 ,
         \35163 , \35164 , \35165 , \35166 , \35167 , \35168 , \35169 , \35170 , \35171 , \35172 ,
         \35173 , \35174 , \35175 , \35176 , \35177 , \35178 , \35179 , \35180 , \35181 , \35182 ,
         \35183 , \35184 , \35185 , \35186 , \35187 , \35188 , \35189 , \35190 , \35191 , \35192 ,
         \35193 , \35194 , \35195 , \35196 , \35197 , \35198 , \35199 , \35200 , \35201 , \35202 ,
         \35203 , \35204 , \35205 , \35206 , \35207 , \35208 , \35209 , \35210 , \35211 , \35212 ,
         \35213 , \35214 , \35215 , \35216 , \35217 , \35218 , \35219 , \35220 , \35221 , \35222 ,
         \35223 , \35224 , \35225 , \35226 , \35227 , \35228 , \35229 , \35230 , \35231 , \35232 ,
         \35233 , \35234 , \35235 , \35236 , \35237 , \35238 , \35239 , \35240 , \35241 , \35242 ,
         \35243 , \35244 , \35245 , \35246 , \35247 , \35248 , \35249 , \35250 , \35251 , \35252 ,
         \35253 , \35254 , \35255 , \35256 , \35257 , \35258 , \35259 , \35260 , \35261 , \35262 ,
         \35263 , \35264 , \35265 , \35266 , \35267 , \35268 , \35269 , \35270 , \35271 , \35272 ,
         \35273 , \35274 , \35275 , \35276 , \35277 , \35278 , \35279 , \35280 , \35281 , \35282 ,
         \35283 , \35284 , \35285 , \35286 , \35287 , \35288 , \35289 , \35290 , \35291 , \35292 ,
         \35293 , \35294 , \35295 , \35296 , \35297 , \35298 , \35299 , \35300 , \35301 , \35302 ,
         \35303 , \35304 , \35305 , \35306 , \35307 , \35308 , \35309 , \35310 , \35311 , \35312 ,
         \35313 , \35314 , \35315 , \35316 , \35317 , \35318 , \35319 , \35320 , \35321 , \35322 ,
         \35323 , \35324 , \35325 , \35326 , \35327 , \35328 , \35329 , \35330 , \35331 , \35332 ,
         \35333 , \35334 , \35335 , \35336 , \35337 , \35338 , \35339 , \35340 , \35341 , \35342 ,
         \35343 , \35344 , \35345 , \35346 , \35347 , \35348 , \35349 , \35350 , \35351 , \35352 ,
         \35353 , \35354 , \35355 , \35356 , \35357 , \35358 , \35359 , \35360 , \35361 , \35362 ,
         \35363 , \35364 , \35365 , \35366 , \35367 , \35368 , \35369 , \35370 , \35371 , \35372 ,
         \35373 , \35374 , \35375 , \35376 , \35377 , \35378 , \35379 , \35380 , \35381 , \35382 ,
         \35383 , \35384 , \35385 , \35386 , \35387 , \35388 , \35389 , \35390 , \35391 , \35392 ,
         \35393 , \35394 , \35395 , \35396 , \35397 , \35398 , \35399 , \35400 , \35401 , \35402 ,
         \35403 , \35404 , \35405 , \35406 , \35407 , \35408 , \35409 , \35410 , \35411 , \35412 ,
         \35413 , \35414 , \35415 , \35416 , \35417 , \35418 , \35419 , \35420 , \35421 , \35422 ,
         \35423 , \35424 , \35425 , \35426 , \35427 , \35428 , \35429 , \35430 , \35431 , \35432 ,
         \35433 , \35434 , \35435 , \35436 , \35437 , \35438 , \35439 , \35440 , \35441 , \35442 ,
         \35443 , \35444 , \35445 , \35446 , \35447 , \35448 , \35449 , \35450 , \35451 , \35452 ,
         \35453 , \35454 , \35455 , \35456 , \35457 , \35458 , \35459 , \35460 , \35461 , \35462 ,
         \35463 , \35464 , \35465 , \35466 , \35467 , \35468 , \35469 , \35470 , \35471 , \35472 ,
         \35473 , \35474 , \35475 , \35476 , \35477 , \35478 , \35479 , \35480 , \35481 , \35482 ,
         \35483 , \35484 , \35485 , \35486 , \35487 , \35488 , \35489 , \35490 , \35491 , \35492 ,
         \35493 , \35494 , \35495 , \35496 , \35497 , \35498 , \35499 , \35500 , \35501 , \35502 ,
         \35503 , \35504 , \35505 , \35506 , \35507 , \35508 , \35509 , \35510 , \35511 , \35512 ,
         \35513 , \35514 , \35515 , \35516 , \35517 , \35518 , \35519 , \35520 , \35521 , \35522 ,
         \35523 , \35524 , \35525 , \35526 , \35527 , \35528 , \35529 , \35530 , \35531 , \35532 ,
         \35533 , \35534 , \35535 , \35536 , \35537 , \35538 , \35539 , \35540 , \35541 , \35542 ,
         \35543 , \35544 , \35545 , \35546 , \35547 , \35548 , \35549 , \35550 , \35551 , \35552 ,
         \35553 , \35554 , \35555 , \35556 , \35557 , \35558 , \35559 , \35560 , \35561 , \35562 ,
         \35563 , \35564 , \35565 , \35566 , \35567 , \35568 , \35569 , \35570 , \35571 , \35572 ,
         \35573 , \35574 , \35575 , \35576 , \35577 , \35578 , \35579 , \35580 , \35581 , \35582 ,
         \35583 , \35584 , \35585 , \35586 , \35587 , \35588 , \35589 , \35590 , \35591 , \35592 ,
         \35593 , \35594 , \35595 , \35596 , \35597 , \35598 , \35599 , \35600 , \35601 , \35602 ,
         \35603 , \35604 , \35605 , \35606 , \35607 , \35608 , \35609 , \35610 , \35611 , \35612 ,
         \35613 , \35614 , \35615 , \35616 , \35617 , \35618 , \35619 , \35620 , \35621 , \35622 ,
         \35623 , \35624 , \35625 , \35626 , \35627 , \35628 , \35629 , \35630 , \35631 , \35632 ,
         \35633 , \35634 , \35635 , \35636 , \35637 , \35638 , \35639 , \35640 , \35641 , \35642 ,
         \35643 , \35644 , \35645 , \35646 , \35647 , \35648 , \35649 , \35650 , \35651 , \35652 ,
         \35653 , \35654 , \35655 , \35656 , \35657 , \35658 , \35659 , \35660 , \35661 , \35662 ,
         \35663 , \35664 , \35665 , \35666 , \35667 , \35668 , \35669 , \35670 , \35671 , \35672 ,
         \35673 , \35674 , \35675 , \35676 , \35677 , \35678 , \35679 , \35680 , \35681 , \35682 ,
         \35683 , \35684 , \35685 , \35686 , \35687 , \35688 , \35689 , \35690 , \35691 , \35692 ,
         \35693 , \35694 , \35695 , \35696 , \35697 , \35698 , \35699 , \35700 , \35701 , \35702 ,
         \35703 , \35704 , \35705 , \35706 , \35707 , \35708 , \35709 , \35710 , \35711 , \35712 ,
         \35713 , \35714 , \35715 , \35716 , \35717 , \35718 , \35719 , \35720 , \35721 , \35722 ,
         \35723 , \35724 , \35725 , \35726 , \35727 , \35728 , \35729 , \35730 , \35731 , \35732 ,
         \35733 , \35734 , \35735 , \35736 , \35737 , \35738 , \35739 , \35740 , \35741 , \35742 ,
         \35743 , \35744 , \35745 , \35746 , \35747 , \35748 , \35749 , \35750 , \35751 , \35752 ,
         \35753 , \35754 , \35755 , \35756 , \35757 , \35758 , \35759 , \35760 , \35761 , \35762 ,
         \35763 , \35764 , \35765 , \35766 , \35767 , \35768 , \35769 , \35770 , \35771 , \35772 ,
         \35773 , \35774 , \35775 , \35776 , \35777 , \35778 , \35779 , \35780 , \35781 , \35782 ,
         \35783 , \35784 , \35785 , \35786 , \35787 , \35788 , \35789 , \35790 , \35791 , \35792 ,
         \35793 , \35794 , \35795 , \35796 , \35797 , \35798 , \35799 , \35800 , \35801 , \35802 ,
         \35803 , \35804 , \35805 , \35806 , \35807 , \35808 , \35809 , \35810 , \35811 , \35812 ,
         \35813 , \35814 , \35815 , \35816 , \35817 , \35818 , \35819 , \35820 , \35821 , \35822 ,
         \35823 , \35824 , \35825 , \35826 , \35827 , \35828 , \35829 , \35830 , \35831 , \35832 ,
         \35833 , \35834 , \35835 , \35836 , \35837 , \35838 , \35839 , \35840 , \35841 , \35842 ,
         \35843 , \35844 , \35845 , \35846 , \35847 , \35848 , \35849 , \35850 , \35851 , \35852 ,
         \35853 , \35854 , \35855 , \35856 , \35857 , \35858 , \35859 , \35860 , \35861 , \35862 ,
         \35863 , \35864 , \35865 , \35866 , \35867 , \35868 , \35869 , \35870 , \35871 , \35872 ,
         \35873 , \35874 , \35875 , \35876 , \35877 , \35878 , \35879 , \35880 , \35881 , \35882 ,
         \35883 , \35884 , \35885 , \35886 , \35887 , \35888 , \35889 , \35890 , \35891 , \35892 ,
         \35893 , \35894 , \35895 , \35896 , \35897 , \35898 , \35899 , \35900 , \35901 , \35902 ,
         \35903 , \35904 , \35905 , \35906 , \35907 , \35908 , \35909 , \35910 , \35911 , \35912 ,
         \35913 , \35914 , \35915 , \35916 , \35917 , \35918 , \35919 , \35920 , \35921 , \35922 ,
         \35923 , \35924 , \35925 , \35926 , \35927 , \35928 , \35929 , \35930 , \35931 , \35932 ,
         \35933 , \35934 , \35935 , \35936 , \35937 , \35938 , \35939 , \35940 , \35941 , \35942 ,
         \35943 , \35944 , \35945 , \35946 , \35947 , \35948 , \35949 , \35950 , \35951 , \35952 ,
         \35953 , \35954 , \35955 , \35956 , \35957 , \35958 , \35959 , \35960 , \35961 , \35962 ,
         \35963 , \35964 , \35965 , \35966 , \35967 , \35968 , \35969 , \35970 , \35971 , \35972 ,
         \35973 , \35974 , \35975 , \35976 , \35977 , \35978 , \35979 , \35980 , \35981 , \35982 ,
         \35983 , \35984 , \35985 , \35986 , \35987 , \35988 , \35989 , \35990 , \35991 , \35992 ,
         \35993 , \35994 , \35995 , \35996 , \35997 , \35998 , \35999 , \36000 , \36001 , \36002 ,
         \36003 , \36004 , \36005 , \36006 , \36007 , \36008 , \36009 , \36010 , \36011 , \36012 ,
         \36013 , \36014 , \36015 , \36016 , \36017 , \36018 , \36019 , \36020 , \36021 , \36022 ,
         \36023 , \36024 , \36025 , \36026 , \36027 , \36028 , \36029 , \36030 , \36031 , \36032 ,
         \36033 , \36034 , \36035 , \36036 , \36037 , \36038 , \36039 , \36040 , \36041 , \36042 ,
         \36043 , \36044 , \36045 , \36046 , \36047 , \36048 , \36049 , \36050 , \36051 , \36052 ,
         \36053 , \36054 , \36055 , \36056 , \36057 , \36058 , \36059 , \36060 , \36061 , \36062 ,
         \36063 , \36064 , \36065 , \36066 , \36067 , \36068 , \36069 , \36070 , \36071 , \36072 ,
         \36073 , \36074 , \36075 , \36076 , \36077 , \36078 , \36079 , \36080 , \36081 , \36082 ,
         \36083 , \36084 , \36085 , \36086 , \36087 , \36088 , \36089 , \36090 , \36091 , \36092 ,
         \36093 , \36094 , \36095 , \36096 , \36097 , \36098 , \36099 , \36100 , \36101 , \36102 ,
         \36103 , \36104 , \36105 , \36106 , \36107 , \36108 , \36109 , \36110 , \36111 , \36112 ,
         \36113 , \36114 , \36115 , \36116 , \36117 , \36118 , \36119 , \36120 , \36121 , \36122 ,
         \36123 , \36124 , \36125 , \36126 , \36127 , \36128 , \36129 , \36130 , \36131 , \36132 ,
         \36133 , \36134 , \36135 , \36136 , \36137 , \36138 , \36139 , \36140 , \36141 , \36142 ,
         \36143 , \36144 , \36145 , \36146 , \36147 , \36148 , \36149 , \36150 , \36151 , \36152 ,
         \36153 , \36154 , \36155 , \36156 , \36157 , \36158 , \36159 , \36160 , \36161 , \36162 ,
         \36163 , \36164 , \36165 , \36166 , \36167 , \36168 , \36169 , \36170 , \36171 , \36172 ,
         \36173 , \36174 , \36175 , \36176 , \36177 , \36178 , \36179 , \36180 , \36181 , \36182 ,
         \36183 , \36184 , \36185 , \36186 , \36187 , \36188 , \36189 , \36190 , \36191 , \36192 ,
         \36193 , \36194 , \36195 , \36196 , \36197 , \36198 , \36199 , \36200 , \36201 , \36202 ,
         \36203 , \36204 , \36205 , \36206 , \36207 , \36208 , \36209 , \36210 , \36211 , \36212 ,
         \36213 , \36214 , \36215 , \36216 , \36217 , \36218 , \36219 , \36220 , \36221 , \36222 ,
         \36223 , \36224 , \36225 , \36226 , \36227 , \36228 , \36229 , \36230 , \36231 , \36232 ,
         \36233 , \36234 , \36235 , \36236 , \36237 , \36238 , \36239 , \36240 , \36241 , \36242 ,
         \36243 , \36244 , \36245 , \36246 , \36247 , \36248 , \36249 , \36250 , \36251 , \36252 ,
         \36253 , \36254 , \36255 , \36256 , \36257 , \36258 , \36259 , \36260 , \36261 , \36262 ,
         \36263 , \36264 , \36265 , \36266 , \36267 , \36268 , \36269 , \36270 , \36271 , \36272 ,
         \36273 , \36274 , \36275 , \36276 , \36277 , \36278 , \36279 , \36280 , \36281 , \36282 ,
         \36283 , \36284 , \36285 , \36286 , \36287 , \36288 , \36289 , \36290 , \36291 , \36292 ,
         \36293 , \36294 , \36295 , \36296 , \36297 , \36298 , \36299 , \36300 , \36301 , \36302 ,
         \36303 , \36304 , \36305 , \36306 , \36307 , \36308 , \36309 , \36310 , \36311 , \36312 ,
         \36313 , \36314 , \36315 , \36316 , \36317 , \36318 , \36319 , \36320 , \36321 , \36322 ,
         \36323 , \36324 , \36325 , \36326 , \36327 , \36328 , \36329 , \36330 , \36331 , \36332 ,
         \36333 , \36334 , \36335 , \36336 , \36337 , \36338 , \36339 , \36340 , \36341 , \36342 ,
         \36343 , \36344 , \36345 , \36346 , \36347 , \36348 , \36349 , \36350 , \36351 , \36352 ,
         \36353 , \36354 , \36355 , \36356 , \36357 , \36358 , \36359 , \36360 , \36361 , \36362 ,
         \36363 , \36364 , \36365 , \36366 , \36367 , \36368 , \36369 , \36370 , \36371 , \36372 ,
         \36373 , \36374 , \36375 , \36376 , \36377 , \36378 , \36379 , \36380 , \36381 , \36382 ,
         \36383 , \36384 , \36385 , \36386 , \36387 , \36388 , \36389 , \36390 , \36391 , \36392 ,
         \36393 , \36394 , \36395 , \36396 , \36397 , \36398 , \36399 , \36400 , \36401 , \36402 ,
         \36403 , \36404 , \36405 , \36406 , \36407 , \36408 , \36409 , \36410 , \36411 , \36412 ,
         \36413 , \36414 , \36415 , \36416 , \36417 , \36418 , \36419 , \36420 , \36421 , \36422 ,
         \36423 , \36424 , \36425 , \36426 , \36427 , \36428 , \36429 , \36430 , \36431 , \36432 ,
         \36433 , \36434 , \36435 , \36436 , \36437 , \36438 , \36439 , \36440 , \36441 , \36442 ,
         \36443 , \36444 , \36445 , \36446 , \36447 , \36448 , \36449 , \36450 , \36451 , \36452 ,
         \36453 , \36454 , \36455 , \36456 , \36457 , \36458 , \36459 , \36460 , \36461 , \36462 ,
         \36463 , \36464 , \36465 , \36466 , \36467 , \36468 , \36469 , \36470 , \36471 , \36472 ,
         \36473 , \36474 , \36475 , \36476 , \36477 , \36478 , \36479 , \36480 , \36481 , \36482 ,
         \36483 , \36484 , \36485 , \36486 , \36487 , \36488 , \36489 , \36490 , \36491 , \36492 ,
         \36493 , \36494 , \36495 , \36496 , \36497 , \36498 , \36499 , \36500 , \36501 , \36502 ,
         \36503 , \36504 , \36505 , \36506 , \36507 , \36508 , \36509 , \36510 , \36511 , \36512 ,
         \36513 , \36514 , \36515 , \36516 , \36517 , \36518 , \36519 , \36520 , \36521 , \36522 ,
         \36523 , \36524 , \36525 , \36526 , \36527 , \36528 , \36529 , \36530 , \36531 , \36532 ,
         \36533 , \36534 , \36535 , \36536 , \36537 , \36538 , \36539 , \36540 , \36541 , \36542 ,
         \36543 , \36544 , \36545 , \36546 , \36547 , \36548 , \36549 , \36550 , \36551 , \36552 ,
         \36553 , \36554 , \36555 , \36556 , \36557 , \36558 , \36559 , \36560 , \36561 , \36562 ,
         \36563 , \36564 , \36565 , \36566 , \36567 , \36568 , \36569 , \36570 , \36571 , \36572 ,
         \36573 , \36574 , \36575 , \36576 , \36577 , \36578 , \36579 , \36580 , \36581 , \36582 ,
         \36583 , \36584 , \36585 , \36586 , \36587 , \36588 , \36589 , \36590 , \36591 , \36592 ,
         \36593 , \36594 , \36595 , \36596 , \36597 , \36598 , \36599 , \36600 , \36601 , \36602 ,
         \36603 , \36604 , \36605 , \36606 , \36607 , \36608 , \36609 , \36610 , \36611 , \36612 ,
         \36613 , \36614 , \36615 , \36616 , \36617 , \36618 , \36619 , \36620 , \36621 , \36622 ,
         \36623 , \36624 , \36625 , \36626 , \36627 , \36628 , \36629 , \36630 , \36631 , \36632 ,
         \36633 , \36634 , \36635 , \36636 , \36637 , \36638 , \36639 , \36640 , \36641 , \36642 ,
         \36643 , \36644 , \36645 , \36646 , \36647 , \36648 , \36649 , \36650 , \36651 , \36652 ,
         \36653 , \36654 , \36655 , \36656 , \36657 , \36658 , \36659 , \36660 , \36661 , \36662 ,
         \36663 , \36664 , \36665 , \36666 , \36667 , \36668 , \36669 , \36670 , \36671 , \36672 ,
         \36673 , \36674 , \36675 , \36676 , \36677 , \36678 , \36679 , \36680 , \36681 , \36682 ,
         \36683 , \36684 , \36685 , \36686 , \36687 , \36688 , \36689 , \36690 , \36691 , \36692 ,
         \36693 , \36694 , \36695 , \36696 , \36697 , \36698 , \36699 , \36700 , \36701 , \36702 ,
         \36703 , \36704 , \36705 , \36706 , \36707 , \36708 , \36709 , \36710 , \36711 , \36712 ,
         \36713 , \36714 , \36715 , \36716 , \36717 , \36718 , \36719 , \36720 , \36721 , \36722 ,
         \36723 , \36724 , \36725 , \36726 , \36727 , \36728 , \36729 , \36730 , \36731 , \36732 ,
         \36733 , \36734 , \36735 , \36736 , \36737 , \36738 , \36739 , \36740 , \36741 , \36742 ,
         \36743 , \36744 , \36745 , \36746 , \36747 , \36748 , \36749 , \36750 , \36751 , \36752 ,
         \36753 , \36754 , \36755 , \36756 , \36757 , \36758 , \36759 , \36760 , \36761 , \36762 ,
         \36763 , \36764 , \36765 , \36766 , \36767 , \36768 , \36769 , \36770 , \36771 , \36772 ,
         \36773 , \36774 , \36775 , \36776 , \36777 , \36778 , \36779 , \36780 , \36781 , \36782 ,
         \36783 , \36784 , \36785 , \36786 , \36787 , \36788 , \36789 , \36790 , \36791 , \36792 ,
         \36793 , \36794 , \36795 , \36796 , \36797 , \36798 , \36799 , \36800 , \36801 , \36802 ,
         \36803 , \36804 , \36805 , \36806 , \36807 , \36808 , \36809 , \36810 , \36811 , \36812 ,
         \36813 , \36814 , \36815 , \36816 , \36817 , \36818 , \36819 , \36820 , \36821 , \36822 ,
         \36823 , \36824 , \36825 , \36826 , \36827 , \36828 , \36829 , \36830 , \36831 , \36832 ,
         \36833 , \36834 , \36835 , \36836 , \36837 , \36838 , \36839 , \36840 , \36841 , \36842 ,
         \36843 , \36844 , \36845 , \36846 , \36847 , \36848 , \36849 , \36850 , \36851 , \36852 ,
         \36853 , \36854 , \36855 , \36856 , \36857 , \36858 , \36859 , \36860 , \36861 , \36862 ,
         \36863 , \36864 , \36865 , \36866 , \36867 , \36868 , \36869 , \36870 , \36871 , \36872 ,
         \36873 , \36874 , \36875 , \36876 , \36877 , \36878 , \36879 , \36880 , \36881 , \36882 ,
         \36883 , \36884 , \36885 , \36886 , \36887 , \36888 , \36889 , \36890 , \36891 , \36892 ,
         \36893 , \36894 , \36895 , \36896 , \36897 , \36898 , \36899 , \36900 , \36901 , \36902 ,
         \36903 , \36904 , \36905 , \36906 , \36907 , \36908 , \36909 , \36910 , \36911 , \36912 ,
         \36913 , \36914 , \36915 , \36916 , \36917 , \36918 , \36919 , \36920 , \36921 , \36922 ,
         \36923 , \36924 , \36925 , \36926 , \36927 , \36928 , \36929 , \36930 , \36931 , \36932 ,
         \36933 , \36934 , \36935 , \36936 , \36937 , \36938 , \36939 , \36940 , \36941 , \36942 ,
         \36943 , \36944 , \36945 , \36946 , \36947 , \36948 , \36949 , \36950 , \36951 , \36952 ,
         \36953 , \36954 , \36955 , \36956 , \36957 , \36958 , \36959 , \36960 , \36961 , \36962 ,
         \36963 , \36964 , \36965 , \36966 , \36967 , \36968 , \36969 , \36970 , \36971 , \36972 ,
         \36973 , \36974 , \36975 , \36976 , \36977 , \36978 , \36979 , \36980 , \36981 , \36982 ,
         \36983 , \36984 , \36985 , \36986 , \36987 , \36988 , \36989 , \36990 , \36991 , \36992 ,
         \36993 , \36994 , \36995 , \36996 , \36997 , \36998 , \36999 , \37000 , \37001 , \37002 ,
         \37003 , \37004 , \37005 , \37006 , \37007 , \37008 , \37009 , \37010 , \37011 , \37012 ,
         \37013 , \37014 , \37015 , \37016 , \37017 , \37018 , \37019 , \37020 , \37021 , \37022 ,
         \37023 , \37024 , \37025 , \37026 , \37027 , \37028 , \37029 , \37030 , \37031 , \37032 ,
         \37033 , \37034 , \37035 , \37036 , \37037 , \37038 , \37039 , \37040 , \37041 , \37042 ,
         \37043 , \37044 , \37045 , \37046 , \37047 , \37048 , \37049 , \37050 , \37051 , \37052 ,
         \37053 , \37054 , \37055 , \37056 , \37057 , \37058 , \37059 , \37060 , \37061 , \37062 ,
         \37063 , \37064 , \37065 , \37066 , \37067 , \37068 , \37069 , \37070 , \37071 , \37072 ,
         \37073 , \37074 , \37075 , \37076 , \37077 , \37078 , \37079 , \37080 , \37081 , \37082 ,
         \37083 , \37084 , \37085 , \37086 , \37087 , \37088 , \37089 , \37090 , \37091 , \37092 ,
         \37093 , \37094 , \37095 , \37096 , \37097 , \37098 , \37099 , \37100 , \37101 , \37102 ,
         \37103 , \37104 , \37105 , \37106 , \37107 , \37108 , \37109 , \37110 , \37111 , \37112 ,
         \37113 , \37114 , \37115 , \37116 , \37117 , \37118 , \37119 , \37120 , \37121 , \37122 ,
         \37123 , \37124 , \37125 , \37126 , \37127 , \37128 , \37129 , \37130 , \37131 , \37132 ,
         \37133 , \37134 , \37135 , \37136 , \37137 , \37138 , \37139 , \37140 , \37141 , \37142 ,
         \37143 , \37144 , \37145 , \37146 , \37147 , \37148 , \37149 , \37150 , \37151 , \37152 ,
         \37153 , \37154 , \37155 , \37156 , \37157 , \37158 , \37159 , \37160 , \37161 , \37162 ,
         \37163 , \37164 , \37165 , \37166 , \37167 , \37168 , \37169 , \37170 , \37171 , \37172 ,
         \37173 , \37174 , \37175 , \37176 , \37177 , \37178 , \37179 , \37180 , \37181 , \37182 ,
         \37183 , \37184 , \37185 , \37186 , \37187 , \37188 , \37189 , \37190 , \37191 , \37192 ,
         \37193 , \37194 , \37195 , \37196 , \37197 , \37198 , \37199 , \37200 , \37201 , \37202 ,
         \37203 , \37204 , \37205 , \37206 , \37207 , \37208 , \37209 , \37210 , \37211 , \37212 ,
         \37213 , \37214 , \37215 , \37216 , \37217 , \37218 , \37219 , \37220 , \37221 , \37222 ,
         \37223 , \37224 , \37225 , \37226 , \37227 , \37228 , \37229 , \37230 , \37231 , \37232 ,
         \37233 , \37234 , \37235 , \37236 , \37237 , \37238 , \37239 , \37240 , \37241 , \37242 ,
         \37243 , \37244 , \37245 , \37246 , \37247 , \37248 , \37249 , \37250 , \37251 , \37252 ,
         \37253 , \37254 , \37255 , \37256 , \37257 , \37258 , \37259 , \37260 , \37261 , \37262 ,
         \37263 , \37264 , \37265 , \37266 , \37267 , \37268 , \37269 , \37270 , \37271 , \37272 ,
         \37273 , \37274 , \37275 , \37276 , \37277 , \37278 , \37279 , \37280 , \37281 , \37282 ,
         \37283 , \37284 , \37285 , \37286 , \37287 , \37288 , \37289 , \37290 , \37291 , \37292 ,
         \37293 , \37294 , \37295 , \37296 , \37297 , \37298 , \37299 , \37300 , \37301 , \37302 ,
         \37303 , \37304 , \37305 , \37306 , \37307 , \37308 , \37309 , \37310 , \37311 , \37312 ,
         \37313 , \37314 , \37315 , \37316 , \37317 , \37318 , \37319 , \37320 , \37321 , \37322 ,
         \37323 , \37324 , \37325 , \37326 , \37327 , \37328 , \37329 , \37330 , \37331 , \37332 ,
         \37333 , \37334 , \37335 , \37336 , \37337 , \37338 , \37339 , \37340 , \37341 , \37342 ,
         \37343 , \37344 , \37345 , \37346 , \37347 , \37348 , \37349 , \37350 , \37351 , \37352 ,
         \37353 , \37354 , \37355 , \37356 , \37357 , \37358 , \37359 , \37360 , \37361 , \37362 ,
         \37363 , \37364 , \37365 , \37366 , \37367 , \37368 , \37369 , \37370 , \37371 , \37372 ,
         \37373 , \37374 , \37375 , \37376 , \37377 , \37378 , \37379 , \37380 , \37381 , \37382 ,
         \37383 , \37384 , \37385 , \37386 , \37387 , \37388 , \37389 , \37390 , \37391 , \37392 ,
         \37393 , \37394 , \37395 , \37396 , \37397 , \37398 , \37399 , \37400 , \37401 , \37402 ,
         \37403 , \37404 , \37405 , \37406 , \37407 , \37408 , \37409 , \37410 , \37411 , \37412 ,
         \37413 , \37414 , \37415 , \37416 , \37417 , \37418 , \37419 , \37420 , \37421 , \37422 ,
         \37423 , \37424 , \37425 , \37426 , \37427 , \37428 , \37429 , \37430 , \37431 , \37432 ,
         \37433 , \37434 , \37435 , \37436 , \37437 , \37438 , \37439 , \37440 , \37441 , \37442 ,
         \37443 , \37444 , \37445 , \37446 , \37447 , \37448 , \37449 , \37450 , \37451 , \37452 ,
         \37453 , \37454 , \37455 , \37456 , \37457 , \37458 , \37459 , \37460 , \37461 , \37462 ,
         \37463 , \37464 , \37465 , \37466 , \37467 , \37468 , \37469 , \37470 , \37471 , \37472 ,
         \37473 , \37474 , \37475 , \37476 , \37477 , \37478 , \37479 , \37480 , \37481 , \37482 ,
         \37483 , \37484 , \37485 , \37486 , \37487 , \37488 , \37489 , \37490 , \37491 , \37492 ,
         \37493 , \37494 , \37495 , \37496 , \37497 , \37498 , \37499 , \37500 , \37501 , \37502 ,
         \37503 , \37504 , \37505 , \37506 , \37507 , \37508 , \37509 , \37510 , \37511 , \37512 ,
         \37513 , \37514 , \37515 , \37516 , \37517 , \37518 , \37519 , \37520 , \37521 , \37522 ,
         \37523 , \37524 , \37525 , \37526 , \37527 , \37528 , \37529 , \37530 , \37531 , \37532 ,
         \37533 , \37534 , \37535 , \37536 , \37537 , \37538 , \37539 , \37540 , \37541 , \37542 ,
         \37543 , \37544 , \37545 , \37546 , \37547 , \37548 , \37549 , \37550 , \37551 , \37552 ,
         \37553 , \37554 , \37555 , \37556 , \37557 , \37558 , \37559 , \37560 , \37561 , \37562 ,
         \37563 , \37564 , \37565 , \37566 , \37567 , \37568 , \37569 , \37570 , \37571 , \37572 ,
         \37573 , \37574 , \37575 , \37576 , \37577 , \37578 , \37579 , \37580 , \37581 , \37582 ,
         \37583 , \37584 , \37585 , \37586 , \37587 , \37588 , \37589 , \37590 , \37591 , \37592 ,
         \37593 , \37594 , \37595 , \37596 , \37597 , \37598 , \37599 , \37600 , \37601 , \37602 ,
         \37603 , \37604 , \37605 , \37606 , \37607 , \37608 , \37609 , \37610 , \37611 , \37612 ,
         \37613 , \37614 , \37615 , \37616 , \37617 , \37618 , \37619 , \37620 , \37621 , \37622 ,
         \37623 , \37624 , \37625 , \37626 , \37627 , \37628 , \37629 , \37630 , \37631 , \37632 ,
         \37633 , \37634 , \37635 , \37636 , \37637 , \37638 , \37639 , \37640 , \37641 , \37642 ,
         \37643 , \37644 , \37645 , \37646 , \37647 , \37648 , \37649 , \37650 , \37651 , \37652 ,
         \37653 , \37654 , \37655 , \37656 , \37657 , \37658 , \37659 , \37660 , \37661 , \37662 ,
         \37663 , \37664 , \37665 , \37666 , \37667 , \37668 , \37669 , \37670 , \37671 , \37672 ,
         \37673 , \37674 , \37675 , \37676 , \37677 , \37678 , \37679 , \37680 , \37681 , \37682 ,
         \37683 , \37684 , \37685 , \37686 , \37687 , \37688 , \37689 , \37690 , \37691 , \37692 ,
         \37693 , \37694 , \37695 , \37696 , \37697 , \37698 , \37699 , \37700 , \37701 , \37702 ,
         \37703 , \37704 , \37705 , \37706 , \37707 , \37708 , \37709 , \37710 , \37711 , \37712 ,
         \37713 , \37714 , \37715 , \37716 , \37717 , \37718 , \37719 , \37720 , \37721 , \37722 ,
         \37723 , \37724 , \37725 , \37726 , \37727 , \37728 , \37729 , \37730 , \37731 , \37732 ,
         \37733 , \37734 , \37735 , \37736 , \37737 , \37738 , \37739 , \37740 , \37741 , \37742 ,
         \37743 , \37744 , \37745 , \37746 , \37747 , \37748 , \37749 , \37750 , \37751 , \37752 ,
         \37753 , \37754 , \37755 , \37756 , \37757 , \37758 , \37759 , \37760 , \37761 , \37762 ,
         \37763 , \37764 , \37765 , \37766 , \37767 , \37768 , \37769 , \37770 , \37771 , \37772 ,
         \37773 , \37774 , \37775 , \37776 , \37777 , \37778 , \37779 , \37780 , \37781 , \37782 ,
         \37783 , \37784 , \37785 , \37786 , \37787 , \37788 , \37789 , \37790 , \37791 , \37792 ,
         \37793 , \37794 , \37795 , \37796 , \37797 , \37798 , \37799 , \37800 , \37801 , \37802 ,
         \37803 , \37804 , \37805 , \37806 , \37807 , \37808 , \37809 , \37810 , \37811 , \37812 ,
         \37813 , \37814 , \37815 , \37816 , \37817 , \37818 , \37819 , \37820 , \37821 , \37822 ,
         \37823 , \37824 , \37825 , \37826 , \37827 , \37828 , \37829 , \37830 , \37831 , \37832 ,
         \37833 , \37834 , \37835 , \37836 , \37837 , \37838 , \37839 , \37840 , \37841 , \37842 ,
         \37843 , \37844 , \37845 , \37846 , \37847 , \37848 , \37849 , \37850 , \37851 , \37852 ,
         \37853 , \37854 , \37855 , \37856 , \37857 , \37858 , \37859 , \37860 , \37861 , \37862 ,
         \37863 , \37864 , \37865 , \37866 , \37867 , \37868 , \37869 , \37870 , \37871 , \37872 ,
         \37873 , \37874 , \37875 , \37876 , \37877 , \37878 , \37879 , \37880 , \37881 , \37882 ,
         \37883 , \37884 , \37885 , \37886 , \37887 , \37888 , \37889 , \37890 , \37891 , \37892 ,
         \37893 , \37894 , \37895 , \37896 , \37897 , \37898 , \37899 , \37900 , \37901 , \37902 ,
         \37903 , \37904 , \37905 , \37906 , \37907 , \37908 , \37909 , \37910 , \37911 , \37912 ,
         \37913 , \37914 , \37915 , \37916 , \37917 , \37918 , \37919 , \37920 , \37921 , \37922 ,
         \37923 , \37924 , \37925 , \37926 , \37927 , \37928 , \37929 , \37930 , \37931 , \37932 ,
         \37933 , \37934 , \37935 , \37936 , \37937 , \37938 , \37939 , \37940 , \37941 , \37942 ,
         \37943 , \37944 , \37945 , \37946 , \37947 , \37948 , \37949 , \37950 , \37951 , \37952 ,
         \37953 , \37954 , \37955 , \37956 , \37957 , \37958 , \37959 , \37960 , \37961 , \37962 ,
         \37963 , \37964 , \37965 , \37966 , \37967 , \37968 , \37969 , \37970 , \37971 , \37972 ,
         \37973 , \37974 , \37975 , \37976 , \37977 , \37978 , \37979 , \37980 , \37981 , \37982 ,
         \37983 , \37984 , \37985 , \37986 , \37987 , \37988 , \37989 , \37990 , \37991 , \37992 ,
         \37993 , \37994 , \37995 , \37996 , \37997 , \37998 , \37999 , \38000 , \38001 , \38002 ,
         \38003 , \38004 , \38005 , \38006 , \38007 , \38008 , \38009 , \38010 , \38011 , \38012 ,
         \38013 , \38014 , \38015 , \38016 , \38017 , \38018 , \38019 , \38020 , \38021 , \38022 ,
         \38023 , \38024 , \38025 , \38026 , \38027 , \38028 , \38029 , \38030 , \38031 , \38032 ,
         \38033 , \38034 , \38035 , \38036 , \38037 , \38038 , \38039 , \38040 , \38041 , \38042 ,
         \38043 , \38044 , \38045 , \38046 , \38047 , \38048 , \38049 , \38050 , \38051 , \38052 ,
         \38053 , \38054 , \38055 , \38056 , \38057 , \38058 , \38059 , \38060 , \38061 , \38062 ,
         \38063 , \38064 , \38065 , \38066 , \38067 , \38068 , \38069 , \38070 , \38071 , \38072 ,
         \38073 , \38074 , \38075 , \38076 , \38077 , \38078 , \38079 , \38080 , \38081 , \38082 ,
         \38083 , \38084 , \38085 , \38086 , \38087 , \38088 , \38089 , \38090 , \38091 , \38092 ,
         \38093 , \38094 , \38095 , \38096 , \38097 , \38098 , \38099 , \38100 , \38101 , \38102 ,
         \38103 , \38104 , \38105 , \38106 , \38107 , \38108 , \38109 , \38110 , \38111 , \38112 ,
         \38113 , \38114 , \38115 , \38116 , \38117 , \38118 , \38119 , \38120 , \38121 , \38122 ,
         \38123 , \38124 , \38125 , \38126 , \38127 , \38128 , \38129 , \38130 , \38131 , \38132 ,
         \38133 , \38134 , \38135 , \38136 , \38137 , \38138 , \38139 , \38140 , \38141 , \38142 ,
         \38143 , \38144 , \38145 , \38146 , \38147 , \38148 , \38149 , \38150 , \38151 , \38152 ,
         \38153 , \38154 , \38155 , \38156 , \38157 , \38158 , \38159 , \38160 , \38161 , \38162 ,
         \38163 , \38164 , \38165 , \38166 , \38167 , \38168 , \38169 , \38170 , \38171 , \38172 ,
         \38173 , \38174 , \38175 , \38176 , \38177 , \38178 , \38179 , \38180 , \38181 , \38182 ,
         \38183 , \38184 , \38185 , \38186 , \38187 , \38188 , \38189 , \38190 , \38191 , \38192 ,
         \38193 , \38194 , \38195 , \38196 , \38197 , \38198 , \38199 , \38200 , \38201 , \38202 ,
         \38203 , \38204 , \38205 , \38206 , \38207 , \38208 , \38209 , \38210 , \38211 , \38212 ,
         \38213 , \38214 , \38215 , \38216 , \38217 , \38218 , \38219 , \38220 , \38221 , \38222 ,
         \38223 , \38224 , \38225 , \38226 , \38227 , \38228 , \38229 , \38230 , \38231 , \38232 ,
         \38233 , \38234 , \38235 , \38236 , \38237 , \38238 , \38239 , \38240 , \38241 , \38242 ,
         \38243 , \38244 , \38245 , \38246 , \38247 , \38248 , \38249 , \38250 , \38251 , \38252 ,
         \38253 , \38254 , \38255 , \38256 , \38257 , \38258 , \38259 , \38260 , \38261 , \38262 ,
         \38263 , \38264 , \38265 , \38266 , \38267 , \38268 , \38269 , \38270 , \38271 , \38272 ,
         \38273 , \38274 , \38275 , \38276 , \38277 , \38278 , \38279 , \38280 , \38281 , \38282 ,
         \38283 , \38284 , \38285 , \38286 , \38287 , \38288 , \38289 , \38290 , \38291 , \38292 ,
         \38293 , \38294 , \38295 , \38296 , \38297 , \38298 , \38299 , \38300 , \38301 , \38302 ,
         \38303 , \38304 , \38305 , \38306 , \38307 , \38308 , \38309 , \38310 , \38311 , \38312 ,
         \38313 , \38314 , \38315 , \38316 , \38317 , \38318 , \38319 , \38320 , \38321 , \38322 ,
         \38323 , \38324 , \38325 , \38326 , \38327 , \38328 , \38329 , \38330 , \38331 , \38332 ,
         \38333 , \38334 , \38335 , \38336 , \38337 , \38338 , \38339 , \38340 , \38341 , \38342 ,
         \38343 , \38344 , \38345 , \38346 , \38347 , \38348 , \38349 , \38350 , \38351 , \38352 ,
         \38353 , \38354 , \38355 , \38356 , \38357 , \38358 , \38359 , \38360 , \38361 , \38362 ,
         \38363 , \38364 , \38365 , \38366 , \38367 , \38368 , \38369 , \38370 , \38371 , \38372 ,
         \38373 , \38374 , \38375 , \38376 , \38377 , \38378 , \38379 , \38380 , \38381 , \38382 ,
         \38383 , \38384 , \38385 , \38386 , \38387 , \38388 , \38389 , \38390 , \38391 , \38392 ,
         \38393 , \38394 , \38395 , \38396 , \38397 , \38398 , \38399 , \38400 , \38401 , \38402 ,
         \38403 , \38404 , \38405 , \38406 , \38407 , \38408 , \38409 , \38410 , \38411 , \38412 ,
         \38413 , \38414 , \38415 , \38416 , \38417 , \38418 , \38419 , \38420 , \38421 , \38422 ,
         \38423 , \38424 , \38425 , \38426 , \38427 , \38428 , \38429 , \38430 , \38431 , \38432 ,
         \38433 , \38434 , \38435 , \38436 , \38437 , \38438 , \38439 , \38440 , \38441 , \38442 ,
         \38443 , \38444 , \38445 , \38446 , \38447 , \38448 , \38449 , \38450 , \38451 , \38452 ,
         \38453 , \38454 , \38455 , \38456 , \38457 , \38458 , \38459 , \38460 , \38461 , \38462 ,
         \38463 , \38464 , \38465 , \38466 , \38467 , \38468 , \38469 , \38470 , \38471 , \38472 ,
         \38473 , \38474 , \38475 , \38476 , \38477 , \38478 , \38479 , \38480 , \38481 , \38482 ,
         \38483 , \38484 , \38485 , \38486 , \38487 , \38488 , \38489 , \38490 , \38491 , \38492 ,
         \38493 , \38494 , \38495 , \38496 , \38497 , \38498 , \38499 , \38500 , \38501 , \38502 ,
         \38503 , \38504 , \38505 , \38506 , \38507 , \38508 , \38509 , \38510 , \38511 , \38512 ,
         \38513 , \38514 , \38515 , \38516 , \38517 , \38518 , \38519 , \38520 , \38521 , \38522 ,
         \38523 , \38524 , \38525 , \38526 , \38527 , \38528 , \38529 , \38530 , \38531 , \38532 ,
         \38533 , \38534 , \38535 , \38536 , \38537 , \38538 , \38539 , \38540 , \38541 , \38542 ,
         \38543 , \38544 , \38545 , \38546 , \38547 , \38548 , \38549 , \38550 , \38551 , \38552 ,
         \38553 , \38554 , \38555 , \38556 , \38557 , \38558 , \38559 , \38560 , \38561 , \38562 ,
         \38563 , \38564 , \38565 , \38566 , \38567 , \38568 , \38569 , \38570 , \38571 , \38572 ,
         \38573 , \38574 , \38575 , \38576 , \38577 , \38578 , \38579 , \38580 , \38581 , \38582 ,
         \38583 , \38584 , \38585 , \38586 , \38587 , \38588 , \38589 , \38590 , \38591 , \38592 ,
         \38593 , \38594 , \38595 , \38596 , \38597 , \38598 , \38599 , \38600 , \38601 , \38602 ,
         \38603 , \38604 , \38605 , \38606 , \38607 , \38608 , \38609 , \38610 , \38611 , \38612 ,
         \38613 , \38614 , \38615 , \38616 , \38617 , \38618 , \38619 , \38620 , \38621 , \38622 ,
         \38623 , \38624 , \38625 , \38626 , \38627 , \38628 , \38629 , \38630 , \38631 , \38632 ,
         \38633 , \38634 , \38635 , \38636 , \38637 , \38638 , \38639 , \38640 , \38641 , \38642 ,
         \38643 , \38644 , \38645 , \38646 , \38647 , \38648 , \38649 , \38650 , \38651 , \38652 ,
         \38653 , \38654 , \38655 , \38656 , \38657 , \38658 , \38659 , \38660 , \38661 , \38662 ,
         \38663 , \38664 , \38665 , \38666 , \38667 , \38668 , \38669 , \38670 , \38671 , \38672 ,
         \38673 , \38674 , \38675 , \38676 , \38677 , \38678 , \38679 , \38680 , \38681 , \38682 ,
         \38683 , \38684 , \38685 , \38686 , \38687 , \38688 , \38689 , \38690 , \38691 , \38692 ,
         \38693 , \38694 , \38695 , \38696 , \38697 , \38698 , \38699 , \38700 , \38701 , \38702 ,
         \38703 , \38704 , \38705 , \38706 , \38707 , \38708 , \38709 , \38710 , \38711 , \38712 ,
         \38713 , \38714 , \38715 , \38716 , \38717 , \38718 , \38719 , \38720 , \38721 , \38722 ,
         \38723 , \38724 , \38725 , \38726 , \38727 , \38728 , \38729 , \38730 , \38731 , \38732 ,
         \38733 , \38734 , \38735 , \38736 , \38737 , \38738 , \38739 , \38740 , \38741 , \38742 ,
         \38743 , \38744 , \38745 , \38746 , \38747 , \38748 , \38749 , \38750 , \38751 , \38752 ,
         \38753 , \38754 , \38755 , \38756 , \38757 , \38758 , \38759 , \38760 , \38761 , \38762 ,
         \38763 , \38764 , \38765 , \38766 , \38767 , \38768 , \38769 , \38770 , \38771 , \38772 ,
         \38773 , \38774 , \38775 , \38776 , \38777 , \38778 , \38779 , \38780 , \38781 , \38782 ,
         \38783 , \38784 , \38785 , \38786 , \38787 , \38788 , \38789 , \38790 , \38791 , \38792 ,
         \38793 , \38794 , \38795 , \38796 , \38797 , \38798 , \38799 , \38800 , \38801 , \38802 ,
         \38803 , \38804 , \38805 , \38806 , \38807 , \38808 , \38809 , \38810 , \38811 , \38812 ,
         \38813 , \38814 , \38815 , \38816 , \38817 , \38818 , \38819 , \38820 , \38821 , \38822 ,
         \38823 , \38824 , \38825 , \38826 , \38827 , \38828 , \38829 , \38830 , \38831 , \38832 ,
         \38833 , \38834 , \38835 , \38836 , \38837 , \38838 , \38839 , \38840 , \38841 , \38842 ,
         \38843 , \38844 , \38845 , \38846 , \38847 , \38848 , \38849 , \38850 , \38851 , \38852 ,
         \38853 , \38854 , \38855 , \38856 , \38857 , \38858 , \38859 , \38860 , \38861 , \38862 ,
         \38863 , \38864 , \38865 , \38866 , \38867 , \38868 , \38869 , \38870 , \38871 , \38872 ,
         \38873 , \38874 , \38875 , \38876 , \38877 , \38878 , \38879 , \38880 , \38881 , \38882 ,
         \38883 , \38884 , \38885 , \38886 , \38887 , \38888 , \38889 , \38890 , \38891 , \38892 ,
         \38893 , \38894 , \38895 , \38896 , \38897 , \38898 , \38899 , \38900 , \38901 , \38902 ,
         \38903 , \38904 , \38905 , \38906 , \38907 , \38908 , \38909 , \38910 , \38911 , \38912 ,
         \38913 , \38914 , \38915 , \38916 , \38917 , \38918 , \38919 , \38920 , \38921 , \38922 ,
         \38923 , \38924 , \38925 , \38926 , \38927 , \38928 , \38929 , \38930 , \38931 , \38932 ,
         \38933 , \38934 , \38935 , \38936 , \38937 , \38938 , \38939 , \38940 , \38941 , \38942 ,
         \38943 , \38944 , \38945 , \38946 , \38947 , \38948 , \38949 , \38950 , \38951 , \38952 ,
         \38953 , \38954 , \38955 , \38956 , \38957 , \38958 , \38959 , \38960 , \38961 , \38962 ,
         \38963 , \38964 , \38965 , \38966 , \38967 , \38968 , \38969 , \38970 , \38971 , \38972 ,
         \38973 , \38974 , \38975 , \38976 , \38977 , \38978 , \38979 , \38980 , \38981 , \38982 ,
         \38983 , \38984 , \38985 , \38986 , \38987 , \38988 , \38989 , \38990 , \38991 , \38992 ,
         \38993 , \38994 , \38995 , \38996 , \38997 , \38998 , \38999 , \39000 , \39001 , \39002 ,
         \39003 , \39004 , \39005 , \39006 , \39007 , \39008 , \39009 , \39010 , \39011 , \39012 ,
         \39013 , \39014 , \39015 , \39016 , \39017 , \39018 , \39019 , \39020 , \39021 , \39022 ,
         \39023 , \39024 , \39025 , \39026 , \39027 , \39028 , \39029 , \39030 , \39031 , \39032 ,
         \39033 , \39034 , \39035 , \39036 , \39037 , \39038 , \39039 , \39040 , \39041 , \39042 ,
         \39043 , \39044 , \39045 , \39046 , \39047 , \39048 , \39049 , \39050 , \39051 , \39052 ,
         \39053 , \39054 , \39055 , \39056 , \39057 , \39058 , \39059 , \39060 , \39061 , \39062 ,
         \39063 , \39064 , \39065 , \39066 , \39067 , \39068 , \39069 , \39070 , \39071 , \39072 ,
         \39073 , \39074 , \39075 , \39076 , \39077 , \39078 , \39079 , \39080 , \39081 , \39082 ,
         \39083 , \39084 , \39085 , \39086 , \39087 , \39088 , \39089 , \39090 , \39091 , \39092 ,
         \39093 , \39094 , \39095 , \39096 , \39097 , \39098 , \39099 , \39100 , \39101 , \39102 ,
         \39103 , \39104 , \39105 , \39106 , \39107 , \39108 , \39109 , \39110 , \39111 , \39112 ,
         \39113 , \39114 , \39115 , \39116 , \39117 , \39118 , \39119 , \39120 , \39121 , \39122 ,
         \39123 , \39124 , \39125 , \39126 , \39127 , \39128 , \39129 , \39130 , \39131 , \39132 ,
         \39133 , \39134 , \39135 , \39136 , \39137 , \39138 , \39139 , \39140 , \39141 , \39142 ,
         \39143 , \39144 , \39145 , \39146 , \39147 , \39148 , \39149 , \39150 , \39151 , \39152 ,
         \39153 , \39154 , \39155 , \39156 , \39157 , \39158 , \39159 , \39160 , \39161 , \39162 ,
         \39163 , \39164 , \39165 , \39166 , \39167 , \39168 , \39169 , \39170 , \39171 , \39172 ,
         \39173 , \39174 , \39175 , \39176 , \39177 , \39178 , \39179 , \39180 , \39181 , \39182 ,
         \39183 , \39184 , \39185 , \39186 , \39187 , \39188 , \39189 , \39190 , \39191 , \39192 ,
         \39193 , \39194 , \39195 , \39196 , \39197 , \39198 , \39199 , \39200 , \39201 , \39202 ,
         \39203 , \39204 , \39205 , \39206 , \39207 , \39208 , \39209 , \39210 , \39211 , \39212 ,
         \39213 , \39214 , \39215 , \39216 , \39217 , \39218 , \39219 , \39220 , \39221 , \39222 ,
         \39223 , \39224 , \39225 , \39226 , \39227 , \39228 , \39229 , \39230 , \39231 , \39232 ,
         \39233 , \39234 , \39235 , \39236 , \39237 , \39238 , \39239 , \39240 , \39241 , \39242 ,
         \39243 , \39244 , \39245 , \39246 , \39247 , \39248 , \39249 , \39250 , \39251 , \39252 ,
         \39253 , \39254 , \39255 , \39256 , \39257 , \39258 , \39259 , \39260 , \39261 , \39262 ,
         \39263 , \39264 , \39265 , \39266 , \39267 , \39268 , \39269 , \39270 , \39271 , \39272 ,
         \39273 , \39274 , \39275 , \39276 , \39277 , \39278 , \39279 , \39280 , \39281 , \39282 ,
         \39283 , \39284 , \39285 , \39286 , \39287 , \39288 , \39289 , \39290 , \39291 , \39292 ,
         \39293 , \39294 , \39295 , \39296 , \39297 , \39298 , \39299 , \39300 , \39301 , \39302 ,
         \39303 , \39304 , \39305 , \39306 , \39307 , \39308 , \39309 , \39310 , \39311 , \39312 ,
         \39313 , \39314 , \39315 , \39316 , \39317 , \39318 , \39319 , \39320 , \39321 , \39322 ,
         \39323 , \39324 , \39325 , \39326 , \39327 , \39328 , \39329 , \39330 , \39331 , \39332 ,
         \39333 , \39334 , \39335 , \39336 , \39337 , \39338 , \39339 , \39340 , \39341 , \39342 ,
         \39343 , \39344 , \39345 , \39346 , \39347 , \39348 , \39349 , \39350 , \39351 , \39352 ,
         \39353 , \39354 , \39355 , \39356 , \39357 , \39358 , \39359 , \39360 , \39361 , \39362 ,
         \39363 , \39364 , \39365 , \39366 , \39367 , \39368 , \39369 , \39370 , \39371 , \39372 ,
         \39373 , \39374 , \39375 , \39376 , \39377 , \39378 , \39379 , \39380 , \39381 , \39382 ,
         \39383 , \39384 , \39385 , \39386 , \39387 , \39388 , \39389 , \39390 , \39391 , \39392 ,
         \39393 , \39394 , \39395 , \39396 , \39397 , \39398 , \39399 , \39400 , \39401 , \39402 ,
         \39403 , \39404 , \39405 , \39406 , \39407 , \39408 , \39409 , \39410 , \39411 , \39412 ,
         \39413 , \39414 , \39415 , \39416 , \39417 , \39418 , \39419 , \39420 , \39421 , \39422 ,
         \39423 , \39424 , \39425 , \39426 , \39427 , \39428 , \39429 , \39430 , \39431 , \39432 ,
         \39433 , \39434 , \39435 , \39436 , \39437 , \39438 , \39439 , \39440 , \39441 , \39442 ,
         \39443 , \39444 , \39445 , \39446 , \39447 , \39448 , \39449 , \39450 , \39451 , \39452 ,
         \39453 , \39454 , \39455 , \39456 , \39457 , \39458 , \39459 , \39460 , \39461 , \39462 ,
         \39463 , \39464 , \39465 , \39466 , \39467 , \39468 , \39469 , \39470 , \39471 , \39472 ,
         \39473 , \39474 , \39475 , \39476 , \39477 , \39478 , \39479 , \39480 , \39481 , \39482 ,
         \39483 , \39484 , \39485 , \39486 , \39487 , \39488 , \39489 , \39490 , \39491 , \39492 ,
         \39493 , \39494 , \39495 , \39496 , \39497 , \39498 , \39499 , \39500 , \39501 , \39502 ,
         \39503 , \39504 , \39505 , \39506 , \39507 , \39508 , \39509 , \39510 , \39511 , \39512 ,
         \39513 , \39514 , \39515 , \39516 , \39517 , \39518 , \39519 , \39520 , \39521 , \39522 ,
         \39523 , \39524 , \39525 , \39526 , \39527 , \39528 , \39529 , \39530 , \39531 , \39532 ,
         \39533 , \39534 , \39535 , \39536 , \39537 , \39538 , \39539 , \39540 , \39541 , \39542 ,
         \39543 , \39544 , \39545 , \39546 , \39547 , \39548 , \39549 , \39550 , \39551 , \39552 ,
         \39553 , \39554 , \39555 , \39556 , \39557 , \39558 , \39559 , \39560 , \39561 , \39562 ,
         \39563 , \39564 , \39565 , \39566 , \39567 , \39568 , \39569 , \39570 , \39571 , \39572 ,
         \39573 , \39574 , \39575 , \39576 , \39577 , \39578 , \39579 , \39580 , \39581 , \39582 ,
         \39583 , \39584 , \39585 , \39586 , \39587 , \39588 , \39589 , \39590 , \39591 , \39592 ,
         \39593 , \39594 , \39595 , \39596 , \39597 , \39598 , \39599 , \39600 , \39601 , \39602 ,
         \39603 , \39604 , \39605 , \39606 , \39607 , \39608 , \39609 , \39610 , \39611 , \39612 ,
         \39613 , \39614 , \39615 , \39616 , \39617 , \39618 , \39619 , \39620 , \39621 , \39622 ,
         \39623 , \39624 , \39625 , \39626 , \39627 , \39628 , \39629 , \39630 , \39631 , \39632 ,
         \39633 , \39634 , \39635 , \39636 , \39637 , \39638 , \39639 , \39640 , \39641 , \39642 ,
         \39643 , \39644 , \39645 , \39646 , \39647 , \39648 , \39649 , \39650 , \39651 , \39652 ,
         \39653 , \39654 , \39655 , \39656 , \39657 , \39658 , \39659 , \39660 , \39661 , \39662 ,
         \39663 , \39664 , \39665 , \39666 , \39667 , \39668 , \39669 , \39670 , \39671 , \39672 ,
         \39673 , \39674 , \39675 , \39676 , \39677 , \39678 , \39679 , \39680 , \39681 , \39682 ,
         \39683 , \39684 , \39685 , \39686 , \39687 , \39688 , \39689 , \39690 , \39691 , \39692 ,
         \39693 , \39694 , \39695 , \39696 , \39697 , \39698 , \39699 , \39700 , \39701 , \39702 ,
         \39703 , \39704 , \39705 , \39706 , \39707 , \39708 , \39709 , \39710 , \39711 , \39712 ,
         \39713 , \39714 , \39715 , \39716 , \39717 , \39718 , \39719 , \39720 , \39721 , \39722 ,
         \39723 , \39724 , \39725 , \39726 , \39727 , \39728 , \39729 , \39730 , \39731 , \39732 ,
         \39733 , \39734 , \39735 , \39736 , \39737 , \39738 , \39739 , \39740 , \39741 , \39742 ,
         \39743 , \39744 , \39745 , \39746 , \39747 , \39748 , \39749 , \39750 , \39751 , \39752 ,
         \39753 , \39754 , \39755 , \39756 , \39757 , \39758 , \39759 , \39760 , \39761 , \39762 ,
         \39763 , \39764 , \39765 , \39766 , \39767 , \39768 , \39769 , \39770 , \39771 , \39772 ,
         \39773 , \39774 , \39775 , \39776 , \39777 , \39778 , \39779 , \39780 , \39781 , \39782 ,
         \39783 , \39784 , \39785 , \39786 , \39787 , \39788 , \39789 , \39790 , \39791 , \39792 ,
         \39793 , \39794 , \39795 , \39796 , \39797 , \39798 , \39799 , \39800 , \39801 , \39802 ,
         \39803 , \39804 , \39805 , \39806 , \39807 , \39808 , \39809 , \39810 , \39811 , \39812 ,
         \39813 , \39814 , \39815 , \39816 , \39817 , \39818 , \39819 , \39820 , \39821 , \39822 ,
         \39823 , \39824 , \39825 , \39826 , \39827 , \39828 , \39829 , \39830 , \39831 , \39832 ,
         \39833 , \39834 , \39835 , \39836 , \39837 , \39838 , \39839 , \39840 , \39841 , \39842 ,
         \39843 , \39844 , \39845 , \39846 , \39847 , \39848 , \39849 , \39850 , \39851 , \39852 ,
         \39853 , \39854 , \39855 , \39856 , \39857 , \39858 , \39859 , \39860 , \39861 , \39862 ,
         \39863 , \39864 , \39865 , \39866 , \39867 , \39868 , \39869 , \39870 , \39871 , \39872 ,
         \39873 , \39874 , \39875 , \39876 , \39877 , \39878 , \39879 , \39880 , \39881 , \39882 ,
         \39883 , \39884 , \39885 , \39886 , \39887 , \39888 , \39889 , \39890 , \39891 , \39892 ,
         \39893 , \39894 , \39895 , \39896 , \39897 , \39898 , \39899 , \39900 , \39901 , \39902 ,
         \39903 , \39904 , \39905 , \39906 , \39907 , \39908 , \39909 , \39910 , \39911 , \39912 ,
         \39913 , \39914 , \39915 , \39916 , \39917 , \39918 , \39919 , \39920 , \39921 , \39922 ,
         \39923 , \39924 , \39925 , \39926 , \39927 , \39928 , \39929 , \39930 , \39931 , \39932 ,
         \39933 , \39934 , \39935 , \39936 , \39937 , \39938 , \39939 , \39940 , \39941 , \39942 ,
         \39943 , \39944 , \39945 , \39946 , \39947 , \39948 , \39949 , \39950 , \39951 , \39952 ,
         \39953 , \39954 , \39955 , \39956 , \39957 , \39958 , \39959 , \39960 , \39961 , \39962 ,
         \39963 , \39964 , \39965 , \39966 , \39967 , \39968 , \39969 , \39970 , \39971 , \39972 ,
         \39973 , \39974 , \39975 , \39976 , \39977 , \39978 , \39979 , \39980 , \39981 , \39982 ,
         \39983 , \39984 , \39985 , \39986 , \39987 , \39988 , \39989 , \39990 , \39991 , \39992 ,
         \39993 , \39994 , \39995 , \39996 , \39997 , \39998 , \39999 , \40000 , \40001 , \40002 ,
         \40003 , \40004 , \40005 , \40006 , \40007 , \40008 , \40009 , \40010 , \40011 , \40012 ,
         \40013 , \40014 , \40015 , \40016 , \40017 , \40018 , \40019 , \40020 , \40021 , \40022 ,
         \40023 , \40024 , \40025 , \40026 , \40027 , \40028 , \40029 , \40030 , \40031 , \40032 ,
         \40033 , \40034 , \40035 , \40036 , \40037 , \40038 , \40039 , \40040 , \40041 , \40042 ,
         \40043 , \40044 , \40045 , \40046 , \40047 , \40048 , \40049 , \40050 , \40051 , \40052 ,
         \40053 , \40054 , \40055 , \40056 , \40057 , \40058 , \40059 , \40060 , \40061 , \40062 ,
         \40063 , \40064 , \40065 , \40066 , \40067 , \40068 , \40069 , \40070 , \40071 , \40072 ,
         \40073 , \40074 , \40075 , \40076 , \40077 , \40078 , \40079 , \40080 , \40081 , \40082 ,
         \40083 , \40084 , \40085 , \40086 , \40087 , \40088 , \40089 , \40090 , \40091 , \40092 ,
         \40093 , \40094 , \40095 , \40096 , \40097 , \40098 , \40099 , \40100 , \40101 , \40102 ,
         \40103 , \40104 , \40105 , \40106 , \40107 , \40108 , \40109 , \40110 , \40111 , \40112 ,
         \40113 , \40114 , \40115 , \40116 , \40117 , \40118 , \40119 , \40120 , \40121 , \40122 ,
         \40123 , \40124 , \40125 , \40126 , \40127 , \40128 , \40129 , \40130 , \40131 , \40132 ,
         \40133 , \40134 , \40135 , \40136 , \40137 , \40138 , \40139 , \40140 , \40141 , \40142 ,
         \40143 , \40144 , \40145 , \40146 , \40147 , \40148 , \40149 , \40150 , \40151 , \40152 ,
         \40153 , \40154 , \40155 , \40156 , \40157 , \40158 , \40159 , \40160 , \40161 , \40162 ,
         \40163 , \40164 , \40165 , \40166 , \40167 , \40168 , \40169 , \40170 , \40171 , \40172 ,
         \40173 , \40174 , \40175 , \40176 , \40177 , \40178 , \40179 , \40180 , \40181 , \40182 ,
         \40183 , \40184 , \40185 , \40186 , \40187 , \40188 , \40189 , \40190 , \40191 , \40192 ,
         \40193 , \40194 , \40195 , \40196 , \40197 , \40198 , \40199 , \40200 , \40201 , \40202 ,
         \40203 , \40204 , \40205 , \40206 , \40207 , \40208 , \40209 , \40210 , \40211 , \40212 ,
         \40213 , \40214 , \40215 , \40216 , \40217 , \40218 , \40219 , \40220 , \40221 , \40222 ,
         \40223 , \40224 , \40225 , \40226 , \40227 , \40228 , \40229 , \40230 , \40231 , \40232 ,
         \40233 , \40234 , \40235 , \40236 , \40237 , \40238 , \40239 , \40240 , \40241 , \40242 ,
         \40243 , \40244 , \40245 , \40246 , \40247 , \40248 , \40249 , \40250 , \40251 , \40252 ,
         \40253 , \40254 , \40255 , \40256 , \40257 , \40258 , \40259 , \40260 , \40261 , \40262 ,
         \40263 , \40264 , \40265 , \40266 , \40267 , \40268 , \40269 , \40270 , \40271 , \40272 ,
         \40273 , \40274 , \40275 , \40276 , \40277 , \40278 , \40279 , \40280 , \40281 , \40282 ,
         \40283 , \40284 , \40285 , \40286 , \40287 , \40288 , \40289 , \40290 , \40291 , \40292 ,
         \40293 , \40294 , \40295 , \40296 , \40297 , \40298 , \40299 , \40300 , \40301 , \40302 ,
         \40303 , \40304 , \40305 , \40306 , \40307 , \40308 , \40309 , \40310 , \40311 , \40312 ,
         \40313 , \40314 , \40315 , \40316 , \40317 , \40318 , \40319 , \40320 , \40321 , \40322 ,
         \40323 , \40324 , \40325 , \40326 , \40327 , \40328 , \40329 , \40330 , \40331 , \40332 ,
         \40333 , \40334 , \40335 , \40336 , \40337 , \40338 , \40339 , \40340 , \40341 , \40342 ,
         \40343 , \40344 , \40345 , \40346 , \40347 , \40348 , \40349 , \40350 , \40351 , \40352 ,
         \40353 , \40354 , \40355 , \40356 , \40357 , \40358 , \40359 , \40360 , \40361 , \40362 ,
         \40363 , \40364 , \40365 , \40366 , \40367 , \40368 , \40369 , \40370 , \40371 , \40372 ,
         \40373 , \40374 , \40375 , \40376 , \40377 , \40378 , \40379 , \40380 , \40381 , \40382 ,
         \40383 , \40384 , \40385 , \40386 , \40387 , \40388 , \40389 , \40390 , \40391 , \40392 ,
         \40393 , \40394 , \40395 , \40396 , \40397 , \40398 , \40399 , \40400 , \40401 , \40402 ,
         \40403 , \40404 , \40405 , \40406 , \40407 , \40408 , \40409 , \40410 , \40411 , \40412 ,
         \40413 , \40414 , \40415 , \40416 , \40417 , \40418 , \40419 , \40420 , \40421 , \40422 ,
         \40423 , \40424 , \40425 , \40426 , \40427 , \40428 , \40429 , \40430 , \40431 , \40432 ,
         \40433 , \40434 , \40435 , \40436 , \40437 , \40438 , \40439 , \40440 , \40441 , \40442 ,
         \40443 , \40444 , \40445 , \40446 , \40447 , \40448 , \40449 , \40450 , \40451 , \40452 ,
         \40453 , \40454 , \40455 , \40456 , \40457 , \40458 , \40459 , \40460 , \40461 , \40462 ,
         \40463 , \40464 , \40465 , \40466 , \40467 , \40468 , \40469 , \40470 , \40471 , \40472 ,
         \40473 , \40474 , \40475 , \40476 , \40477 , \40478 , \40479 , \40480 , \40481 , \40482 ,
         \40483 , \40484 , \40485 , \40486 , \40487 , \40488 , \40489 , \40490 , \40491 , \40492 ,
         \40493 , \40494 , \40495 , \40496 , \40497 , \40498 , \40499 , \40500 , \40501 , \40502 ,
         \40503 , \40504 , \40505 , \40506 , \40507 , \40508 , \40509 , \40510 , \40511 , \40512 ,
         \40513 , \40514 , \40515 , \40516 , \40517 , \40518 , \40519 , \40520 , \40521 , \40522 ,
         \40523 , \40524 , \40525 , \40526 , \40527 , \40528 , \40529 , \40530 , \40531 , \40532 ,
         \40533 , \40534 , \40535 , \40536 , \40537 , \40538 , \40539 , \40540 , \40541 , \40542 ,
         \40543 , \40544 , \40545 , \40546 , \40547 , \40548 , \40549 , \40550 , \40551 , \40552 ,
         \40553 , \40554 , \40555 , \40556 , \40557 , \40558 , \40559 , \40560 , \40561 , \40562 ,
         \40563 , \40564 , \40565 , \40566 , \40567 , \40568 , \40569 , \40570 , \40571 , \40572 ,
         \40573 , \40574 , \40575 , \40576 , \40577 , \40578 , \40579 , \40580 , \40581 , \40582 ,
         \40583 , \40584 , \40585 , \40586 , \40587 , \40588 , \40589 , \40590 , \40591 , \40592 ,
         \40593 , \40594 , \40595 , \40596 , \40597 , \40598 , \40599 , \40600 , \40601 , \40602 ,
         \40603 , \40604 , \40605 , \40606 , \40607 , \40608 , \40609 , \40610 , \40611 , \40612 ,
         \40613 , \40614 , \40615 , \40616 , \40617 , \40618 , \40619 , \40620 , \40621 , \40622 ,
         \40623 , \40624 , \40625 , \40626 , \40627 , \40628 , \40629 , \40630 , \40631 , \40632 ,
         \40633 , \40634 , \40635 , \40636 , \40637 , \40638 , \40639 , \40640 , \40641 , \40642 ,
         \40643 , \40644 , \40645 , \40646 , \40647 , \40648 , \40649 , \40650 , \40651 , \40652 ,
         \40653 , \40654 , \40655 , \40656 , \40657 , \40658 , \40659 , \40660 , \40661 , \40662 ,
         \40663 , \40664 , \40665 , \40666 , \40667 , \40668 , \40669 , \40670 , \40671 , \40672 ,
         \40673 , \40674 , \40675 , \40676 , \40677 , \40678 , \40679 , \40680 , \40681 , \40682 ,
         \40683 , \40684 , \40685 , \40686 , \40687 , \40688 , \40689 , \40690 , \40691 , \40692 ,
         \40693 , \40694 , \40695 , \40696 , \40697 , \40698 , \40699 , \40700 , \40701 , \40702 ,
         \40703 , \40704 , \40705 , \40706 , \40707 , \40708 , \40709 , \40710 , \40711 , \40712 ,
         \40713 , \40714 , \40715 , \40716 , \40717 , \40718 , \40719 , \40720 , \40721 , \40722 ,
         \40723 , \40724 , \40725 , \40726 , \40727 , \40728 , \40729 , \40730 , \40731 , \40732 ,
         \40733 , \40734 , \40735 , \40736 , \40737 , \40738 , \40739 , \40740 , \40741 , \40742 ,
         \40743 , \40744 , \40745 , \40746 , \40747 , \40748 , \40749 , \40750 , \40751 , \40752 ,
         \40753 , \40754 , \40755 , \40756 , \40757 , \40758 , \40759 , \40760 , \40761 , \40762 ,
         \40763 , \40764 , \40765 , \40766 , \40767 , \40768 , \40769 , \40770 , \40771 , \40772 ,
         \40773 , \40774 , \40775 , \40776 , \40777 , \40778 , \40779 , \40780 , \40781 , \40782 ,
         \40783 , \40784 , \40785 , \40786 , \40787 , \40788 , \40789 , \40790 , \40791 , \40792 ,
         \40793 , \40794 , \40795 , \40796 , \40797 , \40798 , \40799 , \40800 , \40801 , \40802 ,
         \40803 , \40804 , \40805 , \40806 , \40807 , \40808 , \40809 , \40810 , \40811 , \40812 ,
         \40813 , \40814 , \40815 , \40816 , \40817 , \40818 , \40819 , \40820 , \40821 , \40822 ,
         \40823 , \40824 , \40825 , \40826 , \40827 , \40828 , \40829 , \40830 , \40831 , \40832 ,
         \40833 , \40834 , \40835 , \40836 , \40837 , \40838 , \40839 , \40840 , \40841 , \40842 ,
         \40843 , \40844 , \40845 , \40846 , \40847 , \40848 , \40849 , \40850 , \40851 , \40852 ,
         \40853 , \40854 , \40855 , \40856 , \40857 , \40858 , \40859 , \40860 , \40861 , \40862 ,
         \40863 , \40864 , \40865 , \40866 , \40867 , \40868 , \40869 , \40870 , \40871 , \40872 ,
         \40873 , \40874 , \40875 , \40876 , \40877 , \40878 , \40879 , \40880 , \40881 , \40882 ,
         \40883 , \40884 , \40885 , \40886 , \40887 , \40888 , \40889 , \40890 , \40891 , \40892 ,
         \40893 , \40894 , \40895 , \40896 , \40897 , \40898 , \40899 , \40900 , \40901 , \40902 ,
         \40903 , \40904 , \40905 , \40906 , \40907 , \40908 , \40909 , \40910 , \40911 , \40912 ,
         \40913 , \40914 , \40915 , \40916 , \40917 , \40918 , \40919 , \40920 , \40921 , \40922 ,
         \40923 , \40924 , \40925 , \40926 , \40927 , \40928 , \40929 , \40930 , \40931 , \40932 ,
         \40933 , \40934 , \40935 , \40936 , \40937 , \40938 , \40939 , \40940 , \40941 , \40942 ,
         \40943 , \40944 , \40945 , \40946 , \40947 , \40948 , \40949 , \40950 , \40951 , \40952 ,
         \40953 , \40954 , \40955 , \40956 , \40957 , \40958 , \40959 , \40960 , \40961 , \40962 ,
         \40963 , \40964 , \40965 , \40966 , \40967 , \40968 , \40969 , \40970 , \40971 , \40972 ,
         \40973 , \40974 , \40975 , \40976 , \40977 , \40978 , \40979 , \40980 , \40981 , \40982 ,
         \40983 , \40984 , \40985 , \40986 , \40987 , \40988 , \40989 , \40990 , \40991 , \40992 ,
         \40993 , \40994 , \40995 , \40996 , \40997 , \40998 , \40999 , \41000 , \41001 , \41002 ,
         \41003 , \41004 , \41005 , \41006 , \41007 , \41008 , \41009 , \41010 , \41011 , \41012 ,
         \41013 , \41014 , \41015 , \41016 , \41017 , \41018 , \41019 , \41020 , \41021 , \41022 ,
         \41023 , \41024 , \41025 , \41026 , \41027 , \41028 , \41029 , \41030 , \41031 , \41032 ,
         \41033 , \41034 , \41035 , \41036 , \41037 , \41038 , \41039 , \41040 , \41041 , \41042 ,
         \41043 , \41044 , \41045 , \41046 , \41047 , \41048 , \41049 , \41050 , \41051 , \41052 ,
         \41053 , \41054 , \41055 , \41056 , \41057 , \41058 , \41059 , \41060 , \41061 , \41062 ,
         \41063 , \41064 , \41065 , \41066 , \41067 , \41068 , \41069 , \41070 , \41071 , \41072 ,
         \41073 , \41074 , \41075 , \41076 , \41077 , \41078 , \41079 , \41080 , \41081 , \41082 ,
         \41083 , \41084 , \41085 , \41086 , \41087 , \41088 , \41089 , \41090 , \41091 , \41092 ,
         \41093 , \41094 , \41095 , \41096 , \41097 , \41098 , \41099 , \41100 , \41101 , \41102 ,
         \41103 , \41104 , \41105 , \41106 , \41107 , \41108 , \41109 , \41110 , \41111 , \41112 ,
         \41113 , \41114 , \41115 , \41116 , \41117 , \41118 , \41119 , \41120 , \41121 , \41122 ,
         \41123 , \41124 , \41125 , \41126 , \41127 , \41128 , \41129 , \41130 , \41131 , \41132 ,
         \41133 , \41134 , \41135 , \41136 , \41137 , \41138 , \41139 , \41140 , \41141 , \41142 ,
         \41143 , \41144 , \41145 , \41146 , \41147 , \41148 , \41149 , \41150 , \41151 , \41152 ,
         \41153 , \41154 , \41155 , \41156 , \41157 , \41158 , \41159 , \41160 , \41161 , \41162 ,
         \41163 , \41164 , \41165 , \41166 , \41167 , \41168 , \41169 , \41170 , \41171 , \41172 ,
         \41173 , \41174 , \41175 , \41176 , \41177 , \41178 , \41179 , \41180 , \41181 , \41182 ,
         \41183 , \41184 , \41185 , \41186 , \41187 , \41188 , \41189 , \41190 , \41191 , \41192 ,
         \41193 , \41194 , \41195 , \41196 , \41197 , \41198 , \41199 , \41200 , \41201 , \41202 ,
         \41203 , \41204 , \41205 , \41206 , \41207 , \41208 , \41209 , \41210 , \41211 , \41212 ,
         \41213 , \41214 , \41215 , \41216 , \41217 , \41218 , \41219 , \41220 , \41221 , \41222 ,
         \41223 , \41224 , \41225 , \41226 , \41227 , \41228 , \41229 , \41230 , \41231 , \41232 ,
         \41233 , \41234 , \41235 , \41236 , \41237 , \41238 , \41239 , \41240 , \41241 , \41242 ,
         \41243 , \41244 , \41245 , \41246 , \41247 , \41248 , \41249 , \41250 , \41251 , \41252 ,
         \41253 , \41254 , \41255 , \41256 , \41257 , \41258 , \41259 , \41260 , \41261 , \41262 ,
         \41263 , \41264 , \41265 , \41266 , \41267 , \41268 , \41269 , \41270 , \41271 , \41272 ,
         \41273 , \41274 , \41275 , \41276 , \41277 , \41278 , \41279 , \41280 , \41281 , \41282 ,
         \41283 , \41284 , \41285 , \41286 , \41287 , \41288 , \41289 , \41290 , \41291 , \41292 ,
         \41293 , \41294 , \41295 , \41296 , \41297 , \41298 , \41299 , \41300 , \41301 , \41302 ,
         \41303 , \41304 , \41305 , \41306 , \41307 , \41308 , \41309 , \41310 , \41311 , \41312 ,
         \41313 , \41314 , \41315 , \41316 , \41317 , \41318 , \41319 , \41320 , \41321 , \41322 ,
         \41323 , \41324 , \41325 , \41326 , \41327 , \41328 , \41329 , \41330 , \41331 , \41332 ,
         \41333 , \41334 , \41335 , \41336 , \41337 , \41338 , \41339 , \41340 , \41341 , \41342 ,
         \41343 , \41344 , \41345 , \41346 , \41347 , \41348 , \41349 , \41350 , \41351 , \41352 ,
         \41353 , \41354 , \41355 , \41356 , \41357 , \41358 , \41359 , \41360 , \41361 , \41362 ,
         \41363 , \41364 , \41365 , \41366 , \41367 , \41368 , \41369 , \41370 , \41371 , \41372 ,
         \41373 , \41374 , \41375 , \41376 , \41377 , \41378 , \41379 , \41380 , \41381 , \41382 ,
         \41383 , \41384 , \41385 , \41386 , \41387 , \41388 , \41389 , \41390 , \41391 , \41392 ,
         \41393 , \41394 , \41395 , \41396 , \41397 , \41398 , \41399 , \41400 , \41401 , \41402 ,
         \41403 , \41404 , \41405 , \41406 , \41407 , \41408 , \41409 , \41410 , \41411 , \41412 ,
         \41413 , \41414 , \41415 , \41416 , \41417 , \41418 , \41419 , \41420 , \41421 , \41422 ,
         \41423 , \41424 , \41425 , \41426 , \41427 , \41428 , \41429 , \41430 , \41431 , \41432 ,
         \41433 , \41434 , \41435 , \41436 , \41437 , \41438 , \41439 , \41440 , \41441 , \41442 ,
         \41443 , \41444 , \41445 , \41446 , \41447 , \41448 , \41449 , \41450 , \41451 , \41452 ,
         \41453 , \41454 , \41455 , \41456 , \41457 , \41458 , \41459 , \41460 , \41461 , \41462 ,
         \41463 , \41464 , \41465 , \41466 , \41467 , \41468 , \41469 , \41470 , \41471 , \41472 ,
         \41473 , \41474 , \41475 , \41476 , \41477 , \41478 , \41479 , \41480 , \41481 , \41482 ,
         \41483 , \41484 , \41485 , \41486 , \41487 , \41488 , \41489 , \41490 , \41491 , \41492 ,
         \41493 , \41494 , \41495 , \41496 , \41497 , \41498 , \41499 , \41500 , \41501 , \41502 ,
         \41503 , \41504 , \41505 , \41506 , \41507 , \41508 , \41509 , \41510 , \41511 , \41512 ,
         \41513 , \41514 , \41515 , \41516 , \41517 , \41518 , \41519 , \41520 , \41521 , \41522 ,
         \41523 , \41524 , \41525 , \41526 , \41527 , \41528 , \41529 , \41530 , \41531 , \41532 ,
         \41533 , \41534 , \41535 , \41536 , \41537 , \41538 , \41539 , \41540 , \41541 , \41542 ,
         \41543 , \41544 , \41545 , \41546 , \41547 , \41548 , \41549 , \41550 , \41551 , \41552 ,
         \41553 , \41554 , \41555 , \41556 , \41557 , \41558 , \41559 , \41560 , \41561 , \41562 ,
         \41563 , \41564 , \41565 , \41566 , \41567 , \41568 , \41569 , \41570 , \41571 , \41572 ,
         \41573 , \41574 , \41575 , \41576 , \41577 , \41578 , \41579 , \41580 , \41581 , \41582 ,
         \41583 , \41584 , \41585 , \41586 , \41587 , \41588 , \41589 , \41590 , \41591 , \41592 ,
         \41593 , \41594 , \41595 , \41596 , \41597 , \41598 , \41599 , \41600 , \41601 , \41602 ,
         \41603 , \41604 , \41605 , \41606 , \41607 , \41608 , \41609 , \41610 , \41611 , \41612 ,
         \41613 , \41614 , \41615 , \41616 , \41617 , \41618 , \41619 , \41620 , \41621 , \41622 ,
         \41623 , \41624 , \41625 , \41626 , \41627 , \41628 , \41629 , \41630 , \41631 , \41632 ,
         \41633 , \41634 , \41635 , \41636 , \41637 , \41638 , \41639 , \41640 , \41641 , \41642 ,
         \41643 , \41644 , \41645 , \41646 , \41647 , \41648 , \41649 , \41650 , \41651 , \41652 ,
         \41653 , \41654 , \41655 , \41656 , \41657 , \41658 , \41659 , \41660 , \41661 , \41662 ,
         \41663 , \41664 , \41665 , \41666 , \41667 , \41668 , \41669 , \41670 , \41671 , \41672 ,
         \41673 , \41674 , \41675 , \41676 , \41677 , \41678 , \41679 , \41680 , \41681 , \41682 ,
         \41683 , \41684 , \41685 , \41686 , \41687 , \41688 , \41689 , \41690 , \41691 , \41692 ,
         \41693 , \41694 , \41695 , \41696 , \41697 , \41698 , \41699 , \41700 , \41701 , \41702 ,
         \41703 , \41704 , \41705 , \41706 , \41707 , \41708 , \41709 , \41710 , \41711 , \41712 ,
         \41713 , \41714 , \41715 , \41716 , \41717 , \41718 , \41719 , \41720 , \41721 , \41722 ,
         \41723 , \41724 , \41725 , \41726 , \41727 , \41728 , \41729 , \41730 , \41731 , \41732 ,
         \41733 , \41734 , \41735 , \41736 , \41737 , \41738 , \41739 , \41740 , \41741 , \41742 ,
         \41743 , \41744 , \41745 , \41746 , \41747 , \41748 , \41749 , \41750 , \41751 , \41752 ,
         \41753 , \41754 , \41755 , \41756 , \41757 , \41758 , \41759 , \41760 , \41761 , \41762 ,
         \41763 , \41764 , \41765 , \41766 , \41767 , \41768 , \41769 , \41770 , \41771 , \41772 ,
         \41773 , \41774 , \41775 , \41776 , \41777 , \41778 , \41779 , \41780 , \41781 , \41782 ,
         \41783 , \41784 , \41785 , \41786 , \41787 , \41788 , \41789 , \41790 , \41791 , \41792 ,
         \41793 , \41794 , \41795 , \41796 , \41797 , \41798 , \41799 , \41800 , \41801 , \41802 ,
         \41803 , \41804 , \41805 , \41806 , \41807 , \41808 , \41809 , \41810 , \41811 , \41812 ,
         \41813 , \41814 , \41815 , \41816 , \41817 , \41818 , \41819 , \41820 , \41821 , \41822 ,
         \41823 , \41824 , \41825 , \41826 , \41827 , \41828 , \41829 , \41830 , \41831 , \41832 ,
         \41833 , \41834 , \41835 , \41836 , \41837 , \41838 , \41839 , \41840 , \41841 , \41842 ,
         \41843 , \41844 , \41845 , \41846 , \41847 , \41848 , \41849 , \41850 , \41851 , \41852 ,
         \41853 , \41854 , \41855 , \41856 , \41857 , \41858 , \41859 , \41860 , \41861 , \41862 ,
         \41863 , \41864 , \41865 , \41866 , \41867 , \41868 , \41869 , \41870 , \41871 , \41872 ,
         \41873 , \41874 , \41875 , \41876 , \41877 , \41878 , \41879 , \41880 , \41881 , \41882 ,
         \41883 , \41884 , \41885 , \41886 , \41887 , \41888 , \41889 , \41890 , \41891 , \41892 ,
         \41893 , \41894 , \41895 , \41896 , \41897 , \41898 , \41899 , \41900 , \41901 , \41902 ,
         \41903 , \41904 , \41905 , \41906 , \41907 , \41908 , \41909 , \41910 , \41911 , \41912 ,
         \41913 , \41914 , \41915 , \41916 , \41917 , \41918 , \41919 , \41920 , \41921 , \41922 ,
         \41923 , \41924 , \41925 , \41926 , \41927 , \41928 , \41929 , \41930 , \41931 , \41932 ,
         \41933_nGfa , \41934_nGf9 , \41935 , \41936 , \41937 , \41938 , \41939 , \41940 , \41941 , \41942 ,
         \41943 , \41944 , \41945 , \41946 , \41947 , \41948 , \41949 , \41950 , \41951 , \41952 ,
         \41953 , \41954 , \41955 , \41956 , \41957 , \41958 , \41959 , \41960 , \41961 , \41962 ,
         \41963 , \41964 , \41965 , \41966 , \41967 , \41968 , \41969 , \41970 , \41971 , \41972 ,
         \41973 , \41974 , \41975 , \41976 , \41977 , \41978 , \41979 , \41980 , \41981 , \41982 ,
         \41983 , \41984 , \41985 , \41986 , \41987 , \41988 , \41989 , \41990 , \41991 , \41992 ,
         \41993 , \41994 , \41995 , \41996 , \41997 , \41998 , \41999 , \42000 , \42001 , \42002 ,
         \42003 , \42004 , \42005 , \42006 , \42007 , \42008 , \42009 , \42010 , \42011 , \42012 ,
         \42013 , \42014 , \42015 , \42016 , \42017 , \42018 , \42019 , \42020 , \42021 , \42022 ,
         \42023 , \42024 , \42025 , \42026 , \42027 , \42028 , \42029 , \42030 , \42031 , \42032 ,
         \42033 , \42034 , \42035 , \42036 , \42037 , \42038 , \42039 , \42040 , \42041 , \42042 ,
         \42043 , \42044 , \42045 , \42046 , \42047 , \42048 , \42049 , \42050 , \42051 , \42052 ,
         \42053 , \42054 , \42055 , \42056 , \42057 , \42058 , \42059 , \42060 , \42061 , \42062 ,
         \42063 , \42064 , \42065 , \42066 , \42067 , \42068 , \42069 , \42070 , \42071 , \42072 ,
         \42073 , \42074 , \42075 , \42076 , \42077 , \42078 , \42079 , \42080 , \42081 , \42082 ,
         \42083 , \42084 , \42085 , \42086 , \42087 , \42088 , \42089 , \42090 , \42091 , \42092 ,
         \42093 , \42094 , \42095 , \42096 , \42097 , \42098 , \42099 , \42100 , \42101 , \42102 ,
         \42103 , \42104 , \42105 , \42106 , \42107 , \42108 , \42109 , \42110 , \42111 , \42112 ,
         \42113 , \42114 , \42115 , \42116 , \42117 , \42118 , \42119 , \42120 , \42121 , \42122 ,
         \42123 , \42124 , \42125 , \42126 , \42127 , \42128 , \42129 , \42130 , \42131 , \42132 ,
         \42133 , \42134 , \42135 , \42136 , \42137 , \42138 , \42139 , \42140 , \42141 , \42142 ,
         \42143 , \42144 , \42145 , \42146 , \42147 , \42148 , \42149 , \42150 , \42151 , \42152 ,
         \42153 , \42154 , \42155 , \42156 , \42157 , \42158 , \42159 , \42160 , \42161 , \42162 ,
         \42163 , \42164 , \42165 , \42166 , \42167 , \42168 , \42169 , \42170 , \42171 , \42172 ,
         \42173 , \42174 , \42175 , \42176 , \42177 , \42178 , \42179 , \42180 , \42181 , \42182 ,
         \42183 , \42184 , \42185 , \42186 , \42187 , \42188 , \42189 , \42190 , \42191 , \42192 ,
         \42193 , \42194 , \42195 , \42196 , \42197 , \42198 , \42199 , \42200 , \42201 , \42202 ,
         \42203 , \42204 , \42205 , \42206 , \42207 , \42208 , \42209 , \42210 , \42211 , \42212 ,
         \42213 , \42214 , \42215 , \42216 , \42217 , \42218 , \42219 , \42220 , \42221 , \42222 ,
         \42223 , \42224 , \42225 , \42226 , \42227 , \42228 , \42229 , \42230 , \42231 , \42232 ,
         \42233 , \42234 , \42235 , \42236 , \42237 , \42238 , \42239 , \42240 , \42241 , \42242 ,
         \42243 , \42244 , \42245 , \42246 , \42247 , \42248 , \42249 , \42250 , \42251 , \42252 ,
         \42253 , \42254 , \42255 , \42256 , \42257 , \42258 , \42259 , \42260 , \42261 , \42262 ,
         \42263 , \42264 , \42265 , \42266 , \42267 , \42268 , \42269 , \42270 , \42271 , \42272 ,
         \42273 , \42274 , \42275 , \42276 , \42277 , \42278 , \42279 , \42280 , \42281 , \42282 ,
         \42283 , \42284 , \42285 , \42286 , \42287 , \42288 , \42289 , \42290 , \42291 , \42292 ,
         \42293 , \42294 , \42295 , \42296 , \42297 , \42298 , \42299 , \42300 , \42301 , \42302 ,
         \42303 , \42304 , \42305 , \42306 , \42307 , \42308 , \42309 , \42310 , \42311 , \42312 ,
         \42313 , \42314 , \42315 , \42316 , \42317 , \42318 , \42319 , \42320 , \42321 , \42322 ,
         \42323 , \42324 , \42325 , \42326 , \42327 , \42328 , \42329 , \42330 , \42331 , \42332 ,
         \42333 , \42334 , \42335 , \42336 , \42337 , \42338 , \42339 , \42340 , \42341 , \42342 ,
         \42343 , \42344 , \42345 , \42346 , \42347 , \42348 , \42349 , \42350 , \42351 , \42352 ,
         \42353 , \42354 , \42355 , \42356 , \42357 , \42358 , \42359 , \42360 , \42361 , \42362 ,
         \42363 , \42364 , \42365 , \42366 , \42367 , \42368 , \42369 , \42370 , \42371 , \42372 ,
         \42373 , \42374 , \42375 , \42376 , \42377 , \42378 , \42379 , \42380 , \42381 , \42382 ,
         \42383 , \42384 , \42385 , \42386 , \42387 , \42388 , \42389 , \42390 , \42391 , \42392 ,
         \42393 , \42394 , \42395 , \42396 , \42397 , \42398 , \42399 , \42400 , \42401 , \42402 ,
         \42403 , \42404 , \42405 , \42406 , \42407 , \42408 , \42409 , \42410 , \42411 , \42412 ,
         \42413 , \42414 , \42415 , \42416 , \42417 , \42418 , \42419 , \42420 , \42421 , \42422 ,
         \42423 , \42424 , \42425 , \42426 , \42427 , \42428 , \42429 , \42430 , \42431 , \42432 ,
         \42433 , \42434 , \42435 , \42436 , \42437 , \42438 , \42439 , \42440 , \42441 , \42442 ,
         \42443 , \42444 , \42445 , \42446 , \42447 , \42448 , \42449 , \42450 , \42451 , \42452 ,
         \42453 , \42454 , \42455 , \42456 , \42457 , \42458 , \42459 , \42460 , \42461 , \42462 ,
         \42463 , \42464 , \42465 , \42466 , \42467 , \42468 , \42469 , \42470 , \42471 , \42472 ,
         \42473 , \42474 , \42475 , \42476 , \42477 , \42478 , \42479 , \42480 , \42481 , \42482 ,
         \42483 , \42484 , \42485 , \42486 , \42487 , \42488 , \42489 , \42490 , \42491 , \42492 ,
         \42493 , \42494 , \42495 , \42496 , \42497 , \42498 , \42499 , \42500 , \42501 , \42502 ,
         \42503 , \42504 , \42505 , \42506 , \42507 , \42508 , \42509 , \42510 , \42511 , \42512 ,
         \42513 , \42514 , \42515 , \42516 , \42517 , \42518 , \42519 , \42520 , \42521 , \42522 ,
         \42523 , \42524 , \42525 , \42526 , \42527 , \42528 , \42529 , \42530 , \42531 , \42532 ,
         \42533 , \42534 , \42535 , \42536 , \42537 , \42538 , \42539 , \42540 , \42541 , \42542 ,
         \42543 , \42544 , \42545 , \42546 , \42547 , \42548 , \42549 , \42550 , \42551 , \42552 ,
         \42553 , \42554 , \42555 , \42556 , \42557 , \42558 , \42559 , \42560 , \42561 , \42562 ,
         \42563 , \42564 , \42565 , \42566 , \42567 , \42568 , \42569 , \42570 , \42571 , \42572 ,
         \42573 , \42574 , \42575 , \42576 , \42577 , \42578 , \42579 , \42580 , \42581 , \42582 ,
         \42583 , \42584 , \42585 , \42586 , \42587 , \42588 , \42589 , \42590 , \42591 , \42592 ,
         \42593 , \42594 , \42595 , \42596 , \42597 , \42598 , \42599 , \42600 , \42601 , \42602 ,
         \42603 , \42604 , \42605 , \42606 , \42607 , \42608 , \42609 , \42610 , \42611 , \42612 ,
         \42613 , \42614 , \42615 , \42616 , \42617 , \42618 , \42619 , \42620 , \42621 , \42622 ,
         \42623 , \42624 , \42625 , \42626 , \42627 , \42628 , \42629 , \42630 , \42631 , \42632 ,
         \42633 , \42634 , \42635 , \42636 , \42637 , \42638 , \42639 , \42640 , \42641 , \42642 ,
         \42643 , \42644 , \42645 , \42646 , \42647 , \42648 , \42649 , \42650 , \42651 , \42652 ,
         \42653 , \42654 , \42655 , \42656 , \42657 , \42658 , \42659 , \42660 , \42661 , \42662 ,
         \42663 , \42664 , \42665 , \42666 , \42667 , \42668 , \42669 , \42670 , \42671 , \42672 ,
         \42673 , \42674 , \42675 , \42676 , \42677 , \42678 , \42679 , \42680 , \42681 , \42682 ,
         \42683 , \42684 , \42685 , \42686 , \42687 , \42688 , \42689 , \42690 , \42691 , \42692 ,
         \42693 , \42694 , \42695 , \42696 , \42697 , \42698 , \42699 , \42700 , \42701 , \42702 ,
         \42703 , \42704 , \42705 , \42706 , \42707 , \42708 , \42709 , \42710 , \42711 , \42712 ,
         \42713 , \42714 , \42715 , \42716 , \42717 , \42718 , \42719 , \42720 , \42721 , \42722 ,
         \42723 , \42724 , \42725 , \42726 , \42727 , \42728 , \42729 , \42730 , \42731 , \42732 ,
         \42733 , \42734 , \42735 , \42736 , \42737 , \42738 , \42739 , \42740 , \42741 , \42742 ,
         \42743 , \42744 , \42745 , \42746 , \42747 , \42748 , \42749 , \42750 , \42751 , \42752 ,
         \42753 , \42754 , \42755 , \42756 , \42757 , \42758 , \42759 , \42760 , \42761 , \42762 ,
         \42763 , \42764 , \42765 , \42766 , \42767 , \42768 , \42769 , \42770 , \42771 , \42772 ,
         \42773 , \42774 , \42775 , \42776 , \42777 , \42778 , \42779 , \42780 , \42781 , \42782 ,
         \42783 , \42784 , \42785 , \42786 , \42787 , \42788 , \42789 , \42790 , \42791 , \42792 ,
         \42793 , \42794 , \42795 , \42796 , \42797 , \42798 , \42799 , \42800 , \42801 , \42802 ,
         \42803 , \42804 , \42805 , \42806 , \42807 , \42808 , \42809 , \42810 , \42811 , \42812 ,
         \42813 , \42814 , \42815 , \42816 , \42817 , \42818 , \42819 , \42820 , \42821 , \42822 ,
         \42823 , \42824 , \42825 , \42826 , \42827 , \42828 , \42829 , \42830 , \42831 , \42832 ,
         \42833 , \42834 , \42835 , \42836 , \42837 , \42838 , \42839 , \42840 , \42841 , \42842 ,
         \42843 , \42844 , \42845 , \42846 , \42847 , \42848 , \42849 , \42850 , \42851 , \42852 ,
         \42853 , \42854 , \42855 , \42856 , \42857 , \42858 , \42859 , \42860 , \42861 , \42862 ,
         \42863 , \42864 , \42865 , \42866 , \42867 , \42868 , \42869 , \42870 , \42871 , \42872 ,
         \42873 , \42874 , \42875 , \42876 , \42877 , \42878 , \42879 , \42880 , \42881 , \42882 ,
         \42883 , \42884 , \42885 , \42886 , \42887 , \42888 , \42889 , \42890 , \42891 , \42892 ,
         \42893 , \42894 , \42895 , \42896 , \42897 , \42898 , \42899 , \42900 , \42901 , \42902 ,
         \42903 , \42904 , \42905 , \42906 , \42907 , \42908 , \42909 , \42910 , \42911 , \42912 ,
         \42913 , \42914 , \42915 , \42916 , \42917 , \42918 , \42919 , \42920 , \42921 , \42922 ,
         \42923 , \42924 , \42925 , \42926 , \42927 , \42928 , \42929 , \42930 , \42931 , \42932 ,
         \42933 , \42934 , \42935 , \42936 , \42937 , \42938 , \42939 , \42940 , \42941 , \42942 ,
         \42943 , \42944 , \42945 , \42946 , \42947 , \42948 , \42949 , \42950 , \42951 , \42952 ,
         \42953 , \42954 , \42955 , \42956 , \42957 , \42958 , \42959 , \42960 , \42961 , \42962 ,
         \42963 , \42964 , \42965 , \42966 , \42967 , \42968 , \42969 , \42970 , \42971 , \42972 ,
         \42973 , \42974 , \42975 , \42976 , \42977 , \42978 , \42979 , \42980 , \42981 , \42982 ,
         \42983 , \42984 , \42985 , \42986 , \42987 , \42988 , \42989 , \42990 , \42991 , \42992 ,
         \42993 , \42994 , \42995 , \42996 , \42997 , \42998 , \42999 , \43000 , \43001 , \43002 ,
         \43003 , \43004 , \43005 , \43006 , \43007 , \43008 , \43009 , \43010 , \43011 , \43012 ,
         \43013 , \43014 , \43015 , \43016 , \43017 , \43018 , \43019 , \43020 , \43021 , \43022 ,
         \43023 , \43024 , \43025 , \43026 , \43027 , \43028 , \43029 , \43030 , \43031 , \43032 ,
         \43033 , \43034 , \43035 , \43036 , \43037 , \43038 , \43039 , \43040 , \43041 , \43042 ,
         \43043 , \43044 , \43045 , \43046 , \43047 , \43048 , \43049 , \43050 , \43051 , \43052 ,
         \43053 , \43054 , \43055 , \43056 , \43057 , \43058 , \43059 , \43060 , \43061 , \43062 ,
         \43063 , \43064 , \43065 , \43066 , \43067 , \43068 , \43069 , \43070 , \43071 , \43072 ,
         \43073 , \43074 , \43075 , \43076 , \43077 , \43078 , \43079 , \43080 , \43081 , \43082 ,
         \43083 , \43084 , \43085 , \43086 , \43087 , \43088 , \43089 , \43090 , \43091 , \43092 ,
         \43093 , \43094 , \43095 , \43096 , \43097 , \43098 , \43099 , \43100 , \43101 , \43102 ,
         \43103 , \43104 , \43105 , \43106 , \43107 , \43108 , \43109 , \43110 , \43111 , \43112 ,
         \43113 , \43114 , \43115 , \43116 , \43117 , \43118 , \43119 , \43120 , \43121 , \43122 ,
         \43123 , \43124 , \43125 , \43126 , \43127 , \43128 , \43129 , \43130 , \43131 , \43132 ,
         \43133 , \43134 , \43135 , \43136 , \43137 , \43138 , \43139 , \43140 , \43141 , \43142 ,
         \43143 , \43144 , \43145 , \43146 , \43147 , \43148 , \43149 , \43150 , \43151 , \43152 ,
         \43153 , \43154 , \43155 , \43156 ;
buf \U$labajz4347 ( R_81_9fc6f08, \42287 );
buf \U$labajz4348 ( R_82_9fc5ea0, \42294 );
buf \U$labajz4349 ( R_83_90f04e0, \42309 );
buf \U$labajz4350 ( R_84_90effa0, \42317 );
buf \U$labajz4351 ( R_85_90e8ad0, \42325 );
buf \U$labajz4352 ( R_86_90e3e08, \42372 );
buf \U$labajz4353 ( R_87_90f1a88, \42380 );
buf \U$labajz4354 ( R_88_90e8638, \42391 );
buf \U$labajz4355 ( R_89_90f1200, \42399 );
buf \U$labajz4356 ( R_8a_90f12a8, \42405 );
buf \U$labajz4357 ( R_8b_90f0cc0, \42421 );
buf \U$labajz4358 ( R_8c_90ef088, \42437 );
buf \U$labajz4359 ( R_8d_90f1158, \42457 );
buf \U$labajz4360 ( R_8e_90e49d8, \42467 );
buf \U$labajz4361 ( R_8f_90e3eb0, \42473 );
buf \U$labajz4362 ( R_90_9fc69c8, \42485 );
buf \U$labajz4363 ( R_91_90e9c88, \42496 );
buf \U$labajz4364 ( R_92_90f0588, \42516 );
buf \U$labajz4365 ( R_93_90eacf0, \42521 );
buf \U$labajz4366 ( R_94_90ebb60, \42527 );
buf \U$labajz4367 ( R_95_90e66b8, \42533 );
buf \U$labajz4368 ( R_96_9fc6d10, \42535 );
buf \U$labajz4369 ( R_97_90ead98, \42542 );
buf \U$labajz4370 ( R_98_90e90b8, \42549 );
buf \U$labajz4371 ( R_99_90eb038, \42551 );
buf \U$labajz4372 ( R_9a_90e9d30, \42553 );
buf \U$labajz4373 ( R_9b_90e7bb8, \42559 );
buf \U$labajz4374 ( R_9c_9fc7b80, \42599 );
buf \U$labajz4375 ( R_9d_90ebd58, \42607 );
buf \U$labajz4376 ( R_9e_90e9a90, \42614 );
buf \U$labajz4377 ( R_9f_90efb08, \42633 );
buf \U$labajz4378 ( R_a0_90e6e98, \42643 );
buf \U$labajz4379 ( R_a1_90f0780, \42663 );
buf \U$labajz4380 ( R_a2_90e2da0, \42670 );
buf \U$labajz4381 ( R_a3_90f0240, \42677 );
buf \U$labajz4382 ( R_a4_9fc7ad8, \42685 );
buf \U$labajz4383 ( R_a5_9fc73a0, \42687 );
buf \U$labajz4384 ( R_a6_9fc6680, \42689 );
buf \U$labajz4385 ( R_a7_90e4f18, \42697 );
buf \U$labajz4386 ( R_a8_90e3388, \42703 );
buf \U$labajz4387 ( R_a9_9fc67d0, \42708 );
buf \U$labajz4388 ( R_aa_90f17e8, \42713 );
buf \U$labajz4389 ( R_ab_90e4888, \42722 );
buf \U$labajz4390 ( R_ac_90e9010, \42729 );
buf \U$labajz4391 ( R_ad_90eee90, \42735 );
buf \U$labajz4392 ( R_ae_90e53b0, \42761 );
buf \U$labajz4393 ( R_af_90ebc08, \42768 );
buf \U$labajz4394 ( R_b0_90e8440, \42785 );
buf \U$labajz4395 ( R_b1_90ea900, \42790 );
buf \U$labajz4396 ( R_b2_90e9400, \42795 );
buf \U$labajz4397 ( R_b3_9fc6bc0, \42802 );
buf \U$labajz4398 ( R_b4_90e4690, \42807 );
buf \U$labajz4399 ( R_b5_90e3778, \42812 );
buf \U$labajz4400 ( R_b6_90e9160, \42818 );
buf \U$labajz4401 ( R_b7_90e29b0, \42824 );
buf \U$labajz4402 ( R_b8_90e2278, \42826 );
buf \U$labajz4403 ( R_b9_9fc6a70, \42828 );
buf \U$labajz4404 ( R_ba_90ebf50, \42830 );
buf \U$labajz4405 ( R_bb_90f0e10, \42849 );
buf \U$labajz4406 ( R_bc_9fc7640, \42854 );
buf \U$labajz4407 ( R_bd_90f1dd0, \42859 );
buf \U$labajz4408 ( R_be_90f0630, \42861 );
buf \U$labajz4409 ( R_bf_90f0eb8, \42866 );
buf \U$labajz4410 ( R_c0_90e34d8, \42868 );
buf \U$labajz4411 ( R_c1_90e9f28, \42900 );
buf \U$labajz4412 ( R_c2_90f0d68, \42908 );
buf \U$labajz4413 ( R_c3_90ea7b0, \42914 );
buf \U$labajz4414 ( R_c4_9fc7448, \42920 );
buf \U$labajz4415 ( R_c5_90eb428, \42926 );
buf \U$labajz4416 ( R_c6_90e81a0, \42932 );
buf \U$labajz4417 ( R_c7_90f0a20, \42940 );
buf \U$labajz4418 ( R_c8_90efda8, \42947 );
buf \U$labajz4419 ( R_c9_90e2c50, \42953 );
buf \U$labajz4420 ( R_ca_90e88d8, \42961 );
buf \U$labajz4421 ( R_cb_9fc6530, \42966 );
buf \U$labajz4422 ( R_cc_90f06d8, \42968 );
buf \U$labajz4423 ( R_cd_90efa60, \42986 );
buf \U$labajz4424 ( R_ce_90e2b00, \42991 );
buf \U$labajz4425 ( R_cf_9fc6920, \43000 );
buf \U$labajz4426 ( R_d0_90f1f20, \43002 );
buf \U$labajz4427 ( R_d1_90e7678, \43004 );
buf \U$labajz4428 ( R_d2_90efd00, \43009 );
buf \U$labajz4429 ( R_d3_90e7e58, \43015 );
buf \U$labajz4430 ( R_d4_90e7d08, \43017 );
buf \U$labajz4431 ( R_d5_90eaa50, \43022 );
buf \U$labajz4432 ( R_d6_90e3040, \43029 );
buf \U$labajz4433 ( R_d7_90efe50, \43031 );
buf \U$labajz4434 ( R_d8_90f1350, \43047 );
buf \U$labajz4435 ( R_d9_9fc71a8, \43050 );
buf \U$labajz4436 ( R_da_9fc9cf8, \43057 );
buf \U$labajz4437 ( R_db_90ef9b8, \43063 );
buf \U$labajz4438 ( R_dc_90e4540, \43065 );
buf \U$labajz4439 ( R_dd_90f0ac8, \43070 );
buf \U$labajz4440 ( R_de_90e30e8, \43072 );
buf \U$labajz4441 ( R_df_9fc6290, \43075 );
buf \U$labajz4442 ( R_e0_9fc78e0, \43077 );
buf \U$labajz4443 ( R_e1_90e5500, \43083 );
buf \U$labajz4444 ( R_e2_90e68b0, \43085 );
buf \U$labajz4445 ( R_e3_90eede8, \43092 );
buf \U$labajz4446 ( R_e4_90e64c0, \43098 );
buf \U$labajz4447 ( R_e5_9fc7100, \43105 );
buf \U$labajz4448 ( R_e6_90e2470, \43121 );
buf \U$labajz4449 ( R_e7_90ebea8, \43123 );
buf \U$labajz4450 ( R_e8_90e4a80, \43125 );
buf \U$labajz4451 ( R_e9_90ef910, \43127 );
buf \U$labajz4452 ( R_ea_9fc7c28, \43132 );
buf \U$labajz4453 ( R_eb_90eb4d0, \43137 );
buf \U$labajz4454 ( R_ec_90f14a0, \43139 );
buf \U$labajz4455 ( R_ed_90ef5c8, \43141 );
buf \U$labajz4456 ( R_ee_90e4498, \43143 );
buf \U$labajz4457 ( R_ef_90e4000, \43145 );
buf \U$labajz4458 ( R_f0_90f0048, \43147 );
buf \U$labajz4459 ( R_f1_90ea3c0, \43149 );
buf \U$labajz4460 ( R_f2_90f1e78, \43151 );
buf \U$labajz4461 ( R_f3_90f00f0, \43156 );
not \U$1 ( \254 , RIbe29380_53);
not \U$2 ( \255 , RIbe27d78_6);
nor \U$3 ( \256 , \254 , \255 );
xnor \U$4 ( \257 , RIbe27ee0_9, RIbe286d8_26);
xor \U$5 ( \258 , RIbe286d8_26, RIbe28570_23);
nor \U$6 ( \259 , \257 , \258 );
buf \U$7 ( \260 , \259 );
buf \U$8 ( \261 , \260 );
and \U$9 ( \262 , \261 , RIbe28e58_42);
buf \U$10 ( \263 , \258 );
buf \U$11 ( \264 , \263 );
and \U$12 ( \265 , \264 , RIbe28de0_41);
nor \U$13 ( \266 , \262 , \265 );
nand \U$14 ( \267 , RIbe286d8_26, RIbe28570_23);
and \U$15 ( \268 , \267 , RIbe27ee0_9);
buf \U$16 ( \269 , \268 );
not \U$17 ( \270 , \269 );
buf \U$18 ( \271 , \270 );
not \U$19 ( \272 , \271 );
and \U$20 ( \273 , \266 , \272 );
not \U$21 ( \274 , \266 );
and \U$22 ( \275 , \274 , \271 );
nor \U$23 ( \276 , \273 , \275 );
not \U$24 ( \277 , \276 );
xnor \U$25 ( \278 , RIbe28570_23, RIbe28840_29);
xor \U$26 ( \279 , RIbe28840_29, RIbe28750_27);
nor \U$27 ( \280 , \278 , \279 );
not \U$28 ( \281 , \280 );
buf \U$29 ( \282 , \281 );
not \U$30 ( \283 , \282 );
and \U$31 ( \284 , \283 , RIbe29920_65);
not \U$32 ( \285 , \279 );
buf \U$33 ( \286 , \285 );
not \U$34 ( \287 , \286 );
and \U$35 ( \288 , \287 , RIbe27b98_2);
nor \U$36 ( \289 , \284 , \288 );
and \U$37 ( \290 , RIbe28840_29, RIbe28750_27);
not \U$38 ( \291 , RIbe28570_23);
nor \U$39 ( \292 , \290 , \291 );
buf \U$40 ( \293 , \292 );
and \U$41 ( \294 , \289 , \293 );
not \U$42 ( \295 , \289 );
not \U$43 ( \296 , RIbe28750_27);
not \U$44 ( \297 , RIbe28840_29);
or \U$45 ( \298 , \296 , \297 );
nand \U$46 ( \299 , \298 , RIbe28570_23);
buf \U$47 ( \300 , \299 );
and \U$48 ( \301 , \295 , \300 );
nor \U$49 ( \302 , \294 , \301 );
and \U$50 ( \303 , RIbe284f8_22, RIbe28318_18);
not \U$51 ( \304 , RIbe28750_27);
nor \U$52 ( \305 , \303 , \304 );
buf \U$53 ( \306 , \305 );
and \U$54 ( \307 , \302 , \306 );
not \U$55 ( \308 , \302 );
not \U$56 ( \309 , RIbe284f8_22);
not \U$57 ( \310 , RIbe28318_18);
or \U$58 ( \311 , \309 , \310 );
nand \U$59 ( \312 , \311 , RIbe28750_27);
buf \U$60 ( \313 , \312 );
and \U$61 ( \314 , \308 , \313 );
nor \U$62 ( \315 , \307 , \314 );
not \U$63 ( \316 , \315 );
or \U$64 ( \317 , \277 , \316 );
or \U$65 ( \318 , \315 , \276 );
nand \U$66 ( \319 , \317 , \318 );
xor \U$67 ( \320 , \256 , \319 );
xnor \U$68 ( \321 , RIbe29380_53, RIbe28048_12);
xor \U$69 ( \322 , RIbe28048_12, RIbe27ee0_9);
nor \U$70 ( \323 , \321 , \322 );
buf \U$71 ( \324 , \323 );
buf \U$72 ( \325 , \324 );
buf \U$73 ( \326 , \325 );
buf \U$74 ( \327 , \326 );
and \U$75 ( \328 , \327 , RIbe27d78_6);
buf \U$76 ( \329 , \322 );
buf \U$77 ( \330 , \329 );
buf \U$78 ( \331 , \330 );
and \U$79 ( \332 , \331 , RIbe27d00_5);
nor \U$80 ( \333 , \328 , \332 );
not \U$81 ( \334 , RIbe27ee0_9);
not \U$82 ( \335 , RIbe28048_12);
or \U$83 ( \336 , \334 , \335 );
nand \U$84 ( \337 , \336 , RIbe29380_53);
not \U$85 ( \338 , \337 );
not \U$86 ( \339 , \338 );
and \U$87 ( \340 , \333 , \339 );
not \U$88 ( \341 , \333 );
not \U$89 ( \342 , \339 );
and \U$90 ( \343 , \341 , \342 );
nor \U$91 ( \344 , \340 , \343 );
not \U$92 ( \345 , RIbe29380_53);
not \U$93 ( \346 , RIbe29a88_68);
nor \U$94 ( \347 , \345 , \346 );
or \U$95 ( \348 , \344 , \347 );
and \U$96 ( \349 , \327 , RIbe27d00_5);
and \U$97 ( \350 , \331 , RIbe27c10_3);
nor \U$98 ( \351 , \349 , \350 );
and \U$99 ( \352 , \351 , \339 );
not \U$100 ( \353 , \351 );
and \U$101 ( \354 , \353 , \342 );
nor \U$102 ( \355 , \352 , \354 );
xor \U$103 ( \356 , \348 , \355 );
and \U$104 ( \357 , \283 , RIbe28de0_41);
and \U$105 ( \358 , \287 , RIbe29920_65);
nor \U$106 ( \359 , \357 , \358 );
and \U$107 ( \360 , \359 , \293 );
not \U$108 ( \361 , \359 );
and \U$109 ( \362 , \361 , \300 );
nor \U$110 ( \363 , \360 , \362 );
and \U$111 ( \364 , \261 , RIbe27c10_3);
and \U$112 ( \365 , \264 , RIbe28e58_42);
nor \U$113 ( \366 , \364 , \365 );
and \U$114 ( \367 , \366 , \272 );
not \U$115 ( \368 , \366 );
and \U$116 ( \369 , \368 , \271 );
nor \U$117 ( \370 , \367 , \369 );
or \U$118 ( \371 , \363 , \370 );
not \U$119 ( \372 , \370 );
not \U$120 ( \373 , \363 );
or \U$121 ( \374 , \372 , \373 );
xnor \U$122 ( \375 , RIbe284f8_22, RIbe28318_18);
not \U$123 ( \376 , RIbe284f8_22);
nand \U$124 ( \377 , \376 , RIbe28750_27);
not \U$125 ( \378 , RIbe28750_27);
nand \U$126 ( \379 , \378 , RIbe284f8_22);
nand \U$127 ( \380 , \377 , \379 );
nand \U$128 ( \381 , \375 , \380 );
buf \U$129 ( \382 , \381 );
not \U$130 ( \383 , \382 );
nand \U$131 ( \384 , \383 , RIbe27b98_2);
and \U$132 ( \385 , \384 , \313 );
not \U$133 ( \386 , \384 );
and \U$134 ( \387 , \386 , \306 );
nor \U$135 ( \388 , \385 , \387 );
nand \U$136 ( \389 , \374 , \388 );
nand \U$137 ( \390 , \371 , \389 );
xor \U$138 ( \391 , \356 , \390 );
and \U$139 ( \392 , \320 , \391 );
not \U$140 ( \393 , \320 );
not \U$141 ( \394 , \391 );
and \U$142 ( \395 , \393 , \394 );
and \U$143 ( \396 , \261 , RIbe27d00_5);
and \U$144 ( \397 , \264 , RIbe27c10_3);
nor \U$145 ( \398 , \396 , \397 );
and \U$146 ( \399 , \398 , \272 );
not \U$147 ( \400 , \398 );
and \U$148 ( \401 , \400 , \271 );
nor \U$149 ( \402 , \399 , \401 );
nand \U$150 ( \403 , RIbe29380_53, RIbe290b0_47);
xor \U$151 ( \404 , \402 , \403 );
and \U$152 ( \405 , \327 , RIbe29a88_68);
and \U$153 ( \406 , \331 , RIbe27d78_6);
nor \U$154 ( \407 , \405 , \406 );
and \U$155 ( \408 , \407 , \342 );
not \U$156 ( \409 , \407 );
and \U$157 ( \410 , \409 , \339 );
nor \U$158 ( \411 , \408 , \410 );
and \U$159 ( \412 , \404 , \411 );
and \U$160 ( \413 , \402 , \403 );
or \U$161 ( \414 , \412 , \413 );
and \U$162 ( \415 , \283 , RIbe28e58_42);
and \U$163 ( \416 , \287 , RIbe28de0_41);
nor \U$164 ( \417 , \415 , \416 );
and \U$165 ( \418 , \417 , \293 );
not \U$166 ( \419 , \417 );
and \U$167 ( \420 , \419 , \300 );
nor \U$168 ( \421 , \418 , \420 );
nand \U$169 ( \422 , RIbe28c78_38, RIbe28c00_37);
nand \U$170 ( \423 , \422 , RIbe28318_18);
buf \U$171 ( \424 , \423 );
not \U$172 ( \425 , \424 );
xor \U$173 ( \426 , \421 , \425 );
and \U$174 ( \427 , \383 , RIbe29920_65);
xor \U$175 ( \428 , RIbe284f8_22, RIbe28318_18);
buf \U$176 ( \429 , \428 );
and \U$177 ( \430 , \429 , RIbe27b98_2);
nor \U$178 ( \431 , \427 , \430 );
and \U$179 ( \432 , \431 , \306 );
not \U$180 ( \433 , \431 );
and \U$181 ( \434 , \433 , \313 );
nor \U$182 ( \435 , \432 , \434 );
and \U$183 ( \436 , \426 , \435 );
and \U$184 ( \437 , \421 , \425 );
or \U$185 ( \438 , \436 , \437 );
xor \U$186 ( \439 , \414 , \438 );
and \U$187 ( \440 , \344 , \347 );
not \U$188 ( \441 , \348 );
nor \U$189 ( \442 , \440 , \441 );
and \U$190 ( \443 , \439 , \442 );
and \U$191 ( \444 , \414 , \438 );
or \U$192 ( \445 , \443 , \444 );
nor \U$193 ( \446 , \395 , \445 );
nor \U$194 ( \447 , \392 , \446 );
not \U$195 ( \448 , \447 );
and \U$196 ( \449 , \256 , \319 );
xor \U$197 ( \450 , \348 , \355 );
and \U$198 ( \451 , \450 , \390 );
and \U$199 ( \452 , \348 , \355 );
or \U$200 ( \453 , \451 , \452 );
xor \U$201 ( \454 , \449 , \453 );
not \U$202 ( \455 , \276 );
not \U$203 ( \456 , \306 );
and \U$204 ( \457 , \455 , \456 );
and \U$205 ( \458 , \276 , \306 );
nor \U$206 ( \459 , \458 , \302 );
nor \U$207 ( \460 , \457 , \459 );
and \U$208 ( \461 , RIbe29380_53, RIbe27d00_5);
and \U$209 ( \462 , \460 , \461 );
nor \U$210 ( \463 , \460 , \461 );
or \U$211 ( \464 , \462 , \463 );
not \U$212 ( \465 , \464 );
and \U$213 ( \466 , \261 , RIbe28de0_41);
and \U$214 ( \467 , \264 , RIbe29920_65);
nor \U$215 ( \468 , \466 , \467 );
and \U$216 ( \469 , \468 , \272 );
not \U$217 ( \470 , \468 );
and \U$218 ( \471 , \470 , \271 );
nor \U$219 ( \472 , \469 , \471 );
nand \U$220 ( \473 , \283 , RIbe27b98_2);
and \U$221 ( \474 , \473 , \293 );
not \U$222 ( \475 , \473 );
and \U$223 ( \476 , \475 , \300 );
nor \U$224 ( \477 , \474 , \476 );
xor \U$225 ( \478 , \472 , \477 );
and \U$226 ( \479 , \327 , RIbe27c10_3);
and \U$227 ( \480 , \331 , RIbe28e58_42);
nor \U$228 ( \481 , \479 , \480 );
and \U$229 ( \482 , \481 , \342 );
not \U$230 ( \483 , \481 );
and \U$231 ( \484 , \483 , \339 );
nor \U$232 ( \485 , \482 , \484 );
xor \U$233 ( \486 , \478 , \485 );
not \U$234 ( \487 , \486 );
and \U$235 ( \488 , \465 , \487 );
and \U$236 ( \489 , \464 , \486 );
nor \U$237 ( \490 , \488 , \489 );
xor \U$238 ( \491 , \454 , \490 );
nand \U$239 ( \492 , \448 , \491 );
not \U$240 ( \493 , \492 );
xor \U$241 ( \494 , \449 , \453 );
and \U$242 ( \495 , \494 , \490 );
and \U$243 ( \496 , \449 , \453 );
or \U$244 ( \497 , \495 , \496 );
not \U$245 ( \498 , \497 );
not \U$246 ( \499 , \461 );
nand \U$247 ( \500 , RIbe29380_53, RIbe27c10_3);
xor \U$248 ( \501 , \499 , \500 );
xor \U$249 ( \502 , \472 , \477 );
and \U$250 ( \503 , \502 , \485 );
and \U$251 ( \504 , \472 , \477 );
or \U$252 ( \505 , \503 , \504 );
xor \U$253 ( \506 , \501 , \505 );
and \U$254 ( \507 , \261 , RIbe29920_65);
and \U$255 ( \508 , \264 , RIbe27b98_2);
nor \U$256 ( \509 , \507 , \508 );
and \U$257 ( \510 , \509 , \272 );
not \U$258 ( \511 , \509 );
and \U$259 ( \512 , \511 , \271 );
nor \U$260 ( \513 , \510 , \512 );
xor \U$261 ( \514 , \513 , \293 );
and \U$262 ( \515 , \327 , RIbe28e58_42);
and \U$263 ( \516 , \331 , RIbe28de0_41);
nor \U$264 ( \517 , \515 , \516 );
and \U$265 ( \518 , \517 , \342 );
not \U$266 ( \519 , \517 );
and \U$267 ( \520 , \519 , \339 );
nor \U$268 ( \521 , \518 , \520 );
xor \U$269 ( \522 , \514 , \521 );
not \U$270 ( \523 , \486 );
not \U$271 ( \524 , \462 );
and \U$272 ( \525 , \523 , \524 );
nor \U$273 ( \526 , \525 , \463 );
xor \U$274 ( \527 , \522 , \526 );
xor \U$275 ( \528 , \506 , \527 );
not \U$276 ( \529 , \528 );
or \U$277 ( \530 , \498 , \529 );
or \U$278 ( \531 , \528 , \497 );
nand \U$279 ( \532 , \530 , \531 );
not \U$280 ( \533 , \532 );
or \U$281 ( \534 , \493 , \533 );
or \U$282 ( \535 , \532 , \492 );
nand \U$283 ( \536 , \534 , \535 );
not \U$284 ( \537 , \536 );
not \U$285 ( \538 , RIbe28318_18);
nand \U$286 ( \539 , \538 , RIbe28c78_38);
and \U$287 ( \540 , RIbe28c00_37, \539 );
not \U$288 ( \541 , RIbe28c00_37);
not \U$289 ( \542 , RIbe28c78_38);
nand \U$290 ( \543 , \542 , RIbe28318_18);
and \U$291 ( \544 , \541 , \543 );
nor \U$292 ( \545 , \540 , \544 );
buf \U$293 ( \546 , \545 );
not \U$294 ( \547 , \546 );
not \U$295 ( \548 , \547 );
buf \U$296 ( \549 , \548 );
and \U$297 ( \550 , \549 , RIbe29920_65);
xor \U$298 ( \551 , RIbe28c78_38, RIbe28c00_37);
buf \U$299 ( \552 , \551 );
buf \U$300 ( \553 , \552 );
buf \U$301 ( \554 , \553 );
and \U$302 ( \555 , \554 , RIbe27b98_2);
nor \U$303 ( \556 , \550 , \555 );
and \U$304 ( \557 , \556 , \424 );
not \U$305 ( \558 , \556 );
and \U$306 ( \559 , \558 , \425 );
nor \U$307 ( \560 , \557 , \559 );
nand \U$308 ( \561 , RIbe29308_52, RIbe293f8_54);
buf \U$309 ( \562 , \561 );
nand \U$310 ( \563 , \562 , RIbe28c00_37);
buf \U$311 ( \564 , \563 );
xor \U$312 ( \565 , \560 , \564 );
and \U$313 ( \566 , \383 , RIbe28e58_42);
and \U$314 ( \567 , \429 , RIbe28de0_41);
nor \U$315 ( \568 , \566 , \567 );
and \U$316 ( \569 , \568 , \313 );
not \U$317 ( \570 , \568 );
and \U$318 ( \571 , \570 , \306 );
nor \U$319 ( \572 , \569 , \571 );
xor \U$320 ( \573 , \565 , \572 );
not \U$321 ( \574 , \573 );
nand \U$322 ( \575 , RIbe29380_53, RIbe29038_46);
nand \U$323 ( \576 , \574 , \575 );
and \U$324 ( \577 , \261 , RIbe29a88_68);
and \U$325 ( \578 , \264 , RIbe27d78_6);
nor \U$326 ( \579 , \577 , \578 );
and \U$327 ( \580 , \579 , \271 );
not \U$328 ( \581 , \579 );
and \U$329 ( \582 , \581 , \272 );
nor \U$330 ( \583 , \580 , \582 );
and \U$331 ( \584 , \283 , RIbe27d00_5);
and \U$332 ( \585 , \287 , RIbe27c10_3);
nor \U$333 ( \586 , \584 , \585 );
and \U$334 ( \587 , \586 , \300 );
not \U$335 ( \588 , \586 );
and \U$336 ( \589 , \588 , \293 );
nor \U$337 ( \590 , \587 , \589 );
xor \U$338 ( \591 , \583 , \590 );
and \U$339 ( \592 , \327 , RIbe28fc0_45);
and \U$340 ( \593 , \331 , RIbe290b0_47);
nor \U$341 ( \594 , \592 , \593 );
and \U$342 ( \595 , \594 , \339 );
not \U$343 ( \596 , \594 );
and \U$344 ( \597 , \596 , \342 );
nor \U$345 ( \598 , \595 , \597 );
xor \U$346 ( \599 , \591 , \598 );
and \U$347 ( \600 , \576 , \599 );
not \U$348 ( \601 , \575 );
and \U$349 ( \602 , \573 , \601 );
nor \U$350 ( \603 , \600 , \602 );
and \U$351 ( \604 , \261 , RIbe27d78_6);
and \U$352 ( \605 , \264 , RIbe27d00_5);
nor \U$353 ( \606 , \604 , \605 );
and \U$354 ( \607 , \606 , \272 );
not \U$355 ( \608 , \606 );
and \U$356 ( \609 , \608 , \271 );
nor \U$357 ( \610 , \607 , \609 );
nand \U$358 ( \611 , RIbe29380_53, RIbe28fc0_45);
xor \U$359 ( \612 , \610 , \611 );
and \U$360 ( \613 , \327 , RIbe290b0_47);
and \U$361 ( \614 , \331 , RIbe29a88_68);
nor \U$362 ( \615 , \613 , \614 );
and \U$363 ( \616 , \615 , \342 );
not \U$364 ( \617 , \615 );
and \U$365 ( \618 , \617 , \339 );
nor \U$366 ( \619 , \616 , \618 );
xor \U$367 ( \620 , \612 , \619 );
xor \U$368 ( \621 , \603 , \620 );
and \U$369 ( \622 , \327 , RIbe29038_46);
and \U$370 ( \623 , \331 , RIbe28fc0_45);
nor \U$371 ( \624 , \622 , \623 );
and \U$372 ( \625 , \624 , \339 );
not \U$373 ( \626 , \624 );
and \U$374 ( \627 , \626 , \342 );
nor \U$375 ( \628 , \625 , \627 );
and \U$376 ( \629 , \283 , RIbe27d78_6);
and \U$377 ( \630 , \287 , RIbe27d00_5);
nor \U$378 ( \631 , \629 , \630 );
and \U$379 ( \632 , \631 , \300 );
not \U$380 ( \633 , \631 );
and \U$381 ( \634 , \633 , \293 );
nor \U$382 ( \635 , \632 , \634 );
xor \U$383 ( \636 , \628 , \635 );
and \U$384 ( \637 , \261 , RIbe290b0_47);
and \U$385 ( \638 , \264 , RIbe29a88_68);
nor \U$386 ( \639 , \637 , \638 );
and \U$387 ( \640 , \639 , \271 );
not \U$388 ( \641 , \639 );
and \U$389 ( \642 , \641 , \272 );
nor \U$390 ( \643 , \640 , \642 );
and \U$391 ( \644 , \636 , \643 );
and \U$392 ( \645 , \628 , \635 );
or \U$393 ( \646 , \644 , \645 );
nand \U$394 ( \647 , RIbe29380_53, RIbe29650_59);
not \U$395 ( \648 , \647 );
and \U$396 ( \649 , \646 , \648 );
not \U$397 ( \650 , \646 );
not \U$398 ( \651 , \648 );
and \U$399 ( \652 , \650 , \651 );
and \U$400 ( \653 , \549 , RIbe28de0_41);
and \U$401 ( \654 , \554 , RIbe29920_65);
nor \U$402 ( \655 , \653 , \654 );
and \U$403 ( \656 , \655 , \424 );
not \U$404 ( \657 , \655 );
and \U$405 ( \658 , \657 , \425 );
nor \U$406 ( \659 , \656 , \658 );
or \U$407 ( \660 , \561 , RIbe28c00_37);
nor \U$408 ( \661 , RIbe29308_52, RIbe293f8_54);
nand \U$409 ( \662 , \661 , RIbe28c00_37);
nand \U$410 ( \663 , \660 , \662 );
buf \U$411 ( \664 , \663 );
not \U$412 ( \665 , \664 );
not \U$413 ( \666 , \665 );
nand \U$414 ( \667 , \666 , RIbe27b98_2);
and \U$415 ( \668 , \667 , \564 );
not \U$416 ( \669 , \667 );
and \U$417 ( \670 , \562 , RIbe28c00_37);
not \U$418 ( \671 , \670 );
not \U$419 ( \672 , \671 );
and \U$420 ( \673 , \669 , \672 );
nor \U$421 ( \674 , \668 , \673 );
xor \U$422 ( \675 , \659 , \674 );
and \U$423 ( \676 , \383 , RIbe27c10_3);
and \U$424 ( \677 , \429 , RIbe28e58_42);
nor \U$425 ( \678 , \676 , \677 );
and \U$426 ( \679 , \678 , \313 );
not \U$427 ( \680 , \678 );
and \U$428 ( \681 , \680 , \306 );
nor \U$429 ( \682 , \679 , \681 );
and \U$430 ( \683 , \675 , \682 );
and \U$431 ( \684 , \659 , \674 );
nor \U$432 ( \685 , \683 , \684 );
nor \U$433 ( \686 , \652 , \685 );
nor \U$434 ( \687 , \649 , \686 );
xor \U$435 ( \688 , \621 , \687 );
xor \U$436 ( \689 , \583 , \590 );
and \U$437 ( \690 , \689 , \598 );
and \U$438 ( \691 , \583 , \590 );
or \U$439 ( \692 , \690 , \691 );
xor \U$440 ( \693 , \560 , \564 );
and \U$441 ( \694 , \693 , \572 );
and \U$442 ( \695 , \560 , \564 );
or \U$443 ( \696 , \694 , \695 );
and \U$444 ( \697 , \692 , \696 );
nor \U$445 ( \698 , \692 , \696 );
nor \U$446 ( \699 , \697 , \698 );
not \U$447 ( \700 , \699 );
not \U$448 ( \701 , \293 );
and \U$449 ( \702 , \283 , RIbe27c10_3);
and \U$450 ( \703 , \287 , RIbe28e58_42);
nor \U$451 ( \704 , \702 , \703 );
not \U$452 ( \705 , \704 );
or \U$453 ( \706 , \701 , \705 );
or \U$454 ( \707 , \704 , \293 );
nand \U$455 ( \708 , \706 , \707 );
nand \U$456 ( \709 , \549 , RIbe27b98_2);
and \U$457 ( \710 , \709 , \424 );
not \U$458 ( \711 , \709 );
and \U$459 ( \712 , \711 , \425 );
nor \U$460 ( \713 , \710 , \712 );
xor \U$461 ( \714 , \708 , \713 );
and \U$462 ( \715 , \383 , RIbe28de0_41);
and \U$463 ( \716 , \429 , RIbe29920_65);
nor \U$464 ( \717 , \715 , \716 );
and \U$465 ( \718 , \717 , \313 );
not \U$466 ( \719 , \717 );
and \U$467 ( \720 , \719 , \306 );
nor \U$468 ( \721 , \718 , \720 );
xor \U$469 ( \722 , \714 , \721 );
not \U$470 ( \723 , \722 );
and \U$471 ( \724 , \700 , \723 );
and \U$472 ( \725 , \699 , \722 );
nor \U$473 ( \726 , \724 , \725 );
or \U$474 ( \727 , \688 , \726 );
not \U$475 ( \728 , \726 );
not \U$476 ( \729 , \688 );
or \U$477 ( \730 , \728 , \729 );
xor \U$478 ( \731 , \659 , \674 );
xor \U$479 ( \732 , \731 , \682 );
xor \U$480 ( \733 , \732 , \647 );
xor \U$481 ( \734 , \628 , \635 );
xor \U$482 ( \735 , \734 , \643 );
and \U$483 ( \736 , \733 , \735 );
and \U$484 ( \737 , \732 , \647 );
or \U$485 ( \738 , \736 , \737 );
and \U$486 ( \739 , \666 , RIbe29920_65);
xor \U$487 ( \740 , RIbe29308_52, RIbe293f8_54);
and \U$488 ( \741 , \740 , RIbe27b98_2);
nor \U$489 ( \742 , \739 , \741 );
and \U$490 ( \743 , \742 , \564 );
not \U$491 ( \744 , \742 );
and \U$492 ( \745 , \744 , \672 );
nor \U$493 ( \746 , \743 , \745 );
not \U$494 ( \747 , RIbe288b8_30);
not \U$495 ( \748 , RIbe28a98_34);
or \U$496 ( \749 , \747 , \748 );
nand \U$497 ( \750 , \749 , RIbe293f8_54);
not \U$498 ( \751 , \750 );
not \U$499 ( \752 , \751 );
xor \U$500 ( \753 , \746 , \752 );
and \U$501 ( \754 , \549 , RIbe28e58_42);
and \U$502 ( \755 , \554 , RIbe28de0_41);
nor \U$503 ( \756 , \754 , \755 );
and \U$504 ( \757 , \756 , \424 );
not \U$505 ( \758 , \756 );
and \U$506 ( \759 , \758 , \425 );
nor \U$507 ( \760 , \757 , \759 );
and \U$508 ( \761 , \753 , \760 );
and \U$509 ( \762 , \746 , \752 );
or \U$510 ( \763 , \761 , \762 );
and \U$511 ( \764 , RIbe296c8_60, RIbe29380_53);
and \U$512 ( \765 , \327 , RIbe29650_59);
and \U$513 ( \766 , \331 , RIbe29038_46);
nor \U$514 ( \767 , \765 , \766 );
and \U$515 ( \768 , \767 , \339 );
not \U$516 ( \769 , \767 );
and \U$517 ( \770 , \769 , \342 );
nor \U$518 ( \771 , \768 , \770 );
and \U$519 ( \772 , \764 , \771 );
xor \U$520 ( \773 , \763 , \772 );
and \U$521 ( \774 , \383 , RIbe27d00_5);
and \U$522 ( \775 , \429 , RIbe27c10_3);
nor \U$523 ( \776 , \774 , \775 );
and \U$524 ( \777 , \776 , \313 );
not \U$525 ( \778 , \776 );
and \U$526 ( \779 , \778 , \306 );
nor \U$527 ( \780 , \777 , \779 );
and \U$528 ( \781 , \261 , RIbe28fc0_45);
and \U$529 ( \782 , \264 , RIbe290b0_47);
nor \U$530 ( \783 , \781 , \782 );
and \U$531 ( \784 , \783 , \271 );
not \U$532 ( \785 , \783 );
and \U$533 ( \786 , \785 , \272 );
nor \U$534 ( \787 , \784 , \786 );
xor \U$535 ( \788 , \780 , \787 );
and \U$536 ( \789 , \283 , RIbe29a88_68);
and \U$537 ( \790 , \287 , RIbe27d78_6);
nor \U$538 ( \791 , \789 , \790 );
and \U$539 ( \792 , \791 , \300 );
not \U$540 ( \793 , \791 );
and \U$541 ( \794 , \793 , \293 );
nor \U$542 ( \795 , \792 , \794 );
and \U$543 ( \796 , \788 , \795 );
and \U$544 ( \797 , \780 , \787 );
or \U$545 ( \798 , \796 , \797 );
and \U$546 ( \799 , \773 , \798 );
and \U$547 ( \800 , \763 , \772 );
or \U$548 ( \801 , \799 , \800 );
xor \U$549 ( \802 , \738 , \801 );
not \U$550 ( \803 , \573 );
not \U$551 ( \804 , \599 );
not \U$552 ( \805 , \575 );
and \U$553 ( \806 , \804 , \805 );
and \U$554 ( \807 , \599 , \575 );
nor \U$555 ( \808 , \806 , \807 );
not \U$556 ( \809 , \808 );
or \U$557 ( \810 , \803 , \809 );
or \U$558 ( \811 , \808 , \573 );
nand \U$559 ( \812 , \810 , \811 );
and \U$560 ( \813 , \802 , \812 );
and \U$561 ( \814 , \738 , \801 );
or \U$562 ( \815 , \813 , \814 );
nand \U$563 ( \816 , \730 , \815 );
nand \U$564 ( \817 , \727 , \816 );
xor \U$565 ( \818 , \421 , \425 );
xor \U$566 ( \819 , \818 , \435 );
xor \U$567 ( \820 , \610 , \611 );
and \U$568 ( \821 , \820 , \619 );
and \U$569 ( \822 , \610 , \611 );
or \U$570 ( \823 , \821 , \822 );
not \U$571 ( \824 , \823 );
xor \U$572 ( \825 , \708 , \713 );
and \U$573 ( \826 , \825 , \721 );
and \U$574 ( \827 , \708 , \713 );
or \U$575 ( \828 , \826 , \827 );
not \U$576 ( \829 , \828 );
or \U$577 ( \830 , \824 , \829 );
or \U$578 ( \831 , \828 , \823 );
nand \U$579 ( \832 , \830 , \831 );
not \U$580 ( \833 , \832 );
xor \U$581 ( \834 , \402 , \403 );
xor \U$582 ( \835 , \834 , \411 );
not \U$583 ( \836 , \835 );
and \U$584 ( \837 , \833 , \836 );
and \U$585 ( \838 , \832 , \835 );
nor \U$586 ( \839 , \837 , \838 );
xor \U$587 ( \840 , \698 , \839 );
xor \U$588 ( \841 , \819 , \840 );
not \U$589 ( \842 , \841 );
not \U$590 ( \843 , \722 );
nor \U$591 ( \844 , \843 , \699 );
not \U$592 ( \845 , \844 );
xor \U$593 ( \846 , \603 , \620 );
and \U$594 ( \847 , \846 , \687 );
and \U$595 ( \848 , \603 , \620 );
or \U$596 ( \849 , \847 , \848 );
not \U$597 ( \850 , \849 );
or \U$598 ( \851 , \845 , \850 );
or \U$599 ( \852 , \849 , \844 );
nand \U$600 ( \853 , \851 , \852 );
not \U$601 ( \854 , \853 );
or \U$602 ( \855 , \842 , \854 );
or \U$603 ( \856 , \853 , \841 );
nand \U$604 ( \857 , \855 , \856 );
and \U$605 ( \858 , \817 , \857 );
not \U$606 ( \859 , \858 );
not \U$607 ( \860 , \388 );
not \U$608 ( \861 , \363 );
or \U$609 ( \862 , \860 , \861 );
or \U$610 ( \863 , \363 , \388 );
nand \U$611 ( \864 , \862 , \863 );
not \U$612 ( \865 , \864 );
not \U$613 ( \866 , \370 );
and \U$614 ( \867 , \865 , \866 );
and \U$615 ( \868 , \864 , \370 );
nor \U$616 ( \869 , \867 , \868 );
not \U$617 ( \870 , \869 );
or \U$618 ( \871 , \835 , \823 );
not \U$619 ( \872 , \823 );
not \U$620 ( \873 , \835 );
or \U$621 ( \874 , \872 , \873 );
nand \U$622 ( \875 , \874 , \828 );
nand \U$623 ( \876 , \871 , \875 );
not \U$624 ( \877 , \876 );
or \U$625 ( \878 , \870 , \877 );
or \U$626 ( \879 , \876 , \869 );
nand \U$627 ( \880 , \878 , \879 );
not \U$628 ( \881 , \880 );
xor \U$629 ( \882 , \414 , \438 );
xor \U$630 ( \883 , \882 , \442 );
not \U$631 ( \884 , \883 );
and \U$632 ( \885 , \881 , \884 );
and \U$633 ( \886 , \880 , \883 );
nor \U$634 ( \887 , \885 , \886 );
xor \U$635 ( \888 , \421 , \425 );
xor \U$636 ( \889 , \888 , \435 );
and \U$637 ( \890 , \698 , \889 );
xor \U$638 ( \891 , \421 , \425 );
xor \U$639 ( \892 , \891 , \435 );
and \U$640 ( \893 , \839 , \892 );
and \U$641 ( \894 , \698 , \839 );
or \U$642 ( \895 , \890 , \893 , \894 );
xor \U$643 ( \896 , \887 , \895 );
not \U$644 ( \897 , \841 );
and \U$645 ( \898 , \897 , \844 );
not \U$646 ( \899 , \897 );
not \U$647 ( \900 , \844 );
and \U$648 ( \901 , \899 , \900 );
nor \U$649 ( \902 , \901 , \849 );
nor \U$650 ( \903 , \898 , \902 );
xor \U$651 ( \904 , \896 , \903 );
not \U$652 ( \905 , \904 );
or \U$653 ( \906 , \859 , \905 );
or \U$654 ( \907 , \904 , \858 );
nand \U$655 ( \908 , \906 , \907 );
not \U$656 ( \909 , \447 );
not \U$657 ( \910 , \491 );
or \U$658 ( \911 , \909 , \910 );
or \U$659 ( \912 , \491 , \447 );
nand \U$660 ( \913 , \911 , \912 );
or \U$661 ( \914 , \883 , \869 );
not \U$662 ( \915 , \869 );
not \U$663 ( \916 , \883 );
or \U$664 ( \917 , \915 , \916 );
nand \U$665 ( \918 , \917 , \876 );
nand \U$666 ( \919 , \914 , \918 );
not \U$667 ( \920 , \391 );
not \U$668 ( \921 , \445 );
or \U$669 ( \922 , \920 , \921 );
or \U$670 ( \923 , \445 , \391 );
nand \U$671 ( \924 , \922 , \923 );
xor \U$672 ( \925 , \320 , \924 );
and \U$673 ( \926 , \919 , \925 );
xor \U$674 ( \927 , \913 , \926 );
not \U$675 ( \928 , \927 );
xor \U$676 ( \929 , \887 , \895 );
and \U$677 ( \930 , \929 , \903 );
and \U$678 ( \931 , \887 , \895 );
or \U$679 ( \932 , \930 , \931 );
not \U$680 ( \933 , \932 );
xor \U$681 ( \934 , \919 , \925 );
not \U$682 ( \935 , \934 );
and \U$683 ( \936 , \933 , \935 );
and \U$684 ( \937 , \932 , \934 );
nor \U$685 ( \938 , \936 , \937 );
nor \U$686 ( \939 , \928 , \938 );
and \U$687 ( \940 , \908 , \939 );
not \U$688 ( \941 , \940 );
not \U$689 ( \942 , \726 );
not \U$690 ( \943 , \815 );
or \U$691 ( \944 , \942 , \943 );
or \U$692 ( \945 , \815 , \726 );
nand \U$693 ( \946 , \944 , \945 );
not \U$694 ( \947 , \946 );
not \U$695 ( \948 , \688 );
and \U$696 ( \949 , \947 , \948 );
and \U$697 ( \950 , \946 , \688 );
nor \U$698 ( \951 , \949 , \950 );
not \U$699 ( \952 , \951 );
not \U$700 ( \953 , \647 );
not \U$701 ( \954 , \685 );
not \U$702 ( \955 , \646 );
or \U$703 ( \956 , \954 , \955 );
or \U$704 ( \957 , \646 , \685 );
nand \U$705 ( \958 , \956 , \957 );
not \U$706 ( \959 , \958 );
or \U$707 ( \960 , \953 , \959 );
or \U$708 ( \961 , \958 , \647 );
nand \U$709 ( \962 , \960 , \961 );
not \U$710 ( \963 , \962 );
xor \U$711 ( \964 , \738 , \801 );
xor \U$712 ( \965 , \964 , \812 );
not \U$713 ( \966 , \965 );
or \U$714 ( \967 , \963 , \966 );
or \U$715 ( \968 , \965 , \962 );
xor \U$716 ( \969 , \764 , \771 );
xor \U$717 ( \970 , \746 , \752 );
xor \U$718 ( \971 , \970 , \760 );
and \U$719 ( \972 , \969 , \971 );
xor \U$720 ( \973 , \780 , \787 );
xor \U$721 ( \974 , \973 , \795 );
xor \U$722 ( \975 , \746 , \752 );
xor \U$723 ( \976 , \975 , \760 );
and \U$724 ( \977 , \974 , \976 );
and \U$725 ( \978 , \969 , \974 );
or \U$726 ( \979 , \972 , \977 , \978 );
and \U$727 ( \980 , \549 , RIbe27c10_3);
and \U$728 ( \981 , \554 , RIbe28e58_42);
nor \U$729 ( \982 , \980 , \981 );
and \U$730 ( \983 , \982 , \425 );
not \U$731 ( \984 , \982 );
and \U$732 ( \985 , \984 , \424 );
nor \U$733 ( \986 , \983 , \985 );
and \U$734 ( \987 , \666 , RIbe28de0_41);
and \U$735 ( \988 , \740 , RIbe29920_65);
nor \U$736 ( \989 , \987 , \988 );
and \U$737 ( \990 , \989 , \672 );
not \U$738 ( \991 , \989 );
and \U$739 ( \992 , \991 , \564 );
nor \U$740 ( \993 , \990 , \992 );
or \U$741 ( \994 , \986 , \993 );
not \U$742 ( \995 , \993 );
not \U$743 ( \996 , \986 );
or \U$744 ( \997 , \995 , \996 );
xor \U$745 ( \998 , RIbe28a98_34, RIbe288b8_30);
not \U$746 ( \999 , \998 );
xor \U$747 ( \1000 , RIbe293f8_54, RIbe28a98_34);
nand \U$748 ( \1001 , \999 , \1000 );
not \U$749 ( \1002 , \1001 );
buf \U$750 ( \1003 , \1002 );
not \U$751 ( \1004 , \1003 );
not \U$752 ( \1005 , \1004 );
nand \U$753 ( \1006 , \1005 , RIbe27b98_2);
and \U$754 ( \1007 , \1006 , \752 );
not \U$755 ( \1008 , \1006 );
nand \U$756 ( \1009 , RIbe28a98_34, RIbe288b8_30);
and \U$757 ( \1010 , \1009 , RIbe293f8_54);
buf \U$758 ( \1011 , \1010 );
and \U$759 ( \1012 , \1008 , \1011 );
nor \U$760 ( \1013 , \1007 , \1012 );
nand \U$761 ( \1014 , \997 , \1013 );
nand \U$762 ( \1015 , \994 , \1014 );
and \U$763 ( \1016 , \327 , RIbe296c8_60);
and \U$764 ( \1017 , \331 , RIbe29650_59);
nor \U$765 ( \1018 , \1016 , \1017 );
and \U$766 ( \1019 , \1018 , \342 );
not \U$767 ( \1020 , \1018 );
and \U$768 ( \1021 , \1020 , \339 );
nor \U$769 ( \1022 , \1019 , \1021 );
nand \U$770 ( \1023 , RIbe29380_53, RIbe29830_63);
nand \U$771 ( \1024 , \1022 , \1023 );
xor \U$772 ( \1025 , \1015 , \1024 );
and \U$773 ( \1026 , \383 , RIbe27d78_6);
and \U$774 ( \1027 , \429 , RIbe27d00_5);
nor \U$775 ( \1028 , \1026 , \1027 );
and \U$776 ( \1029 , \1028 , \306 );
not \U$777 ( \1030 , \1028 );
and \U$778 ( \1031 , \1030 , \313 );
nor \U$779 ( \1032 , \1029 , \1031 );
and \U$780 ( \1033 , \261 , RIbe29038_46);
and \U$781 ( \1034 , \264 , RIbe28fc0_45);
nor \U$782 ( \1035 , \1033 , \1034 );
and \U$783 ( \1036 , \1035 , \272 );
not \U$784 ( \1037 , \1035 );
and \U$785 ( \1038 , \1037 , \271 );
nor \U$786 ( \1039 , \1036 , \1038 );
or \U$787 ( \1040 , \1032 , \1039 );
not \U$788 ( \1041 , \1039 );
not \U$789 ( \1042 , \1032 );
or \U$790 ( \1043 , \1041 , \1042 );
and \U$791 ( \1044 , \283 , RIbe290b0_47);
and \U$792 ( \1045 , \287 , RIbe29a88_68);
nor \U$793 ( \1046 , \1044 , \1045 );
and \U$794 ( \1047 , \1046 , \300 );
not \U$795 ( \1048 , \1046 );
and \U$796 ( \1049 , \1048 , \293 );
nor \U$797 ( \1050 , \1047 , \1049 );
nand \U$798 ( \1051 , \1043 , \1050 );
nand \U$799 ( \1052 , \1040 , \1051 );
and \U$800 ( \1053 , \1025 , \1052 );
and \U$801 ( \1054 , \1015 , \1024 );
or \U$802 ( \1055 , \1053 , \1054 );
xor \U$803 ( \1056 , \979 , \1055 );
xor \U$804 ( \1057 , \732 , \647 );
xor \U$805 ( \1058 , \1057 , \735 );
and \U$806 ( \1059 , \1056 , \1058 );
and \U$807 ( \1060 , \979 , \1055 );
or \U$808 ( \1061 , \1059 , \1060 );
nand \U$809 ( \1062 , \968 , \1061 );
nand \U$810 ( \1063 , \967 , \1062 );
nand \U$811 ( \1064 , \952 , \1063 );
not \U$812 ( \1065 , \1064 );
xor \U$813 ( \1066 , \817 , \857 );
not \U$814 ( \1067 , \1066 );
or \U$815 ( \1068 , \1065 , \1067 );
or \U$816 ( \1069 , \1066 , \1064 );
nand \U$817 ( \1070 , \1068 , \1069 );
not \U$818 ( \1071 , \1070 );
not \U$819 ( \1072 , RIbe291a0_49);
not \U$820 ( \1073 , RIbe295d8_58);
or \U$821 ( \1074 , \1072 , \1073 );
nand \U$822 ( \1075 , \1074 , RIbe29740_61);
buf \U$823 ( \1076 , \1075 );
not \U$824 ( \1077 , RIbe282a0_17);
not \U$825 ( \1078 , RIbe28138_14);
or \U$826 ( \1079 , \1077 , \1078 );
nand \U$827 ( \1080 , \1079 , RIbe29470_55);
not \U$828 ( \1081 , \1080 );
not \U$829 ( \1082 , \1081 );
not \U$830 ( \1083 , \1082 );
not \U$831 ( \1084 , RIbe28e58_42);
not \U$832 ( \1085 , RIbe282a0_17);
nand \U$833 ( \1086 , \1085 , RIbe29470_55);
not \U$834 ( \1087 , \1086 );
not \U$835 ( \1088 , RIbe29470_55);
nand \U$836 ( \1089 , \1088 , RIbe282a0_17);
not \U$837 ( \1090 , \1089 );
or \U$838 ( \1091 , \1087 , \1090 );
xnor \U$839 ( \1092 , RIbe282a0_17, RIbe28138_14);
nand \U$840 ( \1093 , \1091 , \1092 );
not \U$841 ( \1094 , \1093 );
not \U$842 ( \1095 , \1094 );
or \U$843 ( \1096 , \1084 , \1095 );
xor \U$844 ( \1097 , RIbe282a0_17, RIbe28138_14);
buf \U$845 ( \1098 , \1097 );
buf \U$846 ( \1099 , \1098 );
nand \U$847 ( \1100 , \1099 , RIbe28de0_41);
nand \U$848 ( \1101 , \1096 , \1100 );
not \U$849 ( \1102 , \1101 );
or \U$850 ( \1103 , \1083 , \1102 );
or \U$851 ( \1104 , \1101 , \1082 );
nand \U$852 ( \1105 , \1103 , \1104 );
xor \U$853 ( \1106 , \1076 , \1105 );
xor \U$854 ( \1107 , RIbe297b8_62, RIbe29740_61);
not \U$855 ( \1108 , \1107 );
xor \U$856 ( \1109 , RIbe28138_14, RIbe297b8_62);
nand \U$857 ( \1110 , \1108 , \1109 );
not \U$858 ( \1111 , \1110 );
buf \U$859 ( \1112 , \1111 );
buf \U$860 ( \1113 , \1112 );
and \U$861 ( \1114 , \1113 , RIbe29920_65);
not \U$862 ( \1115 , \1107 );
not \U$863 ( \1116 , \1115 );
buf \U$864 ( \1117 , \1116 );
and \U$865 ( \1118 , \1117 , RIbe27b98_2);
nor \U$866 ( \1119 , \1114 , \1118 );
not \U$867 ( \1120 , RIbe29740_61);
not \U$868 ( \1121 , RIbe297b8_62);
or \U$869 ( \1122 , \1120 , \1121 );
nand \U$870 ( \1123 , \1122 , RIbe28138_14);
not \U$871 ( \1124 , \1123 );
not \U$872 ( \1125 , \1124 );
and \U$873 ( \1126 , \1119 , \1125 );
not \U$874 ( \1127 , \1119 );
and \U$875 ( \1128 , RIbe297b8_62, RIbe29740_61);
not \U$876 ( \1129 , RIbe28138_14);
nor \U$877 ( \1130 , \1128 , \1129 );
buf \U$878 ( \1131 , \1130 );
buf \U$879 ( \1132 , \1131 );
and \U$880 ( \1133 , \1127 , \1132 );
nor \U$881 ( \1134 , \1126 , \1133 );
xor \U$882 ( \1135 , \1106 , \1134 );
not \U$883 ( \1136 , \1135 );
not \U$884 ( \1137 , RIbe27d00_5);
xor \U$885 ( \1138 , RIbe294e8_56, RIbe29470_55);
not \U$886 ( \1139 , \1138 );
xor \U$887 ( \1140 , RIbe288b8_30, RIbe294e8_56);
nand \U$888 ( \1141 , \1139 , \1140 );
not \U$889 ( \1142 , \1141 );
buf \U$890 ( \1143 , \1142 );
not \U$891 ( \1144 , \1143 );
or \U$892 ( \1145 , \1137 , \1144 );
buf \U$893 ( \1146 , \1138 );
buf \U$894 ( \1147 , \1146 );
nand \U$895 ( \1148 , \1147 , RIbe27c10_3);
nand \U$896 ( \1149 , \1145 , \1148 );
nand \U$897 ( \1150 , RIbe294e8_56, RIbe29470_55);
nand \U$898 ( \1151 , \1150 , RIbe288b8_30);
buf \U$899 ( \1152 , \1151 );
buf \U$900 ( \1153 , \1152 );
not \U$901 ( \1154 , \1153 );
and \U$902 ( \1155 , \1149 , \1154 );
not \U$903 ( \1156 , \1149 );
buf \U$904 ( \1157 , \1152 );
and \U$905 ( \1158 , \1156 , \1157 );
nor \U$906 ( \1159 , \1155 , \1158 );
buf \U$907 ( \1160 , \1001 );
not \U$908 ( \1161 , \1160 );
and \U$909 ( \1162 , \1161 , RIbe29a88_68);
not \U$910 ( \1163 , \998 );
buf \U$911 ( \1164 , \1163 );
not \U$912 ( \1165 , \1164 );
and \U$913 ( \1166 , \1165 , RIbe27d78_6);
nor \U$914 ( \1167 , \1162 , \1166 );
and \U$915 ( \1168 , \1167 , \1011 );
not \U$916 ( \1169 , \1167 );
and \U$917 ( \1170 , \1169 , \752 );
nor \U$918 ( \1171 , \1168 , \1170 );
and \U$919 ( \1172 , \1159 , \1171 );
not \U$920 ( \1173 , \1159 );
not \U$921 ( \1174 , \1171 );
and \U$922 ( \1175 , \1173 , \1174 );
or \U$923 ( \1176 , \1172 , \1175 );
and \U$924 ( \1177 , \666 , RIbe28fc0_45);
xor \U$925 ( \1178 , RIbe29308_52, RIbe293f8_54);
buf \U$926 ( \1179 , \1178 );
buf \U$927 ( \1180 , \1179 );
and \U$928 ( \1181 , \1180 , RIbe290b0_47);
nor \U$929 ( \1182 , \1177 , \1181 );
and \U$930 ( \1183 , \1182 , \564 );
not \U$931 ( \1184 , \1182 );
and \U$932 ( \1185 , \1184 , \672 );
nor \U$933 ( \1186 , \1183 , \1185 );
xnor \U$934 ( \1187 , \1176 , \1186 );
nor \U$935 ( \1188 , \1136 , \1187 );
not \U$936 ( \1189 , \1188 );
not \U$937 ( \1190 , RIbe27d78_6);
not \U$938 ( \1191 , \1143 );
or \U$939 ( \1192 , \1190 , \1191 );
nand \U$940 ( \1193 , \1147 , RIbe27d00_5);
nand \U$941 ( \1194 , \1192 , \1193 );
not \U$942 ( \1195 , \1194 );
not \U$943 ( \1196 , \1153 );
and \U$944 ( \1197 , \1195 , \1196 );
and \U$945 ( \1198 , \1194 , \1153 );
nor \U$946 ( \1199 , \1197 , \1198 );
not \U$947 ( \1200 , \1199 );
and \U$948 ( \1201 , \1005 , RIbe290b0_47);
not \U$949 ( \1202 , \1163 );
buf \U$950 ( \1203 , \1202 );
and \U$951 ( \1204 , \1203 , RIbe29a88_68);
nor \U$952 ( \1205 , \1201 , \1204 );
and \U$953 ( \1206 , \1205 , \1011 );
not \U$954 ( \1207 , \1205 );
and \U$955 ( \1208 , \1207 , \752 );
nor \U$956 ( \1209 , \1206 , \1208 );
not \U$957 ( \1210 , \1209 );
and \U$958 ( \1211 , \1200 , \1210 );
and \U$959 ( \1212 , \1199 , \1209 );
and \U$960 ( \1213 , \666 , RIbe29038_46);
and \U$961 ( \1214 , \740 , RIbe28fc0_45);
nor \U$962 ( \1215 , \1213 , \1214 );
and \U$963 ( \1216 , \1215 , \672 );
not \U$964 ( \1217 , \1215 );
and \U$965 ( \1218 , \1217 , \564 );
nor \U$966 ( \1219 , \1216 , \1218 );
nor \U$967 ( \1220 , \1212 , \1219 );
nor \U$968 ( \1221 , \1211 , \1220 );
not \U$969 ( \1222 , RIbe280c0_13);
not \U$970 ( \1223 , \382 );
not \U$971 ( \1224 , \1223 );
or \U$972 ( \1225 , \1222 , \1224 );
nand \U$973 ( \1226 , \429 , RIbe29830_63);
nand \U$974 ( \1227 , \1225 , \1226 );
not \U$975 ( \1228 , \1227 );
not \U$976 ( \1229 , \313 );
and \U$977 ( \1230 , \1228 , \1229 );
not \U$978 ( \1231 , \312 );
not \U$979 ( \1232 , \1231 );
and \U$980 ( \1233 , \1227 , \1232 );
nor \U$981 ( \1234 , \1230 , \1233 );
not \U$982 ( \1235 , \1234 );
not \U$983 ( \1236 , RIbe296c8_60);
buf \U$984 ( \1237 , \546 );
not \U$985 ( \1238 , \1237 );
or \U$986 ( \1239 , \1236 , \1238 );
nand \U$987 ( \1240 , \553 , RIbe29650_59);
nand \U$988 ( \1241 , \1239 , \1240 );
not \U$989 ( \1242 , \1241 );
not \U$990 ( \1243 , \424 );
and \U$991 ( \1244 , \1242 , \1243 );
not \U$992 ( \1245 , \424 );
not \U$993 ( \1246 , \1245 );
and \U$994 ( \1247 , \1241 , \1246 );
nor \U$995 ( \1248 , \1244 , \1247 );
not \U$996 ( \1249 , \1248 );
and \U$997 ( \1250 , \1235 , \1249 );
and \U$998 ( \1251 , \1234 , \1248 );
not \U$999 ( \1252 , \281 );
not \U$1000 ( \1253 , \1252 );
not \U$1001 ( \1254 , \1253 );
and \U$1002 ( \1255 , \1254 , RIbe28228_16);
not \U$1003 ( \1256 , \286 );
and \U$1004 ( \1257 , \1256 , RIbe281b0_15);
nor \U$1005 ( \1258 , \1255 , \1257 );
and \U$1006 ( \1259 , \1258 , \293 );
not \U$1007 ( \1260 , \1258 );
and \U$1008 ( \1261 , \1260 , \300 );
nor \U$1009 ( \1262 , \1259 , \1261 );
nor \U$1010 ( \1263 , \1251 , \1262 );
nor \U$1011 ( \1264 , \1250 , \1263 );
xor \U$1012 ( \1265 , \1221 , \1264 );
nand \U$1013 ( \1266 , RIbe295d8_58, RIbe291a0_49);
or \U$1014 ( \1267 , \1266 , RIbe29740_61);
nor \U$1015 ( \1268 , RIbe295d8_58, RIbe291a0_49);
nand \U$1016 ( \1269 , \1268 , RIbe29740_61);
nand \U$1017 ( \1270 , \1267 , \1269 );
not \U$1018 ( \1271 , \1270 );
not \U$1019 ( \1272 , \1271 );
nand \U$1020 ( \1273 , \1272 , RIbe27b98_2);
and \U$1021 ( \1274 , \1266 , RIbe29740_61);
not \U$1022 ( \1275 , \1274 );
not \U$1023 ( \1276 , \1275 );
buf \U$1024 ( \1277 , \1276 );
and \U$1025 ( \1278 , \1273 , \1277 );
not \U$1026 ( \1279 , \1273 );
and \U$1027 ( \1280 , \1279 , \1076 );
nor \U$1028 ( \1281 , \1278 , \1280 );
not \U$1029 ( \1282 , \1281 );
not \U$1030 ( \1283 , \1282 );
buf \U$1031 ( \1284 , \1110 );
buf \U$1032 ( \1285 , \1284 );
not \U$1033 ( \1286 , \1285 );
and \U$1034 ( \1287 , \1286 , RIbe28de0_41);
and \U$1035 ( \1288 , \1117 , RIbe29920_65);
nor \U$1036 ( \1289 , \1287 , \1288 );
and \U$1037 ( \1290 , \1289 , \1132 );
not \U$1038 ( \1291 , \1289 );
and \U$1039 ( \1292 , \1291 , \1125 );
nor \U$1040 ( \1293 , \1290 , \1292 );
not \U$1041 ( \1294 , \1293 );
not \U$1042 ( \1295 , \1294 );
or \U$1043 ( \1296 , \1283 , \1295 );
not \U$1044 ( \1297 , RIbe27c10_3);
not \U$1045 ( \1298 , \1093 );
not \U$1046 ( \1299 , \1298 );
or \U$1047 ( \1300 , \1297 , \1299 );
nand \U$1048 ( \1301 , \1099 , RIbe28e58_42);
nand \U$1049 ( \1302 , \1300 , \1301 );
and \U$1050 ( \1303 , \1302 , \1082 );
not \U$1051 ( \1304 , \1302 );
not \U$1052 ( \1305 , RIbe282a0_17);
not \U$1053 ( \1306 , RIbe28138_14);
or \U$1054 ( \1307 , \1305 , \1306 );
nand \U$1055 ( \1308 , \1307 , RIbe29470_55);
not \U$1056 ( \1309 , \1308 );
and \U$1057 ( \1310 , \1304 , \1309 );
nor \U$1058 ( \1311 , \1303 , \1310 );
not \U$1059 ( \1312 , \1311 );
nand \U$1060 ( \1313 , \1293 , \1281 );
nand \U$1061 ( \1314 , \1312 , \1313 );
nand \U$1062 ( \1315 , \1296 , \1314 );
not \U$1063 ( \1316 , \1315 );
and \U$1064 ( \1317 , \1265 , \1316 );
and \U$1065 ( \1318 , \1221 , \1264 );
or \U$1066 ( \1319 , \1317 , \1318 );
not \U$1067 ( \1320 , \1319 );
not \U$1068 ( \1321 , \1320 );
or \U$1069 ( \1322 , \1189 , \1321 );
or \U$1070 ( \1323 , \1320 , \1188 );
not \U$1071 ( \1324 , RIbe29650_59);
not \U$1072 ( \1325 , \1237 );
or \U$1073 ( \1326 , \1324 , \1325 );
buf \U$1074 ( \1327 , \552 );
nand \U$1075 ( \1328 , \1327 , RIbe29038_46);
nand \U$1076 ( \1329 , \1326 , \1328 );
not \U$1077 ( \1330 , \424 );
and \U$1078 ( \1331 , \1329 , \1330 );
not \U$1079 ( \1332 , \1329 );
not \U$1080 ( \1333 , \1330 );
and \U$1081 ( \1334 , \1332 , \1333 );
nor \U$1082 ( \1335 , \1331 , \1334 );
not \U$1083 ( \1336 , RIbe29830_63);
not \U$1084 ( \1337 , \382 );
not \U$1085 ( \1338 , \1337 );
or \U$1086 ( \1339 , \1336 , \1338 );
nand \U$1087 ( \1340 , \429 , RIbe296c8_60);
nand \U$1088 ( \1341 , \1339 , \1340 );
and \U$1089 ( \1342 , \1341 , \313 );
not \U$1090 ( \1343 , \1341 );
and \U$1091 ( \1344 , \1343 , \306 );
nor \U$1092 ( \1345 , \1342 , \1344 );
xor \U$1093 ( \1346 , \1335 , \1345 );
and \U$1094 ( \1347 , \1254 , RIbe281b0_15);
and \U$1095 ( \1348 , \287 , RIbe280c0_13);
nor \U$1096 ( \1349 , \1347 , \1348 );
and \U$1097 ( \1350 , \1349 , \293 );
not \U$1098 ( \1351 , \1349 );
and \U$1099 ( \1352 , \1351 , \300 );
nor \U$1100 ( \1353 , \1350 , \1352 );
xnor \U$1101 ( \1354 , \1346 , \1353 );
nand \U$1102 ( \1355 , RIbe29380_53, RIbe29290_51);
not \U$1103 ( \1356 , \260 );
not \U$1104 ( \1357 , \1356 );
and \U$1105 ( \1358 , \1357 , RIbe28930_31);
and \U$1106 ( \1359 , \264 , RIbe29560_57);
nor \U$1107 ( \1360 , \1358 , \1359 );
nand \U$1108 ( \1361 , \267 , RIbe27ee0_9);
buf \U$1109 ( \1362 , \1361 );
not \U$1110 ( \1363 , \1362 );
and \U$1111 ( \1364 , \1360 , \1363 );
not \U$1112 ( \1365 , \1360 );
and \U$1113 ( \1366 , \1365 , \270 );
nor \U$1114 ( \1367 , \1364 , \1366 );
xor \U$1115 ( \1368 , \1355 , \1367 );
and \U$1116 ( \1369 , \326 , RIbe28a20_33);
not \U$1117 ( \1370 , \329 );
not \U$1118 ( \1371 , \1370 );
and \U$1119 ( \1372 , \1371 , RIbe289a8_32);
nor \U$1120 ( \1373 , \1369 , \1372 );
buf \U$1121 ( \1374 , \337 );
not \U$1122 ( \1375 , \1374 );
and \U$1123 ( \1376 , \1373 , \1375 );
not \U$1124 ( \1377 , \1373 );
not \U$1125 ( \1378 , \337 );
not \U$1126 ( \1379 , \1378 );
and \U$1127 ( \1380 , \1377 , \1379 );
nor \U$1128 ( \1381 , \1376 , \1380 );
and \U$1129 ( \1382 , \1368 , \1381 );
and \U$1130 ( \1383 , \1355 , \1367 );
or \U$1131 ( \1384 , \1382 , \1383 );
xor \U$1132 ( \1385 , \1354 , \1384 );
and \U$1133 ( \1386 , \326 , RIbe289a8_32);
and \U$1134 ( \1387 , \1371 , RIbe28930_31);
nor \U$1135 ( \1388 , \1386 , \1387 );
and \U$1136 ( \1389 , \1388 , \1378 );
not \U$1137 ( \1390 , \1388 );
and \U$1138 ( \1391 , \1390 , \1374 );
nor \U$1139 ( \1392 , \1389 , \1391 );
not \U$1140 ( \1393 , RIbe29560_57);
not \U$1141 ( \1394 , \261 );
or \U$1142 ( \1395 , \1393 , \1394 );
nand \U$1143 ( \1396 , \264 , RIbe28228_16);
nand \U$1144 ( \1397 , \1395 , \1396 );
not \U$1145 ( \1398 , \1397 );
not \U$1146 ( \1399 , \1362 );
and \U$1147 ( \1400 , \1398 , \1399 );
and \U$1148 ( \1401 , \1397 , \1362 );
nor \U$1149 ( \1402 , \1400 , \1401 );
and \U$1150 ( \1403 , \1392 , \1402 );
not \U$1151 ( \1404 , \1392 );
not \U$1152 ( \1405 , \1402 );
and \U$1153 ( \1406 , \1404 , \1405 );
nor \U$1154 ( \1407 , \1403 , \1406 );
nand \U$1155 ( \1408 , RIbe29380_53, RIbe28a20_33);
and \U$1156 ( \1409 , \1407 , \1408 );
nor \U$1157 ( \1410 , \1407 , \1408 );
nor \U$1158 ( \1411 , \1409 , \1410 );
and \U$1159 ( \1412 , \1385 , \1411 );
and \U$1160 ( \1413 , \1354 , \1384 );
or \U$1161 ( \1414 , \1412 , \1413 );
not \U$1162 ( \1415 , \1414 );
nand \U$1163 ( \1416 , \1323 , \1415 );
nand \U$1164 ( \1417 , \1322 , \1416 );
not \U$1165 ( \1418 , \1417 );
not \U$1166 ( \1419 , RIbe29038_46);
not \U$1167 ( \1420 , \1237 );
or \U$1168 ( \1421 , \1419 , \1420 );
nand \U$1169 ( \1422 , \552 , RIbe28fc0_45);
nand \U$1170 ( \1423 , \1421 , \1422 );
and \U$1171 ( \1424 , \1423 , \425 );
not \U$1172 ( \1425 , \1423 );
and \U$1173 ( \1426 , \1425 , \1333 );
nor \U$1174 ( \1427 , \1424 , \1426 );
and \U$1175 ( \1428 , \664 , RIbe290b0_47);
and \U$1176 ( \1429 , \1180 , RIbe29a88_68);
nor \U$1177 ( \1430 , \1428 , \1429 );
and \U$1178 ( \1431 , \1430 , \564 );
not \U$1179 ( \1432 , \1430 );
and \U$1180 ( \1433 , \1432 , \672 );
nor \U$1181 ( \1434 , \1431 , \1433 );
xor \U$1182 ( \1435 , \1427 , \1434 );
and \U$1183 ( \1436 , \1005 , RIbe27d78_6);
and \U$1184 ( \1437 , \1203 , RIbe27d00_5);
nor \U$1185 ( \1438 , \1436 , \1437 );
and \U$1186 ( \1439 , \1438 , \752 );
not \U$1187 ( \1440 , \1438 );
and \U$1188 ( \1441 , \1440 , \1011 );
nor \U$1189 ( \1442 , \1439 , \1441 );
xor \U$1190 ( \1443 , \1435 , \1442 );
not \U$1191 ( \1444 , \1443 );
nand \U$1192 ( \1445 , \1113 , RIbe27b98_2);
and \U$1193 ( \1446 , \1445 , \1132 );
not \U$1194 ( \1447 , \1445 );
not \U$1195 ( \1448 , \1124 );
and \U$1196 ( \1449 , \1447 , \1448 );
or \U$1197 ( \1450 , \1446 , \1449 );
not \U$1198 ( \1451 , RIbe28de0_41);
not \U$1199 ( \1452 , \1298 );
or \U$1200 ( \1453 , \1451 , \1452 );
buf \U$1201 ( \1454 , \1098 );
buf \U$1202 ( \1455 , \1454 );
nand \U$1203 ( \1456 , \1455 , RIbe29920_65);
nand \U$1204 ( \1457 , \1453 , \1456 );
not \U$1205 ( \1458 , \1081 );
and \U$1206 ( \1459 , \1457 , \1458 );
not \U$1207 ( \1460 , \1457 );
and \U$1208 ( \1461 , \1460 , \1309 );
nor \U$1209 ( \1462 , \1459 , \1461 );
xor \U$1210 ( \1463 , \1450 , \1462 );
and \U$1211 ( \1464 , \1143 , RIbe27c10_3);
and \U$1212 ( \1465 , \1147 , RIbe28e58_42);
nor \U$1213 ( \1466 , \1464 , \1465 );
and \U$1214 ( \1467 , \1466 , \1153 );
not \U$1215 ( \1468 , \1466 );
not \U$1216 ( \1469 , \1157 );
and \U$1217 ( \1470 , \1468 , \1469 );
or \U$1218 ( \1471 , \1467 , \1470 );
xnor \U$1219 ( \1472 , \1463 , \1471 );
not \U$1220 ( \1473 , \1472 );
or \U$1221 ( \1474 , \1444 , \1473 );
or \U$1222 ( \1475 , \1472 , \1443 );
nand \U$1223 ( \1476 , \1474 , \1475 );
not \U$1224 ( \1477 , \1476 );
xor \U$1225 ( \1478 , \1076 , \1105 );
and \U$1226 ( \1479 , \1478 , \1134 );
and \U$1227 ( \1480 , \1076 , \1105 );
or \U$1228 ( \1481 , \1479 , \1480 );
nand \U$1229 ( \1482 , \1345 , \1353 );
and \U$1230 ( \1483 , \1482 , \1335 );
nor \U$1231 ( \1484 , \1345 , \1353 );
nor \U$1232 ( \1485 , \1483 , \1484 );
xnor \U$1233 ( \1486 , \1481 , \1485 );
not \U$1234 ( \1487 , \1174 );
not \U$1235 ( \1488 , \1159 );
or \U$1236 ( \1489 , \1487 , \1488 );
or \U$1237 ( \1490 , \1159 , \1174 );
nand \U$1238 ( \1491 , \1490 , \1186 );
nand \U$1239 ( \1492 , \1489 , \1491 );
xor \U$1240 ( \1493 , \1486 , \1492 );
not \U$1241 ( \1494 , \1493 );
or \U$1242 ( \1495 , \1477 , \1494 );
or \U$1243 ( \1496 , \1493 , \1476 );
or \U$1244 ( \1497 , \1392 , \1408 );
not \U$1245 ( \1498 , \1408 );
not \U$1246 ( \1499 , \1392 );
or \U$1247 ( \1500 , \1498 , \1499 );
nand \U$1248 ( \1501 , \1500 , \1405 );
nand \U$1249 ( \1502 , \1497 , \1501 );
and \U$1250 ( \1503 , \326 , RIbe28930_31);
and \U$1251 ( \1504 , \329 , RIbe29560_57);
nor \U$1252 ( \1505 , \1503 , \1504 );
and \U$1253 ( \1506 , \1505 , \1375 );
not \U$1254 ( \1507 , \1505 );
and \U$1255 ( \1508 , \1507 , \1379 );
nor \U$1256 ( \1509 , \1506 , \1508 );
nand \U$1257 ( \1510 , RIbe29380_53, RIbe289a8_32);
or \U$1258 ( \1511 , \1509 , \1510 );
nand \U$1259 ( \1512 , \1509 , \1510 );
nand \U$1260 ( \1513 , \1511 , \1512 );
xor \U$1261 ( \1514 , \1502 , \1513 );
not \U$1262 ( \1515 , RIbe28228_16);
not \U$1263 ( \1516 , \1356 );
not \U$1264 ( \1517 , \1516 );
or \U$1265 ( \1518 , \1515 , \1517 );
nand \U$1266 ( \1519 , \263 , RIbe281b0_15);
nand \U$1267 ( \1520 , \1518 , \1519 );
not \U$1268 ( \1521 , \1520 );
not \U$1269 ( \1522 , \1362 );
and \U$1270 ( \1523 , \1521 , \1522 );
and \U$1271 ( \1524 , \1520 , \270 );
nor \U$1272 ( \1525 , \1523 , \1524 );
not \U$1273 ( \1526 , \1525 );
not \U$1274 ( \1527 , RIbe280c0_13);
buf \U$1275 ( \1528 , \1252 );
not \U$1276 ( \1529 , \1528 );
or \U$1277 ( \1530 , \1527 , \1529 );
not \U$1278 ( \1531 , \286 );
nand \U$1279 ( \1532 , \1531 , RIbe29830_63);
nand \U$1280 ( \1533 , \1530 , \1532 );
not \U$1281 ( \1534 , \1533 );
not \U$1282 ( \1535 , \300 );
and \U$1283 ( \1536 , \1534 , \1535 );
and \U$1284 ( \1537 , \1533 , \300 );
nor \U$1285 ( \1538 , \1536 , \1537 );
not \U$1286 ( \1539 , \1538 );
not \U$1287 ( \1540 , RIbe296c8_60);
not \U$1288 ( \1541 , \1223 );
or \U$1289 ( \1542 , \1540 , \1541 );
nand \U$1290 ( \1543 , \429 , RIbe29650_59);
nand \U$1291 ( \1544 , \1542 , \1543 );
and \U$1292 ( \1545 , \1544 , \306 );
not \U$1293 ( \1546 , \1544 );
not \U$1294 ( \1547 , \1231 );
and \U$1295 ( \1548 , \1546 , \1547 );
nor \U$1296 ( \1549 , \1545 , \1548 );
not \U$1297 ( \1550 , \1549 );
or \U$1298 ( \1551 , \1539 , \1550 );
or \U$1299 ( \1552 , \1549 , \1538 );
nand \U$1300 ( \1553 , \1551 , \1552 );
not \U$1301 ( \1554 , \1553 );
or \U$1302 ( \1555 , \1526 , \1554 );
or \U$1303 ( \1556 , \1553 , \1525 );
nand \U$1304 ( \1557 , \1555 , \1556 );
xor \U$1305 ( \1558 , \1514 , \1557 );
nand \U$1306 ( \1559 , \1496 , \1558 );
nand \U$1307 ( \1560 , \1495 , \1559 );
not \U$1308 ( \1561 , \1560 );
or \U$1309 ( \1562 , \1418 , \1561 );
or \U$1310 ( \1563 , \1560 , \1417 );
xor \U$1311 ( \1564 , \1427 , \1434 );
and \U$1312 ( \1565 , \1564 , \1442 );
and \U$1313 ( \1566 , \1427 , \1434 );
or \U$1314 ( \1567 , \1565 , \1566 );
nand \U$1315 ( \1568 , \1538 , \1525 );
not \U$1316 ( \1569 , \1568 );
not \U$1317 ( \1570 , \1549 );
or \U$1318 ( \1571 , \1569 , \1570 );
or \U$1319 ( \1572 , \1525 , \1538 );
nand \U$1320 ( \1573 , \1571 , \1572 );
xor \U$1321 ( \1574 , \1567 , \1573 );
or \U$1322 ( \1575 , \1471 , \1462 );
not \U$1323 ( \1576 , \1471 );
not \U$1324 ( \1577 , \1462 );
or \U$1325 ( \1578 , \1576 , \1577 );
nand \U$1326 ( \1579 , \1578 , \1450 );
nand \U$1327 ( \1580 , \1575 , \1579 );
xor \U$1328 ( \1581 , \1574 , \1580 );
and \U$1329 ( \1582 , \327 , RIbe29560_57);
and \U$1330 ( \1583 , \331 , RIbe28228_16);
nor \U$1331 ( \1584 , \1582 , \1583 );
and \U$1332 ( \1585 , \1584 , \339 );
not \U$1333 ( \1586 , \1584 );
and \U$1334 ( \1587 , \1586 , \342 );
nor \U$1335 ( \1588 , \1585 , \1587 );
and \U$1336 ( \1589 , RIbe28930_31, RIbe29380_53);
xor \U$1337 ( \1590 , \1588 , \1589 );
xor \U$1338 ( \1591 , \1590 , \1512 );
not \U$1339 ( \1592 , RIbe28fc0_45);
not \U$1340 ( \1593 , \548 );
or \U$1341 ( \1594 , \1592 , \1593 );
nand \U$1342 ( \1595 , \554 , RIbe290b0_47);
nand \U$1343 ( \1596 , \1594 , \1595 );
not \U$1344 ( \1597 , \1596 );
not \U$1345 ( \1598 , \424 );
and \U$1346 ( \1599 , \1597 , \1598 );
and \U$1347 ( \1600 , \1596 , \424 );
nor \U$1348 ( \1601 , \1599 , \1600 );
not \U$1349 ( \1602 , \1601 );
and \U$1350 ( \1603 , \1161 , RIbe27d00_5);
and \U$1351 ( \1604 , \1165 , RIbe27c10_3);
nor \U$1352 ( \1605 , \1603 , \1604 );
and \U$1353 ( \1606 , \1605 , \1011 );
not \U$1354 ( \1607 , \1605 );
not \U$1355 ( \1608 , \751 );
and \U$1356 ( \1609 , \1607 , \1608 );
nor \U$1357 ( \1610 , \1606 , \1609 );
not \U$1358 ( \1611 , \1180 );
not \U$1359 ( \1612 , \1611 );
not \U$1360 ( \1613 , \255 );
and \U$1361 ( \1614 , \1612 , \1613 );
and \U$1362 ( \1615 , \664 , RIbe29a88_68);
nor \U$1363 ( \1616 , \1614 , \1615 );
not \U$1364 ( \1617 , \563 );
not \U$1365 ( \1618 , \1617 );
and \U$1366 ( \1619 , \1616 , \1618 );
not \U$1367 ( \1620 , \1616 );
not \U$1368 ( \1621 , \671 );
and \U$1369 ( \1622 , \1620 , \1621 );
nor \U$1370 ( \1623 , \1619 , \1622 );
xnor \U$1371 ( \1624 , \1610 , \1623 );
not \U$1372 ( \1625 , \1624 );
or \U$1373 ( \1626 , \1602 , \1625 );
or \U$1374 ( \1627 , \1624 , \1601 );
nand \U$1375 ( \1628 , \1626 , \1627 );
nand \U$1376 ( \1629 , \1086 , \1089 );
nand \U$1377 ( \1630 , \1092 , \1629 );
not \U$1378 ( \1631 , \1630 );
buf \U$1379 ( \1632 , \1631 );
buf \U$1380 ( \1633 , \1632 );
not \U$1381 ( \1634 , \1633 );
not \U$1382 ( \1635 , \1634 );
not \U$1383 ( \1636 , RIbe29920_65);
not \U$1384 ( \1637 , \1636 );
and \U$1385 ( \1638 , \1635 , \1637 );
not \U$1386 ( \1639 , \1099 );
not \U$1387 ( \1640 , RIbe27b98_2);
nor \U$1388 ( \1641 , \1639 , \1640 );
nor \U$1389 ( \1642 , \1638 , \1641 );
and \U$1390 ( \1643 , \1642 , \1458 );
not \U$1391 ( \1644 , \1642 );
and \U$1392 ( \1645 , \1644 , \1309 );
nor \U$1393 ( \1646 , \1643 , \1645 );
and \U$1394 ( \1647 , \1143 , RIbe28e58_42);
and \U$1395 ( \1648 , \1147 , RIbe28de0_41);
nor \U$1396 ( \1649 , \1647 , \1648 );
and \U$1397 ( \1650 , \1649 , \1157 );
not \U$1398 ( \1651 , \1649 );
not \U$1399 ( \1652 , \1152 );
and \U$1400 ( \1653 , \1651 , \1652 );
nor \U$1401 ( \1654 , \1650 , \1653 );
xor \U$1402 ( \1655 , \1646 , \1654 );
xor \U$1403 ( \1656 , \1655 , \1125 );
xor \U$1404 ( \1657 , \1628 , \1656 );
not \U$1405 ( \1658 , \260 );
not \U$1406 ( \1659 , \1658 );
and \U$1407 ( \1660 , \1659 , RIbe281b0_15);
and \U$1408 ( \1661 , \264 , RIbe280c0_13);
nor \U$1409 ( \1662 , \1660 , \1661 );
not \U$1410 ( \1663 , \1362 );
and \U$1411 ( \1664 , \1662 , \1663 );
not \U$1412 ( \1665 , \1662 );
and \U$1413 ( \1666 , \1665 , \1362 );
nor \U$1414 ( \1667 , \1664 , \1666 );
not \U$1415 ( \1668 , \1667 );
not \U$1416 ( \1669 , RIbe29650_59);
not \U$1417 ( \1670 , \1223 );
or \U$1418 ( \1671 , \1669 , \1670 );
nand \U$1419 ( \1672 , \429 , RIbe29038_46);
nand \U$1420 ( \1673 , \1671 , \1672 );
not \U$1421 ( \1674 , \1673 );
not \U$1422 ( \1675 , \313 );
and \U$1423 ( \1676 , \1674 , \1675 );
and \U$1424 ( \1677 , \1673 , \1547 );
nor \U$1425 ( \1678 , \1676 , \1677 );
not \U$1426 ( \1679 , \282 );
and \U$1427 ( \1680 , \1679 , RIbe29830_63);
not \U$1428 ( \1681 , \285 );
buf \U$1429 ( \1682 , \1681 );
and \U$1430 ( \1683 , \1682 , RIbe296c8_60);
nor \U$1431 ( \1684 , \1680 , \1683 );
and \U$1432 ( \1685 , \1684 , \293 );
not \U$1433 ( \1686 , \1684 );
and \U$1434 ( \1687 , \1686 , \300 );
nor \U$1435 ( \1688 , \1685 , \1687 );
xor \U$1436 ( \1689 , \1678 , \1688 );
not \U$1437 ( \1690 , \1689 );
or \U$1438 ( \1691 , \1668 , \1690 );
or \U$1439 ( \1692 , \1689 , \1667 );
nand \U$1440 ( \1693 , \1691 , \1692 );
xor \U$1441 ( \1694 , \1657 , \1693 );
xor \U$1442 ( \1695 , \1591 , \1694 );
xor \U$1443 ( \1696 , \1581 , \1695 );
nand \U$1444 ( \1697 , \1563 , \1696 );
nand \U$1445 ( \1698 , \1562 , \1697 );
xor \U$1446 ( \1699 , \1567 , \1573 );
and \U$1447 ( \1700 , \1699 , \1580 );
and \U$1448 ( \1701 , \1567 , \1573 );
or \U$1449 ( \1702 , \1700 , \1701 );
xor \U$1450 ( \1703 , \1588 , \1589 );
and \U$1451 ( \1704 , \1703 , \1512 );
and \U$1452 ( \1705 , \1588 , \1589 );
or \U$1453 ( \1706 , \1704 , \1705 );
xor \U$1454 ( \1707 , \1702 , \1706 );
xor \U$1455 ( \1708 , \1628 , \1656 );
and \U$1456 ( \1709 , \1708 , \1693 );
and \U$1457 ( \1710 , \1628 , \1656 );
or \U$1458 ( \1711 , \1709 , \1710 );
xor \U$1459 ( \1712 , \1707 , \1711 );
and \U$1460 ( \1713 , \1698 , \1712 );
or \U$1461 ( \1714 , \1698 , \1712 );
xor \U$1462 ( \1715 , \1567 , \1573 );
xor \U$1463 ( \1716 , \1715 , \1580 );
and \U$1464 ( \1717 , \1591 , \1716 );
xor \U$1465 ( \1718 , \1567 , \1573 );
xor \U$1466 ( \1719 , \1718 , \1580 );
and \U$1467 ( \1720 , \1694 , \1719 );
and \U$1468 ( \1721 , \1591 , \1694 );
or \U$1469 ( \1722 , \1717 , \1720 , \1721 );
and \U$1470 ( \1723 , \1481 , \1492 );
not \U$1471 ( \1724 , \1492 );
not \U$1472 ( \1725 , \1481 );
and \U$1473 ( \1726 , \1724 , \1725 );
nor \U$1474 ( \1727 , \1726 , \1485 );
nor \U$1475 ( \1728 , \1723 , \1727 );
not \U$1476 ( \1729 , \1472 );
nand \U$1477 ( \1730 , \1729 , \1443 );
or \U$1478 ( \1731 , \1728 , \1730 );
not \U$1479 ( \1732 , \1730 );
not \U$1480 ( \1733 , \1728 );
or \U$1481 ( \1734 , \1732 , \1733 );
xor \U$1482 ( \1735 , \1502 , \1513 );
and \U$1483 ( \1736 , \1735 , \1557 );
and \U$1484 ( \1737 , \1502 , \1513 );
or \U$1485 ( \1738 , \1736 , \1737 );
nand \U$1486 ( \1739 , \1734 , \1738 );
nand \U$1487 ( \1740 , \1731 , \1739 );
xor \U$1488 ( \1741 , \1722 , \1740 );
not \U$1489 ( \1742 , RIbe27d78_6);
not \U$1490 ( \1743 , \663 );
not \U$1491 ( \1744 , \1743 );
not \U$1492 ( \1745 , \1744 );
or \U$1493 ( \1746 , \1742 , \1745 );
nand \U$1494 ( \1747 , \740 , RIbe27d00_5);
nand \U$1495 ( \1748 , \1746 , \1747 );
not \U$1496 ( \1749 , \1748 );
not \U$1497 ( \1750 , \564 );
and \U$1498 ( \1751 , \1749 , \1750 );
and \U$1499 ( \1752 , \1748 , \1618 );
nor \U$1500 ( \1753 , \1751 , \1752 );
not \U$1501 ( \1754 , \1753 );
not \U$1502 ( \1755 , RIbe290b0_47);
buf \U$1503 ( \1756 , \546 );
not \U$1504 ( \1757 , \1756 );
or \U$1505 ( \1758 , \1755 , \1757 );
nand \U$1506 ( \1759 , \554 , RIbe29a88_68);
nand \U$1507 ( \1760 , \1758 , \1759 );
not \U$1508 ( \1761 , \424 );
and \U$1509 ( \1762 , \1760 , \1761 );
not \U$1510 ( \1763 , \1760 );
not \U$1511 ( \1764 , \1761 );
and \U$1512 ( \1765 , \1763 , \1764 );
nor \U$1513 ( \1766 , \1762 , \1765 );
not \U$1514 ( \1767 , \1766 );
or \U$1515 ( \1768 , \1754 , \1767 );
or \U$1516 ( \1769 , \1753 , \1766 );
nand \U$1517 ( \1770 , \1768 , \1769 );
not \U$1518 ( \1771 , \1770 );
not \U$1519 ( \1772 , RIbe29038_46);
not \U$1520 ( \1773 , \382 );
buf \U$1521 ( \1774 , \1773 );
not \U$1522 ( \1775 , \1774 );
or \U$1523 ( \1776 , \1772 , \1775 );
nand \U$1524 ( \1777 , \429 , RIbe28fc0_45);
nand \U$1525 ( \1778 , \1776 , \1777 );
and \U$1526 ( \1779 , \1778 , \306 );
not \U$1527 ( \1780 , \1778 );
and \U$1528 ( \1781 , \1780 , \313 );
or \U$1529 ( \1782 , \1779 , \1781 );
not \U$1530 ( \1783 , \1782 );
and \U$1531 ( \1784 , \1771 , \1783 );
and \U$1532 ( \1785 , \1770 , \1782 );
nor \U$1533 ( \1786 , \1784 , \1785 );
not \U$1534 ( \1787 , RIbe28de0_41);
not \U$1535 ( \1788 , \1143 );
or \U$1536 ( \1789 , \1787 , \1788 );
nand \U$1537 ( \1790 , \1147 , RIbe29920_65);
nand \U$1538 ( \1791 , \1789 , \1790 );
and \U$1539 ( \1792 , \1791 , \1157 );
not \U$1540 ( \1793 , \1791 );
not \U$1541 ( \1794 , \1153 );
and \U$1542 ( \1795 , \1793 , \1794 );
nor \U$1543 ( \1796 , \1792 , \1795 );
not \U$1544 ( \1797 , \1309 );
not \U$1545 ( \1798 , \1634 );
nand \U$1546 ( \1799 , \1798 , RIbe27b98_2);
not \U$1547 ( \1800 , \1799 );
or \U$1548 ( \1801 , \1797 , \1800 );
or \U$1549 ( \1802 , \1799 , \1309 );
nand \U$1550 ( \1803 , \1801 , \1802 );
xnor \U$1551 ( \1804 , \1796 , \1803 );
not \U$1552 ( \1805 , RIbe27c10_3);
not \U$1553 ( \1806 , \1001 );
buf \U$1554 ( \1807 , \1806 );
not \U$1555 ( \1808 , \1807 );
or \U$1556 ( \1809 , \1805 , \1808 );
nand \U$1557 ( \1810 , \1203 , RIbe28e58_42);
nand \U$1558 ( \1811 , \1809 , \1810 );
not \U$1559 ( \1812 , \1811 );
buf \U$1560 ( \1813 , \750 );
not \U$1561 ( \1814 , \1813 );
and \U$1562 ( \1815 , \1812 , \1814 );
and \U$1563 ( \1816 , \1811 , \752 );
nor \U$1564 ( \1817 , \1815 , \1816 );
xor \U$1565 ( \1818 , \1804 , \1817 );
xor \U$1566 ( \1819 , \1786 , \1818 );
and \U$1567 ( \1820 , \1254 , RIbe296c8_60);
and \U$1568 ( \1821 , \1256 , RIbe29650_59);
nor \U$1569 ( \1822 , \1820 , \1821 );
and \U$1570 ( \1823 , \1822 , \300 );
not \U$1571 ( \1824 , \1822 );
and \U$1572 ( \1825 , \1824 , \293 );
nor \U$1573 ( \1826 , \1823 , \1825 );
not \U$1574 ( \1827 , \1826 );
not \U$1575 ( \1828 , \1827 );
and \U$1576 ( \1829 , \1516 , RIbe280c0_13);
not \U$1577 ( \1830 , \263 );
not \U$1578 ( \1831 , \1830 );
and \U$1579 ( \1832 , \1831 , RIbe29830_63);
nor \U$1580 ( \1833 , \1829 , \1832 );
and \U$1581 ( \1834 , \1833 , \268 );
not \U$1582 ( \1835 , \1833 );
and \U$1583 ( \1836 , \1835 , \1362 );
nor \U$1584 ( \1837 , \1834 , \1836 );
not \U$1585 ( \1838 , \1837 );
not \U$1586 ( \1839 , \1838 );
or \U$1587 ( \1840 , \1828 , \1839 );
nand \U$1588 ( \1841 , \1837 , \1826 );
nand \U$1589 ( \1842 , \1840 , \1841 );
not \U$1590 ( \1843 , \1842 );
and \U$1591 ( \1844 , \326 , RIbe28228_16);
and \U$1592 ( \1845 , \1371 , RIbe281b0_15);
nor \U$1593 ( \1846 , \1844 , \1845 );
and \U$1594 ( \1847 , \1846 , \342 );
not \U$1595 ( \1848 , \1846 );
and \U$1596 ( \1849 , \1848 , \1379 );
nor \U$1597 ( \1850 , \1847 , \1849 );
not \U$1598 ( \1851 , \1850 );
and \U$1599 ( \1852 , \1843 , \1851 );
and \U$1600 ( \1853 , \1842 , \1850 );
nor \U$1601 ( \1854 , \1852 , \1853 );
nand \U$1602 ( \1855 , RIbe29380_53, RIbe29560_57);
or \U$1603 ( \1856 , \1854 , \1855 );
nand \U$1604 ( \1857 , \1854 , \1855 );
nand \U$1605 ( \1858 , \1856 , \1857 );
xor \U$1606 ( \1859 , \1819 , \1858 );
or \U$1607 ( \1860 , \1678 , \1688 );
not \U$1608 ( \1861 , \1688 );
not \U$1609 ( \1862 , \1678 );
or \U$1610 ( \1863 , \1861 , \1862 );
not \U$1611 ( \1864 , \1667 );
nand \U$1612 ( \1865 , \1863 , \1864 );
nand \U$1613 ( \1866 , \1860 , \1865 );
nand \U$1614 ( \1867 , \1610 , \1601 );
not \U$1615 ( \1868 , \1867 );
not \U$1616 ( \1869 , \1623 );
or \U$1617 ( \1870 , \1868 , \1869 );
or \U$1618 ( \1871 , \1610 , \1601 );
nand \U$1619 ( \1872 , \1870 , \1871 );
xor \U$1620 ( \1873 , \1866 , \1872 );
xor \U$1621 ( \1874 , \1646 , \1654 );
and \U$1622 ( \1875 , \1874 , \1125 );
and \U$1623 ( \1876 , \1646 , \1654 );
or \U$1624 ( \1877 , \1875 , \1876 );
xor \U$1625 ( \1878 , \1873 , \1877 );
xor \U$1626 ( \1879 , \1859 , \1878 );
xor \U$1627 ( \1880 , \1741 , \1879 );
and \U$1628 ( \1881 , \1714 , \1880 );
nor \U$1629 ( \1882 , \1713 , \1881 );
not \U$1630 ( \1883 , \1882 );
xor \U$1631 ( \1884 , \1722 , \1740 );
and \U$1632 ( \1885 , \1884 , \1879 );
and \U$1633 ( \1886 , \1722 , \1740 );
or \U$1634 ( \1887 , \1885 , \1886 );
xor \U$1635 ( \1888 , \1866 , \1872 );
and \U$1636 ( \1889 , \1888 , \1877 );
and \U$1637 ( \1890 , \1866 , \1872 );
or \U$1638 ( \1891 , \1889 , \1890 );
not \U$1639 ( \1892 , \1891 );
nor \U$1640 ( \1893 , \1818 , \1786 );
xnor \U$1641 ( \1894 , \1893 , \1857 );
not \U$1642 ( \1895 , \1894 );
or \U$1643 ( \1896 , \1892 , \1895 );
or \U$1644 ( \1897 , \1894 , \1891 );
nand \U$1645 ( \1898 , \1896 , \1897 );
xor \U$1646 ( \1899 , \1887 , \1898 );
xor \U$1647 ( \1900 , \1702 , \1706 );
and \U$1648 ( \1901 , \1900 , \1711 );
and \U$1649 ( \1902 , \1702 , \1706 );
or \U$1650 ( \1903 , \1901 , \1902 );
xor \U$1651 ( \1904 , \1819 , \1858 );
and \U$1652 ( \1905 , \1904 , \1878 );
and \U$1653 ( \1906 , \1819 , \1858 );
or \U$1654 ( \1907 , \1905 , \1906 );
xor \U$1655 ( \1908 , \1903 , \1907 );
not \U$1656 ( \1909 , RIbe29a88_68);
not \U$1657 ( \1910 , \1756 );
or \U$1658 ( \1911 , \1909 , \1910 );
nand \U$1659 ( \1912 , \554 , RIbe27d78_6);
nand \U$1660 ( \1913 , \1911 , \1912 );
and \U$1661 ( \1914 , \1913 , \1330 );
not \U$1662 ( \1915 , \1913 );
and \U$1663 ( \1916 , \1915 , \424 );
nor \U$1664 ( \1917 , \1914 , \1916 );
not \U$1665 ( \1918 , \564 );
not \U$1666 ( \1919 , RIbe27d00_5);
not \U$1667 ( \1920 , \1744 );
or \U$1668 ( \1921 , \1919 , \1920 );
nand \U$1669 ( \1922 , \740 , RIbe27c10_3);
nand \U$1670 ( \1923 , \1921 , \1922 );
not \U$1671 ( \1924 , \1923 );
or \U$1672 ( \1925 , \1918 , \1924 );
or \U$1673 ( \1926 , \1923 , \564 );
nand \U$1674 ( \1927 , \1925 , \1926 );
xor \U$1675 ( \1928 , \1917 , \1927 );
not \U$1676 ( \1929 , \1928 );
not \U$1677 ( \1930 , \382 );
not \U$1678 ( \1931 , RIbe28fc0_45);
not \U$1679 ( \1932 , \1931 );
and \U$1680 ( \1933 , \1930 , \1932 );
and \U$1681 ( \1934 , \429 , RIbe290b0_47);
nor \U$1682 ( \1935 , \1933 , \1934 );
and \U$1683 ( \1936 , \1935 , \306 );
not \U$1684 ( \1937 , \1935 );
and \U$1685 ( \1938 , \1937 , \313 );
nor \U$1686 ( \1939 , \1936 , \1938 );
not \U$1687 ( \1940 , \1939 );
and \U$1688 ( \1941 , \1929 , \1940 );
and \U$1689 ( \1942 , \1928 , \1939 );
nor \U$1690 ( \1943 , \1941 , \1942 );
nand \U$1691 ( \1944 , RIbe29380_53, RIbe28228_16);
xor \U$1692 ( \1945 , \1943 , \1944 );
and \U$1693 ( \1946 , \1516 , RIbe29830_63);
and \U$1694 ( \1947 , \1831 , RIbe296c8_60);
nor \U$1695 ( \1948 , \1946 , \1947 );
and \U$1696 ( \1949 , \1948 , \1363 );
not \U$1697 ( \1950 , \1948 );
and \U$1698 ( \1951 , \1950 , \1362 );
nor \U$1699 ( \1952 , \1949 , \1951 );
not \U$1700 ( \1953 , \1952 );
and \U$1701 ( \1954 , \1254 , RIbe29650_59);
and \U$1702 ( \1955 , \1256 , RIbe29038_46);
nor \U$1703 ( \1956 , \1954 , \1955 );
and \U$1704 ( \1957 , \1956 , \300 );
not \U$1705 ( \1958 , \1956 );
and \U$1706 ( \1959 , \1958 , \293 );
nor \U$1707 ( \1960 , \1957 , \1959 );
not \U$1708 ( \1961 , \1960 );
or \U$1709 ( \1962 , \1953 , \1961 );
or \U$1710 ( \1963 , \1952 , \1960 );
nand \U$1711 ( \1964 , \1962 , \1963 );
not \U$1712 ( \1965 , \1964 );
and \U$1713 ( \1966 , \325 , RIbe281b0_15);
and \U$1714 ( \1967 , \329 , RIbe280c0_13);
nor \U$1715 ( \1968 , \1966 , \1967 );
and \U$1716 ( \1969 , \1968 , \338 );
not \U$1717 ( \1970 , \1968 );
and \U$1718 ( \1971 , \1970 , \1374 );
nor \U$1719 ( \1972 , \1969 , \1971 );
not \U$1720 ( \1973 , \1972 );
and \U$1721 ( \1974 , \1965 , \1973 );
and \U$1722 ( \1975 , \1964 , \1972 );
nor \U$1723 ( \1976 , \1974 , \1975 );
xor \U$1724 ( \1977 , \1945 , \1976 );
not \U$1725 ( \1978 , \1977 );
not \U$1726 ( \1979 , \1827 );
not \U$1727 ( \1980 , \1850 );
or \U$1728 ( \1981 , \1979 , \1980 );
nand \U$1729 ( \1982 , \1981 , \1838 );
not \U$1730 ( \1983 , \1850 );
nand \U$1731 ( \1984 , \1983 , \1826 );
nand \U$1732 ( \1985 , \1982 , \1984 );
nand \U$1733 ( \1986 , \1796 , \1817 );
nand \U$1734 ( \1987 , \1986 , \1803 );
or \U$1735 ( \1988 , \1796 , \1817 );
nand \U$1736 ( \1989 , \1987 , \1988 );
xor \U$1737 ( \1990 , \1985 , \1989 );
not \U$1738 ( \1991 , \1753 );
not \U$1739 ( \1992 , \1766 );
nand \U$1740 ( \1993 , \1992 , \1782 );
nand \U$1741 ( \1994 , \1991 , \1993 );
not \U$1742 ( \1995 , \1782 );
nand \U$1743 ( \1996 , \1995 , \1766 );
nand \U$1744 ( \1997 , \1994 , \1996 );
xor \U$1745 ( \1998 , \1990 , \1997 );
and \U$1746 ( \1999 , \1161 , RIbe28e58_42);
not \U$1747 ( \2000 , \1164 );
and \U$1748 ( \2001 , \2000 , RIbe28de0_41);
nor \U$1749 ( \2002 , \1999 , \2001 );
and \U$1750 ( \2003 , \2002 , \752 );
not \U$1751 ( \2004 , \2002 );
and \U$1752 ( \2005 , \2004 , \1011 );
nor \U$1753 ( \2006 , \2003 , \2005 );
xor \U$1754 ( \2007 , \1458 , \2006 );
not \U$1755 ( \2008 , \1794 );
and \U$1756 ( \2009 , \1143 , RIbe29920_65);
and \U$1757 ( \2010 , \1147 , RIbe27b98_2);
nor \U$1758 ( \2011 , \2009 , \2010 );
not \U$1759 ( \2012 , \2011 );
or \U$1760 ( \2013 , \2008 , \2012 );
or \U$1761 ( \2014 , \2011 , \1469 );
nand \U$1762 ( \2015 , \2013 , \2014 );
xor \U$1763 ( \2016 , \2007 , \2015 );
xor \U$1764 ( \2017 , \1998 , \2016 );
not \U$1765 ( \2018 , \2017 );
or \U$1766 ( \2019 , \1978 , \2018 );
or \U$1767 ( \2020 , \2017 , \1977 );
nand \U$1768 ( \2021 , \2019 , \2020 );
xor \U$1769 ( \2022 , \1908 , \2021 );
xor \U$1770 ( \2023 , \1899 , \2022 );
nand \U$1771 ( \2024 , \1883 , \2023 );
xor \U$1772 ( \2025 , \1887 , \1898 );
and \U$1773 ( \2026 , \2025 , \2022 );
and \U$1774 ( \2027 , \1887 , \1898 );
or \U$1775 ( \2028 , \2026 , \2027 );
not \U$1776 ( \2029 , \2028 );
nand \U$1777 ( \2030 , RIbe29380_53, RIbe281b0_15);
not \U$1778 ( \2031 , \2030 );
and \U$1779 ( \2032 , \1357 , RIbe296c8_60);
and \U$1780 ( \2033 , \264 , RIbe29650_59);
nor \U$1781 ( \2034 , \2032 , \2033 );
and \U$1782 ( \2035 , \2034 , \1363 );
not \U$1783 ( \2036 , \2034 );
and \U$1784 ( \2037 , \2036 , \270 );
nor \U$1785 ( \2038 , \2035 , \2037 );
and \U$1786 ( \2039 , \326 , RIbe280c0_13);
and \U$1787 ( \2040 , \1371 , RIbe29830_63);
nor \U$1788 ( \2041 , \2039 , \2040 );
and \U$1789 ( \2042 , \2041 , \1378 );
not \U$1790 ( \2043 , \2041 );
and \U$1791 ( \2044 , \2043 , \1374 );
nor \U$1792 ( \2045 , \2042 , \2044 );
xor \U$1793 ( \2046 , \2038 , \2045 );
not \U$1794 ( \2047 , \2046 );
or \U$1795 ( \2048 , \2031 , \2047 );
or \U$1796 ( \2049 , \2046 , \2030 );
nand \U$1797 ( \2050 , \2048 , \2049 );
not \U$1798 ( \2051 , RIbe290b0_47);
not \U$1799 ( \2052 , \1223 );
or \U$1800 ( \2053 , \2051 , \2052 );
nand \U$1801 ( \2054 , \429 , RIbe29a88_68);
nand \U$1802 ( \2055 , \2053 , \2054 );
and \U$1803 ( \2056 , \2055 , \306 );
not \U$1804 ( \2057 , \2055 );
and \U$1805 ( \2058 , \2057 , \1547 );
nor \U$1806 ( \2059 , \2056 , \2058 );
and \U$1807 ( \2060 , \1237 , RIbe27d78_6);
and \U$1808 ( \2061 , \554 , RIbe27d00_5);
nor \U$1809 ( \2062 , \2060 , \2061 );
and \U$1810 ( \2063 , \2062 , \1246 );
not \U$1811 ( \2064 , \2062 );
and \U$1812 ( \2065 , \2064 , \1330 );
nor \U$1813 ( \2066 , \2063 , \2065 );
xor \U$1814 ( \2067 , \2059 , \2066 );
and \U$1815 ( \2068 , \283 , RIbe29038_46);
and \U$1816 ( \2069 , \287 , RIbe28fc0_45);
nor \U$1817 ( \2070 , \2068 , \2069 );
and \U$1818 ( \2071 , \2070 , \300 );
not \U$1819 ( \2072 , \2070 );
and \U$1820 ( \2073 , \2072 , \293 );
nor \U$1821 ( \2074 , \2071 , \2073 );
xor \U$1822 ( \2075 , \2067 , \2074 );
and \U$1823 ( \2076 , \2050 , \2075 );
nor \U$1824 ( \2077 , \2050 , \2075 );
nor \U$1825 ( \2078 , \2076 , \2077 );
or \U$1826 ( \2079 , \1893 , \1857 );
and \U$1827 ( \2080 , \2079 , \1891 );
and \U$1828 ( \2081 , \1893 , \1857 );
nor \U$1829 ( \2082 , \2080 , \2081 );
xor \U$1830 ( \2083 , \2078 , \2082 );
and \U$1831 ( \2084 , \1998 , \2016 );
not \U$1832 ( \2085 , \1998 );
not \U$1833 ( \2086 , \2016 );
and \U$1834 ( \2087 , \2085 , \2086 );
nor \U$1835 ( \2088 , \2087 , \1977 );
nor \U$1836 ( \2089 , \2084 , \2088 );
xor \U$1837 ( \2090 , \2083 , \2089 );
xor \U$1838 ( \2091 , \1943 , \1944 );
and \U$1839 ( \2092 , \2091 , \1976 );
and \U$1840 ( \2093 , \1943 , \1944 );
or \U$1841 ( \2094 , \2092 , \2093 );
not \U$1842 ( \2095 , \2094 );
xor \U$1843 ( \2096 , \1985 , \1989 );
and \U$1844 ( \2097 , \2096 , \1997 );
and \U$1845 ( \2098 , \1985 , \1989 );
or \U$1846 ( \2099 , \2097 , \2098 );
and \U$1847 ( \2100 , \1005 , RIbe28de0_41);
and \U$1848 ( \2101 , \1203 , RIbe29920_65);
nor \U$1849 ( \2102 , \2100 , \2101 );
and \U$1850 ( \2103 , \2102 , \752 );
not \U$1851 ( \2104 , \2102 );
and \U$1852 ( \2105 , \2104 , \1011 );
nor \U$1853 ( \2106 , \2103 , \2105 );
and \U$1854 ( \2107 , \666 , RIbe27c10_3);
and \U$1855 ( \2108 , \740 , RIbe28e58_42);
nor \U$1856 ( \2109 , \2107 , \2108 );
and \U$1857 ( \2110 , \2109 , \564 );
not \U$1858 ( \2111 , \2109 );
and \U$1859 ( \2112 , \2111 , \672 );
nor \U$1860 ( \2113 , \2110 , \2112 );
xor \U$1861 ( \2114 , \2106 , \2113 );
nand \U$1862 ( \2115 , \1143 , RIbe27b98_2);
and \U$1863 ( \2116 , \2115 , \1152 );
not \U$1864 ( \2117 , \2115 );
and \U$1865 ( \2118 , \2117 , \1652 );
nor \U$1866 ( \2119 , \2116 , \2118 );
xor \U$1867 ( \2120 , \2114 , \2119 );
xor \U$1868 ( \2121 , \2099 , \2120 );
not \U$1869 ( \2122 , \2121 );
or \U$1870 ( \2123 , \2095 , \2122 );
or \U$1871 ( \2124 , \2121 , \2094 );
nand \U$1872 ( \2125 , \2123 , \2124 );
not \U$1873 ( \2126 , \2125 );
not \U$1874 ( \2127 , \1917 );
nand \U$1875 ( \2128 , \2127 , \1939 );
nand \U$1876 ( \2129 , \2128 , \1927 );
not \U$1877 ( \2130 , \1939 );
nand \U$1878 ( \2131 , \2130 , \1917 );
nand \U$1879 ( \2132 , \2129 , \2131 );
xor \U$1880 ( \2133 , \1458 , \2006 );
and \U$1881 ( \2134 , \2133 , \2015 );
and \U$1882 ( \2135 , \1458 , \2006 );
or \U$1883 ( \2136 , \2134 , \2135 );
xnor \U$1884 ( \2137 , \2132 , \2136 );
not \U$1885 ( \2138 , \2137 );
or \U$1886 ( \2139 , \1972 , \1952 );
not \U$1887 ( \2140 , \1952 );
not \U$1888 ( \2141 , \1972 );
or \U$1889 ( \2142 , \2140 , \2141 );
nand \U$1890 ( \2143 , \2142 , \1960 );
nand \U$1891 ( \2144 , \2139 , \2143 );
not \U$1892 ( \2145 , \2144 );
and \U$1893 ( \2146 , \2138 , \2145 );
and \U$1894 ( \2147 , \2137 , \2144 );
nor \U$1895 ( \2148 , \2146 , \2147 );
not \U$1896 ( \2149 , \2148 );
and \U$1897 ( \2150 , \2126 , \2149 );
and \U$1898 ( \2151 , \2125 , \2148 );
nor \U$1899 ( \2152 , \2150 , \2151 );
xnor \U$1900 ( \2153 , \2090 , \2152 );
not \U$1901 ( \2154 , \2153 );
xor \U$1902 ( \2155 , \1903 , \1907 );
and \U$1903 ( \2156 , \2155 , \2021 );
and \U$1904 ( \2157 , \1903 , \1907 );
or \U$1905 ( \2158 , \2156 , \2157 );
not \U$1906 ( \2159 , \2158 );
and \U$1907 ( \2160 , \2154 , \2159 );
and \U$1908 ( \2161 , \2153 , \2158 );
nor \U$1909 ( \2162 , \2160 , \2161 );
not \U$1910 ( \2163 , \2162 );
or \U$1911 ( \2164 , \2029 , \2163 );
or \U$1912 ( \2165 , \2028 , \2162 );
nand \U$1913 ( \2166 , \2164 , \2165 );
xor \U$1914 ( \2167 , \2024 , \2166 );
and \U$1915 ( \2168 , \2099 , \2120 );
not \U$1916 ( \2169 , \2099 );
not \U$1917 ( \2170 , \2120 );
and \U$1918 ( \2171 , \2169 , \2170 );
nor \U$1919 ( \2172 , \2171 , \2094 );
nor \U$1920 ( \2173 , \2168 , \2172 );
xor \U$1921 ( \2174 , \2059 , \2066 );
and \U$1922 ( \2175 , \2174 , \2074 );
and \U$1923 ( \2176 , \2059 , \2066 );
nor \U$1924 ( \2177 , \2175 , \2176 );
not \U$1925 ( \2178 , \2038 );
not \U$1926 ( \2179 , \2030 );
and \U$1927 ( \2180 , \2178 , \2179 );
and \U$1928 ( \2181 , \2038 , \2030 );
nor \U$1929 ( \2182 , \2181 , \2045 );
nor \U$1930 ( \2183 , \2180 , \2182 );
xor \U$1931 ( \2184 , \2177 , \2183 );
xor \U$1932 ( \2185 , \2106 , \2113 );
and \U$1933 ( \2186 , \2185 , \2119 );
and \U$1934 ( \2187 , \2106 , \2113 );
nor \U$1935 ( \2188 , \2186 , \2187 );
xor \U$1936 ( \2189 , \2184 , \2188 );
xor \U$1937 ( \2190 , \2173 , \2189 );
and \U$1938 ( \2191 , \326 , RIbe29830_63);
and \U$1939 ( \2192 , \1371 , RIbe296c8_60);
nor \U$1940 ( \2193 , \2191 , \2192 );
and \U$1941 ( \2194 , \2193 , \1374 );
not \U$1942 ( \2195 , \2193 );
and \U$1943 ( \2196 , \2195 , \1378 );
or \U$1944 ( \2197 , \2194 , \2196 );
not \U$1945 ( \2198 , \2197 );
and \U$1946 ( \2199 , \1516 , RIbe29650_59);
and \U$1947 ( \2200 , \1831 , RIbe29038_46);
nor \U$1948 ( \2201 , \2199 , \2200 );
and \U$1949 ( \2202 , \2201 , \1362 );
not \U$1950 ( \2203 , \2201 );
and \U$1951 ( \2204 , \2203 , \1663 );
nor \U$1952 ( \2205 , \2202 , \2204 );
not \U$1953 ( \2206 , \2205 );
or \U$1954 ( \2207 , \2198 , \2206 );
or \U$1955 ( \2208 , \2197 , \2205 );
nand \U$1956 ( \2209 , \2207 , \2208 );
not \U$1957 ( \2210 , \2209 );
nand \U$1958 ( \2211 , RIbe29380_53, RIbe280c0_13);
not \U$1959 ( \2212 , \2211 );
and \U$1960 ( \2213 , \2210 , \2212 );
and \U$1961 ( \2214 , \2209 , \2211 );
nor \U$1962 ( \2215 , \2213 , \2214 );
and \U$1963 ( \2216 , \666 , RIbe28e58_42);
and \U$1964 ( \2217 , \1180 , RIbe28de0_41);
nor \U$1965 ( \2218 , \2216 , \2217 );
and \U$1966 ( \2219 , \2218 , \672 );
not \U$1967 ( \2220 , \2218 );
and \U$1968 ( \2221 , \2220 , \564 );
nor \U$1969 ( \2222 , \2219 , \2221 );
xor \U$1970 ( \2223 , \2222 , \1794 );
and \U$1971 ( \2224 , \1005 , RIbe29920_65);
and \U$1972 ( \2225 , \1203 , RIbe27b98_2);
nor \U$1973 ( \2226 , \2224 , \2225 );
and \U$1974 ( \2227 , \2226 , \1011 );
not \U$1975 ( \2228 , \2226 );
and \U$1976 ( \2229 , \2228 , \752 );
nor \U$1977 ( \2230 , \2227 , \2229 );
xor \U$1978 ( \2231 , \2223 , \2230 );
xor \U$1979 ( \2232 , \2215 , \2231 );
and \U$1980 ( \2233 , \283 , RIbe28fc0_45);
and \U$1981 ( \2234 , \287 , RIbe290b0_47);
nor \U$1982 ( \2235 , \2233 , \2234 );
and \U$1983 ( \2236 , \2235 , \293 );
not \U$1984 ( \2237 , \2235 );
and \U$1985 ( \2238 , \2237 , \300 );
nor \U$1986 ( \2239 , \2236 , \2238 );
and \U$1987 ( \2240 , \549 , RIbe27d00_5);
and \U$1988 ( \2241 , \554 , RIbe27c10_3);
nor \U$1989 ( \2242 , \2240 , \2241 );
and \U$1990 ( \2243 , \2242 , \425 );
not \U$1991 ( \2244 , \2242 );
and \U$1992 ( \2245 , \2244 , \424 );
nor \U$1993 ( \2246 , \2243 , \2245 );
xor \U$1994 ( \2247 , \2239 , \2246 );
and \U$1995 ( \2248 , \383 , RIbe29a88_68);
and \U$1996 ( \2249 , \429 , RIbe27d78_6);
nor \U$1997 ( \2250 , \2248 , \2249 );
and \U$1998 ( \2251 , \2250 , \306 );
not \U$1999 ( \2252 , \2250 );
and \U$2000 ( \2253 , \2252 , \313 );
nor \U$2001 ( \2254 , \2251 , \2253 );
xor \U$2002 ( \2255 , \2247 , \2254 );
xor \U$2003 ( \2256 , \2232 , \2255 );
not \U$2004 ( \2257 , \2256 );
not \U$2005 ( \2258 , \2136 );
not \U$2006 ( \2259 , \2144 );
or \U$2007 ( \2260 , \2258 , \2259 );
or \U$2008 ( \2261 , \2144 , \2136 );
nand \U$2009 ( \2262 , \2261 , \2132 );
nand \U$2010 ( \2263 , \2260 , \2262 );
not \U$2011 ( \2264 , \2263 );
not \U$2012 ( \2265 , \2077 );
or \U$2013 ( \2266 , \2264 , \2265 );
or \U$2014 ( \2267 , \2077 , \2263 );
nand \U$2015 ( \2268 , \2266 , \2267 );
not \U$2016 ( \2269 , \2268 );
and \U$2017 ( \2270 , \2257 , \2269 );
and \U$2018 ( \2271 , \2256 , \2268 );
nor \U$2019 ( \2272 , \2270 , \2271 );
xor \U$2020 ( \2273 , \2190 , \2272 );
not \U$2021 ( \2274 , \2148 );
nand \U$2022 ( \2275 , \2274 , \2125 );
xor \U$2023 ( \2276 , \2273 , \2275 );
xor \U$2024 ( \2277 , \2078 , \2082 );
and \U$2025 ( \2278 , \2277 , \2089 );
and \U$2026 ( \2279 , \2078 , \2082 );
nor \U$2027 ( \2280 , \2278 , \2279 );
not \U$2028 ( \2281 , \2280 );
xor \U$2029 ( \2282 , \2276 , \2281 );
not \U$2030 ( \2283 , \2282 );
or \U$2031 ( \2284 , \2152 , \2090 );
not \U$2032 ( \2285 , \2152 );
not \U$2033 ( \2286 , \2090 );
or \U$2034 ( \2287 , \2285 , \2286 );
nand \U$2035 ( \2288 , \2287 , \2158 );
nand \U$2036 ( \2289 , \2284 , \2288 );
not \U$2037 ( \2290 , \2289 );
and \U$2038 ( \2291 , \2283 , \2290 );
and \U$2039 ( \2292 , \2282 , \2289 );
nor \U$2040 ( \2293 , \2291 , \2292 );
not \U$2041 ( \2294 , \2162 );
nand \U$2042 ( \2295 , \2294 , \2028 );
xnor \U$2043 ( \2296 , \2293 , \2295 );
nor \U$2044 ( \2297 , \2167 , \2296 );
not \U$2045 ( \2298 , \1882 );
not \U$2046 ( \2299 , \2023 );
or \U$2047 ( \2300 , \2298 , \2299 );
or \U$2048 ( \2301 , \2023 , \1882 );
nand \U$2049 ( \2302 , \2300 , \2301 );
xnor \U$2050 ( \2303 , \1560 , \1417 );
not \U$2051 ( \2304 , \2303 );
not \U$2052 ( \2305 , \1696 );
and \U$2053 ( \2306 , \2304 , \2305 );
and \U$2054 ( \2307 , \2303 , \1696 );
nor \U$2055 ( \2308 , \2306 , \2307 );
not \U$2056 ( \2309 , \2308 );
xnor \U$2057 ( \2310 , \1728 , \1730 );
not \U$2058 ( \2311 , \2310 );
not \U$2059 ( \2312 , \1738 );
and \U$2060 ( \2313 , \2311 , \2312 );
and \U$2061 ( \2314 , \2310 , \1738 );
nor \U$2062 ( \2315 , \2313 , \2314 );
not \U$2063 ( \2316 , \2315 );
and \U$2064 ( \2317 , \2309 , \2316 );
and \U$2065 ( \2318 , \2308 , \2315 );
xor \U$2066 ( \2319 , \1221 , \1264 );
not \U$2067 ( \2320 , \1315 );
xor \U$2068 ( \2321 , \2319 , \2320 );
not \U$2069 ( \2322 , \1135 );
not \U$2070 ( \2323 , \1187 );
and \U$2071 ( \2324 , \2322 , \2323 );
and \U$2072 ( \2325 , \1187 , \1135 );
nor \U$2073 ( \2326 , \2324 , \2325 );
xor \U$2074 ( \2327 , \2321 , \2326 );
xor \U$2075 ( \2328 , \1354 , \1384 );
xor \U$2076 ( \2329 , \2328 , \1411 );
and \U$2077 ( \2330 , \2327 , \2329 );
and \U$2078 ( \2331 , \2321 , \2326 );
or \U$2079 ( \2332 , \2330 , \2331 );
not \U$2080 ( \2333 , RIbe281b0_15);
not \U$2081 ( \2334 , \1223 );
or \U$2082 ( \2335 , \2333 , \2334 );
nand \U$2083 ( \2336 , \429 , RIbe280c0_13);
nand \U$2084 ( \2337 , \2335 , \2336 );
and \U$2085 ( \2338 , \2337 , \1547 );
not \U$2086 ( \2339 , \2337 );
and \U$2087 ( \2340 , \2339 , \306 );
nor \U$2088 ( \2341 , \2338 , \2340 );
not \U$2089 ( \2342 , RIbe29830_63);
not \U$2090 ( \2343 , \1756 );
or \U$2091 ( \2344 , \2342 , \2343 );
nand \U$2092 ( \2345 , \553 , RIbe296c8_60);
nand \U$2093 ( \2346 , \2344 , \2345 );
and \U$2094 ( \2347 , \2346 , \1330 );
not \U$2095 ( \2348 , \2346 );
and \U$2096 ( \2349 , \2348 , \424 );
nor \U$2097 ( \2350 , \2347 , \2349 );
not \U$2098 ( \2351 , \2350 );
nand \U$2099 ( \2352 , \2341 , \2351 );
not \U$2100 ( \2353 , \2352 );
not \U$2101 ( \2354 , \1611 );
not \U$2102 ( \2355 , RIbe29038_46);
not \U$2103 ( \2356 , \2355 );
and \U$2104 ( \2357 , \2354 , \2356 );
and \U$2105 ( \2358 , \664 , RIbe29650_59);
nor \U$2106 ( \2359 , \2357 , \2358 );
and \U$2107 ( \2360 , \2359 , \1621 );
not \U$2108 ( \2361 , \2359 );
and \U$2109 ( \2362 , \2361 , \564 );
nor \U$2110 ( \2363 , \2360 , \2362 );
not \U$2111 ( \2364 , \2363 );
not \U$2112 ( \2365 , \2364 );
or \U$2113 ( \2366 , \2353 , \2365 );
or \U$2114 ( \2367 , \2351 , \2341 );
nand \U$2115 ( \2368 , \2366 , \2367 );
and \U$2116 ( \2369 , \1113 , RIbe28e58_42);
and \U$2117 ( \2370 , \1117 , RIbe28de0_41);
nor \U$2118 ( \2371 , \2369 , \2370 );
and \U$2119 ( \2372 , \2371 , \1125 );
not \U$2120 ( \2373 , \2371 );
and \U$2121 ( \2374 , \2373 , \1132 );
nor \U$2122 ( \2375 , \2372 , \2374 );
not \U$2123 ( \2376 , \2375 );
nand \U$2124 ( \2377 , RIbe29b00_69, RIbe29128_48);
nand \U$2125 ( \2378 , \2377 , RIbe291a0_49);
buf \U$2126 ( \2379 , \2378 );
not \U$2127 ( \2380 , \2379 );
or \U$2128 ( \2381 , \2376 , \2380 );
or \U$2129 ( \2382 , \2375 , \2379 );
xor \U$2130 ( \2383 , RIbe295d8_58, RIbe291a0_49);
buf \U$2131 ( \2384 , \2383 );
not \U$2132 ( \2385 , \2384 );
not \U$2133 ( \2386 , \2385 );
not \U$2134 ( \2387 , \1640 );
and \U$2135 ( \2388 , \2386 , \2387 );
not \U$2136 ( \2389 , \1270 );
not \U$2137 ( \2390 , \2389 );
buf \U$2138 ( \2391 , \2390 );
and \U$2139 ( \2392 , \2391 , RIbe29920_65);
nor \U$2140 ( \2393 , \2388 , \2392 );
and \U$2141 ( \2394 , \2393 , \1076 );
not \U$2142 ( \2395 , \2393 );
and \U$2143 ( \2396 , \2395 , \1277 );
nor \U$2144 ( \2397 , \2394 , \2396 );
nand \U$2145 ( \2398 , \2382 , \2397 );
nand \U$2146 ( \2399 , \2381 , \2398 );
xor \U$2147 ( \2400 , \2368 , \2399 );
not \U$2148 ( \2401 , RIbe29a88_68);
not \U$2149 ( \2402 , \1143 );
or \U$2150 ( \2403 , \2401 , \2402 );
nand \U$2151 ( \2404 , \1147 , RIbe27d78_6);
nand \U$2152 ( \2405 , \2403 , \2404 );
and \U$2153 ( \2406 , \2405 , \1154 );
not \U$2154 ( \2407 , \2405 );
and \U$2155 ( \2408 , \2407 , \1152 );
nor \U$2156 ( \2409 , \2406 , \2408 );
not \U$2157 ( \2410 , \2409 );
not \U$2158 ( \2411 , RIbe27d00_5);
not \U$2159 ( \2412 , \1094 );
or \U$2160 ( \2413 , \2411 , \2412 );
nand \U$2161 ( \2414 , \1099 , RIbe27c10_3);
nand \U$2162 ( \2415 , \2413 , \2414 );
and \U$2163 ( \2416 , \2415 , \1309 );
not \U$2164 ( \2417 , \2415 );
not \U$2165 ( \2418 , \1081 );
and \U$2166 ( \2419 , \2417 , \2418 );
nor \U$2167 ( \2420 , \2416 , \2419 );
not \U$2168 ( \2421 , \2420 );
or \U$2169 ( \2422 , \2410 , \2421 );
or \U$2170 ( \2423 , \2409 , \2420 );
not \U$2171 ( \2424 , \1001 );
buf \U$2172 ( \2425 , \2424 );
and \U$2173 ( \2426 , \2425 , RIbe28fc0_45);
and \U$2174 ( \2427 , \1203 , RIbe290b0_47);
nor \U$2175 ( \2428 , \2426 , \2427 );
and \U$2176 ( \2429 , \2428 , \1011 );
not \U$2177 ( \2430 , \2428 );
and \U$2178 ( \2431 , \2430 , \752 );
nor \U$2179 ( \2432 , \2429 , \2431 );
not \U$2180 ( \2433 , \2432 );
nand \U$2181 ( \2434 , \2423 , \2433 );
nand \U$2182 ( \2435 , \2422 , \2434 );
and \U$2183 ( \2436 , \2400 , \2435 );
and \U$2184 ( \2437 , \2368 , \2399 );
or \U$2185 ( \2438 , \2436 , \2437 );
xor \U$2186 ( \2439 , \1355 , \1367 );
xor \U$2187 ( \2440 , \2439 , \1381 );
and \U$2188 ( \2441 , \1357 , RIbe289a8_32);
and \U$2189 ( \2442 , \264 , RIbe28930_31);
nor \U$2190 ( \2443 , \2441 , \2442 );
and \U$2191 ( \2444 , \2443 , \1663 );
not \U$2192 ( \2445 , \2443 );
and \U$2193 ( \2446 , \2445 , \1362 );
nor \U$2194 ( \2447 , \2444 , \2446 );
and \U$2195 ( \2448 , \283 , RIbe29560_57);
and \U$2196 ( \2449 , \1682 , RIbe28228_16);
nor \U$2197 ( \2450 , \2448 , \2449 );
and \U$2198 ( \2451 , \2450 , \293 );
not \U$2199 ( \2452 , \2450 );
and \U$2200 ( \2453 , \2452 , \300 );
nor \U$2201 ( \2454 , \2451 , \2453 );
xor \U$2202 ( \2455 , \2447 , \2454 );
and \U$2203 ( \2456 , \326 , RIbe29290_51);
and \U$2204 ( \2457 , \330 , RIbe28a20_33);
nor \U$2205 ( \2458 , \2456 , \2457 );
and \U$2206 ( \2459 , \2458 , \1378 );
not \U$2207 ( \2460 , \2458 );
and \U$2208 ( \2461 , \2460 , \339 );
nor \U$2209 ( \2462 , \2459 , \2461 );
and \U$2210 ( \2463 , \2455 , \2462 );
and \U$2211 ( \2464 , \2447 , \2454 );
or \U$2212 ( \2465 , \2463 , \2464 );
nand \U$2213 ( \2466 , \2440 , \2465 );
xor \U$2214 ( \2467 , \2438 , \2466 );
not \U$2215 ( \2468 , \1311 );
and \U$2216 ( \2469 , \1294 , \1282 );
not \U$2217 ( \2470 , \1294 );
and \U$2218 ( \2471 , \2470 , \1281 );
nor \U$2219 ( \2472 , \2469 , \2471 );
not \U$2220 ( \2473 , \2472 );
or \U$2221 ( \2474 , \2468 , \2473 );
or \U$2222 ( \2475 , \2472 , \1311 );
nand \U$2223 ( \2476 , \2474 , \2475 );
not \U$2224 ( \2477 , \1262 );
xor \U$2225 ( \2478 , \1234 , \1248 );
not \U$2226 ( \2479 , \2478 );
or \U$2227 ( \2480 , \2477 , \2479 );
or \U$2228 ( \2481 , \2478 , \1262 );
nand \U$2229 ( \2482 , \2480 , \2481 );
xor \U$2230 ( \2483 , \2476 , \2482 );
not \U$2231 ( \2484 , \1219 );
xor \U$2232 ( \2485 , \1199 , \1209 );
not \U$2233 ( \2486 , \2485 );
or \U$2234 ( \2487 , \2484 , \2486 );
or \U$2235 ( \2488 , \2485 , \1219 );
nand \U$2236 ( \2489 , \2487 , \2488 );
and \U$2237 ( \2490 , \2483 , \2489 );
and \U$2238 ( \2491 , \2476 , \2482 );
or \U$2239 ( \2492 , \2490 , \2491 );
and \U$2240 ( \2493 , \2467 , \2492 );
and \U$2241 ( \2494 , \2438 , \2466 );
nor \U$2242 ( \2495 , \2493 , \2494 );
xor \U$2243 ( \2496 , \2332 , \2495 );
xnor \U$2244 ( \2497 , \1493 , \1476 );
not \U$2245 ( \2498 , \2497 );
not \U$2246 ( \2499 , \1558 );
and \U$2247 ( \2500 , \2498 , \2499 );
and \U$2248 ( \2501 , \2497 , \1558 );
nor \U$2249 ( \2502 , \2500 , \2501 );
and \U$2250 ( \2503 , \2496 , \2502 );
and \U$2251 ( \2504 , \2332 , \2495 );
or \U$2252 ( \2505 , \2503 , \2504 );
nor \U$2253 ( \2506 , \2318 , \2505 );
nor \U$2254 ( \2507 , \2317 , \2506 );
not \U$2255 ( \2508 , \2507 );
not \U$2256 ( \2509 , \1880 );
xnor \U$2257 ( \2510 , \1698 , \1712 );
not \U$2258 ( \2511 , \2510 );
or \U$2259 ( \2512 , \2509 , \2511 );
or \U$2260 ( \2513 , \2510 , \1880 );
nand \U$2261 ( \2514 , \2512 , \2513 );
nand \U$2262 ( \2515 , \2508 , \2514 );
xor \U$2263 ( \2516 , \2302 , \2515 );
not \U$2264 ( \2517 , \2516 );
xor \U$2265 ( \2518 , \2321 , \2326 );
xor \U$2266 ( \2519 , \2518 , \2329 );
not \U$2267 ( \2520 , RIbe280c0_13);
not \U$2268 ( \2521 , \549 );
or \U$2269 ( \2522 , \2520 , \2521 );
nand \U$2270 ( \2523 , \554 , RIbe29830_63);
nand \U$2271 ( \2524 , \2522 , \2523 );
not \U$2272 ( \2525 , \2524 );
not \U$2273 ( \2526 , \424 );
and \U$2274 ( \2527 , \2525 , \2526 );
and \U$2275 ( \2528 , \2524 , \1333 );
nor \U$2276 ( \2529 , \2527 , \2528 );
not \U$2277 ( \2530 , RIbe296c8_60);
not \U$2278 ( \2531 , \1743 );
not \U$2279 ( \2532 , \2531 );
or \U$2280 ( \2533 , \2530 , \2532 );
nand \U$2281 ( \2534 , \1180 , RIbe29650_59);
nand \U$2282 ( \2535 , \2533 , \2534 );
not \U$2283 ( \2536 , \2535 );
not \U$2284 ( \2537 , \1618 );
and \U$2285 ( \2538 , \2536 , \2537 );
and \U$2286 ( \2539 , \2535 , \1618 );
nor \U$2287 ( \2540 , \2538 , \2539 );
xor \U$2288 ( \2541 , \2529 , \2540 );
not \U$2289 ( \2542 , RIbe28228_16);
not \U$2290 ( \2543 , \1774 );
or \U$2291 ( \2544 , \2542 , \2543 );
nand \U$2292 ( \2545 , \429 , RIbe281b0_15);
nand \U$2293 ( \2546 , \2544 , \2545 );
and \U$2294 ( \2547 , \2546 , \313 );
not \U$2295 ( \2548 , \2546 );
and \U$2296 ( \2549 , \2548 , \306 );
nor \U$2297 ( \2550 , \2547 , \2549 );
and \U$2298 ( \2551 , \2541 , \2550 );
and \U$2299 ( \2552 , \2529 , \2540 );
or \U$2300 ( \2553 , \2551 , \2552 );
not \U$2301 ( \2554 , \1284 );
buf \U$2302 ( \2555 , \2554 );
not \U$2303 ( \2556 , \2555 );
not \U$2304 ( \2557 , \2556 );
and \U$2305 ( \2558 , \2557 , RIbe27c10_3);
and \U$2306 ( \2559 , \1117 , RIbe28e58_42);
nor \U$2307 ( \2560 , \2558 , \2559 );
and \U$2308 ( \2561 , \2560 , \1132 );
not \U$2309 ( \2562 , \2560 );
not \U$2310 ( \2563 , \1124 );
and \U$2311 ( \2564 , \2562 , \2563 );
nor \U$2312 ( \2565 , \2561 , \2564 );
xor \U$2313 ( \2566 , RIbe29128_48, RIbe29b00_69);
not \U$2314 ( \2567 , \2566 );
xor \U$2315 ( \2568 , RIbe29128_48, RIbe291a0_49);
nand \U$2316 ( \2569 , \2567 , \2568 );
buf \U$2317 ( \2570 , \2569 );
not \U$2318 ( \2571 , \2570 );
nand \U$2319 ( \2572 , \2571 , RIbe27b98_2);
not \U$2320 ( \2573 , \2379 );
and \U$2321 ( \2574 , \2572 , \2573 );
not \U$2322 ( \2575 , \2572 );
buf \U$2323 ( \2576 , \2379 );
and \U$2324 ( \2577 , \2575 , \2576 );
nor \U$2325 ( \2578 , \2574 , \2577 );
and \U$2326 ( \2579 , \2565 , \2578 );
not \U$2327 ( \2580 , \2385 );
not \U$2328 ( \2581 , \1636 );
and \U$2329 ( \2582 , \2580 , \2581 );
buf \U$2330 ( \2583 , \1270 );
and \U$2331 ( \2584 , \2583 , RIbe28de0_41);
nor \U$2332 ( \2585 , \2582 , \2584 );
and \U$2333 ( \2586 , \2585 , \1076 );
not \U$2334 ( \2587 , \2585 );
and \U$2335 ( \2588 , \2587 , \1277 );
nor \U$2336 ( \2589 , \2586 , \2588 );
not \U$2337 ( \2590 , \2589 );
nor \U$2338 ( \2591 , \2579 , \2590 );
nor \U$2339 ( \2592 , \2565 , \2578 );
nor \U$2340 ( \2593 , \2591 , \2592 );
xor \U$2341 ( \2594 , \2553 , \2593 );
not \U$2342 ( \2595 , RIbe290b0_47);
buf \U$2343 ( \2596 , \1141 );
not \U$2344 ( \2597 , \2596 );
not \U$2345 ( \2598 , \2597 );
or \U$2346 ( \2599 , \2595 , \2598 );
nand \U$2347 ( \2600 , \1147 , RIbe29a88_68);
nand \U$2348 ( \2601 , \2599 , \2600 );
and \U$2349 ( \2602 , \2601 , \1152 );
not \U$2350 ( \2603 , \2601 );
and \U$2351 ( \2604 , \2603 , \1794 );
nor \U$2352 ( \2605 , \2602 , \2604 );
and \U$2353 ( \2606 , \2425 , RIbe29038_46);
and \U$2354 ( \2607 , \1203 , RIbe28fc0_45);
nor \U$2355 ( \2608 , \2606 , \2607 );
and \U$2356 ( \2609 , \2608 , \1011 );
not \U$2357 ( \2610 , \2608 );
and \U$2358 ( \2611 , \2610 , \1608 );
nor \U$2359 ( \2612 , \2609 , \2611 );
xor \U$2360 ( \2613 , \2605 , \2612 );
not \U$2361 ( \2614 , RIbe27d78_6);
not \U$2362 ( \2615 , \1298 );
or \U$2363 ( \2616 , \2614 , \2615 );
nand \U$2364 ( \2617 , \1099 , RIbe27d00_5);
nand \U$2365 ( \2618 , \2616 , \2617 );
and \U$2366 ( \2619 , \2618 , \1458 );
not \U$2367 ( \2620 , \2618 );
and \U$2368 ( \2621 , \2620 , \1309 );
nor \U$2369 ( \2622 , \2619 , \2621 );
and \U$2370 ( \2623 , \2613 , \2622 );
and \U$2371 ( \2624 , \2605 , \2612 );
or \U$2372 ( \2625 , \2623 , \2624 );
and \U$2373 ( \2626 , \2594 , \2625 );
and \U$2374 ( \2627 , \2553 , \2593 );
or \U$2375 ( \2628 , \2626 , \2627 );
nand \U$2376 ( \2629 , RIbe29380_53, RIbe28b88_36);
nand \U$2377 ( \2630 , RIbe29380_53, RIbe28b10_35);
xor \U$2378 ( \2631 , \2629 , \2630 );
not \U$2379 ( \2632 , RIbe28b88_36);
not \U$2380 ( \2633 , \326 );
or \U$2381 ( \2634 , \2632 , \2633 );
nand \U$2382 ( \2635 , \330 , RIbe29290_51);
nand \U$2383 ( \2636 , \2634 , \2635 );
not \U$2384 ( \2637 , \2636 );
not \U$2385 ( \2638 , \1379 );
and \U$2386 ( \2639 , \2637 , \2638 );
and \U$2387 ( \2640 , \2636 , \339 );
nor \U$2388 ( \2641 , \2639 , \2640 );
not \U$2389 ( \2642 , \2641 );
and \U$2390 ( \2643 , \1254 , RIbe28930_31);
and \U$2391 ( \2644 , \1256 , RIbe29560_57);
nor \U$2392 ( \2645 , \2643 , \2644 );
and \U$2393 ( \2646 , \2645 , \293 );
not \U$2394 ( \2647 , \2645 );
and \U$2395 ( \2648 , \2647 , \300 );
nor \U$2396 ( \2649 , \2646 , \2648 );
not \U$2397 ( \2650 , \2649 );
and \U$2398 ( \2651 , \2642 , \2650 );
and \U$2399 ( \2652 , \2649 , \2641 );
and \U$2400 ( \2653 , \1516 , RIbe28a20_33);
and \U$2401 ( \2654 , \1831 , RIbe289a8_32);
nor \U$2402 ( \2655 , \2653 , \2654 );
and \U$2403 ( \2656 , \2655 , \1362 );
not \U$2404 ( \2657 , \2655 );
and \U$2405 ( \2658 , \2657 , \269 );
nor \U$2406 ( \2659 , \2656 , \2658 );
not \U$2407 ( \2660 , \2659 );
nor \U$2408 ( \2661 , \2652 , \2660 );
nor \U$2409 ( \2662 , \2651 , \2661 );
and \U$2410 ( \2663 , \2631 , \2662 );
and \U$2411 ( \2664 , \2629 , \2630 );
or \U$2412 ( \2665 , \2663 , \2664 );
xor \U$2413 ( \2666 , \2628 , \2665 );
not \U$2414 ( \2667 , \2351 );
not \U$2415 ( \2668 , \2364 );
or \U$2416 ( \2669 , \2667 , \2668 );
nand \U$2417 ( \2670 , \2350 , \2363 );
nand \U$2418 ( \2671 , \2669 , \2670 );
xor \U$2419 ( \2672 , \2671 , \2341 );
xor \U$2420 ( \2673 , \2409 , \2420 );
xor \U$2421 ( \2674 , \2673 , \2432 );
xor \U$2422 ( \2675 , \2672 , \2674 );
xor \U$2423 ( \2676 , \2447 , \2454 );
xor \U$2424 ( \2677 , \2676 , \2462 );
and \U$2425 ( \2678 , \2675 , \2677 );
and \U$2426 ( \2679 , \2672 , \2674 );
or \U$2427 ( \2680 , \2678 , \2679 );
and \U$2428 ( \2681 , \2666 , \2680 );
and \U$2429 ( \2682 , \2628 , \2665 );
or \U$2430 ( \2683 , \2681 , \2682 );
xor \U$2431 ( \2684 , \2519 , \2683 );
xor \U$2432 ( \2685 , \2368 , \2399 );
xor \U$2433 ( \2686 , \2685 , \2435 );
or \U$2434 ( \2687 , \2440 , \2465 );
nand \U$2435 ( \2688 , \2687 , \2466 );
xor \U$2436 ( \2689 , \2686 , \2688 );
xor \U$2437 ( \2690 , \2476 , \2482 );
xor \U$2438 ( \2691 , \2690 , \2489 );
and \U$2439 ( \2692 , \2689 , \2691 );
and \U$2440 ( \2693 , \2686 , \2688 );
or \U$2441 ( \2694 , \2692 , \2693 );
not \U$2442 ( \2695 , \2694 );
and \U$2443 ( \2696 , \2684 , \2695 );
and \U$2444 ( \2697 , \2519 , \2683 );
or \U$2445 ( \2698 , \2696 , \2697 );
xor \U$2446 ( \2699 , \1320 , \1188 );
not \U$2447 ( \2700 , \2699 );
not \U$2448 ( \2701 , \1414 );
and \U$2449 ( \2702 , \2700 , \2701 );
and \U$2450 ( \2703 , \2699 , \1414 );
nor \U$2451 ( \2704 , \2702 , \2703 );
xor \U$2452 ( \2705 , \2698 , \2704 );
xor \U$2453 ( \2706 , \2332 , \2495 );
xor \U$2454 ( \2707 , \2706 , \2502 );
and \U$2455 ( \2708 , \2705 , \2707 );
and \U$2456 ( \2709 , \2698 , \2704 );
or \U$2457 ( \2710 , \2708 , \2709 );
not \U$2458 ( \2711 , \2710 );
not \U$2459 ( \2712 , \2308 );
xor \U$2460 ( \2713 , \2505 , \2315 );
not \U$2461 ( \2714 , \2713 );
or \U$2462 ( \2715 , \2712 , \2714 );
or \U$2463 ( \2716 , \2713 , \2308 );
nand \U$2464 ( \2717 , \2715 , \2716 );
nand \U$2465 ( \2718 , \2711 , \2717 );
not \U$2466 ( \2719 , \2718 );
not \U$2467 ( \2720 , \2507 );
not \U$2468 ( \2721 , \2514 );
or \U$2469 ( \2722 , \2720 , \2721 );
or \U$2470 ( \2723 , \2507 , \2514 );
nand \U$2471 ( \2724 , \2722 , \2723 );
not \U$2472 ( \2725 , \2724 );
and \U$2473 ( \2726 , \2719 , \2725 );
and \U$2474 ( \2727 , \2724 , \2718 );
nor \U$2475 ( \2728 , \2726 , \2727 );
not \U$2476 ( \2729 , \2728 );
xor \U$2477 ( \2730 , \2698 , \2704 );
xor \U$2478 ( \2731 , \2730 , \2707 );
not \U$2479 ( \2732 , \2731 );
and \U$2480 ( \2733 , \2397 , \2379 );
not \U$2481 ( \2734 , \2397 );
and \U$2482 ( \2735 , \2734 , \2380 );
nor \U$2483 ( \2736 , \2733 , \2735 );
not \U$2484 ( \2737 , \2736 );
not \U$2485 ( \2738 , \2376 );
and \U$2486 ( \2739 , \2737 , \2738 );
and \U$2487 ( \2740 , \2736 , \2376 );
nor \U$2488 ( \2741 , \2739 , \2740 );
xor \U$2489 ( \2742 , \2629 , \2630 );
xor \U$2490 ( \2743 , \2742 , \2662 );
and \U$2491 ( \2744 , \2741 , \2743 );
xor \U$2492 ( \2745 , \2672 , \2674 );
xor \U$2493 ( \2746 , \2745 , \2677 );
xor \U$2494 ( \2747 , \2629 , \2630 );
xor \U$2495 ( \2748 , \2747 , \2662 );
and \U$2496 ( \2749 , \2746 , \2748 );
and \U$2497 ( \2750 , \2741 , \2746 );
or \U$2498 ( \2751 , \2744 , \2749 , \2750 );
xor \U$2499 ( \2752 , \2529 , \2540 );
xor \U$2500 ( \2753 , \2752 , \2550 );
not \U$2501 ( \2754 , \2753 );
not \U$2502 ( \2755 , \2754 );
xor \U$2503 ( \2756 , \2605 , \2612 );
xor \U$2504 ( \2757 , \2756 , \2622 );
not \U$2505 ( \2758 , \2757 );
not \U$2506 ( \2759 , \2758 );
or \U$2507 ( \2760 , \2755 , \2759 );
nand \U$2508 ( \2761 , \2757 , \2753 );
and \U$2509 ( \2762 , \2578 , \2589 );
not \U$2510 ( \2763 , \2578 );
and \U$2511 ( \2764 , \2763 , \2590 );
or \U$2512 ( \2765 , \2762 , \2764 );
xnor \U$2513 ( \2766 , \2765 , \2565 );
nand \U$2514 ( \2767 , \2761 , \2766 );
nand \U$2515 ( \2768 , \2760 , \2767 );
and \U$2516 ( \2769 , \2649 , \2659 );
not \U$2517 ( \2770 , \2649 );
and \U$2518 ( \2771 , \2770 , \2660 );
nor \U$2519 ( \2772 , \2769 , \2771 );
xor \U$2520 ( \2773 , \2772 , \2641 );
not \U$2521 ( \2774 , \2773 );
not \U$2522 ( \2775 , \2630 );
and \U$2523 ( \2776 , \1528 , RIbe289a8_32);
and \U$2524 ( \2777 , \1531 , RIbe28930_31);
nor \U$2525 ( \2778 , \2776 , \2777 );
and \U$2526 ( \2779 , \2778 , \293 );
not \U$2527 ( \2780 , \2778 );
and \U$2528 ( \2781 , \2780 , \300 );
nor \U$2529 ( \2782 , \2779 , \2781 );
not \U$2530 ( \2783 , \2782 );
not \U$2531 ( \2784 , RIbe29560_57);
not \U$2532 ( \2785 , \1337 );
or \U$2533 ( \2786 , \2784 , \2785 );
nand \U$2534 ( \2787 , \429 , RIbe28228_16);
nand \U$2535 ( \2788 , \2786 , \2787 );
and \U$2536 ( \2789 , \2788 , \306 );
not \U$2537 ( \2790 , \2788 );
and \U$2538 ( \2791 , \2790 , \313 );
nor \U$2539 ( \2792 , \2789 , \2791 );
not \U$2540 ( \2793 , \2792 );
not \U$2541 ( \2794 , \2793 );
or \U$2542 ( \2795 , \2783 , \2794 );
and \U$2543 ( \2796 , \1516 , RIbe29290_51);
and \U$2544 ( \2797 , \1831 , RIbe28a20_33);
nor \U$2545 ( \2798 , \2796 , \2797 );
and \U$2546 ( \2799 , \2798 , \1362 );
not \U$2547 ( \2800 , \2798 );
and \U$2548 ( \2801 , \2800 , \1663 );
nor \U$2549 ( \2802 , \2799 , \2801 );
nand \U$2550 ( \2803 , \2795 , \2802 );
not \U$2551 ( \2804 , \2782 );
nand \U$2552 ( \2805 , \2792 , \2804 );
nand \U$2553 ( \2806 , \2775 , \2803 , \2805 );
not \U$2554 ( \2807 , \2806 );
or \U$2555 ( \2808 , \2774 , \2807 );
nand \U$2556 ( \2809 , \2803 , \2805 );
nand \U$2557 ( \2810 , \2809 , \2630 );
nand \U$2558 ( \2811 , \2808 , \2810 );
xor \U$2559 ( \2812 , \2768 , \2811 );
not \U$2560 ( \2813 , RIbe29a88_68);
not \U$2561 ( \2814 , \1633 );
or \U$2562 ( \2815 , \2813 , \2814 );
not \U$2563 ( \2816 , \1098 );
not \U$2564 ( \2817 , \2816 );
nand \U$2565 ( \2818 , \2817 , RIbe27d78_6);
nand \U$2566 ( \2819 , \2815 , \2818 );
and \U$2567 ( \2820 , \2819 , \1082 );
not \U$2568 ( \2821 , \2819 );
and \U$2569 ( \2822 , \2821 , \1309 );
nor \U$2570 ( \2823 , \2820 , \2822 );
not \U$2571 ( \2824 , RIbe28fc0_45);
not \U$2572 ( \2825 , \1143 );
or \U$2573 ( \2826 , \2824 , \2825 );
nand \U$2574 ( \2827 , \1147 , RIbe290b0_47);
nand \U$2575 ( \2828 , \2826 , \2827 );
not \U$2576 ( \2829 , \2828 );
not \U$2577 ( \2830 , \1157 );
and \U$2578 ( \2831 , \2829 , \2830 );
and \U$2579 ( \2832 , \2828 , \1157 );
nor \U$2580 ( \2833 , \2831 , \2832 );
nand \U$2581 ( \2834 , \2823 , \2833 );
and \U$2582 ( \2835 , \2557 , RIbe27d00_5);
and \U$2583 ( \2836 , \1117 , RIbe27c10_3);
nor \U$2584 ( \2837 , \2835 , \2836 );
and \U$2585 ( \2838 , \2837 , \2563 );
not \U$2586 ( \2839 , \2837 );
and \U$2587 ( \2840 , \2839 , \1132 );
nor \U$2588 ( \2841 , \2838 , \2840 );
and \U$2589 ( \2842 , \2834 , \2841 );
nor \U$2590 ( \2843 , \2833 , \2823 );
nor \U$2591 ( \2844 , \2842 , \2843 );
not \U$2592 ( \2845 , \2844 );
not \U$2593 ( \2846 , RIbe281b0_15);
not \U$2594 ( \2847 , \548 );
or \U$2595 ( \2848 , \2846 , \2847 );
nand \U$2596 ( \2849 , \554 , RIbe280c0_13);
nand \U$2597 ( \2850 , \2848 , \2849 );
not \U$2598 ( \2851 , \2850 );
not \U$2599 ( \2852 , \1333 );
and \U$2600 ( \2853 , \2851 , \2852 );
and \U$2601 ( \2854 , \2850 , \424 );
nor \U$2602 ( \2855 , \2853 , \2854 );
not \U$2603 ( \2856 , \2855 );
and \U$2604 ( \2857 , \1005 , RIbe29650_59);
and \U$2605 ( \2858 , \1165 , RIbe29038_46);
nor \U$2606 ( \2859 , \2857 , \2858 );
and \U$2607 ( \2860 , \2859 , \1813 );
not \U$2608 ( \2861 , \2859 );
and \U$2609 ( \2862 , \2861 , \1011 );
nor \U$2610 ( \2863 , \2860 , \2862 );
not \U$2611 ( \2864 , \2863 );
not \U$2612 ( \2865 , \2864 );
or \U$2613 ( \2866 , \2856 , \2865 );
not \U$2614 ( \2867 , RIbe29830_63);
not \U$2615 ( \2868 , \664 );
or \U$2616 ( \2869 , \2867 , \2868 );
nand \U$2617 ( \2870 , \1180 , RIbe296c8_60);
nand \U$2618 ( \2871 , \2869 , \2870 );
not \U$2619 ( \2872 , \2871 );
not \U$2620 ( \2873 , \564 );
and \U$2621 ( \2874 , \2872 , \2873 );
and \U$2622 ( \2875 , \2871 , \564 );
nor \U$2623 ( \2876 , \2874 , \2875 );
not \U$2624 ( \2877 , \2876 );
nand \U$2625 ( \2878 , \2866 , \2877 );
not \U$2626 ( \2879 , \2855 );
nand \U$2627 ( \2880 , \2879 , \2863 );
nand \U$2628 ( \2881 , \2878 , \2880 );
or \U$2629 ( \2882 , \2845 , \2881 );
not \U$2630 ( \2883 , RIbe29218_50);
not \U$2631 ( \2884 , RIbe29a10_67);
or \U$2632 ( \2885 , \2883 , \2884 );
nand \U$2633 ( \2886 , \2885 , RIbe29b00_69);
buf \U$2634 ( \2887 , \2886 );
and \U$2635 ( \2888 , \2391 , RIbe28e58_42);
not \U$2636 ( \2889 , \2384 );
not \U$2637 ( \2890 , RIbe28de0_41);
nor \U$2638 ( \2891 , \2889 , \2890 );
nor \U$2639 ( \2892 , \2888 , \2891 );
and \U$2640 ( \2893 , \2892 , \1076 );
not \U$2641 ( \2894 , \2892 );
and \U$2642 ( \2895 , \2894 , \1277 );
nor \U$2643 ( \2896 , \2893 , \2895 );
xor \U$2644 ( \2897 , \2887 , \2896 );
not \U$2645 ( \2898 , \2570 );
and \U$2646 ( \2899 , \2898 , RIbe29920_65);
buf \U$2647 ( \2900 , \2566 );
buf \U$2648 ( \2901 , \2900 );
and \U$2649 ( \2902 , \2901 , RIbe27b98_2);
nor \U$2650 ( \2903 , \2899 , \2902 );
and \U$2651 ( \2904 , \2903 , \2379 );
not \U$2652 ( \2905 , \2903 );
and \U$2653 ( \2906 , \2905 , \2380 );
nor \U$2654 ( \2907 , \2904 , \2906 );
and \U$2655 ( \2908 , \2897 , \2907 );
and \U$2656 ( \2909 , \2887 , \2896 );
or \U$2657 ( \2910 , \2908 , \2909 );
nand \U$2658 ( \2911 , \2882 , \2910 );
nand \U$2659 ( \2912 , \2845 , \2881 );
and \U$2660 ( \2913 , \2911 , \2912 );
not \U$2661 ( \2914 , \2913 );
and \U$2662 ( \2915 , \2812 , \2914 );
and \U$2663 ( \2916 , \2768 , \2811 );
or \U$2664 ( \2917 , \2915 , \2916 );
not \U$2665 ( \2918 , \2917 );
or \U$2666 ( \2919 , \2751 , \2918 );
not \U$2667 ( \2920 , \2918 );
not \U$2668 ( \2921 , \2751 );
or \U$2669 ( \2922 , \2920 , \2921 );
xor \U$2670 ( \2923 , \2686 , \2688 );
xor \U$2671 ( \2924 , \2923 , \2691 );
nand \U$2672 ( \2925 , \2922 , \2924 );
nand \U$2673 ( \2926 , \2919 , \2925 );
xor \U$2674 ( \2927 , \2438 , \2466 );
xor \U$2675 ( \2928 , \2927 , \2492 );
xor \U$2676 ( \2929 , \2926 , \2928 );
xor \U$2677 ( \2930 , \2519 , \2683 );
not \U$2678 ( \2931 , \2694 );
xor \U$2679 ( \2932 , \2930 , \2931 );
not \U$2680 ( \2933 , \2932 );
and \U$2681 ( \2934 , \2929 , \2933 );
and \U$2682 ( \2935 , \2926 , \2928 );
or \U$2683 ( \2936 , \2934 , \2935 );
nand \U$2684 ( \2937 , \2732 , \2936 );
not \U$2685 ( \2938 , \2937 );
not \U$2686 ( \2939 , \2710 );
not \U$2687 ( \2940 , \2717 );
or \U$2688 ( \2941 , \2939 , \2940 );
or \U$2689 ( \2942 , \2717 , \2710 );
nand \U$2690 ( \2943 , \2941 , \2942 );
buf \U$2691 ( \2944 , \2943 );
not \U$2692 ( \2945 , \2944 );
or \U$2693 ( \2946 , \2938 , \2945 );
or \U$2694 ( \2947 , \2937 , \2944 );
nand \U$2695 ( \2948 , \2946 , \2947 );
and \U$2696 ( \2949 , \2297 , \2517 , \2729 , \2948 );
not \U$2697 ( \2950 , \2949 );
not \U$2698 ( \2951 , \951 );
not \U$2699 ( \2952 , \1063 );
and \U$2700 ( \2953 , \2951 , \2952 );
and \U$2701 ( \2954 , \951 , \1063 );
nor \U$2702 ( \2955 , \2953 , \2954 );
xnor \U$2703 ( \2956 , \1061 , \962 );
not \U$2704 ( \2957 , \2956 );
not \U$2705 ( \2958 , \965 );
and \U$2706 ( \2959 , \2957 , \2958 );
and \U$2707 ( \2960 , \2956 , \965 );
nor \U$2708 ( \2961 , \2959 , \2960 );
not \U$2709 ( \2962 , \2961 );
not \U$2710 ( \2963 , \1050 );
not \U$2711 ( \2964 , \1032 );
or \U$2712 ( \2965 , \2963 , \2964 );
or \U$2713 ( \2966 , \1032 , \1050 );
nand \U$2714 ( \2967 , \2965 , \2966 );
not \U$2715 ( \2968 , \2967 );
not \U$2716 ( \2969 , \1039 );
and \U$2717 ( \2970 , \2968 , \2969 );
and \U$2718 ( \2971 , \2967 , \1039 );
nor \U$2719 ( \2972 , \2970 , \2971 );
not \U$2720 ( \2973 , \1013 );
not \U$2721 ( \2974 , \993 );
or \U$2722 ( \2975 , \2973 , \2974 );
or \U$2723 ( \2976 , \993 , \1013 );
nand \U$2724 ( \2977 , \2975 , \2976 );
not \U$2725 ( \2978 , \2977 );
not \U$2726 ( \2979 , \986 );
and \U$2727 ( \2980 , \2978 , \2979 );
and \U$2728 ( \2981 , \2977 , \986 );
nor \U$2729 ( \2982 , \2980 , \2981 );
or \U$2730 ( \2983 , \2972 , \2982 );
not \U$2731 ( \2984 , \2982 );
not \U$2732 ( \2985 , \2972 );
or \U$2733 ( \2986 , \2984 , \2985 );
or \U$2734 ( \2987 , \1022 , \1023 );
nand \U$2735 ( \2988 , \2987 , \1024 );
nand \U$2736 ( \2989 , \2986 , \2988 );
nand \U$2737 ( \2990 , \2983 , \2989 );
xor \U$2738 ( \2991 , \2222 , \1794 );
and \U$2739 ( \2992 , \2991 , \2230 );
and \U$2740 ( \2993 , \2222 , \1794 );
or \U$2741 ( \2994 , \2992 , \2993 );
xor \U$2742 ( \2995 , \2239 , \2246 );
and \U$2743 ( \2996 , \2995 , \2254 );
and \U$2744 ( \2997 , \2239 , \2246 );
or \U$2745 ( \2998 , \2996 , \2997 );
or \U$2746 ( \2999 , \2994 , \2998 );
not \U$2747 ( \3000 , \2998 );
not \U$2748 ( \3001 , \2994 );
or \U$2749 ( \3002 , \3000 , \3001 );
or \U$2750 ( \3003 , \2197 , \2211 );
not \U$2751 ( \3004 , \2211 );
not \U$2752 ( \3005 , \2197 );
or \U$2753 ( \3006 , \3004 , \3005 );
nand \U$2754 ( \3007 , \3006 , \2205 );
nand \U$2755 ( \3008 , \3003 , \3007 );
nand \U$2756 ( \3009 , \3002 , \3008 );
nand \U$2757 ( \3010 , \2999 , \3009 );
xor \U$2758 ( \3011 , \2990 , \3010 );
xor \U$2759 ( \3012 , \746 , \752 );
xor \U$2760 ( \3013 , \3012 , \760 );
xor \U$2761 ( \3014 , \969 , \974 );
xor \U$2762 ( \3015 , \3013 , \3014 );
and \U$2763 ( \3016 , \3011 , \3015 );
and \U$2764 ( \3017 , \2990 , \3010 );
or \U$2765 ( \3018 , \3016 , \3017 );
xor \U$2766 ( \3019 , \763 , \772 );
xor \U$2767 ( \3020 , \3019 , \798 );
xor \U$2768 ( \3021 , \3018 , \3020 );
xor \U$2769 ( \3022 , \979 , \1055 );
xor \U$2770 ( \3023 , \3022 , \1058 );
and \U$2771 ( \3024 , \3021 , \3023 );
and \U$2772 ( \3025 , \3018 , \3020 );
or \U$2773 ( \3026 , \3024 , \3025 );
nand \U$2774 ( \3027 , \2962 , \3026 );
xnor \U$2775 ( \3028 , \2955 , \3027 );
not \U$2776 ( \3029 , \3028 );
xor \U$2777 ( \3030 , \2990 , \3010 );
xor \U$2778 ( \3031 , \3030 , \3015 );
xor \U$2779 ( \3032 , \1015 , \1024 );
xor \U$2780 ( \3033 , \3032 , \1052 );
and \U$2781 ( \3034 , \3031 , \3033 );
not \U$2782 ( \3035 , \3031 );
not \U$2783 ( \3036 , \3033 );
and \U$2784 ( \3037 , \3035 , \3036 );
xor \U$2785 ( \3038 , \2215 , \2231 );
and \U$2786 ( \3039 , \3038 , \2255 );
and \U$2787 ( \3040 , \2215 , \2231 );
or \U$2788 ( \3041 , \3039 , \3040 );
xor \U$2789 ( \3042 , \2177 , \2183 );
and \U$2790 ( \3043 , \3042 , \2188 );
and \U$2791 ( \3044 , \2177 , \2183 );
or \U$2792 ( \3045 , \3043 , \3044 );
xor \U$2793 ( \3046 , \3041 , \3045 );
xnor \U$2794 ( \3047 , \2972 , \2982 );
not \U$2795 ( \3048 , \3047 );
not \U$2796 ( \3049 , \2988 );
and \U$2797 ( \3050 , \3048 , \3049 );
and \U$2798 ( \3051 , \3047 , \2988 );
nor \U$2799 ( \3052 , \3050 , \3051 );
and \U$2800 ( \3053 , \3046 , \3052 );
and \U$2801 ( \3054 , \3041 , \3045 );
or \U$2802 ( \3055 , \3053 , \3054 );
nor \U$2803 ( \3056 , \3037 , \3055 );
nor \U$2804 ( \3057 , \3034 , \3056 );
not \U$2805 ( \3058 , \3057 );
xor \U$2806 ( \3059 , \3018 , \3020 );
xor \U$2807 ( \3060 , \3059 , \3023 );
nand \U$2808 ( \3061 , \3058 , \3060 );
not \U$2809 ( \3062 , \3061 );
not \U$2810 ( \3063 , \3026 );
not \U$2811 ( \3064 , \2961 );
or \U$2812 ( \3065 , \3063 , \3064 );
or \U$2813 ( \3066 , \2961 , \3026 );
nand \U$2814 ( \3067 , \3065 , \3066 );
not \U$2815 ( \3068 , \3067 );
or \U$2816 ( \3069 , \3062 , \3068 );
or \U$2817 ( \3070 , \3067 , \3061 );
nand \U$2818 ( \3071 , \3069 , \3070 );
not \U$2819 ( \3072 , \3057 );
not \U$2820 ( \3073 , \3060 );
or \U$2821 ( \3074 , \3072 , \3073 );
or \U$2822 ( \3075 , \3060 , \3057 );
nand \U$2823 ( \3076 , \3074 , \3075 );
xor \U$2824 ( \3077 , \3041 , \3045 );
xor \U$2825 ( \3078 , \3077 , \3052 );
not \U$2826 ( \3079 , \2994 );
not \U$2827 ( \3080 , \3008 );
or \U$2828 ( \3081 , \3079 , \3080 );
or \U$2829 ( \3082 , \3008 , \2994 );
nand \U$2830 ( \3083 , \3081 , \3082 );
not \U$2831 ( \3084 , \3083 );
not \U$2832 ( \3085 , \2998 );
and \U$2833 ( \3086 , \3084 , \3085 );
and \U$2834 ( \3087 , \3083 , \2998 );
nor \U$2835 ( \3088 , \3086 , \3087 );
or \U$2836 ( \3089 , \3078 , \3088 );
not \U$2837 ( \3090 , \3088 );
not \U$2838 ( \3091 , \3078 );
or \U$2839 ( \3092 , \3090 , \3091 );
or \U$2840 ( \3093 , \2256 , \2077 );
not \U$2841 ( \3094 , \2077 );
not \U$2842 ( \3095 , \2256 );
or \U$2843 ( \3096 , \3094 , \3095 );
nand \U$2844 ( \3097 , \3096 , \2263 );
nand \U$2845 ( \3098 , \3093 , \3097 );
nand \U$2846 ( \3099 , \3092 , \3098 );
nand \U$2847 ( \3100 , \3089 , \3099 );
not \U$2848 ( \3101 , \3031 );
not \U$2849 ( \3102 , \3055 );
not \U$2850 ( \3103 , \3033 );
and \U$2851 ( \3104 , \3102 , \3103 );
and \U$2852 ( \3105 , \3055 , \3033 );
nor \U$2853 ( \3106 , \3104 , \3105 );
not \U$2854 ( \3107 , \3106 );
or \U$2855 ( \3108 , \3101 , \3107 );
or \U$2856 ( \3109 , \3106 , \3031 );
nand \U$2857 ( \3110 , \3108 , \3109 );
and \U$2858 ( \3111 , \3100 , \3110 );
xor \U$2859 ( \3112 , \3076 , \3111 );
nand \U$2860 ( \3113 , \3029 , \3071 , \3112 );
not \U$2861 ( \3114 , \3113 );
not \U$2862 ( \3115 , \3088 );
not \U$2863 ( \3116 , \3098 );
or \U$2864 ( \3117 , \3115 , \3116 );
or \U$2865 ( \3118 , \3098 , \3088 );
nand \U$2866 ( \3119 , \3117 , \3118 );
not \U$2867 ( \3120 , \3119 );
not \U$2868 ( \3121 , \3078 );
and \U$2869 ( \3122 , \3120 , \3121 );
and \U$2870 ( \3123 , \3078 , \3119 );
nor \U$2871 ( \3124 , \3122 , \3123 );
xor \U$2872 ( \3125 , \2173 , \2189 );
and \U$2873 ( \3126 , \3125 , \2272 );
and \U$2874 ( \3127 , \2173 , \2189 );
or \U$2875 ( \3128 , \3126 , \3127 );
xor \U$2876 ( \3129 , \3124 , \3128 );
xor \U$2877 ( \3130 , \2273 , \2275 );
not \U$2878 ( \3131 , \2280 );
and \U$2879 ( \3132 , \3130 , \3131 );
and \U$2880 ( \3133 , \2273 , \2275 );
or \U$2881 ( \3134 , \3132 , \3133 );
xnor \U$2882 ( \3135 , \3129 , \3134 );
not \U$2883 ( \3136 , \2282 );
nand \U$2884 ( \3137 , \3136 , \2289 );
xor \U$2885 ( \3138 , \3135 , \3137 );
not \U$2886 ( \3139 , \3124 );
not \U$2887 ( \3140 , \3128 );
and \U$2888 ( \3141 , \3139 , \3140 );
and \U$2889 ( \3142 , \3124 , \3128 );
nor \U$2890 ( \3143 , \3142 , \3134 );
nor \U$2891 ( \3144 , \3141 , \3143 );
xor \U$2892 ( \3145 , \3100 , \3110 );
xor \U$2893 ( \3146 , \3144 , \3145 );
nor \U$2894 ( \3147 , \3138 , \3146 );
nand \U$2895 ( \3148 , \3114 , \3147 );
nor \U$2896 ( \3149 , \2950 , \3148 );
not \U$2897 ( \3150 , \3149 );
and \U$2898 ( \3151 , \327 , RIbe28b10_35);
and \U$2899 ( \3152 , \1371 , RIbe28b88_36);
nor \U$2900 ( \3153 , \3151 , \3152 );
and \U$2901 ( \3154 , \3153 , \339 );
not \U$2902 ( \3155 , \3153 );
and \U$2903 ( \3156 , \3155 , \342 );
nor \U$2904 ( \3157 , \3154 , \3156 );
and \U$2905 ( \3158 , RIbe29380_53, RIbe28408_20);
not \U$2906 ( \3159 , \3158 );
buf \U$2907 ( \3160 , \324 );
and \U$2908 ( \3161 , \3160 , RIbe28390_19);
and \U$2909 ( \3162 , \1371 , RIbe28b10_35);
nor \U$2910 ( \3163 , \3161 , \3162 );
and \U$2911 ( \3164 , \3163 , \1375 );
not \U$2912 ( \3165 , \3163 );
and \U$2913 ( \3166 , \3165 , \1379 );
nor \U$2914 ( \3167 , \3164 , \3166 );
nand \U$2915 ( \3168 , \3159 , \3167 );
xor \U$2916 ( \3169 , \3157 , \3168 );
not \U$2917 ( \3170 , RIbe28930_31);
not \U$2918 ( \3171 , \1774 );
or \U$2919 ( \3172 , \3170 , \3171 );
nand \U$2920 ( \3173 , \429 , RIbe29560_57);
nand \U$2921 ( \3174 , \3172 , \3173 );
not \U$2922 ( \3175 , \1231 );
and \U$2923 ( \3176 , \3174 , \3175 );
not \U$2924 ( \3177 , \3174 );
and \U$2925 ( \3178 , \3177 , \306 );
nor \U$2926 ( \3179 , \3176 , \3178 );
and \U$2927 ( \3180 , \1516 , RIbe28b88_36);
and \U$2928 ( \3181 , \1831 , RIbe29290_51);
nor \U$2929 ( \3182 , \3180 , \3181 );
and \U$2930 ( \3183 , \3182 , \1663 );
not \U$2931 ( \3184 , \3182 );
and \U$2932 ( \3185 , \3184 , \1362 );
nor \U$2933 ( \3186 , \3183 , \3185 );
or \U$2934 ( \3187 , \3179 , \3186 );
not \U$2935 ( \3188 , \3186 );
not \U$2936 ( \3189 , \3179 );
or \U$2937 ( \3190 , \3188 , \3189 );
and \U$2938 ( \3191 , \1679 , RIbe28a20_33);
and \U$2939 ( \3192 , \1682 , RIbe289a8_32);
nor \U$2940 ( \3193 , \3191 , \3192 );
and \U$2941 ( \3194 , \3193 , \300 );
not \U$2942 ( \3195 , \3193 );
and \U$2943 ( \3196 , \3195 , \293 );
nor \U$2944 ( \3197 , \3194 , \3196 );
nand \U$2945 ( \3198 , \3190 , \3197 );
nand \U$2946 ( \3199 , \3187 , \3198 );
and \U$2947 ( \3200 , \3169 , \3199 );
and \U$2948 ( \3201 , \3157 , \3168 );
or \U$2949 ( \3202 , \3200 , \3201 );
not \U$2950 ( \3203 , \3202 );
and \U$2951 ( \3204 , \1286 , RIbe27d78_6);
and \U$2952 ( \3205 , \1117 , RIbe27d00_5);
nor \U$2953 ( \3206 , \3204 , \3205 );
and \U$2954 ( \3207 , \3206 , \1131 );
not \U$2955 ( \3208 , \3206 );
and \U$2956 ( \3209 , \3208 , \1448 );
nor \U$2957 ( \3210 , \3207 , \3209 );
not \U$2958 ( \3211 , RIbe290b0_47);
not \U$2959 ( \3212 , \1094 );
or \U$2960 ( \3213 , \3211 , \3212 );
nand \U$2961 ( \3214 , \2817 , RIbe29a88_68);
nand \U$2962 ( \3215 , \3213 , \3214 );
and \U$2963 ( \3216 , \3215 , \1309 );
not \U$2964 ( \3217 , \3215 );
and \U$2965 ( \3218 , \3217 , \1082 );
nor \U$2966 ( \3219 , \3216 , \3218 );
not \U$2967 ( \3220 , \3219 );
and \U$2968 ( \3221 , \3210 , \3220 );
not \U$2969 ( \3222 , \1143 );
not \U$2970 ( \3223 , \3222 );
not \U$2971 ( \3224 , \2355 );
and \U$2972 ( \3225 , \3223 , \3224 );
and \U$2973 ( \3226 , \1147 , RIbe28fc0_45);
nor \U$2974 ( \3227 , \3225 , \3226 );
and \U$2975 ( \3228 , \3227 , \1154 );
not \U$2976 ( \3229 , \3227 );
and \U$2977 ( \3230 , \3229 , \1157 );
nor \U$2978 ( \3231 , \3228 , \3230 );
nor \U$2979 ( \3232 , \3221 , \3231 );
nor \U$2980 ( \3233 , \3220 , \3210 );
nor \U$2981 ( \3234 , \3232 , \3233 );
not \U$2982 ( \3235 , \3234 );
and \U$2983 ( \3236 , \2425 , RIbe296c8_60);
and \U$2984 ( \3237 , \2000 , RIbe29650_59);
nor \U$2985 ( \3238 , \3236 , \3237 );
and \U$2986 ( \3239 , \3238 , \1608 );
not \U$2987 ( \3240 , \3238 );
and \U$2988 ( \3241 , \3240 , \1011 );
nor \U$2989 ( \3242 , \3239 , \3241 );
not \U$2990 ( \3243 , \3242 );
not \U$2991 ( \3244 , \547 );
and \U$2992 ( \3245 , \3244 , RIbe28228_16);
and \U$2993 ( \3246 , \553 , RIbe281b0_15);
nor \U$2994 ( \3247 , \3245 , \3246 );
and \U$2995 ( \3248 , \3247 , \1330 );
not \U$2996 ( \3249 , \3247 );
and \U$2997 ( \3250 , \3249 , \1246 );
nor \U$2998 ( \3251 , \3248 , \3250 );
and \U$2999 ( \3252 , \3243 , \3251 );
and \U$3000 ( \3253 , \664 , RIbe280c0_13);
not \U$3001 ( \3254 , RIbe29830_63);
nor \U$3002 ( \3255 , \3254 , \1611 );
nor \U$3003 ( \3256 , \3253 , \3255 );
and \U$3004 ( \3257 , \3256 , \1621 );
not \U$3005 ( \3258 , \3256 );
and \U$3006 ( \3259 , \3258 , \564 );
nor \U$3007 ( \3260 , \3257 , \3259 );
nor \U$3008 ( \3261 , \3252 , \3260 );
nor \U$3009 ( \3262 , \3243 , \3251 );
nor \U$3010 ( \3263 , \3261 , \3262 );
not \U$3011 ( \3264 , \3263 );
and \U$3012 ( \3265 , \3235 , \3264 );
and \U$3013 ( \3266 , \3234 , \3263 );
buf \U$3014 ( \3267 , \2900 );
and \U$3015 ( \3268 , \3267 , RIbe29920_65);
not \U$3016 ( \3269 , \2898 );
nor \U$3017 ( \3270 , \3269 , \2890 );
nor \U$3018 ( \3271 , \3268 , \3270 );
not \U$3019 ( \3272 , \2379 );
and \U$3020 ( \3273 , \3271 , \3272 );
not \U$3021 ( \3274 , \3271 );
not \U$3022 ( \3275 , \3272 );
and \U$3023 ( \3276 , \3274 , \3275 );
nor \U$3024 ( \3277 , \3273 , \3276 );
not \U$3025 ( \3278 , \3277 );
xor \U$3026 ( \3279 , RIbe29a10_67, RIbe29218_50);
not \U$3027 ( \3280 , \3279 );
xor \U$3028 ( \3281 , RIbe29a10_67, RIbe29b00_69);
nand \U$3029 ( \3282 , \3280 , \3281 );
buf \U$3030 ( \3283 , \3282 );
not \U$3031 ( \3284 , \3283 );
buf \U$3032 ( \3285 , \3284 );
nand \U$3033 ( \3286 , \3285 , RIbe27b98_2);
and \U$3034 ( \3287 , RIbe29a10_67, RIbe29218_50);
not \U$3035 ( \3288 , RIbe29b00_69);
nor \U$3036 ( \3289 , \3287 , \3288 );
buf \U$3037 ( \3290 , \3289 );
and \U$3038 ( \3291 , \3286 , \3290 );
not \U$3039 ( \3292 , \3286 );
and \U$3040 ( \3293 , \3292 , \2887 );
nor \U$3041 ( \3294 , \3291 , \3293 );
not \U$3042 ( \3295 , \3294 );
and \U$3043 ( \3296 , \3278 , \3295 );
and \U$3044 ( \3297 , \3277 , \3294 );
not \U$3045 ( \3298 , \2889 );
not \U$3046 ( \3299 , RIbe28e58_42);
not \U$3047 ( \3300 , \3299 );
and \U$3048 ( \3301 , \3298 , \3300 );
not \U$3049 ( \3302 , \2583 );
not \U$3050 ( \3303 , \3302 );
and \U$3051 ( \3304 , \3303 , RIbe27c10_3);
nor \U$3052 ( \3305 , \3301 , \3304 );
and \U$3053 ( \3306 , \3305 , \1277 );
not \U$3054 ( \3307 , \3305 );
and \U$3055 ( \3308 , \3307 , \1076 );
nor \U$3056 ( \3309 , \3306 , \3308 );
nor \U$3057 ( \3310 , \3297 , \3309 );
nor \U$3058 ( \3311 , \3296 , \3310 );
nor \U$3059 ( \3312 , \3266 , \3311 );
nor \U$3060 ( \3313 , \3265 , \3312 );
nand \U$3061 ( \3314 , \3203 , \3313 );
and \U$3062 ( \3315 , RIbe28390_19, RIbe29380_53);
not \U$3063 ( \3316 , \2793 );
not \U$3064 ( \3317 , \2804 );
or \U$3065 ( \3318 , \3316 , \3317 );
nand \U$3066 ( \3319 , \2792 , \2782 );
nand \U$3067 ( \3320 , \3318 , \3319 );
xor \U$3068 ( \3321 , \2802 , \3320 );
xor \U$3069 ( \3322 , \3315 , \3321 );
not \U$3070 ( \3323 , \2855 );
not \U$3071 ( \3324 , \2876 );
not \U$3072 ( \3325 , \2863 );
or \U$3073 ( \3326 , \3324 , \3325 );
or \U$3074 ( \3327 , \2863 , \2876 );
nand \U$3075 ( \3328 , \3326 , \3327 );
not \U$3076 ( \3329 , \3328 );
or \U$3077 ( \3330 , \3323 , \3329 );
or \U$3078 ( \3331 , \3328 , \2855 );
nand \U$3079 ( \3332 , \3330 , \3331 );
and \U$3080 ( \3333 , \3322 , \3332 );
and \U$3081 ( \3334 , \3315 , \3321 );
or \U$3082 ( \3335 , \3333 , \3334 );
and \U$3083 ( \3336 , \3314 , \3335 );
not \U$3084 ( \3337 , \3313 );
and \U$3085 ( \3338 , \3337 , \3202 );
nor \U$3086 ( \3339 , \3336 , \3338 );
xor \U$3087 ( \3340 , \2553 , \2593 );
xor \U$3088 ( \3341 , \3340 , \2625 );
xor \U$3089 ( \3342 , \3339 , \3341 );
nand \U$3090 ( \3343 , \2806 , \2810 );
xor \U$3091 ( \3344 , \3343 , \2773 );
xor \U$3092 ( \3345 , \2881 , \2844 );
xor \U$3093 ( \3346 , \3345 , \2910 );
nand \U$3094 ( \3347 , \3344 , \3346 );
xnor \U$3095 ( \3348 , \2758 , \2766 );
not \U$3096 ( \3349 , \3348 );
not \U$3097 ( \3350 , \2754 );
and \U$3098 ( \3351 , \3349 , \3350 );
and \U$3099 ( \3352 , \3348 , \2754 );
nor \U$3100 ( \3353 , \3351 , \3352 );
not \U$3101 ( \3354 , \3353 );
and \U$3102 ( \3355 , \3347 , \3354 );
nor \U$3103 ( \3356 , \3344 , \3346 );
nor \U$3104 ( \3357 , \3355 , \3356 );
xor \U$3105 ( \3358 , \3342 , \3357 );
xor \U$3106 ( \3359 , \2768 , \2811 );
not \U$3107 ( \3360 , \2913 );
xor \U$3108 ( \3361 , \3359 , \3360 );
xor \U$3109 ( \3362 , \2629 , \2630 );
xor \U$3110 ( \3363 , \3362 , \2662 );
xor \U$3111 ( \3364 , \2741 , \2746 );
xor \U$3112 ( \3365 , \3363 , \3364 );
and \U$3113 ( \3366 , \3361 , \3365 );
nor \U$3114 ( \3367 , \3361 , \3365 );
nor \U$3115 ( \3368 , \3366 , \3367 );
xor \U$3116 ( \3369 , \3358 , \3368 );
xor \U$3117 ( \3370 , \2823 , \2841 );
xor \U$3118 ( \3371 , \3370 , \2833 );
xor \U$3119 ( \3372 , \2887 , \2896 );
xor \U$3120 ( \3373 , \3372 , \2907 );
and \U$3121 ( \3374 , \3371 , \3373 );
xor \U$3122 ( \3375 , \3315 , \3321 );
xor \U$3123 ( \3376 , \3375 , \3332 );
xor \U$3124 ( \3377 , \2887 , \2896 );
xor \U$3125 ( \3378 , \3377 , \2907 );
and \U$3126 ( \3379 , \3376 , \3378 );
and \U$3127 ( \3380 , \3371 , \3376 );
or \U$3128 ( \3381 , \3374 , \3379 , \3380 );
not \U$3129 ( \3382 , \3158 );
not \U$3130 ( \3383 , \3167 );
not \U$3131 ( \3384 , \3383 );
or \U$3132 ( \3385 , \3382 , \3384 );
nand \U$3133 ( \3386 , \3385 , \3168 );
not \U$3134 ( \3387 , RIbe28408_20);
not \U$3135 ( \3388 , \324 );
or \U$3136 ( \3389 , \3387 , \3388 );
nand \U$3137 ( \3390 , \329 , RIbe28390_19);
nand \U$3138 ( \3391 , \3389 , \3390 );
not \U$3139 ( \3392 , \3391 );
not \U$3140 ( \3393 , \1374 );
and \U$3141 ( \3394 , \3392 , \3393 );
and \U$3142 ( \3395 , \3391 , \1379 );
nor \U$3143 ( \3396 , \3394 , \3395 );
nand \U$3144 ( \3397 , RIbe29380_53, RIbe28480_21);
nand \U$3145 ( \3398 , \3396 , \3397 );
and \U$3146 ( \3399 , \1516 , RIbe28b10_35);
and \U$3147 ( \3400 , \264 , RIbe28b88_36);
nor \U$3148 ( \3401 , \3399 , \3400 );
and \U$3149 ( \3402 , \3401 , \1362 );
not \U$3150 ( \3403 , \3401 );
and \U$3151 ( \3404 , \3403 , \269 );
nor \U$3152 ( \3405 , \3402 , \3404 );
nand \U$3153 ( \3406 , \3398 , \3405 );
or \U$3154 ( \3407 , \3397 , \3396 );
nand \U$3155 ( \3408 , \3406 , \3407 );
xor \U$3156 ( \3409 , \3386 , \3408 );
not \U$3157 ( \3410 , RIbe29560_57);
not \U$3158 ( \3411 , \1756 );
or \U$3159 ( \3412 , \3410 , \3411 );
nand \U$3160 ( \3413 , \552 , RIbe28228_16);
nand \U$3161 ( \3414 , \3412 , \3413 );
not \U$3162 ( \3415 , \424 );
and \U$3163 ( \3416 , \3414 , \3415 );
not \U$3164 ( \3417 , \3414 );
and \U$3165 ( \3418 , \3417 , \1333 );
nor \U$3166 ( \3419 , \3416 , \3418 );
not \U$3167 ( \3420 , \382 );
not \U$3168 ( \3421 , RIbe289a8_32);
not \U$3169 ( \3422 , \3421 );
and \U$3170 ( \3423 , \3420 , \3422 );
and \U$3171 ( \3424 , \429 , RIbe28930_31);
nor \U$3172 ( \3425 , \3423 , \3424 );
and \U$3173 ( \3426 , \3425 , \313 );
not \U$3174 ( \3427 , \3425 );
and \U$3175 ( \3428 , \3427 , \306 );
nor \U$3176 ( \3429 , \3426 , \3428 );
xor \U$3177 ( \3430 , \3419 , \3429 );
and \U$3178 ( \3431 , \1254 , RIbe29290_51);
and \U$3179 ( \3432 , \1682 , RIbe28a20_33);
nor \U$3180 ( \3433 , \3431 , \3432 );
and \U$3181 ( \3434 , \3433 , \300 );
not \U$3182 ( \3435 , \3433 );
and \U$3183 ( \3436 , \3435 , \293 );
nor \U$3184 ( \3437 , \3434 , \3436 );
and \U$3185 ( \3438 , \3430 , \3437 );
and \U$3186 ( \3439 , \3419 , \3429 );
or \U$3187 ( \3440 , \3438 , \3439 );
and \U$3188 ( \3441 , \3409 , \3440 );
and \U$3189 ( \3442 , \3386 , \3408 );
or \U$3190 ( \3443 , \3441 , \3442 );
not \U$3191 ( \3444 , RIbe27c88_4);
not \U$3192 ( \3445 , RIbe27df0_7);
or \U$3193 ( \3446 , \3444 , \3445 );
nand \U$3194 ( \3447 , \3446 , RIbe29218_50);
buf \U$3195 ( \3448 , \3447 );
not \U$3196 ( \3449 , \3448 );
not \U$3197 ( \3450 , RIbe29920_65);
not \U$3198 ( \3451 , \3282 );
buf \U$3199 ( \3452 , \3451 );
not \U$3200 ( \3453 , \3452 );
or \U$3201 ( \3454 , \3450 , \3453 );
not \U$3202 ( \3455 , \3279 );
not \U$3203 ( \3456 , \3455 );
buf \U$3204 ( \3457 , \3456 );
buf \U$3205 ( \3458 , \3457 );
nand \U$3206 ( \3459 , \3458 , RIbe27b98_2);
nand \U$3207 ( \3460 , \3454 , \3459 );
buf \U$3208 ( \3461 , \2887 );
and \U$3209 ( \3462 , \3460 , \3461 );
not \U$3210 ( \3463 , \3460 );
and \U$3211 ( \3464 , \3463 , \3290 );
nor \U$3212 ( \3465 , \3462 , \3464 );
not \U$3213 ( \3466 , \3465 );
not \U$3214 ( \3467 , \3466 );
or \U$3215 ( \3468 , \3449 , \3467 );
nand \U$3216 ( \3469 , RIbe27df0_7, RIbe27c88_4);
and \U$3217 ( \3470 , \3469 , RIbe29218_50);
buf \U$3218 ( \3471 , \3470 );
not \U$3219 ( \3472 , \3471 );
not \U$3220 ( \3473 , \3465 );
or \U$3221 ( \3474 , \3472 , \3473 );
not \U$3222 ( \3475 , RIbe28e58_42);
not \U$3223 ( \3476 , \2570 );
not \U$3224 ( \3477 , \3476 );
or \U$3225 ( \3478 , \3475 , \3477 );
nand \U$3226 ( \3479 , \3267 , RIbe28de0_41);
nand \U$3227 ( \3480 , \3478 , \3479 );
not \U$3228 ( \3481 , \2576 );
and \U$3229 ( \3482 , \3480 , \3481 );
not \U$3230 ( \3483 , \3480 );
and \U$3231 ( \3484 , \3483 , \2379 );
nor \U$3232 ( \3485 , \3482 , \3484 );
nand \U$3233 ( \3486 , \3474 , \3485 );
nand \U$3234 ( \3487 , \3468 , \3486 );
and \U$3235 ( \3488 , \1113 , RIbe29a88_68);
and \U$3236 ( \3489 , \1117 , RIbe27d78_6);
nor \U$3237 ( \3490 , \3488 , \3489 );
not \U$3238 ( \3491 , \1124 );
and \U$3239 ( \3492 , \3490 , \3491 );
not \U$3240 ( \3493 , \3490 );
and \U$3241 ( \3494 , \3493 , \1131 );
nor \U$3242 ( \3495 , \3492 , \3494 );
not \U$3243 ( \3496 , \3495 );
not \U$3244 ( \3497 , RIbe28fc0_45);
not \U$3245 ( \3498 , \1094 );
or \U$3246 ( \3499 , \3497 , \3498 );
nand \U$3247 ( \3500 , \1455 , RIbe290b0_47);
nand \U$3248 ( \3501 , \3499 , \3500 );
and \U$3249 ( \3502 , \3501 , \1082 );
not \U$3250 ( \3503 , \3501 );
and \U$3251 ( \3504 , \3503 , \1309 );
nor \U$3252 ( \3505 , \3502 , \3504 );
not \U$3253 ( \3506 , \3505 );
not \U$3254 ( \3507 , \3506 );
or \U$3255 ( \3508 , \3496 , \3507 );
not \U$3256 ( \3509 , RIbe27d00_5);
not \U$3257 ( \3510 , \3303 );
or \U$3258 ( \3511 , \3509 , \3510 );
nand \U$3259 ( \3512 , \2384 , RIbe27c10_3);
nand \U$3260 ( \3513 , \3511 , \3512 );
not \U$3261 ( \3514 , \3513 );
not \U$3262 ( \3515 , \1075 );
not \U$3263 ( \3516 , \3515 );
not \U$3264 ( \3517 , \3516 );
and \U$3265 ( \3518 , \3514 , \3517 );
and \U$3266 ( \3519 , \3513 , \1076 );
nor \U$3267 ( \3520 , \3518 , \3519 );
not \U$3268 ( \3521 , \3520 );
not \U$3269 ( \3522 , \3495 );
nand \U$3270 ( \3523 , \3522 , \3505 );
nand \U$3271 ( \3524 , \3521 , \3523 );
nand \U$3272 ( \3525 , \3508 , \3524 );
or \U$3273 ( \3526 , \3487 , \3525 );
not \U$3274 ( \3527 , RIbe29650_59);
not \U$3275 ( \3528 , \1143 );
or \U$3276 ( \3529 , \3527 , \3528 );
nand \U$3277 ( \3530 , \1147 , RIbe29038_46);
nand \U$3278 ( \3531 , \3529 , \3530 );
and \U$3279 ( \3532 , \3531 , \1652 );
not \U$3280 ( \3533 , \3531 );
and \U$3281 ( \3534 , \3533 , \1152 );
nor \U$3282 ( \3535 , \3532 , \3534 );
not \U$3283 ( \3536 , \1611 );
not \U$3284 ( \3537 , RIbe280c0_13);
not \U$3285 ( \3538 , \3537 );
and \U$3286 ( \3539 , \3536 , \3538 );
and \U$3287 ( \3540 , \664 , RIbe281b0_15);
nor \U$3288 ( \3541 , \3539 , \3540 );
and \U$3289 ( \3542 , \3541 , \672 );
not \U$3290 ( \3543 , \3541 );
and \U$3291 ( \3544 , \3543 , \564 );
or \U$3292 ( \3545 , \3542 , \3544 );
xor \U$3293 ( \3546 , \3535 , \3545 );
and \U$3294 ( \3547 , \1005 , RIbe29830_63);
and \U$3295 ( \3548 , \1203 , RIbe296c8_60);
nor \U$3296 ( \3549 , \3547 , \3548 );
and \U$3297 ( \3550 , \3549 , \752 );
not \U$3298 ( \3551 , \3549 );
and \U$3299 ( \3552 , \3551 , \1011 );
nor \U$3300 ( \3553 , \3550 , \3552 );
and \U$3301 ( \3554 , \3546 , \3553 );
and \U$3302 ( \3555 , \3535 , \3545 );
or \U$3303 ( \3556 , \3554 , \3555 );
nand \U$3304 ( \3557 , \3526 , \3556 );
nand \U$3305 ( \3558 , \3487 , \3525 );
nand \U$3306 ( \3559 , \3557 , \3558 );
xor \U$3307 ( \3560 , \3443 , \3559 );
and \U$3308 ( \3561 , \3210 , \3219 );
not \U$3309 ( \3562 , \3210 );
and \U$3310 ( \3563 , \3562 , \3220 );
or \U$3311 ( \3564 , \3561 , \3563 );
xnor \U$3312 ( \3565 , \3564 , \3231 );
and \U$3313 ( \3566 , \3260 , \3242 );
not \U$3314 ( \3567 , \3260 );
and \U$3315 ( \3568 , \3567 , \3243 );
or \U$3316 ( \3569 , \3566 , \3568 );
xnor \U$3317 ( \3570 , \3569 , \3251 );
xor \U$3318 ( \3571 , \3565 , \3570 );
not \U$3319 ( \3572 , \3186 );
not \U$3320 ( \3573 , \3197 );
not \U$3321 ( \3574 , \3179 );
or \U$3322 ( \3575 , \3573 , \3574 );
or \U$3323 ( \3576 , \3179 , \3197 );
nand \U$3324 ( \3577 , \3575 , \3576 );
not \U$3325 ( \3578 , \3577 );
or \U$3326 ( \3579 , \3572 , \3578 );
or \U$3327 ( \3580 , \3577 , \3186 );
nand \U$3328 ( \3581 , \3579 , \3580 );
and \U$3329 ( \3582 , \3571 , \3581 );
and \U$3330 ( \3583 , \3565 , \3570 );
or \U$3331 ( \3584 , \3582 , \3583 );
and \U$3332 ( \3585 , \3560 , \3584 );
and \U$3333 ( \3586 , \3443 , \3559 );
or \U$3334 ( \3587 , \3585 , \3586 );
xor \U$3335 ( \3588 , \3381 , \3587 );
not \U$3336 ( \3589 , \3356 );
nand \U$3337 ( \3590 , \3589 , \3347 );
not \U$3338 ( \3591 , \3590 );
not \U$3339 ( \3592 , \3353 );
and \U$3340 ( \3593 , \3591 , \3592 );
and \U$3341 ( \3594 , \3590 , \3353 );
nor \U$3342 ( \3595 , \3593 , \3594 );
and \U$3343 ( \3596 , \3588 , \3595 );
and \U$3344 ( \3597 , \3381 , \3587 );
nor \U$3345 ( \3598 , \3596 , \3597 );
and \U$3346 ( \3599 , \3369 , \3598 );
and \U$3347 ( \3600 , \3358 , \3368 );
or \U$3348 ( \3601 , \3599 , \3600 );
xnor \U$3349 ( \3602 , \2918 , \2751 );
and \U$3350 ( \3603 , \3602 , \2924 );
nor \U$3351 ( \3604 , \3602 , \2924 );
nor \U$3352 ( \3605 , \3603 , \3604 );
xor \U$3353 ( \3606 , \3601 , \3605 );
not \U$3354 ( \3607 , \3365 );
nand \U$3355 ( \3608 , \3607 , \3361 );
xor \U$3356 ( \3609 , \2628 , \2665 );
xor \U$3357 ( \3610 , \3609 , \2680 );
xor \U$3358 ( \3611 , \3608 , \3610 );
xor \U$3359 ( \3612 , \3339 , \3341 );
and \U$3360 ( \3613 , \3612 , \3357 );
and \U$3361 ( \3614 , \3339 , \3341 );
or \U$3362 ( \3615 , \3613 , \3614 );
and \U$3363 ( \3616 , \3611 , \3615 );
nor \U$3364 ( \3617 , \3611 , \3615 );
nor \U$3365 ( \3618 , \3616 , \3617 );
xor \U$3366 ( \3619 , \3606 , \3618 );
not \U$3367 ( \3620 , \3619 );
not \U$3368 ( \3621 , \3311 );
xor \U$3369 ( \3622 , \3234 , \3263 );
not \U$3370 ( \3623 , \3622 );
or \U$3371 ( \3624 , \3621 , \3623 );
or \U$3372 ( \3625 , \3622 , \3311 );
nand \U$3373 ( \3626 , \3624 , \3625 );
xor \U$3374 ( \3627 , \2887 , \2896 );
xor \U$3375 ( \3628 , \3627 , \2907 );
xor \U$3376 ( \3629 , \3371 , \3376 );
xor \U$3377 ( \3630 , \3628 , \3629 );
xor \U$3378 ( \3631 , \3626 , \3630 );
xor \U$3379 ( \3632 , \3443 , \3559 );
xor \U$3380 ( \3633 , \3632 , \3584 );
and \U$3381 ( \3634 , \3631 , \3633 );
and \U$3382 ( \3635 , \3626 , \3630 );
or \U$3383 ( \3636 , \3634 , \3635 );
not \U$3384 ( \3637 , \3335 );
xnor \U$3385 ( \3638 , \3337 , \3202 );
not \U$3386 ( \3639 , \3638 );
or \U$3387 ( \3640 , \3637 , \3639 );
or \U$3388 ( \3641 , \3638 , \3335 );
nand \U$3389 ( \3642 , \3640 , \3641 );
xor \U$3390 ( \3643 , \3636 , \3642 );
not \U$3391 ( \3644 , RIbe296c8_60);
not \U$3392 ( \3645 , \1143 );
or \U$3393 ( \3646 , \3644 , \3645 );
nand \U$3394 ( \3647 , \1147 , RIbe29650_59);
nand \U$3395 ( \3648 , \3646 , \3647 );
and \U$3396 ( \3649 , \3648 , \1152 );
not \U$3397 ( \3650 , \3648 );
and \U$3398 ( \3651 , \3650 , \1469 );
nor \U$3399 ( \3652 , \3649 , \3651 );
and \U$3400 ( \3653 , \2425 , RIbe280c0_13);
and \U$3401 ( \3654 , \2000 , RIbe29830_63);
nor \U$3402 ( \3655 , \3653 , \3654 );
and \U$3403 ( \3656 , \3655 , \1608 );
not \U$3404 ( \3657 , \3655 );
and \U$3405 ( \3658 , \3657 , \1011 );
nor \U$3406 ( \3659 , \3656 , \3658 );
not \U$3407 ( \3660 , \3659 );
nand \U$3408 ( \3661 , \3652 , \3660 );
not \U$3409 ( \3662 , \1611 );
not \U$3410 ( \3663 , RIbe281b0_15);
not \U$3411 ( \3664 , \3663 );
and \U$3412 ( \3665 , \3662 , \3664 );
and \U$3413 ( \3666 , \666 , RIbe28228_16);
nor \U$3414 ( \3667 , \3665 , \3666 );
and \U$3415 ( \3668 , \3667 , \564 );
not \U$3416 ( \3669 , \3667 );
and \U$3417 ( \3670 , \3669 , \672 );
nor \U$3418 ( \3671 , \3668 , \3670 );
and \U$3419 ( \3672 , \3661 , \3671 );
nor \U$3420 ( \3673 , \3652 , \3660 );
nor \U$3421 ( \3674 , \3672 , \3673 );
not \U$3422 ( \3675 , RIbe27c10_3);
not \U$3423 ( \3676 , \2898 );
or \U$3424 ( \3677 , \3675 , \3676 );
nand \U$3425 ( \3678 , \2901 , RIbe28e58_42);
nand \U$3426 ( \3679 , \3677 , \3678 );
and \U$3427 ( \3680 , \3679 , \2379 );
not \U$3428 ( \3681 , \3679 );
and \U$3429 ( \3682 , \3681 , \3272 );
nor \U$3430 ( \3683 , \3680 , \3682 );
not \U$3431 ( \3684 , RIbe28de0_41);
not \U$3432 ( \3685 , \3283 );
not \U$3433 ( \3686 , \3685 );
or \U$3434 ( \3687 , \3684 , \3686 );
buf \U$3435 ( \3688 , \3280 );
not \U$3436 ( \3689 , \3688 );
nand \U$3437 ( \3690 , \3689 , RIbe29920_65);
nand \U$3438 ( \3691 , \3687 , \3690 );
and \U$3439 ( \3692 , \3691 , \3461 );
not \U$3440 ( \3693 , \3691 );
and \U$3441 ( \3694 , \3693 , \3290 );
nor \U$3442 ( \3695 , \3692 , \3694 );
nand \U$3443 ( \3696 , \3683 , \3695 );
not \U$3444 ( \3697 , \3447 );
not \U$3445 ( \3698 , \3697 );
not \U$3446 ( \3699 , \3698 );
xnor \U$3447 ( \3700 , RIbe27df0_7, RIbe27c88_4);
xor \U$3448 ( \3701 , RIbe29218_50, RIbe27df0_7);
nand \U$3449 ( \3702 , \3700 , \3701 );
buf \U$3450 ( \3703 , \3702 );
nor \U$3451 ( \3704 , \3703 , \1640 );
not \U$3452 ( \3705 , \3704 );
or \U$3453 ( \3706 , \3699 , \3705 );
or \U$3454 ( \3707 , \3704 , \3448 );
nand \U$3455 ( \3708 , \3706 , \3707 );
and \U$3456 ( \3709 , \3696 , \3708 );
nor \U$3457 ( \3710 , \3683 , \3695 );
nor \U$3458 ( \3711 , \3709 , \3710 );
or \U$3459 ( \3712 , \3674 , \3711 );
not \U$3460 ( \3713 , \3711 );
not \U$3461 ( \3714 , \3674 );
or \U$3462 ( \3715 , \3713 , \3714 );
not \U$3463 ( \3716 , RIbe29038_46);
not \U$3464 ( \3717 , \1094 );
or \U$3465 ( \3718 , \3716 , \3717 );
nand \U$3466 ( \3719 , \1455 , RIbe28fc0_45);
nand \U$3467 ( \3720 , \3718 , \3719 );
and \U$3468 ( \3721 , \3720 , \1082 );
not \U$3469 ( \3722 , \3720 );
and \U$3470 ( \3723 , \3722 , \1309 );
nor \U$3471 ( \3724 , \3721 , \3723 );
not \U$3472 ( \3725 , \3724 );
and \U$3473 ( \3726 , \2557 , RIbe290b0_47);
and \U$3474 ( \3727 , \1117 , RIbe29a88_68);
nor \U$3475 ( \3728 , \3726 , \3727 );
and \U$3476 ( \3729 , \3728 , \2563 );
not \U$3477 ( \3730 , \3728 );
and \U$3478 ( \3731 , \3730 , \1132 );
nor \U$3479 ( \3732 , \3729 , \3731 );
not \U$3480 ( \3733 , \3732 );
not \U$3481 ( \3734 , \3733 );
or \U$3482 ( \3735 , \3725 , \3734 );
and \U$3483 ( \3736 , \1272 , RIbe27d78_6);
not \U$3484 ( \3737 , RIbe27d00_5);
nor \U$3485 ( \3738 , \3737 , \2889 );
nor \U$3486 ( \3739 , \3736 , \3738 );
and \U$3487 ( \3740 , \3739 , \1277 );
not \U$3488 ( \3741 , \3739 );
and \U$3489 ( \3742 , \3741 , \1076 );
nor \U$3490 ( \3743 , \3740 , \3742 );
not \U$3491 ( \3744 , \3743 );
nand \U$3492 ( \3745 , \3735 , \3744 );
not \U$3493 ( \3746 , \3724 );
nand \U$3494 ( \3747 , \3746 , \3732 );
nand \U$3495 ( \3748 , \3745 , \3747 );
nand \U$3496 ( \3749 , \3715 , \3748 );
nand \U$3497 ( \3750 , \3712 , \3749 );
not \U$3498 ( \3751 , RIbe28a20_33);
not \U$3499 ( \3752 , \1774 );
or \U$3500 ( \3753 , \3751 , \3752 );
nand \U$3501 ( \3754 , \429 , RIbe289a8_32);
nand \U$3502 ( \3755 , \3753 , \3754 );
and \U$3503 ( \3756 , \3755 , \313 );
not \U$3504 ( \3757 , \3755 );
and \U$3505 ( \3758 , \3757 , \306 );
nor \U$3506 ( \3759 , \3756 , \3758 );
not \U$3507 ( \3760 , RIbe28b88_36);
not \U$3508 ( \3761 , \1528 );
or \U$3509 ( \3762 , \3760 , \3761 );
nand \U$3510 ( \3763 , \1682 , RIbe29290_51);
nand \U$3511 ( \3764 , \3762 , \3763 );
not \U$3512 ( \3765 , \3764 );
not \U$3513 ( \3766 , \300 );
and \U$3514 ( \3767 , \3765 , \3766 );
and \U$3515 ( \3768 , \3764 , \300 );
nor \U$3516 ( \3769 , \3767 , \3768 );
and \U$3517 ( \3770 , \3759 , \3769 );
not \U$3518 ( \3771 , RIbe28930_31);
not \U$3519 ( \3772 , \548 );
or \U$3520 ( \3773 , \3771 , \3772 );
not \U$3521 ( \3774 , \552 );
not \U$3522 ( \3775 , \3774 );
nand \U$3523 ( \3776 , \3775 , RIbe29560_57);
nand \U$3524 ( \3777 , \3773 , \3776 );
not \U$3525 ( \3778 , \3777 );
not \U$3526 ( \3779 , \1333 );
and \U$3527 ( \3780 , \3778 , \3779 );
and \U$3528 ( \3781 , \3777 , \424 );
nor \U$3529 ( \3782 , \3780 , \3781 );
nor \U$3530 ( \3783 , \3770 , \3782 );
nor \U$3531 ( \3784 , \3759 , \3769 );
nor \U$3532 ( \3785 , \3783 , \3784 );
not \U$3533 ( \3786 , \3785 );
xor \U$3534 ( \3787 , \3397 , \3396 );
xnor \U$3535 ( \3788 , \3787 , \3405 );
not \U$3536 ( \3789 , \3788 );
or \U$3537 ( \3790 , \3786 , \3789 );
nand \U$3538 ( \3791 , RIbe29380_53, RIbe287c8_28);
not \U$3539 ( \3792 , \3791 );
and \U$3540 ( \3793 , \1357 , RIbe28390_19);
and \U$3541 ( \3794 , \264 , RIbe28b10_35);
nor \U$3542 ( \3795 , \3793 , \3794 );
and \U$3543 ( \3796 , \3795 , \1663 );
not \U$3544 ( \3797 , \3795 );
and \U$3545 ( \3798 , \3797 , \1362 );
nor \U$3546 ( \3799 , \3796 , \3798 );
not \U$3547 ( \3800 , \3799 );
or \U$3548 ( \3801 , \3792 , \3800 );
and \U$3549 ( \3802 , \325 , RIbe28480_21);
and \U$3550 ( \3803 , \330 , RIbe28408_20);
nor \U$3551 ( \3804 , \3802 , \3803 );
and \U$3552 ( \3805 , \3804 , \1375 );
not \U$3553 ( \3806 , \3804 );
and \U$3554 ( \3807 , \3806 , \1374 );
nor \U$3555 ( \3808 , \3805 , \3807 );
not \U$3556 ( \3809 , \3808 );
nand \U$3557 ( \3810 , \3801 , \3809 );
not \U$3558 ( \3811 , \3791 );
not \U$3559 ( \3812 , \3799 );
nand \U$3560 ( \3813 , \3811 , \3812 );
nand \U$3561 ( \3814 , \3810 , \3813 );
nand \U$3562 ( \3815 , \3790 , \3814 );
or \U$3563 ( \3816 , \3785 , \3788 );
nand \U$3564 ( \3817 , \3815 , \3816 );
xor \U$3565 ( \3818 , \3750 , \3817 );
xor \U$3566 ( \3819 , \3419 , \3429 );
xor \U$3567 ( \3820 , \3819 , \3437 );
xor \U$3568 ( \3821 , \3535 , \3545 );
xor \U$3569 ( \3822 , \3821 , \3553 );
xor \U$3570 ( \3823 , \3820 , \3822 );
not \U$3571 ( \3824 , \3520 );
not \U$3572 ( \3825 , \3495 );
or \U$3573 ( \3826 , \3824 , \3825 );
or \U$3574 ( \3827 , \3495 , \3520 );
nand \U$3575 ( \3828 , \3826 , \3827 );
and \U$3576 ( \3829 , \3828 , \3506 );
not \U$3577 ( \3830 , \3828 );
and \U$3578 ( \3831 , \3830 , \3505 );
nor \U$3579 ( \3832 , \3829 , \3831 );
and \U$3580 ( \3833 , \3823 , \3832 );
and \U$3581 ( \3834 , \3820 , \3822 );
or \U$3582 ( \3835 , \3833 , \3834 );
and \U$3583 ( \3836 , \3818 , \3835 );
and \U$3584 ( \3837 , \3750 , \3817 );
or \U$3585 ( \3838 , \3836 , \3837 );
xor \U$3586 ( \3839 , \3157 , \3168 );
xor \U$3587 ( \3840 , \3839 , \3199 );
xor \U$3588 ( \3841 , \3838 , \3840 );
not \U$3589 ( \3842 , \3309 );
xor \U$3590 ( \3843 , \3277 , \3294 );
not \U$3591 ( \3844 , \3843 );
or \U$3592 ( \3845 , \3842 , \3844 );
or \U$3593 ( \3846 , \3843 , \3309 );
nand \U$3594 ( \3847 , \3845 , \3846 );
xor \U$3595 ( \3848 , \3386 , \3408 );
xor \U$3596 ( \3849 , \3848 , \3440 );
xor \U$3597 ( \3850 , \3847 , \3849 );
xor \U$3598 ( \3851 , \3565 , \3570 );
xor \U$3599 ( \3852 , \3851 , \3581 );
and \U$3600 ( \3853 , \3850 , \3852 );
and \U$3601 ( \3854 , \3847 , \3849 );
or \U$3602 ( \3855 , \3853 , \3854 );
and \U$3603 ( \3856 , \3841 , \3855 );
and \U$3604 ( \3857 , \3838 , \3840 );
or \U$3605 ( \3858 , \3856 , \3857 );
and \U$3606 ( \3859 , \3643 , \3858 );
and \U$3607 ( \3860 , \3636 , \3642 );
or \U$3608 ( \3861 , \3859 , \3860 );
not \U$3609 ( \3862 , \3861 );
xor \U$3610 ( \3863 , \3358 , \3368 );
xor \U$3611 ( \3864 , \3863 , \3598 );
nand \U$3612 ( \3865 , \3862 , \3864 );
not \U$3613 ( \3866 , \3865 );
xor \U$3614 ( \3867 , \3381 , \3587 );
xor \U$3615 ( \3868 , \3867 , \3595 );
xor \U$3616 ( \3869 , \3636 , \3642 );
xor \U$3617 ( \3870 , \3869 , \3858 );
xor \U$3618 ( \3871 , \3868 , \3870 );
not \U$3619 ( \3872 , \3485 );
xor \U$3620 ( \3873 , \3471 , \3290 );
xor \U$3621 ( \3874 , \3873 , \3460 );
not \U$3622 ( \3875 , \3874 );
or \U$3623 ( \3876 , \3872 , \3875 );
or \U$3624 ( \3877 , \3485 , \3874 );
nand \U$3625 ( \3878 , \3876 , \3877 );
not \U$3626 ( \3879 , \3878 );
xor \U$3627 ( \3880 , \3785 , \3814 );
xnor \U$3628 ( \3881 , \3880 , \3788 );
nand \U$3629 ( \3882 , \3879 , \3881 );
xor \U$3630 ( \3883 , \3820 , \3822 );
xor \U$3631 ( \3884 , \3883 , \3832 );
and \U$3632 ( \3885 , \3882 , \3884 );
not \U$3633 ( \3886 , \3878 );
nor \U$3634 ( \3887 , \3886 , \3881 );
nor \U$3635 ( \3888 , \3885 , \3887 );
xor \U$3636 ( \3889 , \3525 , \3487 );
xnor \U$3637 ( \3890 , \3889 , \3556 );
or \U$3638 ( \3891 , \3888 , \3890 );
not \U$3639 ( \3892 , \3890 );
not \U$3640 ( \3893 , \3888 );
or \U$3641 ( \3894 , \3892 , \3893 );
not \U$3642 ( \3895 , \282 );
and \U$3643 ( \3896 , \3895 , RIbe28b10_35);
not \U$3644 ( \3897 , \286 );
and \U$3645 ( \3898 , \3897 , RIbe28b88_36);
nor \U$3646 ( \3899 , \3896 , \3898 );
and \U$3647 ( \3900 , \3899 , \293 );
not \U$3648 ( \3901 , \3899 );
and \U$3649 ( \3902 , \3901 , \300 );
nor \U$3650 ( \3903 , \3900 , \3902 );
not \U$3651 ( \3904 , \3903 );
not \U$3652 ( \3905 , \3904 );
and \U$3653 ( \3906 , \1659 , RIbe28408_20);
and \U$3654 ( \3907 , \1831 , RIbe28390_19);
nor \U$3655 ( \3908 , \3906 , \3907 );
and \U$3656 ( \3909 , \3908 , \270 );
not \U$3657 ( \3910 , \3908 );
and \U$3658 ( \3911 , \3910 , \1663 );
nor \U$3659 ( \3912 , \3909 , \3911 );
not \U$3660 ( \3913 , \3912 );
or \U$3661 ( \3914 , \3905 , \3913 );
not \U$3662 ( \3915 , \3912 );
nand \U$3663 ( \3916 , \3903 , \3915 );
not \U$3664 ( \3917 , \339 );
not \U$3665 ( \3918 , RIbe287c8_28);
not \U$3666 ( \3919 , \326 );
or \U$3667 ( \3920 , \3918 , \3919 );
nand \U$3668 ( \3921 , \330 , RIbe28480_21);
nand \U$3669 ( \3922 , \3920 , \3921 );
not \U$3670 ( \3923 , \3922 );
or \U$3671 ( \3924 , \3917 , \3923 );
or \U$3672 ( \3925 , \3922 , \339 );
nand \U$3673 ( \3926 , \3924 , \3925 );
nand \U$3674 ( \3927 , \3916 , \3926 );
nand \U$3675 ( \3928 , \3914 , \3927 );
not \U$3676 ( \3929 , \3928 );
not \U$3677 ( \3930 , RIbe29290_51);
not \U$3678 ( \3931 , \1337 );
or \U$3679 ( \3932 , \3930 , \3931 );
nand \U$3680 ( \3933 , \429 , RIbe28a20_33);
nand \U$3681 ( \3934 , \3932 , \3933 );
not \U$3682 ( \3935 , \3934 );
not \U$3683 ( \3936 , \313 );
and \U$3684 ( \3937 , \3935 , \3936 );
and \U$3685 ( \3938 , \3934 , \3175 );
nor \U$3686 ( \3939 , \3937 , \3938 );
not \U$3687 ( \3940 , RIbe289a8_32);
not \U$3688 ( \3941 , \548 );
or \U$3689 ( \3942 , \3940 , \3941 );
nand \U$3690 ( \3943 , \553 , RIbe28930_31);
nand \U$3691 ( \3944 , \3942 , \3943 );
not \U$3692 ( \3945 , \3944 );
not \U$3693 ( \3946 , \1333 );
and \U$3694 ( \3947 , \3945 , \3946 );
and \U$3695 ( \3948 , \3944 , \1764 );
nor \U$3696 ( \3949 , \3947 , \3948 );
and \U$3697 ( \3950 , \3939 , \3949 );
not \U$3698 ( \3951 , \1611 );
not \U$3699 ( \3952 , RIbe28228_16);
not \U$3700 ( \3953 , \3952 );
and \U$3701 ( \3954 , \3951 , \3953 );
and \U$3702 ( \3955 , \666 , RIbe29560_57);
nor \U$3703 ( \3956 , \3954 , \3955 );
and \U$3704 ( \3957 , \3956 , \564 );
not \U$3705 ( \3958 , \3956 );
buf \U$3706 ( \3959 , \670 );
and \U$3707 ( \3960 , \3958 , \3959 );
nor \U$3708 ( \3961 , \3957 , \3960 );
not \U$3709 ( \3962 , \3961 );
nor \U$3710 ( \3963 , \3950 , \3962 );
nor \U$3711 ( \3964 , \3939 , \3949 );
nor \U$3712 ( \3965 , \3963 , \3964 );
nand \U$3713 ( \3966 , \3929 , \3965 );
not \U$3714 ( \3967 , RIbe281b0_15);
not \U$3715 ( \3968 , \2425 );
or \U$3716 ( \3969 , \3967 , \3968 );
nand \U$3717 ( \3970 , \1203 , RIbe280c0_13);
nand \U$3718 ( \3971 , \3969 , \3970 );
not \U$3719 ( \3972 , \3971 );
not \U$3720 ( \3973 , \1813 );
and \U$3721 ( \3974 , \3972 , \3973 );
and \U$3722 ( \3975 , \3971 , \1608 );
nor \U$3723 ( \3976 , \3974 , \3975 );
not \U$3724 ( \3977 , RIbe29650_59);
not \U$3725 ( \3978 , \1094 );
or \U$3726 ( \3979 , \3977 , \3978 );
nand \U$3727 ( \3980 , \1455 , RIbe29038_46);
nand \U$3728 ( \3981 , \3979 , \3980 );
and \U$3729 ( \3982 , \3981 , \1309 );
not \U$3730 ( \3983 , \3981 );
and \U$3731 ( \3984 , \3983 , \1082 );
nor \U$3732 ( \3985 , \3982 , \3984 );
not \U$3733 ( \3986 , \3985 );
and \U$3734 ( \3987 , \3976 , \3986 );
not \U$3735 ( \3988 , RIbe29830_63);
not \U$3736 ( \3989 , \1143 );
or \U$3737 ( \3990 , \3988 , \3989 );
nand \U$3738 ( \3991 , \1147 , RIbe296c8_60);
nand \U$3739 ( \3992 , \3990 , \3991 );
not \U$3740 ( \3993 , \1152 );
not \U$3741 ( \3994 , \3993 );
and \U$3742 ( \3995 , \3992 , \3994 );
not \U$3743 ( \3996 , \3992 );
and \U$3744 ( \3997 , \3996 , \3993 );
nor \U$3745 ( \3998 , \3995 , \3997 );
nor \U$3746 ( \3999 , \3987 , \3998 );
nor \U$3747 ( \4000 , \3986 , \3976 );
nor \U$3748 ( \4001 , \3999 , \4000 );
not \U$3749 ( \4002 , \4001 );
and \U$3750 ( \4003 , RIbe28d68_40, RIbe29998_66);
not \U$3751 ( \4004 , RIbe27c88_4);
nor \U$3752 ( \4005 , \4003 , \4004 );
not \U$3753 ( \4006 , \4005 );
not \U$3754 ( \4007 , \4006 );
not \U$3755 ( \4008 , RIbe28e58_42);
not \U$3756 ( \4009 , \3685 );
or \U$3757 ( \4010 , \4008 , \4009 );
not \U$3758 ( \4011 , \3688 );
nand \U$3759 ( \4012 , \4011 , RIbe28de0_41);
nand \U$3760 ( \4013 , \4010 , \4012 );
not \U$3761 ( \4014 , \4013 );
not \U$3762 ( \4015 , \2887 );
and \U$3763 ( \4016 , \4014 , \4015 );
and \U$3764 ( \4017 , \4013 , \2887 );
nor \U$3765 ( \4018 , \4016 , \4017 );
xor \U$3766 ( \4019 , \4007 , \4018 );
not \U$3767 ( \4020 , RIbe29920_65);
not \U$3768 ( \4021 , \3703 );
not \U$3769 ( \4022 , \4021 );
or \U$3770 ( \4023 , \4020 , \4022 );
xor \U$3771 ( \4024 , RIbe27df0_7, RIbe27c88_4);
not \U$3772 ( \4025 , \4024 );
not \U$3773 ( \4026 , \4025 );
buf \U$3774 ( \4027 , \4026 );
nand \U$3775 ( \4028 , \4027 , RIbe27b98_2);
nand \U$3776 ( \4029 , \4023 , \4028 );
and \U$3777 ( \4030 , \4029 , \3448 );
not \U$3778 ( \4031 , \4029 );
and \U$3779 ( \4032 , \4031 , \3471 );
nor \U$3780 ( \4033 , \4030 , \4032 );
and \U$3781 ( \4034 , \4019 , \4033 );
and \U$3782 ( \4035 , \4007 , \4018 );
or \U$3783 ( \4036 , \4034 , \4035 );
not \U$3784 ( \4037 , \4036 );
or \U$3785 ( \4038 , \4002 , \4037 );
not \U$3786 ( \4039 , RIbe28fc0_45);
not \U$3787 ( \4040 , \1113 );
or \U$3788 ( \4041 , \4039 , \4040 );
nand \U$3789 ( \4042 , \1117 , RIbe290b0_47);
nand \U$3790 ( \4043 , \4041 , \4042 );
not \U$3791 ( \4044 , \4043 );
not \U$3792 ( \4045 , \3491 );
and \U$3793 ( \4046 , \4044 , \4045 );
and \U$3794 ( \4047 , \4043 , \1125 );
nor \U$3795 ( \4048 , \4046 , \4047 );
not \U$3796 ( \4049 , RIbe27d00_5);
not \U$3797 ( \4050 , \2570 );
buf \U$3798 ( \4051 , \4050 );
not \U$3799 ( \4052 , \4051 );
or \U$3800 ( \4053 , \4049 , \4052 );
nand \U$3801 ( \4054 , \3267 , RIbe27c10_3);
nand \U$3802 ( \4055 , \4053 , \4054 );
and \U$3803 ( \4056 , \4055 , \2380 );
not \U$3804 ( \4057 , \4055 );
not \U$3805 ( \4058 , \2379 );
not \U$3806 ( \4059 , \4058 );
and \U$3807 ( \4060 , \4057 , \4059 );
nor \U$3808 ( \4061 , \4056 , \4060 );
not \U$3809 ( \4062 , \4061 );
and \U$3810 ( \4063 , \4048 , \4062 );
not \U$3811 ( \4064 , \2384 );
buf \U$3812 ( \4065 , \4064 );
not \U$3813 ( \4066 , \4065 );
not \U$3814 ( \4067 , \255 );
and \U$3815 ( \4068 , \4066 , \4067 );
and \U$3816 ( \4069 , \2391 , RIbe29a88_68);
nor \U$3817 ( \4070 , \4068 , \4069 );
and \U$3818 ( \4071 , \4070 , \1277 );
not \U$3819 ( \4072 , \4070 );
and \U$3820 ( \4073 , \4072 , \3516 );
nor \U$3821 ( \4074 , \4071 , \4073 );
nor \U$3822 ( \4075 , \4063 , \4074 );
nor \U$3823 ( \4076 , \4048 , \4062 );
nor \U$3824 ( \4077 , \4075 , \4076 );
not \U$3825 ( \4078 , \4077 );
nand \U$3826 ( \4079 , \4038 , \4078 );
or \U$3827 ( \4080 , \4036 , \4001 );
nand \U$3828 ( \4081 , \4079 , \4080 );
xor \U$3829 ( \4082 , \3966 , \4081 );
xor \U$3830 ( \4083 , \3791 , \3808 );
xnor \U$3831 ( \4084 , \4083 , \3812 );
xor \U$3832 ( \4085 , \3782 , \3759 );
xor \U$3833 ( \4086 , \4085 , \3769 );
or \U$3834 ( \4087 , \4084 , \4086 );
not \U$3835 ( \4088 , \4086 );
not \U$3836 ( \4089 , \4084 );
or \U$3837 ( \4090 , \4088 , \4089 );
and \U$3838 ( \4091 , \3652 , \3659 );
not \U$3839 ( \4092 , \3652 );
and \U$3840 ( \4093 , \4092 , \3660 );
or \U$3841 ( \4094 , \4091 , \4093 );
xor \U$3842 ( \4095 , \4094 , \3671 );
nand \U$3843 ( \4096 , \4090 , \4095 );
nand \U$3844 ( \4097 , \4087 , \4096 );
and \U$3845 ( \4098 , \4082 , \4097 );
and \U$3846 ( \4099 , \3966 , \4081 );
or \U$3847 ( \4100 , \4098 , \4099 );
nand \U$3848 ( \4101 , \3894 , \4100 );
nand \U$3849 ( \4102 , \3891 , \4101 );
xor \U$3850 ( \4103 , \3838 , \3840 );
xor \U$3851 ( \4104 , \4103 , \3855 );
xor \U$3852 ( \4105 , \4102 , \4104 );
xor \U$3853 ( \4106 , \3626 , \3630 );
xor \U$3854 ( \4107 , \4106 , \3633 );
and \U$3855 ( \4108 , \4105 , \4107 );
and \U$3856 ( \4109 , \4102 , \4104 );
or \U$3857 ( \4110 , \4108 , \4109 );
and \U$3858 ( \4111 , \3871 , \4110 );
and \U$3859 ( \4112 , \3868 , \3870 );
or \U$3860 ( \4113 , \4111 , \4112 );
not \U$3861 ( \4114 , \4113 );
or \U$3862 ( \4115 , \3866 , \4114 );
not \U$3863 ( \4116 , \3864 );
nand \U$3864 ( \4117 , \4116 , \3861 );
nand \U$3865 ( \4118 , \4115 , \4117 );
not \U$3866 ( \4119 , \4118 );
or \U$3867 ( \4120 , \3620 , \4119 );
or \U$3868 ( \4121 , \4118 , \3619 );
nand \U$3869 ( \4122 , \4120 , \4121 );
not \U$3870 ( \4123 , \2936 );
not \U$3871 ( \4124 , \2731 );
or \U$3872 ( \4125 , \4123 , \4124 );
or \U$3873 ( \4126 , \2731 , \2936 );
nand \U$3874 ( \4127 , \4125 , \4126 );
or \U$3875 ( \4128 , \3608 , \3610 );
and \U$3876 ( \4129 , \3608 , \3610 );
nor \U$3877 ( \4130 , \4129 , \3615 );
not \U$3878 ( \4131 , \4130 );
nand \U$3879 ( \4132 , \4128 , \4131 );
xor \U$3880 ( \4133 , \2926 , \2928 );
xor \U$3881 ( \4134 , \4133 , \2933 );
and \U$3882 ( \4135 , \4132 , \4134 );
xor \U$3883 ( \4136 , \4127 , \4135 );
xor \U$3884 ( \4137 , \4132 , \4134 );
xor \U$3885 ( \4138 , \3601 , \3605 );
and \U$3886 ( \4139 , \4138 , \3618 );
and \U$3887 ( \4140 , \3601 , \3605 );
or \U$3888 ( \4141 , \4139 , \4140 );
xnor \U$3889 ( \4142 , \4137 , \4141 );
nand \U$3890 ( \4143 , \4122 , \4136 , \4142 );
nand \U$3891 ( \4144 , \3915 , \3904 );
nand \U$3892 ( \4145 , \3903 , \3912 );
nand \U$3893 ( \4146 , \4144 , \4145 );
xor \U$3894 ( \4147 , \4146 , \3926 );
not \U$3895 ( \4148 , \4147 );
and \U$3896 ( \4149 , RIbe29380_53, RIbe285e8_24);
not \U$3897 ( \4150 , \4149 );
and \U$3898 ( \4151 , \4148 , \4150 );
xor \U$3899 ( \4152 , \3949 , \3961 );
xnor \U$3900 ( \4153 , \4152 , \3939 );
nor \U$3901 ( \4154 , \4151 , \4153 );
and \U$3902 ( \4155 , \4149 , \4147 );
nor \U$3903 ( \4156 , \4154 , \4155 );
nand \U$3904 ( \4157 , RIbe29380_53, RIbe28660_25);
not \U$3905 ( \4158 , \4157 );
and \U$3906 ( \4159 , \3895 , RIbe28390_19);
and \U$3907 ( \4160 , \1682 , RIbe28b10_35);
nor \U$3908 ( \4161 , \4159 , \4160 );
and \U$3909 ( \4162 , \4161 , \293 );
not \U$3910 ( \4163 , \4161 );
and \U$3911 ( \4164 , \4163 , \300 );
nor \U$3912 ( \4165 , \4162 , \4164 );
not \U$3913 ( \4166 , RIbe285e8_24);
not \U$3914 ( \4167 , \3160 );
or \U$3915 ( \4168 , \4166 , \4167 );
nand \U$3916 ( \4169 , \329 , RIbe287c8_28);
nand \U$3917 ( \4170 , \4168 , \4169 );
not \U$3918 ( \4171 , \4170 );
not \U$3919 ( \4172 , \338 );
not \U$3920 ( \4173 , \4172 );
and \U$3921 ( \4174 , \4171 , \4173 );
and \U$3922 ( \4175 , \4170 , \1374 );
nor \U$3923 ( \4176 , \4174 , \4175 );
nand \U$3924 ( \4177 , \4165 , \4176 );
and \U$3925 ( \4178 , \260 , RIbe28480_21);
and \U$3926 ( \4179 , \264 , RIbe28408_20);
nor \U$3927 ( \4180 , \4178 , \4179 );
and \U$3928 ( \4181 , \4180 , \1362 );
not \U$3929 ( \4182 , \4180 );
and \U$3930 ( \4183 , \4182 , \1663 );
nor \U$3931 ( \4184 , \4181 , \4183 );
and \U$3932 ( \4185 , \4177 , \4184 );
nor \U$3933 ( \4186 , \4165 , \4176 );
nor \U$3934 ( \4187 , \4185 , \4186 );
not \U$3935 ( \4188 , \4187 );
or \U$3936 ( \4189 , \4158 , \4188 );
not \U$3937 ( \4190 , RIbe28a20_33);
not \U$3938 ( \4191 , \3244 );
or \U$3939 ( \4192 , \4190 , \4191 );
nand \U$3940 ( \4193 , \1327 , RIbe289a8_32);
nand \U$3941 ( \4194 , \4192 , \4193 );
and \U$3942 ( \4195 , \4194 , \3415 );
not \U$3943 ( \4196 , \4194 );
and \U$3944 ( \4197 , \4196 , \424 );
nor \U$3945 ( \4198 , \4195 , \4197 );
not \U$3946 ( \4199 , \4198 );
not \U$3947 ( \4200 , RIbe28b88_36);
not \U$3948 ( \4201 , \1223 );
or \U$3949 ( \4202 , \4200 , \4201 );
nand \U$3950 ( \4203 , \429 , RIbe29290_51);
nand \U$3951 ( \4204 , \4202 , \4203 );
not \U$3952 ( \4205 , \4204 );
not \U$3953 ( \4206 , \3175 );
and \U$3954 ( \4207 , \4205 , \4206 );
and \U$3955 ( \4208 , \4204 , \3175 );
nor \U$3956 ( \4209 , \4207 , \4208 );
and \U$3957 ( \4210 , \4199 , \4209 );
not \U$3958 ( \4211 , RIbe28930_31);
not \U$3959 ( \4212 , \664 );
or \U$3960 ( \4213 , \4211 , \4212 );
nand \U$3961 ( \4214 , \1180 , RIbe29560_57);
nand \U$3962 ( \4215 , \4213 , \4214 );
not \U$3963 ( \4216 , \4215 );
not \U$3964 ( \4217 , \1617 );
not \U$3965 ( \4218 , \4217 );
and \U$3966 ( \4219 , \4216 , \4218 );
and \U$3967 ( \4220 , \4215 , \564 );
nor \U$3968 ( \4221 , \4219 , \4220 );
nor \U$3969 ( \4222 , \4210 , \4221 );
nor \U$3970 ( \4223 , \4199 , \4209 );
nor \U$3971 ( \4224 , \4222 , \4223 );
not \U$3972 ( \4225 , \4224 );
nand \U$3973 ( \4226 , \4189 , \4225 );
not \U$3974 ( \4227 , \4187 );
not \U$3975 ( \4228 , \4157 );
nand \U$3976 ( \4229 , \4227 , \4228 );
and \U$3977 ( \4230 , \4226 , \4229 );
nand \U$3978 ( \4231 , \4156 , \4230 );
not \U$3979 ( \4232 , RIbe28228_16);
not \U$3980 ( \4233 , \1807 );
or \U$3981 ( \4234 , \4232 , \4233 );
nand \U$3982 ( \4235 , \1203 , RIbe281b0_15);
nand \U$3983 ( \4236 , \4234 , \4235 );
not \U$3984 ( \4237 , \4236 );
not \U$3985 ( \4238 , \1813 );
and \U$3986 ( \4239 , \4237 , \4238 );
and \U$3987 ( \4240 , \4236 , \1608 );
nor \U$3988 ( \4241 , \4239 , \4240 );
not \U$3989 ( \4242 , \4241 );
not \U$3990 ( \4243 , RIbe296c8_60);
not \U$3991 ( \4244 , \1633 );
or \U$3992 ( \4245 , \4243 , \4244 );
nand \U$3993 ( \4246 , \1099 , RIbe29650_59);
nand \U$3994 ( \4247 , \4245 , \4246 );
not \U$3995 ( \4248 , \4247 );
not \U$3996 ( \4249 , \2418 );
and \U$3997 ( \4250 , \4248 , \4249 );
not \U$3998 ( \4251 , \1081 );
and \U$3999 ( \4252 , \4247 , \4251 );
nor \U$4000 ( \4253 , \4250 , \4252 );
not \U$4001 ( \4254 , \4253 );
or \U$4002 ( \4255 , \4242 , \4254 );
not \U$4003 ( \4256 , RIbe280c0_13);
not \U$4004 ( \4257 , \2596 );
not \U$4005 ( \4258 , \4257 );
or \U$4006 ( \4259 , \4256 , \4258 );
nand \U$4007 ( \4260 , \1147 , RIbe29830_63);
nand \U$4008 ( \4261 , \4259 , \4260 );
and \U$4009 ( \4262 , \4261 , \1469 );
not \U$4010 ( \4263 , \4261 );
and \U$4011 ( \4264 , \4263 , \1157 );
nor \U$4012 ( \4265 , \4262 , \4264 );
nand \U$4013 ( \4266 , \4255 , \4265 );
not \U$4014 ( \4267 , \4253 );
not \U$4015 ( \4268 , \4241 );
nand \U$4016 ( \4269 , \4267 , \4268 );
nand \U$4017 ( \4270 , \4266 , \4269 );
not \U$4018 ( \4271 , \4270 );
not \U$4019 ( \4272 , \4271 );
and \U$4020 ( \4273 , \1286 , RIbe29038_46);
and \U$4021 ( \4274 , \1117 , RIbe28fc0_45);
nor \U$4022 ( \4275 , \4273 , \4274 );
and \U$4023 ( \4276 , \4275 , \1131 );
not \U$4024 ( \4277 , \4275 );
and \U$4025 ( \4278 , \4277 , \1448 );
nor \U$4026 ( \4279 , \4276 , \4278 );
not \U$4027 ( \4280 , \4279 );
not \U$4028 ( \4281 , RIbe27d78_6);
not \U$4029 ( \4282 , \4051 );
or \U$4030 ( \4283 , \4281 , \4282 );
buf \U$4031 ( \4284 , \2900 );
nand \U$4032 ( \4285 , \4284 , RIbe27d00_5);
nand \U$4033 ( \4286 , \4283 , \4285 );
not \U$4034 ( \4287 , \2576 );
and \U$4035 ( \4288 , \4286 , \4287 );
not \U$4036 ( \4289 , \4286 );
and \U$4037 ( \4290 , \4289 , \2576 );
nor \U$4038 ( \4291 , \4288 , \4290 );
not \U$4039 ( \4292 , \4291 );
not \U$4040 ( \4293 , \4292 );
or \U$4041 ( \4294 , \4280 , \4293 );
not \U$4042 ( \4295 , \1271 );
and \U$4043 ( \4296 , \4295 , RIbe290b0_47);
not \U$4044 ( \4297 , RIbe29a88_68);
nor \U$4045 ( \4298 , \4297 , \4065 );
nor \U$4046 ( \4299 , \4296 , \4298 );
and \U$4047 ( \4300 , \4299 , \1277 );
not \U$4048 ( \4301 , \4299 );
and \U$4049 ( \4302 , \4301 , \3516 );
nor \U$4050 ( \4303 , \4300 , \4302 );
not \U$4051 ( \4304 , \4303 );
nand \U$4052 ( \4305 , \4294 , \4304 );
not \U$4053 ( \4306 , \4279 );
nand \U$4054 ( \4307 , \4306 , \4291 );
nand \U$4055 ( \4308 , \4305 , \4307 );
not \U$4056 ( \4309 , \4308 );
not \U$4057 ( \4310 , \4309 );
or \U$4058 ( \4311 , \4272 , \4310 );
xor \U$4059 ( \4312 , RIbe28d68_40, RIbe29998_66);
not \U$4060 ( \4313 , \4312 );
xor \U$4061 ( \4314 , RIbe27c88_4, RIbe28d68_40);
nand \U$4062 ( \4315 , \4313 , \4314 );
buf \U$4063 ( \4316 , \4315 );
not \U$4064 ( \4317 , \4316 );
nand \U$4065 ( \4318 , \4317 , RIbe27b98_2);
not \U$4066 ( \4319 , RIbe29998_66);
not \U$4067 ( \4320 , RIbe28d68_40);
or \U$4068 ( \4321 , \4319 , \4320 );
nand \U$4069 ( \4322 , \4321 , RIbe27c88_4);
buf \U$4070 ( \4323 , \4322 );
and \U$4071 ( \4324 , \4318 , \4323 );
not \U$4072 ( \4325 , \4318 );
not \U$4073 ( \4326 , \4006 );
and \U$4074 ( \4327 , \4325 , \4326 );
nor \U$4075 ( \4328 , \4324 , \4327 );
not \U$4076 ( \4329 , RIbe28de0_41);
not \U$4077 ( \4330 , \4021 );
or \U$4078 ( \4331 , \4329 , \4330 );
not \U$4079 ( \4332 , \4025 );
buf \U$4080 ( \4333 , \4332 );
nand \U$4081 ( \4334 , \4333 , RIbe29920_65);
nand \U$4082 ( \4335 , \4331 , \4334 );
and \U$4083 ( \4336 , \4335 , \3471 );
not \U$4084 ( \4337 , \4335 );
and \U$4085 ( \4338 , \4337 , \3448 );
nor \U$4086 ( \4339 , \4336 , \4338 );
xor \U$4087 ( \4340 , \4328 , \4339 );
not \U$4088 ( \4341 , RIbe27c10_3);
not \U$4089 ( \4342 , \3452 );
or \U$4090 ( \4343 , \4341 , \4342 );
nand \U$4091 ( \4344 , \3458 , RIbe28e58_42);
nand \U$4092 ( \4345 , \4343 , \4344 );
buf \U$4093 ( \4346 , \3289 );
and \U$4094 ( \4347 , \4345 , \4346 );
not \U$4095 ( \4348 , \4345 );
and \U$4096 ( \4349 , \4348 , \2887 );
nor \U$4097 ( \4350 , \4347 , \4349 );
and \U$4098 ( \4351 , \4340 , \4350 );
and \U$4099 ( \4352 , \4328 , \4339 );
or \U$4100 ( \4353 , \4351 , \4352 );
nand \U$4101 ( \4354 , \4311 , \4353 );
nand \U$4102 ( \4355 , \4308 , \4270 );
nand \U$4103 ( \4356 , \4354 , \4355 );
and \U$4104 ( \4357 , \4231 , \4356 );
nor \U$4105 ( \4358 , \4156 , \4230 );
nor \U$4106 ( \4359 , \4357 , \4358 );
xor \U$4107 ( \4360 , \3708 , \3695 );
xnor \U$4108 ( \4361 , \4360 , \3683 );
not \U$4109 ( \4362 , \4361 );
not \U$4110 ( \4363 , \3744 );
not \U$4111 ( \4364 , \3733 );
or \U$4112 ( \4365 , \4363 , \4364 );
nand \U$4113 ( \4366 , \3732 , \3743 );
nand \U$4114 ( \4367 , \4365 , \4366 );
and \U$4115 ( \4368 , \4367 , \3724 );
not \U$4116 ( \4369 , \4367 );
and \U$4117 ( \4370 , \4369 , \3746 );
nor \U$4118 ( \4371 , \4368 , \4370 );
not \U$4119 ( \4372 , \4371 );
and \U$4120 ( \4373 , \4362 , \4372 );
xor \U$4121 ( \4374 , \4007 , \4018 );
xor \U$4122 ( \4375 , \4374 , \4033 );
not \U$4123 ( \4376 , \4375 );
and \U$4124 ( \4377 , \3998 , \3985 );
not \U$4125 ( \4378 , \3998 );
and \U$4126 ( \4379 , \4378 , \3986 );
or \U$4127 ( \4380 , \4377 , \4379 );
xor \U$4128 ( \4381 , \4380 , \3976 );
not \U$4129 ( \4382 , \4381 );
or \U$4130 ( \4383 , \4376 , \4382 );
and \U$4131 ( \4384 , \4074 , \4061 );
not \U$4132 ( \4385 , \4074 );
and \U$4133 ( \4386 , \4385 , \4062 );
or \U$4134 ( \4387 , \4384 , \4386 );
xnor \U$4135 ( \4388 , \4387 , \4048 );
nand \U$4136 ( \4389 , \4383 , \4388 );
or \U$4137 ( \4390 , \4375 , \4381 );
nand \U$4138 ( \4391 , \4389 , \4390 );
nand \U$4139 ( \4392 , \4371 , \4361 );
and \U$4140 ( \4393 , \4391 , \4392 );
nor \U$4141 ( \4394 , \4373 , \4393 );
xor \U$4142 ( \4395 , \4359 , \4394 );
not \U$4143 ( \4396 , \3965 );
not \U$4144 ( \4397 , \4396 );
not \U$4145 ( \4398 , \3928 );
or \U$4146 ( \4399 , \4397 , \4398 );
nand \U$4147 ( \4400 , \4399 , \3966 );
not \U$4148 ( \4401 , \4001 );
and \U$4149 ( \4402 , \4036 , \4078 );
not \U$4150 ( \4403 , \4036 );
and \U$4151 ( \4404 , \4403 , \4077 );
or \U$4152 ( \4405 , \4402 , \4404 );
not \U$4153 ( \4406 , \4405 );
or \U$4154 ( \4407 , \4401 , \4406 );
or \U$4155 ( \4408 , \4405 , \4001 );
nand \U$4156 ( \4409 , \4407 , \4408 );
xor \U$4157 ( \4410 , \4400 , \4409 );
xor \U$4158 ( \4411 , \4084 , \4086 );
xor \U$4159 ( \4412 , \4411 , \4095 );
and \U$4160 ( \4413 , \4410 , \4412 );
and \U$4161 ( \4414 , \4400 , \4409 );
or \U$4162 ( \4415 , \4413 , \4414 );
xnor \U$4163 ( \4416 , \4395 , \4415 );
not \U$4164 ( \4417 , \4224 );
not \U$4165 ( \4418 , \4227 );
or \U$4166 ( \4419 , \4417 , \4418 );
or \U$4167 ( \4420 , \4227 , \4224 );
nand \U$4168 ( \4421 , \4419 , \4420 );
and \U$4169 ( \4422 , \4421 , \4228 );
not \U$4170 ( \4423 , \4421 );
and \U$4171 ( \4424 , \4423 , \4157 );
nor \U$4172 ( \4425 , \4422 , \4424 );
and \U$4173 ( \4426 , \4353 , \4308 );
not \U$4174 ( \4427 , \4353 );
and \U$4175 ( \4428 , \4427 , \4309 );
nor \U$4176 ( \4429 , \4426 , \4428 );
and \U$4177 ( \4430 , \4429 , \4270 );
not \U$4178 ( \4431 , \4429 );
and \U$4179 ( \4432 , \4431 , \4271 );
nor \U$4180 ( \4433 , \4430 , \4432 );
and \U$4181 ( \4434 , \4425 , \4433 );
and \U$4182 ( \4435 , \324 , RIbe28660_25);
and \U$4183 ( \4436 , \1371 , RIbe285e8_24);
nor \U$4184 ( \4437 , \4435 , \4436 );
and \U$4185 ( \4438 , \4437 , \1374 );
not \U$4186 ( \4439 , \4437 );
and \U$4187 ( \4440 , \4439 , \1375 );
nor \U$4188 ( \4441 , \4438 , \4440 );
not \U$4189 ( \4442 , \4441 );
nand \U$4190 ( \4443 , RIbe29380_53, RIbe27e68_8);
nor \U$4191 ( \4444 , \4442 , \4443 );
not \U$4192 ( \4445 , RIbe28408_20);
not \U$4193 ( \4446 , \1679 );
or \U$4194 ( \4447 , \4445 , \4446 );
nand \U$4195 ( \4448 , \3897 , RIbe28390_19);
nand \U$4196 ( \4449 , \4447 , \4448 );
not \U$4197 ( \4450 , \4449 );
not \U$4198 ( \4451 , \300 );
and \U$4199 ( \4452 , \4450 , \4451 );
and \U$4200 ( \4453 , \4449 , \300 );
nor \U$4201 ( \4454 , \4452 , \4453 );
and \U$4202 ( \4455 , \1357 , RIbe287c8_28);
and \U$4203 ( \4456 , \264 , RIbe28480_21);
nor \U$4204 ( \4457 , \4455 , \4456 );
and \U$4205 ( \4458 , \4457 , \1362 );
not \U$4206 ( \4459 , \4457 );
and \U$4207 ( \4460 , \4459 , \269 );
nor \U$4208 ( \4461 , \4458 , \4460 );
not \U$4209 ( \4462 , \4461 );
nand \U$4210 ( \4463 , \4454 , \4462 );
not \U$4211 ( \4464 , \4463 );
not \U$4212 ( \4465 , \1232 );
not \U$4213 ( \4466 , RIbe28b10_35);
not \U$4214 ( \4467 , \1223 );
or \U$4215 ( \4468 , \4466 , \4467 );
nand \U$4216 ( \4469 , \429 , RIbe28b88_36);
nand \U$4217 ( \4470 , \4468 , \4469 );
not \U$4218 ( \4471 , \4470 );
or \U$4219 ( \4472 , \4465 , \4471 );
or \U$4220 ( \4473 , \4470 , \3175 );
nand \U$4221 ( \4474 , \4472 , \4473 );
not \U$4222 ( \4475 , \4474 );
or \U$4223 ( \4476 , \4464 , \4475 );
not \U$4224 ( \4477 , \4454 );
nand \U$4225 ( \4478 , \4477 , \4461 );
nand \U$4226 ( \4479 , \4476 , \4478 );
xor \U$4227 ( \4480 , \4444 , \4479 );
not \U$4228 ( \4481 , RIbe29290_51);
not \U$4229 ( \4482 , \3244 );
or \U$4230 ( \4483 , \4481 , \4482 );
nand \U$4231 ( \4484 , \552 , RIbe28a20_33);
nand \U$4232 ( \4485 , \4483 , \4484 );
and \U$4233 ( \4486 , \4485 , \1245 );
not \U$4234 ( \4487 , \4485 );
and \U$4235 ( \4488 , \4487 , \1333 );
nor \U$4236 ( \4489 , \4486 , \4488 );
and \U$4237 ( \4490 , \1161 , RIbe29560_57);
and \U$4238 ( \4491 , \2000 , RIbe28228_16);
nor \U$4239 ( \4492 , \4490 , \4491 );
and \U$4240 ( \4493 , \4492 , \752 );
not \U$4241 ( \4494 , \4492 );
and \U$4242 ( \4495 , \4494 , \1011 );
nor \U$4243 ( \4496 , \4493 , \4495 );
xor \U$4244 ( \4497 , \4489 , \4496 );
and \U$4245 ( \4498 , \666 , RIbe289a8_32);
and \U$4246 ( \4499 , \1180 , RIbe28930_31);
nor \U$4247 ( \4500 , \4498 , \4499 );
and \U$4248 ( \4501 , \4500 , \564 );
not \U$4249 ( \4502 , \4500 );
and \U$4250 ( \4503 , \4502 , \672 );
nor \U$4251 ( \4504 , \4501 , \4503 );
and \U$4252 ( \4505 , \4497 , \4504 );
and \U$4253 ( \4506 , \4489 , \4496 );
or \U$4254 ( \4507 , \4505 , \4506 );
and \U$4255 ( \4508 , \4480 , \4507 );
and \U$4256 ( \4509 , \4444 , \4479 );
or \U$4257 ( \4510 , \4508 , \4509 );
not \U$4258 ( \4511 , \1153 );
not \U$4259 ( \4512 , RIbe281b0_15);
not \U$4260 ( \4513 , \1143 );
or \U$4261 ( \4514 , \4512 , \4513 );
nand \U$4262 ( \4515 , \1147 , RIbe280c0_13);
nand \U$4263 ( \4516 , \4514 , \4515 );
not \U$4264 ( \4517 , \4516 );
or \U$4265 ( \4518 , \4511 , \4517 );
or \U$4266 ( \4519 , \4516 , \1157 );
nand \U$4267 ( \4520 , \4518 , \4519 );
not \U$4268 ( \4521 , \4520 );
not \U$4269 ( \4522 , RIbe29830_63);
not \U$4270 ( \4523 , \1633 );
or \U$4271 ( \4524 , \4522 , \4523 );
nand \U$4272 ( \4525 , \2817 , RIbe296c8_60);
nand \U$4273 ( \4526 , \4524 , \4525 );
and \U$4274 ( \4527 , \4526 , \1309 );
not \U$4275 ( \4528 , \4526 );
and \U$4276 ( \4529 , \4528 , \1082 );
nor \U$4277 ( \4530 , \4527 , \4529 );
not \U$4278 ( \4531 , \4530 );
or \U$4279 ( \4532 , \4521 , \4531 );
or \U$4280 ( \4533 , \4530 , \4520 );
and \U$4281 ( \4534 , \1286 , RIbe29650_59);
and \U$4282 ( \4535 , \1117 , RIbe29038_46);
nor \U$4283 ( \4536 , \4534 , \4535 );
and \U$4284 ( \4537 , \4536 , \1132 );
not \U$4285 ( \4538 , \4536 );
and \U$4286 ( \4539 , \4538 , \2563 );
nor \U$4287 ( \4540 , \4537 , \4539 );
not \U$4288 ( \4541 , \4540 );
nand \U$4289 ( \4542 , \4533 , \4541 );
nand \U$4290 ( \4543 , \4532 , \4542 );
and \U$4291 ( \4544 , \1272 , RIbe28fc0_45);
not \U$4292 ( \4545 , RIbe290b0_47);
nor \U$4293 ( \4546 , \2889 , \4545 );
nor \U$4294 ( \4547 , \4544 , \4546 );
and \U$4295 ( \4548 , \4547 , \1076 );
not \U$4296 ( \4549 , \4547 );
and \U$4297 ( \4550 , \4549 , \1277 );
nor \U$4298 ( \4551 , \4548 , \4550 );
not \U$4299 ( \4552 , RIbe29a88_68);
not \U$4300 ( \4553 , \3476 );
or \U$4301 ( \4554 , \4552 , \4553 );
nand \U$4302 ( \4555 , \3267 , RIbe27d78_6);
nand \U$4303 ( \4556 , \4554 , \4555 );
and \U$4304 ( \4557 , \4556 , \3272 );
not \U$4305 ( \4558 , \4556 );
and \U$4306 ( \4559 , \4558 , \2576 );
nor \U$4307 ( \4560 , \4557 , \4559 );
xor \U$4308 ( \4561 , \4551 , \4560 );
and \U$4309 ( \4562 , \3285 , RIbe27d00_5);
and \U$4310 ( \4563 , \3458 , RIbe27c10_3);
nor \U$4311 ( \4564 , \4562 , \4563 );
and \U$4312 ( \4565 , \4564 , \2887 );
not \U$4313 ( \4566 , \4564 );
and \U$4314 ( \4567 , \4566 , \4346 );
nor \U$4315 ( \4568 , \4565 , \4567 );
and \U$4316 ( \4569 , \4561 , \4568 );
and \U$4317 ( \4570 , \4551 , \4560 );
or \U$4318 ( \4571 , \4569 , \4570 );
xor \U$4319 ( \4572 , \4543 , \4571 );
not \U$4320 ( \4573 , RIbe28e58_42);
not \U$4321 ( \4574 , \4021 );
or \U$4322 ( \4575 , \4573 , \4574 );
nand \U$4323 ( \4576 , \4027 , RIbe28de0_41);
nand \U$4324 ( \4577 , \4575 , \4576 );
and \U$4325 ( \4578 , \4577 , \3471 );
not \U$4326 ( \4579 , \4577 );
and \U$4327 ( \4580 , \4579 , \3448 );
nor \U$4328 ( \4581 , \4578 , \4580 );
not \U$4329 ( \4582 , \4581 );
and \U$4330 ( \4583 , RIbe298a8_64, RIbe28cf0_39);
not \U$4331 ( \4584 , RIbe29998_66);
nor \U$4332 ( \4585 , \4583 , \4584 );
buf \U$4333 ( \4586 , \4585 );
or \U$4334 ( \4587 , \4582 , \4586 );
not \U$4335 ( \4588 , RIbe28cf0_39);
not \U$4336 ( \4589 , RIbe298a8_64);
or \U$4337 ( \4590 , \4588 , \4589 );
nand \U$4338 ( \4591 , \4590 , RIbe29998_66);
buf \U$4339 ( \4592 , \4591 );
or \U$4340 ( \4593 , \4581 , \4592 );
not \U$4341 ( \4594 , RIbe29920_65);
not \U$4342 ( \4595 , \4316 );
not \U$4343 ( \4596 , \4595 );
or \U$4344 ( \4597 , \4594 , \4596 );
not \U$4345 ( \4598 , \4312 );
not \U$4346 ( \4599 , \4598 );
buf \U$4347 ( \4600 , \4599 );
nand \U$4348 ( \4601 , \4600 , RIbe27b98_2);
nand \U$4349 ( \4602 , \4597 , \4601 );
buf \U$4350 ( \4603 , \4005 );
and \U$4351 ( \4604 , \4602 , \4603 );
not \U$4352 ( \4605 , \4602 );
and \U$4353 ( \4606 , \4605 , \4323 );
nor \U$4354 ( \4607 , \4604 , \4606 );
nand \U$4355 ( \4608 , \4593 , \4607 );
nand \U$4356 ( \4609 , \4587 , \4608 );
and \U$4357 ( \4610 , \4572 , \4609 );
and \U$4358 ( \4611 , \4543 , \4571 );
or \U$4359 ( \4612 , \4610 , \4611 );
xor \U$4360 ( \4613 , \4510 , \4612 );
not \U$4361 ( \4614 , \4165 );
not \U$4362 ( \4615 , \4184 );
or \U$4363 ( \4616 , \4614 , \4615 );
or \U$4364 ( \4617 , \4184 , \4165 );
nand \U$4365 ( \4618 , \4616 , \4617 );
xnor \U$4366 ( \4619 , \4176 , \4618 );
xor \U$4367 ( \4620 , \4157 , \4619 );
not \U$4368 ( \4621 , \4198 );
not \U$4369 ( \4622 , \4221 );
or \U$4370 ( \4623 , \4621 , \4622 );
or \U$4371 ( \4624 , \4221 , \4198 );
nand \U$4372 ( \4625 , \4623 , \4624 );
xnor \U$4373 ( \4626 , \4625 , \4209 );
and \U$4374 ( \4627 , \4620 , \4626 );
and \U$4375 ( \4628 , \4157 , \4619 );
or \U$4376 ( \4629 , \4627 , \4628 );
and \U$4377 ( \4630 , \4613 , \4629 );
and \U$4378 ( \4631 , \4510 , \4612 );
or \U$4379 ( \4632 , \4630 , \4631 );
xor \U$4380 ( \4633 , \4434 , \4632 );
xor \U$4381 ( \4634 , \4328 , \4339 );
xor \U$4382 ( \4635 , \4634 , \4350 );
not \U$4383 ( \4636 , \4304 );
not \U$4384 ( \4637 , \4292 );
or \U$4385 ( \4638 , \4636 , \4637 );
nand \U$4386 ( \4639 , \4291 , \4303 );
nand \U$4387 ( \4640 , \4638 , \4639 );
and \U$4388 ( \4641 , \4640 , \4306 );
not \U$4389 ( \4642 , \4640 );
and \U$4390 ( \4643 , \4642 , \4279 );
nor \U$4391 ( \4644 , \4641 , \4643 );
xor \U$4392 ( \4645 , \4635 , \4644 );
and \U$4393 ( \4646 , \4265 , \4253 );
not \U$4394 ( \4647 , \4265 );
and \U$4395 ( \4648 , \4647 , \4267 );
or \U$4396 ( \4649 , \4646 , \4648 );
and \U$4397 ( \4650 , \4649 , \4268 );
not \U$4398 ( \4651 , \4649 );
and \U$4399 ( \4652 , \4651 , \4241 );
nor \U$4400 ( \4653 , \4650 , \4652 );
and \U$4401 ( \4654 , \4645 , \4653 );
and \U$4402 ( \4655 , \4635 , \4644 );
or \U$4403 ( \4656 , \4654 , \4655 );
not \U$4404 ( \4657 , \4153 );
xor \U$4405 ( \4658 , \4149 , \4147 );
not \U$4406 ( \4659 , \4658 );
or \U$4407 ( \4660 , \4657 , \4659 );
or \U$4408 ( \4661 , \4658 , \4153 );
nand \U$4409 ( \4662 , \4660 , \4661 );
xor \U$4410 ( \4663 , \4656 , \4662 );
not \U$4411 ( \4664 , \4381 );
not \U$4412 ( \4665 , \4388 );
not \U$4413 ( \4666 , \4375 );
or \U$4414 ( \4667 , \4665 , \4666 );
or \U$4415 ( \4668 , \4375 , \4388 );
nand \U$4416 ( \4669 , \4667 , \4668 );
not \U$4417 ( \4670 , \4669 );
or \U$4418 ( \4671 , \4664 , \4670 );
or \U$4419 ( \4672 , \4669 , \4381 );
nand \U$4420 ( \4673 , \4671 , \4672 );
and \U$4421 ( \4674 , \4663 , \4673 );
and \U$4422 ( \4675 , \4656 , \4662 );
or \U$4423 ( \4676 , \4674 , \4675 );
and \U$4424 ( \4677 , \4633 , \4676 );
and \U$4425 ( \4678 , \4434 , \4632 );
or \U$4426 ( \4679 , \4677 , \4678 );
xor \U$4427 ( \4680 , \4361 , \4371 );
xor \U$4428 ( \4681 , \4680 , \4391 );
not \U$4429 ( \4682 , \4156 );
not \U$4430 ( \4683 , \4356 );
not \U$4431 ( \4684 , \4230 );
or \U$4432 ( \4685 , \4683 , \4684 );
or \U$4433 ( \4686 , \4230 , \4356 );
nand \U$4434 ( \4687 , \4685 , \4686 );
not \U$4435 ( \4688 , \4687 );
or \U$4436 ( \4689 , \4682 , \4688 );
or \U$4437 ( \4690 , \4156 , \4687 );
nand \U$4438 ( \4691 , \4689 , \4690 );
xor \U$4439 ( \4692 , \4681 , \4691 );
xor \U$4440 ( \4693 , \4400 , \4409 );
xor \U$4441 ( \4694 , \4693 , \4412 );
and \U$4442 ( \4695 , \4692 , \4694 );
and \U$4443 ( \4696 , \4681 , \4691 );
or \U$4444 ( \4697 , \4695 , \4696 );
xor \U$4445 ( \4698 , \4679 , \4697 );
not \U$4446 ( \4699 , \3674 );
not \U$4447 ( \4700 , \3711 );
not \U$4448 ( \4701 , \3748 );
or \U$4449 ( \4702 , \4700 , \4701 );
or \U$4450 ( \4703 , \3748 , \3711 );
nand \U$4451 ( \4704 , \4702 , \4703 );
not \U$4452 ( \4705 , \4704 );
or \U$4453 ( \4706 , \4699 , \4705 );
or \U$4454 ( \4707 , \4704 , \3674 );
nand \U$4455 ( \4708 , \4706 , \4707 );
xor \U$4456 ( \4709 , \3966 , \4081 );
xor \U$4457 ( \4710 , \4709 , \4097 );
xor \U$4458 ( \4711 , \4708 , \4710 );
not \U$4459 ( \4712 , \3881 );
not \U$4460 ( \4713 , \3878 );
and \U$4461 ( \4714 , \4712 , \4713 );
and \U$4462 ( \4715 , \3881 , \3878 );
nor \U$4463 ( \4716 , \4714 , \4715 );
xnor \U$4464 ( \4717 , \4716 , \3884 );
xor \U$4465 ( \4718 , \4711 , \4717 );
xnor \U$4466 ( \4719 , \4698 , \4718 );
nand \U$4467 ( \4720 , \4416 , \4719 );
not \U$4468 ( \4721 , \4720 );
xor \U$4469 ( \4722 , \4444 , \4479 );
xor \U$4470 ( \4723 , \4722 , \4507 );
xor \U$4471 ( \4724 , \4543 , \4571 );
xor \U$4472 ( \4725 , \4724 , \4609 );
and \U$4473 ( \4726 , \4723 , \4725 );
not \U$4474 ( \4727 , RIbe280c0_13);
not \U$4475 ( \4728 , \1298 );
or \U$4476 ( \4729 , \4727 , \4728 );
buf \U$4477 ( \4730 , \1098 );
nand \U$4478 ( \4731 , \4730 , RIbe29830_63);
nand \U$4479 ( \4732 , \4729 , \4731 );
and \U$4480 ( \4733 , \4732 , \4251 );
not \U$4481 ( \4734 , \4732 );
and \U$4482 ( \4735 , \4734 , \1309 );
nor \U$4483 ( \4736 , \4733 , \4735 );
not \U$4484 ( \4737 , RIbe28228_16);
not \U$4485 ( \4738 , \4257 );
or \U$4486 ( \4739 , \4737 , \4738 );
nand \U$4487 ( \4740 , \1147 , RIbe281b0_15);
nand \U$4488 ( \4741 , \4739 , \4740 );
not \U$4489 ( \4742 , \1652 );
and \U$4490 ( \4743 , \4741 , \4742 );
not \U$4491 ( \4744 , \4741 );
and \U$4492 ( \4745 , \4744 , \1794 );
nor \U$4493 ( \4746 , \4743 , \4745 );
nand \U$4494 ( \4747 , \4736 , \4746 );
not \U$4495 ( \4748 , \1112 );
not \U$4496 ( \4749 , \4748 );
and \U$4497 ( \4750 , \4749 , RIbe296c8_60);
and \U$4498 ( \4751 , \1117 , RIbe29650_59);
nor \U$4499 ( \4752 , \4750 , \4751 );
and \U$4500 ( \4753 , \4752 , \1132 );
not \U$4501 ( \4754 , \4752 );
and \U$4502 ( \4755 , \4754 , \3491 );
nor \U$4503 ( \4756 , \4753 , \4755 );
not \U$4504 ( \4757 , \4756 );
and \U$4505 ( \4758 , \4747 , \4757 );
nor \U$4506 ( \4759 , \4736 , \4746 );
nor \U$4507 ( \4760 , \4758 , \4759 );
not \U$4508 ( \4761 , \4760 );
not \U$4509 ( \4762 , \4761 );
not \U$4510 ( \4763 , RIbe27d78_6);
not \U$4511 ( \4764 , \3283 );
not \U$4512 ( \4765 , \4764 );
or \U$4513 ( \4766 , \4763 , \4765 );
nand \U$4514 ( \4767 , \4011 , RIbe27d00_5);
nand \U$4515 ( \4768 , \4766 , \4767 );
not \U$4516 ( \4769 , \4768 );
not \U$4517 ( \4770 , \3461 );
and \U$4518 ( \4771 , \4769 , \4770 );
and \U$4519 ( \4772 , \4768 , \2887 );
nor \U$4520 ( \4773 , \4771 , \4772 );
not \U$4521 ( \4774 , \4773 );
not \U$4522 ( \4775 , \4774 );
not \U$4523 ( \4776 , RIbe290b0_47);
not \U$4524 ( \4777 , \2898 );
or \U$4525 ( \4778 , \4776 , \4777 );
nand \U$4526 ( \4779 , \4284 , RIbe29a88_68);
nand \U$4527 ( \4780 , \4778 , \4779 );
and \U$4528 ( \4781 , \4780 , \3272 );
not \U$4529 ( \4782 , \4780 );
not \U$4530 ( \4783 , \2380 );
and \U$4531 ( \4784 , \4782 , \4783 );
nor \U$4532 ( \4785 , \4781 , \4784 );
not \U$4533 ( \4786 , \4785 );
or \U$4534 ( \4787 , \4775 , \4786 );
or \U$4535 ( \4788 , \4785 , \4774 );
not \U$4536 ( \4789 , \2889 );
not \U$4537 ( \4790 , \1931 );
and \U$4538 ( \4791 , \4789 , \4790 );
and \U$4539 ( \4792 , \2390 , RIbe29038_46);
nor \U$4540 ( \4793 , \4791 , \4792 );
and \U$4541 ( \4794 , \4793 , \1277 );
not \U$4542 ( \4795 , \4793 );
and \U$4543 ( \4796 , \4795 , \1076 );
or \U$4544 ( \4797 , \4794 , \4796 );
nand \U$4545 ( \4798 , \4788 , \4797 );
nand \U$4546 ( \4799 , \4787 , \4798 );
not \U$4547 ( \4800 , \4799 );
or \U$4548 ( \4801 , \4762 , \4800 );
or \U$4549 ( \4802 , \4799 , \4761 );
not \U$4550 ( \4803 , RIbe28de0_41);
not \U$4551 ( \4804 , \4316 );
not \U$4552 ( \4805 , \4804 );
or \U$4553 ( \4806 , \4803 , \4805 );
buf \U$4554 ( \4807 , \4598 );
not \U$4555 ( \4808 , \4807 );
buf \U$4556 ( \4809 , \4808 );
nand \U$4557 ( \4810 , \4809 , RIbe29920_65);
nand \U$4558 ( \4811 , \4806 , \4810 );
and \U$4559 ( \4812 , \4811 , \4323 );
not \U$4560 ( \4813 , \4811 );
and \U$4561 ( \4814 , \4813 , \4326 );
nor \U$4562 ( \4815 , \4812 , \4814 );
not \U$4563 ( \4816 , RIbe27c10_3);
not \U$4564 ( \4817 , \4021 );
or \U$4565 ( \4818 , \4816 , \4817 );
nand \U$4566 ( \4819 , \4333 , RIbe28e58_42);
nand \U$4567 ( \4820 , \4818 , \4819 );
not \U$4568 ( \4821 , \3697 );
xor \U$4569 ( \4822 , \4820 , \4821 );
and \U$4570 ( \4823 , \4815 , \4822 );
xor \U$4571 ( \4824 , RIbe298a8_64, RIbe28cf0_39);
not \U$4572 ( \4825 , \4824 );
xor \U$4573 ( \4826 , RIbe298a8_64, RIbe29998_66);
nand \U$4574 ( \4827 , \4825 , \4826 );
buf \U$4575 ( \4828 , \4827 );
not \U$4576 ( \4829 , \4828 );
buf \U$4577 ( \4830 , \4829 );
not \U$4578 ( \4831 , \4830 );
not \U$4579 ( \4832 , \4831 );
nand \U$4580 ( \4833 , \4832 , RIbe27b98_2);
and \U$4581 ( \4834 , \4833 , \4586 );
not \U$4582 ( \4835 , \4833 );
and \U$4583 ( \4836 , \4835 , \4592 );
nor \U$4584 ( \4837 , \4834 , \4836 );
nor \U$4585 ( \4838 , \4823 , \4837 );
nor \U$4586 ( \4839 , \4815 , \4822 );
nor \U$4587 ( \4840 , \4838 , \4839 );
not \U$4588 ( \4841 , \4840 );
nand \U$4589 ( \4842 , \4802 , \4841 );
nand \U$4590 ( \4843 , \4801 , \4842 );
not \U$4591 ( \4844 , RIbe27e68_8);
not \U$4592 ( \4845 , \3160 );
or \U$4593 ( \4846 , \4844 , \4845 );
nand \U$4594 ( \4847 , \329 , RIbe28660_25);
nand \U$4595 ( \4848 , \4846 , \4847 );
not \U$4596 ( \4849 , \4848 );
not \U$4597 ( \4850 , \1374 );
and \U$4598 ( \4851 , \4849 , \4850 );
and \U$4599 ( \4852 , \4848 , \339 );
nor \U$4600 ( \4853 , \4851 , \4852 );
nand \U$4601 ( \4854 , RIbe29380_53, RIbe27f58_10);
nand \U$4602 ( \4855 , \4853 , \4854 );
not \U$4603 ( \4856 , RIbe28930_31);
not \U$4604 ( \4857 , \1002 );
not \U$4605 ( \4858 , \4857 );
not \U$4606 ( \4859 , \4858 );
or \U$4607 ( \4860 , \4856 , \4859 );
nand \U$4608 ( \4861 , \1203 , RIbe29560_57);
nand \U$4609 ( \4862 , \4860 , \4861 );
or \U$4610 ( \4863 , \4862 , \750 );
nand \U$4611 ( \4864 , \4862 , \1813 );
nand \U$4612 ( \4865 , \4863 , \4864 );
not \U$4613 ( \4866 , RIbe28b88_36);
not \U$4614 ( \4867 , \548 );
or \U$4615 ( \4868 , \4866 , \4867 );
nand \U$4616 ( \4869 , \1327 , RIbe29290_51);
nand \U$4617 ( \4870 , \4868 , \4869 );
and \U$4618 ( \4871 , \4870 , \1330 );
not \U$4619 ( \4872 , \4870 );
and \U$4620 ( \4873 , \4872 , \1333 );
nor \U$4621 ( \4874 , \4871 , \4873 );
or \U$4622 ( \4875 , \4865 , \4874 );
not \U$4623 ( \4876 , \1611 );
not \U$4624 ( \4877 , \3421 );
and \U$4625 ( \4878 , \4876 , \4877 );
and \U$4626 ( \4879 , \1744 , RIbe28a20_33);
nor \U$4627 ( \4880 , \4878 , \4879 );
and \U$4628 ( \4881 , \4880 , \564 );
not \U$4629 ( \4882 , \4880 );
and \U$4630 ( \4883 , \4882 , \3959 );
nor \U$4631 ( \4884 , \4881 , \4883 );
nand \U$4632 ( \4885 , \4875 , \4884 );
nand \U$4633 ( \4886 , \4865 , \4874 );
nand \U$4634 ( \4887 , \4885 , \4886 );
xor \U$4635 ( \4888 , \4855 , \4887 );
and \U$4636 ( \4889 , \1528 , RIbe28480_21);
and \U$4637 ( \4890 , \1531 , RIbe28408_20);
nor \U$4638 ( \4891 , \4889 , \4890 );
and \U$4639 ( \4892 , \4891 , \300 );
not \U$4640 ( \4893 , \4891 );
and \U$4641 ( \4894 , \4893 , \293 );
nor \U$4642 ( \4895 , \4892 , \4894 );
not \U$4643 ( \4896 , \4895 );
not \U$4644 ( \4897 , \4896 );
and \U$4645 ( \4898 , \1357 , RIbe285e8_24);
and \U$4646 ( \4899 , \264 , RIbe287c8_28);
nor \U$4647 ( \4900 , \4898 , \4899 );
and \U$4648 ( \4901 , \4900 , \268 );
not \U$4649 ( \4902 , \4900 );
and \U$4650 ( \4903 , \4902 , \1362 );
nor \U$4651 ( \4904 , \4901 , \4903 );
not \U$4652 ( \4905 , \4904 );
or \U$4653 ( \4906 , \4897 , \4905 );
not \U$4654 ( \4907 , RIbe28390_19);
not \U$4655 ( \4908 , \383 );
or \U$4656 ( \4909 , \4907 , \4908 );
nand \U$4657 ( \4910 , \429 , RIbe28b10_35);
nand \U$4658 ( \4911 , \4909 , \4910 );
and \U$4659 ( \4912 , \4911 , \313 );
not \U$4660 ( \4913 , \4911 );
and \U$4661 ( \4914 , \4913 , \306 );
nor \U$4662 ( \4915 , \4912 , \4914 );
not \U$4663 ( \4916 , \4915 );
nand \U$4664 ( \4917 , \4906 , \4916 );
not \U$4665 ( \4918 , \4904 );
nand \U$4666 ( \4919 , \4895 , \4918 );
nand \U$4667 ( \4920 , \4917 , \4919 );
and \U$4668 ( \4921 , \4888 , \4920 );
and \U$4669 ( \4922 , \4855 , \4887 );
or \U$4670 ( \4923 , \4921 , \4922 );
xor \U$4671 ( \4924 , \4843 , \4923 );
not \U$4672 ( \4925 , \4443 );
not \U$4673 ( \4926 , \4441 );
or \U$4674 ( \4927 , \4925 , \4926 );
or \U$4675 ( \4928 , \4441 , \4443 );
nand \U$4676 ( \4929 , \4927 , \4928 );
xor \U$4677 ( \4930 , \4462 , \4454 );
xor \U$4678 ( \4931 , \4930 , \4474 );
xor \U$4679 ( \4932 , \4929 , \4931 );
xor \U$4680 ( \4933 , \4489 , \4496 );
xor \U$4681 ( \4934 , \4933 , \4504 );
and \U$4682 ( \4935 , \4932 , \4934 );
and \U$4683 ( \4936 , \4929 , \4931 );
or \U$4684 ( \4937 , \4935 , \4936 );
and \U$4685 ( \4938 , \4924 , \4937 );
and \U$4686 ( \4939 , \4843 , \4923 );
or \U$4687 ( \4940 , \4938 , \4939 );
xor \U$4688 ( \4941 , \4726 , \4940 );
xor \U$4689 ( \4942 , \4551 , \4560 );
xor \U$4690 ( \4943 , \4942 , \4568 );
not \U$4691 ( \4944 , \4943 );
not \U$4692 ( \4945 , \4591 );
not \U$4693 ( \4946 , \4945 );
xor \U$4694 ( \4947 , \4323 , \4946 );
xnor \U$4695 ( \4948 , \4947 , \4602 );
and \U$4696 ( \4949 , \4948 , \4582 );
not \U$4697 ( \4950 , \4948 );
and \U$4698 ( \4951 , \4950 , \4581 );
nor \U$4699 ( \4952 , \4949 , \4951 );
not \U$4700 ( \4953 , \4952 );
not \U$4701 ( \4954 , \4953 );
or \U$4702 ( \4955 , \4944 , \4954 );
or \U$4703 ( \4956 , \4953 , \4943 );
and \U$4704 ( \4957 , \4530 , \4540 );
not \U$4705 ( \4958 , \4530 );
and \U$4706 ( \4959 , \4958 , \4541 );
or \U$4707 ( \4960 , \4957 , \4959 );
xor \U$4708 ( \4961 , \4960 , \4520 );
nand \U$4709 ( \4962 , \4956 , \4961 );
nand \U$4710 ( \4963 , \4955 , \4962 );
xor \U$4711 ( \4964 , \4635 , \4644 );
xor \U$4712 ( \4965 , \4964 , \4653 );
xor \U$4713 ( \4966 , \4963 , \4965 );
xor \U$4714 ( \4967 , \4157 , \4619 );
xor \U$4715 ( \4968 , \4967 , \4626 );
and \U$4716 ( \4969 , \4966 , \4968 );
and \U$4717 ( \4970 , \4963 , \4965 );
or \U$4718 ( \4971 , \4969 , \4970 );
and \U$4719 ( \4972 , \4941 , \4971 );
and \U$4720 ( \4973 , \4726 , \4940 );
or \U$4721 ( \4974 , \4972 , \4973 );
xor \U$4722 ( \4975 , \4425 , \4433 );
xor \U$4723 ( \4976 , \4510 , \4612 );
xor \U$4724 ( \4977 , \4976 , \4629 );
xor \U$4725 ( \4978 , \4975 , \4977 );
xor \U$4726 ( \4979 , \4656 , \4662 );
xor \U$4727 ( \4980 , \4979 , \4673 );
and \U$4728 ( \4981 , \4978 , \4980 );
and \U$4729 ( \4982 , \4975 , \4977 );
or \U$4730 ( \4983 , \4981 , \4982 );
xor \U$4731 ( \4984 , \4974 , \4983 );
xor \U$4732 ( \4985 , \4681 , \4691 );
xor \U$4733 ( \4986 , \4985 , \4694 );
and \U$4734 ( \4987 , \4984 , \4986 );
and \U$4735 ( \4988 , \4974 , \4983 );
or \U$4736 ( \4989 , \4987 , \4988 );
not \U$4737 ( \4990 , \4989 );
or \U$4738 ( \4991 , \4721 , \4990 );
not \U$4739 ( \4992 , \4416 );
not \U$4740 ( \4993 , \4719 );
nand \U$4741 ( \4994 , \4992 , \4993 );
nand \U$4742 ( \4995 , \4991 , \4994 );
xor \U$4743 ( \4996 , \3750 , \3817 );
xor \U$4744 ( \4997 , \4996 , \3835 );
not \U$4745 ( \4998 , \4997 );
xor \U$4746 ( \4999 , \3890 , \4100 );
xnor \U$4747 ( \5000 , \4999 , \3888 );
not \U$4748 ( \5001 , \5000 );
or \U$4749 ( \5002 , \4998 , \5001 );
or \U$4750 ( \5003 , \5000 , \4997 );
nand \U$4751 ( \5004 , \5002 , \5003 );
xor \U$4752 ( \5005 , \3847 , \3849 );
xor \U$4753 ( \5006 , \5005 , \3852 );
xor \U$4754 ( \5007 , \4708 , \4710 );
and \U$4755 ( \5008 , \5007 , \4717 );
and \U$4756 ( \5009 , \4708 , \4710 );
or \U$4757 ( \5010 , \5008 , \5009 );
xor \U$4758 ( \5011 , \5006 , \5010 );
or \U$4759 ( \5012 , \4359 , \4394 );
not \U$4760 ( \5013 , \4394 );
not \U$4761 ( \5014 , \4359 );
or \U$4762 ( \5015 , \5013 , \5014 );
nand \U$4763 ( \5016 , \5015 , \4415 );
nand \U$4764 ( \5017 , \5012 , \5016 );
xor \U$4765 ( \5018 , \5011 , \5017 );
xor \U$4766 ( \5019 , \5004 , \5018 );
not \U$4767 ( \5020 , \4718 );
not \U$4768 ( \5021 , \4679 );
or \U$4769 ( \5022 , \5020 , \5021 );
or \U$4770 ( \5023 , \4718 , \4679 );
nand \U$4771 ( \5024 , \5023 , \4697 );
nand \U$4772 ( \5025 , \5022 , \5024 );
xor \U$4773 ( \5026 , \5019 , \5025 );
xor \U$4774 ( \5027 , \4995 , \5026 );
not \U$4775 ( \5028 , \5027 );
not \U$4776 ( \5029 , \5028 );
xor \U$4777 ( \5030 , \4416 , \4989 );
xor \U$4778 ( \5031 , \5030 , \4993 );
not \U$4779 ( \5032 , \5031 );
xor \U$4780 ( \5033 , \4434 , \4632 );
xor \U$4781 ( \5034 , \5033 , \4676 );
xor \U$4782 ( \5035 , \4855 , \4887 );
xor \U$4783 ( \5036 , \5035 , \4920 );
and \U$4784 ( \5037 , \4840 , \4760 );
not \U$4785 ( \5038 , \4840 );
and \U$4786 ( \5039 , \5038 , \4761 );
nor \U$4787 ( \5040 , \5037 , \5039 );
xor \U$4788 ( \5041 , \5040 , \4799 );
and \U$4789 ( \5042 , \5036 , \5041 );
nand \U$4790 ( \5043 , RIbe27b20_1, RIbe29b78_70);
nand \U$4791 ( \5044 , \5043 , RIbe28cf0_39);
not \U$4792 ( \5045 , \5044 );
not \U$4793 ( \5046 , \5045 );
not \U$4794 ( \5047 , \5046 );
not \U$4795 ( \5048 , RIbe29920_65);
not \U$4796 ( \5049 , \4830 );
or \U$4797 ( \5050 , \5048 , \5049 );
not \U$4798 ( \5051 , \4824 );
not \U$4799 ( \5052 , \5051 );
nand \U$4800 ( \5053 , \5052 , RIbe27b98_2);
nand \U$4801 ( \5054 , \5050 , \5053 );
xnor \U$4802 ( \5055 , \5054 , \4586 );
xor \U$4803 ( \5056 , \5047 , \5055 );
not \U$4804 ( \5057 , RIbe28e58_42);
not \U$4805 ( \5058 , \4316 );
not \U$4806 ( \5059 , \5058 );
or \U$4807 ( \5060 , \5057 , \5059 );
nand \U$4808 ( \5061 , \4600 , RIbe28de0_41);
nand \U$4809 ( \5062 , \5060 , \5061 );
and \U$4810 ( \5063 , \5062 , \4603 );
not \U$4811 ( \5064 , \5062 );
and \U$4812 ( \5065 , \5064 , \4323 );
or \U$4813 ( \5066 , \5063 , \5065 );
and \U$4814 ( \5067 , \5056 , \5066 );
and \U$4815 ( \5068 , \5047 , \5055 );
or \U$4816 ( \5069 , \5067 , \5068 );
not \U$4817 ( \5070 , \5069 );
not \U$4818 ( \5071 , \2887 );
not \U$4819 ( \5072 , RIbe29a88_68);
not \U$4820 ( \5073 , \3685 );
or \U$4821 ( \5074 , \5072 , \5073 );
nand \U$4822 ( \5075 , \4011 , RIbe27d78_6);
nand \U$4823 ( \5076 , \5074 , \5075 );
not \U$4824 ( \5077 , \5076 );
or \U$4825 ( \5078 , \5071 , \5077 );
or \U$4826 ( \5079 , \5076 , \3461 );
nand \U$4827 ( \5080 , \5078 , \5079 );
not \U$4828 ( \5081 , \5080 );
not \U$4829 ( \5082 , RIbe28fc0_45);
not \U$4830 ( \5083 , \4051 );
or \U$4831 ( \5084 , \5082 , \5083 );
nand \U$4832 ( \5085 , \3267 , RIbe290b0_47);
nand \U$4833 ( \5086 , \5084 , \5085 );
not \U$4834 ( \5087 , \5086 );
not \U$4835 ( \5088 , \3275 );
and \U$4836 ( \5089 , \5087 , \5088 );
and \U$4837 ( \5090 , \5086 , \2576 );
nor \U$4838 ( \5091 , \5089 , \5090 );
nand \U$4839 ( \5092 , \5081 , \5091 );
not \U$4840 ( \5093 , RIbe27d00_5);
not \U$4841 ( \5094 , \3703 );
not \U$4842 ( \5095 , \5094 );
or \U$4843 ( \5096 , \5093 , \5095 );
nand \U$4844 ( \5097 , \4333 , RIbe27c10_3);
nand \U$4845 ( \5098 , \5096 , \5097 );
and \U$4846 ( \5099 , \5098 , \4821 );
not \U$4847 ( \5100 , \5098 );
and \U$4848 ( \5101 , \5100 , \3471 );
nor \U$4849 ( \5102 , \5099 , \5101 );
not \U$4850 ( \5103 , \5102 );
and \U$4851 ( \5104 , \5092 , \5103 );
nor \U$4852 ( \5105 , \5081 , \5091 );
nor \U$4853 ( \5106 , \5104 , \5105 );
not \U$4854 ( \5107 , \5106 );
or \U$4855 ( \5108 , \5070 , \5107 );
and \U$4856 ( \5109 , \4749 , RIbe29830_63);
and \U$4857 ( \5110 , \1117 , RIbe296c8_60);
nor \U$4858 ( \5111 , \5109 , \5110 );
and \U$4859 ( \5112 , \5111 , \1448 );
not \U$4860 ( \5113 , \5111 );
and \U$4861 ( \5114 , \5113 , \1132 );
nor \U$4862 ( \5115 , \5112 , \5114 );
not \U$4863 ( \5116 , \5115 );
not \U$4864 ( \5117 , RIbe281b0_15);
not \U$4865 ( \5118 , \1094 );
or \U$4866 ( \5119 , \5117 , \5118 );
nand \U$4867 ( \5120 , \1455 , RIbe280c0_13);
nand \U$4868 ( \5121 , \5119 , \5120 );
not \U$4869 ( \5122 , \5121 );
not \U$4870 ( \5123 , \4251 );
and \U$4871 ( \5124 , \5122 , \5123 );
not \U$4872 ( \5125 , \1081 );
and \U$4873 ( \5126 , \5121 , \5125 );
nor \U$4874 ( \5127 , \5124 , \5126 );
nand \U$4875 ( \5128 , \5116 , \5127 );
and \U$4876 ( \5129 , \3303 , RIbe29650_59);
not \U$4877 ( \5130 , RIbe29038_46);
nor \U$4878 ( \5131 , \5130 , \4065 );
nor \U$4879 ( \5132 , \5129 , \5131 );
and \U$4880 ( \5133 , \5132 , \1277 );
not \U$4881 ( \5134 , \5132 );
and \U$4882 ( \5135 , \5134 , \1076 );
nor \U$4883 ( \5136 , \5133 , \5135 );
not \U$4884 ( \5137 , \5136 );
and \U$4885 ( \5138 , \5128 , \5137 );
nor \U$4886 ( \5139 , \5116 , \5127 );
nor \U$4887 ( \5140 , \5138 , \5139 );
not \U$4888 ( \5141 , \5140 );
nand \U$4889 ( \5142 , \5108 , \5141 );
not \U$4890 ( \5143 , \5069 );
not \U$4891 ( \5144 , \5106 );
nand \U$4892 ( \5145 , \5143 , \5144 );
nand \U$4893 ( \5146 , \5142 , \5145 );
and \U$4894 ( \5147 , RIbe29380_53, RIbe27fd0_11);
and \U$4895 ( \5148 , \325 , RIbe27f58_10);
and \U$4896 ( \5149 , \330 , RIbe27e68_8);
nor \U$4897 ( \5150 , \5148 , \5149 );
not \U$4898 ( \5151 , \338 );
and \U$4899 ( \5152 , \5150 , \5151 );
not \U$4900 ( \5153 , \5150 );
and \U$4901 ( \5154 , \5153 , \1375 );
nor \U$4902 ( \5155 , \5152 , \5154 );
xor \U$4903 ( \5156 , \5147 , \5155 );
and \U$4904 ( \5157 , \260 , RIbe28660_25);
and \U$4905 ( \5158 , \1831 , RIbe285e8_24);
nor \U$4906 ( \5159 , \5157 , \5158 );
and \U$4907 ( \5160 , \5159 , \270 );
not \U$4908 ( \5161 , \5159 );
and \U$4909 ( \5162 , \5161 , \1663 );
nor \U$4910 ( \5163 , \5160 , \5162 );
and \U$4911 ( \5164 , \5156 , \5163 );
and \U$4912 ( \5165 , \5147 , \5155 );
or \U$4913 ( \5166 , \5164 , \5165 );
not \U$4914 ( \5167 , RIbe29560_57);
not \U$4915 ( \5168 , \4257 );
or \U$4916 ( \5169 , \5167 , \5168 );
nand \U$4917 ( \5170 , \1147 , RIbe28228_16);
nand \U$4918 ( \5171 , \5169 , \5170 );
and \U$4919 ( \5172 , \5171 , \1652 );
not \U$4920 ( \5173 , \5171 );
and \U$4921 ( \5174 , \5173 , \1152 );
nor \U$4922 ( \5175 , \5172 , \5174 );
not \U$4923 ( \5176 , \1611 );
not \U$4924 ( \5177 , RIbe28a20_33);
not \U$4925 ( \5178 , \5177 );
and \U$4926 ( \5179 , \5176 , \5178 );
and \U$4927 ( \5180 , \1744 , RIbe29290_51);
nor \U$4928 ( \5181 , \5179 , \5180 );
and \U$4929 ( \5182 , \5181 , \564 );
not \U$4930 ( \5183 , \5181 );
and \U$4931 ( \5184 , \5183 , \1621 );
nor \U$4932 ( \5185 , \5182 , \5184 );
xor \U$4933 ( \5186 , \5175 , \5185 );
and \U$4934 ( \5187 , \1807 , RIbe289a8_32);
and \U$4935 ( \5188 , \1165 , RIbe28930_31);
nor \U$4936 ( \5189 , \5187 , \5188 );
and \U$4937 ( \5190 , \5189 , \1608 );
not \U$4938 ( \5191 , \5189 );
and \U$4939 ( \5192 , \5191 , \1011 );
nor \U$4940 ( \5193 , \5190 , \5192 );
and \U$4941 ( \5194 , \5186 , \5193 );
and \U$4942 ( \5195 , \5175 , \5185 );
or \U$4943 ( \5196 , \5194 , \5195 );
xor \U$4944 ( \5197 , \5166 , \5196 );
not \U$4945 ( \5198 , RIbe28408_20);
not \U$4946 ( \5199 , \1337 );
or \U$4947 ( \5200 , \5198 , \5199 );
nand \U$4948 ( \5201 , \429 , RIbe28390_19);
nand \U$4949 ( \5202 , \5200 , \5201 );
and \U$4950 ( \5203 , \5202 , \306 );
not \U$4951 ( \5204 , \5202 );
and \U$4952 ( \5205 , \5204 , \1547 );
nor \U$4953 ( \5206 , \5203 , \5205 );
not \U$4954 ( \5207 , \5206 );
and \U$4955 ( \5208 , \1528 , RIbe287c8_28);
and \U$4956 ( \5209 , \1531 , RIbe28480_21);
nor \U$4957 ( \5210 , \5208 , \5209 );
and \U$4958 ( \5211 , \5210 , \300 );
not \U$4959 ( \5212 , \5210 );
and \U$4960 ( \5213 , \5212 , \293 );
nor \U$4961 ( \5214 , \5211 , \5213 );
not \U$4962 ( \5215 , \5214 );
or \U$4963 ( \5216 , \5207 , \5215 );
or \U$4964 ( \5217 , \5206 , \5214 );
not \U$4965 ( \5218 , RIbe28b10_35);
not \U$4966 ( \5219 , \548 );
or \U$4967 ( \5220 , \5218 , \5219 );
nand \U$4968 ( \5221 , \3775 , RIbe28b88_36);
nand \U$4969 ( \5222 , \5220 , \5221 );
not \U$4970 ( \5223 , \5222 );
not \U$4971 ( \5224 , \424 );
and \U$4972 ( \5225 , \5223 , \5224 );
and \U$4973 ( \5226 , \5222 , \424 );
nor \U$4974 ( \5227 , \5225 , \5226 );
not \U$4975 ( \5228 , \5227 );
nand \U$4976 ( \5229 , \5217 , \5228 );
nand \U$4977 ( \5230 , \5216 , \5229 );
and \U$4978 ( \5231 , \5197 , \5230 );
and \U$4979 ( \5232 , \5166 , \5196 );
or \U$4980 ( \5233 , \5231 , \5232 );
xor \U$4981 ( \5234 , \5146 , \5233 );
or \U$4982 ( \5235 , \4853 , \4854 );
nand \U$4983 ( \5236 , \5235 , \4855 );
xor \U$4984 ( \5237 , \4865 , \4884 );
xor \U$4985 ( \5238 , \5237 , \4874 );
xor \U$4986 ( \5239 , \5236 , \5238 );
not \U$4987 ( \5240 , \4896 );
not \U$4988 ( \5241 , \4916 );
or \U$4989 ( \5242 , \5240 , \5241 );
nand \U$4990 ( \5243 , \4915 , \4895 );
nand \U$4991 ( \5244 , \5242 , \5243 );
and \U$4992 ( \5245 , \5244 , \4918 );
not \U$4993 ( \5246 , \5244 );
and \U$4994 ( \5247 , \5246 , \4904 );
nor \U$4995 ( \5248 , \5245 , \5247 );
and \U$4996 ( \5249 , \5239 , \5248 );
and \U$4997 ( \5250 , \5236 , \5238 );
or \U$4998 ( \5251 , \5249 , \5250 );
and \U$4999 ( \5252 , \5234 , \5251 );
and \U$5000 ( \5253 , \5146 , \5233 );
or \U$5001 ( \5254 , \5252 , \5253 );
xor \U$5002 ( \5255 , \5042 , \5254 );
and \U$5003 ( \5256 , \4785 , \4773 );
not \U$5004 ( \5257 , \4785 );
and \U$5005 ( \5258 , \5257 , \4774 );
or \U$5006 ( \5259 , \5256 , \5258 );
xor \U$5007 ( \5260 , \5259 , \4797 );
not \U$5008 ( \5261 , \5260 );
and \U$5009 ( \5262 , \4736 , \4757 );
not \U$5010 ( \5263 , \4736 );
and \U$5011 ( \5264 , \5263 , \4756 );
or \U$5012 ( \5265 , \5262 , \5264 );
xnor \U$5013 ( \5266 , \5265 , \4746 );
not \U$5014 ( \5267 , \5266 );
or \U$5015 ( \5268 , \5261 , \5267 );
or \U$5016 ( \5269 , \5266 , \5260 );
xor \U$5017 ( \5270 , \4837 , \4815 );
xnor \U$5018 ( \5271 , \5270 , \4822 );
nand \U$5019 ( \5272 , \5269 , \5271 );
nand \U$5020 ( \5273 , \5268 , \5272 );
xor \U$5021 ( \5274 , \4929 , \4931 );
xor \U$5022 ( \5275 , \5274 , \4934 );
xor \U$5023 ( \5276 , \5273 , \5275 );
and \U$5024 ( \5277 , \4961 , \4952 );
not \U$5025 ( \5278 , \4961 );
and \U$5026 ( \5279 , \5278 , \4953 );
or \U$5027 ( \5280 , \5277 , \5279 );
xor \U$5028 ( \5281 , \5280 , \4943 );
and \U$5029 ( \5282 , \5276 , \5281 );
and \U$5030 ( \5283 , \5273 , \5275 );
or \U$5031 ( \5284 , \5282 , \5283 );
and \U$5032 ( \5285 , \5255 , \5284 );
and \U$5033 ( \5286 , \5042 , \5254 );
or \U$5034 ( \5287 , \5285 , \5286 );
xor \U$5035 ( \5288 , \4723 , \4725 );
xor \U$5036 ( \5289 , \4843 , \4923 );
xor \U$5037 ( \5290 , \5289 , \4937 );
xor \U$5038 ( \5291 , \5288 , \5290 );
xor \U$5039 ( \5292 , \4963 , \4965 );
xor \U$5040 ( \5293 , \5292 , \4968 );
and \U$5041 ( \5294 , \5291 , \5293 );
and \U$5042 ( \5295 , \5288 , \5290 );
or \U$5043 ( \5296 , \5294 , \5295 );
xor \U$5044 ( \5297 , \5287 , \5296 );
xor \U$5045 ( \5298 , \4975 , \4977 );
xor \U$5046 ( \5299 , \5298 , \4980 );
and \U$5047 ( \5300 , \5297 , \5299 );
and \U$5048 ( \5301 , \5287 , \5296 );
or \U$5049 ( \5302 , \5300 , \5301 );
xor \U$5050 ( \5303 , \5034 , \5302 );
xor \U$5051 ( \5304 , \4974 , \4983 );
xor \U$5052 ( \5305 , \5304 , \4986 );
and \U$5053 ( \5306 , \5303 , \5305 );
and \U$5054 ( \5307 , \5034 , \5302 );
or \U$5055 ( \5308 , \5306 , \5307 );
nand \U$5056 ( \5309 , \5032 , \5308 );
not \U$5057 ( \5310 , \5309 );
not \U$5058 ( \5311 , \5310 );
or \U$5059 ( \5312 , \5029 , \5311 );
nand \U$5060 ( \5313 , \5027 , \5309 );
nand \U$5061 ( \5314 , \5312 , \5313 );
and \U$5062 ( \5315 , \4995 , \5026 );
xor \U$5063 ( \5316 , \5004 , \5018 );
and \U$5064 ( \5317 , \5316 , \5025 );
and \U$5065 ( \5318 , \5004 , \5018 );
or \U$5066 ( \5319 , \5317 , \5318 );
xor \U$5067 ( \5320 , \5006 , \5010 );
and \U$5068 ( \5321 , \5320 , \5017 );
and \U$5069 ( \5322 , \5006 , \5010 );
or \U$5070 ( \5323 , \5321 , \5322 );
not \U$5071 ( \5324 , \5000 );
nand \U$5072 ( \5325 , \5324 , \4997 );
not \U$5073 ( \5326 , \5325 );
and \U$5074 ( \5327 , \5323 , \5326 );
not \U$5075 ( \5328 , \5323 );
and \U$5076 ( \5329 , \5328 , \5325 );
nor \U$5077 ( \5330 , \5327 , \5329 );
xor \U$5078 ( \5331 , \4102 , \4104 );
xor \U$5079 ( \5332 , \5331 , \4107 );
and \U$5080 ( \5333 , \5330 , \5332 );
not \U$5081 ( \5334 , \5330 );
not \U$5082 ( \5335 , \5332 );
and \U$5083 ( \5336 , \5334 , \5335 );
nor \U$5084 ( \5337 , \5333 , \5336 );
xor \U$5085 ( \5338 , \5319 , \5337 );
xor \U$5086 ( \5339 , \5315 , \5338 );
and \U$5087 ( \5340 , \5314 , \5339 );
xor \U$5088 ( \5341 , \5031 , \5308 );
xor \U$5089 ( \5342 , \4726 , \4940 );
xor \U$5090 ( \5343 , \5342 , \4971 );
and \U$5091 ( \5344 , \325 , RIbe27fd0_11);
and \U$5092 ( \5345 , \329 , RIbe27f58_10);
nor \U$5093 ( \5346 , \5344 , \5345 );
and \U$5094 ( \5347 , \5346 , \1375 );
not \U$5095 ( \5348 , \5346 );
and \U$5096 ( \5349 , \5348 , \1379 );
nor \U$5097 ( \5350 , \5347 , \5349 );
nand \U$5098 ( \5351 , RIbe29380_53, RIbe28ed0_43);
nand \U$5099 ( \5352 , \5350 , \5351 );
and \U$5100 ( \5353 , \1659 , RIbe27e68_8);
and \U$5101 ( \5354 , \1831 , RIbe28660_25);
nor \U$5102 ( \5355 , \5353 , \5354 );
and \U$5103 ( \5356 , \5355 , \270 );
not \U$5104 ( \5357 , \5355 );
and \U$5105 ( \5358 , \5357 , \1663 );
nor \U$5106 ( \5359 , \5356 , \5358 );
and \U$5107 ( \5360 , \5352 , \5359 );
nor \U$5108 ( \5361 , \5350 , \5351 );
nor \U$5109 ( \5362 , \5360 , \5361 );
not \U$5110 ( \5363 , \5362 );
not \U$5111 ( \5364 , \5363 );
not \U$5112 ( \5365 , \282 );
and \U$5113 ( \5366 , \5365 , RIbe285e8_24);
and \U$5114 ( \5367 , \1682 , RIbe287c8_28);
nor \U$5115 ( \5368 , \5366 , \5367 );
and \U$5116 ( \5369 , \5368 , \293 );
not \U$5117 ( \5370 , \5368 );
and \U$5118 ( \5371 , \5370 , \300 );
nor \U$5119 ( \5372 , \5369 , \5371 );
not \U$5120 ( \5373 , RIbe28390_19);
not \U$5121 ( \5374 , \3244 );
or \U$5122 ( \5375 , \5373 , \5374 );
nand \U$5123 ( \5376 , \3775 , RIbe28b10_35);
nand \U$5124 ( \5377 , \5375 , \5376 );
not \U$5125 ( \5378 , \5377 );
not \U$5126 ( \5379 , \424 );
and \U$5127 ( \5380 , \5378 , \5379 );
and \U$5128 ( \5381 , \5377 , \1333 );
nor \U$5129 ( \5382 , \5380 , \5381 );
and \U$5130 ( \5383 , \5372 , \5382 );
not \U$5131 ( \5384 , RIbe28480_21);
not \U$5132 ( \5385 , \1774 );
or \U$5133 ( \5386 , \5384 , \5385 );
nand \U$5134 ( \5387 , \429 , RIbe28408_20);
nand \U$5135 ( \5388 , \5386 , \5387 );
not \U$5136 ( \5389 , \5388 );
not \U$5137 ( \5390 , \1547 );
and \U$5138 ( \5391 , \5389 , \5390 );
and \U$5139 ( \5392 , \5388 , \1547 );
nor \U$5140 ( \5393 , \5391 , \5392 );
nor \U$5141 ( \5394 , \5383 , \5393 );
nor \U$5142 ( \5395 , \5372 , \5382 );
nor \U$5143 ( \5396 , \5394 , \5395 );
not \U$5144 ( \5397 , \5396 );
not \U$5145 ( \5398 , \5397 );
or \U$5146 ( \5399 , \5364 , \5398 );
nand \U$5147 ( \5400 , \5396 , \5362 );
and \U$5148 ( \5401 , \1807 , RIbe28a20_33);
and \U$5149 ( \5402 , \1203 , RIbe289a8_32);
nor \U$5150 ( \5403 , \5401 , \5402 );
and \U$5151 ( \5404 , \5403 , \1011 );
not \U$5152 ( \5405 , \5403 );
and \U$5153 ( \5406 , \5405 , \1813 );
nor \U$5154 ( \5407 , \5404 , \5406 );
not \U$5155 ( \5408 , \5407 );
not \U$5156 ( \5409 , \5408 );
not \U$5157 ( \5410 , RIbe28930_31);
not \U$5158 ( \5411 , \4257 );
or \U$5159 ( \5412 , \5410 , \5411 );
nand \U$5160 ( \5413 , \1147 , RIbe29560_57);
nand \U$5161 ( \5414 , \5412 , \5413 );
and \U$5162 ( \5415 , \5414 , \1154 );
not \U$5163 ( \5416 , \5414 );
and \U$5164 ( \5417 , \5416 , \1157 );
nor \U$5165 ( \5418 , \5415 , \5417 );
not \U$5166 ( \5419 , \5418 );
or \U$5167 ( \5420 , \5409 , \5419 );
or \U$5168 ( \5421 , \5418 , \5408 );
not \U$5169 ( \5422 , \1611 );
not \U$5170 ( \5423 , RIbe29290_51);
not \U$5171 ( \5424 , \5423 );
and \U$5172 ( \5425 , \5422 , \5424 );
and \U$5173 ( \5426 , \1744 , RIbe28b88_36);
nor \U$5174 ( \5427 , \5425 , \5426 );
and \U$5175 ( \5428 , \5427 , \672 );
not \U$5176 ( \5429 , \5427 );
and \U$5177 ( \5430 , \5429 , \564 );
or \U$5178 ( \5431 , \5428 , \5430 );
nand \U$5179 ( \5432 , \5421 , \5431 );
nand \U$5180 ( \5433 , \5420 , \5432 );
nand \U$5181 ( \5434 , \5400 , \5433 );
nand \U$5182 ( \5435 , \5399 , \5434 );
not \U$5183 ( \5436 , RIbe28de0_41);
not \U$5184 ( \5437 , \4830 );
or \U$5185 ( \5438 , \5436 , \5437 );
nand \U$5186 ( \5439 , \5052 , RIbe29920_65);
nand \U$5187 ( \5440 , \5438 , \5439 );
and \U$5188 ( \5441 , \5440 , \4586 );
not \U$5189 ( \5442 , \5440 );
and \U$5190 ( \5443 , \5442 , \4592 );
nor \U$5191 ( \5444 , \5441 , \5443 );
not \U$5192 ( \5445 , RIbe27c10_3);
not \U$5193 ( \5446 , \4804 );
or \U$5194 ( \5447 , \5445 , \5446 );
nand \U$5195 ( \5448 , \4600 , RIbe28e58_42);
nand \U$5196 ( \5449 , \5447 , \5448 );
xnor \U$5197 ( \5450 , \4323 , \5449 );
or \U$5198 ( \5451 , \5444 , \5450 );
xnor \U$5199 ( \5452 , RIbe27b20_1, RIbe29b78_70);
xor \U$5200 ( \5453 , RIbe28cf0_39, RIbe27b20_1);
nand \U$5201 ( \5454 , \5452 , \5453 );
not \U$5202 ( \5455 , \5454 );
nand \U$5203 ( \5456 , \5455 , RIbe27b98_2);
not \U$5204 ( \5457 , \5045 );
and \U$5205 ( \5458 , \5456 , \5457 );
not \U$5206 ( \5459 , \5456 );
not \U$5207 ( \5460 , \5044 );
and \U$5208 ( \5461 , \5459 , \5460 );
nor \U$5209 ( \5462 , \5458 , \5461 );
nand \U$5210 ( \5463 , \5451 , \5462 );
nand \U$5211 ( \5464 , \5450 , \5444 );
nand \U$5212 ( \5465 , \5463 , \5464 );
and \U$5213 ( \5466 , \4749 , RIbe280c0_13);
buf \U$5214 ( \5467 , \1116 );
and \U$5215 ( \5468 , \5467 , RIbe29830_63);
nor \U$5216 ( \5469 , \5466 , \5468 );
and \U$5217 ( \5470 , \5469 , \1448 );
not \U$5218 ( \5471 , \5469 );
and \U$5219 ( \5472 , \5471 , \1131 );
nor \U$5220 ( \5473 , \5470 , \5472 );
not \U$5221 ( \5474 , \5473 );
not \U$5222 ( \5475 , RIbe28228_16);
not \U$5223 ( \5476 , \1093 );
not \U$5224 ( \5477 , \5476 );
or \U$5225 ( \5478 , \5475 , \5477 );
nand \U$5226 ( \5479 , \1455 , RIbe281b0_15);
nand \U$5227 ( \5480 , \5478 , \5479 );
not \U$5228 ( \5481 , \5480 );
not \U$5229 ( \5482 , \5125 );
and \U$5230 ( \5483 , \5481 , \5482 );
and \U$5231 ( \5484 , \5480 , \4251 );
nor \U$5232 ( \5485 , \5483 , \5484 );
not \U$5233 ( \5486 , \5485 );
not \U$5234 ( \5487 , \5486 );
or \U$5235 ( \5488 , \5474 , \5487 );
not \U$5236 ( \5489 , \5485 );
not \U$5237 ( \5490 , \5473 );
not \U$5238 ( \5491 , \5490 );
or \U$5239 ( \5492 , \5489 , \5491 );
and \U$5240 ( \5493 , \3303 , RIbe296c8_60);
not \U$5241 ( \5494 , RIbe29650_59);
nor \U$5242 ( \5495 , \4065 , \5494 );
nor \U$5243 ( \5496 , \5493 , \5495 );
and \U$5244 ( \5497 , \5496 , \1277 );
not \U$5245 ( \5498 , \5496 );
and \U$5246 ( \5499 , \5498 , \3516 );
nor \U$5247 ( \5500 , \5497 , \5499 );
not \U$5248 ( \5501 , \5500 );
nand \U$5249 ( \5502 , \5492 , \5501 );
nand \U$5250 ( \5503 , \5488 , \5502 );
xor \U$5251 ( \5504 , \5465 , \5503 );
not \U$5252 ( \5505 , RIbe29038_46);
not \U$5253 ( \5506 , \3476 );
or \U$5254 ( \5507 , \5505 , \5506 );
nand \U$5255 ( \5508 , \4284 , RIbe28fc0_45);
nand \U$5256 ( \5509 , \5507 , \5508 );
and \U$5257 ( \5510 , \5509 , \3272 );
not \U$5258 ( \5511 , \5509 );
and \U$5259 ( \5512 , \5511 , \3275 );
nor \U$5260 ( \5513 , \5510 , \5512 );
not \U$5261 ( \5514 , RIbe27d78_6);
not \U$5262 ( \5515 , \5094 );
or \U$5263 ( \5516 , \5514 , \5515 );
nand \U$5264 ( \5517 , \4333 , RIbe27d00_5);
nand \U$5265 ( \5518 , \5516 , \5517 );
and \U$5266 ( \5519 , \5518 , \3471 );
not \U$5267 ( \5520 , \5518 );
and \U$5268 ( \5521 , \5520 , \3448 );
nor \U$5269 ( \5522 , \5519 , \5521 );
xor \U$5270 ( \5523 , \5513 , \5522 );
not \U$5271 ( \5524 , RIbe290b0_47);
not \U$5272 ( \5525 , \3285 );
or \U$5273 ( \5526 , \5524 , \5525 );
nand \U$5274 ( \5527 , \3458 , RIbe29a88_68);
nand \U$5275 ( \5528 , \5526 , \5527 );
and \U$5276 ( \5529 , \5528 , \4346 );
not \U$5277 ( \5530 , \5528 );
and \U$5278 ( \5531 , \5530 , \3461 );
nor \U$5279 ( \5532 , \5529 , \5531 );
and \U$5280 ( \5533 , \5523 , \5532 );
and \U$5281 ( \5534 , \5513 , \5522 );
or \U$5282 ( \5535 , \5533 , \5534 );
and \U$5283 ( \5536 , \5504 , \5535 );
and \U$5284 ( \5537 , \5465 , \5503 );
or \U$5285 ( \5538 , \5536 , \5537 );
xor \U$5286 ( \5539 , \5435 , \5538 );
xor \U$5287 ( \5540 , \5175 , \5185 );
xor \U$5288 ( \5541 , \5540 , \5193 );
not \U$5289 ( \5542 , \5541 );
not \U$5290 ( \5543 , \5542 );
not \U$5291 ( \5544 , \5228 );
not \U$5292 ( \5545 , \5207 );
or \U$5293 ( \5546 , \5544 , \5545 );
nand \U$5294 ( \5547 , \5206 , \5227 );
nand \U$5295 ( \5548 , \5546 , \5547 );
and \U$5296 ( \5549 , \5548 , \5215 );
not \U$5297 ( \5550 , \5548 );
and \U$5298 ( \5551 , \5550 , \5214 );
nor \U$5299 ( \5552 , \5549 , \5551 );
not \U$5300 ( \5553 , \5552 );
or \U$5301 ( \5554 , \5543 , \5553 );
xor \U$5302 ( \5555 , \5147 , \5155 );
xor \U$5303 ( \5556 , \5555 , \5163 );
nand \U$5304 ( \5557 , \5554 , \5556 );
not \U$5305 ( \5558 , \5552 );
nand \U$5306 ( \5559 , \5558 , \5541 );
nand \U$5307 ( \5560 , \5557 , \5559 );
and \U$5308 ( \5561 , \5539 , \5560 );
and \U$5309 ( \5562 , \5435 , \5538 );
or \U$5310 ( \5563 , \5561 , \5562 );
not \U$5311 ( \5564 , \5069 );
not \U$5312 ( \5565 , \5141 );
not \U$5313 ( \5566 , \5106 );
or \U$5314 ( \5567 , \5565 , \5566 );
nand \U$5315 ( \5568 , \5144 , \5140 );
nand \U$5316 ( \5569 , \5567 , \5568 );
not \U$5317 ( \5570 , \5569 );
or \U$5318 ( \5571 , \5564 , \5570 );
or \U$5319 ( \5572 , \5569 , \5069 );
nand \U$5320 ( \5573 , \5571 , \5572 );
xor \U$5321 ( \5574 , \5166 , \5196 );
xor \U$5322 ( \5575 , \5574 , \5230 );
and \U$5323 ( \5576 , \5573 , \5575 );
xor \U$5324 ( \5577 , \5563 , \5576 );
xor \U$5325 ( \5578 , \5047 , \5055 );
xor \U$5326 ( \5579 , \5578 , \5066 );
not \U$5327 ( \5580 , \5579 );
not \U$5328 ( \5581 , \5081 );
not \U$5329 ( \5582 , \5103 );
or \U$5330 ( \5583 , \5581 , \5582 );
nand \U$5331 ( \5584 , \5102 , \5080 );
nand \U$5332 ( \5585 , \5583 , \5584 );
xnor \U$5333 ( \5586 , \5585 , \5091 );
not \U$5334 ( \5587 , \5586 );
not \U$5335 ( \5588 , \5587 );
or \U$5336 ( \5589 , \5580 , \5588 );
not \U$5337 ( \5590 , \5137 );
not \U$5338 ( \5591 , \5116 );
or \U$5339 ( \5592 , \5590 , \5591 );
nand \U$5340 ( \5593 , \5115 , \5136 );
nand \U$5341 ( \5594 , \5592 , \5593 );
xnor \U$5342 ( \5595 , \5594 , \5127 );
nand \U$5343 ( \5596 , \5589 , \5595 );
not \U$5344 ( \5597 , \5579 );
nand \U$5345 ( \5598 , \5597 , \5586 );
nand \U$5346 ( \5599 , \5596 , \5598 );
xor \U$5347 ( \5600 , \5236 , \5238 );
xor \U$5348 ( \5601 , \5600 , \5248 );
xor \U$5349 ( \5602 , \5599 , \5601 );
xor \U$5350 ( \5603 , \5271 , \5266 );
xor \U$5351 ( \5604 , \5603 , \5260 );
and \U$5352 ( \5605 , \5602 , \5604 );
and \U$5353 ( \5606 , \5599 , \5601 );
or \U$5354 ( \5607 , \5605 , \5606 );
and \U$5355 ( \5608 , \5577 , \5607 );
and \U$5356 ( \5609 , \5563 , \5576 );
or \U$5357 ( \5610 , \5608 , \5609 );
xor \U$5358 ( \5611 , \5288 , \5290 );
xor \U$5359 ( \5612 , \5611 , \5293 );
xor \U$5360 ( \5613 , \5610 , \5612 );
xor \U$5361 ( \5614 , \5036 , \5041 );
xor \U$5362 ( \5615 , \5146 , \5233 );
xor \U$5363 ( \5616 , \5615 , \5251 );
xor \U$5364 ( \5617 , \5614 , \5616 );
xor \U$5365 ( \5618 , \5273 , \5275 );
xor \U$5366 ( \5619 , \5618 , \5281 );
and \U$5367 ( \5620 , \5617 , \5619 );
and \U$5368 ( \5621 , \5614 , \5616 );
or \U$5369 ( \5622 , \5620 , \5621 );
and \U$5370 ( \5623 , \5613 , \5622 );
and \U$5371 ( \5624 , \5610 , \5612 );
or \U$5372 ( \5625 , \5623 , \5624 );
xor \U$5373 ( \5626 , \5343 , \5625 );
xor \U$5374 ( \5627 , \5287 , \5296 );
xor \U$5375 ( \5628 , \5627 , \5299 );
and \U$5376 ( \5629 , \5626 , \5628 );
and \U$5377 ( \5630 , \5343 , \5625 );
or \U$5378 ( \5631 , \5629 , \5630 );
xor \U$5379 ( \5632 , \5034 , \5302 );
xor \U$5380 ( \5633 , \5632 , \5305 );
and \U$5381 ( \5634 , \5631 , \5633 );
xor \U$5382 ( \5635 , \5341 , \5634 );
not \U$5383 ( \5636 , \5635 );
xor \U$5384 ( \5637 , \5042 , \5254 );
xor \U$5385 ( \5638 , \5637 , \5284 );
xor \U$5386 ( \5639 , \5465 , \5503 );
xor \U$5387 ( \5640 , \5639 , \5535 );
not \U$5388 ( \5641 , \5640 );
xor \U$5389 ( \5642 , \5362 , \5397 );
xor \U$5390 ( \5643 , \5642 , \5433 );
nor \U$5391 ( \5644 , \5641 , \5643 );
xor \U$5392 ( \5645 , \5350 , \5359 );
xnor \U$5393 ( \5646 , \5645 , \5351 );
xor \U$5394 ( \5647 , \5393 , \5382 );
xor \U$5395 ( \5648 , \5647 , \5372 );
nand \U$5396 ( \5649 , \5646 , \5648 );
not \U$5397 ( \5650 , RIbe28fc0_45);
not \U$5398 ( \5651 , \4764 );
or \U$5399 ( \5652 , \5650 , \5651 );
nand \U$5400 ( \5653 , \3689 , RIbe290b0_47);
nand \U$5401 ( \5654 , \5652 , \5653 );
not \U$5402 ( \5655 , \5654 );
not \U$5403 ( \5656 , \3461 );
and \U$5404 ( \5657 , \5655 , \5656 );
and \U$5405 ( \5658 , \5654 , \3461 );
nor \U$5406 ( \5659 , \5657 , \5658 );
not \U$5407 ( \5660 , \5659 );
not \U$5408 ( \5661 , RIbe27d00_5);
not \U$5409 ( \5662 , \5058 );
or \U$5410 ( \5663 , \5661 , \5662 );
nand \U$5411 ( \5664 , \4809 , RIbe27c10_3);
nand \U$5412 ( \5665 , \5663 , \5664 );
and \U$5413 ( \5666 , \5665 , \4323 );
not \U$5414 ( \5667 , \5665 );
and \U$5415 ( \5668 , \5667 , \4603 );
nor \U$5416 ( \5669 , \5666 , \5668 );
not \U$5417 ( \5670 , \5669 );
or \U$5418 ( \5671 , \5660 , \5670 );
not \U$5419 ( \5672 , RIbe29a88_68);
not \U$5420 ( \5673 , \4021 );
or \U$5421 ( \5674 , \5672 , \5673 );
nand \U$5422 ( \5675 , \4027 , RIbe27d78_6);
nand \U$5423 ( \5676 , \5674 , \5675 );
and \U$5424 ( \5677 , \5676 , \4821 );
not \U$5425 ( \5678 , \5676 );
and \U$5426 ( \5679 , \5678 , \3471 );
nor \U$5427 ( \5680 , \5677 , \5679 );
not \U$5428 ( \5681 , \5680 );
nand \U$5429 ( \5682 , \5671 , \5681 );
not \U$5430 ( \5683 , \5669 );
not \U$5431 ( \5684 , \5659 );
nand \U$5432 ( \5685 , \5683 , \5684 );
and \U$5433 ( \5686 , \5682 , \5685 );
not \U$5434 ( \5687 , \5686 );
not \U$5435 ( \5688 , \5687 );
not \U$5436 ( \5689 , RIbe29650_59);
not \U$5437 ( \5690 , \2898 );
or \U$5438 ( \5691 , \5689 , \5690 );
nand \U$5439 ( \5692 , \4284 , RIbe29038_46);
nand \U$5440 ( \5693 , \5691 , \5692 );
and \U$5441 ( \5694 , \5693 , \2379 );
not \U$5442 ( \5695 , \5693 );
and \U$5443 ( \5696 , \5695 , \4287 );
nor \U$5444 ( \5697 , \5694 , \5696 );
not \U$5445 ( \5698 , \5697 );
not \U$5446 ( \5699 , \5698 );
and \U$5447 ( \5700 , \4749 , RIbe281b0_15);
and \U$5448 ( \5701 , \1117 , RIbe280c0_13);
nor \U$5449 ( \5702 , \5700 , \5701 );
and \U$5450 ( \5703 , \5702 , \1132 );
not \U$5451 ( \5704 , \5702 );
and \U$5452 ( \5705 , \5704 , \3491 );
nor \U$5453 ( \5706 , \5703 , \5705 );
not \U$5454 ( \5707 , \5706 );
not \U$5455 ( \5708 , \5707 );
or \U$5456 ( \5709 , \5699 , \5708 );
not \U$5457 ( \5710 , \5706 );
not \U$5458 ( \5711 , \5697 );
or \U$5459 ( \5712 , \5710 , \5711 );
and \U$5460 ( \5713 , \4295 , RIbe29830_63);
not \U$5461 ( \5714 , RIbe296c8_60);
nor \U$5462 ( \5715 , \5714 , \2889 );
nor \U$5463 ( \5716 , \5713 , \5715 );
and \U$5464 ( \5717 , \5716 , \1277 );
not \U$5465 ( \5718 , \5716 );
and \U$5466 ( \5719 , \5718 , \1076 );
nor \U$5467 ( \5720 , \5717 , \5719 );
not \U$5468 ( \5721 , \5720 );
nand \U$5469 ( \5722 , \5712 , \5721 );
nand \U$5470 ( \5723 , \5709 , \5722 );
not \U$5471 ( \5724 , \5723 );
or \U$5472 ( \5725 , \5688 , \5724 );
not \U$5473 ( \5726 , RIbe28e58_42);
not \U$5474 ( \5727 , \4828 );
not \U$5475 ( \5728 , \5727 );
or \U$5476 ( \5729 , \5726 , \5728 );
buf \U$5477 ( \5730 , \4824 );
buf \U$5478 ( \5731 , \5730 );
nand \U$5479 ( \5732 , \5731 , RIbe28de0_41);
nand \U$5480 ( \5733 , \5729 , \5732 );
and \U$5481 ( \5734 , \5733 , \4592 );
not \U$5482 ( \5735 , \5733 );
and \U$5483 ( \5736 , \5735 , \4586 );
nor \U$5484 ( \5737 , \5734 , \5736 );
nand \U$5485 ( \5738 , RIbe29ce0_73, RIbe29d58_74);
nand \U$5486 ( \5739 , \5738 , RIbe29b78_70);
buf \U$5487 ( \5740 , \5739 );
not \U$5488 ( \5741 , \5740 );
nand \U$5489 ( \5742 , \5737 , \5741 );
not \U$5490 ( \5743 , RIbe29920_65);
not \U$5491 ( \5744 , \5455 );
or \U$5492 ( \5745 , \5743 , \5744 );
xor \U$5493 ( \5746 , RIbe27b20_1, RIbe29b78_70);
not \U$5494 ( \5747 , \5746 );
not \U$5495 ( \5748 , \5747 );
buf \U$5496 ( \5749 , \5748 );
not \U$5497 ( \5750 , \5749 );
not \U$5498 ( \5751 , \5750 );
nand \U$5499 ( \5752 , \5751 , RIbe27b98_2);
nand \U$5500 ( \5753 , \5745 , \5752 );
not \U$5501 ( \5754 , \5460 );
and \U$5502 ( \5755 , \5753 , \5754 );
not \U$5503 ( \5756 , \5753 );
and \U$5504 ( \5757 , \5756 , \5047 );
or \U$5505 ( \5758 , \5755 , \5757 );
and \U$5506 ( \5759 , \5742 , \5758 );
nor \U$5507 ( \5760 , \5737 , \5741 );
nor \U$5508 ( \5761 , \5759 , \5760 );
not \U$5509 ( \5762 , \5761 );
not \U$5510 ( \5763 , \5723 );
nand \U$5511 ( \5764 , \5763 , \5686 );
nand \U$5512 ( \5765 , \5762 , \5764 );
nand \U$5513 ( \5766 , \5725 , \5765 );
xor \U$5514 ( \5767 , \5649 , \5766 );
not \U$5515 ( \5768 , RIbe28408_20);
not \U$5516 ( \5769 , \3244 );
or \U$5517 ( \5770 , \5768 , \5769 );
nand \U$5518 ( \5771 , \3775 , RIbe28390_19);
nand \U$5519 ( \5772 , \5770 , \5771 );
and \U$5520 ( \5773 , \5772 , \3415 );
not \U$5521 ( \5774 , \5772 );
and \U$5522 ( \5775 , \5774 , \424 );
nor \U$5523 ( \5776 , \5773 , \5775 );
not \U$5524 ( \5777 , RIbe287c8_28);
not \U$5525 ( \5778 , \383 );
or \U$5526 ( \5779 , \5777 , \5778 );
nand \U$5527 ( \5780 , \429 , RIbe28480_21);
nand \U$5528 ( \5781 , \5779 , \5780 );
and \U$5529 ( \5782 , \5781 , \306 );
not \U$5530 ( \5783 , \5781 );
and \U$5531 ( \5784 , \5783 , \3175 );
nor \U$5532 ( \5785 , \5782 , \5784 );
or \U$5533 ( \5786 , \5776 , \5785 );
not \U$5534 ( \5787 , RIbe28b10_35);
not \U$5535 ( \5788 , \664 );
or \U$5536 ( \5789 , \5787 , \5788 );
nand \U$5537 ( \5790 , \1180 , RIbe28b88_36);
nand \U$5538 ( \5791 , \5789 , \5790 );
not \U$5539 ( \5792 , \5791 );
not \U$5540 ( \5793 , \564 );
and \U$5541 ( \5794 , \5792 , \5793 );
and \U$5542 ( \5795 , \5791 , \1618 );
nor \U$5543 ( \5796 , \5794 , \5795 );
not \U$5544 ( \5797 , \5796 );
nand \U$5545 ( \5798 , \5786 , \5797 );
nand \U$5546 ( \5799 , \5776 , \5785 );
nand \U$5547 ( \5800 , \5798 , \5799 );
and \U$5548 ( \5801 , \325 , RIbe28ed0_43);
and \U$5549 ( \5802 , \1371 , RIbe27fd0_11);
nor \U$5550 ( \5803 , \5801 , \5802 );
and \U$5551 ( \5804 , \5803 , \1374 );
not \U$5552 ( \5805 , \5803 );
and \U$5553 ( \5806 , \5805 , \1375 );
nor \U$5554 ( \5807 , \5804 , \5806 );
not \U$5555 ( \5808 , \5807 );
and \U$5556 ( \5809 , \283 , RIbe28660_25);
and \U$5557 ( \5810 , \1531 , RIbe285e8_24);
nor \U$5558 ( \5811 , \5809 , \5810 );
and \U$5559 ( \5812 , \5811 , \293 );
not \U$5560 ( \5813 , \5811 );
and \U$5561 ( \5814 , \5813 , \300 );
nor \U$5562 ( \5815 , \5812 , \5814 );
not \U$5563 ( \5816 , \5815 );
not \U$5564 ( \5817 , \5816 );
or \U$5565 ( \5818 , \5808 , \5817 );
or \U$5566 ( \5819 , \5816 , \5807 );
and \U$5567 ( \5820 , \1357 , RIbe27f58_10);
and \U$5568 ( \5821 , \264 , RIbe27e68_8);
nor \U$5569 ( \5822 , \5820 , \5821 );
and \U$5570 ( \5823 , \5822 , \270 );
not \U$5571 ( \5824 , \5822 );
and \U$5572 ( \5825 , \5824 , \1663 );
nor \U$5573 ( \5826 , \5823 , \5825 );
nand \U$5574 ( \5827 , \5819 , \5826 );
nand \U$5575 ( \5828 , \5818 , \5827 );
xor \U$5576 ( \5829 , \5800 , \5828 );
not \U$5577 ( \5830 , RIbe289a8_32);
not \U$5578 ( \5831 , \2597 );
or \U$5579 ( \5832 , \5830 , \5831 );
nand \U$5580 ( \5833 , \1147 , RIbe28930_31);
nand \U$5581 ( \5834 , \5832 , \5833 );
and \U$5582 ( \5835 , \5834 , \1469 );
not \U$5583 ( \5836 , \5834 );
and \U$5584 ( \5837 , \5836 , \1153 );
nor \U$5585 ( \5838 , \5835 , \5837 );
and \U$5586 ( \5839 , \1807 , RIbe29290_51);
and \U$5587 ( \5840 , \1165 , RIbe28a20_33);
nor \U$5588 ( \5841 , \5839 , \5840 );
and \U$5589 ( \5842 , \5841 , \1608 );
not \U$5590 ( \5843 , \5841 );
and \U$5591 ( \5844 , \5843 , \1011 );
nor \U$5592 ( \5845 , \5842 , \5844 );
xor \U$5593 ( \5846 , \5838 , \5845 );
not \U$5594 ( \5847 , RIbe29560_57);
not \U$5595 ( \5848 , \1298 );
or \U$5596 ( \5849 , \5847 , \5848 );
nand \U$5597 ( \5850 , \1455 , RIbe28228_16);
nand \U$5598 ( \5851 , \5849 , \5850 );
and \U$5599 ( \5852 , \5851 , \1309 );
not \U$5600 ( \5853 , \5851 );
and \U$5601 ( \5854 , \5853 , \2418 );
nor \U$5602 ( \5855 , \5852 , \5854 );
and \U$5603 ( \5856 , \5846 , \5855 );
and \U$5604 ( \5857 , \5838 , \5845 );
or \U$5605 ( \5858 , \5856 , \5857 );
and \U$5606 ( \5859 , \5829 , \5858 );
and \U$5607 ( \5860 , \5800 , \5828 );
or \U$5608 ( \5861 , \5859 , \5860 );
and \U$5609 ( \5862 , \5767 , \5861 );
and \U$5610 ( \5863 , \5649 , \5766 );
or \U$5611 ( \5864 , \5862 , \5863 );
xor \U$5612 ( \5865 , \5644 , \5864 );
and \U$5613 ( \5866 , \5418 , \5407 );
not \U$5614 ( \5867 , \5418 );
and \U$5615 ( \5868 , \5867 , \5408 );
or \U$5616 ( \5869 , \5866 , \5868 );
xnor \U$5617 ( \5870 , \5869 , \5431 );
not \U$5618 ( \5871 , \5870 );
not \U$5619 ( \5872 , \5871 );
xor \U$5620 ( \5873 , \5513 , \5522 );
xor \U$5621 ( \5874 , \5873 , \5532 );
not \U$5622 ( \5875 , \5874 );
or \U$5623 ( \5876 , \5872 , \5875 );
not \U$5624 ( \5877 , \5874 );
nand \U$5625 ( \5878 , \5877 , \5870 );
not \U$5626 ( \5879 , \5501 );
not \U$5627 ( \5880 , \5490 );
or \U$5628 ( \5881 , \5879 , \5880 );
nand \U$5629 ( \5882 , \5473 , \5500 );
nand \U$5630 ( \5883 , \5881 , \5882 );
and \U$5631 ( \5884 , \5883 , \5485 );
not \U$5632 ( \5885 , \5883 );
and \U$5633 ( \5886 , \5885 , \5486 );
nor \U$5634 ( \5887 , \5884 , \5886 );
not \U$5635 ( \5888 , \5887 );
nand \U$5636 ( \5889 , \5878 , \5888 );
nand \U$5637 ( \5890 , \5876 , \5889 );
xor \U$5638 ( \5891 , \5552 , \5556 );
xor \U$5639 ( \5892 , \5891 , \5542 );
xor \U$5640 ( \5893 , \5890 , \5892 );
not \U$5641 ( \5894 , \5579 );
and \U$5642 ( \5895 , \5595 , \5587 );
not \U$5643 ( \5896 , \5595 );
and \U$5644 ( \5897 , \5896 , \5586 );
or \U$5645 ( \5898 , \5895 , \5897 );
not \U$5646 ( \5899 , \5898 );
or \U$5647 ( \5900 , \5894 , \5899 );
or \U$5648 ( \5901 , \5898 , \5579 );
nand \U$5649 ( \5902 , \5900 , \5901 );
and \U$5650 ( \5903 , \5893 , \5902 );
and \U$5651 ( \5904 , \5890 , \5892 );
or \U$5652 ( \5905 , \5903 , \5904 );
and \U$5653 ( \5906 , \5865 , \5905 );
and \U$5654 ( \5907 , \5644 , \5864 );
or \U$5655 ( \5908 , \5906 , \5907 );
not \U$5656 ( \5909 , \5908 );
xor \U$5657 ( \5910 , \5599 , \5601 );
xor \U$5658 ( \5911 , \5910 , \5604 );
xor \U$5659 ( \5912 , \5573 , \5575 );
not \U$5660 ( \5913 , \5912 );
xor \U$5661 ( \5914 , \5435 , \5538 );
xor \U$5662 ( \5915 , \5914 , \5560 );
not \U$5663 ( \5916 , \5915 );
nand \U$5664 ( \5917 , \5913 , \5916 );
and \U$5665 ( \5918 , \5911 , \5917 );
and \U$5666 ( \5919 , \5915 , \5912 );
nor \U$5667 ( \5920 , \5918 , \5919 );
not \U$5668 ( \5921 , \5920 );
not \U$5669 ( \5922 , \5921 );
or \U$5670 ( \5923 , \5909 , \5922 );
or \U$5671 ( \5924 , \5921 , \5908 );
xor \U$5672 ( \5925 , \5614 , \5616 );
xor \U$5673 ( \5926 , \5925 , \5619 );
nand \U$5674 ( \5927 , \5924 , \5926 );
nand \U$5675 ( \5928 , \5923 , \5927 );
xor \U$5676 ( \5929 , \5638 , \5928 );
xor \U$5677 ( \5930 , \5610 , \5612 );
xor \U$5678 ( \5931 , \5930 , \5622 );
and \U$5679 ( \5932 , \5929 , \5931 );
and \U$5680 ( \5933 , \5638 , \5928 );
or \U$5681 ( \5934 , \5932 , \5933 );
xor \U$5682 ( \5935 , \5343 , \5625 );
xor \U$5683 ( \5936 , \5935 , \5628 );
and \U$5684 ( \5937 , \5934 , \5936 );
xor \U$5685 ( \5938 , \5631 , \5633 );
xor \U$5686 ( \5939 , \5937 , \5938 );
xor \U$5687 ( \5940 , \5638 , \5928 );
xor \U$5688 ( \5941 , \5940 , \5931 );
xor \U$5689 ( \5942 , \5563 , \5576 );
xor \U$5690 ( \5943 , \5942 , \5607 );
not \U$5691 ( \5944 , \5943 );
xor \U$5692 ( \5945 , \5920 , \5908 );
xor \U$5693 ( \5946 , \5945 , \5926 );
not \U$5694 ( \5947 , \5946 );
not \U$5695 ( \5948 , \5947 );
or \U$5696 ( \5949 , \5944 , \5948 );
not \U$5697 ( \5950 , \5943 );
nand \U$5698 ( \5951 , \5950 , \5946 );
and \U$5699 ( \5952 , \5826 , \5815 );
not \U$5700 ( \5953 , \5826 );
and \U$5701 ( \5954 , \5953 , \5816 );
or \U$5702 ( \5955 , \5952 , \5954 );
not \U$5703 ( \5956 , \5807 );
and \U$5704 ( \5957 , \5955 , \5956 );
not \U$5705 ( \5958 , \5955 );
and \U$5706 ( \5959 , \5958 , \5807 );
nor \U$5707 ( \5960 , \5957 , \5959 );
nand \U$5708 ( \5961 , RIbe29380_53, RIbe28f48_44);
nand \U$5709 ( \5962 , \5960 , \5961 );
not \U$5710 ( \5963 , \5785 );
not \U$5711 ( \5964 , \5963 );
xnor \U$5712 ( \5965 , \5776 , \5796 );
not \U$5713 ( \5966 , \5965 );
or \U$5714 ( \5967 , \5964 , \5966 );
or \U$5715 ( \5968 , \5965 , \5963 );
nand \U$5716 ( \5969 , \5967 , \5968 );
and \U$5717 ( \5970 , \5962 , \5969 );
nor \U$5718 ( \5971 , \5960 , \5961 );
nor \U$5719 ( \5972 , \5970 , \5971 );
not \U$5720 ( \5973 , \1160 );
and \U$5721 ( \5974 , \5973 , RIbe28b88_36);
and \U$5722 ( \5975 , \1165 , RIbe29290_51);
nor \U$5723 ( \5976 , \5974 , \5975 );
and \U$5724 ( \5977 , \5976 , \1011 );
not \U$5725 ( \5978 , \5976 );
and \U$5726 ( \5979 , \5978 , \1813 );
nor \U$5727 ( \5980 , \5977 , \5979 );
not \U$5728 ( \5981 , RIbe28a20_33);
not \U$5729 ( \5982 , \1143 );
or \U$5730 ( \5983 , \5981 , \5982 );
nand \U$5731 ( \5984 , \1147 , RIbe289a8_32);
nand \U$5732 ( \5985 , \5983 , \5984 );
not \U$5733 ( \5986 , \5985 );
not \U$5734 ( \5987 , \1153 );
and \U$5735 ( \5988 , \5986 , \5987 );
and \U$5736 ( \5989 , \5985 , \1152 );
nor \U$5737 ( \5990 , \5988 , \5989 );
and \U$5738 ( \5991 , \5980 , \5990 );
not \U$5739 ( \5992 , RIbe28930_31);
not \U$5740 ( \5993 , \1094 );
or \U$5741 ( \5994 , \5992 , \5993 );
nand \U$5742 ( \5995 , \1455 , RIbe29560_57);
nand \U$5743 ( \5996 , \5994 , \5995 );
and \U$5744 ( \5997 , \5996 , \1309 );
not \U$5745 ( \5998 , \5996 );
and \U$5746 ( \5999 , \5998 , \1082 );
nor \U$5747 ( \6000 , \5997 , \5999 );
not \U$5748 ( \6001 , \6000 );
nor \U$5749 ( \6002 , \5991 , \6001 );
nor \U$5750 ( \6003 , \5980 , \5990 );
nor \U$5751 ( \6004 , \6002 , \6003 );
not \U$5752 ( \6005 , \6004 );
not \U$5753 ( \6006 , RIbe285e8_24);
not \U$5754 ( \6007 , \383 );
or \U$5755 ( \6008 , \6006 , \6007 );
nand \U$5756 ( \6009 , \429 , RIbe287c8_28);
nand \U$5757 ( \6010 , \6008 , \6009 );
and \U$5758 ( \6011 , \6010 , \313 );
not \U$5759 ( \6012 , \6010 );
and \U$5760 ( \6013 , \6012 , \306 );
nor \U$5761 ( \6014 , \6011 , \6013 );
not \U$5762 ( \6015 , RIbe28480_21);
not \U$5763 ( \6016 , \3244 );
or \U$5764 ( \6017 , \6015 , \6016 );
nand \U$5765 ( \6018 , \1327 , RIbe28408_20);
nand \U$5766 ( \6019 , \6017 , \6018 );
not \U$5767 ( \6020 , \6019 );
not \U$5768 ( \6021 , \424 );
and \U$5769 ( \6022 , \6020 , \6021 );
and \U$5770 ( \6023 , \6019 , \1333 );
nor \U$5771 ( \6024 , \6022 , \6023 );
and \U$5772 ( \6025 , \6014 , \6024 );
not \U$5773 ( \6026 , RIbe28390_19);
not \U$5774 ( \6027 , \664 );
or \U$5775 ( \6028 , \6026 , \6027 );
nand \U$5776 ( \6029 , \1180 , RIbe28b10_35);
nand \U$5777 ( \6030 , \6028 , \6029 );
not \U$5778 ( \6031 , \6030 );
not \U$5779 ( \6032 , \564 );
and \U$5780 ( \6033 , \6031 , \6032 );
and \U$5781 ( \6034 , \6030 , \4217 );
nor \U$5782 ( \6035 , \6033 , \6034 );
nor \U$5783 ( \6036 , \6025 , \6035 );
nor \U$5784 ( \6037 , \6014 , \6024 );
nor \U$5785 ( \6038 , \6036 , \6037 );
not \U$5786 ( \6039 , \6038 );
or \U$5787 ( \6040 , \6005 , \6039 );
not \U$5788 ( \6041 , RIbe28f48_44);
not \U$5789 ( \6042 , \3160 );
or \U$5790 ( \6043 , \6041 , \6042 );
nand \U$5791 ( \6044 , \329 , RIbe28ed0_43);
nand \U$5792 ( \6045 , \6043 , \6044 );
not \U$5793 ( \6046 , \6045 );
not \U$5794 ( \6047 , \4172 );
and \U$5795 ( \6048 , \6046 , \6047 );
and \U$5796 ( \6049 , \6045 , \339 );
nor \U$5797 ( \6050 , \6048 , \6049 );
not \U$5798 ( \6051 , \6050 );
not \U$5799 ( \6052 , RIbe27fd0_11);
not \U$5800 ( \6053 , \261 );
or \U$5801 ( \6054 , \6052 , \6053 );
nand \U$5802 ( \6055 , \263 , RIbe27f58_10);
nand \U$5803 ( \6056 , \6054 , \6055 );
not \U$5804 ( \6057 , \6056 );
not \U$5805 ( \6058 , \268 );
not \U$5806 ( \6059 , \6058 );
and \U$5807 ( \6060 , \6057 , \6059 );
and \U$5808 ( \6061 , \6056 , \1362 );
nor \U$5809 ( \6062 , \6060 , \6061 );
not \U$5810 ( \6063 , \6062 );
or \U$5811 ( \6064 , \6051 , \6063 );
not \U$5812 ( \6065 , RIbe27e68_8);
not \U$5813 ( \6066 , \1528 );
or \U$5814 ( \6067 , \6065 , \6066 );
nand \U$5815 ( \6068 , \287 , RIbe28660_25);
nand \U$5816 ( \6069 , \6067 , \6068 );
xnor \U$5817 ( \6070 , \300 , \6069 );
nand \U$5818 ( \6071 , \6064 , \6070 );
or \U$5819 ( \6072 , \6062 , \6050 );
nand \U$5820 ( \6073 , \6071 , \6072 );
nand \U$5821 ( \6074 , \6040 , \6073 );
not \U$5822 ( \6075 , \6038 );
not \U$5823 ( \6076 , \6004 );
nand \U$5824 ( \6077 , \6075 , \6076 );
and \U$5825 ( \6078 , \6074 , \6077 );
nand \U$5826 ( \6079 , \5972 , \6078 );
not \U$5827 ( \6080 , RIbe290b0_47);
not \U$5828 ( \6081 , \5094 );
or \U$5829 ( \6082 , \6080 , \6081 );
nand \U$5830 ( \6083 , \4333 , RIbe29a88_68);
nand \U$5831 ( \6084 , \6082 , \6083 );
and \U$5832 ( \6085 , \6084 , \3448 );
not \U$5833 ( \6086 , \6084 );
and \U$5834 ( \6087 , \6086 , \3471 );
nor \U$5835 ( \6088 , \6085 , \6087 );
not \U$5836 ( \6089 , RIbe29038_46);
not \U$5837 ( \6090 , \3285 );
or \U$5838 ( \6091 , \6089 , \6090 );
nand \U$5839 ( \6092 , \3458 , RIbe28fc0_45);
nand \U$5840 ( \6093 , \6091 , \6092 );
and \U$5841 ( \6094 , \6093 , \3461 );
not \U$5842 ( \6095 , \6093 );
and \U$5843 ( \6096 , \6095 , \4346 );
nor \U$5844 ( \6097 , \6094 , \6096 );
and \U$5845 ( \6098 , \6088 , \6097 );
not \U$5846 ( \6099 , RIbe27d78_6);
not \U$5847 ( \6100 , \4595 );
or \U$5848 ( \6101 , \6099 , \6100 );
nand \U$5849 ( \6102 , \4600 , RIbe27d00_5);
nand \U$5850 ( \6103 , \6101 , \6102 );
and \U$5851 ( \6104 , \6103 , \4323 );
not \U$5852 ( \6105 , \6103 );
and \U$5853 ( \6106 , \6105 , \4007 );
nor \U$5854 ( \6107 , \6104 , \6106 );
nor \U$5855 ( \6108 , \6098 , \6107 );
nor \U$5856 ( \6109 , \6097 , \6088 );
nor \U$5857 ( \6110 , \6108 , \6109 );
not \U$5858 ( \6111 , \6110 );
not \U$5859 ( \6112 , RIbe28de0_41);
not \U$5860 ( \6113 , \5455 );
or \U$5861 ( \6114 , \6112 , \6113 );
nand \U$5862 ( \6115 , \5751 , RIbe29920_65);
nand \U$5863 ( \6116 , \6114 , \6115 );
buf \U$5864 ( \6117 , \5045 );
not \U$5865 ( \6118 , \6117 );
and \U$5866 ( \6119 , \6116 , \6118 );
not \U$5867 ( \6120 , \6116 );
buf \U$5868 ( \6121 , \5460 );
and \U$5869 ( \6122 , \6120 , \6121 );
nor \U$5870 ( \6123 , \6119 , \6122 );
not \U$5871 ( \6124 , RIbe27c10_3);
not \U$5872 ( \6125 , \4830 );
or \U$5873 ( \6126 , \6124 , \6125 );
nand \U$5874 ( \6127 , \5731 , RIbe28e58_42);
nand \U$5875 ( \6128 , \6126 , \6127 );
and \U$5876 ( \6129 , \6128 , \4592 );
not \U$5877 ( \6130 , \6128 );
and \U$5878 ( \6131 , \6130 , \4586 );
nor \U$5879 ( \6132 , \6129 , \6131 );
nand \U$5880 ( \6133 , \6123 , \6132 );
xor \U$5881 ( \6134 , RIbe29b78_70, RIbe29ce0_73);
xor \U$5882 ( \6135 , RIbe29ce0_73, RIbe29d58_74);
not \U$5883 ( \6136 , \6135 );
and \U$5884 ( \6137 , \6134 , \6136 );
buf \U$5885 ( \6138 , \6137 );
buf \U$5886 ( \6139 , \6138 );
nand \U$5887 ( \6140 , \6139 , RIbe27b98_2);
buf \U$5888 ( \6141 , \5740 );
and \U$5889 ( \6142 , \6140 , \6141 );
not \U$5890 ( \6143 , \6140 );
not \U$5891 ( \6144 , \6141 );
and \U$5892 ( \6145 , \6143 , \6144 );
nor \U$5893 ( \6146 , \6142 , \6145 );
and \U$5894 ( \6147 , \6133 , \6146 );
nor \U$5895 ( \6148 , \6123 , \6132 );
nor \U$5896 ( \6149 , \6147 , \6148 );
not \U$5897 ( \6150 , \6149 );
or \U$5898 ( \6151 , \6111 , \6150 );
not \U$5899 ( \6152 , RIbe296c8_60);
not \U$5900 ( \6153 , \4051 );
or \U$5901 ( \6154 , \6152 , \6153 );
nand \U$5902 ( \6155 , \3267 , RIbe29650_59);
nand \U$5903 ( \6156 , \6154 , \6155 );
and \U$5904 ( \6157 , \6156 , \3481 );
not \U$5905 ( \6158 , \6156 );
and \U$5906 ( \6159 , \6158 , \2576 );
nor \U$5907 ( \6160 , \6157 , \6159 );
and \U$5908 ( \6161 , \1272 , RIbe280c0_13);
and \U$5909 ( \6162 , \2384 , RIbe29830_63);
nor \U$5910 ( \6163 , \6161 , \6162 );
and \U$5911 ( \6164 , \6163 , \1076 );
not \U$5912 ( \6165 , \6163 );
and \U$5913 ( \6166 , \6165 , \1277 );
nor \U$5914 ( \6167 , \6164 , \6166 );
xor \U$5915 ( \6168 , \6160 , \6167 );
and \U$5916 ( \6169 , \1113 , RIbe28228_16);
and \U$5917 ( \6170 , \1117 , RIbe281b0_15);
nor \U$5918 ( \6171 , \6169 , \6170 );
and \U$5919 ( \6172 , \6171 , \1125 );
not \U$5920 ( \6173 , \6171 );
and \U$5921 ( \6174 , \6173 , \1132 );
nor \U$5922 ( \6175 , \6172 , \6174 );
and \U$5923 ( \6176 , \6168 , \6175 );
and \U$5924 ( \6177 , \6160 , \6167 );
or \U$5925 ( \6178 , \6176 , \6177 );
nand \U$5926 ( \6179 , \6151 , \6178 );
not \U$5927 ( \6180 , \6110 );
not \U$5928 ( \6181 , \6149 );
nand \U$5929 ( \6182 , \6180 , \6181 );
nand \U$5930 ( \6183 , \6179 , \6182 );
and \U$5931 ( \6184 , \6079 , \6183 );
nor \U$5932 ( \6185 , \5972 , \6078 );
nor \U$5933 ( \6186 , \6184 , \6185 );
xor \U$5934 ( \6187 , \5800 , \5828 );
xor \U$5935 ( \6188 , \6187 , \5858 );
not \U$5936 ( \6189 , \6188 );
or \U$5937 ( \6190 , \5646 , \5648 );
and \U$5938 ( \6191 , \5649 , \6190 );
and \U$5939 ( \6192 , \6189 , \6191 );
xor \U$5940 ( \6193 , \5723 , \5761 );
xor \U$5941 ( \6194 , \6193 , \5687 );
nor \U$5942 ( \6195 , \6192 , \6194 );
nor \U$5943 ( \6196 , \6189 , \6191 );
nor \U$5944 ( \6197 , \6195 , \6196 );
nand \U$5945 ( \6198 , \6186 , \6197 );
not \U$5946 ( \6199 , \6198 );
xor \U$5947 ( \6200 , \5444 , \5462 );
xor \U$5948 ( \6201 , \5450 , \6200 );
xor \U$5949 ( \6202 , \5838 , \5845 );
xor \U$5950 ( \6203 , \6202 , \5855 );
not \U$5951 ( \6204 , \6203 );
not \U$5952 ( \6205 , \5669 );
not \U$5953 ( \6206 , \5681 );
or \U$5954 ( \6207 , \6205 , \6206 );
nand \U$5955 ( \6208 , \5680 , \5683 );
nand \U$5956 ( \6209 , \6207 , \6208 );
and \U$5957 ( \6210 , \6209 , \5659 );
not \U$5958 ( \6211 , \6209 );
and \U$5959 ( \6212 , \6211 , \5684 );
nor \U$5960 ( \6213 , \6210 , \6212 );
not \U$5961 ( \6214 , \6213 );
not \U$5962 ( \6215 , \6214 );
or \U$5963 ( \6216 , \6204 , \6215 );
not \U$5964 ( \6217 , \5721 );
not \U$5965 ( \6218 , \5697 );
or \U$5966 ( \6219 , \6217 , \6218 );
nand \U$5967 ( \6220 , \5698 , \5720 );
nand \U$5968 ( \6221 , \6219 , \6220 );
and \U$5969 ( \6222 , \6221 , \5706 );
not \U$5970 ( \6223 , \6221 );
and \U$5971 ( \6224 , \6223 , \5707 );
nor \U$5972 ( \6225 , \6222 , \6224 );
not \U$5973 ( \6226 , \6225 );
not \U$5974 ( \6227 , \6203 );
nand \U$5975 ( \6228 , \6227 , \6213 );
nand \U$5976 ( \6229 , \6226 , \6228 );
nand \U$5977 ( \6230 , \6216 , \6229 );
xor \U$5978 ( \6231 , \6201 , \6230 );
and \U$5979 ( \6232 , \5874 , \5887 );
not \U$5980 ( \6233 , \5874 );
and \U$5981 ( \6234 , \6233 , \5888 );
nor \U$5982 ( \6235 , \6232 , \6234 );
and \U$5983 ( \6236 , \6235 , \5870 );
not \U$5984 ( \6237 , \6235 );
and \U$5985 ( \6238 , \6237 , \5871 );
nor \U$5986 ( \6239 , \6236 , \6238 );
and \U$5987 ( \6240 , \6231 , \6239 );
and \U$5988 ( \6241 , \6201 , \6230 );
or \U$5989 ( \6242 , \6240 , \6241 );
not \U$5990 ( \6243 , \6242 );
or \U$5991 ( \6244 , \6199 , \6243 );
not \U$5992 ( \6245 , \6186 );
not \U$5993 ( \6246 , \6197 );
nand \U$5994 ( \6247 , \6245 , \6246 );
nand \U$5995 ( \6248 , \6244 , \6247 );
xnor \U$5996 ( \6249 , \5640 , \5643 );
xor \U$5997 ( \6250 , \5649 , \5766 );
xor \U$5998 ( \6251 , \6250 , \5861 );
xor \U$5999 ( \6252 , \6249 , \6251 );
xor \U$6000 ( \6253 , \5890 , \5892 );
xor \U$6001 ( \6254 , \6253 , \5902 );
and \U$6002 ( \6255 , \6252 , \6254 );
and \U$6003 ( \6256 , \6249 , \6251 );
or \U$6004 ( \6257 , \6255 , \6256 );
xor \U$6005 ( \6258 , \6248 , \6257 );
and \U$6006 ( \6259 , \5912 , \5916 );
not \U$6007 ( \6260 , \5912 );
and \U$6008 ( \6261 , \6260 , \5915 );
nor \U$6009 ( \6262 , \6259 , \6261 );
not \U$6010 ( \6263 , \6262 );
not \U$6011 ( \6264 , \5911 );
or \U$6012 ( \6265 , \6263 , \6264 );
or \U$6013 ( \6266 , \5911 , \6262 );
nand \U$6014 ( \6267 , \6265 , \6266 );
and \U$6015 ( \6268 , \6258 , \6267 );
and \U$6016 ( \6269 , \6248 , \6257 );
or \U$6017 ( \6270 , \6268 , \6269 );
nand \U$6018 ( \6271 , \5951 , \6270 );
nand \U$6019 ( \6272 , \5949 , \6271 );
nand \U$6020 ( \6273 , \5941 , \6272 );
not \U$6021 ( \6274 , \6273 );
xor \U$6022 ( \6275 , \5934 , \5936 );
not \U$6023 ( \6276 , \6275 );
or \U$6024 ( \6277 , \6274 , \6276 );
or \U$6025 ( \6278 , \6275 , \6273 );
nand \U$6026 ( \6279 , \6277 , \6278 );
and \U$6027 ( \6280 , \5340 , \5636 , \5939 , \6279 );
xor \U$6028 ( \6281 , \3861 , \3864 );
xor \U$6029 ( \6282 , \6281 , \4113 );
not \U$6030 ( \6283 , \5323 );
nand \U$6031 ( \6284 , \6283 , \5325 );
and \U$6032 ( \6285 , \6284 , \5332 );
and \U$6033 ( \6286 , \5323 , \5326 );
nor \U$6034 ( \6287 , \6285 , \6286 );
not \U$6035 ( \6288 , \6287 );
xor \U$6036 ( \6289 , \3868 , \3870 );
xor \U$6037 ( \6290 , \6289 , \4110 );
nand \U$6038 ( \6291 , \6288 , \6290 );
xor \U$6039 ( \6292 , \6282 , \6291 );
and \U$6040 ( \6293 , \5319 , \5337 );
xnor \U$6041 ( \6294 , \6287 , \6290 );
xor \U$6042 ( \6295 , \6293 , \6294 );
nand \U$6043 ( \6296 , \6280 , \6292 , \6295 );
nor \U$6044 ( \6297 , \4143 , \6296 );
not \U$6045 ( \6298 , \6297 );
and \U$6046 ( \6299 , RIbe2a2f8_86, RIbe29380_53);
not \U$6047 ( \6300 , RIbe29bf0_71);
not \U$6048 ( \6301 , \1223 );
or \U$6049 ( \6302 , \6300 , \6301 );
nand \U$6050 ( \6303 , \429 , RIbe28f48_44);
nand \U$6051 ( \6304 , \6302 , \6303 );
and \U$6052 ( \6305 , \6304 , \306 );
not \U$6053 ( \6306 , \6304 );
and \U$6054 ( \6307 , \6306 , \1232 );
nor \U$6055 ( \6308 , \6305 , \6307 );
not \U$6056 ( \6309 , \6308 );
not \U$6057 ( \6310 , RIbe29dd0_75);
not \U$6058 ( \6311 , \282 );
not \U$6059 ( \6312 , \6311 );
or \U$6060 ( \6313 , \6310 , \6312 );
nand \U$6061 ( \6314 , \1256 , RIbe29c68_72);
nand \U$6062 ( \6315 , \6313 , \6314 );
and \U$6063 ( \6316 , \6315 , \300 );
not \U$6064 ( \6317 , \6315 );
and \U$6065 ( \6318 , \6317 , \293 );
nor \U$6066 ( \6319 , \6316 , \6318 );
not \U$6067 ( \6320 , \6319 );
or \U$6068 ( \6321 , \6309 , \6320 );
or \U$6069 ( \6322 , \6308 , \6319 );
nand \U$6070 ( \6323 , \6321 , \6322 );
and \U$6071 ( \6324 , \1659 , RIbe29fb0_79);
buf \U$6072 ( \6325 , \263 );
and \U$6073 ( \6326 , \6325 , RIbe29e48_76);
nor \U$6074 ( \6327 , \6324 , \6326 );
and \U$6075 ( \6328 , \6327 , \269 );
not \U$6076 ( \6329 , \6327 );
and \U$6077 ( \6330 , \6329 , \1362 );
nor \U$6078 ( \6331 , \6328 , \6330 );
xnor \U$6079 ( \6332 , \6323 , \6331 );
xor \U$6080 ( \6333 , \6299 , \6332 );
not \U$6081 ( \6334 , RIbe28ed0_43);
not \U$6082 ( \6335 , \548 );
or \U$6083 ( \6336 , \6334 , \6335 );
nand \U$6084 ( \6337 , \1327 , RIbe27fd0_11);
nand \U$6085 ( \6338 , \6336 , \6337 );
not \U$6086 ( \6339 , \6338 );
not \U$6087 ( \6340 , \3415 );
not \U$6088 ( \6341 , \6340 );
and \U$6089 ( \6342 , \6339 , \6341 );
and \U$6090 ( \6343 , \6338 , \424 );
nor \U$6091 ( \6344 , \6342 , \6343 );
not \U$6092 ( \6345 , \1179 );
not \U$6093 ( \6346 , \6345 );
not \U$6094 ( \6347 , RIbe27e68_8);
not \U$6095 ( \6348 , \6347 );
and \U$6096 ( \6349 , \6346 , \6348 );
not \U$6097 ( \6350 , \1743 );
and \U$6098 ( \6351 , \6350 , RIbe27f58_10);
nor \U$6099 ( \6352 , \6349 , \6351 );
and \U$6100 ( \6353 , \6352 , \1618 );
not \U$6101 ( \6354 , \6352 );
and \U$6102 ( \6355 , \6354 , \1621 );
nor \U$6103 ( \6356 , \6353 , \6355 );
xor \U$6104 ( \6357 , \6344 , \6356 );
and \U$6105 ( \6358 , \1807 , RIbe28660_25);
and \U$6106 ( \6359 , \2000 , RIbe285e8_24);
nor \U$6107 ( \6360 , \6358 , \6359 );
and \U$6108 ( \6361 , \6360 , \1011 );
not \U$6109 ( \6362 , \6360 );
and \U$6110 ( \6363 , \6362 , \1813 );
nor \U$6111 ( \6364 , \6361 , \6363 );
xor \U$6112 ( \6365 , \6357 , \6364 );
and \U$6113 ( \6366 , \6333 , \6365 );
and \U$6114 ( \6367 , \6299 , \6332 );
or \U$6115 ( \6368 , \6366 , \6367 );
not \U$6116 ( \6369 , RIbe28408_20);
not \U$6117 ( \6370 , \1633 );
or \U$6118 ( \6371 , \6369 , \6370 );
nand \U$6119 ( \6372 , \4730 , RIbe28390_19);
nand \U$6120 ( \6373 , \6371 , \6372 );
and \U$6121 ( \6374 , \6373 , \5125 );
not \U$6122 ( \6375 , \6373 );
and \U$6123 ( \6376 , \6375 , \1309 );
nor \U$6124 ( \6377 , \6374 , \6376 );
not \U$6125 ( \6378 , \6377 );
not \U$6126 ( \6379 , \6378 );
not \U$6127 ( \6380 , \1284 );
and \U$6128 ( \6381 , \6380 , RIbe28b10_35);
buf \U$6129 ( \6382 , \1115 );
not \U$6130 ( \6383 , \6382 );
and \U$6131 ( \6384 , \6383 , RIbe28b88_36);
nor \U$6132 ( \6385 , \6381 , \6384 );
and \U$6133 ( \6386 , \6385 , \3491 );
not \U$6134 ( \6387 , \6385 );
and \U$6135 ( \6388 , \6387 , \1131 );
nor \U$6136 ( \6389 , \6386 , \6388 );
not \U$6137 ( \6390 , \6389 );
not \U$6138 ( \6391 , \6390 );
or \U$6139 ( \6392 , \6379 , \6391 );
nand \U$6140 ( \6393 , \6389 , \6377 );
nand \U$6141 ( \6394 , \6392 , \6393 );
not \U$6142 ( \6395 , RIbe287c8_28);
not \U$6143 ( \6396 , \1143 );
or \U$6144 ( \6397 , \6395 , \6396 );
nand \U$6145 ( \6398 , \1147 , RIbe28480_21);
nand \U$6146 ( \6399 , \6397 , \6398 );
and \U$6147 ( \6400 , \6399 , \1469 );
not \U$6148 ( \6401 , \6399 );
and \U$6149 ( \6402 , \6401 , \1153 );
nor \U$6150 ( \6403 , \6400 , \6402 );
not \U$6151 ( \6404 , \6403 );
and \U$6152 ( \6405 , \6394 , \6404 );
not \U$6153 ( \6406 , \6394 );
and \U$6154 ( \6407 , \6406 , \6403 );
nor \U$6155 ( \6408 , \6405 , \6407 );
not \U$6156 ( \6409 , \6408 );
not \U$6157 ( \6410 , \6409 );
not \U$6158 ( \6411 , \4323 );
not \U$6159 ( \6412 , RIbe29830_63);
not \U$6160 ( \6413 , \4316 );
buf \U$6161 ( \6414 , \6413 );
not \U$6162 ( \6415 , \6414 );
or \U$6163 ( \6416 , \6412 , \6415 );
not \U$6164 ( \6417 , \4599 );
not \U$6165 ( \6418 , \6417 );
nand \U$6166 ( \6419 , \6418 , RIbe296c8_60);
nand \U$6167 ( \6420 , \6416 , \6419 );
not \U$6168 ( \6421 , \6420 );
or \U$6169 ( \6422 , \6411 , \6421 );
or \U$6170 ( \6423 , \6420 , \4323 );
nand \U$6171 ( \6424 , \6422 , \6423 );
not \U$6172 ( \6425 , \6424 );
not \U$6173 ( \6426 , RIbe29650_59);
not \U$6174 ( \6427 , \4828 );
not \U$6175 ( \6428 , \6427 );
or \U$6176 ( \6429 , \6426 , \6428 );
nand \U$6177 ( \6430 , \5052 , RIbe29038_46);
nand \U$6178 ( \6431 , \6429 , \6430 );
and \U$6179 ( \6432 , \6431 , \4592 );
not \U$6180 ( \6433 , \6431 );
and \U$6181 ( \6434 , \6433 , \4586 );
nor \U$6182 ( \6435 , \6432 , \6434 );
not \U$6183 ( \6436 , \6435 );
or \U$6184 ( \6437 , \6425 , \6436 );
or \U$6185 ( \6438 , \6435 , \6424 );
nand \U$6186 ( \6439 , \6437 , \6438 );
not \U$6187 ( \6440 , RIbe281b0_15);
not \U$6188 ( \6441 , \4021 );
or \U$6189 ( \6442 , \6440 , \6441 );
nand \U$6190 ( \6443 , \4333 , RIbe280c0_13);
nand \U$6191 ( \6444 , \6442 , \6443 );
and \U$6192 ( \6445 , \6444 , \3698 );
not \U$6193 ( \6446 , \6444 );
and \U$6194 ( \6447 , \6446 , \3471 );
nor \U$6195 ( \6448 , \6445 , \6447 );
xnor \U$6196 ( \6449 , \6439 , \6448 );
not \U$6197 ( \6450 , \6449 );
or \U$6198 ( \6451 , \6410 , \6450 );
not \U$6199 ( \6452 , RIbe29560_57);
not \U$6200 ( \6453 , \3452 );
or \U$6201 ( \6454 , \6452 , \6453 );
nand \U$6202 ( \6455 , \3458 , RIbe28228_16);
nand \U$6203 ( \6456 , \6454 , \6455 );
and \U$6204 ( \6457 , \6456 , \2887 );
not \U$6205 ( \6458 , \6456 );
and \U$6206 ( \6459 , \6458 , \3290 );
nor \U$6207 ( \6460 , \6457 , \6459 );
not \U$6208 ( \6461 , RIbe289a8_32);
not \U$6209 ( \6462 , \4051 );
or \U$6210 ( \6463 , \6461 , \6462 );
nand \U$6211 ( \6464 , \3267 , RIbe28930_31);
nand \U$6212 ( \6465 , \6463 , \6464 );
and \U$6213 ( \6466 , \6465 , \4287 );
not \U$6214 ( \6467 , \6465 );
not \U$6215 ( \6468 , \4287 );
and \U$6216 ( \6469 , \6467 , \6468 );
nor \U$6217 ( \6470 , \6466 , \6469 );
and \U$6218 ( \6471 , \6460 , \6470 );
not \U$6219 ( \6472 , \6460 );
not \U$6220 ( \6473 , \6470 );
and \U$6221 ( \6474 , \6472 , \6473 );
or \U$6222 ( \6475 , \6471 , \6474 );
not \U$6223 ( \6476 , RIbe29290_51);
not \U$6224 ( \6477 , \3303 );
or \U$6225 ( \6478 , \6476 , \6477 );
not \U$6226 ( \6479 , \4065 );
nand \U$6227 ( \6480 , \6479 , RIbe28a20_33);
nand \U$6228 ( \6481 , \6478 , \6480 );
xnor \U$6229 ( \6482 , \6481 , \1076 );
xnor \U$6230 ( \6483 , \6475 , \6482 );
not \U$6231 ( \6484 , \6483 );
not \U$6232 ( \6485 , \6449 );
nand \U$6233 ( \6486 , \6485 , \6408 );
nand \U$6234 ( \6487 , \6484 , \6486 );
nand \U$6235 ( \6488 , \6451 , \6487 );
xor \U$6236 ( \6489 , \6368 , \6488 );
not \U$6237 ( \6490 , RIbe280c0_13);
not \U$6238 ( \6491 , \4021 );
or \U$6239 ( \6492 , \6490 , \6491 );
nand \U$6240 ( \6493 , \4027 , RIbe29830_63);
nand \U$6241 ( \6494 , \6492 , \6493 );
and \U$6242 ( \6495 , \6494 , \3471 );
not \U$6243 ( \6496 , \6494 );
and \U$6244 ( \6497 , \6496 , \4821 );
nor \U$6245 ( \6498 , \6495 , \6497 );
not \U$6246 ( \6499 , \6498 );
not \U$6247 ( \6500 , \6499 );
not \U$6248 ( \6501 , RIbe296c8_60);
not \U$6249 ( \6502 , \5058 );
or \U$6250 ( \6503 , \6501 , \6502 );
nand \U$6251 ( \6504 , \4600 , RIbe29650_59);
nand \U$6252 ( \6505 , \6503 , \6504 );
and \U$6253 ( \6506 , \6505 , \4323 );
not \U$6254 ( \6507 , \6505 );
and \U$6255 ( \6508 , \6507 , \4326 );
nor \U$6256 ( \6509 , \6506 , \6508 );
not \U$6257 ( \6510 , \6509 );
not \U$6258 ( \6511 , \6510 );
or \U$6259 ( \6512 , \6500 , \6511 );
nand \U$6260 ( \6513 , \6509 , \6498 );
nand \U$6261 ( \6514 , \6512 , \6513 );
not \U$6262 ( \6515 , RIbe28228_16);
not \U$6263 ( \6516 , \3285 );
or \U$6264 ( \6517 , \6515 , \6516 );
nand \U$6265 ( \6518 , \3458 , RIbe281b0_15);
nand \U$6266 ( \6519 , \6517 , \6518 );
and \U$6267 ( \6520 , \6519 , \3290 );
not \U$6268 ( \6521 , \6519 );
and \U$6269 ( \6522 , \6521 , \3461 );
nor \U$6270 ( \6523 , \6520 , \6522 );
not \U$6271 ( \6524 , \6523 );
and \U$6272 ( \6525 , \6514 , \6524 );
not \U$6273 ( \6526 , \6514 );
and \U$6274 ( \6527 , \6526 , \6523 );
nor \U$6275 ( \6528 , \6525 , \6527 );
not \U$6276 ( \6529 , RIbe29f38_78);
not \U$6277 ( \6530 , RIbe29ec0_77);
nand \U$6278 ( \6531 , \6529 , \6530 , RIbe29d58_74);
not \U$6279 ( \6532 , RIbe29d58_74);
nand \U$6280 ( \6533 , \6532 , RIbe29f38_78, RIbe29ec0_77);
nand \U$6281 ( \6534 , \6531 , \6533 );
buf \U$6282 ( \6535 , \6534 );
buf \U$6283 ( \6536 , \6535 );
buf \U$6284 ( \6537 , \6536 );
and \U$6285 ( \6538 , \6537 , RIbe27c10_3);
xor \U$6286 ( \6539 , RIbe29ec0_77, RIbe29f38_78);
buf \U$6287 ( \6540 , \6539 );
not \U$6288 ( \6541 , \6540 );
nor \U$6289 ( \6542 , \6541 , \3299 );
nor \U$6290 ( \6543 , \6538 , \6542 );
nand \U$6291 ( \6544 , RIbe29ec0_77, RIbe29f38_78);
nand \U$6292 ( \6545 , \6544 , RIbe29d58_74);
not \U$6293 ( \6546 , \6545 );
buf \U$6294 ( \6547 , \6546 );
not \U$6295 ( \6548 , \6547 );
and \U$6296 ( \6549 , \6543 , \6548 );
not \U$6297 ( \6550 , \6543 );
not \U$6298 ( \6551 , \6546 );
not \U$6299 ( \6552 , \6551 );
and \U$6300 ( \6553 , \6550 , \6552 );
nor \U$6301 ( \6554 , \6549 , \6553 );
xor \U$6302 ( \6555 , RIbe2aa00_101, RIbe2a898_98);
not \U$6303 ( \6556 , \6555 );
xor \U$6304 ( \6557 , RIbe2aa78_102, RIbe2aa00_101);
nand \U$6305 ( \6558 , \6556 , \6557 );
buf \U$6306 ( \6559 , \6558 );
not \U$6307 ( \6560 , \6559 );
buf \U$6308 ( \6561 , \6560 );
not \U$6309 ( \6562 , \6561 );
nor \U$6310 ( \6563 , \6562 , \1640 );
not \U$6311 ( \6564 , \6563 );
not \U$6312 ( \6565 , RIbe2aa00_101);
not \U$6313 ( \6566 , RIbe2a898_98);
or \U$6314 ( \6567 , \6565 , \6566 );
nand \U$6315 ( \6568 , \6567 , RIbe2aa78_102);
buf \U$6316 ( \6569 , \6568 );
not \U$6317 ( \6570 , \6569 );
and \U$6318 ( \6571 , \6564 , \6570 );
buf \U$6319 ( \6572 , \6568 );
and \U$6320 ( \6573 , \6563 , \6572 );
nor \U$6321 ( \6574 , \6571 , \6573 );
and \U$6322 ( \6575 , \6554 , \6574 );
not \U$6323 ( \6576 , \6554 );
not \U$6324 ( \6577 , \6574 );
and \U$6325 ( \6578 , \6576 , \6577 );
or \U$6326 ( \6579 , \6575 , \6578 );
nand \U$6327 ( \6580 , RIbe2b6a8_128, RIbe2aa78_102);
and \U$6328 ( \6581 , \6580 , RIbe29f38_78);
buf \U$6329 ( \6582 , \6581 );
not \U$6330 ( \6583 , \6582 );
not \U$6331 ( \6584 , \6583 );
not \U$6332 ( \6585 , RIbe28de0_41);
xor \U$6333 ( \6586 , RIbe2b6a8_128, RIbe2aa78_102);
not \U$6334 ( \6587 , \6586 );
xor \U$6335 ( \6588 , RIbe29f38_78, RIbe2b6a8_128);
nand \U$6336 ( \6589 , \6587 , \6588 );
buf \U$6337 ( \6590 , \6589 );
not \U$6338 ( \6591 , \6590 );
buf \U$6339 ( \6592 , \6591 );
not \U$6340 ( \6593 , \6592 );
or \U$6341 ( \6594 , \6585 , \6593 );
not \U$6342 ( \6595 , \6587 );
buf \U$6343 ( \6596 , \6595 );
nand \U$6344 ( \6597 , \6596 , RIbe29920_65);
nand \U$6345 ( \6598 , \6594 , \6597 );
not \U$6346 ( \6599 , \6598 );
or \U$6347 ( \6600 , \6584 , \6599 );
buf \U$6348 ( \6601 , \6581 );
not \U$6349 ( \6602 , \6601 );
or \U$6350 ( \6603 , \6598 , \6602 );
nand \U$6351 ( \6604 , \6600 , \6603 );
xnor \U$6352 ( \6605 , \6579 , \6604 );
not \U$6353 ( \6606 , \6605 );
and \U$6354 ( \6607 , \6528 , \6606 );
not \U$6355 ( \6608 , \6528 );
and \U$6356 ( \6609 , \6608 , \6605 );
nor \U$6357 ( \6610 , \6607 , \6609 );
not \U$6358 ( \6611 , RIbe27d78_6);
not \U$6359 ( \6612 , \6139 );
or \U$6360 ( \6613 , \6611 , \6612 );
not \U$6361 ( \6614 , \6135 );
buf \U$6362 ( \6615 , \6614 );
not \U$6363 ( \6616 , \6615 );
buf \U$6364 ( \6617 , \6616 );
nand \U$6365 ( \6618 , \6617 , RIbe27d00_5);
nand \U$6366 ( \6619 , \6613 , \6618 );
not \U$6367 ( \6620 , \5740 );
and \U$6368 ( \6621 , \6619 , \6620 );
not \U$6369 ( \6622 , \6619 );
not \U$6370 ( \6623 , \5740 );
not \U$6371 ( \6624 , \6623 );
and \U$6372 ( \6625 , \6622 , \6624 );
nor \U$6373 ( \6626 , \6621 , \6625 );
not \U$6374 ( \6627 , RIbe290b0_47);
not \U$6375 ( \6628 , \5746 );
nand \U$6376 ( \6629 , \6628 , \5453 );
not \U$6377 ( \6630 , \6629 );
not \U$6378 ( \6631 , \6630 );
or \U$6379 ( \6632 , \6627 , \6631 );
not \U$6380 ( \6633 , \5747 );
buf \U$6381 ( \6634 , \6633 );
nand \U$6382 ( \6635 , \6634 , RIbe29a88_68);
nand \U$6383 ( \6636 , \6632 , \6635 );
not \U$6384 ( \6637 , \6117 );
and \U$6385 ( \6638 , \6636 , \6637 );
not \U$6386 ( \6639 , \6636 );
buf \U$6387 ( \6640 , \5044 );
buf \U$6388 ( \6641 , \6640 );
not \U$6389 ( \6642 , \6641 );
and \U$6390 ( \6643 , \6639 , \6642 );
nor \U$6391 ( \6644 , \6638 , \6643 );
and \U$6392 ( \6645 , \6626 , \6644 );
not \U$6393 ( \6646 , \6626 );
not \U$6394 ( \6647 , \6644 );
and \U$6395 ( \6648 , \6646 , \6647 );
or \U$6396 ( \6649 , \6645 , \6648 );
not \U$6397 ( \6650 , RIbe29038_46);
nor \U$6398 ( \6651 , \6650 , \4831 );
and \U$6399 ( \6652 , \5731 , RIbe28fc0_45);
nor \U$6400 ( \6653 , \6651 , \6652 );
xnor \U$6401 ( \6654 , \4586 , \6653 );
not \U$6402 ( \6655 , \6654 );
and \U$6403 ( \6656 , \6649 , \6655 );
not \U$6404 ( \6657 , \6649 );
and \U$6405 ( \6658 , \6657 , \6654 );
nor \U$6406 ( \6659 , \6656 , \6658 );
xor \U$6407 ( \6660 , \6610 , \6659 );
xor \U$6408 ( \6661 , \6489 , \6660 );
nand \U$6409 ( \6662 , RIbe29380_53, RIbe2b5b8_126);
not \U$6410 ( \6663 , RIbe2a3e8_88);
not \U$6411 ( \6664 , \325 );
or \U$6412 ( \6665 , \6663 , \6664 );
nand \U$6413 ( \6666 , \330 , RIbe2a370_87);
nand \U$6414 ( \6667 , \6665 , \6666 );
xnor \U$6415 ( \6668 , \6667 , \1375 );
xor \U$6416 ( \6669 , \6662 , \6668 );
and \U$6417 ( \6670 , \260 , RIbe2a2f8_86);
and \U$6418 ( \6671 , \264 , RIbe2acd0_107);
nor \U$6419 ( \6672 , \6670 , \6671 );
and \U$6420 ( \6673 , \6672 , \270 );
not \U$6421 ( \6674 , \6672 );
and \U$6422 ( \6675 , \6674 , \1663 );
or \U$6423 ( \6676 , \6673 , \6675 );
and \U$6424 ( \6677 , \6669 , \6676 );
and \U$6425 ( \6678 , \6662 , \6668 );
or \U$6426 ( \6679 , \6677 , \6678 );
not \U$6427 ( \6680 , \6679 );
not \U$6428 ( \6681 , \6680 );
and \U$6429 ( \6682 , \1756 , RIbe29c68_72);
and \U$6430 ( \6683 , \1327 , RIbe29bf0_71);
nor \U$6431 ( \6684 , \6682 , \6683 );
and \U$6432 ( \6685 , \6684 , \3415 );
not \U$6433 ( \6686 , \6684 );
and \U$6434 ( \6687 , \6686 , \424 );
nor \U$6435 ( \6688 , \6685 , \6687 );
and \U$6436 ( \6689 , \1528 , RIbe2a028_80);
and \U$6437 ( \6690 , \1531 , RIbe29fb0_79);
nor \U$6438 ( \6691 , \6689 , \6690 );
and \U$6439 ( \6692 , \6691 , \293 );
not \U$6440 ( \6693 , \6691 );
and \U$6441 ( \6694 , \6693 , \300 );
nor \U$6442 ( \6695 , \6692 , \6694 );
nand \U$6443 ( \6696 , \6688 , \6695 );
not \U$6444 ( \6697 , RIbe29e48_76);
not \U$6445 ( \6698 , \1774 );
or \U$6446 ( \6699 , \6697 , \6698 );
nand \U$6447 ( \6700 , \429 , RIbe29dd0_75);
nand \U$6448 ( \6701 , \6699 , \6700 );
and \U$6449 ( \6702 , \6701 , \1232 );
not \U$6450 ( \6703 , \6701 );
and \U$6451 ( \6704 , \6703 , \306 );
nor \U$6452 ( \6705 , \6702 , \6704 );
not \U$6453 ( \6706 , \6705 );
and \U$6454 ( \6707 , \6696 , \6706 );
nor \U$6455 ( \6708 , \6695 , \6688 );
nor \U$6456 ( \6709 , \6707 , \6708 );
not \U$6457 ( \6710 , \6709 );
not \U$6458 ( \6711 , \6710 );
or \U$6459 ( \6712 , \6681 , \6711 );
not \U$6460 ( \6713 , \6709 );
not \U$6461 ( \6714 , \6679 );
or \U$6462 ( \6715 , \6713 , \6714 );
nand \U$6463 ( \6716 , RIbe29380_53, RIbe2a3e8_88);
not \U$6464 ( \6717 , RIbe2a370_87);
not \U$6465 ( \6718 , \324 );
or \U$6466 ( \6719 , \6717 , \6718 );
nand \U$6467 ( \6720 , \329 , RIbe2a2f8_86);
nand \U$6468 ( \6721 , \6719 , \6720 );
xor \U$6469 ( \6722 , \6721 , \5151 );
not \U$6470 ( \6723 , \6722 );
xor \U$6471 ( \6724 , \6716 , \6723 );
not \U$6472 ( \6725 , \6058 );
not \U$6473 ( \6726 , RIbe2acd0_107);
not \U$6474 ( \6727 , \1516 );
or \U$6475 ( \6728 , \6726 , \6727 );
nand \U$6476 ( \6729 , \264 , RIbe2a028_80);
nand \U$6477 ( \6730 , \6728 , \6729 );
not \U$6478 ( \6731 , \6730 );
or \U$6479 ( \6732 , \6725 , \6731 );
or \U$6480 ( \6733 , \6730 , \270 );
nand \U$6481 ( \6734 , \6732 , \6733 );
xnor \U$6482 ( \6735 , \6724 , \6734 );
nand \U$6483 ( \6736 , \6715 , \6735 );
nand \U$6484 ( \6737 , \6712 , \6736 );
not \U$6485 ( \6738 , RIbe27e68_8);
not \U$6486 ( \6739 , \1143 );
or \U$6487 ( \6740 , \6738 , \6739 );
nand \U$6488 ( \6741 , \1147 , RIbe28660_25);
nand \U$6489 ( \6742 , \6740 , \6741 );
and \U$6490 ( \6743 , \6742 , \1152 );
not \U$6491 ( \6744 , \6742 );
and \U$6492 ( \6745 , \6744 , \1652 );
nor \U$6493 ( \6746 , \6743 , \6745 );
not \U$6494 ( \6747 , \1001 );
and \U$6495 ( \6748 , \6747 , RIbe27fd0_11);
and \U$6496 ( \6749 , \2000 , RIbe27f58_10);
nor \U$6497 ( \6750 , \6748 , \6749 );
and \U$6498 ( \6751 , \6750 , \1011 );
not \U$6499 ( \6752 , \6750 );
and \U$6500 ( \6753 , \6752 , \752 );
nor \U$6501 ( \6754 , \6751 , \6753 );
nand \U$6502 ( \6755 , \6746 , \6754 );
not \U$6503 ( \6756 , \1611 );
not \U$6504 ( \6757 , RIbe28ed0_43);
not \U$6505 ( \6758 , \6757 );
and \U$6506 ( \6759 , \6756 , \6758 );
buf \U$6507 ( \6760 , \664 );
and \U$6508 ( \6761 , \6760 , RIbe28f48_44);
nor \U$6509 ( \6762 , \6759 , \6761 );
and \U$6510 ( \6763 , \6762 , \3959 );
not \U$6511 ( \6764 , \6762 );
and \U$6512 ( \6765 , \6764 , \4217 );
nor \U$6513 ( \6766 , \6763 , \6765 );
not \U$6514 ( \6767 , \6766 );
and \U$6515 ( \6768 , \6755 , \6767 );
nor \U$6516 ( \6769 , \6746 , \6754 );
nor \U$6517 ( \6770 , \6768 , \6769 );
not \U$6518 ( \6771 , \6770 );
not \U$6519 ( \6772 , \6771 );
not \U$6520 ( \6773 , RIbe28b88_36);
not \U$6521 ( \6774 , \3476 );
or \U$6522 ( \6775 , \6773 , \6774 );
nand \U$6523 ( \6776 , \4284 , RIbe29290_51);
nand \U$6524 ( \6777 , \6775 , \6776 );
and \U$6525 ( \6778 , \6777 , \3275 );
not \U$6526 ( \6779 , \6777 );
and \U$6527 ( \6780 , \6779 , \4287 );
nor \U$6528 ( \6781 , \6778 , \6780 );
not \U$6529 ( \6782 , RIbe28930_31);
not \U$6530 ( \6783 , \3703 );
not \U$6531 ( \6784 , \6783 );
or \U$6532 ( \6785 , \6782 , \6784 );
not \U$6533 ( \6786 , \4024 );
not \U$6534 ( \6787 , \6786 );
nand \U$6535 ( \6788 , \6787 , RIbe29560_57);
nand \U$6536 ( \6789 , \6785 , \6788 );
and \U$6537 ( \6790 , \6789 , \3471 );
not \U$6538 ( \6791 , \6789 );
and \U$6539 ( \6792 , \6791 , \3698 );
nor \U$6540 ( \6793 , \6790 , \6792 );
not \U$6541 ( \6794 , \6793 );
nand \U$6542 ( \6795 , \6781 , \6794 );
not \U$6543 ( \6796 , RIbe28a20_33);
not \U$6544 ( \6797 , \3282 );
not \U$6545 ( \6798 , \6797 );
or \U$6546 ( \6799 , \6796 , \6798 );
not \U$6547 ( \6800 , \3455 );
nand \U$6548 ( \6801 , \6800 , RIbe289a8_32);
nand \U$6549 ( \6802 , \6799 , \6801 );
and \U$6550 ( \6803 , \6802 , \2887 );
not \U$6551 ( \6804 , \6802 );
and \U$6552 ( \6805 , \6804 , \3290 );
nor \U$6553 ( \6806 , \6803 , \6805 );
not \U$6554 ( \6807 , \6806 );
and \U$6555 ( \6808 , \6795 , \6807 );
nor \U$6556 ( \6809 , \6781 , \6794 );
nor \U$6557 ( \6810 , \6808 , \6809 );
not \U$6558 ( \6811 , \6810 );
not \U$6559 ( \6812 , \6811 );
or \U$6560 ( \6813 , \6772 , \6812 );
not \U$6561 ( \6814 , \6770 );
not \U$6562 ( \6815 , \6810 );
or \U$6563 ( \6816 , \6814 , \6815 );
not \U$6564 ( \6817 , RIbe28390_19);
not \U$6565 ( \6818 , \4295 );
or \U$6566 ( \6819 , \6817 , \6818 );
nand \U$6567 ( \6820 , \2384 , RIbe28b10_35);
nand \U$6568 ( \6821 , \6819 , \6820 );
not \U$6569 ( \6822 , \6821 );
not \U$6570 ( \6823 , \3516 );
and \U$6571 ( \6824 , \6822 , \6823 );
and \U$6572 ( \6825 , \6821 , \1076 );
nor \U$6573 ( \6826 , \6824 , \6825 );
not \U$6574 ( \6827 , \6826 );
and \U$6575 ( \6828 , \2554 , RIbe28480_21);
and \U$6576 ( \6829 , \5467 , RIbe28408_20);
nor \U$6577 ( \6830 , \6828 , \6829 );
not \U$6578 ( \6831 , \1124 );
and \U$6579 ( \6832 , \6830 , \6831 );
not \U$6580 ( \6833 , \6830 );
and \U$6581 ( \6834 , \6833 , \1131 );
nor \U$6582 ( \6835 , \6832 , \6834 );
not \U$6583 ( \6836 , \6835 );
not \U$6584 ( \6837 , RIbe285e8_24);
not \U$6585 ( \6838 , \5476 );
or \U$6586 ( \6839 , \6837 , \6838 );
nand \U$6587 ( \6840 , \2817 , RIbe287c8_28);
nand \U$6588 ( \6841 , \6839 , \6840 );
and \U$6589 ( \6842 , \6841 , \2418 );
not \U$6590 ( \6843 , \6841 );
and \U$6591 ( \6844 , \6843 , \1309 );
nor \U$6592 ( \6845 , \6842 , \6844 );
nand \U$6593 ( \6846 , \6836 , \6845 );
nand \U$6594 ( \6847 , \6827 , \6846 );
not \U$6595 ( \6848 , \6845 );
nand \U$6596 ( \6849 , \6848 , \6835 );
nand \U$6597 ( \6850 , \6847 , \6849 );
nand \U$6598 ( \6851 , \6816 , \6850 );
nand \U$6599 ( \6852 , \6813 , \6851 );
or \U$6600 ( \6853 , \6737 , \6852 );
not \U$6601 ( \6854 , RIbe29038_46);
not \U$6602 ( \6855 , \6137 );
not \U$6603 ( \6856 , \6855 );
not \U$6604 ( \6857 , \6856 );
or \U$6605 ( \6858 , \6854 , \6857 );
not \U$6606 ( \6859 , \6615 );
nand \U$6607 ( \6860 , \6859 , RIbe28fc0_45);
nand \U$6608 ( \6861 , \6858 , \6860 );
not \U$6609 ( \6862 , \6861 );
not \U$6610 ( \6863 , \6624 );
and \U$6611 ( \6864 , \6862 , \6863 );
and \U$6612 ( \6865 , \6861 , \5740 );
nor \U$6613 ( \6866 , \6864 , \6865 );
not \U$6614 ( \6867 , RIbe27d78_6);
not \U$6615 ( \6868 , \6590 );
not \U$6616 ( \6869 , \6868 );
or \U$6617 ( \6870 , \6867 , \6869 );
nand \U$6618 ( \6871 , \6596 , RIbe27d00_5);
nand \U$6619 ( \6872 , \6870 , \6871 );
not \U$6620 ( \6873 , \6601 );
and \U$6621 ( \6874 , \6872 , \6873 );
not \U$6622 ( \6875 , \6872 );
and \U$6623 ( \6876 , \6875 , \6601 );
nor \U$6624 ( \6877 , \6874 , \6876 );
nand \U$6625 ( \6878 , \6866 , \6877 );
not \U$6626 ( \6879 , RIbe290b0_47);
buf \U$6627 ( \6880 , \6535 );
not \U$6628 ( \6881 , \6880 );
or \U$6629 ( \6882 , \6879 , \6881 );
not \U$6630 ( \6883 , \6539 );
not \U$6631 ( \6884 , \6883 );
nand \U$6632 ( \6885 , \6884 , RIbe29a88_68);
nand \U$6633 ( \6886 , \6882 , \6885 );
not \U$6634 ( \6887 , \6886 );
not \U$6635 ( \6888 , \6546 );
not \U$6636 ( \6889 , \6888 );
and \U$6637 ( \6890 , \6887 , \6889 );
buf \U$6638 ( \6891 , \6545 );
and \U$6639 ( \6892 , \6886 , \6891 );
nor \U$6640 ( \6893 , \6890 , \6892 );
not \U$6641 ( \6894 , \6893 );
and \U$6642 ( \6895 , \6878 , \6894 );
nor \U$6643 ( \6896 , \6877 , \6866 );
nor \U$6644 ( \6897 , \6895 , \6896 );
not \U$6645 ( \6898 , \6897 );
not \U$6646 ( \6899 , \6898 );
not \U$6647 ( \6900 , RIbe296c8_60);
not \U$6648 ( \6901 , \5455 );
or \U$6649 ( \6902 , \6900 , \6901 );
nand \U$6650 ( \6903 , \6634 , RIbe29650_59);
nand \U$6651 ( \6904 , \6902 , \6903 );
and \U$6652 ( \6905 , \6904 , \5754 );
not \U$6653 ( \6906 , \6904 );
not \U$6654 ( \6907 , \5457 );
and \U$6655 ( \6908 , \6906 , \6907 );
nor \U$6656 ( \6909 , \6905 , \6908 );
not \U$6657 ( \6910 , RIbe28228_16);
not \U$6658 ( \6911 , \4317 );
or \U$6659 ( \6912 , \6910 , \6911 );
nand \U$6660 ( \6913 , \4600 , RIbe281b0_15);
nand \U$6661 ( \6914 , \6912 , \6913 );
and \U$6662 ( \6915 , \6914 , \4323 );
not \U$6663 ( \6916 , \6914 );
and \U$6664 ( \6917 , \6916 , \4007 );
nor \U$6665 ( \6918 , \6915 , \6917 );
nand \U$6666 ( \6919 , \6909 , \6918 );
not \U$6667 ( \6920 , \4592 );
not \U$6668 ( \6921 , RIbe280c0_13);
not \U$6669 ( \6922 , \5727 );
or \U$6670 ( \6923 , \6921 , \6922 );
nand \U$6671 ( \6924 , \5731 , RIbe29830_63);
nand \U$6672 ( \6925 , \6923 , \6924 );
not \U$6673 ( \6926 , \6925 );
or \U$6674 ( \6927 , \6920 , \6926 );
or \U$6675 ( \6928 , \6925 , \4592 );
nand \U$6676 ( \6929 , \6927 , \6928 );
and \U$6677 ( \6930 , \6919 , \6929 );
nor \U$6678 ( \6931 , \6909 , \6918 );
nor \U$6679 ( \6932 , \6930 , \6931 );
not \U$6680 ( \6933 , \6932 );
not \U$6681 ( \6934 , \6933 );
or \U$6682 ( \6935 , \6899 , \6934 );
not \U$6683 ( \6936 , \6932 );
not \U$6684 ( \6937 , \6897 );
or \U$6685 ( \6938 , \6936 , \6937 );
xor \U$6686 ( \6939 , RIbe2a118_82, RIbe2a0a0_81);
xnor \U$6687 ( \6940 , RIbe2a0a0_81, RIbe2b360_121);
nand \U$6688 ( \6941 , \6939 , \6940 );
not \U$6689 ( \6942 , \6941 );
nand \U$6690 ( \6943 , \6942 , RIbe27b98_2);
not \U$6691 ( \6944 , RIbe2b360_121);
not \U$6692 ( \6945 , RIbe2a0a0_81);
or \U$6693 ( \6946 , \6944 , \6945 );
nand \U$6694 ( \6947 , \6946 , RIbe2a118_82);
buf \U$6695 ( \6948 , \6947 );
buf \U$6696 ( \6949 , \6948 );
not \U$6697 ( \6950 , \6949 );
and \U$6698 ( \6951 , \6943 , \6950 );
not \U$6699 ( \6952 , \6943 );
and \U$6700 ( \6953 , \6952 , \6948 );
nor \U$6701 ( \6954 , \6951 , \6953 );
not \U$6702 ( \6955 , \6954 );
not \U$6703 ( \6956 , \6955 );
not \U$6704 ( \6957 , RIbe27c10_3);
not \U$6705 ( \6958 , \6559 );
not \U$6706 ( \6959 , \6958 );
or \U$6707 ( \6960 , \6957 , \6959 );
buf \U$6708 ( \6961 , \6555 );
buf \U$6709 ( \6962 , \6961 );
buf \U$6710 ( \6963 , \6962 );
nand \U$6711 ( \6964 , \6963 , RIbe28e58_42);
nand \U$6712 ( \6965 , \6960 , \6964 );
xor \U$6713 ( \6966 , \6965 , \6572 );
not \U$6714 ( \6967 , \6966 );
not \U$6715 ( \6968 , \6967 );
or \U$6716 ( \6969 , \6956 , \6968 );
not \U$6717 ( \6970 , \6966 );
not \U$6718 ( \6971 , \6954 );
or \U$6719 ( \6972 , \6970 , \6971 );
not \U$6720 ( \6973 , RIbe28de0_41);
not \U$6721 ( \6974 , RIbe2a118_82);
not \U$6722 ( \6975 , RIbe2a820_97);
nand \U$6723 ( \6976 , \6974 , \6975 , RIbe2a898_98);
not \U$6724 ( \6977 , RIbe2a898_98);
nand \U$6725 ( \6978 , \6977 , RIbe2a118_82, RIbe2a820_97);
nand \U$6726 ( \6979 , \6976 , \6978 );
buf \U$6727 ( \6980 , \6979 );
not \U$6728 ( \6981 , \6980 );
or \U$6729 ( \6982 , \6973 , \6981 );
xor \U$6730 ( \6983 , RIbe2a820_97, RIbe2a118_82);
not \U$6731 ( \6984 , \6983 );
not \U$6732 ( \6985 , \6984 );
nand \U$6733 ( \6986 , \6985 , RIbe29920_65);
nand \U$6734 ( \6987 , \6982 , \6986 );
not \U$6735 ( \6988 , RIbe2a118_82);
not \U$6736 ( \6989 , RIbe2a820_97);
or \U$6737 ( \6990 , \6988 , \6989 );
nand \U$6738 ( \6991 , \6990 , RIbe2a898_98);
buf \U$6739 ( \6992 , \6991 );
not \U$6740 ( \6993 , \6992 );
and \U$6741 ( \6994 , \6987 , \6993 );
not \U$6742 ( \6995 , \6987 );
and \U$6743 ( \6996 , \6995 , \6992 );
nor \U$6744 ( \6997 , \6994 , \6996 );
nand \U$6745 ( \6998 , \6972 , \6997 );
nand \U$6746 ( \6999 , \6969 , \6998 );
nand \U$6747 ( \7000 , \6938 , \6999 );
nand \U$6748 ( \7001 , \6935 , \7000 );
nand \U$6749 ( \7002 , \6853 , \7001 );
nand \U$6750 ( \7003 , \6737 , \6852 );
and \U$6751 ( \7004 , \7002 , \7003 );
not \U$6752 ( \7005 , \7004 );
not \U$6753 ( \7006 , RIbe28a20_33);
not \U$6754 ( \7007 , \2570 );
not \U$6755 ( \7008 , \7007 );
or \U$6756 ( \7009 , \7006 , \7008 );
not \U$6757 ( \7010 , \3421 );
nand \U$6758 ( \7011 , \7010 , \3267 );
nand \U$6759 ( \7012 , \7009 , \7011 );
and \U$6760 ( \7013 , \7012 , \3272 );
not \U$6761 ( \7014 , \7012 );
and \U$6762 ( \7015 , \7014 , \2576 );
nor \U$6763 ( \7016 , \7013 , \7015 );
not \U$6764 ( \7017 , \7016 );
not \U$6765 ( \7018 , \7017 );
not \U$6766 ( \7019 , RIbe28930_31);
not \U$6767 ( \7020 , \6797 );
or \U$6768 ( \7021 , \7019 , \7020 );
nand \U$6769 ( \7022 , \6800 , RIbe29560_57);
nand \U$6770 ( \7023 , \7021 , \7022 );
and \U$6771 ( \7024 , \7023 , \3461 );
not \U$6772 ( \7025 , \7023 );
and \U$6773 ( \7026 , \7025 , \3290 );
nor \U$6774 ( \7027 , \7024 , \7026 );
not \U$6775 ( \7028 , \7027 );
not \U$6776 ( \7029 , \7028 );
or \U$6777 ( \7030 , \7018 , \7029 );
nand \U$6778 ( \7031 , \7027 , \7016 );
nand \U$6779 ( \7032 , \7030 , \7031 );
not \U$6780 ( \7033 , \4065 );
not \U$6781 ( \7034 , \5423 );
and \U$6782 ( \7035 , \7033 , \7034 );
and \U$6783 ( \7036 , \1272 , RIbe28b88_36);
nor \U$6784 ( \7037 , \7035 , \7036 );
not \U$6785 ( \7038 , \3515 );
and \U$6786 ( \7039 , \7037 , \7038 );
not \U$6787 ( \7040 , \7037 );
and \U$6788 ( \7041 , \7040 , \1277 );
nor \U$6789 ( \7042 , \7039 , \7041 );
xnor \U$6790 ( \7043 , \7032 , \7042 );
not \U$6791 ( \7044 , RIbe280c0_13);
not \U$6792 ( \7045 , \4804 );
or \U$6793 ( \7046 , \7044 , \7045 );
nand \U$6794 ( \7047 , \6418 , RIbe29830_63);
nand \U$6795 ( \7048 , \7046 , \7047 );
and \U$6796 ( \7049 , \7048 , \4326 );
not \U$6797 ( \7050 , \7048 );
and \U$6798 ( \7051 , \7050 , \4323 );
nor \U$6799 ( \7052 , \7049 , \7051 );
not \U$6800 ( \7053 , RIbe296c8_60);
not \U$6801 ( \7054 , \6427 );
or \U$6802 ( \7055 , \7053 , \7054 );
buf \U$6803 ( \7056 , \5730 );
nand \U$6804 ( \7057 , \7056 , RIbe29650_59);
nand \U$6805 ( \7058 , \7055 , \7057 );
and \U$6806 ( \7059 , \7058 , \4586 );
not \U$6807 ( \7060 , \7058 );
and \U$6808 ( \7061 , \7060 , \4592 );
nor \U$6809 ( \7062 , \7059 , \7061 );
xor \U$6810 ( \7063 , \7052 , \7062 );
not \U$6811 ( \7064 , RIbe28228_16);
not \U$6812 ( \7065 , \4021 );
or \U$6813 ( \7066 , \7064 , \7065 );
nand \U$6814 ( \7067 , \4333 , RIbe281b0_15);
nand \U$6815 ( \7068 , \7066 , \7067 );
and \U$6816 ( \7069 , \7068 , \3471 );
not \U$6817 ( \7070 , \7068 );
and \U$6818 ( \7071 , \7070 , \4821 );
nor \U$6819 ( \7072 , \7069 , \7071 );
xor \U$6820 ( \7073 , \7063 , \7072 );
xor \U$6821 ( \7074 , \7043 , \7073 );
not \U$6822 ( \7075 , \6883 );
buf \U$6823 ( \7076 , \7075 );
and \U$6824 ( \7077 , \7076 , RIbe27d00_5);
and \U$6825 ( \7078 , \6536 , RIbe27d78_6);
nor \U$6826 ( \7079 , \7077 , \7078 );
and \U$6827 ( \7080 , \7079 , \6891 );
not \U$6828 ( \7081 , \7079 );
and \U$6829 ( \7082 , \7081 , \6546 );
nor \U$6830 ( \7083 , \7080 , \7082 );
not \U$6831 ( \7084 , RIbe290b0_47);
not \U$6832 ( \7085 , \6139 );
or \U$6833 ( \7086 , \7084 , \7085 );
not \U$6834 ( \7087 , \6615 );
nand \U$6835 ( \7088 , \7087 , RIbe29a88_68);
nand \U$6836 ( \7089 , \7086 , \7088 );
and \U$6837 ( \7090 , \7089 , \6144 );
not \U$6838 ( \7091 , \7089 );
and \U$6839 ( \7092 , \7091 , \5740 );
nor \U$6840 ( \7093 , \7090 , \7092 );
xor \U$6841 ( \7094 , \7083 , \7093 );
not \U$6842 ( \7095 , RIbe29038_46);
not \U$6843 ( \7096 , \6630 );
or \U$6844 ( \7097 , \7095 , \7096 );
buf \U$6845 ( \7098 , \5747 );
not \U$6846 ( \7099 , \7098 );
buf \U$6847 ( \7100 , \7099 );
nand \U$6848 ( \7101 , \7100 , RIbe28fc0_45);
nand \U$6849 ( \7102 , \7097 , \7101 );
and \U$6850 ( \7103 , \7102 , \5047 );
not \U$6851 ( \7104 , \7102 );
and \U$6852 ( \7105 , \7104 , \5754 );
nor \U$6853 ( \7106 , \7103 , \7105 );
xor \U$6854 ( \7107 , \7094 , \7106 );
xor \U$6855 ( \7108 , \7074 , \7107 );
nand \U$6856 ( \7109 , \6722 , \6716 );
and \U$6857 ( \7110 , \7109 , \6734 );
nor \U$6858 ( \7111 , \6722 , \6716 );
nor \U$6859 ( \7112 , \7110 , \7111 );
not \U$6860 ( \7113 , \7112 );
not \U$6861 ( \7114 , \7113 );
and \U$6862 ( \7115 , \1679 , RIbe29fb0_79);
not \U$6863 ( \7116 , \285 );
and \U$6864 ( \7117 , \7116 , RIbe29e48_76);
nor \U$6865 ( \7118 , \7115 , \7117 );
and \U$6866 ( \7119 , \7118 , \293 );
not \U$6867 ( \7120 , \7118 );
and \U$6868 ( \7121 , \7120 , \300 );
nor \U$6869 ( \7122 , \7119 , \7121 );
not \U$6870 ( \7123 , \424 );
not \U$6871 ( \7124 , \7123 );
not \U$6872 ( \7125 , \7124 );
not \U$6873 ( \7126 , RIbe29bf0_71);
not \U$6874 ( \7127 , \546 );
or \U$6875 ( \7128 , \7126 , \7127 );
nand \U$6876 ( \7129 , \1327 , RIbe28f48_44);
nand \U$6877 ( \7130 , \7128 , \7129 );
not \U$6878 ( \7131 , \7130 );
and \U$6879 ( \7132 , \7125 , \7131 );
and \U$6880 ( \7133 , \7130 , \424 );
nor \U$6881 ( \7134 , \7132 , \7133 );
nand \U$6882 ( \7135 , \7122 , \7134 );
not \U$6883 ( \7136 , RIbe29dd0_75);
not \U$6884 ( \7137 , \1773 );
or \U$6885 ( \7138 , \7136 , \7137 );
nand \U$6886 ( \7139 , \429 , RIbe29c68_72);
nand \U$6887 ( \7140 , \7138 , \7139 );
and \U$6888 ( \7141 , \7140 , \306 );
not \U$6889 ( \7142 , \7140 );
and \U$6890 ( \7143 , \7142 , \1232 );
nor \U$6891 ( \7144 , \7141 , \7143 );
and \U$6892 ( \7145 , \7135 , \7144 );
nor \U$6893 ( \7146 , \7122 , \7134 );
nor \U$6894 ( \7147 , \7145 , \7146 );
not \U$6895 ( \7148 , \7147 );
or \U$6896 ( \7149 , \7114 , \7148 );
not \U$6897 ( \7150 , \7147 );
nand \U$6898 ( \7151 , \7150 , \7112 );
nand \U$6899 ( \7152 , \7149 , \7151 );
and \U$6900 ( \7153 , RIbe29380_53, RIbe2a370_87);
not \U$6901 ( \7154 , \7153 );
not \U$6902 ( \7155 , RIbe2a2f8_86);
not \U$6903 ( \7156 , \3160 );
or \U$6904 ( \7157 , \7155 , \7156 );
nand \U$6905 ( \7158 , \329 , RIbe2acd0_107);
nand \U$6906 ( \7159 , \7157 , \7158 );
xnor \U$6907 ( \7160 , \7159 , \1375 );
not \U$6908 ( \7161 , \7160 );
not \U$6909 ( \7162 , \7161 );
or \U$6910 ( \7163 , \7154 , \7162 );
not \U$6911 ( \7164 , \7153 );
nand \U$6912 ( \7165 , \7164 , \7160 );
nand \U$6913 ( \7166 , \7163 , \7165 );
xor \U$6914 ( \7167 , \7152 , \7166 );
not \U$6915 ( \7168 , \7167 );
nand \U$6916 ( \7169 , \7108 , \7168 );
and \U$6917 ( \7170 , \1756 , RIbe28f48_44);
and \U$6918 ( \7171 , \552 , RIbe28ed0_43);
nor \U$6919 ( \7172 , \7170 , \7171 );
not \U$6920 ( \7173 , \7172 );
not \U$6921 ( \7174 , \425 );
and \U$6922 ( \7175 , \7173 , \7174 );
and \U$6923 ( \7176 , \7172 , \1761 );
nor \U$6924 ( \7177 , \7175 , \7176 );
not \U$6925 ( \7178 , \7177 );
not \U$6926 ( \7179 , \1611 );
not \U$6927 ( \7180 , RIbe27f58_10);
not \U$6928 ( \7181 , \7180 );
and \U$6929 ( \7182 , \7179 , \7181 );
and \U$6930 ( \7183 , \2531 , RIbe27fd0_11);
nor \U$6931 ( \7184 , \7182 , \7183 );
and \U$6932 ( \7185 , \7184 , \3959 );
not \U$6933 ( \7186 , \7184 );
and \U$6934 ( \7187 , \7186 , \1618 );
nor \U$6935 ( \7188 , \7185 , \7187 );
xor \U$6936 ( \7189 , \7178 , \7188 );
and \U$6937 ( \7190 , \5973 , RIbe27e68_8);
and \U$6938 ( \7191 , \1203 , RIbe28660_25);
nor \U$6939 ( \7192 , \7190 , \7191 );
and \U$6940 ( \7193 , \7192 , \1011 );
not \U$6941 ( \7194 , \7192 );
and \U$6942 ( \7195 , \7194 , \1813 );
nor \U$6943 ( \7196 , \7193 , \7195 );
and \U$6944 ( \7197 , \7189 , \7196 );
not \U$6945 ( \7198 , \7189 );
not \U$6946 ( \7199 , \7196 );
and \U$6947 ( \7200 , \7198 , \7199 );
nor \U$6948 ( \7201 , \7197 , \7200 );
not \U$6949 ( \7202 , \7201 );
not \U$6950 ( \7203 , \7202 );
not \U$6951 ( \7204 , RIbe29c68_72);
not \U$6952 ( \7205 , \1773 );
or \U$6953 ( \7206 , \7204 , \7205 );
nand \U$6954 ( \7207 , \429 , RIbe29bf0_71);
nand \U$6955 ( \7208 , \7206 , \7207 );
and \U$6956 ( \7209 , \7208 , \306 );
not \U$6957 ( \7210 , \7208 );
and \U$6958 ( \7211 , \7210 , \1232 );
nor \U$6959 ( \7212 , \7209 , \7211 );
and \U$6960 ( \7213 , \1252 , RIbe29e48_76);
and \U$6961 ( \7214 , \1531 , RIbe29dd0_75);
nor \U$6962 ( \7215 , \7213 , \7214 );
and \U$6963 ( \7216 , \7215 , \300 );
not \U$6964 ( \7217 , \7215 );
and \U$6965 ( \7218 , \7217 , \293 );
nor \U$6966 ( \7219 , \7216 , \7218 );
xor \U$6967 ( \7220 , \7212 , \7219 );
and \U$6968 ( \7221 , \260 , RIbe2a028_80);
and \U$6969 ( \7222 , \264 , RIbe29fb0_79);
nor \U$6970 ( \7223 , \7221 , \7222 );
and \U$6971 ( \7224 , \7223 , \1362 );
not \U$6972 ( \7225 , \7223 );
and \U$6973 ( \7226 , \7225 , \1363 );
nor \U$6974 ( \7227 , \7224 , \7226 );
xor \U$6975 ( \7228 , \7220 , \7227 );
not \U$6976 ( \7229 , \7228 );
and \U$6977 ( \7230 , \2555 , RIbe28390_19);
and \U$6978 ( \7231 , \1117 , RIbe28b10_35);
nor \U$6979 ( \7232 , \7230 , \7231 );
and \U$6980 ( \7233 , \7232 , \1448 );
not \U$6981 ( \7234 , \7232 );
and \U$6982 ( \7235 , \7234 , \1132 );
nor \U$6983 ( \7236 , \7233 , \7235 );
not \U$6984 ( \7237 , RIbe28480_21);
not \U$6985 ( \7238 , \1633 );
or \U$6986 ( \7239 , \7237 , \7238 );
nand \U$6987 ( \7240 , \1455 , RIbe28408_20);
nand \U$6988 ( \7241 , \7239 , \7240 );
and \U$6989 ( \7242 , \7241 , \2418 );
not \U$6990 ( \7243 , \7241 );
and \U$6991 ( \7244 , \7243 , \1309 );
nor \U$6992 ( \7245 , \7242 , \7244 );
xor \U$6993 ( \7246 , \7236 , \7245 );
not \U$6994 ( \7247 , \1157 );
not \U$6995 ( \7248 , RIbe285e8_24);
not \U$6996 ( \7249 , \2597 );
or \U$6997 ( \7250 , \7248 , \7249 );
nand \U$6998 ( \7251 , \1147 , RIbe287c8_28);
nand \U$6999 ( \7252 , \7250 , \7251 );
not \U$7000 ( \7253 , \7252 );
or \U$7001 ( \7254 , \7247 , \7253 );
or \U$7002 ( \7255 , \7252 , \1157 );
nand \U$7003 ( \7256 , \7254 , \7255 );
xor \U$7004 ( \7257 , \7246 , \7256 );
not \U$7005 ( \7258 , \7257 );
or \U$7006 ( \7259 , \7229 , \7258 );
or \U$7007 ( \7260 , \7257 , \7228 );
nand \U$7008 ( \7261 , \7259 , \7260 );
not \U$7009 ( \7262 , \7261 );
or \U$7010 ( \7263 , \7203 , \7262 );
or \U$7011 ( \7264 , \7261 , \7202 );
nand \U$7012 ( \7265 , \7263 , \7264 );
and \U$7013 ( \7266 , \7169 , \7265 );
nor \U$7014 ( \7267 , \7108 , \7168 );
nor \U$7015 ( \7268 , \7266 , \7267 );
not \U$7016 ( \7269 , \7268 );
or \U$7017 ( \7270 , \7005 , \7269 );
not \U$7018 ( \7271 , \6582 );
not \U$7019 ( \7272 , \7271 );
not \U$7020 ( \7273 , RIbe27c10_3);
not \U$7021 ( \7274 , \6590 );
not \U$7022 ( \7275 , \7274 );
or \U$7023 ( \7276 , \7273 , \7275 );
buf \U$7024 ( \7277 , \6586 );
buf \U$7025 ( \7278 , \7277 );
nand \U$7026 ( \7279 , \7278 , RIbe28e58_42);
nand \U$7027 ( \7280 , \7276 , \7279 );
not \U$7028 ( \7281 , \7280 );
or \U$7029 ( \7282 , \7272 , \7281 );
or \U$7030 ( \7283 , \7280 , \6873 );
nand \U$7031 ( \7284 , \7282 , \7283 );
not \U$7032 ( \7285 , RIbe28de0_41);
not \U$7033 ( \7286 , \6561 );
or \U$7034 ( \7287 , \7285 , \7286 );
nand \U$7035 ( \7288 , \6963 , RIbe29920_65);
nand \U$7036 ( \7289 , \7287 , \7288 );
and \U$7037 ( \7290 , RIbe2aa00_101, RIbe2a898_98);
not \U$7038 ( \7291 , RIbe2aa78_102);
nor \U$7039 ( \7292 , \7290 , \7291 );
buf \U$7040 ( \7293 , \7292 );
and \U$7041 ( \7294 , \7289 , \7293 );
not \U$7042 ( \7295 , \7289 );
and \U$7043 ( \7296 , \7295 , \6572 );
nor \U$7044 ( \7297 , \7294 , \7296 );
buf \U$7045 ( \7298 , \6979 );
buf \U$7046 ( \7299 , \7298 );
nand \U$7047 ( \7300 , \7299 , RIbe27b98_2);
buf \U$7048 ( \7301 , \6991 );
and \U$7049 ( \7302 , \7300 , \7301 );
not \U$7050 ( \7303 , \7300 );
not \U$7051 ( \7304 , \6992 );
and \U$7052 ( \7305 , \7303 , \7304 );
nor \U$7053 ( \7306 , \7302 , \7305 );
xor \U$7054 ( \7307 , \7297 , \7306 );
xnor \U$7055 ( \7308 , \7284 , \7307 );
not \U$7056 ( \7309 , \7308 );
not \U$7057 ( \7310 , \7134 );
not \U$7058 ( \7311 , \7144 );
or \U$7059 ( \7312 , \7310 , \7311 );
or \U$7060 ( \7313 , \7144 , \7134 );
nand \U$7061 ( \7314 , \7312 , \7313 );
xor \U$7062 ( \7315 , \7314 , \7122 );
not \U$7063 ( \7316 , \7315 );
not \U$7064 ( \7317 , RIbe28408_20);
not \U$7065 ( \7318 , \2554 );
or \U$7066 ( \7319 , \7317 , \7318 );
nand \U$7067 ( \7320 , \5467 , RIbe28390_19);
nand \U$7068 ( \7321 , \7319 , \7320 );
not \U$7069 ( \7322 , \7321 );
not \U$7070 ( \7323 , \1448 );
and \U$7071 ( \7324 , \7322 , \7323 );
and \U$7072 ( \7325 , \7321 , \6831 );
nor \U$7073 ( \7326 , \7324 , \7325 );
not \U$7074 ( \7327 , RIbe28b10_35);
not \U$7075 ( \7328 , \4295 );
or \U$7076 ( \7329 , \7327 , \7328 );
nand \U$7077 ( \7330 , \2384 , RIbe28b88_36);
nand \U$7078 ( \7331 , \7329 , \7330 );
not \U$7079 ( \7332 , \7331 );
not \U$7080 ( \7333 , \3516 );
and \U$7081 ( \7334 , \7332 , \7333 );
and \U$7082 ( \7335 , \7331 , \7038 );
nor \U$7083 ( \7336 , \7334 , \7335 );
xor \U$7084 ( \7337 , \7326 , \7336 );
not \U$7085 ( \7338 , RIbe287c8_28);
not \U$7086 ( \7339 , \1633 );
or \U$7087 ( \7340 , \7338 , \7339 );
nand \U$7088 ( \7341 , \4730 , RIbe28480_21);
nand \U$7089 ( \7342 , \7340 , \7341 );
and \U$7090 ( \7343 , \7342 , \2418 );
not \U$7091 ( \7344 , \7342 );
and \U$7092 ( \7345 , \7344 , \1309 );
nor \U$7093 ( \7346 , \7343 , \7345 );
xor \U$7094 ( \7347 , \7337 , \7346 );
not \U$7095 ( \7348 , \7347 );
or \U$7096 ( \7349 , \7316 , \7348 );
not \U$7097 ( \7350 , RIbe28660_25);
not \U$7098 ( \7351 , \1143 );
or \U$7099 ( \7352 , \7350 , \7351 );
nand \U$7100 ( \7353 , \1147 , RIbe285e8_24);
nand \U$7101 ( \7354 , \7352 , \7353 );
and \U$7102 ( \7355 , \7354 , \1469 );
not \U$7103 ( \7356 , \7354 );
and \U$7104 ( \7357 , \7356 , \1152 );
nor \U$7105 ( \7358 , \7355 , \7357 );
not \U$7106 ( \7359 , \6345 );
not \U$7107 ( \7360 , RIbe27fd0_11);
not \U$7108 ( \7361 , \7360 );
and \U$7109 ( \7362 , \7359 , \7361 );
not \U$7110 ( \7363 , \1743 );
and \U$7111 ( \7364 , \7363 , RIbe28ed0_43);
nor \U$7112 ( \7365 , \7362 , \7364 );
and \U$7113 ( \7366 , \7365 , \564 );
not \U$7114 ( \7367 , \7365 );
and \U$7115 ( \7368 , \7367 , \1621 );
nor \U$7116 ( \7369 , \7366 , \7368 );
xor \U$7117 ( \7370 , \7358 , \7369 );
and \U$7118 ( \7371 , \1807 , RIbe27f58_10);
and \U$7119 ( \7372 , \2000 , RIbe27e68_8);
nor \U$7120 ( \7373 , \7371 , \7372 );
and \U$7121 ( \7374 , \7373 , \752 );
not \U$7122 ( \7375 , \7373 );
and \U$7123 ( \7376 , \7375 , \1011 );
nor \U$7124 ( \7377 , \7374 , \7376 );
xor \U$7125 ( \7378 , \7370 , \7377 );
nand \U$7126 ( \7379 , \7349 , \7378 );
not \U$7127 ( \7380 , \7347 );
not \U$7128 ( \7381 , \7315 );
nand \U$7129 ( \7382 , \7380 , \7381 );
nand \U$7130 ( \7383 , \7379 , \7382 );
not \U$7131 ( \7384 , \7383 );
not \U$7132 ( \7385 , \7384 );
or \U$7133 ( \7386 , \7309 , \7385 );
not \U$7134 ( \7387 , \4592 );
not \U$7135 ( \7388 , RIbe29830_63);
not \U$7136 ( \7389 , \5727 );
or \U$7137 ( \7390 , \7388 , \7389 );
nand \U$7138 ( \7391 , \7056 , RIbe296c8_60);
nand \U$7139 ( \7392 , \7390 , \7391 );
not \U$7140 ( \7393 , \7392 );
or \U$7141 ( \7394 , \7387 , \7393 );
or \U$7142 ( \7395 , \7392 , \4592 );
nand \U$7143 ( \7396 , \7394 , \7395 );
not \U$7144 ( \7397 , \7396 );
not \U$7145 ( \7398 , \5754 );
not \U$7146 ( \7399 , RIbe29650_59);
not \U$7147 ( \7400 , \5455 );
or \U$7148 ( \7401 , \7399 , \7400 );
nand \U$7149 ( \7402 , \5751 , RIbe29038_46);
nand \U$7150 ( \7403 , \7401 , \7402 );
not \U$7151 ( \7404 , \7403 );
and \U$7152 ( \7405 , \7398 , \7404 );
and \U$7153 ( \7406 , \7403 , \6641 );
nor \U$7154 ( \7407 , \7405 , \7406 );
not \U$7155 ( \7408 , \7407 );
or \U$7156 ( \7409 , \7397 , \7408 );
or \U$7157 ( \7410 , \7407 , \7396 );
nand \U$7158 ( \7411 , \7409 , \7410 );
not \U$7159 ( \7412 , \4323 );
not \U$7160 ( \7413 , RIbe281b0_15);
not \U$7161 ( \7414 , \5058 );
or \U$7162 ( \7415 , \7413 , \7414 );
nand \U$7163 ( \7416 , \4809 , RIbe280c0_13);
nand \U$7164 ( \7417 , \7415 , \7416 );
not \U$7165 ( \7418 , \7417 );
or \U$7166 ( \7419 , \7412 , \7418 );
or \U$7167 ( \7420 , \7417 , \4323 );
nand \U$7168 ( \7421 , \7419 , \7420 );
xnor \U$7169 ( \7422 , \7411 , \7421 );
not \U$7170 ( \7423 , \7422 );
not \U$7171 ( \7424 , RIbe289a8_32);
not \U$7172 ( \7425 , \4764 );
or \U$7173 ( \7426 , \7424 , \7425 );
nand \U$7174 ( \7427 , \4011 , RIbe28930_31);
nand \U$7175 ( \7428 , \7426 , \7427 );
and \U$7176 ( \7429 , \7428 , \3290 );
not \U$7177 ( \7430 , \7428 );
and \U$7178 ( \7431 , \7430 , \2887 );
nor \U$7179 ( \7432 , \7429 , \7431 );
not \U$7180 ( \7433 , \7432 );
not \U$7181 ( \7434 , \7433 );
not \U$7182 ( \7435 , RIbe29560_57);
not \U$7183 ( \7436 , \4021 );
or \U$7184 ( \7437 , \7435 , \7436 );
not \U$7185 ( \7438 , \4025 );
nand \U$7186 ( \7439 , \7438 , RIbe28228_16);
nand \U$7187 ( \7440 , \7437 , \7439 );
and \U$7188 ( \7441 , \7440 , \4821 );
not \U$7189 ( \7442 , \7440 );
and \U$7190 ( \7443 , \7442 , \3471 );
nor \U$7191 ( \7444 , \7441 , \7443 );
not \U$7192 ( \7445 , \7444 );
not \U$7193 ( \7446 , \7445 );
or \U$7194 ( \7447 , \7434 , \7446 );
nand \U$7195 ( \7448 , \7432 , \7444 );
nand \U$7196 ( \7449 , \7447 , \7448 );
not \U$7197 ( \7450 , RIbe29290_51);
not \U$7198 ( \7451 , \4050 );
or \U$7199 ( \7452 , \7450 , \7451 );
nand \U$7200 ( \7453 , \3267 , RIbe28a20_33);
nand \U$7201 ( \7454 , \7452 , \7453 );
and \U$7202 ( \7455 , \7454 , \2576 );
not \U$7203 ( \7456 , \7454 );
not \U$7204 ( \7457 , \2379 );
and \U$7205 ( \7458 , \7456 , \7457 );
nor \U$7206 ( \7459 , \7455 , \7458 );
and \U$7207 ( \7460 , \7449 , \7459 );
not \U$7208 ( \7461 , \7449 );
not \U$7209 ( \7462 , \7459 );
and \U$7210 ( \7463 , \7461 , \7462 );
nor \U$7211 ( \7464 , \7460 , \7463 );
not \U$7212 ( \7465 , \7464 );
or \U$7213 ( \7466 , \7423 , \7465 );
not \U$7214 ( \7467 , RIbe29a88_68);
not \U$7215 ( \7468 , \6536 );
or \U$7216 ( \7469 , \7467 , \7468 );
nand \U$7217 ( \7470 , \6540 , RIbe27d78_6);
nand \U$7218 ( \7471 , \7469 , \7470 );
not \U$7219 ( \7472 , \7471 );
not \U$7220 ( \7473 , \6548 );
and \U$7221 ( \7474 , \7472 , \7473 );
and \U$7222 ( \7475 , \7471 , \6891 );
nor \U$7223 ( \7476 , \7474 , \7475 );
not \U$7224 ( \7477 , \7476 );
not \U$7225 ( \7478 , \7477 );
not \U$7226 ( \7479 , RIbe27d00_5);
not \U$7227 ( \7480 , \6592 );
or \U$7228 ( \7481 , \7479 , \7480 );
not \U$7229 ( \7482 , \7277 );
not \U$7230 ( \7483 , \7482 );
nand \U$7231 ( \7484 , \7483 , RIbe27c10_3);
nand \U$7232 ( \7485 , \7481 , \7484 );
and \U$7233 ( \7486 , \7485 , \6582 );
not \U$7234 ( \7487 , \7485 );
not \U$7235 ( \7488 , \6582 );
and \U$7236 ( \7489 , \7487 , \7488 );
nor \U$7237 ( \7490 , \7486 , \7489 );
not \U$7238 ( \7491 , \7490 );
not \U$7239 ( \7492 , \7491 );
or \U$7240 ( \7493 , \7478 , \7492 );
nand \U$7241 ( \7494 , \7490 , \7476 );
nand \U$7242 ( \7495 , \7493 , \7494 );
not \U$7243 ( \7496 , RIbe28fc0_45);
not \U$7244 ( \7497 , \6139 );
or \U$7245 ( \7498 , \7496 , \7497 );
nand \U$7246 ( \7499 , \7087 , RIbe290b0_47);
nand \U$7247 ( \7500 , \7498 , \7499 );
not \U$7248 ( \7501 , \5740 );
and \U$7249 ( \7502 , \7500 , \7501 );
not \U$7250 ( \7503 , \7500 );
and \U$7251 ( \7504 , \7503 , \5740 );
nor \U$7252 ( \7505 , \7502 , \7504 );
not \U$7253 ( \7506 , \7505 );
and \U$7254 ( \7507 , \7495 , \7506 );
not \U$7255 ( \7508 , \7495 );
and \U$7256 ( \7509 , \7508 , \7505 );
nor \U$7257 ( \7510 , \7507 , \7509 );
not \U$7258 ( \7511 , \7510 );
nand \U$7259 ( \7512 , \7466 , \7511 );
not \U$7260 ( \7513 , \7464 );
not \U$7261 ( \7514 , \7422 );
nand \U$7262 ( \7515 , \7513 , \7514 );
nand \U$7263 ( \7516 , \7512 , \7515 );
nand \U$7264 ( \7517 , \7386 , \7516 );
not \U$7265 ( \7518 , \7308 );
nand \U$7266 ( \7519 , \7518 , \7383 );
nand \U$7267 ( \7520 , \7517 , \7519 );
nand \U$7268 ( \7521 , \7270 , \7520 );
or \U$7269 ( \7522 , \7268 , \7004 );
nand \U$7270 ( \7523 , \7521 , \7522 );
xor \U$7271 ( \7524 , \6661 , \7523 );
not \U$7272 ( \7525 , RIbe29a88_68);
not \U$7273 ( \7526 , \6139 );
or \U$7274 ( \7527 , \7525 , \7526 );
not \U$7275 ( \7528 , \6615 );
nand \U$7276 ( \7529 , \7528 , RIbe27d78_6);
nand \U$7277 ( \7530 , \7527 , \7529 );
not \U$7278 ( \7531 , \7530 );
not \U$7279 ( \7532 , \5740 );
and \U$7280 ( \7533 , \7531 , \7532 );
not \U$7281 ( \7534 , \5740 );
not \U$7282 ( \7535 , \7534 );
and \U$7283 ( \7536 , \7530 , \7535 );
nor \U$7284 ( \7537 , \7533 , \7536 );
not \U$7285 ( \7538 , RIbe27d00_5);
not \U$7286 ( \7539 , \6537 );
or \U$7287 ( \7540 , \7538 , \7539 );
nand \U$7288 ( \7541 , \6540 , RIbe27c10_3);
nand \U$7289 ( \7542 , \7540 , \7541 );
not \U$7290 ( \7543 , \7542 );
not \U$7291 ( \7544 , \6551 );
and \U$7292 ( \7545 , \7543 , \7544 );
not \U$7293 ( \7546 , \6546 );
and \U$7294 ( \7547 , \7542 , \7546 );
nor \U$7295 ( \7548 , \7545 , \7547 );
not \U$7296 ( \7549 , \7548 );
and \U$7297 ( \7550 , \7537 , \7549 );
not \U$7298 ( \7551 , \7537 );
and \U$7299 ( \7552 , \7551 , \7548 );
or \U$7300 ( \7553 , \7550 , \7552 );
not \U$7301 ( \7554 , RIbe28fc0_45);
not \U$7302 ( \7555 , \5455 );
or \U$7303 ( \7556 , \7554 , \7555 );
nand \U$7304 ( \7557 , \7100 , RIbe290b0_47);
nand \U$7305 ( \7558 , \7556 , \7557 );
and \U$7306 ( \7559 , \7558 , \5457 );
not \U$7307 ( \7560 , \7558 );
and \U$7308 ( \7561 , \7560 , \6117 );
nor \U$7309 ( \7562 , \7559 , \7561 );
not \U$7310 ( \7563 , \7562 );
and \U$7311 ( \7564 , \7553 , \7563 );
not \U$7312 ( \7565 , \7553 );
and \U$7313 ( \7566 , \7565 , \7562 );
nor \U$7314 ( \7567 , \7564 , \7566 );
not \U$7315 ( \7568 , \7043 );
not \U$7316 ( \7569 , \7568 );
not \U$7317 ( \7570 , \7073 );
or \U$7318 ( \7571 , \7569 , \7570 );
or \U$7319 ( \7572 , \7073 , \7568 );
nand \U$7320 ( \7573 , \7572 , \7107 );
nand \U$7321 ( \7574 , \7571 , \7573 );
xor \U$7322 ( \7575 , \7567 , \7574 );
not \U$7323 ( \7576 , \7228 );
not \U$7324 ( \7577 , \7257 );
not \U$7325 ( \7578 , \7577 );
or \U$7326 ( \7579 , \7576 , \7578 );
or \U$7327 ( \7580 , \7577 , \7228 );
nand \U$7328 ( \7581 , \7580 , \7201 );
nand \U$7329 ( \7582 , \7579 , \7581 );
xor \U$7330 ( \7583 , \7575 , \7582 );
and \U$7331 ( \7584 , \326 , RIbe2acd0_107);
and \U$7332 ( \7585 , \330 , RIbe2a028_80);
nor \U$7333 ( \7586 , \7584 , \7585 );
and \U$7334 ( \7587 , \7586 , \339 );
not \U$7335 ( \7588 , \7586 );
and \U$7336 ( \7589 , \7588 , \342 );
nor \U$7337 ( \7590 , \7587 , \7589 );
xor \U$7338 ( \7591 , \7590 , \7165 );
xor \U$7339 ( \7592 , \7212 , \7219 );
and \U$7340 ( \7593 , \7592 , \7227 );
and \U$7341 ( \7594 , \7212 , \7219 );
or \U$7342 ( \7595 , \7593 , \7594 );
xor \U$7343 ( \7596 , \7591 , \7595 );
not \U$7344 ( \7597 , \7017 );
not \U$7345 ( \7598 , \7027 );
or \U$7346 ( \7599 , \7597 , \7598 );
nand \U$7347 ( \7600 , \7599 , \7042 );
nand \U$7348 ( \7601 , \7028 , \7016 );
nand \U$7349 ( \7602 , \7600 , \7601 );
not \U$7350 ( \7603 , \7199 );
not \U$7351 ( \7604 , \7178 );
or \U$7352 ( \7605 , \7603 , \7604 );
not \U$7353 ( \7606 , \7188 );
nand \U$7354 ( \7607 , \7177 , \7196 );
nand \U$7355 ( \7608 , \7606 , \7607 );
nand \U$7356 ( \7609 , \7605 , \7608 );
xor \U$7357 ( \7610 , \7602 , \7609 );
not \U$7358 ( \7611 , \7256 );
not \U$7359 ( \7612 , \7245 );
not \U$7360 ( \7613 , \7612 );
or \U$7361 ( \7614 , \7611 , \7613 );
or \U$7362 ( \7615 , \7612 , \7256 );
nand \U$7363 ( \7616 , \7615 , \7236 );
nand \U$7364 ( \7617 , \7614 , \7616 );
xor \U$7365 ( \7618 , \7610 , \7617 );
xor \U$7366 ( \7619 , \7596 , \7618 );
not \U$7367 ( \7620 , \7306 );
not \U$7368 ( \7621 , \7284 );
or \U$7369 ( \7622 , \7620 , \7621 );
or \U$7370 ( \7623 , \7284 , \7306 );
nand \U$7371 ( \7624 , \7623 , \7297 );
nand \U$7372 ( \7625 , \7622 , \7624 );
xor \U$7373 ( \7626 , \7052 , \7062 );
and \U$7374 ( \7627 , \7626 , \7072 );
and \U$7375 ( \7628 , \7052 , \7062 );
or \U$7376 ( \7629 , \7627 , \7628 );
xor \U$7377 ( \7630 , \7625 , \7629 );
xor \U$7378 ( \7631 , \7083 , \7093 );
and \U$7379 ( \7632 , \7631 , \7106 );
and \U$7380 ( \7633 , \7083 , \7093 );
or \U$7381 ( \7634 , \7632 , \7633 );
xor \U$7382 ( \7635 , \7630 , \7634 );
xor \U$7383 ( \7636 , \7619 , \7635 );
xor \U$7384 ( \7637 , \7583 , \7636 );
not \U$7385 ( \7638 , RIbe28e58_42);
not \U$7386 ( \7639 , \6592 );
or \U$7387 ( \7640 , \7638 , \7639 );
nand \U$7388 ( \7641 , \7278 , RIbe28de0_41);
nand \U$7389 ( \7642 , \7640 , \7641 );
not \U$7390 ( \7643 , \7642 );
not \U$7391 ( \7644 , \6602 );
and \U$7392 ( \7645 , \7643 , \7644 );
not \U$7393 ( \7646 , \6582 );
and \U$7394 ( \7647 , \7642 , \7646 );
nor \U$7395 ( \7648 , \7645 , \7647 );
not \U$7396 ( \7649 , \7648 );
not \U$7397 ( \7650 , RIbe29920_65);
not \U$7398 ( \7651 , \6561 );
or \U$7399 ( \7652 , \7650 , \7651 );
buf \U$7400 ( \7653 , \6963 );
nand \U$7401 ( \7654 , \7653 , RIbe27b98_2);
nand \U$7402 ( \7655 , \7652 , \7654 );
and \U$7403 ( \7656 , \7655 , \7293 );
not \U$7404 ( \7657 , \7655 );
and \U$7405 ( \7658 , \7657 , \6572 );
nor \U$7406 ( \7659 , \7656 , \7658 );
not \U$7407 ( \7660 , \7301 );
not \U$7408 ( \7661 , \7660 );
and \U$7409 ( \7662 , \7659 , \7661 );
not \U$7410 ( \7663 , \7659 );
and \U$7411 ( \7664 , \7663 , \7660 );
nor \U$7412 ( \7665 , \7662 , \7664 );
not \U$7413 ( \7666 , \7665 );
or \U$7414 ( \7667 , \7649 , \7666 );
or \U$7415 ( \7668 , \7665 , \7648 );
nand \U$7416 ( \7669 , \7667 , \7668 );
xor \U$7417 ( \7670 , \6299 , \6332 );
xor \U$7418 ( \7671 , \7670 , \6365 );
xor \U$7419 ( \7672 , \7669 , \7671 );
not \U$7420 ( \7673 , \6483 );
not \U$7421 ( \7674 , \6449 );
or \U$7422 ( \7675 , \7673 , \7674 );
or \U$7423 ( \7676 , \6449 , \6483 );
nand \U$7424 ( \7677 , \7675 , \7676 );
and \U$7425 ( \7678 , \7677 , \6409 );
not \U$7426 ( \7679 , \7677 );
and \U$7427 ( \7680 , \7679 , \6408 );
nor \U$7428 ( \7681 , \7678 , \7680 );
xor \U$7429 ( \7682 , \7672 , \7681 );
and \U$7430 ( \7683 , \7637 , \7682 );
and \U$7431 ( \7684 , \7583 , \7636 );
or \U$7432 ( \7685 , \7683 , \7684 );
xor \U$7433 ( \7686 , \7524 , \7685 );
and \U$7434 ( \7687 , \6877 , \6894 );
not \U$7435 ( \7688 , \6877 );
and \U$7436 ( \7689 , \7688 , \6893 );
or \U$7437 ( \7690 , \7687 , \7689 );
xor \U$7438 ( \7691 , \7690 , \6866 );
and \U$7439 ( \7692 , \6997 , \6954 );
not \U$7440 ( \7693 , \6997 );
and \U$7441 ( \7694 , \7693 , \6955 );
or \U$7442 ( \7695 , \7692 , \7694 );
and \U$7443 ( \7696 , \7695 , \6966 );
not \U$7444 ( \7697 , \7695 );
and \U$7445 ( \7698 , \7697 , \6967 );
nor \U$7446 ( \7699 , \7696 , \7698 );
nor \U$7447 ( \7700 , \7691 , \7699 );
xor \U$7448 ( \7701 , \6826 , \6835 );
xnor \U$7449 ( \7702 , \7701 , \6845 );
not \U$7450 ( \7703 , \7702 );
not \U$7451 ( \7704 , \6794 );
not \U$7452 ( \7705 , \6807 );
or \U$7453 ( \7706 , \7704 , \7705 );
nand \U$7454 ( \7707 , \6793 , \6806 );
nand \U$7455 ( \7708 , \7706 , \7707 );
not \U$7456 ( \7709 , \6781 );
and \U$7457 ( \7710 , \7708 , \7709 );
not \U$7458 ( \7711 , \7708 );
and \U$7459 ( \7712 , \7711 , \6781 );
nor \U$7460 ( \7713 , \7710 , \7712 );
not \U$7461 ( \7714 , \7713 );
not \U$7462 ( \7715 , \6929 );
not \U$7463 ( \7716 , \6909 );
or \U$7464 ( \7717 , \7715 , \7716 );
or \U$7465 ( \7718 , \6929 , \6909 );
nand \U$7466 ( \7719 , \7717 , \7718 );
xor \U$7467 ( \7720 , \7719 , \6918 );
nand \U$7468 ( \7721 , \7714 , \7720 );
nand \U$7469 ( \7722 , \7703 , \7721 );
not \U$7470 ( \7723 , \7720 );
nand \U$7471 ( \7724 , \7723 , \7713 );
nand \U$7472 ( \7725 , \7722 , \7724 );
xor \U$7473 ( \7726 , \7700 , \7725 );
xor \U$7474 ( \7727 , \6662 , \6668 );
xor \U$7475 ( \7728 , \7727 , \6676 );
not \U$7476 ( \7729 , \7728 );
not \U$7477 ( \7730 , \7729 );
not \U$7478 ( \7731 , \6688 );
not \U$7479 ( \7732 , \6706 );
or \U$7480 ( \7733 , \7731 , \7732 );
not \U$7481 ( \7734 , \6688 );
nand \U$7482 ( \7735 , \7734 , \6705 );
nand \U$7483 ( \7736 , \7733 , \7735 );
xor \U$7484 ( \7737 , \7736 , \6695 );
not \U$7485 ( \7738 , \7737 );
not \U$7486 ( \7739 , \7738 );
or \U$7487 ( \7740 , \7730 , \7739 );
not \U$7488 ( \7741 , \7728 );
not \U$7489 ( \7742 , \7737 );
or \U$7490 ( \7743 , \7741 , \7742 );
not \U$7491 ( \7744 , \6746 );
not \U$7492 ( \7745 , \6767 );
or \U$7493 ( \7746 , \7744 , \7745 );
not \U$7494 ( \7747 , \6746 );
nand \U$7495 ( \7748 , \7747 , \6766 );
nand \U$7496 ( \7749 , \7746 , \7748 );
xnor \U$7497 ( \7750 , \7749 , \6754 );
nand \U$7498 ( \7751 , \7743 , \7750 );
nand \U$7499 ( \7752 , \7740 , \7751 );
xor \U$7500 ( \7753 , \7726 , \7752 );
not \U$7501 ( \7754 , RIbe29fb0_79);
not \U$7502 ( \7755 , \1774 );
or \U$7503 ( \7756 , \7754 , \7755 );
nand \U$7504 ( \7757 , \429 , RIbe29e48_76);
nand \U$7505 ( \7758 , \7756 , \7757 );
and \U$7506 ( \7759 , \7758 , \1232 );
not \U$7507 ( \7760 , \7758 );
and \U$7508 ( \7761 , \7760 , \306 );
nor \U$7509 ( \7762 , \7759 , \7761 );
not \U$7510 ( \7763 , RIbe29dd0_75);
not \U$7511 ( \7764 , \3244 );
or \U$7512 ( \7765 , \7763 , \7764 );
nand \U$7513 ( \7766 , \1327 , RIbe29c68_72);
nand \U$7514 ( \7767 , \7765 , \7766 );
not \U$7515 ( \7768 , \7767 );
not \U$7516 ( \7769 , \424 );
and \U$7517 ( \7770 , \7768 , \7769 );
and \U$7518 ( \7771 , \7767 , \424 );
nor \U$7519 ( \7772 , \7770 , \7771 );
and \U$7520 ( \7773 , \7762 , \7772 );
not \U$7521 ( \7774 , \1611 );
not \U$7522 ( \7775 , RIbe28f48_44);
not \U$7523 ( \7776 , \7775 );
and \U$7524 ( \7777 , \7774 , \7776 );
and \U$7525 ( \7778 , \6760 , RIbe29bf0_71);
nor \U$7526 ( \7779 , \7777 , \7778 );
and \U$7527 ( \7780 , \7779 , \1618 );
not \U$7528 ( \7781 , \7779 );
and \U$7529 ( \7782 , \7781 , \3959 );
nor \U$7530 ( \7783 , \7780 , \7782 );
not \U$7531 ( \7784 , \7783 );
nor \U$7532 ( \7785 , \7773 , \7784 );
nor \U$7533 ( \7786 , \7762 , \7772 );
nor \U$7534 ( \7787 , \7785 , \7786 );
not \U$7535 ( \7788 , RIbe2b5b8_126);
not \U$7536 ( \7789 , \325 );
or \U$7537 ( \7790 , \7788 , \7789 );
nand \U$7538 ( \7791 , \329 , RIbe2a3e8_88);
nand \U$7539 ( \7792 , \7790 , \7791 );
not \U$7540 ( \7793 , \7792 );
not \U$7541 ( \7794 , \5151 );
and \U$7542 ( \7795 , \7793 , \7794 );
and \U$7543 ( \7796 , \7792 , \339 );
nor \U$7544 ( \7797 , \7795 , \7796 );
and \U$7545 ( \7798 , \1528 , RIbe2acd0_107);
and \U$7546 ( \7799 , \1531 , RIbe2a028_80);
nor \U$7547 ( \7800 , \7798 , \7799 );
and \U$7548 ( \7801 , \7800 , \293 );
not \U$7549 ( \7802 , \7800 );
and \U$7550 ( \7803 , \7802 , \300 );
nor \U$7551 ( \7804 , \7801 , \7803 );
and \U$7552 ( \7805 , \7797 , \7804 );
and \U$7553 ( \7806 , \260 , RIbe2a370_87);
and \U$7554 ( \7807 , \264 , RIbe2a2f8_86);
nor \U$7555 ( \7808 , \7806 , \7807 );
and \U$7556 ( \7809 , \7808 , \1362 );
not \U$7557 ( \7810 , \7808 );
and \U$7558 ( \7811 , \7810 , \1663 );
nor \U$7559 ( \7812 , \7809 , \7811 );
not \U$7560 ( \7813 , \7812 );
nor \U$7561 ( \7814 , \7805 , \7813 );
nor \U$7562 ( \7815 , \7797 , \7804 );
nor \U$7563 ( \7816 , \7814 , \7815 );
nand \U$7564 ( \7817 , \7787 , \7816 );
and \U$7565 ( \7818 , \2555 , RIbe287c8_28);
and \U$7566 ( \7819 , \1117 , RIbe28480_21);
nor \U$7567 ( \7820 , \7818 , \7819 );
and \U$7568 ( \7821 , \7820 , \1125 );
not \U$7569 ( \7822 , \7820 );
and \U$7570 ( \7823 , \7822 , \1131 );
nor \U$7571 ( \7824 , \7821 , \7823 );
not \U$7572 ( \7825 , \7824 );
not \U$7573 ( \7826 , RIbe28b10_35);
not \U$7574 ( \7827 , \2570 );
not \U$7575 ( \7828 , \7827 );
or \U$7576 ( \7829 , \7826 , \7828 );
nand \U$7577 ( \7830 , \2900 , RIbe28b88_36);
nand \U$7578 ( \7831 , \7829 , \7830 );
and \U$7579 ( \7832 , \7831 , \2573 );
not \U$7580 ( \7833 , \7831 );
and \U$7581 ( \7834 , \7833 , \2379 );
nor \U$7582 ( \7835 , \7832 , \7834 );
not \U$7583 ( \7836 , \7835 );
or \U$7584 ( \7837 , \7825 , \7836 );
or \U$7585 ( \7838 , \7835 , \7824 );
not \U$7586 ( \7839 , RIbe28408_20);
not \U$7587 ( \7840 , \2583 );
or \U$7588 ( \7841 , \7839 , \7840 );
nand \U$7589 ( \7842 , \2384 , RIbe28390_19);
nand \U$7590 ( \7843 , \7841 , \7842 );
not \U$7591 ( \7844 , \7843 );
not \U$7592 ( \7845 , \1076 );
and \U$7593 ( \7846 , \7844 , \7845 );
and \U$7594 ( \7847 , \7843 , \1076 );
nor \U$7595 ( \7848 , \7846 , \7847 );
not \U$7596 ( \7849 , \7848 );
nand \U$7597 ( \7850 , \7838 , \7849 );
nand \U$7598 ( \7851 , \7837 , \7850 );
not \U$7599 ( \7852 , \7851 );
not \U$7600 ( \7853 , \7852 );
not \U$7601 ( \7854 , RIbe29560_57);
not \U$7602 ( \7855 , \6413 );
or \U$7603 ( \7856 , \7854 , \7855 );
buf \U$7604 ( \7857 , \4312 );
buf \U$7605 ( \7858 , \7857 );
nand \U$7606 ( \7859 , \7858 , RIbe28228_16);
nand \U$7607 ( \7860 , \7856 , \7859 );
not \U$7608 ( \7861 , \7860 );
not \U$7609 ( \7862 , \4323 );
and \U$7610 ( \7863 , \7861 , \7862 );
not \U$7611 ( \7864 , \4322 );
not \U$7612 ( \7865 , \7864 );
and \U$7613 ( \7866 , \7860 , \7865 );
nor \U$7614 ( \7867 , \7863 , \7866 );
not \U$7615 ( \7868 , RIbe29290_51);
not \U$7616 ( \7869 , \3452 );
or \U$7617 ( \7870 , \7868 , \7869 );
nand \U$7618 ( \7871 , \3458 , RIbe28a20_33);
nand \U$7619 ( \7872 , \7870 , \7871 );
not \U$7620 ( \7873 , \7872 );
not \U$7621 ( \7874 , \2887 );
and \U$7622 ( \7875 , \7873 , \7874 );
and \U$7623 ( \7876 , \7872 , \3461 );
nor \U$7624 ( \7877 , \7875 , \7876 );
nand \U$7625 ( \7878 , \7867 , \7877 );
not \U$7626 ( \7879 , RIbe289a8_32);
not \U$7627 ( \7880 , \3703 );
not \U$7628 ( \7881 , \7880 );
or \U$7629 ( \7882 , \7879 , \7881 );
nand \U$7630 ( \7883 , \7438 , RIbe28930_31);
nand \U$7631 ( \7884 , \7882 , \7883 );
and \U$7632 ( \7885 , \7884 , \3471 );
not \U$7633 ( \7886 , \7884 );
and \U$7634 ( \7887 , \7886 , \3448 );
nor \U$7635 ( \7888 , \7885 , \7887 );
and \U$7636 ( \7889 , \7878 , \7888 );
nor \U$7637 ( \7890 , \7877 , \7867 );
nor \U$7638 ( \7891 , \7889 , \7890 );
not \U$7639 ( \7892 , \7891 );
or \U$7640 ( \7893 , \7853 , \7892 );
not \U$7641 ( \7894 , RIbe27f58_10);
not \U$7642 ( \7895 , \2597 );
or \U$7643 ( \7896 , \7894 , \7895 );
nand \U$7644 ( \7897 , \1147 , RIbe27e68_8);
nand \U$7645 ( \7898 , \7896 , \7897 );
not \U$7646 ( \7899 , \1152 );
and \U$7647 ( \7900 , \7898 , \7899 );
not \U$7648 ( \7901 , \7898 );
and \U$7649 ( \7902 , \7901 , \3994 );
nor \U$7650 ( \7903 , \7900 , \7902 );
and \U$7651 ( \7904 , \5973 , RIbe28ed0_43);
not \U$7652 ( \7905 , \1164 );
and \U$7653 ( \7906 , \7905 , RIbe27fd0_11);
nor \U$7654 ( \7907 , \7904 , \7906 );
and \U$7655 ( \7908 , \7907 , \750 );
not \U$7656 ( \7909 , \7907 );
and \U$7657 ( \7910 , \7909 , \1011 );
nor \U$7658 ( \7911 , \7908 , \7910 );
xor \U$7659 ( \7912 , \7903 , \7911 );
not \U$7660 ( \7913 , RIbe28660_25);
not \U$7661 ( \7914 , \1633 );
or \U$7662 ( \7915 , \7913 , \7914 );
nand \U$7663 ( \7916 , \1455 , RIbe285e8_24);
nand \U$7664 ( \7917 , \7915 , \7916 );
and \U$7665 ( \7918 , \7917 , \1309 );
not \U$7666 ( \7919 , \7917 );
and \U$7667 ( \7920 , \7919 , \1082 );
nor \U$7668 ( \7921 , \7918 , \7920 );
and \U$7669 ( \7922 , \7912 , \7921 );
and \U$7670 ( \7923 , \7903 , \7911 );
or \U$7671 ( \7924 , \7922 , \7923 );
nand \U$7672 ( \7925 , \7893 , \7924 );
not \U$7673 ( \7926 , \7891 );
nand \U$7674 ( \7927 , \7926 , \7851 );
nand \U$7675 ( \7928 , \7925 , \7927 );
xor \U$7676 ( \7929 , \7817 , \7928 );
not \U$7677 ( \7930 , RIbe28fc0_45);
not \U$7678 ( \7931 , \6535 );
or \U$7679 ( \7932 , \7930 , \7931 );
nand \U$7680 ( \7933 , \7075 , RIbe290b0_47);
nand \U$7681 ( \7934 , \7932 , \7933 );
not \U$7682 ( \7935 , \7546 );
and \U$7683 ( \7936 , \7934 , \7935 );
not \U$7684 ( \7937 , \7934 );
and \U$7685 ( \7938 , \7937 , \6548 );
nor \U$7686 ( \7939 , \7936 , \7938 );
not \U$7687 ( \7940 , RIbe29a88_68);
not \U$7688 ( \7941 , \6590 );
not \U$7689 ( \7942 , \7941 );
or \U$7690 ( \7943 , \7940 , \7942 );
nand \U$7691 ( \7944 , \6596 , RIbe27d78_6);
nand \U$7692 ( \7945 , \7943 , \7944 );
and \U$7693 ( \7946 , \7945 , \6601 );
not \U$7694 ( \7947 , \7945 );
buf \U$7695 ( \7948 , \6581 );
not \U$7696 ( \7949 , \7948 );
and \U$7697 ( \7950 , \7947 , \7949 );
nor \U$7698 ( \7951 , \7946 , \7950 );
xor \U$7699 ( \7952 , \7939 , \7951 );
not \U$7700 ( \7953 , RIbe27d00_5);
not \U$7701 ( \7954 , \6559 );
not \U$7702 ( \7955 , \7954 );
or \U$7703 ( \7956 , \7953 , \7955 );
not \U$7704 ( \7957 , \6556 );
buf \U$7705 ( \7958 , \7957 );
nand \U$7706 ( \7959 , \7958 , RIbe27c10_3);
nand \U$7707 ( \7960 , \7956 , \7959 );
and \U$7708 ( \7961 , \7960 , \7293 );
not \U$7709 ( \7962 , \7960 );
and \U$7710 ( \7963 , \7962 , \6572 );
nor \U$7711 ( \7964 , \7961 , \7963 );
and \U$7712 ( \7965 , \7952 , \7964 );
and \U$7713 ( \7966 , \7939 , \7951 );
or \U$7714 ( \7967 , \7965 , \7966 );
nand \U$7715 ( \7968 , RIbe2b2e8_120, RIbe2a4d8_90);
nand \U$7716 ( \7969 , \7968 , RIbe2b360_121);
not \U$7717 ( \7970 , \7969 );
not \U$7718 ( \7971 , \7970 );
not \U$7719 ( \7972 , \7971 );
not \U$7720 ( \7973 , RIbe29920_65);
not \U$7721 ( \7974 , \6941 );
buf \U$7722 ( \7975 , \7974 );
not \U$7723 ( \7976 , \7975 );
or \U$7724 ( \7977 , \7973 , \7976 );
xor \U$7725 ( \7978 , RIbe2a0a0_81, RIbe2b360_121);
not \U$7726 ( \7979 , \7978 );
buf \U$7727 ( \7980 , \7979 );
not \U$7728 ( \7981 , \7980 );
nand \U$7729 ( \7982 , \7981 , RIbe27b98_2);
nand \U$7730 ( \7983 , \7977 , \7982 );
buf \U$7731 ( \7984 , \6948 );
not \U$7732 ( \7985 , \7984 );
and \U$7733 ( \7986 , \7983 , \7985 );
not \U$7734 ( \7987 , \7983 );
not \U$7735 ( \7988 , \6948 );
not \U$7736 ( \7989 , \7988 );
and \U$7737 ( \7990 , \7987 , \7989 );
nor \U$7738 ( \7991 , \7986 , \7990 );
not \U$7739 ( \7992 , \7991 );
or \U$7740 ( \7993 , \7972 , \7992 );
not \U$7741 ( \7994 , \7991 );
nand \U$7742 ( \7995 , \7994 , \7970 );
not \U$7743 ( \7996 , RIbe28e58_42);
not \U$7744 ( \7997 , \7298 );
or \U$7745 ( \7998 , \7996 , \7997 );
nand \U$7746 ( \7999 , \6983 , RIbe28de0_41);
nand \U$7747 ( \8000 , \7998 , \7999 );
not \U$7748 ( \8001 , RIbe2a820_97);
not \U$7749 ( \8002 , RIbe2a118_82);
or \U$7750 ( \8003 , \8001 , \8002 );
nand \U$7751 ( \8004 , \8003 , RIbe2a898_98);
nor \U$7752 ( \8005 , \8000 , \8004 );
not \U$7753 ( \8006 , \8005 );
nand \U$7754 ( \8007 , \8000 , \7301 );
nand \U$7755 ( \8008 , \8006 , \8007 );
nand \U$7756 ( \8009 , \7995 , \8008 );
nand \U$7757 ( \8010 , \7993 , \8009 );
xor \U$7758 ( \8011 , \7967 , \8010 );
not \U$7759 ( \8012 , RIbe29650_59);
not \U$7760 ( \8013 , \6856 );
or \U$7761 ( \8014 , \8012 , \8013 );
nand \U$7762 ( \8015 , \6617 , RIbe29038_46);
nand \U$7763 ( \8016 , \8014 , \8015 );
and \U$7764 ( \8017 , \8016 , \7501 );
not \U$7765 ( \8018 , \8016 );
and \U$7766 ( \8019 , \8018 , \6624 );
nor \U$7767 ( \8020 , \8017 , \8019 );
not \U$7768 ( \8021 , \8020 );
not \U$7769 ( \8022 , RIbe281b0_15);
not \U$7770 ( \8023 , \5727 );
or \U$7771 ( \8024 , \8022 , \8023 );
nand \U$7772 ( \8025 , \5731 , RIbe280c0_13);
nand \U$7773 ( \8026 , \8024 , \8025 );
and \U$7774 ( \8027 , \8026 , \4586 );
not \U$7775 ( \8028 , \8026 );
and \U$7776 ( \8029 , \8028 , \4592 );
nor \U$7777 ( \8030 , \8027 , \8029 );
not \U$7778 ( \8031 , \8030 );
or \U$7779 ( \8032 , \8021 , \8031 );
or \U$7780 ( \8033 , \8030 , \8020 );
not \U$7781 ( \8034 , RIbe29830_63);
not \U$7782 ( \8035 , \5455 );
or \U$7783 ( \8036 , \8034 , \8035 );
nand \U$7784 ( \8037 , \6634 , RIbe296c8_60);
nand \U$7785 ( \8038 , \8036 , \8037 );
and \U$7786 ( \8039 , \8038 , \6641 );
not \U$7787 ( \8040 , \8038 );
and \U$7788 ( \8041 , \8040 , \6907 );
nor \U$7789 ( \8042 , \8039 , \8041 );
not \U$7790 ( \8043 , \8042 );
nand \U$7791 ( \8044 , \8033 , \8043 );
nand \U$7792 ( \8045 , \8032 , \8044 );
and \U$7793 ( \8046 , \8011 , \8045 );
and \U$7794 ( \8047 , \7967 , \8010 );
or \U$7795 ( \8048 , \8046 , \8047 );
xor \U$7796 ( \8049 , \7929 , \8048 );
nand \U$7797 ( \8050 , \7753 , \8049 );
and \U$7798 ( \8051 , \7804 , \7812 );
not \U$7799 ( \8052 , \7804 );
and \U$7800 ( \8053 , \8052 , \7813 );
or \U$7801 ( \8054 , \8051 , \8053 );
xor \U$7802 ( \8055 , \8054 , \7797 );
nand \U$7803 ( \8056 , RIbe29380_53, RIbe2a910_99);
nand \U$7804 ( \8057 , \8055 , \8056 );
not \U$7805 ( \8058 , \7772 );
not \U$7806 ( \8059 , \7783 );
or \U$7807 ( \8060 , \8058 , \8059 );
or \U$7808 ( \8061 , \7772 , \7783 );
nand \U$7809 ( \8062 , \8060 , \8061 );
not \U$7810 ( \8063 , \7762 );
and \U$7811 ( \8064 , \8062 , \8063 );
not \U$7812 ( \8065 , \8062 );
and \U$7813 ( \8066 , \8065 , \7762 );
nor \U$7814 ( \8067 , \8064 , \8066 );
and \U$7815 ( \8068 , \8057 , \8067 );
nor \U$7816 ( \8069 , \8055 , \8056 );
nor \U$7817 ( \8070 , \8068 , \8069 );
not \U$7818 ( \8071 , \8070 );
and \U$7819 ( \8072 , \8020 , \8042 );
not \U$7820 ( \8073 , \8020 );
and \U$7821 ( \8074 , \8073 , \8043 );
nor \U$7822 ( \8075 , \8072 , \8074 );
xor \U$7823 ( \8076 , \8075 , \8030 );
buf \U$7824 ( \8077 , \7969 );
xor \U$7825 ( \8078 , \8077 , \8008 );
xnor \U$7826 ( \8079 , \8078 , \7991 );
and \U$7827 ( \8080 , \8076 , \8079 );
xor \U$7828 ( \8081 , \7939 , \7951 );
xor \U$7829 ( \8082 , \8081 , \7964 );
not \U$7830 ( \8083 , \8082 );
nor \U$7831 ( \8084 , \8080 , \8083 );
nor \U$7832 ( \8085 , \8076 , \8079 );
nor \U$7833 ( \8086 , \8084 , \8085 );
not \U$7834 ( \8087 , \8086 );
or \U$7835 ( \8088 , \8071 , \8087 );
not \U$7836 ( \8089 , \7867 );
not \U$7837 ( \8090 , \7888 );
or \U$7838 ( \8091 , \8089 , \8090 );
or \U$7839 ( \8092 , \7888 , \7867 );
nand \U$7840 ( \8093 , \8091 , \8092 );
xor \U$7841 ( \8094 , \8093 , \7877 );
not \U$7842 ( \8095 , \8094 );
not \U$7843 ( \8096 , \8095 );
xor \U$7844 ( \8097 , \7903 , \7911 );
xor \U$7845 ( \8098 , \8097 , \7921 );
not \U$7846 ( \8099 , \8098 );
or \U$7847 ( \8100 , \8096 , \8099 );
not \U$7848 ( \8101 , \8094 );
not \U$7849 ( \8102 , \8098 );
not \U$7850 ( \8103 , \8102 );
or \U$7851 ( \8104 , \8101 , \8103 );
xor \U$7852 ( \8105 , \7848 , \7835 );
xor \U$7853 ( \8106 , \8105 , \7824 );
not \U$7854 ( \8107 , \8106 );
nand \U$7855 ( \8108 , \8104 , \8107 );
nand \U$7856 ( \8109 , \8100 , \8108 );
nand \U$7857 ( \8110 , \8088 , \8109 );
or \U$7858 ( \8111 , \8070 , \8086 );
nand \U$7859 ( \8112 , \8110 , \8111 );
not \U$7860 ( \8113 , \8112 );
and \U$7861 ( \8114 , RIbe29380_53, RIbe2a988_100);
not \U$7862 ( \8115 , \1362 );
not \U$7863 ( \8116 , RIbe2a3e8_88);
not \U$7864 ( \8117 , \260 );
or \U$7865 ( \8118 , \8116 , \8117 );
nand \U$7866 ( \8119 , \263 , RIbe2a370_87);
nand \U$7867 ( \8120 , \8118 , \8119 );
not \U$7868 ( \8121 , \8120 );
or \U$7869 ( \8122 , \8115 , \8121 );
or \U$7870 ( \8123 , \8120 , \1362 );
nand \U$7871 ( \8124 , \8122 , \8123 );
not \U$7872 ( \8125 , RIbe2a910_99);
not \U$7873 ( \8126 , \324 );
or \U$7874 ( \8127 , \8125 , \8126 );
nand \U$7875 ( \8128 , \330 , RIbe2b5b8_126);
nand \U$7876 ( \8129 , \8127 , \8128 );
xnor \U$7877 ( \8130 , \8129 , \1374 );
xor \U$7878 ( \8131 , \8124 , \8130 );
not \U$7879 ( \8132 , \300 );
not \U$7880 ( \8133 , RIbe2a2f8_86);
not \U$7881 ( \8134 , \1528 );
or \U$7882 ( \8135 , \8133 , \8134 );
nand \U$7883 ( \8136 , \1531 , RIbe2acd0_107);
nand \U$7884 ( \8137 , \8135 , \8136 );
not \U$7885 ( \8138 , \8137 );
or \U$7886 ( \8139 , \8132 , \8138 );
or \U$7887 ( \8140 , \8137 , \300 );
nand \U$7888 ( \8141 , \8139 , \8140 );
and \U$7889 ( \8142 , \8131 , \8141 );
and \U$7890 ( \8143 , \8124 , \8130 );
or \U$7891 ( \8144 , \8142 , \8143 );
xor \U$7892 ( \8145 , \8114 , \8144 );
not \U$7893 ( \8146 , RIbe29e48_76);
not \U$7894 ( \8147 , \1237 );
or \U$7895 ( \8148 , \8146 , \8147 );
nand \U$7896 ( \8149 , \553 , RIbe29dd0_75);
nand \U$7897 ( \8150 , \8148 , \8149 );
not \U$7898 ( \8151 , \8150 );
not \U$7899 ( \8152 , \424 );
and \U$7900 ( \8153 , \8151 , \8152 );
and \U$7901 ( \8154 , \8150 , \424 );
nor \U$7902 ( \8155 , \8153 , \8154 );
not \U$7903 ( \8156 , \8155 );
not \U$7904 ( \8157 , \8156 );
not \U$7905 ( \8158 , RIbe2a028_80);
not \U$7906 ( \8159 , \1337 );
or \U$7907 ( \8160 , \8158 , \8159 );
nand \U$7908 ( \8161 , \429 , RIbe29fb0_79);
nand \U$7909 ( \8162 , \8160 , \8161 );
and \U$7910 ( \8163 , \8162 , \1547 );
not \U$7911 ( \8164 , \8162 );
and \U$7912 ( \8165 , \8164 , \306 );
nor \U$7913 ( \8166 , \8163 , \8165 );
not \U$7914 ( \8167 , \8166 );
not \U$7915 ( \8168 , \8167 );
or \U$7916 ( \8169 , \8157 , \8168 );
not \U$7917 ( \8170 , \8166 );
not \U$7918 ( \8171 , \8155 );
or \U$7919 ( \8172 , \8170 , \8171 );
not \U$7920 ( \8173 , \740 );
not \U$7921 ( \8174 , \8173 );
not \U$7922 ( \8175 , RIbe29bf0_71);
not \U$7923 ( \8176 , \8175 );
and \U$7924 ( \8177 , \8174 , \8176 );
and \U$7925 ( \8178 , \7363 , RIbe29c68_72);
nor \U$7926 ( \8179 , \8177 , \8178 );
and \U$7927 ( \8180 , \8179 , \564 );
not \U$7928 ( \8181 , \8179 );
and \U$7929 ( \8182 , \8181 , \1621 );
nor \U$7930 ( \8183 , \8180 , \8182 );
nand \U$7931 ( \8184 , \8172 , \8183 );
nand \U$7932 ( \8185 , \8169 , \8184 );
and \U$7933 ( \8186 , \8145 , \8185 );
and \U$7934 ( \8187 , \8114 , \8144 );
or \U$7935 ( \8188 , \8186 , \8187 );
not \U$7936 ( \8189 , RIbe290b0_47);
not \U$7937 ( \8190 , \7274 );
or \U$7938 ( \8191 , \8189 , \8190 );
nand \U$7939 ( \8192 , \6596 , RIbe29a88_68);
nand \U$7940 ( \8193 , \8191 , \8192 );
and \U$7941 ( \8194 , \8193 , \6873 );
not \U$7942 ( \8195 , \8193 );
and \U$7943 ( \8196 , \8195 , \6582 );
nor \U$7944 ( \8197 , \8194 , \8196 );
not \U$7945 ( \8198 , RIbe27d78_6);
not \U$7946 ( \8199 , \6559 );
not \U$7947 ( \8200 , \8199 );
or \U$7948 ( \8201 , \8198 , \8200 );
buf \U$7949 ( \8202 , \6962 );
nand \U$7950 ( \8203 , \8202 , RIbe27d00_5);
nand \U$7951 ( \8204 , \8201 , \8203 );
and \U$7952 ( \8205 , \8204 , \6572 );
not \U$7953 ( \8206 , \8204 );
and \U$7954 ( \8207 , \8206 , \7293 );
nor \U$7955 ( \8208 , \8205 , \8207 );
and \U$7956 ( \8209 , \8197 , \8208 );
not \U$7957 ( \8210 , RIbe29038_46);
not \U$7958 ( \8211 , \6880 );
or \U$7959 ( \8212 , \8210 , \8211 );
nand \U$7960 ( \8213 , \6540 , RIbe28fc0_45);
nand \U$7961 ( \8214 , \8212 , \8213 );
not \U$7962 ( \8215 , \8214 );
not \U$7963 ( \8216 , \7546 );
and \U$7964 ( \8217 , \8215 , \8216 );
and \U$7965 ( \8218 , \8214 , \6888 );
nor \U$7966 ( \8219 , \8217 , \8218 );
nor \U$7967 ( \8220 , \8209 , \8219 );
nor \U$7968 ( \8221 , \8197 , \8208 );
nor \U$7969 ( \8222 , \8220 , \8221 );
not \U$7970 ( \8223 , \8222 );
not \U$7971 ( \8224 , RIbe28228_16);
not \U$7972 ( \8225 , \5727 );
or \U$7973 ( \8226 , \8224 , \8225 );
nand \U$7974 ( \8227 , \5052 , RIbe281b0_15);
nand \U$7975 ( \8228 , \8226 , \8227 );
xor \U$7976 ( \8229 , \8228 , \4946 );
not \U$7977 ( \8230 , RIbe296c8_60);
buf \U$7978 ( \8231 , \6138 );
not \U$7979 ( \8232 , \8231 );
or \U$7980 ( \8233 , \8230 , \8232 );
not \U$7981 ( \8234 , \6614 );
buf \U$7982 ( \8235 , \8234 );
nand \U$7983 ( \8236 , \8235 , RIbe29650_59);
nand \U$7984 ( \8237 , \8233 , \8236 );
and \U$7985 ( \8238 , \8237 , \5740 );
not \U$7986 ( \8239 , \8237 );
and \U$7987 ( \8240 , \8239 , \7501 );
nor \U$7988 ( \8241 , \8238 , \8240 );
and \U$7989 ( \8242 , \8229 , \8241 );
not \U$7990 ( \8243 , RIbe280c0_13);
not \U$7991 ( \8244 , \5455 );
or \U$7992 ( \8245 , \8243 , \8244 );
not \U$7993 ( \8246 , \7098 );
buf \U$7994 ( \8247 , \8246 );
nand \U$7995 ( \8248 , \8247 , RIbe29830_63);
nand \U$7996 ( \8249 , \8245 , \8248 );
and \U$7997 ( \8250 , \8249 , \5046 );
not \U$7998 ( \8251 , \8249 );
not \U$7999 ( \8252 , \5045 );
not \U$8000 ( \8253 , \8252 );
and \U$8001 ( \8254 , \8251 , \8253 );
nor \U$8002 ( \8255 , \8250 , \8254 );
nor \U$8003 ( \8256 , \8242 , \8255 );
not \U$8004 ( \8257 , \8228 );
not \U$8005 ( \8258 , \4946 );
and \U$8006 ( \8259 , \8257 , \8258 );
and \U$8007 ( \8260 , \8228 , \4946 );
nor \U$8008 ( \8261 , \8259 , \8260 );
nor \U$8009 ( \8262 , \8261 , \8241 );
nor \U$8010 ( \8263 , \8256 , \8262 );
not \U$8011 ( \8264 , \8263 );
or \U$8012 ( \8265 , \8223 , \8264 );
not \U$8013 ( \8266 , RIbe28de0_41);
not \U$8014 ( \8267 , \7975 );
or \U$8015 ( \8268 , \8266 , \8267 );
not \U$8016 ( \8269 , \7980 );
nand \U$8017 ( \8270 , \8269 , RIbe29920_65);
nand \U$8018 ( \8271 , \8268 , \8270 );
xor \U$8019 ( \8272 , \8271 , \7984 );
xnor \U$8020 ( \8273 , RIbe2b360_121, RIbe2b2e8_120);
xor \U$8021 ( \8274 , RIbe2b2e8_120, RIbe2a4d8_90);
nor \U$8022 ( \8275 , \8273 , \8274 );
buf \U$8023 ( \8276 , \8275 );
not \U$8024 ( \8277 , \8276 );
not \U$8025 ( \8278 , \8277 );
nand \U$8026 ( \8279 , \8278 , RIbe27b98_2);
and \U$8027 ( \8280 , \8279 , \8077 );
not \U$8028 ( \8281 , \8279 );
and \U$8029 ( \8282 , \8281 , \7970 );
or \U$8030 ( \8283 , \8280 , \8282 );
and \U$8031 ( \8284 , \8272 , \8283 );
and \U$8032 ( \8285 , \7299 , RIbe27c10_3);
not \U$8033 ( \8286 , \6983 );
not \U$8034 ( \8287 , \8286 );
not \U$8035 ( \8288 , \8287 );
nor \U$8036 ( \8289 , \8288 , \3299 );
nor \U$8037 ( \8290 , \8285 , \8289 );
and \U$8038 ( \8291 , \8290 , \6993 );
not \U$8039 ( \8292 , \8290 );
and \U$8040 ( \8293 , \8292 , \7661 );
nor \U$8041 ( \8294 , \8291 , \8293 );
nor \U$8042 ( \8295 , \8284 , \8294 );
nor \U$8043 ( \8296 , \8272 , \8283 );
nor \U$8044 ( \8297 , \8295 , \8296 );
not \U$8045 ( \8298 , \8297 );
nand \U$8046 ( \8299 , \8265 , \8298 );
or \U$8047 ( \8300 , \8263 , \8222 );
nand \U$8048 ( \8301 , \8299 , \8300 );
xor \U$8049 ( \8302 , \8188 , \8301 );
and \U$8050 ( \8303 , \5973 , RIbe28f48_44);
and \U$8051 ( \8304 , \1203 , RIbe28ed0_43);
nor \U$8052 ( \8305 , \8303 , \8304 );
and \U$8053 ( \8306 , \8305 , \750 );
not \U$8054 ( \8307 , \8305 );
and \U$8055 ( \8308 , \8307 , \1011 );
nor \U$8056 ( \8309 , \8306 , \8308 );
not \U$8057 ( \8310 , RIbe27e68_8);
not \U$8058 ( \8311 , \1298 );
or \U$8059 ( \8312 , \8310 , \8311 );
nand \U$8060 ( \8313 , \1454 , RIbe28660_25);
nand \U$8061 ( \8314 , \8312 , \8313 );
and \U$8062 ( \8315 , \8314 , \1309 );
not \U$8063 ( \8316 , \8314 );
and \U$8064 ( \8317 , \8316 , \5125 );
nor \U$8065 ( \8318 , \8315 , \8317 );
or \U$8066 ( \8319 , \8309 , \8318 );
not \U$8067 ( \8320 , RIbe27fd0_11);
not \U$8068 ( \8321 , \1143 );
or \U$8069 ( \8322 , \8320 , \8321 );
nand \U$8070 ( \8323 , \1147 , RIbe27f58_10);
nand \U$8071 ( \8324 , \8322 , \8323 );
and \U$8072 ( \8325 , \8324 , \1469 );
not \U$8073 ( \8326 , \8324 );
not \U$8074 ( \8327 , \7899 );
and \U$8075 ( \8328 , \8326 , \8327 );
nor \U$8076 ( \8329 , \8325 , \8328 );
nand \U$8077 ( \8330 , \8319 , \8329 );
nand \U$8078 ( \8331 , \8318 , \8309 );
nand \U$8079 ( \8332 , \8330 , \8331 );
and \U$8080 ( \8333 , \1113 , RIbe285e8_24);
and \U$8081 ( \8334 , \1117 , RIbe287c8_28);
nor \U$8082 ( \8335 , \8333 , \8334 );
and \U$8083 ( \8336 , \8335 , \1125 );
not \U$8084 ( \8337 , \8335 );
and \U$8085 ( \8338 , \8337 , \1131 );
nor \U$8086 ( \8339 , \8336 , \8338 );
not \U$8087 ( \8340 , \8339 );
not \U$8088 ( \8341 , RIbe28390_19);
not \U$8089 ( \8342 , \2570 );
not \U$8090 ( \8343 , \8342 );
or \U$8091 ( \8344 , \8341 , \8343 );
nand \U$8092 ( \8345 , \4284 , RIbe28b10_35);
nand \U$8093 ( \8346 , \8344 , \8345 );
and \U$8094 ( \8347 , \8346 , \7457 );
not \U$8095 ( \8348 , \8346 );
and \U$8096 ( \8349 , \8348 , \4783 );
nor \U$8097 ( \8350 , \8347 , \8349 );
not \U$8098 ( \8351 , \8350 );
or \U$8099 ( \8352 , \8340 , \8351 );
or \U$8100 ( \8353 , \8350 , \8339 );
not \U$8101 ( \8354 , RIbe28480_21);
not \U$8102 ( \8355 , \2583 );
or \U$8103 ( \8356 , \8354 , \8355 );
nand \U$8104 ( \8357 , \2384 , RIbe28408_20);
nand \U$8105 ( \8358 , \8356 , \8357 );
xor \U$8106 ( \8359 , \8358 , \1076 );
not \U$8107 ( \8360 , \8359 );
nand \U$8108 ( \8361 , \8353 , \8360 );
nand \U$8109 ( \8362 , \8352 , \8361 );
xor \U$8110 ( \8363 , \8332 , \8362 );
not \U$8111 ( \8364 , RIbe28a20_33);
not \U$8112 ( \8365 , \4021 );
or \U$8113 ( \8366 , \8364 , \8365 );
buf \U$8114 ( \8367 , \4025 );
not \U$8115 ( \8368 , \8367 );
nand \U$8116 ( \8369 , \8368 , RIbe289a8_32);
nand \U$8117 ( \8370 , \8366 , \8369 );
and \U$8118 ( \8371 , \8370 , \3471 );
not \U$8119 ( \8372 , \8370 );
and \U$8120 ( \8373 , \8372 , \3448 );
nor \U$8121 ( \8374 , \8371 , \8373 );
not \U$8122 ( \8375 , RIbe28b88_36);
not \U$8123 ( \8376 , \3284 );
or \U$8124 ( \8377 , \8375 , \8376 );
nand \U$8125 ( \8378 , \4011 , RIbe29290_51);
nand \U$8126 ( \8379 , \8377 , \8378 );
and \U$8127 ( \8380 , \8379 , \4346 );
not \U$8128 ( \8381 , \8379 );
and \U$8129 ( \8382 , \8381 , \3461 );
nor \U$8130 ( \8383 , \8380 , \8382 );
xor \U$8131 ( \8384 , \8374 , \8383 );
not \U$8132 ( \8385 , RIbe28930_31);
not \U$8133 ( \8386 , \5058 );
or \U$8134 ( \8387 , \8385 , \8386 );
nand \U$8135 ( \8388 , \4600 , RIbe29560_57);
nand \U$8136 ( \8389 , \8387 , \8388 );
and \U$8137 ( \8390 , \8389 , \4007 );
not \U$8138 ( \8391 , \8389 );
and \U$8139 ( \8392 , \8391 , \4323 );
nor \U$8140 ( \8393 , \8390 , \8392 );
and \U$8141 ( \8394 , \8384 , \8393 );
and \U$8142 ( \8395 , \8374 , \8383 );
or \U$8143 ( \8396 , \8394 , \8395 );
and \U$8144 ( \8397 , \8363 , \8396 );
and \U$8145 ( \8398 , \8332 , \8362 );
or \U$8146 ( \8399 , \8397 , \8398 );
and \U$8147 ( \8400 , \8302 , \8399 );
and \U$8148 ( \8401 , \8188 , \8301 );
or \U$8149 ( \8402 , \8400 , \8401 );
not \U$8150 ( \8403 , \8402 );
and \U$8151 ( \8404 , \8113 , \8403 );
not \U$8152 ( \8405 , \7750 );
not \U$8153 ( \8406 , \8405 );
not \U$8154 ( \8407 , \7738 );
or \U$8155 ( \8408 , \8406 , \8407 );
nand \U$8156 ( \8409 , \7737 , \7750 );
nand \U$8157 ( \8410 , \8408 , \8409 );
and \U$8158 ( \8411 , \8410 , \7728 );
not \U$8159 ( \8412 , \8410 );
and \U$8160 ( \8413 , \8412 , \7729 );
nor \U$8161 ( \8414 , \8411 , \8413 );
not \U$8162 ( \8415 , \7691 );
xor \U$8163 ( \8416 , \7699 , \8415 );
buf \U$8164 ( \8417 , \8416 );
nand \U$8165 ( \8418 , \8414 , \8417 );
not \U$8166 ( \8419 , \7723 );
not \U$8167 ( \8420 , \8419 );
not \U$8168 ( \8421 , \7702 );
not \U$8169 ( \8422 , \7713 );
or \U$8170 ( \8423 , \8421 , \8422 );
or \U$8171 ( \8424 , \7713 , \7702 );
nand \U$8172 ( \8425 , \8423 , \8424 );
not \U$8173 ( \8426 , \8425 );
or \U$8174 ( \8427 , \8420 , \8426 );
or \U$8175 ( \8428 , \8425 , \8419 );
nand \U$8176 ( \8429 , \8427 , \8428 );
and \U$8177 ( \8430 , \8418 , \8429 );
nor \U$8178 ( \8431 , \8414 , \8417 );
nor \U$8179 ( \8432 , \8430 , \8431 );
nor \U$8180 ( \8433 , \8404 , \8432 );
and \U$8181 ( \8434 , \8112 , \8402 );
nor \U$8182 ( \8435 , \8433 , \8434 );
xor \U$8183 ( \8436 , \8050 , \8435 );
not \U$8184 ( \8437 , \6999 );
not \U$8185 ( \8438 , \6897 );
or \U$8186 ( \8439 , \8437 , \8438 );
not \U$8187 ( \8440 , \6999 );
nand \U$8188 ( \8441 , \8440 , \6898 );
nand \U$8189 ( \8442 , \8439 , \8441 );
and \U$8190 ( \8443 , \8442 , \6933 );
not \U$8191 ( \8444 , \8442 );
and \U$8192 ( \8445 , \8444 , \6932 );
nor \U$8193 ( \8446 , \8443 , \8445 );
xor \U$8194 ( \8447 , \6850 , \6810 );
xor \U$8195 ( \8448 , \8447 , \6770 );
xor \U$8196 ( \8449 , \8446 , \8448 );
and \U$8197 ( \8450 , \6710 , \6679 );
not \U$8198 ( \8451 , \6710 );
and \U$8199 ( \8452 , \8451 , \6680 );
nor \U$8200 ( \8453 , \8450 , \8452 );
xnor \U$8201 ( \8454 , \8453 , \6735 );
xnor \U$8202 ( \8455 , \8449 , \8454 );
or \U$8203 ( \8456 , \7816 , \7787 );
nand \U$8204 ( \8457 , \8456 , \7817 );
and \U$8205 ( \8458 , \7891 , \7852 );
not \U$8206 ( \8459 , \7891 );
and \U$8207 ( \8460 , \8459 , \7851 );
or \U$8208 ( \8461 , \8458 , \8460 );
xnor \U$8209 ( \8462 , \8461 , \7924 );
xor \U$8210 ( \8463 , \8457 , \8462 );
xor \U$8211 ( \8464 , \7967 , \8010 );
xor \U$8212 ( \8465 , \8464 , \8045 );
and \U$8213 ( \8466 , \8463 , \8465 );
and \U$8214 ( \8467 , \8457 , \8462 );
or \U$8215 ( \8468 , \8466 , \8467 );
not \U$8216 ( \8469 , \8468 );
nand \U$8217 ( \8470 , \8455 , \8469 );
not \U$8218 ( \8471 , RIbe29920_65);
not \U$8219 ( \8472 , \7299 );
or \U$8220 ( \8473 , \8471 , \8472 );
nand \U$8221 ( \8474 , \6985 , RIbe27b98_2);
nand \U$8222 ( \8475 , \8473 , \8474 );
and \U$8223 ( \8476 , \8475 , \6993 );
not \U$8224 ( \8477 , \8475 );
and \U$8225 ( \8478 , \8477 , \7301 );
nor \U$8226 ( \8479 , \8476 , \8478 );
not \U$8227 ( \8480 , \6949 );
and \U$8228 ( \8481 , \8479 , \8480 );
not \U$8229 ( \8482 , \8479 );
and \U$8230 ( \8483 , \8482 , \7989 );
nor \U$8231 ( \8484 , \8481 , \8483 );
not \U$8232 ( \8485 , \8484 );
not \U$8233 ( \8486 , RIbe28e58_42);
not \U$8234 ( \8487 , \6561 );
or \U$8235 ( \8488 , \8486 , \8487 );
nand \U$8236 ( \8489 , \7653 , RIbe28de0_41);
nand \U$8237 ( \8490 , \8488 , \8489 );
xor \U$8238 ( \8491 , \8490 , \6572 );
not \U$8239 ( \8492 , \8491 );
not \U$8240 ( \8493 , \8492 );
and \U$8241 ( \8494 , \8485 , \8493 );
and \U$8242 ( \8495 , \8484 , \8492 );
nor \U$8243 ( \8496 , \8494 , \8495 );
xor \U$8244 ( \8497 , \7347 , \7378 );
xor \U$8245 ( \8498 , \8497 , \7381 );
xor \U$8246 ( \8499 , \8496 , \8498 );
not \U$8247 ( \8500 , \7464 );
not \U$8248 ( \8501 , \7510 );
not \U$8249 ( \8502 , \8501 );
or \U$8250 ( \8503 , \8500 , \8502 );
nand \U$8251 ( \8504 , \7513 , \7510 );
nand \U$8252 ( \8505 , \8503 , \8504 );
and \U$8253 ( \8506 , \8505 , \7422 );
not \U$8254 ( \8507 , \8505 );
and \U$8255 ( \8508 , \8507 , \7514 );
nor \U$8256 ( \8509 , \8506 , \8508 );
xor \U$8257 ( \8510 , \8499 , \8509 );
not \U$8258 ( \8511 , \8510 );
and \U$8259 ( \8512 , \8470 , \8511 );
nor \U$8260 ( \8513 , \8455 , \8469 );
nor \U$8261 ( \8514 , \8512 , \8513 );
and \U$8262 ( \8515 , \8436 , \8514 );
and \U$8263 ( \8516 , \8050 , \8435 );
or \U$8264 ( \8517 , \8515 , \8516 );
not \U$8265 ( \8518 , \8517 );
not \U$8266 ( \8519 , \7004 );
not \U$8267 ( \8520 , \7520 );
or \U$8268 ( \8521 , \8519 , \8520 );
or \U$8269 ( \8522 , \7004 , \7520 );
nand \U$8270 ( \8523 , \8521 , \8522 );
not \U$8271 ( \8524 , \8523 );
not \U$8272 ( \8525 , \7268 );
and \U$8273 ( \8526 , \8524 , \8525 );
and \U$8274 ( \8527 , \7268 , \8523 );
nor \U$8275 ( \8528 , \8526 , \8527 );
not \U$8276 ( \8529 , \8528 );
not \U$8277 ( \8530 , \7112 );
not \U$8278 ( \8531 , \7147 );
or \U$8279 ( \8532 , \8530 , \8531 );
nand \U$8280 ( \8533 , \8532 , \7166 );
nand \U$8281 ( \8534 , \7150 , \7113 );
nand \U$8282 ( \8535 , \8533 , \8534 );
xor \U$8283 ( \8536 , \7326 , \7336 );
and \U$8284 ( \8537 , \8536 , \7346 );
and \U$8285 ( \8538 , \7326 , \7336 );
or \U$8286 ( \8539 , \8537 , \8538 );
not \U$8287 ( \8540 , \8539 );
and \U$8288 ( \8541 , \7459 , \7433 );
nor \U$8289 ( \8542 , \8541 , \7444 );
nor \U$8290 ( \8543 , \7459 , \7433 );
nor \U$8291 ( \8544 , \8542 , \8543 );
not \U$8292 ( \8545 , \8544 );
or \U$8293 ( \8546 , \8540 , \8545 );
xor \U$8294 ( \8547 , \7358 , \7369 );
and \U$8295 ( \8548 , \8547 , \7377 );
and \U$8296 ( \8549 , \7358 , \7369 );
or \U$8297 ( \8550 , \8548 , \8549 );
nand \U$8298 ( \8551 , \8546 , \8550 );
not \U$8299 ( \8552 , \8544 );
not \U$8300 ( \8553 , \8539 );
nand \U$8301 ( \8554 , \8552 , \8553 );
nand \U$8302 ( \8555 , \8551 , \8554 );
xor \U$8303 ( \8556 , \8535 , \8555 );
not \U$8304 ( \8557 , \7989 );
not \U$8305 ( \8558 , \8492 );
or \U$8306 ( \8559 , \8557 , \8558 );
not \U$8307 ( \8560 , \8491 );
not \U$8308 ( \8561 , \8480 );
or \U$8309 ( \8562 , \8560 , \8561 );
nand \U$8310 ( \8563 , \8562 , \8479 );
nand \U$8311 ( \8564 , \8559 , \8563 );
not \U$8312 ( \8565 , \7505 );
not \U$8313 ( \8566 , \7490 );
or \U$8314 ( \8567 , \8565 , \8566 );
or \U$8315 ( \8568 , \7490 , \7505 );
nand \U$8316 ( \8569 , \8568 , \7477 );
nand \U$8317 ( \8570 , \8567 , \8569 );
xor \U$8318 ( \8571 , \8564 , \8570 );
not \U$8319 ( \8572 , \7421 );
not \U$8320 ( \8573 , \7407 );
not \U$8321 ( \8574 , \8573 );
or \U$8322 ( \8575 , \8572 , \8574 );
or \U$8323 ( \8576 , \8573 , \7421 );
nand \U$8324 ( \8577 , \8576 , \7396 );
nand \U$8325 ( \8578 , \8575 , \8577 );
and \U$8326 ( \8579 , \8571 , \8578 );
and \U$8327 ( \8580 , \8564 , \8570 );
or \U$8328 ( \8581 , \8579 , \8580 );
xor \U$8329 ( \8582 , \8556 , \8581 );
not \U$8330 ( \8583 , \8582 );
and \U$8331 ( \8584 , \8529 , \8583 );
and \U$8332 ( \8585 , \8528 , \8582 );
nor \U$8333 ( \8586 , \8584 , \8585 );
not \U$8334 ( \8587 , \8586 );
xor \U$8335 ( \8588 , \7583 , \7636 );
xor \U$8336 ( \8589 , \8588 , \7682 );
not \U$8337 ( \8590 , \8589 );
and \U$8338 ( \8591 , \8587 , \8590 );
and \U$8339 ( \8592 , \8586 , \8589 );
nor \U$8340 ( \8593 , \8591 , \8592 );
not \U$8341 ( \8594 , \8593 );
or \U$8342 ( \8595 , \8518 , \8594 );
xor \U$8343 ( \8596 , \8544 , \8553 );
xor \U$8344 ( \8597 , \8596 , \8550 );
not \U$8345 ( \8598 , \8597 );
xor \U$8346 ( \8599 , \8564 , \8570 );
xor \U$8347 ( \8600 , \8599 , \8578 );
not \U$8348 ( \8601 , \8600 );
and \U$8349 ( \8602 , \8598 , \8601 );
and \U$8350 ( \8603 , \8597 , \8600 );
nor \U$8351 ( \8604 , \8602 , \8603 );
not \U$8352 ( \8605 , \8604 );
not \U$8353 ( \8606 , \8454 );
buf \U$8354 ( \8607 , \8446 );
not \U$8355 ( \8608 , \8607 );
or \U$8356 ( \8609 , \8606 , \8608 );
or \U$8357 ( \8610 , \8607 , \8454 );
nand \U$8358 ( \8611 , \8610 , \8448 );
nand \U$8359 ( \8612 , \8609 , \8611 );
not \U$8360 ( \8613 , \8612 );
or \U$8361 ( \8614 , \8605 , \8613 );
or \U$8362 ( \8615 , \8612 , \8604 );
nand \U$8363 ( \8616 , \8614 , \8615 );
not \U$8364 ( \8617 , \8616 );
xor \U$8365 ( \8618 , \8496 , \8498 );
and \U$8366 ( \8619 , \8618 , \8509 );
and \U$8367 ( \8620 , \8496 , \8498 );
or \U$8368 ( \8621 , \8619 , \8620 );
not \U$8369 ( \8622 , \8621 );
xor \U$8370 ( \8623 , \7700 , \7725 );
and \U$8371 ( \8624 , \8623 , \7752 );
and \U$8372 ( \8625 , \7700 , \7725 );
or \U$8373 ( \8626 , \8624 , \8625 );
not \U$8374 ( \8627 , \8626 );
xor \U$8375 ( \8628 , \7817 , \7928 );
and \U$8376 ( \8629 , \8628 , \8048 );
and \U$8377 ( \8630 , \7817 , \7928 );
or \U$8378 ( \8631 , \8629 , \8630 );
not \U$8379 ( \8632 , \8631 );
not \U$8380 ( \8633 , \8632 );
and \U$8381 ( \8634 , \8627 , \8633 );
and \U$8382 ( \8635 , \8626 , \8632 );
nor \U$8383 ( \8636 , \8634 , \8635 );
not \U$8384 ( \8637 , \8636 );
not \U$8385 ( \8638 , \8637 );
or \U$8386 ( \8639 , \8622 , \8638 );
not \U$8387 ( \8640 , \8621 );
nand \U$8388 ( \8641 , \8640 , \8636 );
nand \U$8389 ( \8642 , \8639 , \8641 );
not \U$8390 ( \8643 , \8642 );
or \U$8391 ( \8644 , \8617 , \8643 );
or \U$8392 ( \8645 , \8616 , \8642 );
not \U$8393 ( \8646 , \6737 );
not \U$8394 ( \8647 , \8646 );
xor \U$8395 ( \8648 , \7001 , \6852 );
not \U$8396 ( \8649 , \8648 );
or \U$8397 ( \8650 , \8647 , \8649 );
or \U$8398 ( \8651 , \8648 , \8646 );
nand \U$8399 ( \8652 , \8650 , \8651 );
xor \U$8400 ( \8653 , \7308 , \7383 );
xnor \U$8401 ( \8654 , \8653 , \7516 );
xor \U$8402 ( \8655 , \8652 , \8654 );
xor \U$8403 ( \8656 , \7167 , \7108 );
xnor \U$8404 ( \8657 , \8656 , \7265 );
xor \U$8405 ( \8658 , \8655 , \8657 );
nand \U$8406 ( \8659 , \8645 , \8658 );
nand \U$8407 ( \8660 , \8644 , \8659 );
nand \U$8408 ( \8661 , \8595 , \8660 );
not \U$8409 ( \8662 , \8517 );
not \U$8410 ( \8663 , \8593 );
nand \U$8411 ( \8664 , \8662 , \8663 );
nand \U$8412 ( \8665 , \8661 , \8664 );
or \U$8413 ( \8666 , \7686 , \8665 );
not \U$8414 ( \8667 , \8600 );
nand \U$8415 ( \8668 , \8667 , \8597 );
and \U$8416 ( \8669 , \8612 , \8668 );
not \U$8417 ( \8670 , \8600 );
nor \U$8418 ( \8671 , \8670 , \8597 );
nor \U$8419 ( \8672 , \8669 , \8671 );
not \U$8420 ( \8673 , \8672 );
not \U$8421 ( \8674 , \8673 );
not \U$8422 ( \8675 , \8626 );
and \U$8423 ( \8676 , \8675 , \8632 );
nor \U$8424 ( \8677 , \8676 , \8621 );
nor \U$8425 ( \8678 , \8675 , \8632 );
nor \U$8426 ( \8679 , \8677 , \8678 );
not \U$8427 ( \8680 , \8679 );
not \U$8428 ( \8681 , \8680 );
or \U$8429 ( \8682 , \8674 , \8681 );
not \U$8430 ( \8683 , \8679 );
not \U$8431 ( \8684 , \8672 );
or \U$8432 ( \8685 , \8683 , \8684 );
xor \U$8433 ( \8686 , \8652 , \8654 );
and \U$8434 ( \8687 , \8686 , \8657 );
and \U$8435 ( \8688 , \8652 , \8654 );
or \U$8436 ( \8689 , \8687 , \8688 );
nand \U$8437 ( \8690 , \8685 , \8689 );
nand \U$8438 ( \8691 , \8682 , \8690 );
not \U$8439 ( \8692 , \8582 );
nand \U$8440 ( \8693 , \8692 , \8528 );
not \U$8441 ( \8694 , \8693 );
not \U$8442 ( \8695 , \8589 );
or \U$8443 ( \8696 , \8694 , \8695 );
not \U$8444 ( \8697 , \8528 );
nand \U$8445 ( \8698 , \8697 , \8582 );
nand \U$8446 ( \8699 , \8696 , \8698 );
xor \U$8447 ( \8700 , \8691 , \8699 );
xor \U$8448 ( \8701 , \7590 , \7165 );
and \U$8449 ( \8702 , \8701 , \7595 );
and \U$8450 ( \8703 , \7590 , \7165 );
or \U$8451 ( \8704 , \8702 , \8703 );
xor \U$8452 ( \8705 , \7602 , \7609 );
and \U$8453 ( \8706 , \8705 , \7617 );
and \U$8454 ( \8707 , \7602 , \7609 );
or \U$8455 ( \8708 , \8706 , \8707 );
xor \U$8456 ( \8709 , \8704 , \8708 );
xor \U$8457 ( \8710 , \7625 , \7629 );
and \U$8458 ( \8711 , \8710 , \7634 );
and \U$8459 ( \8712 , \7625 , \7629 );
or \U$8460 ( \8713 , \8711 , \8712 );
xor \U$8461 ( \8714 , \8709 , \8713 );
xor \U$8462 ( \8715 , \8535 , \8555 );
and \U$8463 ( \8716 , \8715 , \8581 );
and \U$8464 ( \8717 , \8535 , \8555 );
or \U$8465 ( \8718 , \8716 , \8717 );
xor \U$8466 ( \8719 , \7567 , \7574 );
and \U$8467 ( \8720 , \8719 , \7582 );
and \U$8468 ( \8721 , \7567 , \7574 );
or \U$8469 ( \8722 , \8720 , \8721 );
xor \U$8470 ( \8723 , \8718 , \8722 );
xor \U$8471 ( \8724 , \7669 , \7671 );
and \U$8472 ( \8725 , \8724 , \7681 );
and \U$8473 ( \8726 , \7669 , \7671 );
or \U$8474 ( \8727 , \8725 , \8726 );
xor \U$8475 ( \8728 , \8723 , \8727 );
xor \U$8476 ( \8729 , \8714 , \8728 );
nand \U$8477 ( \8730 , \7562 , \7537 );
and \U$8478 ( \8731 , \8730 , \7549 );
nor \U$8479 ( \8732 , \7537 , \7562 );
nor \U$8480 ( \8733 , \8731 , \8732 );
not \U$8481 ( \8734 , \8733 );
not \U$8482 ( \8735 , \7660 );
not \U$8483 ( \8736 , \7648 );
or \U$8484 ( \8737 , \8735 , \8736 );
nand \U$8485 ( \8738 , \8737 , \7659 );
not \U$8486 ( \8739 , \7648 );
nand \U$8487 ( \8740 , \8739 , \7661 );
nand \U$8488 ( \8741 , \8738 , \8740 );
not \U$8489 ( \8742 , \8741 );
not \U$8490 ( \8743 , \6424 );
and \U$8491 ( \8744 , \6448 , \8743 );
nor \U$8492 ( \8745 , \8744 , \6435 );
nor \U$8493 ( \8746 , \6448 , \8743 );
nor \U$8494 ( \8747 , \8745 , \8746 );
not \U$8495 ( \8748 , \8747 );
or \U$8496 ( \8749 , \8742 , \8748 );
or \U$8497 ( \8750 , \8747 , \8741 );
nand \U$8498 ( \8751 , \8749 , \8750 );
not \U$8499 ( \8752 , \8751 );
or \U$8500 ( \8753 , \8734 , \8752 );
or \U$8501 ( \8754 , \8751 , \8733 );
nand \U$8502 ( \8755 , \8753 , \8754 );
xor \U$8503 ( \8756 , \7596 , \7618 );
and \U$8504 ( \8757 , \8756 , \7635 );
and \U$8505 ( \8758 , \7596 , \7618 );
or \U$8506 ( \8759 , \8757 , \8758 );
xor \U$8507 ( \8760 , \8755 , \8759 );
nand \U$8508 ( \8761 , \6319 , \6331 );
and \U$8509 ( \8762 , \8761 , \6308 );
nor \U$8510 ( \8763 , \6331 , \6319 );
nor \U$8511 ( \8764 , \8762 , \8763 );
and \U$8512 ( \8765 , RIbe29380_53, RIbe2acd0_107);
nor \U$8513 ( \8766 , \8764 , \8765 );
not \U$8514 ( \8767 , \8766 );
nand \U$8515 ( \8768 , \8764 , \8765 );
nand \U$8516 ( \8769 , \8767 , \8768 );
and \U$8517 ( \8770 , \260 , RIbe29e48_76);
and \U$8518 ( \8771 , \264 , RIbe29dd0_75);
nor \U$8519 ( \8772 , \8770 , \8771 );
and \U$8520 ( \8773 , \8772 , \1362 );
not \U$8521 ( \8774 , \8772 );
and \U$8522 ( \8775 , \8774 , \1663 );
nor \U$8523 ( \8776 , \8773 , \8775 );
and \U$8524 ( \8777 , \1528 , RIbe29c68_72);
and \U$8525 ( \8778 , \1256 , RIbe29bf0_71);
nor \U$8526 ( \8779 , \8777 , \8778 );
and \U$8527 ( \8780 , \8779 , \293 );
not \U$8528 ( \8781 , \8779 );
and \U$8529 ( \8782 , \8781 , \300 );
nor \U$8530 ( \8783 , \8780 , \8782 );
buf \U$8531 ( \8784 , \8783 );
xor \U$8532 ( \8785 , \8776 , \8784 );
not \U$8533 ( \8786 , RIbe2a028_80);
not \U$8534 ( \8787 , \324 );
or \U$8535 ( \8788 , \8786 , \8787 );
nand \U$8536 ( \8789 , \329 , RIbe29fb0_79);
nand \U$8537 ( \8790 , \8788 , \8789 );
not \U$8538 ( \8791 , \8790 );
not \U$8539 ( \8792 , \1379 );
and \U$8540 ( \8793 , \8791 , \8792 );
and \U$8541 ( \8794 , \8790 , \1374 );
nor \U$8542 ( \8795 , \8793 , \8794 );
xnor \U$8543 ( \8796 , \8785 , \8795 );
xor \U$8544 ( \8797 , \8769 , \8796 );
not \U$8545 ( \8798 , \6378 );
not \U$8546 ( \8799 , \6403 );
or \U$8547 ( \8800 , \8798 , \8799 );
or \U$8548 ( \8801 , \6403 , \6378 );
nand \U$8549 ( \8802 , \8801 , \6389 );
nand \U$8550 ( \8803 , \8800 , \8802 );
nand \U$8551 ( \8804 , \6460 , \6473 );
and \U$8552 ( \8805 , \8804 , \6482 );
nor \U$8553 ( \8806 , \6460 , \6473 );
nor \U$8554 ( \8807 , \8805 , \8806 );
not \U$8555 ( \8808 , \8807 );
and \U$8556 ( \8809 , \8803 , \8808 );
not \U$8557 ( \8810 , \8803 );
and \U$8558 ( \8811 , \8810 , \8807 );
nor \U$8559 ( \8812 , \8809 , \8811 );
nand \U$8560 ( \8813 , \6344 , \6364 );
and \U$8561 ( \8814 , \8813 , \6356 );
nor \U$8562 ( \8815 , \6344 , \6364 );
nor \U$8563 ( \8816 , \8814 , \8815 );
and \U$8564 ( \8817 , \8812 , \8816 );
not \U$8565 ( \8818 , \8812 );
not \U$8566 ( \8819 , \8816 );
and \U$8567 ( \8820 , \8818 , \8819 );
or \U$8568 ( \8821 , \8817 , \8820 );
xor \U$8569 ( \8822 , \8797 , \8821 );
not \U$8570 ( \8823 , \1284 );
and \U$8571 ( \8824 , \8823 , RIbe28b88_36);
and \U$8572 ( \8825 , \6383 , RIbe29290_51);
nor \U$8573 ( \8826 , \8824 , \8825 );
and \U$8574 ( \8827 , \8826 , \1131 );
not \U$8575 ( \8828 , \8826 );
and \U$8576 ( \8829 , \8828 , \3491 );
nor \U$8577 ( \8830 , \8827 , \8829 );
not \U$8578 ( \8831 , \8830 );
not \U$8579 ( \8832 , RIbe28a20_33);
not \U$8580 ( \8833 , \1271 );
not \U$8581 ( \8834 , \8833 );
or \U$8582 ( \8835 , \8832 , \8834 );
nand \U$8583 ( \8836 , \2384 , RIbe289a8_32);
nand \U$8584 ( \8837 , \8835 , \8836 );
not \U$8585 ( \8838 , \8837 );
not \U$8586 ( \8839 , \1076 );
and \U$8587 ( \8840 , \8838 , \8839 );
and \U$8588 ( \8841 , \8837 , \1076 );
nor \U$8589 ( \8842 , \8840 , \8841 );
not \U$8590 ( \8843 , RIbe28930_31);
not \U$8591 ( \8844 , \4050 );
or \U$8592 ( \8845 , \8843 , \8844 );
nand \U$8593 ( \8846 , \3267 , RIbe29560_57);
nand \U$8594 ( \8847 , \8845 , \8846 );
and \U$8595 ( \8848 , \8847 , \2576 );
not \U$8596 ( \8849 , \8847 );
and \U$8597 ( \8850 , \8849 , \4287 );
nor \U$8598 ( \8851 , \8848 , \8850 );
xor \U$8599 ( \8852 , \8842 , \8851 );
not \U$8600 ( \8853 , \8852 );
or \U$8601 ( \8854 , \8831 , \8853 );
or \U$8602 ( \8855 , \8852 , \8830 );
nand \U$8603 ( \8856 , \8854 , \8855 );
not \U$8604 ( \8857 , RIbe28480_21);
not \U$8605 ( \8858 , \1143 );
or \U$8606 ( \8859 , \8857 , \8858 );
nand \U$8607 ( \8860 , \1147 , RIbe28408_20);
nand \U$8608 ( \8861 , \8859 , \8860 );
not \U$8609 ( \8862 , \8861 );
not \U$8610 ( \8863 , \1153 );
and \U$8611 ( \8864 , \8862 , \8863 );
and \U$8612 ( \8865 , \8861 , \3994 );
nor \U$8613 ( \8866 , \8864 , \8865 );
not \U$8614 ( \8867 , RIbe28390_19);
not \U$8615 ( \8868 , \1093 );
not \U$8616 ( \8869 , \8868 );
or \U$8617 ( \8870 , \8867 , \8869 );
nand \U$8618 ( \8871 , \1455 , RIbe28b10_35);
nand \U$8619 ( \8872 , \8870 , \8871 );
and \U$8620 ( \8873 , \8872 , \1309 );
not \U$8621 ( \8874 , \8872 );
and \U$8622 ( \8875 , \8874 , \4251 );
nor \U$8623 ( \8876 , \8873 , \8875 );
xor \U$8624 ( \8877 , \8866 , \8876 );
and \U$8625 ( \8878 , \1003 , RIbe285e8_24);
and \U$8626 ( \8879 , \1203 , RIbe287c8_28);
nor \U$8627 ( \8880 , \8878 , \8879 );
and \U$8628 ( \8881 , \8880 , \1813 );
not \U$8629 ( \8882 , \8880 );
and \U$8630 ( \8883 , \8882 , \1011 );
nor \U$8631 ( \8884 , \8881 , \8883 );
xor \U$8632 ( \8885 , \8877 , \8884 );
not \U$8633 ( \8886 , \8885 );
not \U$8634 ( \8887 , \8886 );
and \U$8635 ( \8888 , \1756 , RIbe27fd0_11);
and \U$8636 ( \8889 , \1327 , RIbe27f58_10);
nor \U$8637 ( \8890 , \8888 , \8889 );
and \U$8638 ( \8891 , \8890 , \1333 );
not \U$8639 ( \8892 , \8890 );
and \U$8640 ( \8893 , \8892 , \1245 );
nor \U$8641 ( \8894 , \8891 , \8893 );
not \U$8642 ( \8895 , RIbe27e68_8);
not \U$8643 ( \8896 , \6350 );
or \U$8644 ( \8897 , \8895 , \8896 );
nand \U$8645 ( \8898 , \740 , RIbe28660_25);
nand \U$8646 ( \8899 , \8897 , \8898 );
not \U$8647 ( \8900 , \8899 );
not \U$8648 ( \8901 , \564 );
and \U$8649 ( \8902 , \8900 , \8901 );
and \U$8650 ( \8903 , \8899 , \564 );
nor \U$8651 ( \8904 , \8902 , \8903 );
xor \U$8652 ( \8905 , \8894 , \8904 );
not \U$8653 ( \8906 , RIbe28f48_44);
not \U$8654 ( \8907 , \1774 );
or \U$8655 ( \8908 , \8906 , \8907 );
nand \U$8656 ( \8909 , \429 , RIbe28ed0_43);
nand \U$8657 ( \8910 , \8908 , \8909 );
not \U$8658 ( \8911 , \8910 );
not \U$8659 ( \8912 , \313 );
and \U$8660 ( \8913 , \8911 , \8912 );
and \U$8661 ( \8914 , \8910 , \1547 );
nor \U$8662 ( \8915 , \8913 , \8914 );
not \U$8663 ( \8916 , \8915 );
and \U$8664 ( \8917 , \8905 , \8916 );
not \U$8665 ( \8918 , \8905 );
and \U$8666 ( \8919 , \8918 , \8915 );
nor \U$8667 ( \8920 , \8917 , \8919 );
not \U$8668 ( \8921 , \8920 );
or \U$8669 ( \8922 , \8887 , \8921 );
not \U$8670 ( \8923 , \8920 );
nand \U$8671 ( \8924 , \8885 , \8923 );
nand \U$8672 ( \8925 , \8922 , \8924 );
xor \U$8673 ( \8926 , \8856 , \8925 );
xor \U$8674 ( \8927 , \8822 , \8926 );
xor \U$8675 ( \8928 , \8760 , \8927 );
xor \U$8676 ( \8929 , \8729 , \8928 );
xor \U$8677 ( \8930 , \8700 , \8929 );
and \U$8678 ( \8931 , \8666 , \8930 );
and \U$8679 ( \8932 , \7686 , \8665 );
nor \U$8680 ( \8933 , \8931 , \8932 );
not \U$8681 ( \8934 , \8933 );
xor \U$8682 ( \8935 , \8755 , \8759 );
and \U$8683 ( \8936 , \8935 , \8927 );
and \U$8684 ( \8937 , \8755 , \8759 );
or \U$8685 ( \8938 , \8936 , \8937 );
xor \U$8686 ( \8939 , \8718 , \8722 );
and \U$8687 ( \8940 , \8939 , \8727 );
and \U$8688 ( \8941 , \8718 , \8722 );
or \U$8689 ( \8942 , \8940 , \8941 );
xor \U$8690 ( \8943 , \8938 , \8942 );
not \U$8691 ( \8944 , RIbe28e58_42);
not \U$8692 ( \8945 , \6537 );
or \U$8693 ( \8946 , \8944 , \8945 );
nand \U$8694 ( \8947 , \7076 , RIbe28de0_41);
nand \U$8695 ( \8948 , \8946 , \8947 );
and \U$8696 ( \8949 , \8948 , \7546 );
not \U$8697 ( \8950 , \8948 );
and \U$8698 ( \8951 , \8950 , \6546 );
or \U$8699 ( \8952 , \8949 , \8951 );
xor \U$8700 ( \8953 , \6572 , \8952 );
and \U$8701 ( \8954 , \6592 , RIbe29920_65);
and \U$8702 ( \8955 , \6596 , RIbe27b98_2);
nor \U$8703 ( \8956 , \8954 , \8955 );
not \U$8704 ( \8957 , \6601 );
and \U$8705 ( \8958 , \8956 , \8957 );
not \U$8706 ( \8959 , \8956 );
and \U$8707 ( \8960 , \8959 , \6601 );
nor \U$8708 ( \8961 , \8958 , \8960 );
xor \U$8709 ( \8962 , \8953 , \8961 );
not \U$8710 ( \8963 , \8886 );
not \U$8711 ( \8964 , \8923 );
or \U$8712 ( \8965 , \8963 , \8964 );
not \U$8713 ( \8966 , \8920 );
not \U$8714 ( \8967 , \8885 );
or \U$8715 ( \8968 , \8966 , \8967 );
nand \U$8716 ( \8969 , \8968 , \8856 );
nand \U$8717 ( \8970 , \8965 , \8969 );
xor \U$8718 ( \8971 , \8962 , \8970 );
not \U$8719 ( \8972 , \6528 );
not \U$8720 ( \8973 , \6659 );
or \U$8721 ( \8974 , \8972 , \8973 );
nand \U$8722 ( \8975 , \8974 , \6606 );
or \U$8723 ( \8976 , \6528 , \6659 );
nand \U$8724 ( \8977 , \8975 , \8976 );
xor \U$8725 ( \8978 , \8971 , \8977 );
xor \U$8726 ( \8979 , \8943 , \8978 );
xor \U$8727 ( \8980 , \8691 , \8699 );
and \U$8728 ( \8981 , \8980 , \8929 );
and \U$8729 ( \8982 , \8691 , \8699 );
or \U$8730 ( \8983 , \8981 , \8982 );
xor \U$8731 ( \8984 , \8979 , \8983 );
not \U$8732 ( \8985 , \8796 );
and \U$8733 ( \8986 , \8985 , \8768 );
nor \U$8734 ( \8987 , \8986 , \8766 );
buf \U$8735 ( \8988 , \8987 );
not \U$8736 ( \8989 , \8988 );
not \U$8737 ( \8990 , \8819 );
not \U$8738 ( \8991 , \8808 );
or \U$8739 ( \8992 , \8990 , \8991 );
not \U$8740 ( \8993 , \8816 );
not \U$8741 ( \8994 , \8807 );
or \U$8742 ( \8995 , \8993 , \8994 );
nand \U$8743 ( \8996 , \8995 , \8803 );
nand \U$8744 ( \8997 , \8992 , \8996 );
not \U$8745 ( \8998 , \8997 );
nand \U$8746 ( \8999 , \8733 , \8747 );
and \U$8747 ( \9000 , \8999 , \8741 );
nor \U$8748 ( \9001 , \8747 , \8733 );
nor \U$8749 ( \9002 , \9000 , \9001 );
not \U$8750 ( \9003 , \9002 );
or \U$8751 ( \9004 , \8998 , \9003 );
or \U$8752 ( \9005 , \9002 , \8997 );
nand \U$8753 ( \9006 , \9004 , \9005 );
not \U$8754 ( \9007 , \9006 );
or \U$8755 ( \9008 , \8989 , \9007 );
or \U$8756 ( \9009 , \8988 , \9006 );
nand \U$8757 ( \9010 , \9008 , \9009 );
not \U$8758 ( \9011 , \8866 );
not \U$8759 ( \9012 , \9011 );
not \U$8760 ( \9013 , \8884 );
or \U$8761 ( \9014 , \9012 , \9013 );
or \U$8762 ( \9015 , \9011 , \8884 );
nand \U$8763 ( \9016 , \9015 , \8876 );
nand \U$8764 ( \9017 , \9014 , \9016 );
not \U$8765 ( \9018 , \9017 );
not \U$8766 ( \9019 , \9018 );
and \U$8767 ( \9020 , \8830 , \8851 );
nor \U$8768 ( \9021 , \9020 , \8842 );
nor \U$8769 ( \9022 , \8851 , \8830 );
nor \U$8770 ( \9023 , \9021 , \9022 );
not \U$8771 ( \9024 , \9023 );
not \U$8772 ( \9025 , \8916 );
not \U$8773 ( \9026 , \8894 );
or \U$8774 ( \9027 , \9025 , \9026 );
not \U$8775 ( \9028 , \8904 );
not \U$8776 ( \9029 , \8894 );
nand \U$8777 ( \9030 , \9029 , \8915 );
nand \U$8778 ( \9031 , \9028 , \9030 );
nand \U$8779 ( \9032 , \9027 , \9031 );
not \U$8780 ( \9033 , \9032 );
and \U$8781 ( \9034 , \9024 , \9033 );
and \U$8782 ( \9035 , \9023 , \9032 );
nor \U$8783 ( \9036 , \9034 , \9035 );
not \U$8784 ( \9037 , \9036 );
not \U$8785 ( \9038 , \9037 );
or \U$8786 ( \9039 , \9019 , \9038 );
not \U$8787 ( \9040 , \9018 );
nand \U$8788 ( \9041 , \9040 , \9036 );
nand \U$8789 ( \9042 , \9039 , \9041 );
not \U$8790 ( \9043 , \6499 );
not \U$8791 ( \9044 , \6524 );
or \U$8792 ( \9045 , \9043 , \9044 );
nand \U$8793 ( \9046 , \9045 , \6510 );
nand \U$8794 ( \9047 , \6523 , \6498 );
nand \U$8795 ( \9048 , \9046 , \9047 );
not \U$8796 ( \9049 , \6577 );
not \U$8797 ( \9050 , \6604 );
or \U$8798 ( \9051 , \9049 , \9050 );
or \U$8799 ( \9052 , \6604 , \6577 );
nand \U$8800 ( \9053 , \9052 , \6554 );
nand \U$8801 ( \9054 , \9051 , \9053 );
xor \U$8802 ( \9055 , \9048 , \9054 );
not \U$8803 ( \9056 , \6654 );
not \U$8804 ( \9057 , \6647 );
or \U$8805 ( \9058 , \9056 , \9057 );
or \U$8806 ( \9059 , \6654 , \6647 );
nand \U$8807 ( \9060 , \9059 , \6626 );
nand \U$8808 ( \9061 , \9058 , \9060 );
xor \U$8809 ( \9062 , \9055 , \9061 );
xnor \U$8810 ( \9063 , \9042 , \9062 );
not \U$8811 ( \9064 , \9063 );
not \U$8812 ( \9065 , \9064 );
not \U$8813 ( \9066 , RIbe29560_57);
not \U$8814 ( \9067 , \4050 );
or \U$8815 ( \9068 , \9066 , \9067 );
nand \U$8816 ( \9069 , \3267 , RIbe28228_16);
nand \U$8817 ( \9070 , \9068 , \9069 );
and \U$8818 ( \9071 , \9070 , \4287 );
not \U$8819 ( \9072 , \9070 );
and \U$8820 ( \9073 , \9072 , \4059 );
nor \U$8821 ( \9074 , \9071 , \9073 );
not \U$8822 ( \9075 , \9074 );
not \U$8823 ( \9076 , \9075 );
not \U$8824 ( \9077 , \4065 );
not \U$8825 ( \9078 , RIbe28930_31);
not \U$8826 ( \9079 , \9078 );
and \U$8827 ( \9080 , \9077 , \9079 );
and \U$8828 ( \9081 , \3303 , RIbe289a8_32);
nor \U$8829 ( \9082 , \9080 , \9081 );
not \U$8830 ( \9083 , \1275 );
and \U$8831 ( \9084 , \9082 , \9083 );
not \U$8832 ( \9085 , \9082 );
and \U$8833 ( \9086 , \9085 , \1076 );
nor \U$8834 ( \9087 , \9084 , \9086 );
not \U$8835 ( \9088 , \9087 );
not \U$8836 ( \9089 , \9088 );
or \U$8837 ( \9090 , \9076 , \9089 );
nand \U$8838 ( \9091 , \9074 , \9087 );
nand \U$8839 ( \9092 , \9090 , \9091 );
and \U$8840 ( \9093 , \8823 , RIbe29290_51);
and \U$8841 ( \9094 , \6383 , RIbe28a20_33);
nor \U$8842 ( \9095 , \9093 , \9094 );
and \U$8843 ( \9096 , \9095 , \1131 );
not \U$8844 ( \9097 , \9095 );
and \U$8845 ( \9098 , \9097 , \3491 );
nor \U$8846 ( \9099 , \9096 , \9098 );
buf \U$8847 ( \9100 , \9099 );
xor \U$8848 ( \9101 , \9092 , \9100 );
not \U$8849 ( \9102 , RIbe29830_63);
not \U$8850 ( \9103 , \4021 );
or \U$8851 ( \9104 , \9102 , \9103 );
nand \U$8852 ( \9105 , \7438 , RIbe296c8_60);
nand \U$8853 ( \9106 , \9104 , \9105 );
and \U$8854 ( \9107 , \9106 , \3471 );
not \U$8855 ( \9108 , \9106 );
and \U$8856 ( \9109 , \9108 , \4821 );
nor \U$8857 ( \9110 , \9107 , \9109 );
not \U$8858 ( \9111 , RIbe29650_59);
not \U$8859 ( \9112 , \5058 );
or \U$8860 ( \9113 , \9111 , \9112 );
nand \U$8861 ( \9114 , \4600 , RIbe29038_46);
nand \U$8862 ( \9115 , \9113 , \9114 );
and \U$8863 ( \9116 , \9115 , \4326 );
not \U$8864 ( \9117 , \9115 );
and \U$8865 ( \9118 , \9117 , \4323 );
nor \U$8866 ( \9119 , \9116 , \9118 );
xor \U$8867 ( \9120 , \9110 , \9119 );
not \U$8868 ( \9121 , RIbe281b0_15);
not \U$8869 ( \9122 , \4764 );
or \U$8870 ( \9123 , \9121 , \9122 );
nand \U$8871 ( \9124 , \3689 , RIbe280c0_13);
nand \U$8872 ( \9125 , \9123 , \9124 );
and \U$8873 ( \9126 , \9125 , \3290 );
not \U$8874 ( \9127 , \9125 );
and \U$8875 ( \9128 , \9127 , \2887 );
nor \U$8876 ( \9129 , \9126 , \9128 );
xor \U$8877 ( \9130 , \9120 , \9129 );
xor \U$8878 ( \9131 , \9101 , \9130 );
not \U$8879 ( \9132 , RIbe27d00_5);
not \U$8880 ( \9133 , \6856 );
or \U$8881 ( \9134 , \9132 , \9133 );
nand \U$8882 ( \9135 , \6617 , RIbe27c10_3);
nand \U$8883 ( \9136 , \9134 , \9135 );
and \U$8884 ( \9137 , \9136 , \6624 );
not \U$8885 ( \9138 , \9136 );
and \U$8886 ( \9139 , \9138 , \6620 );
nor \U$8887 ( \9140 , \9137 , \9139 );
not \U$8888 ( \9141 , \9140 );
not \U$8889 ( \9142 , \9141 );
not \U$8890 ( \9143 , RIbe29a88_68);
not \U$8891 ( \9144 , \5455 );
or \U$8892 ( \9145 , \9143 , \9144 );
nand \U$8893 ( \9146 , \8247 , RIbe27d78_6);
nand \U$8894 ( \9147 , \9145 , \9146 );
and \U$8895 ( \9148 , \9147 , \6117 );
not \U$8896 ( \9149 , \9147 );
and \U$8897 ( \9150 , \9149 , \5754 );
nor \U$8898 ( \9151 , \9148 , \9150 );
not \U$8899 ( \9152 , \9151 );
not \U$8900 ( \9153 , \9152 );
or \U$8901 ( \9154 , \9142 , \9153 );
nand \U$8902 ( \9155 , \9151 , \9140 );
nand \U$8903 ( \9156 , \9154 , \9155 );
not \U$8904 ( \9157 , RIbe28fc0_45);
not \U$8905 ( \9158 , \4830 );
or \U$8906 ( \9159 , \9157 , \9158 );
nand \U$8907 ( \9160 , \5731 , RIbe290b0_47);
nand \U$8908 ( \9161 , \9159 , \9160 );
and \U$8909 ( \9162 , \9161 , \4946 );
not \U$8910 ( \9163 , \9161 );
and \U$8911 ( \9164 , \9163 , \4586 );
nor \U$8912 ( \9165 , \9162 , \9164 );
xor \U$8913 ( \9166 , \9156 , \9165 );
not \U$8914 ( \9167 , \9166 );
and \U$8915 ( \9168 , \9131 , \9167 );
not \U$8916 ( \9169 , \9131 );
and \U$8917 ( \9170 , \9169 , \9166 );
nor \U$8918 ( \9171 , \9168 , \9170 );
not \U$8919 ( \9172 , \9171 );
not \U$8920 ( \9173 , \9172 );
and \U$8921 ( \9174 , \1659 , RIbe29dd0_75);
and \U$8922 ( \9175 , \6325 , RIbe29c68_72);
nor \U$8923 ( \9176 , \9174 , \9175 );
and \U$8924 ( \9177 , \9176 , \1363 );
not \U$8925 ( \9178 , \9176 );
and \U$8926 ( \9179 , \9178 , \270 );
nor \U$8927 ( \9180 , \9177 , \9179 );
not \U$8928 ( \9181 , RIbe29fb0_79);
not \U$8929 ( \9182 , \325 );
or \U$8930 ( \9183 , \9181 , \9182 );
nand \U$8931 ( \9184 , \330 , RIbe29e48_76);
nand \U$8932 ( \9185 , \9183 , \9184 );
not \U$8933 ( \9186 , \9185 );
not \U$8934 ( \9187 , \1379 );
and \U$8935 ( \9188 , \9186 , \9187 );
and \U$8936 ( \9189 , \9185 , \1379 );
nor \U$8937 ( \9190 , \9188 , \9189 );
xor \U$8938 ( \9191 , \9180 , \9190 );
and \U$8939 ( \9192 , \3895 , RIbe29bf0_71);
and \U$8940 ( \9193 , \1256 , RIbe28f48_44);
nor \U$8941 ( \9194 , \9192 , \9193 );
and \U$8942 ( \9195 , \9194 , \293 );
not \U$8943 ( \9196 , \9194 );
and \U$8944 ( \9197 , \9196 , \300 );
nor \U$8945 ( \9198 , \9195 , \9197 );
xor \U$8946 ( \9199 , \9191 , \9198 );
not \U$8947 ( \9200 , \9199 );
not \U$8948 ( \9201 , RIbe287c8_28);
not \U$8949 ( \9202 , \1003 );
or \U$8950 ( \9203 , \9201 , \9202 );
nand \U$8951 ( \9204 , \1203 , RIbe28480_21);
nand \U$8952 ( \9205 , \9203 , \9204 );
not \U$8953 ( \9206 , \9205 );
not \U$8954 ( \9207 , \1813 );
and \U$8955 ( \9208 , \9206 , \9207 );
and \U$8956 ( \9209 , \9205 , \1608 );
nor \U$8957 ( \9210 , \9208 , \9209 );
not \U$8958 ( \9211 , \9210 );
not \U$8959 ( \9212 , RIbe28408_20);
not \U$8960 ( \9213 , \4257 );
or \U$8961 ( \9214 , \9212 , \9213 );
nand \U$8962 ( \9215 , \1147 , RIbe28390_19);
nand \U$8963 ( \9216 , \9214 , \9215 );
xor \U$8964 ( \9217 , \9216 , \4742 );
not \U$8965 ( \9218 , \9217 );
not \U$8966 ( \9219 , \1080 );
not \U$8967 ( \9220 , RIbe28b10_35);
not \U$8968 ( \9221 , \8868 );
or \U$8969 ( \9222 , \9220 , \9221 );
nand \U$8970 ( \9223 , \4730 , RIbe28b88_36);
nand \U$8971 ( \9224 , \9222 , \9223 );
not \U$8972 ( \9225 , \9224 );
or \U$8973 ( \9226 , \9219 , \9225 );
or \U$8974 ( \9227 , \9224 , \2418 );
nand \U$8975 ( \9228 , \9226 , \9227 );
not \U$8976 ( \9229 , \9228 );
or \U$8977 ( \9230 , \9218 , \9229 );
or \U$8978 ( \9231 , \9228 , \9217 );
nand \U$8979 ( \9232 , \9230 , \9231 );
not \U$8980 ( \9233 , \9232 );
or \U$8981 ( \9234 , \9211 , \9233 );
or \U$8982 ( \9235 , \9232 , \9210 );
nand \U$8983 ( \9236 , \9234 , \9235 );
not \U$8984 ( \9237 , \9236 );
not \U$8985 ( \9238 , RIbe28ed0_43);
and \U$8986 ( \9239 , \375 , \380 );
not \U$8987 ( \9240 , \9239 );
or \U$8988 ( \9241 , \9238 , \9240 );
nand \U$8989 ( \9242 , \428 , RIbe27fd0_11);
nand \U$8990 ( \9243 , \9241 , \9242 );
not \U$8991 ( \9244 , \9243 );
not \U$8992 ( \9245 , \312 );
and \U$8993 ( \9246 , \9244 , \9245 );
and \U$8994 ( \9247 , \9243 , \313 );
nor \U$8995 ( \9248 , \9246 , \9247 );
and \U$8996 ( \9249 , \2531 , RIbe28660_25);
and \U$8997 ( \9250 , \1179 , RIbe285e8_24);
nor \U$8998 ( \9251 , \9249 , \9250 );
not \U$8999 ( \9252 , \9251 );
not \U$9000 ( \9253 , \3959 );
and \U$9001 ( \9254 , \9252 , \9253 );
and \U$9002 ( \9255 , \672 , \9251 );
nor \U$9003 ( \9256 , \9254 , \9255 );
xor \U$9004 ( \9257 , \9248 , \9256 );
not \U$9005 ( \9258 , RIbe27f58_10);
not \U$9006 ( \9259 , \3244 );
or \U$9007 ( \9260 , \9258 , \9259 );
nand \U$9008 ( \9261 , \1327 , RIbe27e68_8);
nand \U$9009 ( \9262 , \9260 , \9261 );
not \U$9010 ( \9263 , \9262 );
not \U$9011 ( \9264 , \424 );
and \U$9012 ( \9265 , \9263 , \9264 );
and \U$9013 ( \9266 , \9262 , \1333 );
nor \U$9014 ( \9267 , \9265 , \9266 );
xor \U$9015 ( \9268 , \9257 , \9267 );
not \U$9016 ( \9269 , \9268 );
or \U$9017 ( \9270 , \9237 , \9269 );
or \U$9018 ( \9271 , \9236 , \9268 );
nand \U$9019 ( \9272 , \9270 , \9271 );
not \U$9020 ( \9273 , \9272 );
or \U$9021 ( \9274 , \9200 , \9273 );
or \U$9022 ( \9275 , \9272 , \9199 );
nand \U$9023 ( \9276 , \9274 , \9275 );
not \U$9024 ( \9277 , \9276 );
nand \U$9025 ( \9278 , \8783 , \8795 );
and \U$9026 ( \9279 , \9278 , \8776 );
nor \U$9027 ( \9280 , \8783 , \8795 );
nor \U$9028 ( \9281 , \9279 , \9280 );
and \U$9029 ( \9282 , RIbe29380_53, RIbe2a028_80);
xnor \U$9030 ( \9283 , \9282 , \8765 );
xnor \U$9031 ( \9284 , \9281 , \9283 );
not \U$9032 ( \9285 , \9284 );
and \U$9033 ( \9286 , \9277 , \9285 );
and \U$9034 ( \9287 , \9276 , \9284 );
nor \U$9035 ( \9288 , \9286 , \9287 );
not \U$9036 ( \9289 , \9288 );
or \U$9037 ( \9290 , \9173 , \9289 );
or \U$9038 ( \9291 , \9288 , \9172 );
nand \U$9039 ( \9292 , \9290 , \9291 );
not \U$9040 ( \9293 , \9292 );
not \U$9041 ( \9294 , \9293 );
or \U$9042 ( \9295 , \9065 , \9294 );
nand \U$9043 ( \9296 , \9292 , \9063 );
nand \U$9044 ( \9297 , \9295 , \9296 );
xor \U$9045 ( \9298 , \9010 , \9297 );
xor \U$9046 ( \9299 , \8704 , \8708 );
and \U$9047 ( \9300 , \9299 , \8713 );
and \U$9048 ( \9301 , \8704 , \8708 );
or \U$9049 ( \9302 , \9300 , \9301 );
xor \U$9050 ( \9303 , \6368 , \6488 );
and \U$9051 ( \9304 , \9303 , \6660 );
and \U$9052 ( \9305 , \6368 , \6488 );
or \U$9053 ( \9306 , \9304 , \9305 );
xor \U$9054 ( \9307 , \9302 , \9306 );
xor \U$9055 ( \9308 , \8797 , \8821 );
and \U$9056 ( \9309 , \9308 , \8926 );
and \U$9057 ( \9310 , \8797 , \8821 );
or \U$9058 ( \9311 , \9309 , \9310 );
xor \U$9059 ( \9312 , \9307 , \9311 );
xnor \U$9060 ( \9313 , \9298 , \9312 );
not \U$9061 ( \9314 , \9313 );
xor \U$9062 ( \9315 , \8714 , \8728 );
and \U$9063 ( \9316 , \9315 , \8928 );
and \U$9064 ( \9317 , \8714 , \8728 );
or \U$9065 ( \9318 , \9316 , \9317 );
xor \U$9066 ( \9319 , \6661 , \7523 );
and \U$9067 ( \9320 , \9319 , \7685 );
and \U$9068 ( \9321 , \6661 , \7523 );
or \U$9069 ( \9322 , \9320 , \9321 );
and \U$9070 ( \9323 , \9318 , \9322 );
not \U$9071 ( \9324 , \9318 );
not \U$9072 ( \9325 , \9322 );
and \U$9073 ( \9326 , \9324 , \9325 );
nor \U$9074 ( \9327 , \9323 , \9326 );
not \U$9075 ( \9328 , \9327 );
or \U$9076 ( \9329 , \9314 , \9328 );
or \U$9077 ( \9330 , \9313 , \9327 );
nand \U$9078 ( \9331 , \9329 , \9330 );
xor \U$9079 ( \9332 , \8984 , \9331 );
nand \U$9080 ( \9333 , \8934 , \9332 );
not \U$9081 ( \9334 , \9333 );
not \U$9082 ( \9335 , \9334 );
xor \U$9083 ( \9336 , \8979 , \8983 );
and \U$9084 ( \9337 , \9336 , \9331 );
and \U$9085 ( \9338 , \8979 , \8983 );
or \U$9086 ( \9339 , \9337 , \9338 );
not \U$9087 ( \9340 , \9339 );
xor \U$9088 ( \9341 , \8962 , \8970 );
and \U$9089 ( \9342 , \9341 , \8977 );
and \U$9090 ( \9343 , \8962 , \8970 );
or \U$9091 ( \9344 , \9342 , \9343 );
not \U$9092 ( \9345 , \8997 );
not \U$9093 ( \9346 , \9002 );
not \U$9094 ( \9347 , \9346 );
or \U$9095 ( \9348 , \9345 , \9347 );
not \U$9096 ( \9349 , \8987 );
not \U$9097 ( \9350 , \8997 );
nand \U$9098 ( \9351 , \9350 , \9002 );
nand \U$9099 ( \9352 , \9349 , \9351 );
nand \U$9100 ( \9353 , \9348 , \9352 );
xor \U$9101 ( \9354 , \9344 , \9353 );
nand \U$9102 ( \9355 , \9171 , \9284 );
and \U$9103 ( \9356 , \9355 , \9276 );
nor \U$9104 ( \9357 , \9171 , \9284 );
nor \U$9105 ( \9358 , \9356 , \9357 );
xnor \U$9106 ( \9359 , \9354 , \9358 );
not \U$9107 ( \9360 , \9042 );
not \U$9108 ( \9361 , \9062 );
or \U$9109 ( \9362 , \9360 , \9361 );
or \U$9110 ( \9363 , \9062 , \9042 );
nand \U$9111 ( \9364 , \9363 , \9292 );
nand \U$9112 ( \9365 , \9362 , \9364 );
not \U$9113 ( \9366 , \9365 );
xor \U$9114 ( \9367 , \9359 , \9366 );
xor \U$9115 ( \9368 , \9302 , \9306 );
and \U$9116 ( \9369 , \9368 , \9311 );
and \U$9117 ( \9370 , \9302 , \9306 );
or \U$9118 ( \9371 , \9369 , \9370 );
not \U$9119 ( \9372 , \9282 );
not \U$9120 ( \9373 , \8765 );
or \U$9121 ( \9374 , \9372 , \9373 );
not \U$9122 ( \9375 , \9281 );
or \U$9123 ( \9376 , \8765 , \9282 );
nand \U$9124 ( \9377 , \9375 , \9376 );
nand \U$9125 ( \9378 , \9374 , \9377 );
not \U$9126 ( \9379 , \9032 );
not \U$9127 ( \9380 , \9023 );
not \U$9128 ( \9381 , \9380 );
or \U$9129 ( \9382 , \9379 , \9381 );
or \U$9130 ( \9383 , \9380 , \9032 );
nand \U$9131 ( \9384 , \9383 , \9017 );
nand \U$9132 ( \9385 , \9382 , \9384 );
xor \U$9133 ( \9386 , \9378 , \9385 );
xor \U$9134 ( \9387 , \9048 , \9054 );
and \U$9135 ( \9388 , \9387 , \9061 );
and \U$9136 ( \9389 , \9048 , \9054 );
or \U$9137 ( \9390 , \9388 , \9389 );
xor \U$9138 ( \9391 , \9386 , \9390 );
not \U$9139 ( \9392 , \9391 );
and \U$9140 ( \9393 , \9371 , \9392 );
not \U$9141 ( \9394 , \9371 );
and \U$9142 ( \9395 , \9394 , \9391 );
nor \U$9143 ( \9396 , \9393 , \9395 );
xnor \U$9144 ( \9397 , \9367 , \9396 );
not \U$9145 ( \9398 , \9397 );
not \U$9146 ( \9399 , \9398 );
xor \U$9147 ( \9400 , \9110 , \9119 );
and \U$9148 ( \9401 , \9400 , \9129 );
and \U$9149 ( \9402 , \9110 , \9119 );
or \U$9150 ( \9403 , \9401 , \9402 );
xor \U$9151 ( \9404 , \6572 , \8952 );
and \U$9152 ( \9405 , \9404 , \8961 );
and \U$9153 ( \9406 , \6572 , \8952 );
or \U$9154 ( \9407 , \9405 , \9406 );
xor \U$9155 ( \9408 , \9403 , \9407 );
or \U$9156 ( \9409 , \9165 , \9152 );
not \U$9157 ( \9410 , \9152 );
not \U$9158 ( \9411 , \9165 );
or \U$9159 ( \9412 , \9410 , \9411 );
nand \U$9160 ( \9413 , \9412 , \9141 );
nand \U$9161 ( \9414 , \9409 , \9413 );
xor \U$9162 ( \9415 , \9408 , \9414 );
nand \U$9163 ( \9416 , RIbe29380_53, RIbe29fb0_79);
and \U$9164 ( \9417 , \325 , RIbe29e48_76);
and \U$9165 ( \9418 , \329 , RIbe29dd0_75);
nor \U$9166 ( \9419 , \9417 , \9418 );
and \U$9167 ( \9420 , \9419 , \1375 );
not \U$9168 ( \9421 , \9419 );
and \U$9169 ( \9422 , \9421 , \1374 );
nor \U$9170 ( \9423 , \9420 , \9422 );
xor \U$9171 ( \9424 , \9416 , \9423 );
not \U$9172 ( \9425 , \269 );
and \U$9173 ( \9426 , \261 , RIbe29c68_72);
and \U$9174 ( \9427 , \1831 , RIbe29bf0_71);
nor \U$9175 ( \9428 , \9426 , \9427 );
not \U$9176 ( \9429 , \9428 );
or \U$9177 ( \9430 , \9425 , \9429 );
or \U$9178 ( \9431 , \9428 , \269 );
nand \U$9179 ( \9432 , \9430 , \9431 );
xnor \U$9180 ( \9433 , \9424 , \9432 );
xor \U$9181 ( \9434 , \9180 , \9190 );
and \U$9182 ( \9435 , \9434 , \9198 );
and \U$9183 ( \9436 , \9180 , \9190 );
or \U$9184 ( \9437 , \9435 , \9436 );
nor \U$9185 ( \9438 , \9433 , \9437 );
not \U$9186 ( \9439 , \9438 );
nand \U$9187 ( \9440 , \9433 , \9437 );
nand \U$9188 ( \9441 , \9439 , \9440 );
not \U$9189 ( \9442 , \9441 );
not \U$9190 ( \9443 , \9442 );
and \U$9191 ( \9444 , \9099 , \9075 );
nor \U$9192 ( \9445 , \9444 , \9087 );
nor \U$9193 ( \9446 , \9075 , \9099 );
nor \U$9194 ( \9447 , \9445 , \9446 );
xor \U$9195 ( \9448 , \9248 , \9256 );
and \U$9196 ( \9449 , \9448 , \9267 );
and \U$9197 ( \9450 , \9248 , \9256 );
or \U$9198 ( \9451 , \9449 , \9450 );
xor \U$9199 ( \9452 , \9447 , \9451 );
not \U$9200 ( \9453 , \9210 );
not \U$9201 ( \9454 , \9217 );
and \U$9202 ( \9455 , \9453 , \9454 );
and \U$9203 ( \9456 , \9210 , \9217 );
not \U$9204 ( \9457 , \9228 );
nor \U$9205 ( \9458 , \9456 , \9457 );
nor \U$9206 ( \9459 , \9455 , \9458 );
xor \U$9207 ( \9460 , \9452 , \9459 );
not \U$9208 ( \9461 , \9460 );
not \U$9209 ( \9462 , \9461 );
or \U$9210 ( \9463 , \9443 , \9462 );
nand \U$9211 ( \9464 , \9460 , \9441 );
nand \U$9212 ( \9465 , \9463 , \9464 );
not \U$9213 ( \9466 , RIbe27fd0_11);
not \U$9214 ( \9467 , \1223 );
or \U$9215 ( \9468 , \9466 , \9467 );
nand \U$9216 ( \9469 , \429 , RIbe27f58_10);
nand \U$9217 ( \9470 , \9468 , \9469 );
and \U$9218 ( \9471 , \9470 , \306 );
not \U$9219 ( \9472 , \9470 );
and \U$9220 ( \9473 , \9472 , \313 );
nor \U$9221 ( \9474 , \9471 , \9473 );
not \U$9222 ( \9475 , RIbe27e68_8);
not \U$9223 ( \9476 , \1756 );
or \U$9224 ( \9477 , \9475 , \9476 );
nand \U$9225 ( \9478 , \1327 , RIbe28660_25);
nand \U$9226 ( \9479 , \9477 , \9478 );
not \U$9227 ( \9480 , \9479 );
not \U$9228 ( \9481 , \424 );
and \U$9229 ( \9482 , \9480 , \9481 );
and \U$9230 ( \9483 , \9479 , \6340 );
nor \U$9231 ( \9484 , \9482 , \9483 );
and \U$9232 ( \9485 , \9474 , \9484 );
not \U$9233 ( \9486 , \9474 );
not \U$9234 ( \9487 , \9484 );
and \U$9235 ( \9488 , \9486 , \9487 );
or \U$9236 ( \9489 , \9485 , \9488 );
and \U$9237 ( \9490 , \283 , RIbe28f48_44);
and \U$9238 ( \9491 , \1531 , RIbe28ed0_43);
nor \U$9239 ( \9492 , \9490 , \9491 );
and \U$9240 ( \9493 , \9492 , \293 );
not \U$9241 ( \9494 , \9492 );
and \U$9242 ( \9495 , \9494 , \300 );
nor \U$9243 ( \9496 , \9493 , \9495 );
not \U$9244 ( \9497 , \9496 );
and \U$9245 ( \9498 , \9489 , \9497 );
not \U$9246 ( \9499 , \9489 );
and \U$9247 ( \9500 , \9499 , \9496 );
nor \U$9248 ( \9501 , \9498 , \9500 );
and \U$9249 ( \9502 , \5973 , RIbe28480_21);
and \U$9250 ( \9503 , \1203 , RIbe28408_20);
nor \U$9251 ( \9504 , \9502 , \9503 );
and \U$9252 ( \9505 , \9504 , \1011 );
not \U$9253 ( \9506 , \9504 );
and \U$9254 ( \9507 , \9506 , \1813 );
nor \U$9255 ( \9508 , \9505 , \9507 );
not \U$9256 ( \9509 , RIbe285e8_24);
not \U$9257 ( \9510 , \664 );
or \U$9258 ( \9511 , \9509 , \9510 );
nand \U$9259 ( \9512 , \1179 , RIbe287c8_28);
nand \U$9260 ( \9513 , \9511 , \9512 );
not \U$9261 ( \9514 , \9513 );
not \U$9262 ( \9515 , \4217 );
and \U$9263 ( \9516 , \9514 , \9515 );
and \U$9264 ( \9517 , \9513 , \4217 );
nor \U$9265 ( \9518 , \9516 , \9517 );
not \U$9266 ( \9519 , \9518 );
not \U$9267 ( \9520 , \9519 );
not \U$9268 ( \9521 , RIbe28390_19);
not \U$9269 ( \9522 , \2597 );
or \U$9270 ( \9523 , \9521 , \9522 );
nand \U$9271 ( \9524 , \1147 , RIbe28b10_35);
nand \U$9272 ( \9525 , \9523 , \9524 );
and \U$9273 ( \9526 , \9525 , \1652 );
not \U$9274 ( \9527 , \9525 );
and \U$9275 ( \9528 , \9527 , \1157 );
nor \U$9276 ( \9529 , \9526 , \9528 );
not \U$9277 ( \9530 , \9529 );
not \U$9278 ( \9531 , \9530 );
or \U$9279 ( \9532 , \9520 , \9531 );
nand \U$9280 ( \9533 , \9529 , \9518 );
nand \U$9281 ( \9534 , \9532 , \9533 );
xnor \U$9282 ( \9535 , \9508 , \9534 );
xor \U$9283 ( \9536 , \9501 , \9535 );
not \U$9284 ( \9537 , RIbe28b88_36);
not \U$9285 ( \9538 , \1633 );
or \U$9286 ( \9539 , \9537 , \9538 );
nand \U$9287 ( \9540 , \1455 , RIbe29290_51);
nand \U$9288 ( \9541 , \9539 , \9540 );
not \U$9289 ( \9542 , \9541 );
not \U$9290 ( \9543 , \5125 );
and \U$9291 ( \9544 , \9542 , \9543 );
and \U$9292 ( \9545 , \9541 , \5125 );
nor \U$9293 ( \9546 , \9544 , \9545 );
not \U$9294 ( \9547 , RIbe28930_31);
not \U$9295 ( \9548 , \1272 );
or \U$9296 ( \9549 , \9547 , \9548 );
nand \U$9297 ( \9550 , \2384 , RIbe29560_57);
nand \U$9298 ( \9551 , \9549 , \9550 );
not \U$9299 ( \9552 , \9551 );
not \U$9300 ( \9553 , \3516 );
and \U$9301 ( \9554 , \9552 , \9553 );
and \U$9302 ( \9555 , \9551 , \1076 );
nor \U$9303 ( \9556 , \9554 , \9555 );
not \U$9304 ( \9557 , \9556 );
not \U$9305 ( \9558 , \9557 );
and \U$9306 ( \9559 , \1113 , RIbe28a20_33);
and \U$9307 ( \9560 , \1117 , RIbe289a8_32);
nor \U$9308 ( \9561 , \9559 , \9560 );
and \U$9309 ( \9562 , \9561 , \1448 );
not \U$9310 ( \9563 , \9561 );
and \U$9311 ( \9564 , \9563 , \1131 );
nor \U$9312 ( \9565 , \9562 , \9564 );
not \U$9313 ( \9566 , \9565 );
not \U$9314 ( \9567 , \9566 );
or \U$9315 ( \9568 , \9558 , \9567 );
nand \U$9316 ( \9569 , \9565 , \9556 );
nand \U$9317 ( \9570 , \9568 , \9569 );
xnor \U$9318 ( \9571 , \9546 , \9570 );
xor \U$9319 ( \9572 , \9536 , \9571 );
xnor \U$9320 ( \9573 , \9465 , \9572 );
not \U$9321 ( \9574 , \9573 );
xor \U$9322 ( \9575 , \9415 , \9574 );
not \U$9323 ( \9576 , \9236 );
and \U$9324 ( \9577 , \9576 , \9199 );
nor \U$9325 ( \9578 , \9577 , \9268 );
nor \U$9326 ( \9579 , \9576 , \9199 );
nor \U$9327 ( \9580 , \9578 , \9579 );
not \U$9328 ( \9581 , \9580 );
not \U$9329 ( \9582 , \9130 );
and \U$9330 ( \9583 , \9582 , \9166 );
nor \U$9331 ( \9584 , \9583 , \9101 );
nor \U$9332 ( \9585 , \9166 , \9582 );
nor \U$9333 ( \9586 , \9584 , \9585 );
not \U$9334 ( \9587 , \9586 );
not \U$9335 ( \9588 , \9587 );
or \U$9336 ( \9589 , \9581 , \9588 );
not \U$9337 ( \9590 , \9580 );
nand \U$9338 ( \9591 , \9586 , \9590 );
nand \U$9339 ( \9592 , \9589 , \9591 );
not \U$9340 ( \9593 , \6582 );
nand \U$9341 ( \9594 , \6592 , RIbe27b98_2);
not \U$9342 ( \9595 , \9594 );
or \U$9343 ( \9596 , \9593 , \9595 );
or \U$9344 ( \9597 , \9594 , \6601 );
nand \U$9345 ( \9598 , \9596 , \9597 );
not \U$9346 ( \9599 , RIbe28de0_41);
not \U$9347 ( \9600 , \6537 );
or \U$9348 ( \9601 , \9599 , \9600 );
nand \U$9349 ( \9602 , \7076 , RIbe29920_65);
nand \U$9350 ( \9603 , \9601 , \9602 );
and \U$9351 ( \9604 , \9603 , \6547 );
not \U$9352 ( \9605 , \9603 );
and \U$9353 ( \9606 , \9605 , \6551 );
nor \U$9354 ( \9607 , \9604 , \9606 );
xor \U$9355 ( \9608 , \9598 , \9607 );
not \U$9356 ( \9609 , RIbe27c10_3);
not \U$9357 ( \9610 , \6139 );
or \U$9358 ( \9611 , \9609 , \9610 );
nand \U$9359 ( \9612 , \6617 , RIbe28e58_42);
nand \U$9360 ( \9613 , \9611 , \9612 );
and \U$9361 ( \9614 , \9613 , \6144 );
not \U$9362 ( \9615 , \9613 );
and \U$9363 ( \9616 , \9615 , \6141 );
nor \U$9364 ( \9617 , \9614 , \9616 );
xor \U$9365 ( \9618 , \9608 , \9617 );
not \U$9366 ( \9619 , RIbe280c0_13);
not \U$9367 ( \9620 , \4764 );
or \U$9368 ( \9621 , \9619 , \9620 );
nand \U$9369 ( \9622 , \3689 , RIbe29830_63);
nand \U$9370 ( \9623 , \9621 , \9622 );
and \U$9371 ( \9624 , \9623 , \4346 );
not \U$9372 ( \9625 , \9623 );
and \U$9373 ( \9626 , \9625 , \2887 );
nor \U$9374 ( \9627 , \9624 , \9626 );
not \U$9375 ( \9628 , \9627 );
not \U$9376 ( \9629 , \9628 );
not \U$9377 ( \9630 , RIbe296c8_60);
not \U$9378 ( \9631 , \5094 );
or \U$9379 ( \9632 , \9630 , \9631 );
nand \U$9380 ( \9633 , \4027 , RIbe29650_59);
nand \U$9381 ( \9634 , \9632 , \9633 );
not \U$9382 ( \9635 , \9634 );
not \U$9383 ( \9636 , \3448 );
and \U$9384 ( \9637 , \9635 , \9636 );
and \U$9385 ( \9638 , \9634 , \3448 );
nor \U$9386 ( \9639 , \9637 , \9638 );
not \U$9387 ( \9640 , \9639 );
not \U$9388 ( \9641 , \9640 );
or \U$9389 ( \9642 , \9629 , \9641 );
nand \U$9390 ( \9643 , \9639 , \9627 );
nand \U$9391 ( \9644 , \9642 , \9643 );
not \U$9392 ( \9645 , RIbe28228_16);
not \U$9393 ( \9646 , \2898 );
or \U$9394 ( \9647 , \9645 , \9646 );
nand \U$9395 ( \9648 , \4284 , RIbe281b0_15);
nand \U$9396 ( \9649 , \9647 , \9648 );
not \U$9397 ( \9650 , \9649 );
not \U$9398 ( \9651 , \2379 );
and \U$9399 ( \9652 , \9650 , \9651 );
and \U$9400 ( \9653 , \9649 , \2379 );
nor \U$9401 ( \9654 , \9652 , \9653 );
xnor \U$9402 ( \9655 , \9644 , \9654 );
xor \U$9403 ( \9656 , \9618 , \9655 );
not \U$9404 ( \9657 , RIbe27d78_6);
not \U$9405 ( \9658 , \6630 );
or \U$9406 ( \9659 , \9657 , \9658 );
nand \U$9407 ( \9660 , \6634 , RIbe27d00_5);
nand \U$9408 ( \9661 , \9659 , \9660 );
not \U$9409 ( \9662 , \9661 );
not \U$9410 ( \9663 , \8252 );
and \U$9411 ( \9664 , \9662 , \9663 );
and \U$9412 ( \9665 , \9661 , \5457 );
nor \U$9413 ( \9666 , \9664 , \9665 );
not \U$9414 ( \9667 , RIbe290b0_47);
not \U$9415 ( \9668 , \4830 );
or \U$9416 ( \9669 , \9667 , \9668 );
nand \U$9417 ( \9670 , \5731 , RIbe29a88_68);
nand \U$9418 ( \9671 , \9669 , \9670 );
and \U$9419 ( \9672 , \9671 , \4586 );
not \U$9420 ( \9673 , \9671 );
and \U$9421 ( \9674 , \9673 , \4592 );
nor \U$9422 ( \9675 , \9672 , \9674 );
and \U$9423 ( \9676 , \9666 , \9675 );
not \U$9424 ( \9677 , \9666 );
not \U$9425 ( \9678 , \9675 );
and \U$9426 ( \9679 , \9677 , \9678 );
or \U$9427 ( \9680 , \9676 , \9679 );
not \U$9428 ( \9681 , RIbe29038_46);
not \U$9429 ( \9682 , \4317 );
or \U$9430 ( \9683 , \9681 , \9682 );
nand \U$9431 ( \9684 , \4809 , RIbe28fc0_45);
nand \U$9432 ( \9685 , \9683 , \9684 );
not \U$9433 ( \9686 , \9685 );
not \U$9434 ( \9687 , \4323 );
and \U$9435 ( \9688 , \9686 , \9687 );
and \U$9436 ( \9689 , \9685 , \4323 );
nor \U$9437 ( \9690 , \9688 , \9689 );
xnor \U$9438 ( \9691 , \9680 , \9690 );
xor \U$9439 ( \9692 , \9656 , \9691 );
not \U$9440 ( \9693 , \9692 );
xor \U$9441 ( \9694 , \9592 , \9693 );
xnor \U$9442 ( \9695 , \9575 , \9694 );
not \U$9443 ( \9696 , \8978 );
not \U$9444 ( \9697 , \8942 );
or \U$9445 ( \9698 , \9696 , \9697 );
or \U$9446 ( \9699 , \8942 , \8978 );
nand \U$9447 ( \9700 , \9699 , \8938 );
nand \U$9448 ( \9701 , \9698 , \9700 );
xor \U$9449 ( \9702 , \9695 , \9701 );
not \U$9450 ( \9703 , \9010 );
not \U$9451 ( \9704 , \9297 );
or \U$9452 ( \9705 , \9703 , \9704 );
not \U$9453 ( \9706 , \9010 );
not \U$9454 ( \9707 , \9297 );
nand \U$9455 ( \9708 , \9706 , \9707 );
nand \U$9456 ( \9709 , \9312 , \9708 );
nand \U$9457 ( \9710 , \9705 , \9709 );
xor \U$9458 ( \9711 , \9702 , \9710 );
not \U$9459 ( \9712 , \9711 );
not \U$9460 ( \9713 , \9712 );
or \U$9461 ( \9714 , \9399 , \9713 );
nand \U$9462 ( \9715 , \9711 , \9397 );
nand \U$9463 ( \9716 , \9714 , \9715 );
nand \U$9464 ( \9717 , \9313 , \9325 );
buf \U$9465 ( \9718 , \9318 );
and \U$9466 ( \9719 , \9717 , \9718 );
nor \U$9467 ( \9720 , \9313 , \9325 );
nor \U$9468 ( \9721 , \9719 , \9720 );
not \U$9469 ( \9722 , \9721 );
not \U$9470 ( \9723 , \9722 );
and \U$9471 ( \9724 , \9716 , \9723 );
not \U$9472 ( \9725 , \9716 );
and \U$9473 ( \9726 , \9725 , \9722 );
nor \U$9474 ( \9727 , \9724 , \9726 );
not \U$9475 ( \9728 , \9727 );
or \U$9476 ( \9729 , \9340 , \9728 );
or \U$9477 ( \9730 , \9727 , \9339 );
nand \U$9478 ( \9731 , \9729 , \9730 );
not \U$9479 ( \9732 , \9731 );
not \U$9480 ( \9733 , \9732 );
or \U$9481 ( \9734 , \9335 , \9733 );
nand \U$9482 ( \9735 , \9731 , \9333 );
nand \U$9483 ( \9736 , \9734 , \9735 );
xor \U$9484 ( \9737 , \8680 , \8673 );
xnor \U$9485 ( \9738 , \9737 , \8689 );
xor \U$9486 ( \9739 , \8114 , \8144 );
xor \U$9487 ( \9740 , \9739 , \8185 );
and \U$9488 ( \9741 , \8222 , \8297 );
not \U$9489 ( \9742 , \8222 );
and \U$9490 ( \9743 , \9742 , \8298 );
nor \U$9491 ( \9744 , \9741 , \9743 );
not \U$9492 ( \9745 , \9744 );
not \U$9493 ( \9746 , \8263 );
and \U$9494 ( \9747 , \9745 , \9746 );
and \U$9495 ( \9748 , \9744 , \8263 );
nor \U$9496 ( \9749 , \9747 , \9748 );
not \U$9497 ( \9750 , \9749 );
or \U$9498 ( \9751 , \9740 , \9750 );
xor \U$9499 ( \9752 , \8332 , \8362 );
xor \U$9500 ( \9753 , \9752 , \8396 );
nand \U$9501 ( \9754 , \9751 , \9753 );
nand \U$9502 ( \9755 , \9750 , \9740 );
nand \U$9503 ( \9756 , \9754 , \9755 );
xor \U$9504 ( \9757 , \8457 , \8462 );
xor \U$9505 ( \9758 , \9757 , \8465 );
xor \U$9506 ( \9759 , \9756 , \9758 );
xor \U$9507 ( \9760 , \8429 , \8417 );
buf \U$9508 ( \9761 , \8414 );
and \U$9509 ( \9762 , \9760 , \9761 );
not \U$9510 ( \9763 , \9760 );
not \U$9511 ( \9764 , \9761 );
and \U$9512 ( \9765 , \9763 , \9764 );
nor \U$9513 ( \9766 , \9762 , \9765 );
and \U$9514 ( \9767 , \9759 , \9766 );
and \U$9515 ( \9768 , \9756 , \9758 );
or \U$9516 ( \9769 , \9767 , \9768 );
not \U$9517 ( \9770 , RIbe2a988_100);
not \U$9518 ( \9771 , \325 );
or \U$9519 ( \9772 , \9770 , \9771 );
nand \U$9520 ( \9773 , RIbe2a910_99, \330 );
nand \U$9521 ( \9774 , \9772 , \9773 );
not \U$9522 ( \9775 , \9774 );
nand \U$9523 ( \9776 , \338 , \9775 );
nand \U$9524 ( \9777 , \9774 , \1374 );
and \U$9525 ( \9778 , \9776 , \9777 );
nand \U$9526 ( \9779 , RIbe29380_53, RIbe2a550_91);
nor \U$9527 ( \9780 , \9778 , \9779 );
not \U$9528 ( \9781 , RIbe29fb0_79);
not \U$9529 ( \9782 , \546 );
or \U$9530 ( \9783 , \9781 , \9782 );
nand \U$9531 ( \9784 , \553 , RIbe29e48_76);
nand \U$9532 ( \9785 , \9783 , \9784 );
xor \U$9533 ( \9786 , \9785 , \424 );
not \U$9534 ( \9787 , \9786 );
and \U$9535 ( \9788 , \1161 , RIbe29bf0_71);
and \U$9536 ( \9789 , \1165 , RIbe28f48_44);
nor \U$9537 ( \9790 , \9788 , \9789 );
and \U$9538 ( \9791 , \9790 , \1011 );
not \U$9539 ( \9792 , \9790 );
and \U$9540 ( \9793 , \9792 , \1813 );
nor \U$9541 ( \9794 , \9791 , \9793 );
not \U$9542 ( \9795 , \9794 );
nand \U$9543 ( \9796 , \9787 , \9795 );
not \U$9544 ( \9797 , \9794 );
not \U$9545 ( \9798 , \9786 );
or \U$9546 ( \9799 , \9797 , \9798 );
not \U$9547 ( \9800 , \8173 );
not \U$9548 ( \9801 , RIbe29c68_72);
not \U$9549 ( \9802 , \9801 );
and \U$9550 ( \9803 , \9800 , \9802 );
and \U$9551 ( \9804 , \2531 , RIbe29dd0_75);
nor \U$9552 ( \9805 , \9803 , \9804 );
and \U$9553 ( \9806 , \9805 , \564 );
not \U$9554 ( \9807 , \9805 );
and \U$9555 ( \9808 , \9807 , \3959 );
nor \U$9556 ( \9809 , \9806 , \9808 );
nand \U$9557 ( \9810 , \9799 , \9809 );
nand \U$9558 ( \9811 , \9796 , \9810 );
xor \U$9559 ( \9812 , \9780 , \9811 );
not \U$9560 ( \9813 , RIbe2a370_87);
not \U$9561 ( \9814 , \1252 );
or \U$9562 ( \9815 , \9813 , \9814 );
not \U$9563 ( \9816 , \285 );
nand \U$9564 ( \9817 , \9816 , RIbe2a2f8_86);
nand \U$9565 ( \9818 , \9815 , \9817 );
not \U$9566 ( \9819 , \9818 );
not \U$9567 ( \9820 , \300 );
and \U$9568 ( \9821 , \9819 , \9820 );
and \U$9569 ( \9822 , \9818 , \300 );
nor \U$9570 ( \9823 , \9821 , \9822 );
not \U$9571 ( \9824 , \9823 );
and \U$9572 ( \9825 , \260 , RIbe2b5b8_126);
and \U$9573 ( \9826 , \264 , RIbe2a3e8_88);
nor \U$9574 ( \9827 , \9825 , \9826 );
and \U$9575 ( \9828 , \9827 , \1363 );
not \U$9576 ( \9829 , \9827 );
and \U$9577 ( \9830 , \9829 , \1362 );
nor \U$9578 ( \9831 , \9828 , \9830 );
not \U$9579 ( \9832 , \9831 );
or \U$9580 ( \9833 , \9824 , \9832 );
not \U$9581 ( \9834 , RIbe2acd0_107);
not \U$9582 ( \9835 , \1773 );
or \U$9583 ( \9836 , \9834 , \9835 );
nand \U$9584 ( \9837 , \429 , RIbe2a028_80);
nand \U$9585 ( \9838 , \9836 , \9837 );
and \U$9586 ( \9839 , \9838 , \306 );
not \U$9587 ( \9840 , \9838 );
and \U$9588 ( \9841 , \9840 , \1547 );
nor \U$9589 ( \9842 , \9839 , \9841 );
nand \U$9590 ( \9843 , \9833 , \9842 );
not \U$9591 ( \9844 , \9823 );
not \U$9592 ( \9845 , \9831 );
nand \U$9593 ( \9846 , \9844 , \9845 );
nand \U$9594 ( \9847 , \9843 , \9846 );
and \U$9595 ( \9848 , \9812 , \9847 );
and \U$9596 ( \9849 , \9780 , \9811 );
or \U$9597 ( \9850 , \9848 , \9849 );
not \U$9598 ( \9851 , RIbe29a88_68);
not \U$9599 ( \9852 , \8199 );
or \U$9600 ( \9853 , \9851 , \9852 );
nand \U$9601 ( \9854 , \7958 , RIbe27d78_6);
nand \U$9602 ( \9855 , \9853 , \9854 );
and \U$9603 ( \9856 , \9855 , \6572 );
not \U$9604 ( \9857 , \9855 );
and \U$9605 ( \9858 , \9857 , \7293 );
nor \U$9606 ( \9859 , \9856 , \9858 );
not \U$9607 ( \9860 , RIbe28fc0_45);
not \U$9608 ( \9861 , \6592 );
or \U$9609 ( \9862 , \9860 , \9861 );
nand \U$9610 ( \9863 , \7278 , RIbe290b0_47);
nand \U$9611 ( \9864 , \9862 , \9863 );
not \U$9612 ( \9865 , \9864 );
not \U$9613 ( \9866 , \6602 );
and \U$9614 ( \9867 , \9865 , \9866 );
not \U$9615 ( \9868 , \6601 );
and \U$9616 ( \9869 , \9864 , \9868 );
nor \U$9617 ( \9870 , \9867 , \9869 );
nand \U$9618 ( \9871 , \9859 , \9870 );
not \U$9619 ( \9872 , RIbe27d00_5);
not \U$9620 ( \9873 , \7299 );
or \U$9621 ( \9874 , \9872 , \9873 );
not \U$9622 ( \9875 , \6984 );
nand \U$9623 ( \9876 , \9875 , RIbe27c10_3);
nand \U$9624 ( \9877 , \9874 , \9876 );
not \U$9625 ( \9878 , \9877 );
not \U$9626 ( \9879 , \6992 );
and \U$9627 ( \9880 , \9878 , \9879 );
and \U$9628 ( \9881 , \9877 , \6992 );
nor \U$9629 ( \9882 , \9880 , \9881 );
not \U$9630 ( \9883 , \9882 );
and \U$9631 ( \9884 , \9871 , \9883 );
nor \U$9632 ( \9885 , \9859 , \9870 );
nor \U$9633 ( \9886 , \9884 , \9885 );
not \U$9634 ( \9887 , \9886 );
not \U$9635 ( \9888 , RIbe28e58_42);
not \U$9636 ( \9889 , \7975 );
or \U$9637 ( \9890 , \9888 , \9889 );
not \U$9638 ( \9891 , \7980 );
nand \U$9639 ( \9892 , \9891 , RIbe28de0_41);
nand \U$9640 ( \9893 , \9890 , \9892 );
and \U$9641 ( \9894 , \9893 , \6948 );
not \U$9642 ( \9895 , \9893 );
not \U$9643 ( \9896 , \6948 );
and \U$9644 ( \9897 , \9895 , \9896 );
nor \U$9645 ( \9898 , \9894 , \9897 );
nand \U$9646 ( \9899 , RIbe2a460_89, RIbe2adc0_109);
nand \U$9647 ( \9900 , \9899 , RIbe2a4d8_90);
not \U$9648 ( \9901 , \9900 );
buf \U$9649 ( \9902 , \9901 );
not \U$9650 ( \9903 , \9902 );
not \U$9651 ( \9904 , \9903 );
nand \U$9652 ( \9905 , \9898 , \9904 );
not \U$9653 ( \9906 , \8077 );
not \U$9654 ( \9907 , RIbe29920_65);
not \U$9655 ( \9908 , \8276 );
not \U$9656 ( \9909 , \9908 );
not \U$9657 ( \9910 , \9909 );
or \U$9658 ( \9911 , \9907 , \9910 );
buf \U$9659 ( \9912 , \8274 );
buf \U$9660 ( \9913 , \9912 );
buf \U$9661 ( \9914 , \9913 );
nand \U$9662 ( \9915 , \9914 , RIbe27b98_2);
nand \U$9663 ( \9916 , \9911 , \9915 );
not \U$9664 ( \9917 , \9916 );
or \U$9665 ( \9918 , \9906 , \9917 );
or \U$9666 ( \9919 , \9916 , \8077 );
nand \U$9667 ( \9920 , \9918 , \9919 );
and \U$9668 ( \9921 , \9905 , \9920 );
nor \U$9669 ( \9922 , \9898 , \9904 );
nor \U$9670 ( \9923 , \9921 , \9922 );
not \U$9671 ( \9924 , \9923 );
or \U$9672 ( \9925 , \9887 , \9924 );
not \U$9673 ( \9926 , RIbe29650_59);
not \U$9674 ( \9927 , \6536 );
or \U$9675 ( \9928 , \9926 , \9927 );
nand \U$9676 ( \9929 , \6540 , RIbe29038_46);
nand \U$9677 ( \9930 , \9928 , \9929 );
and \U$9678 ( \9931 , \9930 , \6552 );
not \U$9679 ( \9932 , \9930 );
not \U$9680 ( \9933 , \6546 );
and \U$9681 ( \9934 , \9932 , \9933 );
nor \U$9682 ( \9935 , \9931 , \9934 );
not \U$9683 ( \9936 , RIbe29830_63);
not \U$9684 ( \9937 , \8231 );
or \U$9685 ( \9938 , \9936 , \9937 );
not \U$9686 ( \9939 , \6615 );
nand \U$9687 ( \9940 , \9939 , RIbe296c8_60);
nand \U$9688 ( \9941 , \9938 , \9940 );
and \U$9689 ( \9942 , \9941 , \7501 );
not \U$9690 ( \9943 , \9941 );
not \U$9691 ( \9944 , \6620 );
and \U$9692 ( \9945 , \9943 , \9944 );
nor \U$9693 ( \9946 , \9942 , \9945 );
xor \U$9694 ( \9947 , \9935 , \9946 );
not \U$9695 ( \9948 , RIbe281b0_15);
not \U$9696 ( \9949 , \5455 );
or \U$9697 ( \9950 , \9948 , \9949 );
nand \U$9698 ( \9951 , \7100 , RIbe280c0_13);
nand \U$9699 ( \9952 , \9950 , \9951 );
and \U$9700 ( \9953 , \9952 , \6117 );
not \U$9701 ( \9954 , \9952 );
and \U$9702 ( \9955 , \9954 , \6637 );
nor \U$9703 ( \9956 , \9953 , \9955 );
and \U$9704 ( \9957 , \9947 , \9956 );
and \U$9705 ( \9958 , \9935 , \9946 );
or \U$9706 ( \9959 , \9957 , \9958 );
nand \U$9707 ( \9960 , \9925 , \9959 );
not \U$9708 ( \9961 , \9923 );
not \U$9709 ( \9962 , \9886 );
nand \U$9710 ( \9963 , \9961 , \9962 );
nand \U$9711 ( \9964 , \9960 , \9963 );
xor \U$9712 ( \9965 , \9850 , \9964 );
not \U$9713 ( \9966 , RIbe28ed0_43);
not \U$9714 ( \9967 , \1143 );
or \U$9715 ( \9968 , \9966 , \9967 );
nand \U$9716 ( \9969 , \1147 , RIbe27fd0_11);
nand \U$9717 ( \9970 , \9968 , \9969 );
and \U$9718 ( \9971 , \9970 , \3993 );
not \U$9719 ( \9972 , \9970 );
and \U$9720 ( \9973 , \9972 , \1157 );
nor \U$9721 ( \9974 , \9971 , \9973 );
not \U$9722 ( \9975 , RIbe27f58_10);
not \U$9723 ( \9976 , \5476 );
or \U$9724 ( \9977 , \9975 , \9976 );
nand \U$9725 ( \9978 , \1454 , RIbe27e68_8);
nand \U$9726 ( \9979 , \9977 , \9978 );
and \U$9727 ( \9980 , \9979 , \1309 );
not \U$9728 ( \9981 , \9979 );
and \U$9729 ( \9982 , \9981 , \1458 );
nor \U$9730 ( \9983 , \9980 , \9982 );
or \U$9731 ( \9984 , \9974 , \9983 );
not \U$9732 ( \9985 , RIbe28660_25);
not \U$9733 ( \9986 , \1112 );
or \U$9734 ( \9987 , \9985 , \9986 );
nand \U$9735 ( \9988 , \5467 , RIbe285e8_24);
nand \U$9736 ( \9989 , \9987 , \9988 );
not \U$9737 ( \9990 , \9989 );
not \U$9738 ( \9991 , \6831 );
and \U$9739 ( \9992 , \9990 , \9991 );
and \U$9740 ( \9993 , \9989 , \2563 );
nor \U$9741 ( \9994 , \9992 , \9993 );
not \U$9742 ( \9995 , \9994 );
nand \U$9743 ( \9996 , \9984 , \9995 );
nand \U$9744 ( \9997 , \9974 , \9983 );
nand \U$9745 ( \9998 , \9996 , \9997 );
not \U$9746 ( \9999 , RIbe28b10_35);
not \U$9747 ( \10000 , \3685 );
or \U$9748 ( \10001 , \9999 , \10000 );
nand \U$9749 ( \10002 , \3689 , RIbe28b88_36);
nand \U$9750 ( \10003 , \10001 , \10002 );
and \U$9751 ( \10004 , \10003 , \3290 );
not \U$9752 ( \10005 , \10003 );
and \U$9753 ( \10006 , \10005 , \2887 );
nor \U$9754 ( \10007 , \10004 , \10006 );
not \U$9755 ( \10008 , \10007 );
not \U$9756 ( \10009 , RIbe28408_20);
not \U$9757 ( \10010 , \2570 );
not \U$9758 ( \10011 , \10010 );
or \U$9759 ( \10012 , \10009 , \10011 );
nand \U$9760 ( \10013 , \2901 , RIbe28390_19);
nand \U$9761 ( \10014 , \10012 , \10013 );
not \U$9762 ( \10015 , \10014 );
not \U$9763 ( \10016 , \2576 );
and \U$9764 ( \10017 , \10015 , \10016 );
and \U$9765 ( \10018 , \10014 , \2379 );
nor \U$9766 ( \10019 , \10017 , \10018 );
not \U$9767 ( \10020 , \10019 );
not \U$9768 ( \10021 , \10020 );
or \U$9769 ( \10022 , \10008 , \10021 );
or \U$9770 ( \10023 , \10020 , \10007 );
not \U$9771 ( \10024 , \4065 );
not \U$9772 ( \10025 , RIbe28480_21);
not \U$9773 ( \10026 , \10025 );
and \U$9774 ( \10027 , \10024 , \10026 );
and \U$9775 ( \10028 , \4295 , RIbe287c8_28);
nor \U$9776 ( \10029 , \10027 , \10028 );
and \U$9777 ( \10030 , \10029 , \3516 );
not \U$9778 ( \10031 , \10029 );
and \U$9779 ( \10032 , \10031 , \1277 );
nor \U$9780 ( \10033 , \10030 , \10032 );
nand \U$9781 ( \10034 , \10023 , \10033 );
nand \U$9782 ( \10035 , \10022 , \10034 );
xor \U$9783 ( \10036 , \9998 , \10035 );
not \U$9784 ( \10037 , RIbe29290_51);
not \U$9785 ( \10038 , \5094 );
or \U$9786 ( \10039 , \10037 , \10038 );
nand \U$9787 ( \10040 , \7438 , RIbe28a20_33);
nand \U$9788 ( \10041 , \10039 , \10040 );
and \U$9789 ( \10042 , \10041 , \3471 );
not \U$9790 ( \10043 , \10041 );
and \U$9791 ( \10044 , \10043 , \3448 );
nor \U$9792 ( \10045 , \10042 , \10044 );
not \U$9793 ( \10046 , RIbe29560_57);
not \U$9794 ( \10047 , \5727 );
or \U$9795 ( \10048 , \10046 , \10047 );
nand \U$9796 ( \10049 , \5052 , RIbe28228_16);
nand \U$9797 ( \10050 , \10048 , \10049 );
and \U$9798 ( \10051 , \10050 , \4586 );
not \U$9799 ( \10052 , \10050 );
and \U$9800 ( \10053 , \10052 , \4592 );
nor \U$9801 ( \10054 , \10051 , \10053 );
xor \U$9802 ( \10055 , \10045 , \10054 );
not \U$9803 ( \10056 , RIbe289a8_32);
not \U$9804 ( \10057 , \4317 );
or \U$9805 ( \10058 , \10056 , \10057 );
nand \U$9806 ( \10059 , \4600 , RIbe28930_31);
nand \U$9807 ( \10060 , \10058 , \10059 );
and \U$9808 ( \10061 , \10060 , \4007 );
not \U$9809 ( \10062 , \10060 );
and \U$9810 ( \10063 , \10062 , \4323 );
nor \U$9811 ( \10064 , \10061 , \10063 );
and \U$9812 ( \10065 , \10055 , \10064 );
and \U$9813 ( \10066 , \10045 , \10054 );
or \U$9814 ( \10067 , \10065 , \10066 );
and \U$9815 ( \10068 , \10036 , \10067 );
and \U$9816 ( \10069 , \9998 , \10035 );
or \U$9817 ( \10070 , \10068 , \10069 );
and \U$9818 ( \10071 , \9965 , \10070 );
and \U$9819 ( \10072 , \9850 , \9964 );
or \U$9820 ( \10073 , \10071 , \10072 );
xor \U$9821 ( \10074 , \8124 , \8130 );
xor \U$9822 ( \10075 , \10074 , \8141 );
not \U$9823 ( \10076 , \8114 );
or \U$9824 ( \10077 , \10075 , \10076 );
not \U$9825 ( \10078 , \8183 );
not \U$9826 ( \10079 , \10078 );
not \U$9827 ( \10080 , \8156 );
or \U$9828 ( \10081 , \10079 , \10080 );
nand \U$9829 ( \10082 , \8155 , \8183 );
nand \U$9830 ( \10083 , \10081 , \10082 );
and \U$9831 ( \10084 , \10083 , \8167 );
not \U$9832 ( \10085 , \10083 );
and \U$9833 ( \10086 , \10085 , \8166 );
nor \U$9834 ( \10087 , \10084 , \10086 );
nand \U$9835 ( \10088 , \10077 , \10087 );
nand \U$9836 ( \10089 , \10075 , \10076 );
nand \U$9837 ( \10090 , \10088 , \10089 );
not \U$9838 ( \10091 , \10090 );
not \U$9839 ( \10092 , \10091 );
not \U$9840 ( \10093 , \10092 );
xor \U$9841 ( \10094 , \8208 , \8197 );
xor \U$9842 ( \10095 , \10094 , \8219 );
xor \U$9843 ( \10096 , \8261 , \8255 );
xor \U$9844 ( \10097 , \10096 , \8241 );
nand \U$9845 ( \10098 , \10095 , \10097 );
xor \U$9846 ( \10099 , \8283 , \8294 );
xnor \U$9847 ( \10100 , \10099 , \8272 );
and \U$9848 ( \10101 , \10098 , \10100 );
nor \U$9849 ( \10102 , \10095 , \10097 );
nor \U$9850 ( \10103 , \10101 , \10102 );
not \U$9851 ( \10104 , \10103 );
not \U$9852 ( \10105 , \10104 );
or \U$9853 ( \10106 , \10093 , \10105 );
not \U$9854 ( \10107 , \10091 );
not \U$9855 ( \10108 , \10103 );
or \U$9856 ( \10109 , \10107 , \10108 );
xor \U$9857 ( \10110 , \8374 , \8383 );
xor \U$9858 ( \10111 , \10110 , \8393 );
xor \U$9859 ( \10112 , \8329 , \8318 );
buf \U$9860 ( \10113 , \8309 );
xor \U$9861 ( \10114 , \10112 , \10113 );
or \U$9862 ( \10115 , \10111 , \10114 );
xor \U$9863 ( \10116 , \8359 , \8350 );
xor \U$9864 ( \10117 , \10116 , \8339 );
not \U$9865 ( \10118 , \10117 );
nand \U$9866 ( \10119 , \10115 , \10118 );
nand \U$9867 ( \10120 , \10111 , \10114 );
nand \U$9868 ( \10121 , \10119 , \10120 );
nand \U$9869 ( \10122 , \10109 , \10121 );
nand \U$9870 ( \10123 , \10106 , \10122 );
xor \U$9871 ( \10124 , \10073 , \10123 );
not \U$9872 ( \10125 , \8082 );
not \U$9873 ( \10126 , \8079 );
or \U$9874 ( \10127 , \10125 , \10126 );
or \U$9875 ( \10128 , \8082 , \8079 );
nand \U$9876 ( \10129 , \10127 , \10128 );
xor \U$9877 ( \10130 , \10129 , \8076 );
not \U$9878 ( \10131 , \10130 );
xor \U$9879 ( \10132 , \8056 , \8063 );
xnor \U$9880 ( \10133 , \10132 , \8062 );
xnor \U$9881 ( \10134 , \10133 , \8055 );
or \U$9882 ( \10135 , \10131 , \10134 );
not \U$9883 ( \10136 , \8098 );
not \U$9884 ( \10137 , \8106 );
or \U$9885 ( \10138 , \10136 , \10137 );
or \U$9886 ( \10139 , \8106 , \8098 );
nand \U$9887 ( \10140 , \10138 , \10139 );
and \U$9888 ( \10141 , \10140 , \8095 );
not \U$9889 ( \10142 , \10140 );
and \U$9890 ( \10143 , \10142 , \8094 );
nor \U$9891 ( \10144 , \10141 , \10143 );
nand \U$9892 ( \10145 , \10135 , \10144 );
nand \U$9893 ( \10146 , \10131 , \10134 );
nand \U$9894 ( \10147 , \10145 , \10146 );
and \U$9895 ( \10148 , \10124 , \10147 );
and \U$9896 ( \10149 , \10073 , \10123 );
or \U$9897 ( \10150 , \10148 , \10149 );
not \U$9898 ( \10151 , \10150 );
xor \U$9899 ( \10152 , \8109 , \8086 );
xnor \U$9900 ( \10153 , \10152 , \8070 );
not \U$9901 ( \10154 , \10153 );
xor \U$9902 ( \10155 , \8188 , \8301 );
xor \U$9903 ( \10156 , \10155 , \8399 );
nand \U$9904 ( \10157 , \10154 , \10156 );
nand \U$9905 ( \10158 , \10151 , \10157 );
and \U$9906 ( \10159 , \9769 , \10158 );
not \U$9907 ( \10160 , \10150 );
nor \U$9908 ( \10161 , \10160 , \10157 );
nor \U$9909 ( \10162 , \10159 , \10161 );
xor \U$9910 ( \10163 , \8402 , \8112 );
xnor \U$9911 ( \10164 , \10163 , \8432 );
xor \U$9912 ( \10165 , \8049 , \7753 );
or \U$9913 ( \10166 , \10164 , \10165 );
not \U$9914 ( \10167 , \8469 );
not \U$9915 ( \10168 , \8511 );
or \U$9916 ( \10169 , \10167 , \10168 );
nand \U$9917 ( \10170 , \8510 , \8468 );
nand \U$9918 ( \10171 , \10169 , \10170 );
xnor \U$9919 ( \10172 , \10171 , \8455 );
and \U$9920 ( \10173 , \10166 , \10172 );
and \U$9921 ( \10174 , \10165 , \10164 );
nor \U$9922 ( \10175 , \10173 , \10174 );
xor \U$9923 ( \10176 , \10162 , \10175 );
xor \U$9924 ( \10177 , \8616 , \8642 );
xnor \U$9925 ( \10178 , \10177 , \8658 );
and \U$9926 ( \10179 , \10176 , \10178 );
and \U$9927 ( \10180 , \10162 , \10175 );
or \U$9928 ( \10181 , \10179 , \10180 );
xor \U$9929 ( \10182 , \9738 , \10181 );
not \U$9930 ( \10183 , \8517 );
not \U$9931 ( \10184 , \8660 );
or \U$9932 ( \10185 , \10183 , \10184 );
or \U$9933 ( \10186 , \8660 , \8517 );
nand \U$9934 ( \10187 , \10185 , \10186 );
and \U$9935 ( \10188 , \10187 , \8663 );
not \U$9936 ( \10189 , \10187 );
and \U$9937 ( \10190 , \10189 , \8593 );
or \U$9938 ( \10191 , \10188 , \10190 );
and \U$9939 ( \10192 , \10182 , \10191 );
and \U$9940 ( \10193 , \9738 , \10181 );
or \U$9941 ( \10194 , \10192 , \10193 );
not \U$9942 ( \10195 , \10194 );
xor \U$9943 ( \10196 , \7686 , \8665 );
and \U$9944 ( \10197 , \10196 , \8930 );
not \U$9945 ( \10198 , \10196 );
not \U$9946 ( \10199 , \8930 );
and \U$9947 ( \10200 , \10198 , \10199 );
nor \U$9948 ( \10201 , \10197 , \10200 );
nand \U$9949 ( \10202 , \10195 , \10201 );
not \U$9950 ( \10203 , \10202 );
not \U$9951 ( \10204 , \10203 );
not \U$9952 ( \10205 , \8933 );
not \U$9953 ( \10206 , \9332 );
or \U$9954 ( \10207 , \10205 , \10206 );
or \U$9955 ( \10208 , \9332 , \8933 );
nand \U$9956 ( \10209 , \10207 , \10208 );
not \U$9957 ( \10210 , \10209 );
not \U$9958 ( \10211 , \10210 );
or \U$9959 ( \10212 , \10204 , \10211 );
nand \U$9960 ( \10213 , \10209 , \10202 );
nand \U$9961 ( \10214 , \10212 , \10213 );
not \U$9962 ( \10215 , \9727 );
nand \U$9963 ( \10216 , \10215 , \9339 );
not \U$9964 ( \10217 , \9398 );
not \U$9965 ( \10218 , \9722 );
or \U$9966 ( \10219 , \10217 , \10218 );
not \U$9967 ( \10220 , \9397 );
not \U$9968 ( \10221 , \9721 );
or \U$9969 ( \10222 , \10220 , \10221 );
nand \U$9970 ( \10223 , \10222 , \9711 );
nand \U$9971 ( \10224 , \10219 , \10223 );
and \U$9972 ( \10225 , \9396 , \9366 );
not \U$9973 ( \10226 , \9396 );
and \U$9974 ( \10227 , \10226 , \9365 );
nor \U$9975 ( \10228 , \10225 , \10227 );
and \U$9976 ( \10229 , \10228 , \9359 );
xor \U$9977 ( \10230 , \9695 , \9701 );
and \U$9978 ( \10231 , \10230 , \9710 );
and \U$9979 ( \10232 , \9695 , \9701 );
or \U$9980 ( \10233 , \10231 , \10232 );
xor \U$9981 ( \10234 , \10229 , \10233 );
not \U$9982 ( \10235 , \9391 );
not \U$9983 ( \10236 , \9371 );
or \U$9984 ( \10237 , \10235 , \10236 );
or \U$9985 ( \10238 , \9391 , \9371 );
nand \U$9986 ( \10239 , \10238 , \9365 );
nand \U$9987 ( \10240 , \10237 , \10239 );
not \U$9988 ( \10241 , \9415 );
not \U$9989 ( \10242 , \9574 );
or \U$9990 ( \10243 , \10241 , \10242 );
not \U$9991 ( \10244 , \9694 );
not \U$9992 ( \10245 , \9415 );
nand \U$9993 ( \10246 , \10245 , \9573 );
nand \U$9994 ( \10247 , \10244 , \10246 );
nand \U$9995 ( \10248 , \10243 , \10247 );
not \U$9996 ( \10249 , \10248 );
not \U$9997 ( \10250 , \9358 );
nor \U$9998 ( \10251 , \9344 , \9353 );
not \U$9999 ( \10252 , \10251 );
and \U$10000 ( \10253 , \10250 , \10252 );
and \U$10001 ( \10254 , \9344 , \9353 );
nor \U$10002 ( \10255 , \10253 , \10254 );
not \U$10003 ( \10256 , \10255 );
not \U$10004 ( \10257 , RIbe28fc0_45);
not \U$10005 ( \10258 , \5058 );
or \U$10006 ( \10259 , \10257 , \10258 );
nand \U$10007 ( \10260 , \4600 , RIbe290b0_47);
nand \U$10008 ( \10261 , \10259 , \10260 );
and \U$10009 ( \10262 , \10261 , \4603 );
not \U$10010 ( \10263 , \10261 );
and \U$10011 ( \10264 , \10263 , \4323 );
nor \U$10012 ( \10265 , \10262 , \10264 );
not \U$10013 ( \10266 , RIbe27d00_5);
not \U$10014 ( \10267 , \5455 );
or \U$10015 ( \10268 , \10266 , \10267 );
buf \U$10016 ( \10269 , \5749 );
nand \U$10017 ( \10270 , \10269 , RIbe27c10_3);
nand \U$10018 ( \10271 , \10268 , \10270 );
not \U$10019 ( \10272 , \5754 );
and \U$10020 ( \10273 , \10271 , \10272 );
not \U$10021 ( \10274 , \10271 );
and \U$10022 ( \10275 , \10274 , \5754 );
nor \U$10023 ( \10276 , \10273 , \10275 );
not \U$10024 ( \10277 , RIbe29a88_68);
not \U$10025 ( \10278 , \5727 );
or \U$10026 ( \10279 , \10277 , \10278 );
nand \U$10027 ( \10280 , \5731 , RIbe27d78_6);
nand \U$10028 ( \10281 , \10279 , \10280 );
and \U$10029 ( \10282 , \10281 , \4586 );
not \U$10030 ( \10283 , \10281 );
and \U$10031 ( \10284 , \10283 , \4592 );
nor \U$10032 ( \10285 , \10282 , \10284 );
xor \U$10033 ( \10286 , \10276 , \10285 );
xor \U$10034 ( \10287 , \10265 , \10286 );
xor \U$10035 ( \10288 , \9501 , \9535 );
and \U$10036 ( \10289 , \10288 , \9571 );
and \U$10037 ( \10290 , \9501 , \9535 );
or \U$10038 ( \10291 , \10289 , \10290 );
xor \U$10039 ( \10292 , \10287 , \10291 );
xor \U$10040 ( \10293 , \9618 , \9655 );
and \U$10041 ( \10294 , \10293 , \9691 );
and \U$10042 ( \10295 , \9618 , \9655 );
or \U$10043 ( \10296 , \10294 , \10295 );
xor \U$10044 ( \10297 , \10292 , \10296 );
not \U$10045 ( \10298 , \10297 );
and \U$10046 ( \10299 , \10256 , \10298 );
and \U$10047 ( \10300 , \10255 , \10297 );
nor \U$10048 ( \10301 , \10299 , \10300 );
not \U$10049 ( \10302 , \10301 );
or \U$10050 ( \10303 , \10249 , \10302 );
or \U$10051 ( \10304 , \10248 , \10301 );
nand \U$10052 ( \10305 , \10303 , \10304 );
xor \U$10053 ( \10306 , \10240 , \10305 );
not \U$10054 ( \10307 , \9440 );
xor \U$10055 ( \10308 , \9403 , \9407 );
and \U$10056 ( \10309 , \10308 , \9414 );
and \U$10057 ( \10310 , \9403 , \9407 );
or \U$10058 ( \10311 , \10309 , \10310 );
xor \U$10059 ( \10312 , \10307 , \10311 );
xor \U$10060 ( \10313 , \9447 , \9451 );
and \U$10061 ( \10314 , \10313 , \9459 );
and \U$10062 ( \10315 , \9447 , \9451 );
or \U$10063 ( \10316 , \10314 , \10315 );
xor \U$10064 ( \10317 , \10312 , \10316 );
not \U$10065 ( \10318 , \10317 );
xor \U$10066 ( \10319 , \9378 , \9385 );
and \U$10067 ( \10320 , \10319 , \9390 );
and \U$10068 ( \10321 , \9378 , \9385 );
or \U$10069 ( \10322 , \10320 , \10321 );
not \U$10070 ( \10323 , \9590 );
not \U$10071 ( \10324 , \9587 );
or \U$10072 ( \10325 , \10323 , \10324 );
not \U$10073 ( \10326 , \9580 );
not \U$10074 ( \10327 , \9586 );
or \U$10075 ( \10328 , \10326 , \10327 );
nand \U$10076 ( \10329 , \10328 , \9692 );
nand \U$10077 ( \10330 , \10325 , \10329 );
xor \U$10078 ( \10331 , \10322 , \10330 );
not \U$10079 ( \10332 , \9441 );
not \U$10080 ( \10333 , \9461 );
or \U$10081 ( \10334 , \10332 , \10333 );
or \U$10082 ( \10335 , \9461 , \9441 );
nand \U$10083 ( \10336 , \10335 , \9572 );
nand \U$10084 ( \10337 , \10334 , \10336 );
xor \U$10085 ( \10338 , \10331 , \10337 );
not \U$10086 ( \10339 , \10338 );
not \U$10087 ( \10340 , \10339 );
or \U$10088 ( \10341 , \10318 , \10340 );
not \U$10089 ( \10342 , \10317 );
nand \U$10090 ( \10343 , \10342 , \10338 );
nand \U$10091 ( \10344 , \10341 , \10343 );
not \U$10092 ( \10345 , RIbe29920_65);
not \U$10093 ( \10346 , \6536 );
or \U$10094 ( \10347 , \10345 , \10346 );
buf \U$10095 ( \10348 , \6884 );
nand \U$10096 ( \10349 , \10348 , RIbe27b98_2);
nand \U$10097 ( \10350 , \10347 , \10349 );
or \U$10098 ( \10351 , \10350 , \7546 );
nand \U$10099 ( \10352 , \10350 , \6551 );
nand \U$10100 ( \10353 , \10351 , \10352 );
and \U$10101 ( \10354 , \10353 , \8957 );
not \U$10102 ( \10355 , \10353 );
and \U$10103 ( \10356 , \10355 , \6601 );
nor \U$10104 ( \10357 , \10354 , \10356 );
not \U$10105 ( \10358 , \10357 );
not \U$10106 ( \10359 , RIbe28e58_42);
not \U$10107 ( \10360 , \6139 );
or \U$10108 ( \10361 , \10359 , \10360 );
nand \U$10109 ( \10362 , \9939 , RIbe28de0_41);
nand \U$10110 ( \10363 , \10361 , \10362 );
and \U$10111 ( \10364 , \10363 , \6144 );
not \U$10112 ( \10365 , \10363 );
and \U$10113 ( \10366 , \10365 , \6624 );
nor \U$10114 ( \10367 , \10364 , \10366 );
not \U$10115 ( \10368 , \10367 );
not \U$10116 ( \10369 , \10368 );
and \U$10117 ( \10370 , \10358 , \10369 );
and \U$10118 ( \10371 , \10357 , \10368 );
nor \U$10119 ( \10372 , \10370 , \10371 );
not \U$10120 ( \10373 , RIbe29650_59);
not \U$10121 ( \10374 , \4021 );
or \U$10122 ( \10375 , \10373 , \10374 );
nand \U$10123 ( \10376 , \4027 , RIbe29038_46);
nand \U$10124 ( \10377 , \10375 , \10376 );
and \U$10125 ( \10378 , \10377 , \3471 );
not \U$10126 ( \10379 , \10377 );
and \U$10127 ( \10380 , \10379 , \3448 );
nor \U$10128 ( \10381 , \10378 , \10380 );
not \U$10129 ( \10382 , RIbe29830_63);
not \U$10130 ( \10383 , \3452 );
or \U$10131 ( \10384 , \10382 , \10383 );
nand \U$10132 ( \10385 , \3458 , RIbe296c8_60);
nand \U$10133 ( \10386 , \10384 , \10385 );
and \U$10134 ( \10387 , \10386 , \2887 );
not \U$10135 ( \10388 , \10386 );
and \U$10136 ( \10389 , \10388 , \3290 );
nor \U$10137 ( \10390 , \10387 , \10389 );
and \U$10138 ( \10391 , \10381 , \10390 );
not \U$10139 ( \10392 , \10381 );
not \U$10140 ( \10393 , \10390 );
and \U$10141 ( \10394 , \10392 , \10393 );
or \U$10142 ( \10395 , \10391 , \10394 );
not \U$10143 ( \10396 , \2379 );
not \U$10144 ( \10397 , RIbe281b0_15);
not \U$10145 ( \10398 , \2898 );
or \U$10146 ( \10399 , \10397 , \10398 );
nand \U$10147 ( \10400 , \4284 , RIbe280c0_13);
nand \U$10148 ( \10401 , \10399 , \10400 );
not \U$10149 ( \10402 , \10401 );
or \U$10150 ( \10403 , \10396 , \10402 );
or \U$10151 ( \10404 , \10401 , \2379 );
nand \U$10152 ( \10405 , \10403 , \10404 );
xor \U$10153 ( \10406 , \10395 , \10405 );
xor \U$10154 ( \10407 , \10372 , \10406 );
not \U$10155 ( \10408 , RIbe28b10_35);
not \U$10156 ( \10409 , \1143 );
or \U$10157 ( \10410 , \10408 , \10409 );
nand \U$10158 ( \10411 , \1147 , RIbe28b88_36);
nand \U$10159 ( \10412 , \10410 , \10411 );
and \U$10160 ( \10413 , \10412 , \1652 );
not \U$10161 ( \10414 , \10412 );
and \U$10162 ( \10415 , \10414 , \3994 );
nor \U$10163 ( \10416 , \10413 , \10415 );
not \U$10164 ( \10417 , \6345 );
not \U$10165 ( \10418 , \10025 );
and \U$10166 ( \10419 , \10417 , \10418 );
and \U$10167 ( \10420 , \1744 , RIbe287c8_28);
nor \U$10168 ( \10421 , \10419 , \10420 );
and \U$10169 ( \10422 , \10421 , \1618 );
not \U$10170 ( \10423 , \10421 );
and \U$10171 ( \10424 , \10423 , \3959 );
nor \U$10172 ( \10425 , \10422 , \10424 );
xor \U$10173 ( \10426 , \10416 , \10425 );
and \U$10174 ( \10427 , \1807 , RIbe28408_20);
and \U$10175 ( \10428 , \1165 , RIbe28390_19);
nor \U$10176 ( \10429 , \10427 , \10428 );
and \U$10177 ( \10430 , \10429 , \1608 );
not \U$10178 ( \10431 , \10429 );
and \U$10179 ( \10432 , \10431 , \1011 );
nor \U$10180 ( \10433 , \10430 , \10432 );
xor \U$10181 ( \10434 , \10426 , \10433 );
not \U$10182 ( \10435 , \4065 );
not \U$10183 ( \10436 , \3952 );
and \U$10184 ( \10437 , \10435 , \10436 );
and \U$10185 ( \10438 , \3303 , RIbe29560_57);
nor \U$10186 ( \10439 , \10437 , \10438 );
and \U$10187 ( \10440 , \10439 , \1277 );
not \U$10188 ( \10441 , \10439 );
and \U$10189 ( \10442 , \10441 , \3516 );
nor \U$10190 ( \10443 , \10440 , \10442 );
not \U$10191 ( \10444 , \10443 );
not \U$10192 ( \10445 , \10444 );
and \U$10193 ( \10446 , \6380 , RIbe289a8_32);
and \U$10194 ( \10447 , \5467 , RIbe28930_31);
nor \U$10195 ( \10448 , \10446 , \10447 );
and \U$10196 ( \10449 , \10448 , \3491 );
not \U$10197 ( \10450 , \10448 );
and \U$10198 ( \10451 , \10450 , \1131 );
or \U$10199 ( \10452 , \10449 , \10451 );
not \U$10200 ( \10453 , \10452 );
or \U$10201 ( \10454 , \10445 , \10453 );
not \U$10202 ( \10455 , \10452 );
nand \U$10203 ( \10456 , \10455 , \10443 );
nand \U$10204 ( \10457 , \10454 , \10456 );
not \U$10205 ( \10458 , RIbe29290_51);
not \U$10206 ( \10459 , \1633 );
or \U$10207 ( \10460 , \10458 , \10459 );
nand \U$10208 ( \10461 , \2817 , RIbe28a20_33);
nand \U$10209 ( \10462 , \10460 , \10461 );
and \U$10210 ( \10463 , \10462 , \5125 );
not \U$10211 ( \10464 , \10462 );
and \U$10212 ( \10465 , \10464 , \1309 );
nor \U$10213 ( \10466 , \10463 , \10465 );
not \U$10214 ( \10467 , \10466 );
not \U$10215 ( \10468 , \10467 );
and \U$10216 ( \10469 , \10457 , \10468 );
not \U$10217 ( \10470 , \10457 );
and \U$10218 ( \10471 , \10470 , \10467 );
nor \U$10219 ( \10472 , \10469 , \10471 );
and \U$10220 ( \10473 , \10434 , \10472 );
not \U$10221 ( \10474 , \10434 );
not \U$10222 ( \10475 , \10472 );
and \U$10223 ( \10476 , \10474 , \10475 );
or \U$10224 ( \10477 , \10473 , \10476 );
xnor \U$10225 ( \10478 , \10407 , \10477 );
nand \U$10226 ( \10479 , \9423 , \9416 );
nand \U$10227 ( \10480 , \10479 , \9432 );
or \U$10228 ( \10481 , \9416 , \9423 );
nand \U$10229 ( \10482 , \10480 , \10481 );
and \U$10230 ( \10483 , RIbe29380_53, RIbe29e48_76);
and \U$10231 ( \10484 , \324 , RIbe29dd0_75);
and \U$10232 ( \10485 , \329 , RIbe29c68_72);
nor \U$10233 ( \10486 , \10484 , \10485 );
and \U$10234 ( \10487 , \10486 , \1374 );
not \U$10235 ( \10488 , \10486 );
and \U$10236 ( \10489 , \10488 , \338 );
nor \U$10237 ( \10490 , \10487 , \10489 );
xor \U$10238 ( \10491 , \10483 , \10490 );
and \U$10239 ( \10492 , \260 , RIbe29bf0_71);
and \U$10240 ( \10493 , \1831 , RIbe28f48_44);
nor \U$10241 ( \10494 , \10492 , \10493 );
and \U$10242 ( \10495 , \10494 , \1362 );
not \U$10243 ( \10496 , \10494 );
and \U$10244 ( \10497 , \10496 , \1363 );
nor \U$10245 ( \10498 , \10495 , \10497 );
xor \U$10246 ( \10499 , \10491 , \10498 );
xor \U$10247 ( \10500 , \10482 , \10499 );
not \U$10248 ( \10501 , RIbe28660_25);
not \U$10249 ( \10502 , \548 );
or \U$10250 ( \10503 , \10501 , \10502 );
nand \U$10251 ( \10504 , \552 , RIbe285e8_24);
nand \U$10252 ( \10505 , \10503 , \10504 );
and \U$10253 ( \10506 , \10505 , \1330 );
not \U$10254 ( \10507 , \10505 );
and \U$10255 ( \10508 , \10507 , \424 );
nor \U$10256 ( \10509 , \10506 , \10508 );
not \U$10257 ( \10510 , RIbe27f58_10);
not \U$10258 ( \10511 , \1774 );
or \U$10259 ( \10512 , \10510 , \10511 );
nand \U$10260 ( \10513 , \429 , RIbe27e68_8);
nand \U$10261 ( \10514 , \10512 , \10513 );
and \U$10262 ( \10515 , \10514 , \306 );
not \U$10263 ( \10516 , \10514 );
and \U$10264 ( \10517 , \10516 , \3175 );
nor \U$10265 ( \10518 , \10515 , \10517 );
xor \U$10266 ( \10519 , \10509 , \10518 );
and \U$10267 ( \10520 , \1254 , RIbe28ed0_43);
and \U$10268 ( \10521 , \1531 , RIbe27fd0_11);
nor \U$10269 ( \10522 , \10520 , \10521 );
and \U$10270 ( \10523 , \10522 , \300 );
not \U$10271 ( \10524 , \10522 );
and \U$10272 ( \10525 , \10524 , \293 );
nor \U$10273 ( \10526 , \10523 , \10525 );
xor \U$10274 ( \10527 , \10519 , \10526 );
xnor \U$10275 ( \10528 , \10500 , \10527 );
not \U$10276 ( \10529 , \10528 );
and \U$10277 ( \10530 , \10478 , \10529 );
not \U$10278 ( \10531 , \10478 );
and \U$10279 ( \10532 , \10531 , \10528 );
nor \U$10280 ( \10533 , \10530 , \10532 );
not \U$10281 ( \10534 , \10533 );
xor \U$10282 ( \10535 , \9598 , \9607 );
and \U$10283 ( \10536 , \10535 , \9617 );
and \U$10284 ( \10537 , \9598 , \9607 );
or \U$10285 ( \10538 , \10536 , \10537 );
and \U$10286 ( \10539 , \9690 , \9678 );
nor \U$10287 ( \10540 , \10539 , \9666 );
nor \U$10288 ( \10541 , \9690 , \9678 );
nor \U$10289 ( \10542 , \10540 , \10541 );
xor \U$10290 ( \10543 , \10538 , \10542 );
nand \U$10291 ( \10544 , \9628 , \9654 );
and \U$10292 ( \10545 , \10544 , \9640 );
nor \U$10293 ( \10546 , \9654 , \9628 );
nor \U$10294 ( \10547 , \10545 , \10546 );
xnor \U$10295 ( \10548 , \10543 , \10547 );
not \U$10296 ( \10549 , \10548 );
not \U$10297 ( \10550 , \9530 );
not \U$10298 ( \10551 , \9508 );
or \U$10299 ( \10552 , \10550 , \10551 );
nand \U$10300 ( \10553 , \10552 , \9519 );
not \U$10301 ( \10554 , \9508 );
nand \U$10302 ( \10555 , \10554 , \9529 );
nand \U$10303 ( \10556 , \10553 , \10555 );
not \U$10304 ( \10557 , \9487 );
not \U$10305 ( \10558 , \9497 );
or \U$10306 ( \10559 , \10557 , \10558 );
nand \U$10307 ( \10560 , \9496 , \9484 );
nand \U$10308 ( \10561 , \10560 , \9474 );
nand \U$10309 ( \10562 , \10559 , \10561 );
not \U$10310 ( \10563 , \10562 );
and \U$10311 ( \10564 , \9566 , \9546 );
nor \U$10312 ( \10565 , \10564 , \9556 );
nor \U$10313 ( \10566 , \9546 , \9566 );
nor \U$10314 ( \10567 , \10565 , \10566 );
not \U$10315 ( \10568 , \10567 );
or \U$10316 ( \10569 , \10563 , \10568 );
or \U$10317 ( \10570 , \10567 , \10562 );
nand \U$10318 ( \10571 , \10569 , \10570 );
xor \U$10319 ( \10572 , \10556 , \10571 );
not \U$10320 ( \10573 , \10572 );
and \U$10321 ( \10574 , \10549 , \10573 );
and \U$10322 ( \10575 , \10572 , \10548 );
nor \U$10323 ( \10576 , \10574 , \10575 );
not \U$10324 ( \10577 , \10576 );
and \U$10325 ( \10578 , \10534 , \10577 );
and \U$10326 ( \10579 , \10533 , \10576 );
nor \U$10327 ( \10580 , \10578 , \10579 );
xnor \U$10328 ( \10581 , \10344 , \10580 );
xor \U$10329 ( \10582 , \10306 , \10581 );
xor \U$10330 ( \10583 , \10234 , \10582 );
xor \U$10331 ( \10584 , \10224 , \10583 );
xnor \U$10332 ( \10585 , \10216 , \10584 );
not \U$10333 ( \10586 , \10194 );
not \U$10334 ( \10587 , \10201 );
or \U$10335 ( \10588 , \10586 , \10587 );
or \U$10336 ( \10589 , \10201 , \10194 );
nand \U$10337 ( \10590 , \10588 , \10589 );
xor \U$10338 ( \10591 , \9738 , \10181 );
xor \U$10339 ( \10592 , \10591 , \10191 );
xor \U$10340 ( \10593 , \8050 , \8435 );
xor \U$10341 ( \10594 , \10593 , \8514 );
not \U$10342 ( \10595 , \10144 );
not \U$10343 ( \10596 , \10130 );
or \U$10344 ( \10597 , \10595 , \10596 );
or \U$10345 ( \10598 , \10144 , \10130 );
nand \U$10346 ( \10599 , \10597 , \10598 );
not \U$10347 ( \10600 , \10134 );
and \U$10348 ( \10601 , \10599 , \10600 );
not \U$10349 ( \10602 , \10599 );
and \U$10350 ( \10603 , \10602 , \10134 );
nor \U$10351 ( \10604 , \10601 , \10603 );
xor \U$10352 ( \10605 , \9780 , \9811 );
xor \U$10353 ( \10606 , \10605 , \9847 );
xor \U$10354 ( \10607 , \9998 , \10035 );
xor \U$10355 ( \10608 , \10607 , \10067 );
xor \U$10356 ( \10609 , \10606 , \10608 );
and \U$10357 ( \10610 , \9923 , \9886 );
not \U$10358 ( \10611 , \9923 );
and \U$10359 ( \10612 , \10611 , \9962 );
nor \U$10360 ( \10613 , \10610 , \10612 );
xor \U$10361 ( \10614 , \10613 , \9959 );
and \U$10362 ( \10615 , \10609 , \10614 );
and \U$10363 ( \10616 , \10606 , \10608 );
or \U$10364 ( \10617 , \10615 , \10616 );
not \U$10365 ( \10618 , \10617 );
nand \U$10366 ( \10619 , \10604 , \10618 );
xor \U$10367 ( \10620 , \9753 , \9749 );
xor \U$10368 ( \10621 , \10620 , \9740 );
not \U$10369 ( \10622 , \10621 );
and \U$10370 ( \10623 , \10619 , \10622 );
nor \U$10371 ( \10624 , \10604 , \10618 );
nor \U$10372 ( \10625 , \10623 , \10624 );
not \U$10373 ( \10626 , \9823 );
not \U$10374 ( \10627 , \9842 );
or \U$10375 ( \10628 , \10626 , \10627 );
or \U$10376 ( \10629 , \9842 , \9823 );
nand \U$10377 ( \10630 , \10628 , \10629 );
and \U$10378 ( \10631 , \10630 , \9831 );
not \U$10379 ( \10632 , \10630 );
and \U$10380 ( \10633 , \10632 , \9845 );
nor \U$10381 ( \10634 , \10631 , \10633 );
not \U$10382 ( \10635 , \10634 );
not \U$10383 ( \10636 , \10635 );
xor \U$10384 ( \10637 , \9779 , \1378 );
xnor \U$10385 ( \10638 , \10637 , \9775 );
not \U$10386 ( \10639 , \10638 );
not \U$10387 ( \10640 , \10639 );
or \U$10388 ( \10641 , \10636 , \10640 );
not \U$10389 ( \10642 , \10634 );
not \U$10390 ( \10643 , \10638 );
or \U$10391 ( \10644 , \10642 , \10643 );
xor \U$10392 ( \10645 , \9786 , \9809 );
and \U$10393 ( \10646 , \10645 , \9794 );
not \U$10394 ( \10647 , \10645 );
and \U$10395 ( \10648 , \10647 , \9795 );
nor \U$10396 ( \10649 , \10646 , \10648 );
nand \U$10397 ( \10650 , \10644 , \10649 );
nand \U$10398 ( \10651 , \10641 , \10650 );
not \U$10399 ( \10652 , \10651 );
not \U$10400 ( \10653 , \10652 );
xor \U$10401 ( \10654 , \9983 , \9994 );
xor \U$10402 ( \10655 , \10654 , \9974 );
not \U$10403 ( \10656 , \10655 );
xor \U$10404 ( \10657 , \10019 , \10007 );
xor \U$10405 ( \10658 , \10657 , \10033 );
not \U$10406 ( \10659 , \10658 );
or \U$10407 ( \10660 , \10656 , \10659 );
xor \U$10408 ( \10661 , \10045 , \10054 );
xor \U$10409 ( \10662 , \10661 , \10064 );
nand \U$10410 ( \10663 , \10660 , \10662 );
not \U$10411 ( \10664 , \10658 );
not \U$10412 ( \10665 , \10655 );
nand \U$10413 ( \10666 , \10664 , \10665 );
nand \U$10414 ( \10667 , \10663 , \10666 );
not \U$10415 ( \10668 , \10667 );
not \U$10416 ( \10669 , \10668 );
or \U$10417 ( \10670 , \10653 , \10669 );
xor \U$10418 ( \10671 , \9935 , \9946 );
xor \U$10419 ( \10672 , \10671 , \9956 );
not \U$10420 ( \10673 , \10672 );
xor \U$10421 ( \10674 , \7969 , \9902 );
xor \U$10422 ( \10675 , \10674 , \9916 );
xnor \U$10423 ( \10676 , \10675 , \9898 );
buf \U$10424 ( \10677 , \10676 );
not \U$10425 ( \10678 , \10677 );
or \U$10426 ( \10679 , \10673 , \10678 );
or \U$10427 ( \10680 , \10677 , \10672 );
not \U$10428 ( \10681 , \9859 );
not \U$10429 ( \10682 , \9883 );
or \U$10430 ( \10683 , \10681 , \10682 );
not \U$10431 ( \10684 , \9859 );
nand \U$10432 ( \10685 , \10684 , \9882 );
nand \U$10433 ( \10686 , \10683 , \10685 );
xnor \U$10434 ( \10687 , \10686 , \9870 );
nand \U$10435 ( \10688 , \10680 , \10687 );
nand \U$10436 ( \10689 , \10679 , \10688 );
nand \U$10437 ( \10690 , \10670 , \10689 );
nand \U$10438 ( \10691 , \10667 , \10651 );
nand \U$10439 ( \10692 , \10690 , \10691 );
not \U$10440 ( \10693 , \10692 );
and \U$10441 ( \10694 , \325 , RIbe2a550_91);
and \U$10442 ( \10695 , \330 , RIbe2a988_100);
nor \U$10443 ( \10696 , \10694 , \10695 );
and \U$10444 ( \10697 , \10696 , \1375 );
not \U$10445 ( \10698 , \10696 );
and \U$10446 ( \10699 , \10698 , \1379 );
nor \U$10447 ( \10700 , \10697 , \10699 );
nand \U$10448 ( \10701 , RIbe29380_53, RIbe2a5c8_92);
nand \U$10449 ( \10702 , \10700 , \10701 );
and \U$10450 ( \10703 , \6311 , RIbe2a3e8_88);
and \U$10451 ( \10704 , \9816 , RIbe2a370_87);
nor \U$10452 ( \10705 , \10703 , \10704 );
and \U$10453 ( \10706 , \10705 , \300 );
not \U$10454 ( \10707 , \10705 );
and \U$10455 ( \10708 , \10707 , \293 );
nor \U$10456 ( \10709 , \10706 , \10708 );
not \U$10457 ( \10710 , RIbe2a2f8_86);
not \U$10458 ( \10711 , \1773 );
or \U$10459 ( \10712 , \10710 , \10711 );
nand \U$10460 ( \10713 , \429 , RIbe2acd0_107);
nand \U$10461 ( \10714 , \10712 , \10713 );
and \U$10462 ( \10715 , \10714 , \306 );
not \U$10463 ( \10716 , \10714 );
and \U$10464 ( \10717 , \10716 , \313 );
nor \U$10465 ( \10718 , \10715 , \10717 );
xor \U$10466 ( \10719 , \10709 , \10718 );
and \U$10467 ( \10720 , \261 , RIbe2a910_99);
and \U$10468 ( \10721 , \263 , RIbe2b5b8_126);
nor \U$10469 ( \10722 , \10720 , \10721 );
and \U$10470 ( \10723 , \10722 , \270 );
not \U$10471 ( \10724 , \10722 );
and \U$10472 ( \10725 , \10724 , \1363 );
nor \U$10473 ( \10726 , \10723 , \10725 );
and \U$10474 ( \10727 , \10719 , \10726 );
and \U$10475 ( \10728 , \10709 , \10718 );
or \U$10476 ( \10729 , \10727 , \10728 );
xor \U$10477 ( \10730 , \10702 , \10729 );
not \U$10478 ( \10731 , RIbe2a028_80);
not \U$10479 ( \10732 , \1756 );
or \U$10480 ( \10733 , \10731 , \10732 );
nand \U$10481 ( \10734 , \1327 , RIbe29fb0_79);
nand \U$10482 ( \10735 , \10733 , \10734 );
xnor \U$10483 ( \10736 , \10735 , \424 );
and \U$10484 ( \10737 , \1807 , RIbe29c68_72);
and \U$10485 ( \10738 , \1203 , RIbe29bf0_71);
nor \U$10486 ( \10739 , \10737 , \10738 );
and \U$10487 ( \10740 , \10739 , \1813 );
not \U$10488 ( \10741 , \10739 );
and \U$10489 ( \10742 , \10741 , \1011 );
nor \U$10490 ( \10743 , \10740 , \10742 );
or \U$10491 ( \10744 , \10736 , \10743 );
not \U$10492 ( \10745 , RIbe29e48_76);
not \U$10493 ( \10746 , \1744 );
or \U$10494 ( \10747 , \10745 , \10746 );
nand \U$10495 ( \10748 , \1180 , RIbe29dd0_75);
nand \U$10496 ( \10749 , \10747 , \10748 );
xor \U$10497 ( \10750 , \10749 , \564 );
not \U$10498 ( \10751 , \10750 );
nand \U$10499 ( \10752 , \10744 , \10751 );
nand \U$10500 ( \10753 , \10736 , \10743 );
nand \U$10501 ( \10754 , \10752 , \10753 );
and \U$10502 ( \10755 , \10730 , \10754 );
and \U$10503 ( \10756 , \10702 , \10729 );
or \U$10504 ( \10757 , \10755 , \10756 );
not \U$10505 ( \10758 , \10757 );
not \U$10506 ( \10759 , \1284 );
and \U$10507 ( \10760 , \10759 , RIbe27e68_8);
not \U$10508 ( \10761 , \6382 );
and \U$10509 ( \10762 , \10761 , RIbe28660_25);
nor \U$10510 ( \10763 , \10760 , \10762 );
and \U$10511 ( \10764 , \10763 , \2563 );
not \U$10512 ( \10765 , \10763 );
and \U$10513 ( \10766 , \10765 , \1131 );
nor \U$10514 ( \10767 , \10764 , \10766 );
not \U$10515 ( \10768 , \10767 );
not \U$10516 ( \10769 , RIbe28f48_44);
not \U$10517 ( \10770 , \1143 );
or \U$10518 ( \10771 , \10769 , \10770 );
nand \U$10519 ( \10772 , \1147 , RIbe28ed0_43);
nand \U$10520 ( \10773 , \10771 , \10772 );
and \U$10521 ( \10774 , \10773 , \1153 );
not \U$10522 ( \10775 , \10773 );
and \U$10523 ( \10776 , \10775 , \1469 );
nor \U$10524 ( \10777 , \10774 , \10776 );
nand \U$10525 ( \10778 , \10768 , \10777 );
not \U$10526 ( \10779 , RIbe27fd0_11);
not \U$10527 ( \10780 , \8868 );
or \U$10528 ( \10781 , \10779 , \10780 );
nand \U$10529 ( \10782 , \2817 , RIbe27f58_10);
nand \U$10530 ( \10783 , \10781 , \10782 );
and \U$10531 ( \10784 , \10783 , \1082 );
not \U$10532 ( \10785 , \10783 );
and \U$10533 ( \10786 , \10785 , \1309 );
nor \U$10534 ( \10787 , \10784 , \10786 );
not \U$10535 ( \10788 , \10787 );
and \U$10536 ( \10789 , \10778 , \10788 );
nor \U$10537 ( \10790 , \10768 , \10777 );
nor \U$10538 ( \10791 , \10789 , \10790 );
not \U$10539 ( \10792 , \10791 );
not \U$10540 ( \10793 , RIbe28b88_36);
not \U$10541 ( \10794 , \5094 );
or \U$10542 ( \10795 , \10793 , \10794 );
nand \U$10543 ( \10796 , \7438 , RIbe29290_51);
nand \U$10544 ( \10797 , \10795 , \10796 );
and \U$10545 ( \10798 , \10797 , \4821 );
not \U$10546 ( \10799 , \10797 );
and \U$10547 ( \10800 , \10799 , \3471 );
nor \U$10548 ( \10801 , \10798 , \10800 );
not \U$10549 ( \10802 , RIbe28a20_33);
not \U$10550 ( \10803 , \6414 );
or \U$10551 ( \10804 , \10802 , \10803 );
nand \U$10552 ( \10805 , \4600 , RIbe289a8_32);
nand \U$10553 ( \10806 , \10804 , \10805 );
and \U$10554 ( \10807 , \10806 , \4323 );
not \U$10555 ( \10808 , \10806 );
and \U$10556 ( \10809 , \10808 , \4326 );
nor \U$10557 ( \10810 , \10807 , \10809 );
nand \U$10558 ( \10811 , \10801 , \10810 );
not \U$10559 ( \10812 , RIbe28930_31);
not \U$10560 ( \10813 , \6427 );
or \U$10561 ( \10814 , \10812 , \10813 );
nand \U$10562 ( \10815 , \7056 , RIbe29560_57);
nand \U$10563 ( \10816 , \10814 , \10815 );
and \U$10564 ( \10817 , \10816 , \4586 );
not \U$10565 ( \10818 , \10816 );
and \U$10566 ( \10819 , \10818 , \4592 );
nor \U$10567 ( \10820 , \10817 , \10819 );
and \U$10568 ( \10821 , \10811 , \10820 );
nor \U$10569 ( \10822 , \10801 , \10810 );
nor \U$10570 ( \10823 , \10821 , \10822 );
not \U$10571 ( \10824 , \10823 );
or \U$10572 ( \10825 , \10792 , \10824 );
not \U$10573 ( \10826 , RIbe28480_21);
not \U$10574 ( \10827 , \7827 );
or \U$10575 ( \10828 , \10826 , \10827 );
nand \U$10576 ( \10829 , \3267 , RIbe28408_20);
nand \U$10577 ( \10830 , \10828 , \10829 );
not \U$10578 ( \10831 , \10830 );
not \U$10579 ( \10832 , \2379 );
and \U$10580 ( \10833 , \10831 , \10832 );
and \U$10581 ( \10834 , \10830 , \2379 );
nor \U$10582 ( \10835 , \10833 , \10834 );
not \U$10583 ( \10836 , \10835 );
not \U$10584 ( \10837 , \10836 );
not \U$10585 ( \10838 , RIbe28390_19);
not \U$10586 ( \10839 , \3284 );
or \U$10587 ( \10840 , \10838 , \10839 );
nand \U$10588 ( \10841 , \4011 , RIbe28b10_35);
nand \U$10589 ( \10842 , \10840 , \10841 );
and \U$10590 ( \10843 , \10842 , \4346 );
not \U$10591 ( \10844 , \10842 );
and \U$10592 ( \10845 , \10844 , \3461 );
nor \U$10593 ( \10846 , \10843 , \10845 );
not \U$10594 ( \10847 , \10846 );
or \U$10595 ( \10848 , \10837 , \10847 );
not \U$10596 ( \10849 , \10835 );
not \U$10597 ( \10850 , \10846 );
not \U$10598 ( \10851 , \10850 );
or \U$10599 ( \10852 , \10849 , \10851 );
not \U$10600 ( \10853 , \4065 );
not \U$10601 ( \10854 , RIbe287c8_28);
not \U$10602 ( \10855 , \10854 );
and \U$10603 ( \10856 , \10853 , \10855 );
and \U$10604 ( \10857 , \1272 , RIbe285e8_24);
nor \U$10605 ( \10858 , \10856 , \10857 );
and \U$10606 ( \10859 , \10858 , \3516 );
not \U$10607 ( \10860 , \10858 );
and \U$10608 ( \10861 , \10860 , \1277 );
nor \U$10609 ( \10862 , \10859 , \10861 );
nand \U$10610 ( \10863 , \10852 , \10862 );
nand \U$10611 ( \10864 , \10848 , \10863 );
nand \U$10612 ( \10865 , \10825 , \10864 );
not \U$10613 ( \10866 , \10823 );
not \U$10614 ( \10867 , \10791 );
nand \U$10615 ( \10868 , \10866 , \10867 );
nand \U$10616 ( \10869 , \10865 , \10868 );
not \U$10617 ( \10870 , \10869 );
or \U$10618 ( \10871 , \10758 , \10870 );
or \U$10619 ( \10872 , \10869 , \10757 );
not \U$10620 ( \10873 , RIbe290b0_47);
not \U$10621 ( \10874 , \7954 );
or \U$10622 ( \10875 , \10873 , \10874 );
nand \U$10623 ( \10876 , \7958 , RIbe29a88_68);
nand \U$10624 ( \10877 , \10875 , \10876 );
and \U$10625 ( \10878 , \10877 , \7293 );
not \U$10626 ( \10879 , \10877 );
and \U$10627 ( \10880 , \10879 , \6572 );
nor \U$10628 ( \10881 , \10878 , \10880 );
not \U$10629 ( \10882 , \10881 );
not \U$10630 ( \10883 , RIbe29038_46);
not \U$10631 ( \10884 , \6592 );
or \U$10632 ( \10885 , \10883 , \10884 );
nand \U$10633 ( \10886 , \7483 , RIbe28fc0_45);
nand \U$10634 ( \10887 , \10885 , \10886 );
not \U$10635 ( \10888 , \7948 );
and \U$10636 ( \10889 , \10887 , \10888 );
not \U$10637 ( \10890 , \10887 );
and \U$10638 ( \10891 , \10890 , \7948 );
nor \U$10639 ( \10892 , \10889 , \10891 );
nand \U$10640 ( \10893 , \10882 , \10892 );
not \U$10641 ( \10894 , RIbe27d78_6);
not \U$10642 ( \10895 , \7298 );
or \U$10643 ( \10896 , \10894 , \10895 );
not \U$10644 ( \10897 , \6983 );
not \U$10645 ( \10898 , \10897 );
nand \U$10646 ( \10899 , \10898 , RIbe27d00_5);
nand \U$10647 ( \10900 , \10896 , \10899 );
not \U$10648 ( \10901 , \10900 );
buf \U$10649 ( \10902 , \6992 );
not \U$10650 ( \10903 , \10902 );
and \U$10651 ( \10904 , \10901 , \10903 );
and \U$10652 ( \10905 , \10900 , \7661 );
nor \U$10653 ( \10906 , \10904 , \10905 );
not \U$10654 ( \10907 , \10906 );
and \U$10655 ( \10908 , \10893 , \10907 );
nor \U$10656 ( \10909 , \10882 , \10892 );
nor \U$10657 ( \10910 , \10908 , \10909 );
not \U$10658 ( \10911 , \10910 );
not \U$10659 ( \10912 , \7970 );
not \U$10660 ( \10913 , \10912 );
not \U$10661 ( \10914 , RIbe28de0_41);
buf \U$10662 ( \10915 , \8276 );
buf \U$10663 ( \10916 , \10915 );
not \U$10664 ( \10917 , \10916 );
or \U$10665 ( \10918 , \10914 , \10917 );
buf \U$10666 ( \10919 , \9912 );
not \U$10667 ( \10920 , \10919 );
not \U$10668 ( \10921 , \10920 );
nand \U$10669 ( \10922 , \10921 , RIbe29920_65);
nand \U$10670 ( \10923 , \10918 , \10922 );
not \U$10671 ( \10924 , \10923 );
or \U$10672 ( \10925 , \10913 , \10924 );
not \U$10673 ( \10926 , \8077 );
not \U$10674 ( \10927 , \10926 );
or \U$10675 ( \10928 , \10927 , \10923 );
nand \U$10676 ( \10929 , \10925 , \10928 );
nand \U$10677 ( \10930 , RIbe2a4d8_90, RIbe2a460_89);
nor \U$10678 ( \10931 , RIbe2a4d8_90, RIbe2adc0_109);
not \U$10679 ( \10932 , \10931 );
not \U$10680 ( \10933 , RIbe2a460_89);
nand \U$10681 ( \10934 , \10933 , RIbe2adc0_109);
and \U$10682 ( \10935 , \10930 , \10932 , \10934 );
buf \U$10683 ( \10936 , \10935 );
not \U$10684 ( \10937 , \10936 );
not \U$10685 ( \10938 , \10937 );
nand \U$10686 ( \10939 , \10938 , RIbe27b98_2);
not \U$10687 ( \10940 , \9902 );
and \U$10688 ( \10941 , \10939 , \10940 );
not \U$10689 ( \10942 , \10939 );
not \U$10690 ( \10943 , \9901 );
not \U$10691 ( \10944 , \10943 );
and \U$10692 ( \10945 , \10942 , \10944 );
nor \U$10693 ( \10946 , \10941 , \10945 );
or \U$10694 ( \10947 , \10929 , \10946 );
not \U$10695 ( \10948 , RIbe27c10_3);
buf \U$10696 ( \10949 , \7974 );
not \U$10697 ( \10950 , \10949 );
or \U$10698 ( \10951 , \10948 , \10950 );
not \U$10699 ( \10952 , \7980 );
nand \U$10700 ( \10953 , \10952 , RIbe28e58_42);
nand \U$10701 ( \10954 , \10951 , \10953 );
and \U$10702 ( \10955 , \10954 , \7988 );
not \U$10703 ( \10956 , \10954 );
and \U$10704 ( \10957 , \10956 , \7989 );
nor \U$10705 ( \10958 , \10955 , \10957 );
and \U$10706 ( \10959 , \10947 , \10958 );
and \U$10707 ( \10960 , \10946 , \10929 );
nor \U$10708 ( \10961 , \10959 , \10960 );
not \U$10709 ( \10962 , \10961 );
or \U$10710 ( \10963 , \10911 , \10962 );
not \U$10711 ( \10964 , RIbe280c0_13);
not \U$10712 ( \10965 , \6139 );
or \U$10713 ( \10966 , \10964 , \10965 );
nand \U$10714 ( \10967 , \7528 , RIbe29830_63);
nand \U$10715 ( \10968 , \10966 , \10967 );
not \U$10716 ( \10969 , \6141 );
and \U$10717 ( \10970 , \10968 , \10969 );
not \U$10718 ( \10971 , \10968 );
not \U$10719 ( \10972 , \5741 );
and \U$10720 ( \10973 , \10971 , \10972 );
nor \U$10721 ( \10974 , \10970 , \10973 );
not \U$10722 ( \10975 , \10974 );
not \U$10723 ( \10976 , \5754 );
not \U$10724 ( \10977 , RIbe28228_16);
not \U$10725 ( \10978 , \5455 );
or \U$10726 ( \10979 , \10977 , \10978 );
nand \U$10727 ( \10980 , \10269 , RIbe281b0_15);
nand \U$10728 ( \10981 , \10979 , \10980 );
not \U$10729 ( \10982 , \10981 );
or \U$10730 ( \10983 , \10976 , \10982 );
not \U$10731 ( \10984 , \6121 );
or \U$10732 ( \10985 , \10981 , \10984 );
nand \U$10733 ( \10986 , \10983 , \10985 );
not \U$10734 ( \10987 , \10986 );
or \U$10735 ( \10988 , \10975 , \10987 );
or \U$10736 ( \10989 , \10986 , \10974 );
not \U$10737 ( \10990 , RIbe296c8_60);
not \U$10738 ( \10991 , \6537 );
or \U$10739 ( \10992 , \10990 , \10991 );
nand \U$10740 ( \10993 , \6540 , RIbe29650_59);
nand \U$10741 ( \10994 , \10992 , \10993 );
and \U$10742 ( \10995 , \10994 , \6546 );
not \U$10743 ( \10996 , \10994 );
and \U$10744 ( \10997 , \10996 , \6551 );
nor \U$10745 ( \10998 , \10995 , \10997 );
nand \U$10746 ( \10999 , \10989 , \10998 );
nand \U$10747 ( \11000 , \10988 , \10999 );
nand \U$10748 ( \11001 , \10963 , \11000 );
not \U$10749 ( \11002 , \10961 );
not \U$10750 ( \11003 , \10910 );
nand \U$10751 ( \11004 , \11002 , \11003 );
nand \U$10752 ( \11005 , \11001 , \11004 );
nand \U$10753 ( \11006 , \10872 , \11005 );
nand \U$10754 ( \11007 , \10871 , \11006 );
not \U$10755 ( \11008 , \11007 );
nand \U$10756 ( \11009 , \10693 , \11008 );
not \U$10757 ( \11010 , \11009 );
not \U$10758 ( \11011 , \10075 );
not \U$10759 ( \11012 , \11011 );
xor \U$10760 ( \11013 , \8114 , \8167 );
xnor \U$10761 ( \11014 , \11013 , \10083 );
not \U$10762 ( \11015 , \11014 );
or \U$10763 ( \11016 , \11012 , \11015 );
or \U$10764 ( \11017 , \11014 , \11011 );
nand \U$10765 ( \11018 , \11016 , \11017 );
not \U$10766 ( \11019 , \10114 );
not \U$10767 ( \11020 , \11019 );
not \U$10768 ( \11021 , \10117 );
not \U$10769 ( \11022 , \10111 );
or \U$10770 ( \11023 , \11021 , \11022 );
or \U$10771 ( \11024 , \10111 , \10117 );
nand \U$10772 ( \11025 , \11023 , \11024 );
not \U$10773 ( \11026 , \11025 );
or \U$10774 ( \11027 , \11020 , \11026 );
or \U$10775 ( \11028 , \11025 , \11019 );
nand \U$10776 ( \11029 , \11027 , \11028 );
xor \U$10777 ( \11030 , \11018 , \11029 );
not \U$10778 ( \11031 , \10097 );
not \U$10779 ( \11032 , \10100 );
not \U$10780 ( \11033 , \10095 );
or \U$10781 ( \11034 , \11032 , \11033 );
or \U$10782 ( \11035 , \10095 , \10100 );
nand \U$10783 ( \11036 , \11034 , \11035 );
not \U$10784 ( \11037 , \11036 );
or \U$10785 ( \11038 , \11031 , \11037 );
or \U$10786 ( \11039 , \11036 , \10097 );
nand \U$10787 ( \11040 , \11038 , \11039 );
and \U$10788 ( \11041 , \11030 , \11040 );
and \U$10789 ( \11042 , \11018 , \11029 );
or \U$10790 ( \11043 , \11041 , \11042 );
not \U$10791 ( \11044 , \11043 );
or \U$10792 ( \11045 , \11010 , \11044 );
not \U$10793 ( \11046 , \11008 );
nand \U$10794 ( \11047 , \11046 , \10692 );
nand \U$10795 ( \11048 , \11045 , \11047 );
xor \U$10796 ( \11049 , \10090 , \10121 );
xnor \U$10797 ( \11050 , \11049 , \10104 );
not \U$10798 ( \11051 , \11050 );
xor \U$10799 ( \11052 , \9850 , \9964 );
xor \U$10800 ( \11053 , \11052 , \10070 );
nand \U$10801 ( \11054 , \11051 , \11053 );
not \U$10802 ( \11055 , \11054 );
nor \U$10803 ( \11056 , \11048 , \11055 );
or \U$10804 ( \11057 , \10625 , \11056 );
nand \U$10805 ( \11058 , \11048 , \11055 );
nand \U$10806 ( \11059 , \11057 , \11058 );
not \U$10807 ( \11060 , \11059 );
not \U$10808 ( \11061 , \11060 );
xor \U$10809 ( \11062 , \10073 , \10123 );
xor \U$10810 ( \11063 , \11062 , \10147 );
not \U$10811 ( \11064 , \11063 );
not \U$10812 ( \11065 , \10153 );
not \U$10813 ( \11066 , \10156 );
and \U$10814 ( \11067 , \11065 , \11066 );
and \U$10815 ( \11068 , \10153 , \10156 );
nor \U$10816 ( \11069 , \11067 , \11068 );
nand \U$10817 ( \11070 , \11064 , \11069 );
xor \U$10818 ( \11071 , \9756 , \9758 );
xor \U$10819 ( \11072 , \11071 , \9766 );
and \U$10820 ( \11073 , \11070 , \11072 );
nor \U$10821 ( \11074 , \11064 , \11069 );
nor \U$10822 ( \11075 , \11073 , \11074 );
not \U$10823 ( \11076 , \11075 );
or \U$10824 ( \11077 , \11061 , \11076 );
xor \U$10825 ( \11078 , \10165 , \10164 );
xor \U$10826 ( \11079 , \11078 , \10172 );
nand \U$10827 ( \11080 , \11077 , \11079 );
or \U$10828 ( \11081 , \11060 , \11075 );
and \U$10829 ( \11082 , \11080 , \11081 );
xor \U$10830 ( \11083 , \10594 , \11082 );
xor \U$10831 ( \11084 , \10162 , \10175 );
xor \U$10832 ( \11085 , \11084 , \10178 );
and \U$10833 ( \11086 , \11083 , \11085 );
and \U$10834 ( \11087 , \10594 , \11082 );
or \U$10835 ( \11088 , \11086 , \11087 );
nor \U$10836 ( \11089 , \10592 , \11088 );
xor \U$10837 ( \11090 , \10590 , \11089 );
and \U$10838 ( \11091 , \9736 , \10214 , \10585 , \11090 );
buf \U$10839 ( \11092 , \11091 );
xor \U$10840 ( \11093 , \10229 , \10233 );
and \U$10841 ( \11094 , \11093 , \10582 );
and \U$10842 ( \11095 , \10229 , \10233 );
or \U$10843 ( \11096 , \11094 , \11095 );
not \U$10844 ( \11097 , \11096 );
not \U$10845 ( \11098 , \10556 );
not \U$10846 ( \11099 , \10562 );
or \U$10847 ( \11100 , \11098 , \11099 );
or \U$10848 ( \11101 , \10562 , \10556 );
not \U$10849 ( \11102 , \10567 );
nand \U$10850 ( \11103 , \11101 , \11102 );
nand \U$10851 ( \11104 , \11100 , \11103 );
not \U$10852 ( \11105 , \10547 );
not \U$10853 ( \11106 , \10542 );
or \U$10854 ( \11107 , \11105 , \11106 );
nand \U$10855 ( \11108 , \11107 , \10538 );
or \U$10856 ( \11109 , \10542 , \10547 );
nand \U$10857 ( \11110 , \11108 , \11109 );
xor \U$10858 ( \11111 , \11104 , \11110 );
not \U$10859 ( \11112 , \10499 );
not \U$10860 ( \11113 , \10527 );
or \U$10861 ( \11114 , \11112 , \11113 );
or \U$10862 ( \11115 , \10499 , \10527 );
nand \U$10863 ( \11116 , \11115 , \10482 );
nand \U$10864 ( \11117 , \11114 , \11116 );
xor \U$10865 ( \11118 , \11111 , \11117 );
not \U$10866 ( \11119 , RIbe29038_46);
not \U$10867 ( \11120 , \4021 );
or \U$10868 ( \11121 , \11119 , \11120 );
nand \U$10869 ( \11122 , \4027 , RIbe28fc0_45);
nand \U$10870 ( \11123 , \11121 , \11122 );
and \U$10871 ( \11124 , \11123 , \4821 );
not \U$10872 ( \11125 , \11123 );
and \U$10873 ( \11126 , \11125 , \3471 );
nor \U$10874 ( \11127 , \11124 , \11126 );
not \U$10875 ( \11128 , \4946 );
not \U$10876 ( \11129 , RIbe27d78_6);
not \U$10877 ( \11130 , \5727 );
or \U$10878 ( \11131 , \11129 , \11130 );
nand \U$10879 ( \11132 , \5731 , RIbe27d00_5);
nand \U$10880 ( \11133 , \11131 , \11132 );
not \U$10881 ( \11134 , \11133 );
or \U$10882 ( \11135 , \11128 , \11134 );
or \U$10883 ( \11136 , \11133 , \4592 );
nand \U$10884 ( \11137 , \11135 , \11136 );
xor \U$10885 ( \11138 , \11127 , \11137 );
not \U$10886 ( \11139 , RIbe290b0_47);
not \U$10887 ( \11140 , \4804 );
or \U$10888 ( \11141 , \11139 , \11140 );
nand \U$10889 ( \11142 , \4809 , RIbe29a88_68);
nand \U$10890 ( \11143 , \11141 , \11142 );
not \U$10891 ( \11144 , \11143 );
not \U$10892 ( \11145 , \4323 );
and \U$10893 ( \11146 , \11144 , \11145 );
and \U$10894 ( \11147 , \11143 , \4323 );
nor \U$10895 ( \11148 , \11146 , \11147 );
xor \U$10896 ( \11149 , \11138 , \11148 );
nand \U$10897 ( \11150 , \6537 , RIbe27b98_2);
and \U$10898 ( \11151 , \11150 , \7546 );
not \U$10899 ( \11152 , \11150 );
and \U$10900 ( \11153 , \11152 , \6546 );
nor \U$10901 ( \11154 , \11151 , \11153 );
not \U$10902 ( \11155 , RIbe28de0_41);
not \U$10903 ( \11156 , \8231 );
or \U$10904 ( \11157 , \11155 , \11156 );
nand \U$10905 ( \11158 , \6617 , RIbe29920_65);
nand \U$10906 ( \11159 , \11157 , \11158 );
and \U$10907 ( \11160 , \11159 , \6144 );
not \U$10908 ( \11161 , \11159 );
and \U$10909 ( \11162 , \11161 , \10972 );
nor \U$10910 ( \11163 , \11160 , \11162 );
xor \U$10911 ( \11164 , \11154 , \11163 );
and \U$10912 ( \11165 , \5455 , RIbe27c10_3);
and \U$10913 ( \11166 , \5751 , RIbe28e58_42);
nor \U$10914 ( \11167 , \11165 , \11166 );
and \U$10915 ( \11168 , \11167 , \5754 );
not \U$10916 ( \11169 , \11167 );
and \U$10917 ( \11170 , \11169 , \10272 );
nor \U$10918 ( \11171 , \11168 , \11170 );
xor \U$10919 ( \11172 , \11164 , \11171 );
xor \U$10920 ( \11173 , \11149 , \11172 );
not \U$10921 ( \11174 , \10475 );
not \U$10922 ( \11175 , \10406 );
or \U$10923 ( \11176 , \11174 , \11175 );
or \U$10924 ( \11177 , \10406 , \10475 );
nand \U$10925 ( \11178 , \11177 , \10434 );
nand \U$10926 ( \11179 , \11176 , \11178 );
xor \U$10927 ( \11180 , \11173 , \11179 );
not \U$10928 ( \11181 , RIbe28480_21);
not \U$10929 ( \11182 , \2531 );
or \U$10930 ( \11183 , \11181 , \11182 );
nand \U$10931 ( \11184 , \1180 , RIbe28408_20);
nand \U$10932 ( \11185 , \11183 , \11184 );
and \U$10933 ( \11186 , \11185 , \1621 );
not \U$10934 ( \11187 , \11185 );
and \U$10935 ( \11188 , \11187 , \1618 );
nor \U$10936 ( \11189 , \11186 , \11188 );
not \U$10937 ( \11190 , \11189 );
and \U$10938 ( \11191 , \5973 , RIbe28390_19);
and \U$10939 ( \11192 , \1203 , RIbe28b10_35);
nor \U$10940 ( \11193 , \11191 , \11192 );
and \U$10941 ( \11194 , \11193 , \1011 );
not \U$10942 ( \11195 , \11193 );
and \U$10943 ( \11196 , \11195 , \1813 );
nor \U$10944 ( \11197 , \11194 , \11196 );
not \U$10945 ( \11198 , \11197 );
or \U$10946 ( \11199 , \11190 , \11198 );
not \U$10947 ( \11200 , \11189 );
not \U$10948 ( \11201 , \11197 );
nand \U$10949 ( \11202 , \11200 , \11201 );
nand \U$10950 ( \11203 , \11199 , \11202 );
not \U$10951 ( \11204 , RIbe285e8_24);
not \U$10952 ( \11205 , \1237 );
or \U$10953 ( \11206 , \11204 , \11205 );
nand \U$10954 ( \11207 , \552 , RIbe287c8_28);
nand \U$10955 ( \11208 , \11206 , \11207 );
not \U$10956 ( \11209 , \11208 );
not \U$10957 ( \11210 , \1246 );
and \U$10958 ( \11211 , \11209 , \11210 );
and \U$10959 ( \11212 , \11208 , \1764 );
nor \U$10960 ( \11213 , \11211 , \11212 );
and \U$10961 ( \11214 , \11203 , \11213 );
not \U$10962 ( \11215 , \11203 );
not \U$10963 ( \11216 , \11213 );
and \U$10964 ( \11217 , \11215 , \11216 );
nor \U$10965 ( \11218 , \11214 , \11217 );
not \U$10966 ( \11219 , \11218 );
not \U$10967 ( \11220 , \11219 );
not \U$10968 ( \11221 , RIbe28a20_33);
not \U$10969 ( \11222 , \5476 );
or \U$10970 ( \11223 , \11221 , \11222 );
nand \U$10971 ( \11224 , \1455 , RIbe289a8_32);
nand \U$10972 ( \11225 , \11223 , \11224 );
and \U$10973 ( \11226 , \11225 , \1309 );
not \U$10974 ( \11227 , \11225 );
and \U$10975 ( \11228 , \11227 , \5125 );
nor \U$10976 ( \11229 , \11226 , \11228 );
not \U$10977 ( \11230 , RIbe28b88_36);
not \U$10978 ( \11231 , \1143 );
or \U$10979 ( \11232 , \11230 , \11231 );
nand \U$10980 ( \11233 , \1147 , RIbe29290_51);
nand \U$10981 ( \11234 , \11232 , \11233 );
and \U$10982 ( \11235 , \11234 , \7899 );
not \U$10983 ( \11236 , \11234 );
and \U$10984 ( \11237 , \11236 , \3994 );
nor \U$10985 ( \11238 , \11235 , \11237 );
xor \U$10986 ( \11239 , \11229 , \11238 );
and \U$10987 ( \11240 , \2557 , RIbe28930_31);
and \U$10988 ( \11241 , \1117 , RIbe29560_57);
nor \U$10989 ( \11242 , \11240 , \11241 );
and \U$10990 ( \11243 , \11242 , \1125 );
not \U$10991 ( \11244 , \11242 );
and \U$10992 ( \11245 , \11244 , \1132 );
nor \U$10993 ( \11246 , \11243 , \11245 );
xor \U$10994 ( \11247 , \11239 , \11246 );
not \U$10995 ( \11248 , \11247 );
not \U$10996 ( \11249 , \11248 );
or \U$10997 ( \11250 , \11220 , \11249 );
nand \U$10998 ( \11251 , \11247 , \11218 );
nand \U$10999 ( \11252 , \11250 , \11251 );
not \U$11000 ( \11253 , RIbe296c8_60);
not \U$11001 ( \11254 , \3685 );
or \U$11002 ( \11255 , \11253 , \11254 );
nand \U$11003 ( \11256 , \4011 , RIbe29650_59);
nand \U$11004 ( \11257 , \11255 , \11256 );
and \U$11005 ( \11258 , \11257 , \3290 );
not \U$11006 ( \11259 , \11257 );
and \U$11007 ( \11260 , \11259 , \3461 );
nor \U$11008 ( \11261 , \11258 , \11260 );
not \U$11009 ( \11262 , \11261 );
not \U$11010 ( \11263 , \11262 );
not \U$11011 ( \11264 , RIbe280c0_13);
not \U$11012 ( \11265 , \3476 );
or \U$11013 ( \11266 , \11264 , \11265 );
nand \U$11014 ( \11267 , \2901 , RIbe29830_63);
nand \U$11015 ( \11268 , \11266 , \11267 );
not \U$11016 ( \11269 , \11268 );
not \U$11017 ( \11270 , \2379 );
and \U$11018 ( \11271 , \11269 , \11270 );
and \U$11019 ( \11272 , \11268 , \2379 );
nor \U$11020 ( \11273 , \11271 , \11272 );
not \U$11021 ( \11274 , \11273 );
not \U$11022 ( \11275 , \11274 );
or \U$11023 ( \11276 , \11263 , \11275 );
nand \U$11024 ( \11277 , \11261 , \11273 );
nand \U$11025 ( \11278 , \11276 , \11277 );
not \U$11026 ( \11279 , \2385 );
not \U$11027 ( \11280 , \3663 );
and \U$11028 ( \11281 , \11279 , \11280 );
and \U$11029 ( \11282 , \8833 , RIbe28228_16);
nor \U$11030 ( \11283 , \11281 , \11282 );
and \U$11031 ( \11284 , \11283 , \1277 );
not \U$11032 ( \11285 , \11283 );
and \U$11033 ( \11286 , \11285 , \1076 );
or \U$11034 ( \11287 , \11284 , \11286 );
xnor \U$11035 ( \11288 , \11278 , \11287 );
not \U$11036 ( \11289 , \11288 );
and \U$11037 ( \11290 , \11252 , \11289 );
not \U$11038 ( \11291 , \11252 );
and \U$11039 ( \11292 , \11291 , \11288 );
nor \U$11040 ( \11293 , \11290 , \11292 );
xor \U$11041 ( \11294 , \11180 , \11293 );
xor \U$11042 ( \11295 , \11118 , \11294 );
xor \U$11043 ( \11296 , \10483 , \10490 );
and \U$11044 ( \11297 , \11296 , \10498 );
and \U$11045 ( \11298 , \10483 , \10490 );
or \U$11046 ( \11299 , \11297 , \11298 );
nand \U$11047 ( \11300 , RIbe29380_53, RIbe29dd0_75);
and \U$11048 ( \11301 , \325 , RIbe29c68_72);
and \U$11049 ( \11302 , \329 , RIbe29bf0_71);
nor \U$11050 ( \11303 , \11301 , \11302 );
and \U$11051 ( \11304 , \11303 , \1375 );
not \U$11052 ( \11305 , \11303 );
and \U$11053 ( \11306 , \11305 , \339 );
nor \U$11054 ( \11307 , \11304 , \11306 );
or \U$11055 ( \11308 , \11300 , \11307 );
nand \U$11056 ( \11309 , \11307 , \11300 );
nand \U$11057 ( \11310 , \11308 , \11309 );
xor \U$11058 ( \11311 , \11299 , \11310 );
and \U$11059 ( \11312 , \5365 , RIbe27fd0_11);
and \U$11060 ( \11313 , \3897 , RIbe27f58_10);
nor \U$11061 ( \11314 , \11312 , \11313 );
and \U$11062 ( \11315 , \11314 , \300 );
not \U$11063 ( \11316 , \11314 );
and \U$11064 ( \11317 , \11316 , \293 );
nor \U$11065 ( \11318 , \11315 , \11317 );
and \U$11066 ( \11319 , \261 , RIbe28f48_44);
and \U$11067 ( \11320 , \264 , RIbe28ed0_43);
nor \U$11068 ( \11321 , \11319 , \11320 );
and \U$11069 ( \11322 , \11321 , \1362 );
not \U$11070 ( \11323 , \11321 );
and \U$11071 ( \11324 , \11323 , \269 );
nor \U$11072 ( \11325 , \11322 , \11324 );
xor \U$11073 ( \11326 , \11318 , \11325 );
not \U$11074 ( \11327 , RIbe27e68_8);
not \U$11075 ( \11328 , \383 );
or \U$11076 ( \11329 , \11327 , \11328 );
nand \U$11077 ( \11330 , \429 , RIbe28660_25);
nand \U$11078 ( \11331 , \11329 , \11330 );
and \U$11079 ( \11332 , \11331 , \306 );
not \U$11080 ( \11333 , \11331 );
and \U$11081 ( \11334 , \11333 , \3175 );
nor \U$11082 ( \11335 , \11332 , \11334 );
xor \U$11083 ( \11336 , \11326 , \11335 );
xor \U$11084 ( \11337 , \11311 , \11336 );
or \U$11085 ( \11338 , \10367 , \6602 );
nand \U$11086 ( \11339 , \11338 , \10353 );
nand \U$11087 ( \11340 , \10367 , \8957 );
nand \U$11088 ( \11341 , \11339 , \11340 );
or \U$11089 ( \11342 , \10285 , \10265 );
nand \U$11090 ( \11343 , \11342 , \10276 );
nand \U$11091 ( \11344 , \10265 , \10285 );
nand \U$11092 ( \11345 , \11343 , \11344 );
xor \U$11093 ( \11346 , \11341 , \11345 );
not \U$11094 ( \11347 , \10393 );
not \U$11095 ( \11348 , \10405 );
or \U$11096 ( \11349 , \11347 , \11348 );
or \U$11097 ( \11350 , \10405 , \10393 );
nand \U$11098 ( \11351 , \11350 , \10381 );
nand \U$11099 ( \11352 , \11349 , \11351 );
xor \U$11100 ( \11353 , \11346 , \11352 );
xor \U$11101 ( \11354 , \11337 , \11353 );
not \U$11102 ( \11355 , \10452 );
not \U$11103 ( \11356 , \10466 );
or \U$11104 ( \11357 , \11355 , \11356 );
nand \U$11105 ( \11358 , \11357 , \10444 );
nand \U$11106 ( \11359 , \10467 , \10455 );
nand \U$11107 ( \11360 , \11358 , \11359 );
xor \U$11108 ( \11361 , \10416 , \10425 );
and \U$11109 ( \11362 , \11361 , \10433 );
and \U$11110 ( \11363 , \10416 , \10425 );
or \U$11111 ( \11364 , \11362 , \11363 );
xor \U$11112 ( \11365 , \11360 , \11364 );
xor \U$11113 ( \11366 , \10509 , \10518 );
and \U$11114 ( \11367 , \11366 , \10526 );
and \U$11115 ( \11368 , \10509 , \10518 );
or \U$11116 ( \11369 , \11367 , \11368 );
xor \U$11117 ( \11370 , \11365 , \11369 );
xor \U$11118 ( \11371 , \11354 , \11370 );
xor \U$11119 ( \11372 , \11295 , \11371 );
not \U$11120 ( \11373 , \10572 );
nand \U$11121 ( \11374 , \11373 , \10548 );
not \U$11122 ( \11375 , \11374 );
not \U$11123 ( \11376 , \10533 );
or \U$11124 ( \11377 , \11375 , \11376 );
not \U$11125 ( \11378 , \10548 );
nand \U$11126 ( \11379 , \11378 , \10572 );
nand \U$11127 ( \11380 , \11377 , \11379 );
xor \U$11128 ( \11381 , \10322 , \10330 );
and \U$11129 ( \11382 , \11381 , \10337 );
and \U$11130 ( \11383 , \10322 , \10330 );
or \U$11131 ( \11384 , \11382 , \11383 );
and \U$11132 ( \11385 , \11380 , \11384 );
not \U$11133 ( \11386 , \11380 );
not \U$11134 ( \11387 , \11384 );
and \U$11135 ( \11388 , \11386 , \11387 );
nor \U$11136 ( \11389 , \11385 , \11388 );
xnor \U$11137 ( \11390 , \11372 , \11389 );
or \U$11138 ( \11391 , \10305 , \10240 );
and \U$11139 ( \11392 , \11391 , \10581 );
and \U$11140 ( \11393 , \10240 , \10305 );
nor \U$11141 ( \11394 , \11392 , \11393 );
xor \U$11142 ( \11395 , \11390 , \11394 );
not \U$11143 ( \11396 , \10307 );
not \U$11144 ( \11397 , \10316 );
or \U$11145 ( \11398 , \11396 , \11397 );
nand \U$11146 ( \11399 , \11398 , \10311 );
or \U$11147 ( \11400 , \10316 , \10307 );
and \U$11148 ( \11401 , \11399 , \11400 );
not \U$11149 ( \11402 , \11401 );
xor \U$11150 ( \11403 , \10287 , \10291 );
and \U$11151 ( \11404 , \11403 , \10296 );
and \U$11152 ( \11405 , \10287 , \10291 );
or \U$11153 ( \11406 , \11404 , \11405 );
not \U$11154 ( \11407 , \11406 );
or \U$11155 ( \11408 , \11402 , \11407 );
or \U$11156 ( \11409 , \11406 , \11401 );
nand \U$11157 ( \11410 , \11408 , \11409 );
not \U$11158 ( \11411 , \11410 );
and \U$11159 ( \11412 , \10528 , \10372 );
xnor \U$11160 ( \11413 , \10477 , \10406 );
nor \U$11161 ( \11414 , \11412 , \11413 );
nor \U$11162 ( \11415 , \10528 , \10372 );
nor \U$11163 ( \11416 , \11414 , \11415 );
not \U$11164 ( \11417 , \11416 );
and \U$11165 ( \11418 , \11411 , \11417 );
and \U$11166 ( \11419 , \11410 , \11416 );
nor \U$11167 ( \11420 , \11418 , \11419 );
or \U$11168 ( \11421 , \10248 , \10297 );
not \U$11169 ( \11422 , \10255 );
nand \U$11170 ( \11423 , \11421 , \11422 );
nand \U$11171 ( \11424 , \10248 , \10297 );
and \U$11172 ( \11425 , \11423 , \11424 );
xor \U$11173 ( \11426 , \11420 , \11425 );
not \U$11174 ( \11427 , \10317 );
and \U$11175 ( \11428 , \10580 , \11427 );
nor \U$11176 ( \11429 , \11428 , \10339 );
nor \U$11177 ( \11430 , \10580 , \11427 );
nor \U$11178 ( \11431 , \11429 , \11430 );
xor \U$11179 ( \11432 , \11426 , \11431 );
xor \U$11180 ( \11433 , \11395 , \11432 );
nor \U$11181 ( \11434 , \11097 , \11433 );
not \U$11182 ( \11435 , \11434 );
xor \U$11183 ( \11436 , \11420 , \11425 );
and \U$11184 ( \11437 , \11436 , \11431 );
and \U$11185 ( \11438 , \11420 , \11425 );
or \U$11186 ( \11439 , \11437 , \11438 );
xor \U$11187 ( \11440 , \11104 , \11110 );
and \U$11188 ( \11441 , \11440 , \11117 );
and \U$11189 ( \11442 , \11104 , \11110 );
or \U$11190 ( \11443 , \11441 , \11442 );
xor \U$11191 ( \11444 , \11337 , \11353 );
and \U$11192 ( \11445 , \11444 , \11370 );
and \U$11193 ( \11446 , \11337 , \11353 );
or \U$11194 ( \11447 , \11445 , \11446 );
xor \U$11195 ( \11448 , \11443 , \11447 );
xor \U$11196 ( \11449 , \11173 , \11179 );
and \U$11197 ( \11450 , \11449 , \11293 );
and \U$11198 ( \11451 , \11173 , \11179 );
or \U$11199 ( \11452 , \11450 , \11451 );
xor \U$11200 ( \11453 , \11448 , \11452 );
not \U$11201 ( \11454 , \11274 );
not \U$11202 ( \11455 , \11261 );
or \U$11203 ( \11456 , \11454 , \11455 );
nand \U$11204 ( \11457 , \11262 , \11273 );
nand \U$11205 ( \11458 , \11457 , \11287 );
nand \U$11206 ( \11459 , \11456 , \11458 );
xor \U$11207 ( \11460 , \11154 , \11163 );
and \U$11208 ( \11461 , \11460 , \11171 );
and \U$11209 ( \11462 , \11154 , \11163 );
or \U$11210 ( \11463 , \11461 , \11462 );
not \U$11211 ( \11464 , \11148 );
not \U$11212 ( \11465 , \11127 );
or \U$11213 ( \11466 , \11464 , \11465 );
nand \U$11214 ( \11467 , \11466 , \11137 );
or \U$11215 ( \11468 , \11127 , \11148 );
nand \U$11216 ( \11469 , \11467 , \11468 );
xor \U$11217 ( \11470 , \11463 , \11469 );
xor \U$11218 ( \11471 , \11459 , \11470 );
and \U$11219 ( \11472 , \326 , RIbe29bf0_71);
and \U$11220 ( \11473 , \330 , RIbe28f48_44);
nor \U$11221 ( \11474 , \11472 , \11473 );
and \U$11222 ( \11475 , \11474 , \1379 );
not \U$11223 ( \11476 , \11474 );
and \U$11224 ( \11477 , \11476 , \1378 );
nor \U$11225 ( \11478 , \11475 , \11477 );
and \U$11226 ( \11479 , RIbe29380_53, RIbe29c68_72);
xor \U$11227 ( \11480 , \11478 , \11479 );
xor \U$11228 ( \11481 , \11480 , \11309 );
not \U$11229 ( \11482 , \11213 );
not \U$11230 ( \11483 , \11197 );
or \U$11231 ( \11484 , \11482 , \11483 );
nand \U$11232 ( \11485 , \11484 , \11189 );
nand \U$11233 ( \11486 , \11201 , \11216 );
nand \U$11234 ( \11487 , \11485 , \11486 );
xor \U$11235 ( \11488 , \11229 , \11238 );
and \U$11236 ( \11489 , \11488 , \11246 );
and \U$11237 ( \11490 , \11229 , \11238 );
or \U$11238 ( \11491 , \11489 , \11490 );
xor \U$11239 ( \11492 , \11487 , \11491 );
xor \U$11240 ( \11493 , \11318 , \11325 );
and \U$11241 ( \11494 , \11493 , \11335 );
and \U$11242 ( \11495 , \11318 , \11325 );
or \U$11243 ( \11496 , \11494 , \11495 );
xor \U$11244 ( \11497 , \11492 , \11496 );
xor \U$11245 ( \11498 , \11481 , \11497 );
not \U$11246 ( \11499 , RIbe289a8_32);
not \U$11247 ( \11500 , \1633 );
or \U$11248 ( \11501 , \11499 , \11500 );
nand \U$11249 ( \11502 , \1099 , RIbe28930_31);
nand \U$11250 ( \11503 , \11501 , \11502 );
and \U$11251 ( \11504 , \11503 , \1309 );
not \U$11252 ( \11505 , \11503 );
and \U$11253 ( \11506 , \11505 , \5125 );
nor \U$11254 ( \11507 , \11504 , \11506 );
and \U$11255 ( \11508 , \6380 , RIbe29560_57);
and \U$11256 ( \11509 , \5467 , RIbe28228_16);
nor \U$11257 ( \11510 , \11508 , \11509 );
and \U$11258 ( \11511 , \11510 , \1131 );
not \U$11259 ( \11512 , \11510 );
and \U$11260 ( \11513 , \11512 , \3491 );
nor \U$11261 ( \11514 , \11511 , \11513 );
and \U$11262 ( \11515 , \11507 , \11514 );
not \U$11263 ( \11516 , \11507 );
not \U$11264 ( \11517 , \11514 );
and \U$11265 ( \11518 , \11516 , \11517 );
or \U$11266 ( \11519 , \11515 , \11518 );
not \U$11267 ( \11520 , RIbe29290_51);
not \U$11268 ( \11521 , \1143 );
or \U$11269 ( \11522 , \11520 , \11521 );
nand \U$11270 ( \11523 , \1147 , RIbe28a20_33);
nand \U$11271 ( \11524 , \11522 , \11523 );
not \U$11272 ( \11525 , \11524 );
not \U$11273 ( \11526 , \1152 );
and \U$11274 ( \11527 , \11525 , \11526 );
and \U$11275 ( \11528 , \11524 , \8327 );
nor \U$11276 ( \11529 , \11527 , \11528 );
not \U$11277 ( \11530 , \11529 );
and \U$11278 ( \11531 , \11519 , \11530 );
not \U$11279 ( \11532 , \11519 );
and \U$11280 ( \11533 , \11532 , \11529 );
nor \U$11281 ( \11534 , \11531 , \11533 );
not \U$11282 ( \11535 , RIbe28408_20);
not \U$11283 ( \11536 , \7363 );
or \U$11284 ( \11537 , \11535 , \11536 );
nand \U$11285 ( \11538 , \1180 , RIbe28390_19);
nand \U$11286 ( \11539 , \11537 , \11538 );
xor \U$11287 ( \11540 , \11539 , \564 );
not \U$11288 ( \11541 , \11540 );
not \U$11289 ( \11542 , \11541 );
and \U$11290 ( \11543 , \1807 , RIbe28b10_35);
and \U$11291 ( \11544 , \1165 , RIbe28b88_36);
nor \U$11292 ( \11545 , \11543 , \11544 );
and \U$11293 ( \11546 , \11545 , \1608 );
not \U$11294 ( \11547 , \11545 );
and \U$11295 ( \11548 , \11547 , \1011 );
nor \U$11296 ( \11549 , \11546 , \11548 );
not \U$11297 ( \11550 , \11549 );
not \U$11298 ( \11551 , \11550 );
or \U$11299 ( \11552 , \11542 , \11551 );
nand \U$11300 ( \11553 , \11549 , \11540 );
nand \U$11301 ( \11554 , \11552 , \11553 );
not \U$11302 ( \11555 , RIbe287c8_28);
not \U$11303 ( \11556 , \3244 );
or \U$11304 ( \11557 , \11555 , \11556 );
nand \U$11305 ( \11558 , \553 , RIbe28480_21);
nand \U$11306 ( \11559 , \11557 , \11558 );
not \U$11307 ( \11560 , \11559 );
not \U$11308 ( \11561 , \1333 );
and \U$11309 ( \11562 , \11560 , \11561 );
and \U$11310 ( \11563 , \11559 , \1333 );
nor \U$11311 ( \11564 , \11562 , \11563 );
xnor \U$11312 ( \11565 , \11554 , \11564 );
xor \U$11313 ( \11566 , \11534 , \11565 );
and \U$11314 ( \11567 , \1254 , RIbe27f58_10);
and \U$11315 ( \11568 , \287 , RIbe27e68_8);
nor \U$11316 ( \11569 , \11567 , \11568 );
and \U$11317 ( \11570 , \11569 , \300 );
not \U$11318 ( \11571 , \11569 );
and \U$11319 ( \11572 , \11571 , \293 );
nor \U$11320 ( \11573 , \11570 , \11572 );
not \U$11321 ( \11574 , RIbe28660_25);
not \U$11322 ( \11575 , \1337 );
or \U$11323 ( \11576 , \11574 , \11575 );
nand \U$11324 ( \11577 , \429 , RIbe285e8_24);
nand \U$11325 ( \11578 , \11576 , \11577 );
not \U$11326 ( \11579 , \11578 );
not \U$11327 ( \11580 , \3175 );
and \U$11328 ( \11581 , \11579 , \11580 );
and \U$11329 ( \11582 , \11578 , \3175 );
nor \U$11330 ( \11583 , \11581 , \11582 );
not \U$11331 ( \11584 , \11583 );
and \U$11332 ( \11585 , \11573 , \11584 );
not \U$11333 ( \11586 , \11573 );
and \U$11334 ( \11587 , \11586 , \11583 );
nor \U$11335 ( \11588 , \11585 , \11587 );
and \U$11336 ( \11589 , \1659 , RIbe28ed0_43);
and \U$11337 ( \11590 , \1831 , RIbe27fd0_11);
nor \U$11338 ( \11591 , \11589 , \11590 );
and \U$11339 ( \11592 , \11591 , \269 );
not \U$11340 ( \11593 , \11591 );
and \U$11341 ( \11594 , \11593 , \1362 );
nor \U$11342 ( \11595 , \11592 , \11594 );
not \U$11343 ( \11596 , \11595 );
and \U$11344 ( \11597 , \11588 , \11596 );
not \U$11345 ( \11598 , \11588 );
and \U$11346 ( \11599 , \11598 , \11595 );
nor \U$11347 ( \11600 , \11597 , \11599 );
xor \U$11348 ( \11601 , \11566 , \11600 );
xor \U$11349 ( \11602 , \11498 , \11601 );
xor \U$11350 ( \11603 , \11471 , \11602 );
not \U$11351 ( \11604 , \11288 );
not \U$11352 ( \11605 , \11248 );
or \U$11353 ( \11606 , \11604 , \11605 );
nand \U$11354 ( \11607 , \11606 , \11219 );
nand \U$11355 ( \11608 , \11247 , \11289 );
nand \U$11356 ( \11609 , \11607 , \11608 );
and \U$11357 ( \11610 , \11149 , \11172 );
xor \U$11358 ( \11611 , \11609 , \11610 );
not \U$11359 ( \11612 , RIbe29920_65);
not \U$11360 ( \11613 , \8231 );
or \U$11361 ( \11614 , \11612 , \11613 );
nand \U$11362 ( \11615 , \7087 , RIbe27b98_2);
nand \U$11363 ( \11616 , \11614 , \11615 );
and \U$11364 ( \11617 , \11616 , \5741 );
not \U$11365 ( \11618 , \11616 );
and \U$11366 ( \11619 , \11618 , \6141 );
nor \U$11367 ( \11620 , \11617 , \11619 );
xor \U$11368 ( \11621 , \7546 , \11620 );
not \U$11369 ( \11622 , RIbe28e58_42);
not \U$11370 ( \11623 , \5455 );
or \U$11371 ( \11624 , \11622 , \11623 );
nand \U$11372 ( \11625 , \10269 , RIbe28de0_41);
nand \U$11373 ( \11626 , \11624 , \11625 );
and \U$11374 ( \11627 , \11626 , \10272 );
not \U$11375 ( \11628 , \11626 );
and \U$11376 ( \11629 , \11628 , \10984 );
nor \U$11377 ( \11630 , \11627 , \11629 );
xor \U$11378 ( \11631 , \11621 , \11630 );
not \U$11379 ( \11632 , RIbe29a88_68);
not \U$11380 ( \11633 , \4804 );
or \U$11381 ( \11634 , \11632 , \11633 );
nand \U$11382 ( \11635 , \4809 , RIbe27d78_6);
nand \U$11383 ( \11636 , \11634 , \11635 );
xnor \U$11384 ( \11637 , \11636 , \4323 );
not \U$11385 ( \11638 , RIbe27d00_5);
not \U$11386 ( \11639 , \4830 );
or \U$11387 ( \11640 , \11638 , \11639 );
nand \U$11388 ( \11641 , \5052 , RIbe27c10_3);
nand \U$11389 ( \11642 , \11640 , \11641 );
xor \U$11390 ( \11643 , \11642 , \4592 );
xor \U$11391 ( \11644 , \11637 , \11643 );
not \U$11392 ( \11645 , RIbe28fc0_45);
not \U$11393 ( \11646 , \4021 );
or \U$11394 ( \11647 , \11645 , \11646 );
nand \U$11395 ( \11648 , \4027 , RIbe290b0_47);
nand \U$11396 ( \11649 , \11647 , \11648 );
and \U$11397 ( \11650 , \11649 , \4821 );
not \U$11398 ( \11651 , \11649 );
and \U$11399 ( \11652 , \11651 , \3471 );
nor \U$11400 ( \11653 , \11650 , \11652 );
xnor \U$11401 ( \11654 , \11644 , \11653 );
xor \U$11402 ( \11655 , \11631 , \11654 );
not \U$11403 ( \11656 , RIbe29830_63);
not \U$11404 ( \11657 , \2898 );
or \U$11405 ( \11658 , \11656 , \11657 );
nand \U$11406 ( \11659 , \4284 , RIbe296c8_60);
nand \U$11407 ( \11660 , \11658 , \11659 );
and \U$11408 ( \11661 , \11660 , \2380 );
not \U$11409 ( \11662 , \11660 );
and \U$11410 ( \11663 , \11662 , \2379 );
nor \U$11411 ( \11664 , \11661 , \11663 );
not \U$11412 ( \11665 , RIbe29650_59);
not \U$11413 ( \11666 , \3452 );
or \U$11414 ( \11667 , \11665 , \11666 );
nand \U$11415 ( \11668 , \3458 , RIbe29038_46);
nand \U$11416 ( \11669 , \11667 , \11668 );
and \U$11417 ( \11670 , \11669 , \3461 );
not \U$11418 ( \11671 , \11669 );
and \U$11419 ( \11672 , \11671 , \4346 );
nor \U$11420 ( \11673 , \11670 , \11672 );
and \U$11421 ( \11674 , \11664 , \11673 );
not \U$11422 ( \11675 , \11664 );
not \U$11423 ( \11676 , \11673 );
and \U$11424 ( \11677 , \11675 , \11676 );
or \U$11425 ( \11678 , \11674 , \11677 );
not \U$11426 ( \11679 , \2889 );
not \U$11427 ( \11680 , \3537 );
and \U$11428 ( \11681 , \11679 , \11680 );
and \U$11429 ( \11682 , \3303 , RIbe281b0_15);
nor \U$11430 ( \11683 , \11681 , \11682 );
and \U$11431 ( \11684 , \11683 , \1076 );
not \U$11432 ( \11685 , \11683 );
and \U$11433 ( \11686 , \11685 , \1277 );
nor \U$11434 ( \11687 , \11684 , \11686 );
xor \U$11435 ( \11688 , \11678 , \11687 );
xnor \U$11436 ( \11689 , \11655 , \11688 );
xor \U$11437 ( \11690 , \11611 , \11689 );
xor \U$11438 ( \11691 , \11603 , \11690 );
xor \U$11439 ( \11692 , \11453 , \11691 );
not \U$11440 ( \11693 , \11384 );
not \U$11441 ( \11694 , \11380 );
or \U$11442 ( \11695 , \11693 , \11694 );
not \U$11443 ( \11696 , \11380 );
nand \U$11444 ( \11697 , \11696 , \11387 );
nand \U$11445 ( \11698 , \11372 , \11697 );
nand \U$11446 ( \11699 , \11695 , \11698 );
xor \U$11447 ( \11700 , \11692 , \11699 );
xor \U$11448 ( \11701 , \11341 , \11345 );
and \U$11449 ( \11702 , \11701 , \11352 );
and \U$11450 ( \11703 , \11341 , \11345 );
or \U$11451 ( \11704 , \11702 , \11703 );
xor \U$11452 ( \11705 , \11360 , \11364 );
and \U$11453 ( \11706 , \11705 , \11369 );
and \U$11454 ( \11707 , \11360 , \11364 );
or \U$11455 ( \11708 , \11706 , \11707 );
xor \U$11456 ( \11709 , \11704 , \11708 );
xor \U$11457 ( \11710 , \11299 , \11310 );
and \U$11458 ( \11711 , \11710 , \11336 );
and \U$11459 ( \11712 , \11299 , \11310 );
or \U$11460 ( \11713 , \11711 , \11712 );
xor \U$11461 ( \11714 , \11709 , \11713 );
not \U$11462 ( \11715 , \11401 );
not \U$11463 ( \11716 , \11416 );
or \U$11464 ( \11717 , \11715 , \11716 );
nand \U$11465 ( \11718 , \11717 , \11406 );
or \U$11466 ( \11719 , \11416 , \11401 );
nand \U$11467 ( \11720 , \11718 , \11719 );
xor \U$11468 ( \11721 , \11714 , \11720 );
xor \U$11469 ( \11722 , \11118 , \11294 );
and \U$11470 ( \11723 , \11722 , \11371 );
and \U$11471 ( \11724 , \11118 , \11294 );
or \U$11472 ( \11725 , \11723 , \11724 );
xor \U$11473 ( \11726 , \11721 , \11725 );
not \U$11474 ( \11727 , \11726 );
xor \U$11475 ( \11728 , \11700 , \11727 );
xor \U$11476 ( \11729 , \11439 , \11728 );
xor \U$11477 ( \11730 , \11390 , \11394 );
and \U$11478 ( \11731 , \11730 , \11432 );
and \U$11479 ( \11732 , \11390 , \11394 );
or \U$11480 ( \11733 , \11731 , \11732 );
xor \U$11481 ( \11734 , \11729 , \11733 );
not \U$11482 ( \11735 , \11734 );
or \U$11483 ( \11736 , \11435 , \11735 );
or \U$11484 ( \11737 , \11734 , \11434 );
nand \U$11485 ( \11738 , \11736 , \11737 );
buf \U$11486 ( \11739 , \11738 );
and \U$11487 ( \11740 , \10224 , \10583 );
not \U$11488 ( \11741 , \11096 );
not \U$11489 ( \11742 , \11433 );
or \U$11490 ( \11743 , \11741 , \11742 );
or \U$11491 ( \11744 , \11433 , \11096 );
nand \U$11492 ( \11745 , \11743 , \11744 );
xor \U$11493 ( \11746 , \11740 , \11745 );
not \U$11494 ( \11747 , \6097 );
xor \U$11495 ( \11748 , \6088 , \6107 );
not \U$11496 ( \11749 , \11748 );
or \U$11497 ( \11750 , \11747 , \11749 );
or \U$11498 ( \11751 , \11748 , \6097 );
nand \U$11499 ( \11752 , \11750 , \11751 );
not \U$11500 ( \11753 , \11688 );
not \U$11501 ( \11754 , \11631 );
or \U$11502 ( \11755 , \11753 , \11754 );
or \U$11503 ( \11756 , \11688 , \11631 );
not \U$11504 ( \11757 , \11654 );
nand \U$11505 ( \11758 , \11756 , \11757 );
nand \U$11506 ( \11759 , \11755 , \11758 );
xor \U$11507 ( \11760 , \11752 , \11759 );
xor \U$11508 ( \11761 , \11534 , \11565 );
and \U$11509 ( \11762 , \11761 , \11600 );
and \U$11510 ( \11763 , \11534 , \11565 );
or \U$11511 ( \11764 , \11762 , \11763 );
xor \U$11512 ( \11765 , \11760 , \11764 );
xor \U$11513 ( \11766 , \11443 , \11447 );
and \U$11514 ( \11767 , \11766 , \11452 );
and \U$11515 ( \11768 , \11443 , \11447 );
or \U$11516 ( \11769 , \11767 , \11768 );
xor \U$11517 ( \11770 , \11765 , \11769 );
xor \U$11518 ( \11771 , \11471 , \11602 );
and \U$11519 ( \11772 , \11771 , \11690 );
and \U$11520 ( \11773 , \11471 , \11602 );
or \U$11521 ( \11774 , \11772 , \11773 );
xor \U$11522 ( \11775 , \11770 , \11774 );
not \U$11523 ( \11776 , \11699 );
not \U$11524 ( \11777 , \11692 );
or \U$11525 ( \11778 , \11776 , \11777 );
or \U$11526 ( \11779 , \11692 , \11699 );
nand \U$11527 ( \11780 , \11779 , \11726 );
nand \U$11528 ( \11781 , \11778 , \11780 );
xor \U$11529 ( \11782 , \11775 , \11781 );
and \U$11530 ( \11783 , \11453 , \11691 );
xor \U$11531 ( \11784 , \11714 , \11720 );
and \U$11532 ( \11785 , \11784 , \11725 );
and \U$11533 ( \11786 , \11714 , \11720 );
or \U$11534 ( \11787 , \11785 , \11786 );
xor \U$11535 ( \11788 , \11783 , \11787 );
xor \U$11536 ( \11789 , \11478 , \11479 );
and \U$11537 ( \11790 , \11789 , \11309 );
and \U$11538 ( \11791 , \11478 , \11479 );
or \U$11539 ( \11792 , \11790 , \11791 );
or \U$11540 ( \11793 , \11469 , \11459 );
nand \U$11541 ( \11794 , \11793 , \11463 );
nand \U$11542 ( \11795 , \11469 , \11459 );
nand \U$11543 ( \11796 , \11794 , \11795 );
xor \U$11544 ( \11797 , \11792 , \11796 );
xor \U$11545 ( \11798 , \11487 , \11491 );
and \U$11546 ( \11799 , \11798 , \11496 );
and \U$11547 ( \11800 , \11487 , \11491 );
or \U$11548 ( \11801 , \11799 , \11800 );
xor \U$11549 ( \11802 , \11797 , \11801 );
not \U$11550 ( \11803 , \11676 );
not \U$11551 ( \11804 , \11664 );
or \U$11552 ( \11805 , \11803 , \11804 );
or \U$11553 ( \11806 , \11664 , \11676 );
nand \U$11554 ( \11807 , \11806 , \11687 );
nand \U$11555 ( \11808 , \11805 , \11807 );
xor \U$11556 ( \11809 , \7546 , \11620 );
and \U$11557 ( \11810 , \11809 , \11630 );
and \U$11558 ( \11811 , \7546 , \11620 );
or \U$11559 ( \11812 , \11810 , \11811 );
xor \U$11560 ( \11813 , \11808 , \11812 );
or \U$11561 ( \11814 , \11653 , \11643 );
not \U$11562 ( \11815 , \11643 );
not \U$11563 ( \11816 , \11653 );
or \U$11564 ( \11817 , \11815 , \11816 );
nand \U$11565 ( \11818 , \11817 , \11637 );
nand \U$11566 ( \11819 , \11814 , \11818 );
xor \U$11567 ( \11820 , \11813 , \11819 );
nand \U$11568 ( \11821 , \11550 , \11564 );
and \U$11569 ( \11822 , \11821 , \11541 );
nor \U$11570 ( \11823 , \11564 , \11550 );
nor \U$11571 ( \11824 , \11822 , \11823 );
not \U$11572 ( \11825 , \11824 );
not \U$11573 ( \11826 , \11517 );
not \U$11574 ( \11827 , \11530 );
or \U$11575 ( \11828 , \11826 , \11827 );
nand \U$11576 ( \11829 , \11514 , \11529 );
nand \U$11577 ( \11830 , \11829 , \11507 );
nand \U$11578 ( \11831 , \11828 , \11830 );
not \U$11579 ( \11832 , \11831 );
or \U$11580 ( \11833 , \11825 , \11832 );
or \U$11581 ( \11834 , \11831 , \11824 );
nand \U$11582 ( \11835 , \11833 , \11834 );
not \U$11583 ( \11836 , \11596 );
not \U$11584 ( \11837 , \11584 );
or \U$11585 ( \11838 , \11836 , \11837 );
nand \U$11586 ( \11839 , \11583 , \11595 );
nand \U$11587 ( \11840 , \11839 , \11573 );
nand \U$11588 ( \11841 , \11838 , \11840 );
xor \U$11589 ( \11842 , \11835 , \11841 );
xor \U$11590 ( \11843 , \11820 , \11842 );
xor \U$11591 ( \11844 , \6062 , \6070 );
xnor \U$11592 ( \11845 , \11844 , \6050 );
nand \U$11593 ( \11846 , RIbe29380_53, RIbe29bf0_71);
or \U$11594 ( \11847 , \11845 , \11846 );
nand \U$11595 ( \11848 , \11845 , \11846 );
nand \U$11596 ( \11849 , \11847 , \11848 );
not \U$11597 ( \11850 , \6132 );
not \U$11598 ( \11851 , \6146 );
not \U$11599 ( \11852 , \6123 );
or \U$11600 ( \11853 , \11851 , \11852 );
or \U$11601 ( \11854 , \6123 , \6146 );
nand \U$11602 ( \11855 , \11853 , \11854 );
not \U$11603 ( \11856 , \11855 );
or \U$11604 ( \11857 , \11850 , \11856 );
or \U$11605 ( \11858 , \11855 , \6132 );
nand \U$11606 ( \11859 , \11857 , \11858 );
xor \U$11607 ( \11860 , \11849 , \11859 );
xor \U$11608 ( \11861 , \6160 , \6167 );
xor \U$11609 ( \11862 , \11861 , \6175 );
and \U$11610 ( \11863 , \5990 , \6000 );
not \U$11611 ( \11864 , \5990 );
and \U$11612 ( \11865 , \11864 , \6001 );
or \U$11613 ( \11866 , \11863 , \11865 );
xor \U$11614 ( \11867 , \11866 , \5980 );
and \U$11615 ( \11868 , \11862 , \11867 );
not \U$11616 ( \11869 , \11862 );
not \U$11617 ( \11870 , \11867 );
and \U$11618 ( \11871 , \11869 , \11870 );
or \U$11619 ( \11872 , \11868 , \11871 );
xor \U$11620 ( \11873 , \6024 , \6035 );
xnor \U$11621 ( \11874 , \11873 , \6014 );
xor \U$11622 ( \11875 , \11872 , \11874 );
xor \U$11623 ( \11876 , \11860 , \11875 );
xor \U$11624 ( \11877 , \11843 , \11876 );
xor \U$11625 ( \11878 , \11802 , \11877 );
xor \U$11626 ( \11879 , \11704 , \11708 );
and \U$11627 ( \11880 , \11879 , \11713 );
and \U$11628 ( \11881 , \11704 , \11708 );
or \U$11629 ( \11882 , \11880 , \11881 );
xor \U$11630 ( \11883 , \11481 , \11497 );
and \U$11631 ( \11884 , \11883 , \11601 );
and \U$11632 ( \11885 , \11481 , \11497 );
or \U$11633 ( \11886 , \11884 , \11885 );
xor \U$11634 ( \11887 , \11882 , \11886 );
xor \U$11635 ( \11888 , \11609 , \11610 );
and \U$11636 ( \11889 , \11888 , \11689 );
and \U$11637 ( \11890 , \11609 , \11610 );
or \U$11638 ( \11891 , \11889 , \11890 );
xor \U$11639 ( \11892 , \11887 , \11891 );
xor \U$11640 ( \11893 , \11878 , \11892 );
xor \U$11641 ( \11894 , \11788 , \11893 );
xnor \U$11642 ( \11895 , \11782 , \11894 );
not \U$11643 ( \11896 , \11895 );
not \U$11644 ( \11897 , \11896 );
xor \U$11645 ( \11898 , \11439 , \11728 );
and \U$11646 ( \11899 , \11898 , \11733 );
and \U$11647 ( \11900 , \11439 , \11728 );
or \U$11648 ( \11901 , \11899 , \11900 );
not \U$11649 ( \11902 , \11901 );
or \U$11650 ( \11903 , \11897 , \11902 );
not \U$11651 ( \11904 , \11901 );
nand \U$11652 ( \11905 , \11904 , \11895 );
nand \U$11653 ( \11906 , \11903 , \11905 );
not \U$11654 ( \11907 , \11775 );
not \U$11655 ( \11908 , \11781 );
or \U$11656 ( \11909 , \11907 , \11908 );
or \U$11657 ( \11910 , \11781 , \11775 );
nand \U$11658 ( \11911 , \11910 , \11894 );
nand \U$11659 ( \11912 , \11909 , \11911 );
not \U$11660 ( \11913 , \11912 );
xor \U$11661 ( \11914 , \11882 , \11886 );
and \U$11662 ( \11915 , \11914 , \11891 );
and \U$11663 ( \11916 , \11882 , \11886 );
or \U$11664 ( \11917 , \11915 , \11916 );
xor \U$11665 ( \11918 , \11820 , \11842 );
and \U$11666 ( \11919 , \11918 , \11876 );
and \U$11667 ( \11920 , \11820 , \11842 );
or \U$11668 ( \11921 , \11919 , \11920 );
xor \U$11669 ( \11922 , \11917 , \11921 );
not \U$11670 ( \11923 , \11841 );
not \U$11671 ( \11924 , \11831 );
or \U$11672 ( \11925 , \11923 , \11924 );
or \U$11673 ( \11926 , \11831 , \11841 );
not \U$11674 ( \11927 , \11824 );
nand \U$11675 ( \11928 , \11926 , \11927 );
nand \U$11676 ( \11929 , \11925 , \11928 );
xor \U$11677 ( \11930 , \11848 , \11929 );
xor \U$11678 ( \11931 , \11808 , \11812 );
and \U$11679 ( \11932 , \11931 , \11819 );
and \U$11680 ( \11933 , \11808 , \11812 );
or \U$11681 ( \11934 , \11932 , \11933 );
xor \U$11682 ( \11935 , \11930 , \11934 );
and \U$11683 ( \11936 , \6073 , \6076 );
not \U$11684 ( \11937 , \6073 );
and \U$11685 ( \11938 , \11937 , \6004 );
nor \U$11686 ( \11939 , \11936 , \11938 );
and \U$11687 ( \11940 , \11939 , \6075 );
not \U$11688 ( \11941 , \11939 );
and \U$11689 ( \11942 , \11941 , \6038 );
nor \U$11690 ( \11943 , \11940 , \11942 );
not \U$11691 ( \11944 , \6110 );
not \U$11692 ( \11945 , \6178 );
or \U$11693 ( \11946 , \11944 , \11945 );
or \U$11694 ( \11947 , \6178 , \6110 );
nand \U$11695 ( \11948 , \11946 , \11947 );
and \U$11696 ( \11949 , \11948 , \6181 );
not \U$11697 ( \11950 , \11948 );
and \U$11698 ( \11951 , \11950 , \6149 );
nor \U$11699 ( \11952 , \11949 , \11951 );
xor \U$11700 ( \11953 , \11943 , \11952 );
not \U$11701 ( \11954 , \5969 );
xor \U$11702 ( \11955 , \5961 , \5956 );
xnor \U$11703 ( \11956 , \11955 , \5955 );
not \U$11704 ( \11957 , \11956 );
or \U$11705 ( \11958 , \11954 , \11957 );
or \U$11706 ( \11959 , \11956 , \5969 );
nand \U$11707 ( \11960 , \11958 , \11959 );
xor \U$11708 ( \11961 , \11953 , \11960 );
xor \U$11709 ( \11962 , \11935 , \11961 );
not \U$11710 ( \11963 , \5737 );
and \U$11711 ( \11964 , \5758 , \10972 );
not \U$11712 ( \11965 , \5758 );
and \U$11713 ( \11966 , \11965 , \5741 );
nor \U$11714 ( \11967 , \11964 , \11966 );
not \U$11715 ( \11968 , \11967 );
or \U$11716 ( \11969 , \11963 , \11968 );
or \U$11717 ( \11970 , \11967 , \5737 );
nand \U$11718 ( \11971 , \11969 , \11970 );
not \U$11719 ( \11972 , \11874 );
not \U$11720 ( \11973 , \11870 );
or \U$11721 ( \11974 , \11972 , \11973 );
or \U$11722 ( \11975 , \11874 , \11870 );
nand \U$11723 ( \11976 , \11975 , \11862 );
nand \U$11724 ( \11977 , \11974 , \11976 );
xor \U$11725 ( \11978 , \11971 , \11977 );
not \U$11726 ( \11979 , \6203 );
not \U$11727 ( \11980 , \6225 );
or \U$11728 ( \11981 , \11979 , \11980 );
or \U$11729 ( \11982 , \6225 , \6203 );
nand \U$11730 ( \11983 , \11981 , \11982 );
and \U$11731 ( \11984 , \11983 , \6214 );
not \U$11732 ( \11985 , \11983 );
and \U$11733 ( \11986 , \11985 , \6213 );
nor \U$11734 ( \11987 , \11984 , \11986 );
xor \U$11735 ( \11988 , \11978 , \11987 );
xor \U$11736 ( \11989 , \11962 , \11988 );
xor \U$11737 ( \11990 , \11922 , \11989 );
xor \U$11738 ( \11991 , \11783 , \11787 );
and \U$11739 ( \11992 , \11991 , \11893 );
and \U$11740 ( \11993 , \11783 , \11787 );
or \U$11741 ( \11994 , \11992 , \11993 );
xor \U$11742 ( \11995 , \11990 , \11994 );
xor \U$11743 ( \11996 , \11792 , \11796 );
and \U$11744 ( \11997 , \11996 , \11801 );
and \U$11745 ( \11998 , \11792 , \11796 );
or \U$11746 ( \11999 , \11997 , \11998 );
xor \U$11747 ( \12000 , \11752 , \11759 );
and \U$11748 ( \12001 , \12000 , \11764 );
and \U$11749 ( \12002 , \11752 , \11759 );
or \U$11750 ( \12003 , \12001 , \12002 );
xor \U$11751 ( \12004 , \11999 , \12003 );
xor \U$11752 ( \12005 , \11849 , \11859 );
and \U$11753 ( \12006 , \12005 , \11875 );
and \U$11754 ( \12007 , \11849 , \11859 );
or \U$11755 ( \12008 , \12006 , \12007 );
xor \U$11756 ( \12009 , \12004 , \12008 );
xor \U$11757 ( \12010 , \11765 , \11769 );
and \U$11758 ( \12011 , \12010 , \11774 );
and \U$11759 ( \12012 , \11765 , \11769 );
or \U$11760 ( \12013 , \12011 , \12012 );
xor \U$11761 ( \12014 , \12009 , \12013 );
xor \U$11762 ( \12015 , \11802 , \11877 );
and \U$11763 ( \12016 , \12015 , \11892 );
and \U$11764 ( \12017 , \11802 , \11877 );
or \U$11765 ( \12018 , \12016 , \12017 );
xor \U$11766 ( \12019 , \12014 , \12018 );
xor \U$11767 ( \12020 , \11995 , \12019 );
not \U$11768 ( \12021 , \12020 );
not \U$11769 ( \12022 , \12021 );
or \U$11770 ( \12023 , \11913 , \12022 );
not \U$11771 ( \12024 , \11912 );
nand \U$11772 ( \12025 , \12024 , \12020 );
nand \U$11773 ( \12026 , \12023 , \12025 );
and \U$11774 ( \12027 , \11739 , \11746 , \11906 , \12026 );
xor \U$11775 ( \12028 , \10594 , \11082 );
xor \U$11776 ( \12029 , \12028 , \11085 );
not \U$11777 ( \12030 , \12029 );
not \U$11778 ( \12031 , \10150 );
not \U$11779 ( \12032 , \10157 );
or \U$11780 ( \12033 , \12031 , \12032 );
or \U$11781 ( \12034 , \10157 , \10150 );
nand \U$11782 ( \12035 , \12033 , \12034 );
xor \U$11783 ( \12036 , \12035 , \9769 );
xor \U$11784 ( \12037 , \11018 , \11029 );
xor \U$11785 ( \12038 , \12037 , \11040 );
not \U$11786 ( \12039 , \12038 );
xor \U$11787 ( \12040 , \10702 , \10729 );
xor \U$11788 ( \12041 , \12040 , \10754 );
not \U$11789 ( \12042 , \10823 );
not \U$11790 ( \12043 , \10867 );
not \U$11791 ( \12044 , \10864 );
not \U$11792 ( \12045 , \12044 );
or \U$11793 ( \12046 , \12043 , \12045 );
nand \U$11794 ( \12047 , \10864 , \10791 );
nand \U$11795 ( \12048 , \12046 , \12047 );
not \U$11796 ( \12049 , \12048 );
or \U$11797 ( \12050 , \12042 , \12049 );
or \U$11798 ( \12051 , \12048 , \10823 );
nand \U$11799 ( \12052 , \12050 , \12051 );
xor \U$11800 ( \12053 , \12041 , \12052 );
not \U$11801 ( \12054 , \10961 );
not \U$11802 ( \12055 , \10910 );
not \U$11803 ( \12056 , \11000 );
or \U$11804 ( \12057 , \12055 , \12056 );
or \U$11805 ( \12058 , \11000 , \10910 );
nand \U$11806 ( \12059 , \12057 , \12058 );
not \U$11807 ( \12060 , \12059 );
or \U$11808 ( \12061 , \12054 , \12060 );
or \U$11809 ( \12062 , \12059 , \10961 );
nand \U$11810 ( \12063 , \12061 , \12062 );
and \U$11811 ( \12064 , \12053 , \12063 );
and \U$11812 ( \12065 , \12041 , \12052 );
or \U$11813 ( \12066 , \12064 , \12065 );
not \U$11814 ( \12067 , \12066 );
nand \U$11815 ( \12068 , \12039 , \12067 );
xor \U$11816 ( \12069 , \10606 , \10608 );
xor \U$11817 ( \12070 , \12069 , \10614 );
and \U$11818 ( \12071 , \12068 , \12070 );
nor \U$11819 ( \12072 , \12039 , \12067 );
nor \U$11820 ( \12073 , \12071 , \12072 );
xor \U$11821 ( \12074 , \10667 , \10689 );
buf \U$11822 ( \12075 , \10652 );
and \U$11823 ( \12076 , \12074 , \12075 );
not \U$11824 ( \12077 , \12074 );
not \U$11825 ( \12078 , \12075 );
and \U$11826 ( \12079 , \12077 , \12078 );
nor \U$11827 ( \12080 , \12076 , \12079 );
not \U$11828 ( \12081 , \12080 );
not \U$11829 ( \12082 , \10757 );
not \U$11830 ( \12083 , \12082 );
xor \U$11831 ( \12084 , \11005 , \10869 );
not \U$11832 ( \12085 , \12084 );
or \U$11833 ( \12086 , \12083 , \12085 );
or \U$11834 ( \12087 , \12084 , \12082 );
nand \U$11835 ( \12088 , \12086 , \12087 );
nand \U$11836 ( \12089 , \12081 , \12088 );
not \U$11837 ( \12090 , \12089 );
and \U$11838 ( \12091 , \2555 , RIbe27f58_10);
and \U$11839 ( \12092 , \6383 , RIbe27e68_8);
nor \U$11840 ( \12093 , \12091 , \12092 );
and \U$11841 ( \12094 , \12093 , \6831 );
not \U$11842 ( \12095 , \12093 );
and \U$11843 ( \12096 , \12095 , \1131 );
nor \U$11844 ( \12097 , \12094 , \12096 );
not \U$11845 ( \12098 , \12097 );
not \U$11846 ( \12099 , RIbe28ed0_43);
not \U$11847 ( \12100 , \1633 );
or \U$11848 ( \12101 , \12099 , \12100 );
nand \U$11849 ( \12102 , \4730 , RIbe27fd0_11);
nand \U$11850 ( \12103 , \12101 , \12102 );
and \U$11851 ( \12104 , \12103 , \5125 );
not \U$11852 ( \12105 , \12103 );
and \U$11853 ( \12106 , \12105 , \1309 );
nor \U$11854 ( \12107 , \12104 , \12106 );
nand \U$11855 ( \12108 , \12098 , \12107 );
and \U$11856 ( \12109 , \1272 , RIbe28660_25);
not \U$11857 ( \12110 , RIbe285e8_24);
nor \U$11858 ( \12111 , \12110 , \2385 );
nor \U$11859 ( \12112 , \12109 , \12111 );
and \U$11860 ( \12113 , \12112 , \1277 );
not \U$11861 ( \12114 , \12112 );
and \U$11862 ( \12115 , \12114 , \3516 );
nor \U$11863 ( \12116 , \12113 , \12115 );
not \U$11864 ( \12117 , \12116 );
and \U$11865 ( \12118 , \12108 , \12117 );
nor \U$11866 ( \12119 , \12098 , \12107 );
nor \U$11867 ( \12120 , \12118 , \12119 );
not \U$11868 ( \12121 , \12120 );
not \U$11869 ( \12122 , \4592 );
not \U$11870 ( \12123 , RIbe289a8_32);
not \U$11871 ( \12124 , \5727 );
or \U$11872 ( \12125 , \12123 , \12124 );
nand \U$11873 ( \12126 , \5731 , RIbe28930_31);
nand \U$11874 ( \12127 , \12125 , \12126 );
not \U$11875 ( \12128 , \12127 );
or \U$11876 ( \12129 , \12122 , \12128 );
or \U$11877 ( \12130 , \12127 , \4946 );
nand \U$11878 ( \12131 , \12129 , \12130 );
not \U$11879 ( \12132 , RIbe29290_51);
not \U$11880 ( \12133 , \6414 );
or \U$11881 ( \12134 , \12132 , \12133 );
nand \U$11882 ( \12135 , \4600 , RIbe28a20_33);
nand \U$11883 ( \12136 , \12134 , \12135 );
and \U$11884 ( \12137 , \12136 , \4326 );
not \U$11885 ( \12138 , \12136 );
and \U$11886 ( \12139 , \12138 , \7865 );
nor \U$11887 ( \12140 , \12137 , \12139 );
xor \U$11888 ( \12141 , \12131 , \12140 );
not \U$11889 ( \12142 , RIbe29560_57);
not \U$11890 ( \12143 , \5455 );
or \U$11891 ( \12144 , \12142 , \12143 );
nand \U$11892 ( \12145 , \6634 , RIbe28228_16);
nand \U$11893 ( \12146 , \12144 , \12145 );
xnor \U$11894 ( \12147 , \12146 , \8252 );
and \U$11895 ( \12148 , \12141 , \12147 );
and \U$11896 ( \12149 , \12131 , \12140 );
or \U$11897 ( \12150 , \12148 , \12149 );
not \U$11898 ( \12151 , \12150 );
not \U$11899 ( \12152 , \12151 );
or \U$11900 ( \12153 , \12121 , \12152 );
not \U$11901 ( \12154 , RIbe28408_20);
not \U$11902 ( \12155 , \3284 );
or \U$11903 ( \12156 , \12154 , \12155 );
nand \U$11904 ( \12157 , \3457 , RIbe28390_19);
nand \U$11905 ( \12158 , \12156 , \12157 );
and \U$11906 ( \12159 , \12158 , \3290 );
not \U$11907 ( \12160 , \12158 );
and \U$11908 ( \12161 , \12160 , \2887 );
or \U$11909 ( \12162 , \12159 , \12161 );
not \U$11910 ( \12163 , \12162 );
not \U$11911 ( \12164 , RIbe287c8_28);
not \U$11912 ( \12165 , \2898 );
or \U$11913 ( \12166 , \12164 , \12165 );
nand \U$11914 ( \12167 , \2901 , RIbe28480_21);
nand \U$11915 ( \12168 , \12166 , \12167 );
and \U$11916 ( \12169 , \12168 , \2379 );
not \U$11917 ( \12170 , \12168 );
and \U$11918 ( \12171 , \12170 , \4287 );
nor \U$11919 ( \12172 , \12169 , \12171 );
not \U$11920 ( \12173 , \12172 );
or \U$11921 ( \12174 , \12163 , \12173 );
not \U$11922 ( \12175 , RIbe28b10_35);
not \U$11923 ( \12176 , \4021 );
or \U$11924 ( \12177 , \12175 , \12176 );
nand \U$11925 ( \12178 , \4332 , RIbe28b88_36);
nand \U$11926 ( \12179 , \12177 , \12178 );
and \U$11927 ( \12180 , \12179 , \3471 );
not \U$11928 ( \12181 , \12179 );
and \U$11929 ( \12182 , \12181 , \3448 );
nor \U$11930 ( \12183 , \12180 , \12182 );
nand \U$11931 ( \12184 , \12174 , \12183 );
or \U$11932 ( \12185 , \12162 , \12172 );
nand \U$11933 ( \12186 , \12184 , \12185 );
nand \U$11934 ( \12187 , \12153 , \12186 );
not \U$11935 ( \12188 , \12120 );
nand \U$11936 ( \12189 , \12188 , \12150 );
nand \U$11937 ( \12190 , \12187 , \12189 );
not \U$11938 ( \12191 , \12190 );
and \U$11939 ( \12192 , RIbe2ad48_108, RIbe2b540_125);
not \U$11940 ( \12193 , RIbe2adc0_109);
nor \U$11941 ( \12194 , \12192 , \12193 );
buf \U$11942 ( \12195 , \12194 );
not \U$11943 ( \12196 , RIbe28e58_42);
not \U$11944 ( \12197 , \10916 );
or \U$11945 ( \12198 , \12196 , \12197 );
nand \U$11946 ( \12199 , \10921 , RIbe28de0_41);
nand \U$11947 ( \12200 , \12198 , \12199 );
not \U$11948 ( \12201 , \12200 );
not \U$11949 ( \12202 , \7970 );
not \U$11950 ( \12203 , \12202 );
and \U$11951 ( \12204 , \12201 , \12203 );
and \U$11952 ( \12205 , \12200 , \10927 );
nor \U$11953 ( \12206 , \12204 , \12205 );
xor \U$11954 ( \12207 , \12195 , \12206 );
not \U$11955 ( \12208 , RIbe29920_65);
not \U$11956 ( \12209 , \10936 );
or \U$11957 ( \12210 , \12208 , \12209 );
xor \U$11958 ( \12211 , RIbe2a460_89, RIbe2adc0_109);
buf \U$11959 ( \12212 , \12211 );
buf \U$11960 ( \12213 , \12212 );
nand \U$11961 ( \12214 , \12213 , RIbe27b98_2);
nand \U$11962 ( \12215 , \12210 , \12214 );
and \U$11963 ( \12216 , \12215 , \9902 );
not \U$11964 ( \12217 , \12215 );
not \U$11965 ( \12218 , \9902 );
buf \U$11966 ( \12219 , \12218 );
and \U$11967 ( \12220 , \12217 , \12219 );
or \U$11968 ( \12221 , \12216 , \12220 );
and \U$11969 ( \12222 , \12207 , \12221 );
and \U$11970 ( \12223 , \12195 , \12206 );
or \U$11971 ( \12224 , \12222 , \12223 );
not \U$11972 ( \12225 , \12224 );
not \U$11973 ( \12226 , \12225 );
not \U$11974 ( \12227 , RIbe27d00_5);
not \U$11975 ( \12228 , \10949 );
or \U$11976 ( \12229 , \12227 , \12228 );
nand \U$11977 ( \12230 , \9891 , RIbe27c10_3);
nand \U$11978 ( \12231 , \12229 , \12230 );
and \U$11979 ( \12232 , \12231 , \6949 );
not \U$11980 ( \12233 , \12231 );
not \U$11981 ( \12234 , \7984 );
and \U$11982 ( \12235 , \12233 , \12234 );
nor \U$11983 ( \12236 , \12232 , \12235 );
not \U$11984 ( \12237 , RIbe28fc0_45);
not \U$11985 ( \12238 , \6561 );
or \U$11986 ( \12239 , \12237 , \12238 );
nand \U$11987 ( \12240 , \7958 , RIbe290b0_47);
nand \U$11988 ( \12241 , \12239 , \12240 );
and \U$11989 ( \12242 , \12241 , \6572 );
not \U$11990 ( \12243 , \12241 );
and \U$11991 ( \12244 , \12243 , \7293 );
nor \U$11992 ( \12245 , \12242 , \12244 );
nand \U$11993 ( \12246 , \12236 , \12245 );
not \U$11994 ( \12247 , \7661 );
not \U$11995 ( \12248 , RIbe29a88_68);
not \U$11996 ( \12249 , \6980 );
or \U$11997 ( \12250 , \12248 , \12249 );
buf \U$11998 ( \12251 , \10898 );
nand \U$11999 ( \12252 , \12251 , RIbe27d78_6);
nand \U$12000 ( \12253 , \12250 , \12252 );
not \U$12001 ( \12254 , \12253 );
or \U$12002 ( \12255 , \12247 , \12254 );
or \U$12003 ( \12256 , \12253 , \6992 );
nand \U$12004 ( \12257 , \12255 , \12256 );
and \U$12005 ( \12258 , \12246 , \12257 );
nor \U$12006 ( \12259 , \12236 , \12245 );
nor \U$12007 ( \12260 , \12258 , \12259 );
not \U$12008 ( \12261 , \12260 );
not \U$12009 ( \12262 , \12261 );
or \U$12010 ( \12263 , \12226 , \12262 );
not \U$12011 ( \12264 , \12260 );
not \U$12012 ( \12265 , \12224 );
or \U$12013 ( \12266 , \12264 , \12265 );
not \U$12014 ( \12267 , RIbe281b0_15);
not \U$12015 ( \12268 , \6855 );
not \U$12016 ( \12269 , \12268 );
or \U$12017 ( \12270 , \12267 , \12269 );
nand \U$12018 ( \12271 , \7528 , RIbe280c0_13);
nand \U$12019 ( \12272 , \12270 , \12271 );
not \U$12020 ( \12273 , \12272 );
not \U$12021 ( \12274 , \7535 );
and \U$12022 ( \12275 , \12273 , \12274 );
and \U$12023 ( \12276 , \12272 , \6141 );
nor \U$12024 ( \12277 , \12275 , \12276 );
not \U$12025 ( \12278 , \12277 );
not \U$12026 ( \12279 , RIbe29650_59);
not \U$12027 ( \12280 , \6592 );
or \U$12028 ( \12281 , \12279 , \12280 );
nand \U$12029 ( \12282 , \7278 , RIbe29038_46);
nand \U$12030 ( \12283 , \12281 , \12282 );
not \U$12031 ( \12284 , \12283 );
not \U$12032 ( \12285 , \7488 );
and \U$12033 ( \12286 , \12284 , \12285 );
and \U$12034 ( \12287 , \12283 , \7949 );
nor \U$12035 ( \12288 , \12286 , \12287 );
not \U$12036 ( \12289 , \12288 );
or \U$12037 ( \12290 , \12278 , \12289 );
not \U$12038 ( \12291 , \6891 );
not \U$12039 ( \12292 , RIbe29830_63);
not \U$12040 ( \12293 , \6536 );
or \U$12041 ( \12294 , \12292 , \12293 );
nand \U$12042 ( \12295 , \6540 , RIbe296c8_60);
nand \U$12043 ( \12296 , \12294 , \12295 );
not \U$12044 ( \12297 , \12296 );
or \U$12045 ( \12298 , \12291 , \12297 );
or \U$12046 ( \12299 , \12296 , \6891 );
nand \U$12047 ( \12300 , \12298 , \12299 );
nand \U$12048 ( \12301 , \12290 , \12300 );
or \U$12049 ( \12302 , \12288 , \12277 );
nand \U$12050 ( \12303 , \12301 , \12302 );
nand \U$12051 ( \12304 , \12266 , \12303 );
nand \U$12052 ( \12305 , \12263 , \12304 );
not \U$12053 ( \12306 , \12305 );
or \U$12054 ( \12307 , \12191 , \12306 );
or \U$12055 ( \12308 , \12305 , \12190 );
nand \U$12056 ( \12309 , RIbe29380_53, RIbe2a190_83);
not \U$12057 ( \12310 , \12309 );
not \U$12058 ( \12311 , RIbe2a5c8_92);
nor \U$12059 ( \12312 , \322 , \321 );
not \U$12060 ( \12313 , \12312 );
or \U$12061 ( \12314 , \12311 , \12313 );
nand \U$12062 ( \12315 , \329 , RIbe2a550_91);
nand \U$12063 ( \12316 , \12314 , \12315 );
not \U$12064 ( \12317 , \12316 );
not \U$12065 ( \12318 , RIbe28048_12);
not \U$12066 ( \12319 , RIbe27ee0_9);
or \U$12067 ( \12320 , \12318 , \12319 );
nand \U$12068 ( \12321 , \12320 , RIbe29380_53);
not \U$12069 ( \12322 , \12321 );
and \U$12070 ( \12323 , \12317 , \12322 );
and \U$12071 ( \12324 , \12316 , \12321 );
nor \U$12072 ( \12325 , \12323 , \12324 );
not \U$12073 ( \12326 , \12325 );
or \U$12074 ( \12327 , \12310 , \12326 );
and \U$12075 ( \12328 , \261 , RIbe2a988_100);
and \U$12076 ( \12329 , \264 , RIbe2a910_99);
nor \U$12077 ( \12330 , \12328 , \12329 );
and \U$12078 ( \12331 , \12330 , \270 );
not \U$12079 ( \12332 , \12330 );
and \U$12080 ( \12333 , \12332 , \269 );
nor \U$12081 ( \12334 , \12331 , \12333 );
nand \U$12082 ( \12335 , \12327 , \12334 );
or \U$12083 ( \12336 , \12309 , \12325 );
nand \U$12084 ( \12337 , \12335 , \12336 );
and \U$12085 ( \12338 , \546 , RIbe2acd0_107);
and \U$12086 ( \12339 , \552 , RIbe2a028_80);
nor \U$12087 ( \12340 , \12338 , \12339 );
not \U$12088 ( \12341 , \12340 );
not \U$12089 ( \12342 , \425 );
and \U$12090 ( \12343 , \12341 , \12342 );
and \U$12091 ( \12344 , \12340 , \425 );
nor \U$12092 ( \12345 , \12343 , \12344 );
not \U$12093 ( \12346 , \12345 );
not \U$12094 ( \12347 , \12346 );
and \U$12095 ( \12348 , \3895 , RIbe2b5b8_126);
and \U$12096 ( \12349 , \3897 , RIbe2a3e8_88);
nor \U$12097 ( \12350 , \12348 , \12349 );
and \U$12098 ( \12351 , \12350 , \300 );
not \U$12099 ( \12352 , \12350 );
and \U$12100 ( \12353 , \12352 , \293 );
nor \U$12101 ( \12354 , \12351 , \12353 );
not \U$12102 ( \12355 , \12354 );
or \U$12103 ( \12356 , \12347 , \12355 );
or \U$12104 ( \12357 , \12354 , \12346 );
not \U$12105 ( \12358 , RIbe2a370_87);
not \U$12106 ( \12359 , \1223 );
or \U$12107 ( \12360 , \12358 , \12359 );
nand \U$12108 ( \12361 , \429 , RIbe2a2f8_86);
nand \U$12109 ( \12362 , \12360 , \12361 );
and \U$12110 ( \12363 , \12362 , \306 );
not \U$12111 ( \12364 , \12362 );
and \U$12112 ( \12365 , \12364 , \1232 );
nor \U$12113 ( \12366 , \12363 , \12365 );
nand \U$12114 ( \12367 , \12357 , \12366 );
nand \U$12115 ( \12368 , \12356 , \12367 );
xor \U$12116 ( \12369 , \12337 , \12368 );
not \U$12117 ( \12370 , RIbe29bf0_71);
not \U$12118 ( \12371 , \1143 );
or \U$12119 ( \12372 , \12370 , \12371 );
nand \U$12120 ( \12373 , \1147 , RIbe28f48_44);
nand \U$12121 ( \12374 , \12372 , \12373 );
and \U$12122 ( \12375 , \12374 , \1469 );
not \U$12123 ( \12376 , \12374 );
and \U$12124 ( \12377 , \12376 , \1152 );
nor \U$12125 ( \12378 , \12375 , \12377 );
not \U$12126 ( \12379 , \8173 );
not \U$12127 ( \12380 , RIbe29e48_76);
not \U$12128 ( \12381 , \12380 );
and \U$12129 ( \12382 , \12379 , \12381 );
and \U$12130 ( \12383 , \664 , RIbe29fb0_79);
nor \U$12131 ( \12384 , \12382 , \12383 );
and \U$12132 ( \12385 , \12384 , \564 );
not \U$12133 ( \12386 , \12384 );
and \U$12134 ( \12387 , \12386 , \3959 );
nor \U$12135 ( \12388 , \12385 , \12387 );
xor \U$12136 ( \12389 , \12378 , \12388 );
and \U$12137 ( \12390 , \2425 , RIbe29dd0_75);
and \U$12138 ( \12391 , \1203 , RIbe29c68_72);
nor \U$12139 ( \12392 , \12390 , \12391 );
and \U$12140 ( \12393 , \12392 , \752 );
not \U$12141 ( \12394 , \12392 );
and \U$12142 ( \12395 , \12394 , \1011 );
nor \U$12143 ( \12396 , \12393 , \12395 );
and \U$12144 ( \12397 , \12389 , \12396 );
and \U$12145 ( \12398 , \12378 , \12388 );
or \U$12146 ( \12399 , \12397 , \12398 );
and \U$12147 ( \12400 , \12369 , \12399 );
and \U$12148 ( \12401 , \12337 , \12368 );
or \U$12149 ( \12402 , \12400 , \12401 );
nand \U$12150 ( \12403 , \12308 , \12402 );
nand \U$12151 ( \12404 , \12307 , \12403 );
or \U$12152 ( \12405 , \10701 , \10700 );
nand \U$12153 ( \12406 , \12405 , \10702 );
xor \U$12154 ( \12407 , \10709 , \10718 );
xor \U$12155 ( \12408 , \12407 , \10726 );
xor \U$12156 ( \12409 , \12406 , \12408 );
not \U$12157 ( \12410 , \10743 );
not \U$12158 ( \12411 , \12410 );
not \U$12159 ( \12412 , \10736 );
not \U$12160 ( \12413 , \10750 );
or \U$12161 ( \12414 , \12412 , \12413 );
or \U$12162 ( \12415 , \10750 , \10736 );
nand \U$12163 ( \12416 , \12414 , \12415 );
not \U$12164 ( \12417 , \12416 );
or \U$12165 ( \12418 , \12411 , \12417 );
or \U$12166 ( \12419 , \12416 , \12410 );
nand \U$12167 ( \12420 , \12418 , \12419 );
and \U$12168 ( \12421 , \12409 , \12420 );
and \U$12169 ( \12422 , \12406 , \12408 );
or \U$12170 ( \12423 , \12421 , \12422 );
not \U$12171 ( \12424 , \10835 );
not \U$12172 ( \12425 , \10846 );
or \U$12173 ( \12426 , \12424 , \12425 );
or \U$12174 ( \12427 , \10846 , \10835 );
nand \U$12175 ( \12428 , \12426 , \12427 );
xnor \U$12176 ( \12429 , \12428 , \10862 );
not \U$12177 ( \12430 , \12429 );
not \U$12178 ( \12431 , \10810 );
not \U$12179 ( \12432 , \10820 );
or \U$12180 ( \12433 , \12431 , \12432 );
or \U$12181 ( \12434 , \10820 , \10810 );
nand \U$12182 ( \12435 , \12433 , \12434 );
and \U$12183 ( \12436 , \12435 , \10801 );
not \U$12184 ( \12437 , \12435 );
not \U$12185 ( \12438 , \10801 );
and \U$12186 ( \12439 , \12437 , \12438 );
nor \U$12187 ( \12440 , \12436 , \12439 );
not \U$12188 ( \12441 , \12440 );
or \U$12189 ( \12442 , \12430 , \12441 );
not \U$12190 ( \12443 , \10768 );
not \U$12191 ( \12444 , \10788 );
or \U$12192 ( \12445 , \12443 , \12444 );
nand \U$12193 ( \12446 , \10787 , \10767 );
nand \U$12194 ( \12447 , \12445 , \12446 );
xnor \U$12195 ( \12448 , \12447 , \10777 );
nand \U$12196 ( \12449 , \12442 , \12448 );
not \U$12197 ( \12450 , \12429 );
not \U$12198 ( \12451 , \12440 );
nand \U$12199 ( \12452 , \12450 , \12451 );
nand \U$12200 ( \12453 , \12449 , \12452 );
xor \U$12201 ( \12454 , \12423 , \12453 );
not \U$12202 ( \12455 , \10907 );
not \U$12203 ( \12456 , \10882 );
or \U$12204 ( \12457 , \12455 , \12456 );
nand \U$12205 ( \12458 , \10881 , \10906 );
nand \U$12206 ( \12459 , \12457 , \12458 );
buf \U$12207 ( \12460 , \10892 );
xnor \U$12208 ( \12461 , \12459 , \12460 );
xor \U$12209 ( \12462 , \10974 , \10998 );
xor \U$12210 ( \12463 , \12462 , \10986 );
xor \U$12211 ( \12464 , \12461 , \12463 );
xor \U$12212 ( \12465 , \10946 , \10929 );
xor \U$12213 ( \12466 , \12465 , \10958 );
and \U$12214 ( \12467 , \12464 , \12466 );
and \U$12215 ( \12468 , \12461 , \12463 );
or \U$12216 ( \12469 , \12467 , \12468 );
and \U$12217 ( \12470 , \12454 , \12469 );
and \U$12218 ( \12471 , \12423 , \12453 );
or \U$12219 ( \12472 , \12470 , \12471 );
xor \U$12220 ( \12473 , \12404 , \12472 );
xnor \U$12221 ( \12474 , \10658 , \10662 );
and \U$12222 ( \12475 , \12474 , \10655 );
not \U$12223 ( \12476 , \12474 );
and \U$12224 ( \12477 , \12476 , \10665 );
nor \U$12225 ( \12478 , \12475 , \12477 );
not \U$12226 ( \12479 , \12478 );
and \U$12227 ( \12480 , \10649 , \10634 );
not \U$12228 ( \12481 , \10649 );
and \U$12229 ( \12482 , \12481 , \10635 );
or \U$12230 ( \12483 , \12480 , \12482 );
and \U$12231 ( \12484 , \12483 , \10638 );
not \U$12232 ( \12485 , \12483 );
and \U$12233 ( \12486 , \12485 , \10639 );
nor \U$12234 ( \12487 , \12484 , \12486 );
not \U$12235 ( \12488 , \12487 );
or \U$12236 ( \12489 , \12479 , \12488 );
xor \U$12237 ( \12490 , \10676 , \10687 );
xnor \U$12238 ( \12491 , \12490 , \10672 );
not \U$12239 ( \12492 , \12491 );
nand \U$12240 ( \12493 , \12489 , \12492 );
not \U$12241 ( \12494 , \12487 );
not \U$12242 ( \12495 , \12478 );
nand \U$12243 ( \12496 , \12494 , \12495 );
nand \U$12244 ( \12497 , \12493 , \12496 );
and \U$12245 ( \12498 , \12473 , \12497 );
and \U$12246 ( \12499 , \12404 , \12472 );
or \U$12247 ( \12500 , \12498 , \12499 );
nor \U$12248 ( \12501 , \12090 , \12500 );
or \U$12249 ( \12502 , \12073 , \12501 );
not \U$12250 ( \12503 , \12089 );
nand \U$12251 ( \12504 , \12503 , \12500 );
nand \U$12252 ( \12505 , \12502 , \12504 );
not \U$12253 ( \12506 , \12505 );
not \U$12254 ( \12507 , \12506 );
and \U$12255 ( \12508 , \10621 , \10617 );
not \U$12256 ( \12509 , \10621 );
and \U$12257 ( \12510 , \12509 , \10618 );
nor \U$12258 ( \12511 , \12508 , \12510 );
xor \U$12259 ( \12512 , \12511 , \10604 );
not \U$12260 ( \12513 , \10692 );
not \U$12261 ( \12514 , \11008 );
and \U$12262 ( \12515 , \12513 , \12514 );
and \U$12263 ( \12516 , \10692 , \11008 );
nor \U$12264 ( \12517 , \12515 , \12516 );
not \U$12265 ( \12518 , \12517 );
not \U$12266 ( \12519 , \11043 );
and \U$12267 ( \12520 , \12518 , \12519 );
and \U$12268 ( \12521 , \12517 , \11043 );
nor \U$12269 ( \12522 , \12520 , \12521 );
not \U$12270 ( \12523 , \11050 );
not \U$12271 ( \12524 , \11053 );
and \U$12272 ( \12525 , \12523 , \12524 );
and \U$12273 ( \12526 , \11050 , \11053 );
nor \U$12274 ( \12527 , \12525 , \12526 );
nand \U$12275 ( \12528 , \12522 , \12527 );
and \U$12276 ( \12529 , \12512 , \12528 );
nor \U$12277 ( \12530 , \12522 , \12527 );
nor \U$12278 ( \12531 , \12529 , \12530 );
not \U$12279 ( \12532 , \12531 );
or \U$12280 ( \12533 , \12507 , \12532 );
not \U$12281 ( \12534 , \11064 );
xor \U$12282 ( \12535 , \11069 , \12534 );
xnor \U$12283 ( \12536 , \12535 , \11072 );
nand \U$12284 ( \12537 , \12533 , \12536 );
or \U$12285 ( \12538 , \12506 , \12531 );
nand \U$12286 ( \12539 , \12537 , \12538 );
xor \U$12287 ( \12540 , \12036 , \12539 );
nor \U$12288 ( \12541 , \11075 , \11059 );
not \U$12289 ( \12542 , \12541 );
nand \U$12290 ( \12543 , \11075 , \11059 );
nand \U$12291 ( \12544 , \12542 , \12543 );
xor \U$12292 ( \12545 , \12544 , \11079 );
and \U$12293 ( \12546 , \12540 , \12545 );
and \U$12294 ( \12547 , \12036 , \12539 );
or \U$12295 ( \12548 , \12546 , \12547 );
nand \U$12296 ( \12549 , \12030 , \12548 );
not \U$12297 ( \12550 , \12549 );
xor \U$12298 ( \12551 , \10592 , \11088 );
not \U$12299 ( \12552 , \12551 );
or \U$12300 ( \12553 , \12550 , \12552 );
or \U$12301 ( \12554 , \12551 , \12549 );
nand \U$12302 ( \12555 , \12553 , \12554 );
xor \U$12303 ( \12556 , \12009 , \12013 );
and \U$12304 ( \12557 , \12556 , \12018 );
and \U$12305 ( \12558 , \12009 , \12013 );
or \U$12306 ( \12559 , \12557 , \12558 );
xor \U$12307 ( \12560 , \11848 , \11929 );
and \U$12308 ( \12561 , \12560 , \11934 );
and \U$12309 ( \12562 , \11848 , \11929 );
or \U$12310 ( \12563 , \12561 , \12562 );
xor \U$12311 ( \12564 , \11971 , \11977 );
and \U$12312 ( \12565 , \12564 , \11987 );
and \U$12313 ( \12566 , \11971 , \11977 );
or \U$12314 ( \12567 , \12565 , \12566 );
xor \U$12315 ( \12568 , \12563 , \12567 );
xor \U$12316 ( \12569 , \11943 , \11952 );
and \U$12317 ( \12570 , \12569 , \11960 );
and \U$12318 ( \12571 , \11943 , \11952 );
or \U$12319 ( \12572 , \12570 , \12571 );
xor \U$12320 ( \12573 , \12568 , \12572 );
xor \U$12321 ( \12574 , \11917 , \11921 );
and \U$12322 ( \12575 , \12574 , \11989 );
and \U$12323 ( \12576 , \11917 , \11921 );
or \U$12324 ( \12577 , \12575 , \12576 );
xor \U$12325 ( \12578 , \12573 , \12577 );
xor \U$12326 ( \12579 , \11999 , \12003 );
and \U$12327 ( \12580 , \12579 , \12008 );
and \U$12328 ( \12581 , \11999 , \12003 );
or \U$12329 ( \12582 , \12580 , \12581 );
xor \U$12330 ( \12583 , \11935 , \11961 );
and \U$12331 ( \12584 , \12583 , \11988 );
and \U$12332 ( \12585 , \11935 , \11961 );
or \U$12333 ( \12586 , \12584 , \12585 );
xor \U$12334 ( \12587 , \12582 , \12586 );
not \U$12335 ( \12588 , \6191 );
not \U$12336 ( \12589 , \6188 );
not \U$12337 ( \12590 , \6194 );
or \U$12338 ( \12591 , \12589 , \12590 );
or \U$12339 ( \12592 , \6194 , \6188 );
nand \U$12340 ( \12593 , \12591 , \12592 );
not \U$12341 ( \12594 , \12593 );
or \U$12342 ( \12595 , \12588 , \12594 );
or \U$12343 ( \12596 , \12593 , \6191 );
nand \U$12344 ( \12597 , \12595 , \12596 );
xor \U$12345 ( \12598 , \5972 , \6183 );
xor \U$12346 ( \12599 , \12598 , \6078 );
xor \U$12347 ( \12600 , \12597 , \12599 );
xor \U$12348 ( \12601 , \6201 , \6230 );
xor \U$12349 ( \12602 , \12601 , \6239 );
xor \U$12350 ( \12603 , \12600 , \12602 );
xor \U$12351 ( \12604 , \12587 , \12603 );
xor \U$12352 ( \12605 , \12578 , \12604 );
xor \U$12353 ( \12606 , \12559 , \12605 );
xor \U$12354 ( \12607 , \11990 , \11994 );
and \U$12355 ( \12608 , \12607 , \12019 );
and \U$12356 ( \12609 , \11990 , \11994 );
or \U$12357 ( \12610 , \12608 , \12609 );
xor \U$12358 ( \12611 , \12606 , \12610 );
and \U$12359 ( \12612 , \12027 , \12555 , \12611 );
not \U$12360 ( \12613 , \6246 );
not \U$12361 ( \12614 , \6242 );
not \U$12362 ( \12615 , \6186 );
and \U$12363 ( \12616 , \12614 , \12615 );
and \U$12364 ( \12617 , \6186 , \6242 );
nor \U$12365 ( \12618 , \12616 , \12617 );
not \U$12366 ( \12619 , \12618 );
or \U$12367 ( \12620 , \12613 , \12619 );
or \U$12368 ( \12621 , \12618 , \6246 );
nand \U$12369 ( \12622 , \12620 , \12621 );
xor \U$12370 ( \12623 , \12582 , \12586 );
and \U$12371 ( \12624 , \12623 , \12603 );
and \U$12372 ( \12625 , \12582 , \12586 );
or \U$12373 ( \12626 , \12624 , \12625 );
xor \U$12374 ( \12627 , \12622 , \12626 );
xor \U$12375 ( \12628 , \12563 , \12567 );
and \U$12376 ( \12629 , \12628 , \12572 );
and \U$12377 ( \12630 , \12563 , \12567 );
or \U$12378 ( \12631 , \12629 , \12630 );
xor \U$12379 ( \12632 , \6249 , \6251 );
xor \U$12380 ( \12633 , \12632 , \6254 );
xor \U$12381 ( \12634 , \12631 , \12633 );
xor \U$12382 ( \12635 , \12597 , \12599 );
and \U$12383 ( \12636 , \12635 , \12602 );
and \U$12384 ( \12637 , \12597 , \12599 );
or \U$12385 ( \12638 , \12636 , \12637 );
xor \U$12386 ( \12639 , \12634 , \12638 );
xor \U$12387 ( \12640 , \12627 , \12639 );
xor \U$12388 ( \12641 , \12573 , \12577 );
and \U$12389 ( \12642 , \12641 , \12604 );
and \U$12390 ( \12643 , \12573 , \12577 );
or \U$12391 ( \12644 , \12642 , \12643 );
and \U$12392 ( \12645 , \12640 , \12644 );
not \U$12393 ( \12646 , \12640 );
not \U$12394 ( \12647 , \12644 );
and \U$12395 ( \12648 , \12646 , \12647 );
nor \U$12396 ( \12649 , \12645 , \12648 );
and \U$12397 ( \12650 , \12559 , \12605 );
xnor \U$12398 ( \12651 , \12649 , \12650 );
not \U$12399 ( \12652 , \12640 );
nor \U$12400 ( \12653 , \12652 , \12647 );
xor \U$12401 ( \12654 , \5644 , \5864 );
xor \U$12402 ( \12655 , \12654 , \5905 );
xor \U$12403 ( \12656 , \12631 , \12633 );
and \U$12404 ( \12657 , \12656 , \12638 );
and \U$12405 ( \12658 , \12631 , \12633 );
or \U$12406 ( \12659 , \12657 , \12658 );
xor \U$12407 ( \12660 , \12655 , \12659 );
xor \U$12408 ( \12661 , \6248 , \6257 );
xor \U$12409 ( \12662 , \12661 , \6267 );
xor \U$12410 ( \12663 , \12660 , \12662 );
xor \U$12411 ( \12664 , \12622 , \12626 );
and \U$12412 ( \12665 , \12664 , \12639 );
and \U$12413 ( \12666 , \12622 , \12626 );
or \U$12414 ( \12667 , \12665 , \12666 );
xor \U$12415 ( \12668 , \12663 , \12667 );
xnor \U$12416 ( \12669 , \12653 , \12668 );
nor \U$12417 ( \12670 , \12651 , \12669 );
not \U$12418 ( \12671 , \12670 );
and \U$12419 ( \12672 , \12663 , \12667 );
xnor \U$12420 ( \12673 , \6270 , \5943 );
not \U$12421 ( \12674 , \12673 );
not \U$12422 ( \12675 , \5947 );
and \U$12423 ( \12676 , \12674 , \12675 );
and \U$12424 ( \12677 , \12673 , \5947 );
nor \U$12425 ( \12678 , \12676 , \12677 );
not \U$12426 ( \12679 , \12678 );
xor \U$12427 ( \12680 , \12655 , \12659 );
and \U$12428 ( \12681 , \12680 , \12662 );
and \U$12429 ( \12682 , \12655 , \12659 );
or \U$12430 ( \12683 , \12681 , \12682 );
not \U$12431 ( \12684 , \12683 );
or \U$12432 ( \12685 , \12679 , \12684 );
or \U$12433 ( \12686 , \12683 , \12678 );
nand \U$12434 ( \12687 , \12685 , \12686 );
xor \U$12435 ( \12688 , \12672 , \12687 );
not \U$12436 ( \12689 , \12678 );
nand \U$12437 ( \12690 , \12689 , \12683 );
xor \U$12438 ( \12691 , \5941 , \6272 );
not \U$12439 ( \12692 , \12691 );
and \U$12440 ( \12693 , \12690 , \12692 );
not \U$12441 ( \12694 , \12690 );
and \U$12442 ( \12695 , \12694 , \12691 );
nor \U$12443 ( \12696 , \12693 , \12695 );
nand \U$12444 ( \12697 , \12688 , \12696 );
nor \U$12445 ( \12698 , \12671 , \12697 );
and \U$12446 ( \12699 , \11092 , \12612 , \12698 );
not \U$12447 ( \12700 , \12699 );
not \U$12448 ( \12701 , RIbe2acd0_107);
xor \U$12449 ( \12702 , RIbe2a640_93, RIbe2ac58_106);
not \U$12450 ( \12703 , \12702 );
xor \U$12451 ( \12704 , RIbe2a640_93, RIbe2a6b8_94);
nand \U$12452 ( \12705 , \12703 , \12704 );
buf \U$12453 ( \12706 , \12705 );
not \U$12454 ( \12707 , \12706 );
not \U$12455 ( \12708 , \12707 );
or \U$12456 ( \12709 , \12701 , \12708 );
buf \U$12457 ( \12710 , \12702 );
buf \U$12458 ( \12711 , \12710 );
nand \U$12459 ( \12712 , \12711 , RIbe2a028_80);
nand \U$12460 ( \12713 , \12709 , \12712 );
nand \U$12461 ( \12714 , RIbe2a640_93, RIbe2ac58_106);
and \U$12462 ( \12715 , \12714 , RIbe2a6b8_94);
buf \U$12463 ( \12716 , \12715 );
and \U$12464 ( \12717 , \12713 , \12716 );
not \U$12465 ( \12718 , \12713 );
not \U$12466 ( \12719 , RIbe2ac58_106);
not \U$12467 ( \12720 , RIbe2a640_93);
or \U$12468 ( \12721 , \12719 , \12720 );
nand \U$12469 ( \12722 , \12721 , RIbe2a6b8_94);
buf \U$12470 ( \12723 , \12722 );
and \U$12471 ( \12724 , \12718 , \12723 );
nor \U$12472 ( \12725 , \12717 , \12724 );
not \U$12473 ( \12726 , RIbe29fb0_79);
xor \U$12474 ( \12727 , RIbe2abe0_105, RIbe2a7a8_96);
not \U$12475 ( \12728 , \12727 );
xor \U$12476 ( \12729 , RIbe2abe0_105, RIbe2ac58_106);
nand \U$12477 ( \12730 , \12728 , \12729 );
buf \U$12478 ( \12731 , \12730 );
not \U$12479 ( \12732 , \12731 );
not \U$12480 ( \12733 , \12732 );
or \U$12481 ( \12734 , \12726 , \12733 );
buf \U$12482 ( \12735 , \12727 );
nand \U$12483 ( \12736 , \12735 , RIbe29e48_76);
nand \U$12484 ( \12737 , \12734 , \12736 );
not \U$12485 ( \12738 , RIbe2a7a8_96);
not \U$12486 ( \12739 , RIbe2abe0_105);
or \U$12487 ( \12740 , \12738 , \12739 );
nand \U$12488 ( \12741 , \12740 , RIbe2ac58_106);
buf \U$12489 ( \12742 , \12741 );
not \U$12490 ( \12743 , \12742 );
and \U$12491 ( \12744 , \12737 , \12743 );
not \U$12492 ( \12745 , \12737 );
buf \U$12493 ( \12746 , \12741 );
and \U$12494 ( \12747 , \12745 , \12746 );
nor \U$12495 ( \12748 , \12744 , \12747 );
xor \U$12496 ( \12749 , \12725 , \12748 );
xor \U$12497 ( \12750 , RIbe2b4c8_124, RIbe2a6b8_94);
not \U$12498 ( \12751 , \12750 );
buf \U$12499 ( \12752 , \12751 );
buf \U$12500 ( \12753 , \12752 );
not \U$12501 ( \12754 , \12753 );
not \U$12502 ( \12755 , RIbe2a2f8_86);
not \U$12503 ( \12756 , \12755 );
and \U$12504 ( \12757 , \12754 , \12756 );
nand \U$12505 ( \12758 , RIbe2b4c8_124, RIbe2a6b8_94);
or \U$12506 ( \12759 , \12758 , RIbe2b540_125);
nor \U$12507 ( \12760 , RIbe2b4c8_124, RIbe2a6b8_94);
nand \U$12508 ( \12761 , \12760 , RIbe2b540_125);
nand \U$12509 ( \12762 , \12759 , \12761 );
not \U$12510 ( \12763 , \12762 );
not \U$12511 ( \12764 , \12763 );
buf \U$12512 ( \12765 , \12764 );
and \U$12513 ( \12766 , \12765 , RIbe2a370_87);
nor \U$12514 ( \12767 , \12757 , \12766 );
nand \U$12515 ( \12768 , \12758 , RIbe2b540_125);
buf \U$12516 ( \12769 , \12768 );
buf \U$12517 ( \12770 , \12769 );
and \U$12518 ( \12771 , \12767 , \12770 );
not \U$12519 ( \12772 , \12767 );
and \U$12520 ( \12773 , \12758 , RIbe2b540_125);
buf \U$12521 ( \12774 , \12773 );
and \U$12522 ( \12775 , \12772 , \12774 );
nor \U$12523 ( \12776 , \12771 , \12775 );
xnor \U$12524 ( \12777 , \12749 , \12776 );
not \U$12525 ( \12778 , \12777 );
not \U$12526 ( \12779 , RIbe29bf0_71);
and \U$12527 ( \12780 , RIbe2b450_123, RIbe2b3d8_122);
nor \U$12528 ( \12781 , RIbe2b450_123, RIbe2aeb0_111);
nor \U$12529 ( \12782 , \12780 , \12781 );
not \U$12530 ( \12783 , RIbe2b3d8_122);
nand \U$12531 ( \12784 , \12783 , RIbe2aeb0_111);
nand \U$12532 ( \12785 , \12782 , \12784 );
not \U$12533 ( \12786 , \12785 );
buf \U$12534 ( \12787 , \12786 );
not \U$12535 ( \12788 , \12787 );
or \U$12536 ( \12789 , \12779 , \12788 );
and \U$12537 ( \12790 , RIbe2aeb0_111, RIbe2b3d8_122);
not \U$12538 ( \12791 , RIbe2aeb0_111);
and \U$12539 ( \12792 , \12791 , \12783 );
nor \U$12540 ( \12793 , \12790 , \12792 );
buf \U$12541 ( \12794 , \12793 );
nand \U$12542 ( \12795 , \12794 , RIbe28f48_44);
nand \U$12543 ( \12796 , \12789 , \12795 );
not \U$12544 ( \12797 , RIbe2b3d8_122);
not \U$12545 ( \12798 , RIbe2aeb0_111);
or \U$12546 ( \12799 , \12797 , \12798 );
nand \U$12547 ( \12800 , \12799 , RIbe2b450_123);
buf \U$12548 ( \12801 , \12800 );
and \U$12549 ( \12802 , \12796 , \12801 );
not \U$12550 ( \12803 , \12796 );
not \U$12551 ( \12804 , \12800 );
and \U$12552 ( \12805 , \12803 , \12804 );
nor \U$12553 ( \12806 , \12802 , \12805 );
not \U$12554 ( \12807 , RIbe28ed0_43);
not \U$12555 ( \12808 , RIbe2ae38_110);
nand \U$12556 ( \12809 , \12808 , RIbe2aeb0_111);
buf \U$12557 ( \12810 , \12809 );
not \U$12558 ( \12811 , \12810 );
not \U$12559 ( \12812 , \12811 );
or \U$12560 ( \12813 , \12807 , \12812 );
nand \U$12561 ( \12814 , RIbe27fd0_11, RIbe2ae38_110);
nand \U$12562 ( \12815 , \12813 , \12814 );
not \U$12563 ( \12816 , RIbe2aeb0_111);
xor \U$12564 ( \12817 , \12815 , \12816 );
xor \U$12565 ( \12818 , \12806 , \12817 );
not \U$12566 ( \12819 , RIbe2b450_123);
not \U$12567 ( \12820 , RIbe2a730_95);
or \U$12568 ( \12821 , \12819 , \12820 );
nand \U$12569 ( \12822 , \12821 , RIbe2a7a8_96);
buf \U$12570 ( \12823 , \12822 );
not \U$12571 ( \12824 , \12823 );
not \U$12572 ( \12825 , RIbe29dd0_75);
xor \U$12573 ( \12826 , RIbe2a730_95, RIbe2b450_123);
not \U$12574 ( \12827 , \12826 );
xor \U$12575 ( \12828 , RIbe2a730_95, RIbe2a7a8_96);
nand \U$12576 ( \12829 , \12827 , \12828 );
buf \U$12577 ( \12830 , \12829 );
not \U$12578 ( \12831 , \12830 );
not \U$12579 ( \12832 , \12831 );
or \U$12580 ( \12833 , \12825 , \12832 );
buf \U$12581 ( \12834 , \12826 );
buf \U$12582 ( \12835 , \12834 );
nand \U$12583 ( \12836 , \12835 , RIbe29c68_72);
nand \U$12584 ( \12837 , \12833 , \12836 );
not \U$12585 ( \12838 , \12837 );
or \U$12586 ( \12839 , \12824 , \12838 );
or \U$12587 ( \12840 , \12837 , \12823 );
nand \U$12588 ( \12841 , \12839 , \12840 );
xnor \U$12589 ( \12842 , \12818 , \12841 );
not \U$12590 ( \12843 , \12842 );
and \U$12591 ( \12844 , \12778 , \12843 );
not \U$12592 ( \12845 , RIbe2a028_80);
buf \U$12593 ( \12846 , \12731 );
not \U$12594 ( \12847 , \12846 );
not \U$12595 ( \12848 , \12847 );
or \U$12596 ( \12849 , \12845 , \12848 );
nand \U$12597 ( \12850 , \12735 , RIbe29fb0_79);
nand \U$12598 ( \12851 , \12849 , \12850 );
not \U$12599 ( \12852 , \12746 );
and \U$12600 ( \12853 , \12851 , \12852 );
not \U$12601 ( \12854 , \12851 );
and \U$12602 ( \12855 , \12854 , \12746 );
nor \U$12603 ( \12856 , \12853 , \12855 );
not \U$12604 ( \12857 , RIbe29e48_76);
not \U$12605 ( \12858 , \12830 );
not \U$12606 ( \12859 , \12858 );
or \U$12607 ( \12860 , \12857 , \12859 );
nand \U$12608 ( \12861 , RIbe29dd0_75, \12834 );
nand \U$12609 ( \12862 , \12860 , \12861 );
buf \U$12610 ( \12863 , \12822 );
and \U$12611 ( \12864 , \12862 , \12863 );
not \U$12612 ( \12865 , \12862 );
not \U$12613 ( \12866 , \12823 );
and \U$12614 ( \12867 , \12865 , \12866 );
nor \U$12615 ( \12868 , \12864 , \12867 );
xor \U$12616 ( \12869 , \12856 , \12868 );
not \U$12617 ( \12870 , RIbe2a2f8_86);
not \U$12618 ( \12871 , \12706 );
not \U$12619 ( \12872 , \12871 );
or \U$12620 ( \12873 , \12870 , \12872 );
nand \U$12621 ( \12874 , \12711 , RIbe2acd0_107);
nand \U$12622 ( \12875 , \12873 , \12874 );
and \U$12623 ( \12876 , \12875 , \12723 );
not \U$12624 ( \12877 , \12875 );
not \U$12625 ( \12878 , \12715 );
not \U$12626 ( \12879 , \12878 );
and \U$12627 ( \12880 , \12877 , \12879 );
nor \U$12628 ( \12881 , \12876 , \12880 );
xnor \U$12629 ( \12882 , \12869 , \12881 );
not \U$12630 ( \12883 , \12882 );
not \U$12631 ( \12884 , \12883 );
not \U$12632 ( \12885 , RIbe29c68_72);
buf \U$12633 ( \12886 , \12785 );
not \U$12634 ( \12887 , \12886 );
not \U$12635 ( \12888 , \12887 );
or \U$12636 ( \12889 , \12885 , \12888 );
buf \U$12637 ( \12890 , \12794 );
nand \U$12638 ( \12891 , \12890 , RIbe29bf0_71);
nand \U$12639 ( \12892 , \12889 , \12891 );
buf \U$12640 ( \12893 , \12800 );
xnor \U$12641 ( \12894 , \12892 , \12893 );
not \U$12642 ( \12895 , \12894 );
not \U$12643 ( \12896 , RIbe28f48_44);
not \U$12644 ( \12897 , \12811 );
or \U$12645 ( \12898 , \12896 , \12897 );
nand \U$12646 ( \12899 , RIbe28ed0_43, RIbe2ae38_110);
nand \U$12647 ( \12900 , \12898 , \12899 );
xor \U$12648 ( \12901 , \12900 , RIbe2aeb0_111);
and \U$12649 ( \12902 , \12901 , \6118 );
not \U$12650 ( \12903 , \12901 );
and \U$12651 ( \12904 , \12903 , \10272 );
nor \U$12652 ( \12905 , \12902 , \12904 );
not \U$12653 ( \12906 , \12905 );
and \U$12654 ( \12907 , \12895 , \12906 );
and \U$12655 ( \12908 , \12894 , \12905 );
nor \U$12656 ( \12909 , \12907 , \12908 );
not \U$12657 ( \12910 , \12909 );
not \U$12658 ( \12911 , \12910 );
or \U$12659 ( \12912 , \12884 , \12911 );
not \U$12660 ( \12913 , \12909 );
not \U$12661 ( \12914 , \12882 );
or \U$12662 ( \12915 , \12913 , \12914 );
not \U$12663 ( \12916 , \12751 );
not \U$12664 ( \12917 , RIbe2a370_87);
not \U$12665 ( \12918 , \12917 );
and \U$12666 ( \12919 , \12916 , \12918 );
buf \U$12667 ( \12920 , \12762 );
buf \U$12668 ( \12921 , \12920 );
and \U$12669 ( \12922 , \12921 , RIbe2a3e8_88);
nor \U$12670 ( \12923 , \12919 , \12922 );
buf \U$12671 ( \12924 , \12769 );
and \U$12672 ( \12925 , \12923 , \12924 );
not \U$12673 ( \12926 , \12923 );
buf \U$12674 ( \12927 , \12773 );
and \U$12675 ( \12928 , \12926 , \12927 );
nor \U$12676 ( \12929 , \12925 , \12928 );
not \U$12677 ( \12930 , \12929 );
not \U$12678 ( \12931 , \12930 );
not \U$12679 ( \12932 , RIbe2a910_99);
not \U$12680 ( \12933 , RIbe2b540_125);
not \U$12681 ( \12934 , \12933 );
not \U$12682 ( \12935 , RIbe2adc0_109);
nor \U$12683 ( \12936 , \12935 , RIbe2ad48_108);
not \U$12684 ( \12937 , \12936 );
or \U$12685 ( \12938 , \12934 , \12937 );
not \U$12686 ( \12939 , RIbe2adc0_109);
nand \U$12687 ( \12940 , \12939 , RIbe2b540_125, RIbe2ad48_108);
nand \U$12688 ( \12941 , \12938 , \12940 );
buf \U$12689 ( \12942 , \12941 );
buf \U$12690 ( \12943 , \12942 );
not \U$12691 ( \12944 , \12943 );
or \U$12692 ( \12945 , \12932 , \12944 );
xor \U$12693 ( \12946 , RIbe2ad48_108, RIbe2b540_125);
buf \U$12694 ( \12947 , \12946 );
buf \U$12695 ( \12948 , \12947 );
nand \U$12696 ( \12949 , \12948 , RIbe2b5b8_126);
nand \U$12697 ( \12950 , \12945 , \12949 );
not \U$12698 ( \12951 , \12950 );
not \U$12699 ( \12952 , RIbe2b540_125);
not \U$12700 ( \12953 , RIbe2ad48_108);
or \U$12701 ( \12954 , \12952 , \12953 );
nand \U$12702 ( \12955 , \12954 , RIbe2adc0_109);
buf \U$12703 ( \12956 , \12955 );
buf \U$12704 ( \12957 , \12956 );
not \U$12705 ( \12958 , \12957 );
and \U$12706 ( \12959 , \12951 , \12958 );
buf \U$12707 ( \12960 , \12956 );
and \U$12708 ( \12961 , \12950 , \12960 );
nor \U$12709 ( \12962 , \12959 , \12961 );
not \U$12710 ( \12963 , \12962 );
not \U$12711 ( \12964 , \12963 );
or \U$12712 ( \12965 , \12931 , \12964 );
nand \U$12713 ( \12966 , \12962 , \12929 );
nand \U$12714 ( \12967 , \12965 , \12966 );
not \U$12715 ( \12968 , RIbe2a550_91);
not \U$12716 ( \12969 , \10936 );
or \U$12717 ( \12970 , \12968 , \12969 );
buf \U$12718 ( \12971 , \12212 );
nand \U$12719 ( \12972 , \12971 , RIbe2a988_100);
nand \U$12720 ( \12973 , \12970 , \12972 );
not \U$12721 ( \12974 , \12973 );
not \U$12722 ( \12975 , \12219 );
and \U$12723 ( \12976 , \12974 , \12975 );
and \U$12724 ( \12977 , \12973 , \10940 );
nor \U$12725 ( \12978 , \12976 , \12977 );
and \U$12726 ( \12979 , \12967 , \12978 );
not \U$12727 ( \12980 , \12967 );
not \U$12728 ( \12981 , \12978 );
and \U$12729 ( \12982 , \12980 , \12981 );
nor \U$12730 ( \12983 , \12979 , \12982 );
not \U$12731 ( \12984 , \12983 );
nand \U$12732 ( \12985 , \12915 , \12984 );
nand \U$12733 ( \12986 , \12912 , \12985 );
nand \U$12734 ( \12987 , \12777 , \12842 );
and \U$12735 ( \12988 , \12986 , \12987 );
nor \U$12736 ( \12989 , \12844 , \12988 );
not \U$12737 ( \12990 , RIbe29dd0_75);
not \U$12738 ( \12991 , \12787 );
or \U$12739 ( \12992 , \12990 , \12991 );
nand \U$12740 ( \12993 , \12890 , RIbe29c68_72);
nand \U$12741 ( \12994 , \12992 , \12993 );
not \U$12742 ( \12995 , \12893 );
and \U$12743 ( \12996 , \12994 , \12995 );
not \U$12744 ( \12997 , \12994 );
not \U$12745 ( \12998 , \12804 );
and \U$12746 ( \12999 , \12997 , \12998 );
nor \U$12747 ( \13000 , \12996 , \12999 );
not \U$12748 ( \13001 , \13000 );
not \U$12749 ( \13002 , \12809 );
buf \U$12750 ( \13003 , \13002 );
buf \U$12751 ( \13004 , \13003 );
and \U$12752 ( \13005 , \13004 , RIbe29bf0_71);
and \U$12753 ( \13006 , RIbe28f48_44, RIbe2ae38_110);
nor \U$12754 ( \13007 , \13005 , \13006 );
xor \U$12755 ( \13008 , \13007 , RIbe2aeb0_111);
nand \U$12756 ( \13009 , \13001 , \13008 );
not \U$12757 ( \13010 , \12830 );
nand \U$12758 ( \13011 , \13010 , RIbe29fb0_79);
not \U$12759 ( \13012 , \12827 );
nand \U$12760 ( \13013 , \13012 , RIbe29e48_76);
and \U$12761 ( \13014 , \13011 , \13013 );
and \U$12762 ( \13015 , \13014 , \12823 );
not \U$12763 ( \13016 , \13014 );
and \U$12764 ( \13017 , \13016 , \12866 );
nor \U$12765 ( \13018 , \13015 , \13017 );
and \U$12766 ( \13019 , \13009 , \13018 );
nor \U$12767 ( \13020 , \13001 , \13008 );
nor \U$12768 ( \13021 , \13019 , \13020 );
not \U$12769 ( \13022 , \13021 );
not \U$12770 ( \13023 , RIbe2a5c8_92);
buf \U$12771 ( \13024 , \10935 );
not \U$12772 ( \13025 , \13024 );
or \U$12773 ( \13026 , \13023 , \13025 );
nand \U$12774 ( \13027 , \12212 , RIbe2a550_91);
nand \U$12775 ( \13028 , \13026 , \13027 );
not \U$12776 ( \13029 , \13028 );
not \U$12777 ( \13030 , \9902 );
not \U$12778 ( \13031 , \13030 );
and \U$12779 ( \13032 , \13029 , \13031 );
not \U$12780 ( \13033 , \9901 );
and \U$12781 ( \13034 , \13028 , \13033 );
nor \U$12782 ( \13035 , \13032 , \13034 );
not \U$12783 ( \13036 , \8277 );
and \U$12784 ( \13037 , \13036 , RIbe2a208_84);
buf \U$12785 ( \13038 , \9912 );
not \U$12786 ( \13039 , \13038 );
not \U$12787 ( \13040 , \13039 );
and \U$12788 ( \13041 , \13040 , RIbe2a190_83);
nor \U$12789 ( \13042 , \13037 , \13041 );
and \U$12790 ( \13043 , \13042 , \10926 );
not \U$12791 ( \13044 , \13042 );
and \U$12792 ( \13045 , \13044 , \8077 );
nor \U$12793 ( \13046 , \13043 , \13045 );
nand \U$12794 ( \13047 , \13035 , \13046 );
not \U$12795 ( \13048 , \12195 );
buf \U$12796 ( \13049 , \12942 );
and \U$12797 ( \13050 , \13049 , RIbe2a988_100);
and \U$12798 ( \13051 , \12947 , RIbe2a910_99);
nor \U$12799 ( \13052 , \13050 , \13051 );
not \U$12800 ( \13053 , \13052 );
or \U$12801 ( \13054 , \13048 , \13053 );
or \U$12802 ( \13055 , \13052 , \12195 );
nand \U$12803 ( \13056 , \13054 , \13055 );
and \U$12804 ( \13057 , \13047 , \13056 );
nor \U$12805 ( \13058 , \13035 , \13046 );
nor \U$12806 ( \13059 , \13057 , \13058 );
not \U$12807 ( \13060 , \13059 );
or \U$12808 ( \13061 , \13022 , \13060 );
not \U$12809 ( \13062 , RIbe2a370_87);
not \U$12810 ( \13063 , \12706 );
not \U$12811 ( \13064 , \13063 );
or \U$12812 ( \13065 , \13062 , \13064 );
nand \U$12813 ( \13066 , \12711 , RIbe2a2f8_86);
nand \U$12814 ( \13067 , \13065 , \13066 );
not \U$12815 ( \13068 , \12878 );
and \U$12816 ( \13069 , \13067 , \13068 );
not \U$12817 ( \13070 , \13067 );
and \U$12818 ( \13071 , \13070 , \12723 );
nor \U$12819 ( \13072 , \13069 , \13071 );
not \U$12820 ( \13073 , RIbe2acd0_107);
not \U$12821 ( \13074 , \12731 );
not \U$12822 ( \13075 , \13074 );
or \U$12823 ( \13076 , \13073 , \13075 );
buf \U$12824 ( \13077 , \12735 );
nand \U$12825 ( \13078 , \13077 , RIbe2a028_80);
nand \U$12826 ( \13079 , \13076 , \13078 );
and \U$12827 ( \13080 , \13079 , \12852 );
not \U$12828 ( \13081 , \13079 );
and \U$12829 ( \13082 , \13081 , \12746 );
nor \U$12830 ( \13083 , \13080 , \13082 );
xor \U$12831 ( \13084 , \13072 , \13083 );
not \U$12832 ( \13085 , \12750 );
not \U$12833 ( \13086 , \13085 );
not \U$12834 ( \13087 , \13086 );
not \U$12835 ( \13088 , \13087 );
not \U$12836 ( \13089 , RIbe2a3e8_88);
not \U$12837 ( \13090 , \13089 );
and \U$12838 ( \13091 , \13088 , \13090 );
not \U$12839 ( \13092 , \12763 );
and \U$12840 ( \13093 , \13092 , RIbe2b5b8_126);
nor \U$12841 ( \13094 , \13091 , \13093 );
and \U$12842 ( \13095 , \13094 , \12924 );
not \U$12843 ( \13096 , \13094 );
and \U$12844 ( \13097 , \13096 , \12927 );
nor \U$12845 ( \13098 , \13095 , \13097 );
and \U$12846 ( \13099 , \13084 , \13098 );
and \U$12847 ( \13100 , \13072 , \13083 );
or \U$12848 ( \13101 , \13099 , \13100 );
nand \U$12849 ( \13102 , \13061 , \13101 );
or \U$12850 ( \13103 , \13021 , \13059 );
nand \U$12851 ( \13104 , \13102 , \13103 );
not \U$12852 ( \13105 , \13104 );
not \U$12853 ( \13106 , RIbe2b180_117);
not \U$12854 ( \13107 , \6561 );
or \U$12855 ( \13108 , \13106 , \13107 );
not \U$12856 ( \13109 , RIbe2b270_119);
not \U$12857 ( \13110 , \13109 );
nand \U$12858 ( \13111 , \13110 , \7653 );
nand \U$12859 ( \13112 , \13108 , \13111 );
not \U$12860 ( \13113 , \13112 );
not \U$12861 ( \13114 , \6569 );
and \U$12862 ( \13115 , \13113 , \13114 );
and \U$12863 ( \13116 , \13112 , \6569 );
nor \U$12864 ( \13117 , \13115 , \13116 );
not \U$12865 ( \13118 , \13117 );
not \U$12866 ( \13119 , \13118 );
not \U$12867 ( \13120 , RIbe2af28_112);
not \U$12868 ( \13121 , \7274 );
or \U$12869 ( \13122 , \13120 , \13121 );
nand \U$12870 ( \13123 , \7483 , RIbe2b1f8_118);
nand \U$12871 ( \13124 , \13122 , \13123 );
and \U$12872 ( \13125 , \13124 , \8957 );
not \U$12873 ( \13126 , \13124 );
and \U$12874 ( \13127 , \13126 , \6601 );
nor \U$12875 ( \13128 , \13125 , \13127 );
not \U$12876 ( \13129 , \13128 );
or \U$12877 ( \13130 , \13119 , \13129 );
not \U$12878 ( \13131 , \13128 );
nand \U$12879 ( \13132 , \13131 , \13117 );
nand \U$12880 ( \13133 , \13130 , \13132 );
not \U$12881 ( \13134 , \6548 );
not \U$12882 ( \13135 , RIbe2b018_114);
not \U$12883 ( \13136 , \6537 );
or \U$12884 ( \13137 , \13135 , \13136 );
nand \U$12885 ( \13138 , \6540 , RIbe2afa0_113);
nand \U$12886 ( \13139 , \13137 , \13138 );
not \U$12887 ( \13140 , \13139 );
or \U$12888 ( \13141 , \13134 , \13140 );
or \U$12889 ( \13142 , \13139 , \6551 );
nand \U$12890 ( \13143 , \13141 , \13142 );
xor \U$12891 ( \13144 , \13133 , \13143 );
and \U$12892 ( \13145 , \10915 , RIbe2a190_83);
and \U$12893 ( \13146 , \9914 , RIbe2a5c8_92);
nor \U$12894 ( \13147 , \13145 , \13146 );
not \U$12895 ( \13148 , \10912 );
and \U$12896 ( \13149 , \13147 , \13148 );
not \U$12897 ( \13150 , \13147 );
and \U$12898 ( \13151 , \13150 , \8077 );
nor \U$12899 ( \13152 , \13149 , \13151 );
not \U$12900 ( \13153 , RIbe2a280_85);
not \U$12901 ( \13154 , \10949 );
or \U$12902 ( \13155 , \13153 , \13154 );
not \U$12903 ( \13156 , RIbe2a208_84);
not \U$12904 ( \13157 , \13156 );
not \U$12905 ( \13158 , \7980 );
nand \U$12906 ( \13159 , \13157 , \13158 );
nand \U$12907 ( \13160 , \13155 , \13159 );
not \U$12908 ( \13161 , \13160 );
not \U$12909 ( \13162 , \6948 );
and \U$12910 ( \13163 , \13161 , \13162 );
and \U$12911 ( \13164 , \13160 , \7984 );
nor \U$12912 ( \13165 , \13163 , \13164 );
xor \U$12913 ( \13166 , \13152 , \13165 );
not \U$12914 ( \13167 , \6992 );
not \U$12915 ( \13168 , \13167 );
not \U$12916 ( \13169 , \13168 );
not \U$12917 ( \13170 , RIbe2b108_116);
buf \U$12918 ( \13171 , \6980 );
not \U$12919 ( \13172 , \13171 );
or \U$12920 ( \13173 , \13170 , \13172 );
nand \U$12921 ( \13174 , \9875 , RIbe2b090_115);
nand \U$12922 ( \13175 , \13173 , \13174 );
not \U$12923 ( \13176 , \13175 );
or \U$12924 ( \13177 , \13169 , \13176 );
or \U$12925 ( \13178 , \13175 , \6992 );
nand \U$12926 ( \13179 , \13177 , \13178 );
xnor \U$12927 ( \13180 , \13166 , \13179 );
nand \U$12928 ( \13181 , \5751 , RIbe2ab68_104);
and \U$12929 ( \13182 , \13181 , \6117 );
not \U$12930 ( \13183 , \13181 );
and \U$12931 ( \13184 , \13183 , \5046 );
nor \U$12932 ( \13185 , \13182 , \13184 );
nand \U$12933 ( \13186 , \13180 , \13185 );
and \U$12934 ( \13187 , \13144 , \13186 );
nor \U$12935 ( \13188 , \13180 , \13185 );
nor \U$12936 ( \13189 , \13187 , \13188 );
and \U$12937 ( \13190 , \13105 , \13189 );
not \U$12938 ( \13191 , \8231 );
not \U$12939 ( \13192 , RIbe2aaf0_103);
nor \U$12940 ( \13193 , \13191 , \13192 );
and \U$12941 ( \13194 , \6617 , RIbe2b630_127);
nor \U$12942 ( \13195 , \13193 , \13194 );
and \U$12943 ( \13196 , \13195 , \6141 );
not \U$12944 ( \13197 , \13195 );
and \U$12945 ( \13198 , \13197 , \6144 );
nor \U$12946 ( \13199 , \13196 , \13198 );
not \U$12947 ( \13200 , \13199 );
not \U$12948 ( \13201 , \13200 );
not \U$12949 ( \13202 , RIbe2b090_115);
not \U$12950 ( \13203 , \10949 );
or \U$12951 ( \13204 , \13202 , \13203 );
nand \U$12952 ( \13205 , \7981 , RIbe2a280_85);
nand \U$12953 ( \13206 , \13204 , \13205 );
and \U$12954 ( \13207 , \13206 , \7984 );
not \U$12955 ( \13208 , \13206 );
and \U$12956 ( \13209 , \13208 , \7985 );
nor \U$12957 ( \13210 , \13207 , \13209 );
not \U$12958 ( \13211 , RIbe2b1f8_118);
not \U$12959 ( \13212 , \6958 );
or \U$12960 ( \13213 , \13211 , \13212 );
nand \U$12961 ( \13214 , \6963 , RIbe2b180_117);
nand \U$12962 ( \13215 , \13213 , \13214 );
and \U$12963 ( \13216 , \13215 , \6572 );
not \U$12964 ( \13217 , \13215 );
and \U$12965 ( \13218 , \13217 , \7293 );
nor \U$12966 ( \13219 , \13216 , \13218 );
nand \U$12967 ( \13220 , \13210 , \13219 );
not \U$12968 ( \13221 , RIbe2b270_119);
not \U$12969 ( \13222 , \6980 );
or \U$12970 ( \13223 , \13221 , \13222 );
not \U$12971 ( \13224 , \8286 );
nand \U$12972 ( \13225 , \13224 , RIbe2b108_116);
nand \U$12973 ( \13226 , \13223 , \13225 );
not \U$12974 ( \13227 , \7301 );
and \U$12975 ( \13228 , \13226 , \13227 );
not \U$12976 ( \13229 , \13226 );
and \U$12977 ( \13230 , \13229 , \6992 );
nor \U$12978 ( \13231 , \13228 , \13230 );
and \U$12979 ( \13232 , \13220 , \13231 );
nor \U$12980 ( \13233 , \13210 , \13219 );
nor \U$12981 ( \13234 , \13232 , \13233 );
not \U$12982 ( \13235 , \13234 );
or \U$12983 ( \13236 , \13201 , \13235 );
not \U$12984 ( \13237 , RIbe2afa0_113);
not \U$12985 ( \13238 , \6590 );
not \U$12986 ( \13239 , \13238 );
or \U$12987 ( \13240 , \13237 , \13239 );
nand \U$12988 ( \13241 , \6596 , RIbe2af28_112);
nand \U$12989 ( \13242 , \13240 , \13241 );
and \U$12990 ( \13243 , \13242 , \6582 );
not \U$12991 ( \13244 , \13242 );
and \U$12992 ( \13245 , \13244 , \8957 );
nor \U$12993 ( \13246 , \13243 , \13245 );
and \U$12994 ( \13247 , \6536 , RIbe2b630_127);
and \U$12995 ( \13248 , \6884 , RIbe2b018_114);
nor \U$12996 ( \13249 , \13247 , \13248 );
and \U$12997 ( \13250 , \13249 , \6551 );
not \U$12998 ( \13251 , \13249 );
and \U$12999 ( \13252 , \13251 , \6547 );
nor \U$13000 ( \13253 , \13250 , \13252 );
xor \U$13001 ( \13254 , \13246 , \13253 );
not \U$13002 ( \13255 , RIbe2ab68_104);
not \U$13003 ( \13256 , \8231 );
or \U$13004 ( \13257 , \13255 , \13256 );
nand \U$13005 ( \13258 , \7528 , RIbe2aaf0_103);
nand \U$13006 ( \13259 , \13257 , \13258 );
and \U$13007 ( \13260 , \13259 , \6144 );
not \U$13008 ( \13261 , \13259 );
and \U$13009 ( \13262 , \13261 , \5740 );
nor \U$13010 ( \13263 , \13260 , \13262 );
and \U$13011 ( \13264 , \13254 , \13263 );
and \U$13012 ( \13265 , \13246 , \13253 );
or \U$13013 ( \13266 , \13264 , \13265 );
nand \U$13014 ( \13267 , \13236 , \13266 );
not \U$13015 ( \13268 , \13234 );
nand \U$13016 ( \13269 , \13268 , \13199 );
and \U$13017 ( \13270 , \13267 , \13269 );
nor \U$13018 ( \13271 , \13190 , \13270 );
nor \U$13019 ( \13272 , \13105 , \13189 );
nor \U$13020 ( \13273 , \13271 , \13272 );
xor \U$13021 ( \13274 , \12989 , \13273 );
not \U$13022 ( \13275 , \5046 );
not \U$13023 ( \13276 , RIbe2ab68_104);
not \U$13024 ( \13277 , \5455 );
or \U$13025 ( \13278 , \13276 , \13277 );
nand \U$13026 ( \13279 , \7100 , RIbe2aaf0_103);
nand \U$13027 ( \13280 , \13278 , \13279 );
not \U$13028 ( \13281 , \13280 );
or \U$13029 ( \13282 , \13275 , \13281 );
or \U$13030 ( \13283 , \13280 , \6118 );
nand \U$13031 ( \13284 , \13282 , \13283 );
not \U$13032 ( \13285 , \13152 );
not \U$13033 ( \13286 , \13165 );
or \U$13034 ( \13287 , \13285 , \13286 );
nand \U$13035 ( \13288 , \13287 , \13179 );
or \U$13036 ( \13289 , \13152 , \13165 );
nand \U$13037 ( \13290 , \13288 , \13289 );
xor \U$13038 ( \13291 , \13284 , \13290 );
not \U$13039 ( \13292 , \13118 );
not \U$13040 ( \13293 , \13131 );
or \U$13041 ( \13294 , \13292 , \13293 );
not \U$13042 ( \13295 , \13128 );
not \U$13043 ( \13296 , \13117 );
or \U$13044 ( \13297 , \13295 , \13296 );
nand \U$13045 ( \13298 , \13297 , \13143 );
nand \U$13046 ( \13299 , \13294 , \13298 );
xor \U$13047 ( \13300 , \13291 , \13299 );
or \U$13048 ( \13301 , \12901 , \6121 );
and \U$13049 ( \13302 , \12894 , \13301 );
not \U$13050 ( \13303 , \12901 );
nor \U$13051 ( \13304 , \13303 , \10984 );
nor \U$13052 ( \13305 , \13302 , \13304 );
not \U$13053 ( \13306 , \13305 );
nor \U$13054 ( \13307 , \12881 , \12868 );
not \U$13055 ( \13308 , \13307 );
not \U$13056 ( \13309 , \12881 );
not \U$13057 ( \13310 , \12868 );
or \U$13058 ( \13311 , \13309 , \13310 );
buf \U$13059 ( \13312 , \12856 );
nand \U$13060 ( \13313 , \13311 , \13312 );
nand \U$13061 ( \13314 , \13308 , \13313 );
xor \U$13062 ( \13315 , \13306 , \13314 );
not \U$13063 ( \13316 , \12981 );
not \U$13064 ( \13317 , \12929 );
or \U$13065 ( \13318 , \13316 , \13317 );
not \U$13066 ( \13319 , \12930 );
not \U$13067 ( \13320 , \12978 );
or \U$13068 ( \13321 , \13319 , \13320 );
nand \U$13069 ( \13322 , \13321 , \12963 );
nand \U$13070 ( \13323 , \13318 , \13322 );
xor \U$13071 ( \13324 , \13315 , \13323 );
or \U$13072 ( \13325 , \13300 , \13324 );
not \U$13073 ( \13326 , RIbe2b270_119);
not \U$13074 ( \13327 , \6559 );
not \U$13075 ( \13328 , \13327 );
or \U$13076 ( \13329 , \13326 , \13328 );
nand \U$13077 ( \13330 , \8202 , RIbe2b108_116);
nand \U$13078 ( \13331 , \13329 , \13330 );
and \U$13079 ( \13332 , \13331 , \6572 );
not \U$13080 ( \13333 , \13331 );
and \U$13081 ( \13334 , \13333 , \7293 );
nor \U$13082 ( \13335 , \13332 , \13334 );
not \U$13083 ( \13336 , RIbe2a208_84);
not \U$13084 ( \13337 , \6942 );
or \U$13085 ( \13338 , \13336 , \13337 );
not \U$13086 ( \13339 , \7980 );
nand \U$13087 ( \13340 , \13339 , RIbe2a190_83);
nand \U$13088 ( \13341 , \13338 , \13340 );
and \U$13089 ( \13342 , \13341 , \6948 );
not \U$13090 ( \13343 , \13341 );
and \U$13091 ( \13344 , \13343 , \12234 );
nor \U$13092 ( \13345 , \13342 , \13344 );
xor \U$13093 ( \13346 , \13335 , \13345 );
and \U$13094 ( \13347 , RIbe2b090_115, \13171 );
not \U$13095 ( \13348 , RIbe2a280_85);
nor \U$13096 ( \13349 , \13348 , \10897 );
nor \U$13097 ( \13350 , \13347 , \13349 );
and \U$13098 ( \13351 , \13350 , \6992 );
not \U$13099 ( \13352 , \13350 );
not \U$13100 ( \13353 , \10902 );
and \U$13101 ( \13354 , \13352 , \13353 );
nor \U$13102 ( \13355 , \13351 , \13354 );
not \U$13103 ( \13356 , \13355 );
xor \U$13104 ( \13357 , \13346 , \13356 );
not \U$13105 ( \13358 , \12957 );
not \U$13106 ( \13359 , RIbe2b5b8_126);
not \U$13107 ( \13360 , \13049 );
or \U$13108 ( \13361 , \13359 , \13360 );
nand \U$13109 ( \13362 , \12948 , RIbe2a3e8_88);
nand \U$13110 ( \13363 , \13361 , \13362 );
not \U$13111 ( \13364 , \13363 );
or \U$13112 ( \13365 , \13358 , \13364 );
or \U$13113 ( \13366 , \13363 , \12957 );
nand \U$13114 ( \13367 , \13365 , \13366 );
not \U$13115 ( \13368 , RIbe2a988_100);
not \U$13116 ( \13369 , \13024 );
or \U$13117 ( \13370 , \13368 , \13369 );
nand \U$13118 ( \13371 , \12213 , RIbe2a910_99);
nand \U$13119 ( \13372 , \13370 , \13371 );
and \U$13120 ( \13373 , \13372 , \13033 );
not \U$13121 ( \13374 , \13372 );
and \U$13122 ( \13375 , \13374 , \9904 );
nor \U$13123 ( \13376 , \13373 , \13375 );
xor \U$13124 ( \13377 , \13367 , \13376 );
and \U$13125 ( \13378 , \8278 , RIbe2a5c8_92);
not \U$13126 ( \13379 , \10919 );
not \U$13127 ( \13380 , \13379 );
and \U$13128 ( \13381 , \13380 , RIbe2a550_91);
nor \U$13129 ( \13382 , \13378 , \13381 );
not \U$13130 ( \13383 , \7970 );
not \U$13131 ( \13384 , \13383 );
and \U$13132 ( \13385 , \13382 , \13384 );
not \U$13133 ( \13386 , \13382 );
and \U$13134 ( \13387 , \13386 , \8077 );
nor \U$13135 ( \13388 , \13385 , \13387 );
xnor \U$13136 ( \13389 , \13377 , \13388 );
not \U$13137 ( \13390 , \13389 );
and \U$13138 ( \13391 , \13357 , \13390 );
not \U$13139 ( \13392 , \13357 );
and \U$13140 ( \13393 , \13392 , \13389 );
nor \U$13141 ( \13394 , \13391 , \13393 );
not \U$13142 ( \13395 , RIbe2b630_127);
not \U$13143 ( \13396 , \8231 );
or \U$13144 ( \13397 , \13395 , \13396 );
nand \U$13145 ( \13398 , \6859 , RIbe2b018_114);
nand \U$13146 ( \13399 , \13397 , \13398 );
not \U$13147 ( \13400 , \13399 );
not \U$13148 ( \13401 , \10972 );
and \U$13149 ( \13402 , \13400 , \13401 );
and \U$13150 ( \13403 , \13399 , \5740 );
nor \U$13151 ( \13404 , \13402 , \13403 );
not \U$13152 ( \13405 , RIbe2afa0_113);
not \U$13153 ( \13406 , \6536 );
or \U$13154 ( \13407 , \13405 , \13406 );
nand \U$13155 ( \13408 , \7076 , RIbe2af28_112);
nand \U$13156 ( \13409 , \13407 , \13408 );
and \U$13157 ( \13410 , \13409 , \6547 );
not \U$13158 ( \13411 , \13409 );
not \U$13159 ( \13412 , \6546 );
and \U$13160 ( \13413 , \13411 , \13412 );
nor \U$13161 ( \13414 , \13410 , \13413 );
xor \U$13162 ( \13415 , \13404 , \13414 );
not \U$13163 ( \13416 , RIbe2b1f8_118);
not \U$13164 ( \13417 , \7274 );
or \U$13165 ( \13418 , \13416 , \13417 );
nand \U$13166 ( \13419 , \6596 , RIbe2b180_117);
nand \U$13167 ( \13420 , \13418 , \13419 );
and \U$13168 ( \13421 , \13420 , \6583 );
not \U$13169 ( \13422 , \13420 );
and \U$13170 ( \13423 , \13422 , \6601 );
nor \U$13171 ( \13424 , \13421 , \13423 );
xor \U$13172 ( \13425 , \13415 , \13424 );
not \U$13173 ( \13426 , \13425 );
xor \U$13174 ( \13427 , \13394 , \13426 );
and \U$13175 ( \13428 , \13325 , \13427 );
and \U$13176 ( \13429 , \13300 , \13324 );
nor \U$13177 ( \13430 , \13428 , \13429 );
xor \U$13178 ( \13431 , \13274 , \13430 );
not \U$13179 ( \13432 , \13431 );
not \U$13180 ( \13433 , RIbe2b018_114);
not \U$13181 ( \13434 , \7941 );
or \U$13182 ( \13435 , \13433 , \13434 );
buf \U$13183 ( \13436 , \7277 );
nand \U$13184 ( \13437 , \13436 , RIbe2afa0_113);
nand \U$13185 ( \13438 , \13435 , \13437 );
and \U$13186 ( \13439 , \13438 , \9868 );
not \U$13187 ( \13440 , \13438 );
and \U$13188 ( \13441 , \13440 , \6582 );
nor \U$13189 ( \13442 , \13439 , \13441 );
not \U$13190 ( \13443 , \13442 );
not \U$13191 ( \13444 , RIbe2af28_112);
not \U$13192 ( \13445 , \7954 );
or \U$13193 ( \13446 , \13444 , \13445 );
nand \U$13194 ( \13447 , \7958 , RIbe2b1f8_118);
nand \U$13195 ( \13448 , \13446 , \13447 );
and \U$13196 ( \13449 , \13448 , \7293 );
not \U$13197 ( \13450 , \13448 );
and \U$13198 ( \13451 , \13450 , \6572 );
nor \U$13199 ( \13452 , \13449 , \13451 );
or \U$13200 ( \13453 , \13443 , \13452 );
not \U$13201 ( \13454 , RIbe2aaf0_103);
not \U$13202 ( \13455 , \6536 );
or \U$13203 ( \13456 , \13454 , \13455 );
nand \U$13204 ( \13457 , \10348 , RIbe2b630_127);
nand \U$13205 ( \13458 , \13456 , \13457 );
and \U$13206 ( \13459 , \13458 , \7935 );
not \U$13207 ( \13460 , \13458 );
and \U$13208 ( \13461 , \13460 , \6891 );
nor \U$13209 ( \13462 , \13459 , \13461 );
nand \U$13210 ( \13463 , \13453 , \13462 );
nand \U$13211 ( \13464 , \13443 , \13452 );
nand \U$13212 ( \13465 , \13463 , \13464 );
not \U$13213 ( \13466 , RIbe2b108_116);
not \U$13214 ( \13467 , \10949 );
or \U$13215 ( \13468 , \13466 , \13467 );
nand \U$13216 ( \13469 , \9891 , RIbe2b090_115);
nand \U$13217 ( \13470 , \13468 , \13469 );
and \U$13218 ( \13471 , \13470 , \9896 );
not \U$13219 ( \13472 , \13470 );
and \U$13220 ( \13473 , \13472 , \6948 );
nor \U$13221 ( \13474 , \13471 , \13473 );
not \U$13222 ( \13475 , \13474 );
not \U$13223 ( \13476 , RIbe2a280_85);
not \U$13224 ( \13477 , \8276 );
not \U$13225 ( \13478 , \13477 );
not \U$13226 ( \13479 , \13478 );
or \U$13227 ( \13480 , \13476 , \13479 );
nand \U$13228 ( \13481 , \13038 , RIbe2a208_84);
nand \U$13229 ( \13482 , \13480 , \13481 );
not \U$13230 ( \13483 , \13482 );
not \U$13231 ( \13484 , \8077 );
and \U$13232 ( \13485 , \13483 , \13484 );
and \U$13233 ( \13486 , \13482 , \8077 );
nor \U$13234 ( \13487 , \13485 , \13486 );
not \U$13235 ( \13488 , \13487 );
not \U$13236 ( \13489 , \13488 );
or \U$13237 ( \13490 , \13475 , \13489 );
or \U$13238 ( \13491 , \13488 , \13474 );
not \U$13239 ( \13492 , RIbe2b180_117);
not \U$13240 ( \13493 , \6980 );
or \U$13241 ( \13494 , \13492 , \13493 );
nand \U$13242 ( \13495 , \8287 , RIbe2b270_119);
nand \U$13243 ( \13496 , \13494 , \13495 );
and \U$13244 ( \13497 , \13496 , \7304 );
not \U$13245 ( \13498 , \13496 );
and \U$13246 ( \13499 , \13498 , \6992 );
nor \U$13247 ( \13500 , \13497 , \13499 );
nand \U$13248 ( \13501 , \13491 , \13500 );
nand \U$13249 ( \13502 , \13490 , \13501 );
xor \U$13250 ( \13503 , \13465 , \13502 );
xor \U$13251 ( \13504 , \13246 , \13253 );
xor \U$13252 ( \13505 , \13504 , \13263 );
and \U$13253 ( \13506 , \13503 , \13505 );
and \U$13254 ( \13507 , \13465 , \13502 );
or \U$13255 ( \13508 , \13506 , \13507 );
not \U$13256 ( \13509 , RIbe29c68_72);
not \U$13257 ( \13510 , \13004 );
or \U$13258 ( \13511 , \13509 , \13510 );
nand \U$13259 ( \13512 , RIbe29bf0_71, RIbe2ae38_110);
nand \U$13260 ( \13513 , \13511 , \13512 );
xor \U$13261 ( \13514 , \13513 , RIbe2aeb0_111);
xor \U$13262 ( \13515 , \7501 , \13514 );
not \U$13263 ( \13516 , \12801 );
not \U$13264 ( \13517 , RIbe29e48_76);
not \U$13265 ( \13518 , \12886 );
not \U$13266 ( \13519 , \13518 );
or \U$13267 ( \13520 , \13517 , \13519 );
nand \U$13268 ( \13521 , \12890 , RIbe29dd0_75);
nand \U$13269 ( \13522 , \13520 , \13521 );
not \U$13270 ( \13523 , \13522 );
or \U$13271 ( \13524 , \13516 , \13523 );
or \U$13272 ( \13525 , \13522 , \12998 );
nand \U$13273 ( \13526 , \13524 , \13525 );
and \U$13274 ( \13527 , \13515 , \13526 );
and \U$13275 ( \13528 , \7501 , \13514 );
or \U$13276 ( \13529 , \13527 , \13528 );
not \U$13277 ( \13530 , \12752 );
not \U$13278 ( \13531 , RIbe2b5b8_126);
not \U$13279 ( \13532 , \13531 );
and \U$13280 ( \13533 , \13530 , \13532 );
and \U$13281 ( \13534 , \13092 , RIbe2a910_99);
nor \U$13282 ( \13535 , \13533 , \13534 );
and \U$13283 ( \13536 , \13535 , \12770 );
not \U$13284 ( \13537 , \13535 );
and \U$13285 ( \13538 , \13537 , \12927 );
nor \U$13286 ( \13539 , \13536 , \13538 );
not \U$13287 ( \13540 , RIbe2a190_83);
not \U$13288 ( \13541 , \10936 );
or \U$13289 ( \13542 , \13540 , \13541 );
nand \U$13290 ( \13543 , \12971 , RIbe2a5c8_92);
nand \U$13291 ( \13544 , \13542 , \13543 );
and \U$13292 ( \13545 , \13544 , \9904 );
not \U$13293 ( \13546 , \13544 );
and \U$13294 ( \13547 , \13546 , \9903 );
nor \U$13295 ( \13548 , \13545 , \13547 );
xor \U$13296 ( \13549 , \13539 , \13548 );
and \U$13297 ( \13550 , \12943 , RIbe2a550_91);
not \U$13298 ( \13551 , \12948 );
not \U$13299 ( \13552 , RIbe2a988_100);
nor \U$13300 ( \13553 , \13551 , \13552 );
nor \U$13301 ( \13554 , \13550 , \13553 );
and \U$13302 ( \13555 , \13554 , \12956 );
not \U$13303 ( \13556 , \13554 );
and \U$13304 ( \13557 , \13556 , \12195 );
nor \U$13305 ( \13558 , \13555 , \13557 );
and \U$13306 ( \13559 , \13549 , \13558 );
and \U$13307 ( \13560 , \13539 , \13548 );
or \U$13308 ( \13561 , \13559 , \13560 );
xor \U$13309 ( \13562 , \13529 , \13561 );
not \U$13310 ( \13563 , RIbe2a2f8_86);
not \U$13311 ( \13564 , \13074 );
or \U$13312 ( \13565 , \13563 , \13564 );
nand \U$13313 ( \13566 , \12735 , RIbe2acd0_107);
nand \U$13314 ( \13567 , \13565 , \13566 );
and \U$13315 ( \13568 , \13567 , \12746 );
not \U$13316 ( \13569 , \13567 );
not \U$13317 ( \13570 , \12746 );
and \U$13318 ( \13571 , \13569 , \13570 );
nor \U$13319 ( \13572 , \13568 , \13571 );
not \U$13320 ( \13573 , \13572 );
not \U$13321 ( \13574 , \13573 );
not \U$13322 ( \13575 , RIbe2a3e8_88);
not \U$13323 ( \13576 , \13063 );
or \U$13324 ( \13577 , \13575 , \13576 );
nand \U$13325 ( \13578 , \12711 , RIbe2a370_87);
nand \U$13326 ( \13579 , \13577 , \13578 );
and \U$13327 ( \13580 , \13579 , \13068 );
not \U$13328 ( \13581 , \13579 );
not \U$13329 ( \13582 , \12723 );
not \U$13330 ( \13583 , \13582 );
and \U$13331 ( \13584 , \13581 , \13583 );
nor \U$13332 ( \13585 , \13580 , \13584 );
not \U$13333 ( \13586 , \13585 );
or \U$13334 ( \13587 , \13574 , \13586 );
or \U$13335 ( \13588 , \13585 , \13573 );
not \U$13336 ( \13589 , RIbe2a028_80);
not \U$13337 ( \13590 , \12830 );
not \U$13338 ( \13591 , \13590 );
or \U$13339 ( \13592 , \13589 , \13591 );
nand \U$13340 ( \13593 , \12835 , RIbe29fb0_79);
nand \U$13341 ( \13594 , \13592 , \13593 );
not \U$13342 ( \13595 , \12822 );
and \U$13343 ( \13596 , \13594 , \13595 );
not \U$13344 ( \13597 , \13594 );
and \U$13345 ( \13598 , \13597 , \12863 );
nor \U$13346 ( \13599 , \13596 , \13598 );
nand \U$13347 ( \13600 , \13588 , \13599 );
nand \U$13348 ( \13601 , \13587 , \13600 );
and \U$13349 ( \13602 , \13562 , \13601 );
and \U$13350 ( \13603 , \13529 , \13561 );
or \U$13351 ( \13604 , \13602 , \13603 );
xor \U$13352 ( \13605 , \13508 , \13604 );
xor \U$13353 ( \13606 , \13072 , \13083 );
xor \U$13354 ( \13607 , \13606 , \13098 );
xor \U$13355 ( \13608 , \13056 , \13035 );
xor \U$13356 ( \13609 , \13608 , \13046 );
xor \U$13357 ( \13610 , \13607 , \13609 );
xor \U$13358 ( \13611 , \13231 , \13210 );
xor \U$13359 ( \13612 , \13611 , \13219 );
and \U$13360 ( \13613 , \13610 , \13612 );
and \U$13361 ( \13614 , \13607 , \13609 );
or \U$13362 ( \13615 , \13613 , \13614 );
and \U$13363 ( \13616 , \13605 , \13615 );
and \U$13364 ( \13617 , \13508 , \13604 );
or \U$13365 ( \13618 , \13616 , \13617 );
xor \U$13366 ( \13619 , \13199 , \13234 );
xnor \U$13367 ( \13620 , \13619 , \13266 );
xor \U$13368 ( \13621 , \13185 , \13180 );
xor \U$13369 ( \13622 , \13621 , \13144 );
xor \U$13370 ( \13623 , \13620 , \13622 );
and \U$13371 ( \13624 , \12983 , \12883 );
not \U$13372 ( \13625 , \12983 );
and \U$13373 ( \13626 , \13625 , \12882 );
nor \U$13374 ( \13627 , \13624 , \13626 );
and \U$13375 ( \13628 , \13627 , \12909 );
not \U$13376 ( \13629 , \13627 );
and \U$13377 ( \13630 , \13629 , \12910 );
nor \U$13378 ( \13631 , \13628 , \13630 );
and \U$13379 ( \13632 , \13623 , \13631 );
and \U$13380 ( \13633 , \13620 , \13622 );
or \U$13381 ( \13634 , \13632 , \13633 );
xor \U$13382 ( \13635 , \13618 , \13634 );
xor \U$13383 ( \13636 , \13300 , \13324 );
xor \U$13384 ( \13637 , \13636 , \13427 );
xor \U$13385 ( \13638 , \13635 , \13637 );
xor \U$13386 ( \13639 , \13021 , \13059 );
xor \U$13387 ( \13640 , \13639 , \13101 );
and \U$13388 ( \13641 , \13478 , RIbe2b090_115);
not \U$13389 ( \13642 , \9913 );
not \U$13390 ( \13643 , \13642 );
and \U$13391 ( \13644 , \13643 , RIbe2a280_85);
nor \U$13392 ( \13645 , \13641 , \13644 );
not \U$13393 ( \13646 , \12202 );
and \U$13394 ( \13647 , \13645 , \13646 );
not \U$13395 ( \13648 , \13645 );
not \U$13396 ( \13649 , \8077 );
not \U$13397 ( \13650 , \13649 );
and \U$13398 ( \13651 , \13648 , \13650 );
nor \U$13399 ( \13652 , \13647 , \13651 );
not \U$13400 ( \13653 , RIbe2a208_84);
not \U$13401 ( \13654 , \13024 );
or \U$13402 ( \13655 , \13653 , \13654 );
nand \U$13403 ( \13656 , \12212 , RIbe2a190_83);
nand \U$13404 ( \13657 , \13655 , \13656 );
not \U$13405 ( \13658 , \13657 );
not \U$13406 ( \13659 , \12218 );
and \U$13407 ( \13660 , \13658 , \13659 );
not \U$13408 ( \13661 , \9902 );
and \U$13409 ( \13662 , \13657 , \13661 );
nor \U$13410 ( \13663 , \13660 , \13662 );
nand \U$13411 ( \13664 , \13652 , \13663 );
not \U$13412 ( \13665 , \12960 );
not \U$13413 ( \13666 , RIbe2a5c8_92);
not \U$13414 ( \13667 , \12942 );
or \U$13415 ( \13668 , \13666 , \13667 );
buf \U$13416 ( \13669 , \12947 );
nand \U$13417 ( \13670 , \13669 , RIbe2a550_91);
nand \U$13418 ( \13671 , \13668 , \13670 );
not \U$13419 ( \13672 , \13671 );
or \U$13420 ( \13673 , \13665 , \13672 );
or \U$13421 ( \13674 , \13671 , \12960 );
nand \U$13422 ( \13675 , \13673 , \13674 );
and \U$13423 ( \13676 , \13664 , \13675 );
nor \U$13424 ( \13677 , \13663 , \13652 );
nor \U$13425 ( \13678 , \13676 , \13677 );
not \U$13426 ( \13679 , \13678 );
not \U$13427 ( \13680 , RIbe29fb0_79);
not \U$13428 ( \13681 , \13518 );
or \U$13429 ( \13682 , \13680 , \13681 );
nand \U$13430 ( \13683 , \12794 , RIbe29e48_76);
nand \U$13431 ( \13684 , \13682 , \13683 );
and \U$13432 ( \13685 , \13684 , \12801 );
not \U$13433 ( \13686 , \13684 );
and \U$13434 ( \13687 , \13686 , \12995 );
nor \U$13435 ( \13688 , \13685 , \13687 );
not \U$13436 ( \13689 , RIbe29dd0_75);
not \U$13437 ( \13690 , \12810 );
not \U$13438 ( \13691 , \13690 );
or \U$13439 ( \13692 , \13689 , \13691 );
nand \U$13440 ( \13693 , RIbe29c68_72, RIbe2ae38_110);
nand \U$13441 ( \13694 , \13692 , \13693 );
xnor \U$13442 ( \13695 , \13694 , RIbe2aeb0_111);
nand \U$13443 ( \13696 , \13688 , \13695 );
not \U$13444 ( \13697 , \12863 );
not \U$13445 ( \13698 , RIbe2acd0_107);
not \U$13446 ( \13699 , \13590 );
or \U$13447 ( \13700 , \13698 , \13699 );
nand \U$13448 ( \13701 , \13012 , RIbe2a028_80);
nand \U$13449 ( \13702 , \13700 , \13701 );
not \U$13450 ( \13703 , \13702 );
or \U$13451 ( \13704 , \13697 , \13703 );
buf \U$13452 ( \13705 , \13595 );
not \U$13453 ( \13706 , \13705 );
or \U$13454 ( \13707 , \13702 , \13706 );
nand \U$13455 ( \13708 , \13704 , \13707 );
and \U$13456 ( \13709 , \13696 , \13708 );
nor \U$13457 ( \13710 , \13688 , \13695 );
nor \U$13458 ( \13711 , \13709 , \13710 );
not \U$13459 ( \13712 , \13711 );
or \U$13460 ( \13713 , \13679 , \13712 );
not \U$13461 ( \13714 , RIbe2a370_87);
not \U$13462 ( \13715 , \12847 );
or \U$13463 ( \13716 , \13714 , \13715 );
nand \U$13464 ( \13717 , \13077 , RIbe2a2f8_86);
nand \U$13465 ( \13718 , \13716 , \13717 );
and \U$13466 ( \13719 , \13718 , \12746 );
not \U$13467 ( \13720 , \13718 );
and \U$13468 ( \13721 , \13720 , \13570 );
nor \U$13469 ( \13722 , \13719 , \13721 );
not \U$13470 ( \13723 , \13722 );
not \U$13471 ( \13724 , RIbe2b5b8_126);
not \U$13472 ( \13725 , \13063 );
or \U$13473 ( \13726 , \13724 , \13725 );
not \U$13474 ( \13727 , \12703 );
buf \U$13475 ( \13728 , \13727 );
nand \U$13476 ( \13729 , \13728 , RIbe2a3e8_88);
nand \U$13477 ( \13730 , \13726 , \13729 );
and \U$13478 ( \13731 , \13730 , \12723 );
not \U$13479 ( \13732 , \13730 );
and \U$13480 ( \13733 , \13732 , \12716 );
nor \U$13481 ( \13734 , \13731 , \13733 );
not \U$13482 ( \13735 , \13734 );
or \U$13483 ( \13736 , \13723 , \13735 );
not \U$13484 ( \13737 , RIbe2a988_100);
buf \U$13485 ( \13738 , \12920 );
not \U$13486 ( \13739 , \13738 );
or \U$13487 ( \13740 , \13737 , \13739 );
nand \U$13488 ( \13741 , \13086 , RIbe2a910_99);
nand \U$13489 ( \13742 , \13740 , \13741 );
xnor \U$13490 ( \13743 , \13742 , \12924 );
nand \U$13491 ( \13744 , \13736 , \13743 );
not \U$13492 ( \13745 , \13722 );
not \U$13493 ( \13746 , \13734 );
nand \U$13494 ( \13747 , \13745 , \13746 );
nand \U$13495 ( \13748 , \13744 , \13747 );
nand \U$13496 ( \13749 , \13713 , \13748 );
not \U$13497 ( \13750 , \13711 );
not \U$13498 ( \13751 , \13678 );
nand \U$13499 ( \13752 , \13750 , \13751 );
nand \U$13500 ( \13753 , \13749 , \13752 );
nand \U$13501 ( \13754 , \7087 , RIbe2ab68_104);
and \U$13502 ( \13755 , \13754 , \10972 );
not \U$13503 ( \13756 , \13754 );
and \U$13504 ( \13757 , \13756 , \10969 );
nor \U$13505 ( \13758 , \13755 , \13757 );
not \U$13506 ( \13759 , \13758 );
xor \U$13507 ( \13760 , \13452 , \13442 );
xor \U$13508 ( \13761 , \13760 , \13462 );
not \U$13509 ( \13762 , \13761 );
not \U$13510 ( \13763 , \13762 );
or \U$13511 ( \13764 , \13759 , \13763 );
not \U$13512 ( \13765 , \13758 );
nand \U$13513 ( \13766 , \13765 , \13761 );
not \U$13514 ( \13767 , RIbe2afa0_113);
not \U$13515 ( \13768 , \6561 );
or \U$13516 ( \13769 , \13767 , \13768 );
nand \U$13517 ( \13770 , \7958 , RIbe2af28_112);
nand \U$13518 ( \13771 , \13769 , \13770 );
and \U$13519 ( \13772 , \13771 , \7293 );
not \U$13520 ( \13773 , \13771 );
and \U$13521 ( \13774 , \13773 , \6572 );
nor \U$13522 ( \13775 , \13772 , \13774 );
not \U$13523 ( \13776 , \13775 );
not \U$13524 ( \13777 , RIbe2b270_119);
not \U$13525 ( \13778 , \7975 );
or \U$13526 ( \13779 , \13777 , \13778 );
nand \U$13527 ( \13780 , \9891 , RIbe2b108_116);
nand \U$13528 ( \13781 , \13779 , \13780 );
and \U$13529 ( \13782 , \13781 , \8480 );
not \U$13530 ( \13783 , \13781 );
and \U$13531 ( \13784 , \13783 , \6949 );
nor \U$13532 ( \13785 , \13782 , \13784 );
not \U$13533 ( \13786 , \13785 );
or \U$13534 ( \13787 , \13776 , \13786 );
or \U$13535 ( \13788 , \13785 , \13775 );
not \U$13536 ( \13789 , RIbe2b1f8_118);
not \U$13537 ( \13790 , \7298 );
or \U$13538 ( \13791 , \13789 , \13790 );
not \U$13539 ( \13792 , \10897 );
nand \U$13540 ( \13793 , \13792 , RIbe2b180_117);
nand \U$13541 ( \13794 , \13791 , \13793 );
and \U$13542 ( \13795 , \13794 , \13167 );
not \U$13543 ( \13796 , \13794 );
and \U$13544 ( \13797 , \13796 , \7301 );
or \U$13545 ( \13798 , \13795 , \13797 );
not \U$13546 ( \13799 , \13798 );
nand \U$13547 ( \13800 , \13788 , \13799 );
nand \U$13548 ( \13801 , \13787 , \13800 );
nand \U$13549 ( \13802 , \13766 , \13801 );
nand \U$13550 ( \13803 , \13764 , \13802 );
xor \U$13551 ( \13804 , \13753 , \13803 );
and \U$13552 ( \13805 , \13599 , \13572 );
not \U$13553 ( \13806 , \13599 );
and \U$13554 ( \13807 , \13806 , \13573 );
or \U$13555 ( \13808 , \13805 , \13807 );
xnor \U$13556 ( \13809 , \13808 , \13585 );
not \U$13557 ( \13810 , \13809 );
xor \U$13558 ( \13811 , \13474 , \13487 );
xor \U$13559 ( \13812 , \13811 , \13500 );
not \U$13560 ( \13813 , \13812 );
or \U$13561 ( \13814 , \13810 , \13813 );
xor \U$13562 ( \13815 , \13539 , \13548 );
xor \U$13563 ( \13816 , \13815 , \13558 );
nand \U$13564 ( \13817 , \13814 , \13816 );
not \U$13565 ( \13818 , \13809 );
not \U$13566 ( \13819 , \13812 );
nand \U$13567 ( \13820 , \13818 , \13819 );
nand \U$13568 ( \13821 , \13817 , \13820 );
and \U$13569 ( \13822 , \13804 , \13821 );
and \U$13570 ( \13823 , \13753 , \13803 );
or \U$13571 ( \13824 , \13822 , \13823 );
xor \U$13572 ( \13825 , \13640 , \13824 );
xor \U$13573 ( \13826 , \13000 , \13008 );
xnor \U$13574 ( \13827 , \13826 , \13018 );
xor \U$13575 ( \13828 , \13465 , \13502 );
xor \U$13576 ( \13829 , \13828 , \13505 );
xor \U$13577 ( \13830 , \13827 , \13829 );
xor \U$13578 ( \13831 , \13607 , \13609 );
xor \U$13579 ( \13832 , \13831 , \13612 );
and \U$13580 ( \13833 , \13830 , \13832 );
and \U$13581 ( \13834 , \13827 , \13829 );
or \U$13582 ( \13835 , \13833 , \13834 );
and \U$13583 ( \13836 , \13825 , \13835 );
and \U$13584 ( \13837 , \13640 , \13824 );
or \U$13585 ( \13838 , \13836 , \13837 );
xor \U$13586 ( \13839 , \12842 , \12777 );
xor \U$13587 ( \13840 , \13839 , \12986 );
not \U$13588 ( \13841 , \13189 );
and \U$13589 ( \13842 , \13270 , \13105 );
not \U$13590 ( \13843 , \13270 );
and \U$13591 ( \13844 , \13843 , \13104 );
nor \U$13592 ( \13845 , \13842 , \13844 );
not \U$13593 ( \13846 , \13845 );
or \U$13594 ( \13847 , \13841 , \13846 );
or \U$13595 ( \13848 , \13845 , \13189 );
nand \U$13596 ( \13849 , \13847 , \13848 );
xor \U$13597 ( \13850 , \13840 , \13849 );
or \U$13598 ( \13851 , \13838 , \13850 );
and \U$13599 ( \13852 , \13638 , \13851 );
and \U$13600 ( \13853 , \13838 , \13850 );
nor \U$13601 ( \13854 , \13852 , \13853 );
not \U$13602 ( \13855 , \13854 );
or \U$13603 ( \13856 , \13432 , \13855 );
and \U$13604 ( \13857 , \13840 , \13849 );
not \U$13605 ( \13858 , \13306 );
not \U$13606 ( \13859 , \13314 );
or \U$13607 ( \13860 , \13858 , \13859 );
not \U$13608 ( \13861 , \13305 );
nand \U$13609 ( \13862 , \12881 , \12868 );
and \U$13610 ( \13863 , \13312 , \13862 );
nor \U$13611 ( \13864 , \13863 , \13307 );
not \U$13612 ( \13865 , \13864 );
or \U$13613 ( \13866 , \13861 , \13865 );
nand \U$13614 ( \13867 , \13866 , \13323 );
nand \U$13615 ( \13868 , \13860 , \13867 );
xor \U$13616 ( \13869 , \13284 , \13290 );
and \U$13617 ( \13870 , \13869 , \13299 );
and \U$13618 ( \13871 , \13284 , \13290 );
or \U$13619 ( \13872 , \13870 , \13871 );
xor \U$13620 ( \13873 , \13868 , \13872 );
not \U$13621 ( \13874 , \13390 );
not \U$13622 ( \13875 , \13357 );
not \U$13623 ( \13876 , \13875 );
or \U$13624 ( \13877 , \13874 , \13876 );
not \U$13625 ( \13878 , \13357 );
not \U$13626 ( \13879 , \13389 );
or \U$13627 ( \13880 , \13878 , \13879 );
nand \U$13628 ( \13881 , \13880 , \13425 );
nand \U$13629 ( \13882 , \13877 , \13881 );
xor \U$13630 ( \13883 , \13873 , \13882 );
nand \U$13631 ( \13884 , \13345 , \13335 );
and \U$13632 ( \13885 , \13884 , \13355 );
nor \U$13633 ( \13886 , \13345 , \13335 );
nor \U$13634 ( \13887 , \13885 , \13886 );
nand \U$13635 ( \13888 , \13424 , \13404 );
and \U$13636 ( \13889 , \13888 , \13414 );
nor \U$13637 ( \13890 , \13424 , \13404 );
nor \U$13638 ( \13891 , \13889 , \13890 );
xor \U$13639 ( \13892 , \13887 , \13891 );
not \U$13640 ( \13893 , RIbe2b018_114);
not \U$13641 ( \13894 , \6855 );
not \U$13642 ( \13895 , \13894 );
or \U$13643 ( \13896 , \13893 , \13895 );
nand \U$13644 ( \13897 , \7528 , RIbe2afa0_113);
nand \U$13645 ( \13898 , \13896 , \13897 );
and \U$13646 ( \13899 , \13898 , \7501 );
not \U$13647 ( \13900 , \13898 );
and \U$13648 ( \13901 , \13900 , \10972 );
nor \U$13649 ( \13902 , \13899 , \13901 );
not \U$13650 ( \13903 , RIbe2aaf0_103);
not \U$13651 ( \13904 , \6630 );
or \U$13652 ( \13905 , \13903 , \13904 );
nand \U$13653 ( \13906 , \6634 , RIbe2b630_127);
nand \U$13654 ( \13907 , \13905 , \13906 );
and \U$13655 ( \13908 , \13907 , \8252 );
not \U$13656 ( \13909 , \13907 );
and \U$13657 ( \13910 , \13909 , \6121 );
nor \U$13658 ( \13911 , \13908 , \13910 );
xor \U$13659 ( \13912 , \13902 , \13911 );
and \U$13660 ( \13913 , \5052 , RIbe2ab68_104);
and \U$13661 ( \13914 , \13913 , \4592 );
not \U$13662 ( \13915 , \13913 );
and \U$13663 ( \13916 , \13915 , \4586 );
nor \U$13664 ( \13917 , \13914 , \13916 );
not \U$13665 ( \13918 , \13917 );
xor \U$13666 ( \13919 , \13912 , \13918 );
xor \U$13667 ( \13920 , \13892 , \13919 );
or \U$13668 ( \13921 , \12725 , \12748 );
nand \U$13669 ( \13922 , \13921 , \12776 );
nand \U$13670 ( \13923 , \12748 , \12725 );
nand \U$13671 ( \13924 , \13922 , \13923 );
not \U$13672 ( \13925 , \13924 );
nand \U$13673 ( \13926 , \13376 , \13388 );
and \U$13674 ( \13927 , \13926 , \13367 );
nor \U$13675 ( \13928 , \13376 , \13388 );
nor \U$13676 ( \13929 , \13927 , \13928 );
not \U$13677 ( \13930 , \13929 );
or \U$13678 ( \13931 , \13925 , \13930 );
not \U$13679 ( \13932 , \13924 );
not \U$13680 ( \13933 , \13929 );
nand \U$13681 ( \13934 , \13932 , \13933 );
nand \U$13682 ( \13935 , \13931 , \13934 );
nand \U$13683 ( \13936 , \12806 , \12817 );
and \U$13684 ( \13937 , \13936 , \12841 );
nor \U$13685 ( \13938 , \12806 , \12817 );
nor \U$13686 ( \13939 , \13937 , \13938 );
not \U$13687 ( \13940 , \13939 );
and \U$13688 ( \13941 , \13935 , \13940 );
not \U$13689 ( \13942 , \13935 );
and \U$13690 ( \13943 , \13942 , \13939 );
nor \U$13691 ( \13944 , \13941 , \13943 );
xnor \U$13692 ( \13945 , \13920 , \13944 );
not \U$13693 ( \13946 , \13945 );
and \U$13694 ( \13947 , \13883 , \13946 );
not \U$13695 ( \13948 , \13883 );
and \U$13696 ( \13949 , \13948 , \13945 );
nor \U$13697 ( \13950 , \13947 , \13949 );
not \U$13698 ( \13951 , RIbe2b180_117);
not \U$13699 ( \13952 , \7941 );
or \U$13700 ( \13953 , \13951 , \13952 );
nand \U$13701 ( \13954 , \13436 , RIbe2b270_119);
nand \U$13702 ( \13955 , \13953 , \13954 );
not \U$13703 ( \13956 , \6582 );
and \U$13704 ( \13957 , \13955 , \13956 );
not \U$13705 ( \13958 , \13955 );
and \U$13706 ( \13959 , \13958 , \6601 );
nor \U$13707 ( \13960 , \13957 , \13959 );
not \U$13708 ( \13961 , RIbe2b108_116);
not \U$13709 ( \13962 , \6958 );
or \U$13710 ( \13963 , \13961 , \13962 );
nand \U$13711 ( \13964 , \8202 , RIbe2b090_115);
nand \U$13712 ( \13965 , \13963 , \13964 );
and \U$13713 ( \13966 , \13965 , \6572 );
not \U$13714 ( \13967 , \13965 );
and \U$13715 ( \13968 , \13967 , \7293 );
nor \U$13716 ( \13969 , \13966 , \13968 );
not \U$13717 ( \13970 , \13969 );
and \U$13718 ( \13971 , \13960 , \13970 );
not \U$13719 ( \13972 , \13960 );
and \U$13720 ( \13973 , \13972 , \13969 );
or \U$13721 ( \13974 , \13971 , \13973 );
not \U$13722 ( \13975 , \7546 );
not \U$13723 ( \13976 , RIbe2af28_112);
not \U$13724 ( \13977 , \6880 );
or \U$13725 ( \13978 , \13976 , \13977 );
nand \U$13726 ( \13979 , \6540 , RIbe2b1f8_118);
nand \U$13727 ( \13980 , \13978 , \13979 );
not \U$13728 ( \13981 , \13980 );
or \U$13729 ( \13982 , \13975 , \13981 );
or \U$13730 ( \13983 , \13980 , \13412 );
nand \U$13731 ( \13984 , \13982 , \13983 );
not \U$13732 ( \13985 , \13984 );
and \U$13733 ( \13986 , \13974 , \13985 );
not \U$13734 ( \13987 , \13974 );
and \U$13735 ( \13988 , \13987 , \13984 );
nor \U$13736 ( \13989 , \13986 , \13988 );
not \U$13737 ( \13990 , \13989 );
not \U$13738 ( \13991 , RIbe2a2f8_86);
not \U$13739 ( \13992 , \12921 );
or \U$13740 ( \13993 , \13991 , \13992 );
nand \U$13741 ( \13994 , \13086 , RIbe2acd0_107);
nand \U$13742 ( \13995 , \13993 , \13994 );
not \U$13743 ( \13996 , \13995 );
not \U$13744 ( \13997 , \12769 );
and \U$13745 ( \13998 , \13996 , \13997 );
not \U$13746 ( \13999 , \12769 );
not \U$13747 ( \14000 , \13999 );
and \U$13748 ( \14001 , \13995 , \14000 );
nor \U$13749 ( \14002 , \13998 , \14001 );
and \U$13750 ( \14003 , \12943 , RIbe2a3e8_88);
and \U$13751 ( \14004 , \13669 , RIbe2a370_87);
nor \U$13752 ( \14005 , \14003 , \14004 );
not \U$13753 ( \14006 , \14005 );
not \U$13754 ( \14007 , \12195 );
and \U$13755 ( \14008 , \14006 , \14007 );
and \U$13756 ( \14009 , \14005 , \12195 );
nor \U$13757 ( \14010 , \14008 , \14009 );
xor \U$13758 ( \14011 , \14002 , \14010 );
not \U$13759 ( \14012 , RIbe2a910_99);
not \U$13760 ( \14013 , \10936 );
or \U$13761 ( \14014 , \14012 , \14013 );
nand \U$13762 ( \14015 , \12971 , RIbe2b5b8_126);
nand \U$13763 ( \14016 , \14014 , \14015 );
not \U$13764 ( \14017 , \14016 );
not \U$13765 ( \14018 , \13030 );
and \U$13766 ( \14019 , \14017 , \14018 );
and \U$13767 ( \14020 , \14016 , \12218 );
nor \U$13768 ( \14021 , \14019 , \14020 );
xor \U$13769 ( \14022 , \14011 , \14021 );
not \U$13770 ( \14023 , \14022 );
not \U$13771 ( \14024 , \14023 );
or \U$13772 ( \14025 , \13990 , \14024 );
not \U$13773 ( \14026 , \13989 );
nand \U$13774 ( \14027 , \14022 , \14026 );
nand \U$13775 ( \14028 , \14025 , \14027 );
and \U$13776 ( \14029 , \8278 , RIbe2a550_91);
and \U$13777 ( \14030 , \13380 , RIbe2a988_100);
nor \U$13778 ( \14031 , \14029 , \14030 );
and \U$13779 ( \14032 , \14031 , \13148 );
not \U$13780 ( \14033 , \14031 );
and \U$13781 ( \14034 , \14033 , \12202 );
nor \U$13782 ( \14035 , \14032 , \14034 );
not \U$13783 ( \14036 , RIbe2a280_85);
not \U$13784 ( \14037 , \6980 );
or \U$13785 ( \14038 , \14036 , \14037 );
nand \U$13786 ( \14039 , \10898 , RIbe2a208_84);
nand \U$13787 ( \14040 , \14038 , \14039 );
not \U$13788 ( \14041 , \14040 );
not \U$13789 ( \14042 , \7301 );
and \U$13790 ( \14043 , \14041 , \14042 );
and \U$13791 ( \14044 , \14040 , \7301 );
nor \U$13792 ( \14045 , \14043 , \14044 );
xor \U$13793 ( \14046 , \14035 , \14045 );
not \U$13794 ( \14047 , RIbe2a190_83);
not \U$13795 ( \14048 , \10949 );
or \U$13796 ( \14049 , \14047 , \14048 );
nand \U$13797 ( \14050 , \10952 , RIbe2a5c8_92);
nand \U$13798 ( \14051 , \14049 , \14050 );
not \U$13799 ( \14052 , \14051 );
not \U$13800 ( \14053 , \6949 );
and \U$13801 ( \14054 , \14052 , \14053 );
and \U$13802 ( \14055 , \14051 , \7989 );
nor \U$13803 ( \14056 , \14054 , \14055 );
xor \U$13804 ( \14057 , \14046 , \14056 );
not \U$13805 ( \14058 , \14057 );
and \U$13806 ( \14059 , \14028 , \14058 );
not \U$13807 ( \14060 , \14028 );
and \U$13808 ( \14061 , \14060 , \14057 );
nor \U$13809 ( \14062 , \14059 , \14061 );
not \U$13810 ( \14063 , \14062 );
not \U$13811 ( \14064 , RIbe29c68_72);
not \U$13812 ( \14065 , \13010 );
or \U$13813 ( \14066 , \14064 , \14065 );
nand \U$13814 ( \14067 , \12835 , RIbe29bf0_71);
nand \U$13815 ( \14068 , \14066 , \14067 );
xor \U$13816 ( \14069 , \14068 , \12823 );
not \U$13817 ( \14070 , RIbe29e48_76);
not \U$13818 ( \14071 , \12731 );
not \U$13819 ( \14072 , \14071 );
or \U$13820 ( \14073 , \14070 , \14072 );
buf \U$13821 ( \14074 , \12735 );
nand \U$13822 ( \14075 , \14074 , RIbe29dd0_75);
nand \U$13823 ( \14076 , \14073 , \14075 );
not \U$13824 ( \14077 , \12746 );
and \U$13825 ( \14078 , \14076 , \14077 );
not \U$13826 ( \14079 , \14076 );
and \U$13827 ( \14080 , \14079 , \12742 );
nor \U$13828 ( \14081 , \14078 , \14080 );
and \U$13829 ( \14082 , \14069 , \14081 );
not \U$13830 ( \14083 , \14069 );
not \U$13831 ( \14084 , \14081 );
and \U$13832 ( \14085 , \14083 , \14084 );
or \U$13833 ( \14086 , \14082 , \14085 );
not \U$13834 ( \14087 , RIbe2a028_80);
not \U$13835 ( \14088 , \13063 );
or \U$13836 ( \14089 , \14087 , \14088 );
nand \U$13837 ( \14090 , \12711 , RIbe29fb0_79);
nand \U$13838 ( \14091 , \14089 , \14090 );
not \U$13839 ( \14092 , \14091 );
not \U$13840 ( \14093 , \12723 );
and \U$13841 ( \14094 , \14092 , \14093 );
and \U$13842 ( \14095 , \14091 , \13583 );
nor \U$13843 ( \14096 , \14094 , \14095 );
xor \U$13844 ( \14097 , \14086 , \14096 );
not \U$13845 ( \14098 , RIbe28f48_44);
not \U$13846 ( \14099 , \13518 );
or \U$13847 ( \14100 , \14098 , \14099 );
nand \U$13848 ( \14101 , \12890 , RIbe28ed0_43);
nand \U$13849 ( \14102 , \14100 , \14101 );
not \U$13850 ( \14103 , \12801 );
and \U$13851 ( \14104 , \14102 , \14103 );
not \U$13852 ( \14105 , \14102 );
and \U$13853 ( \14106 , \14105 , \12801 );
nor \U$13854 ( \14107 , \14104 , \14106 );
not \U$13855 ( \14108 , \4946 );
not \U$13856 ( \14109 , RIbe27fd0_11);
not \U$13857 ( \14110 , \13004 );
or \U$13858 ( \14111 , \14109 , \14110 );
nand \U$13859 ( \14112 , RIbe27f58_10, RIbe2ae38_110);
nand \U$13860 ( \14113 , \14111 , \14112 );
xnor \U$13861 ( \14114 , \14113 , RIbe2aeb0_111);
not \U$13862 ( \14115 , \14114 );
not \U$13863 ( \14116 , \14115 );
or \U$13864 ( \14117 , \14108 , \14116 );
nand \U$13865 ( \14118 , \14114 , \4586 );
nand \U$13866 ( \14119 , \14117 , \14118 );
xnor \U$13867 ( \14120 , \14107 , \14119 );
xnor \U$13868 ( \14121 , \14097 , \14120 );
not \U$13869 ( \14122 , \14121 );
and \U$13870 ( \14123 , \14063 , \14122 );
and \U$13871 ( \14124 , \14121 , \14062 );
nor \U$13872 ( \14125 , \14123 , \14124 );
xor \U$13873 ( \14126 , \13950 , \14125 );
xor \U$13874 ( \14127 , \13857 , \14126 );
xor \U$13875 ( \14128 , \13618 , \13634 );
and \U$13876 ( \14129 , \14128 , \13637 );
and \U$13877 ( \14130 , \13618 , \13634 );
or \U$13878 ( \14131 , \14129 , \14130 );
xor \U$13879 ( \14132 , \14127 , \14131 );
nand \U$13880 ( \14133 , \13856 , \14132 );
or \U$13881 ( \14134 , \13854 , \13431 );
nand \U$13882 ( \14135 , \14133 , \14134 );
not \U$13883 ( \14136 , \13920 );
nand \U$13884 ( \14137 , \14136 , \13944 );
or \U$13885 ( \14138 , \13872 , \13868 );
and \U$13886 ( \14139 , \13882 , \14138 );
and \U$13887 ( \14140 , \13868 , \13872 );
nor \U$13888 ( \14141 , \14139 , \14140 );
not \U$13889 ( \14142 , \14141 );
xor \U$13890 ( \14143 , \14137 , \14142 );
nand \U$13891 ( \14144 , \14097 , \14120 );
not \U$13892 ( \14145 , \14144 );
not \U$13893 ( \14146 , \14062 );
or \U$13894 ( \14147 , \14145 , \14146 );
or \U$13895 ( \14148 , \14097 , \14120 );
nand \U$13896 ( \14149 , \14147 , \14148 );
xor \U$13897 ( \14150 , \14143 , \14149 );
xor \U$13898 ( \14151 , \13857 , \14126 );
and \U$13899 ( \14152 , \14151 , \14131 );
and \U$13900 ( \14153 , \13857 , \14126 );
or \U$13901 ( \14154 , \14152 , \14153 );
xor \U$13902 ( \14155 , \14150 , \14154 );
not \U$13903 ( \14156 , \13946 );
not \U$13904 ( \14157 , \14125 );
or \U$13905 ( \14158 , \14156 , \14157 );
nand \U$13906 ( \14159 , \14158 , \13883 );
not \U$13907 ( \14160 , \14125 );
nand \U$13908 ( \14161 , \14160 , \13945 );
nand \U$13909 ( \14162 , \14159 , \14161 );
not \U$13910 ( \14163 , \14162 );
xor \U$13911 ( \14164 , \12989 , \13273 );
and \U$13912 ( \14165 , \14164 , \13430 );
and \U$13913 ( \14166 , \12989 , \13273 );
or \U$13914 ( \14167 , \14165 , \14166 );
not \U$13915 ( \14168 , \14167 );
and \U$13916 ( \14169 , \14163 , \14168 );
and \U$13917 ( \14170 , \14162 , \14167 );
nor \U$13918 ( \14171 , \14169 , \14170 );
not \U$13919 ( \14172 , \14171 );
xor \U$13920 ( \14173 , \14002 , \14010 );
and \U$13921 ( \14174 , \14173 , \14021 );
and \U$13922 ( \14175 , \14002 , \14010 );
or \U$13923 ( \14176 , \14174 , \14175 );
not \U$13924 ( \14177 , \4586 );
not \U$13925 ( \14178 , \14115 );
or \U$13926 ( \14179 , \14177 , \14178 );
nand \U$13927 ( \14180 , \14114 , \4592 );
nand \U$13928 ( \14181 , \14107 , \14180 );
nand \U$13929 ( \14182 , \14179 , \14181 );
and \U$13930 ( \14183 , \14176 , \14182 );
not \U$13931 ( \14184 , \14176 );
not \U$13932 ( \14185 , \14182 );
and \U$13933 ( \14186 , \14184 , \14185 );
nor \U$13934 ( \14187 , \14183 , \14186 );
not \U$13935 ( \14188 , \14096 );
not \U$13936 ( \14189 , \14084 );
and \U$13937 ( \14190 , \14188 , \14189 );
and \U$13938 ( \14191 , \14084 , \14096 );
nor \U$13939 ( \14192 , \14191 , \14069 );
nor \U$13940 ( \14193 , \14190 , \14192 );
xor \U$13941 ( \14194 , \14187 , \14193 );
not \U$13942 ( \14195 , \14058 );
not \U$13943 ( \14196 , \14026 );
or \U$13944 ( \14197 , \14195 , \14196 );
not \U$13945 ( \14198 , \13989 );
not \U$13946 ( \14199 , \14057 );
or \U$13947 ( \14200 , \14198 , \14199 );
nand \U$13948 ( \14201 , \14200 , \14023 );
nand \U$13949 ( \14202 , \14197 , \14201 );
not \U$13950 ( \14203 , \14202 );
not \U$13951 ( \14204 , \14203 );
xor \U$13952 ( \14205 , \13887 , \13891 );
and \U$13953 ( \14206 , \14205 , \13919 );
and \U$13954 ( \14207 , \13887 , \13891 );
or \U$13955 ( \14208 , \14206 , \14207 );
not \U$13956 ( \14209 , \13940 );
not \U$13957 ( \14210 , \13933 );
or \U$13958 ( \14211 , \14209 , \14210 );
not \U$13959 ( \14212 , \13939 );
not \U$13960 ( \14213 , \13929 );
or \U$13961 ( \14214 , \14212 , \14213 );
nand \U$13962 ( \14215 , \14214 , \13924 );
nand \U$13963 ( \14216 , \14211 , \14215 );
not \U$13964 ( \14217 , \14216 );
and \U$13965 ( \14218 , \14208 , \14217 );
not \U$13966 ( \14219 , \14208 );
and \U$13967 ( \14220 , \14219 , \14216 );
nor \U$13968 ( \14221 , \14218 , \14220 );
not \U$13969 ( \14222 , \14221 );
or \U$13970 ( \14223 , \14204 , \14222 );
or \U$13971 ( \14224 , \14221 , \14203 );
nand \U$13972 ( \14225 , \14223 , \14224 );
xor \U$13973 ( \14226 , \14194 , \14225 );
not \U$13974 ( \14227 , RIbe2ab68_104);
not \U$13975 ( \14228 , \5727 );
or \U$13976 ( \14229 , \14227 , \14228 );
nand \U$13977 ( \14230 , \5052 , RIbe2aaf0_103);
nand \U$13978 ( \14231 , \14229 , \14230 );
and \U$13979 ( \14232 , \14231 , \4586 );
not \U$13980 ( \14233 , \14231 );
and \U$13981 ( \14234 , \14233 , \4592 );
nor \U$13982 ( \14235 , \14232 , \14234 );
not \U$13983 ( \14236 , RIbe2b630_127);
not \U$13984 ( \14237 , \5455 );
or \U$13985 ( \14238 , \14236 , \14237 );
not \U$13986 ( \14239 , \5750 );
nand \U$13987 ( \14240 , \14239 , RIbe2b018_114);
nand \U$13988 ( \14241 , \14238 , \14240 );
and \U$13989 ( \14242 , \14241 , \6642 );
not \U$13990 ( \14243 , \14241 );
and \U$13991 ( \14244 , \14243 , \5754 );
nor \U$13992 ( \14245 , \14242 , \14244 );
xor \U$13993 ( \14246 , \14235 , \14245 );
not \U$13994 ( \14247 , \6883 );
not \U$13995 ( \14248 , RIbe2b180_117);
not \U$13996 ( \14249 , \14248 );
and \U$13997 ( \14250 , \14247 , \14249 );
and \U$13998 ( \14251 , \6535 , RIbe2b1f8_118);
nor \U$13999 ( \14252 , \14250 , \14251 );
and \U$14000 ( \14253 , \14252 , \9933 );
not \U$14001 ( \14254 , \14252 );
and \U$14002 ( \14255 , \14254 , \6546 );
nor \U$14003 ( \14256 , \14253 , \14255 );
not \U$14004 ( \14257 , RIbe2b270_119);
not \U$14005 ( \14258 , \6591 );
or \U$14006 ( \14259 , \14257 , \14258 );
nand \U$14007 ( \14260 , RIbe2b108_116, \13436 );
nand \U$14008 ( \14261 , \14259 , \14260 );
not \U$14009 ( \14262 , \6601 );
and \U$14010 ( \14263 , \14261 , \14262 );
not \U$14011 ( \14264 , \14261 );
and \U$14012 ( \14265 , \14264 , \7948 );
nor \U$14013 ( \14266 , \14263 , \14265 );
and \U$14014 ( \14267 , \14256 , \14266 );
not \U$14015 ( \14268 , \14256 );
not \U$14016 ( \14269 , \14266 );
and \U$14017 ( \14270 , \14268 , \14269 );
or \U$14018 ( \14271 , \14267 , \14270 );
not \U$14019 ( \14272 , \7535 );
not \U$14020 ( \14273 , RIbe2afa0_113);
not \U$14021 ( \14274 , \12268 );
or \U$14022 ( \14275 , \14273 , \14274 );
nand \U$14023 ( \14276 , \7087 , RIbe2af28_112);
nand \U$14024 ( \14277 , \14275 , \14276 );
not \U$14025 ( \14278 , \14277 );
or \U$14026 ( \14279 , \14272 , \14278 );
or \U$14027 ( \14280 , \14277 , \6141 );
nand \U$14028 ( \14281 , \14279 , \14280 );
xor \U$14029 ( \14282 , \14271 , \14281 );
xor \U$14030 ( \14283 , \14246 , \14282 );
and \U$14031 ( \14284 , \13171 , RIbe2a208_84);
not \U$14032 ( \14285 , RIbe2a190_83);
nor \U$14033 ( \14286 , \10897 , \14285 );
nor \U$14034 ( \14287 , \14284 , \14286 );
and \U$14035 ( \14288 , \14287 , \6993 );
not \U$14036 ( \14289 , \14287 );
and \U$14037 ( \14290 , \14289 , \7301 );
nor \U$14038 ( \14291 , \14288 , \14290 );
not \U$14039 ( \14292 , \14291 );
not \U$14040 ( \14293 , \14292 );
not \U$14041 ( \14294 , RIbe2a5c8_92);
not \U$14042 ( \14295 , \10949 );
or \U$14043 ( \14296 , \14294 , \14295 );
nand \U$14044 ( \14297 , \9891 , RIbe2a550_91);
nand \U$14045 ( \14298 , \14296 , \14297 );
not \U$14046 ( \14299 , \6948 );
and \U$14047 ( \14300 , \14298 , \14299 );
not \U$14048 ( \14301 , \14298 );
not \U$14049 ( \14302 , \7985 );
and \U$14050 ( \14303 , \14301 , \14302 );
nor \U$14051 ( \14304 , \14300 , \14303 );
not \U$14052 ( \14305 , \14304 );
not \U$14053 ( \14306 , \14305 );
or \U$14054 ( \14307 , \14293 , \14306 );
nand \U$14055 ( \14308 , \14304 , \14291 );
nand \U$14056 ( \14309 , \14307 , \14308 );
not \U$14057 ( \14310 , RIbe2b090_115);
not \U$14058 ( \14311 , \13327 );
or \U$14059 ( \14312 , \14310 , \14311 );
nand \U$14060 ( \14313 , \7653 , RIbe2a280_85);
nand \U$14061 ( \14314 , \14312 , \14313 );
and \U$14062 ( \14315 , \14314 , \7293 );
not \U$14063 ( \14316 , \14314 );
and \U$14064 ( \14317 , \14316 , \6569 );
nor \U$14065 ( \14318 , \14315 , \14317 );
xnor \U$14066 ( \14319 , \14309 , \14318 );
xnor \U$14067 ( \14320 , \14283 , \14319 );
not \U$14068 ( \14321 , RIbe27f58_10);
not \U$14069 ( \14322 , \12811 );
or \U$14070 ( \14323 , \14321 , \14322 );
nand \U$14071 ( \14324 , RIbe27e68_8, RIbe2ae38_110);
nand \U$14072 ( \14325 , \14323 , \14324 );
xor \U$14073 ( \14326 , \14325 , RIbe2aeb0_111);
not \U$14074 ( \14327 , RIbe28ed0_43);
not \U$14075 ( \14328 , \12786 );
or \U$14076 ( \14329 , \14327 , \14328 );
nand \U$14077 ( \14330 , \12794 , RIbe27fd0_11);
nand \U$14078 ( \14331 , \14329 , \14330 );
not \U$14079 ( \14332 , RIbe2aeb0_111);
not \U$14080 ( \14333 , RIbe2b3d8_122);
or \U$14081 ( \14334 , \14332 , \14333 );
nand \U$14082 ( \14335 , \14334 , RIbe2b450_123);
not \U$14083 ( \14336 , \14335 );
and \U$14084 ( \14337 , \14331 , \14336 );
not \U$14085 ( \14338 , \14331 );
and \U$14086 ( \14339 , \14338 , \14335 );
nor \U$14087 ( \14340 , \14337 , \14339 );
xor \U$14088 ( \14341 , \14326 , \14340 );
not \U$14089 ( \14342 , RIbe29bf0_71);
not \U$14090 ( \14343 , \12858 );
or \U$14091 ( \14344 , \14342 , \14343 );
nand \U$14092 ( \14345 , \12835 , RIbe28f48_44);
nand \U$14093 ( \14346 , \14344 , \14345 );
and \U$14094 ( \14347 , \14346 , \13705 );
not \U$14095 ( \14348 , \14346 );
and \U$14096 ( \14349 , \14348 , \12823 );
nor \U$14097 ( \14350 , \14347 , \14349 );
xnor \U$14098 ( \14351 , \14341 , \14350 );
not \U$14099 ( \14352 , RIbe29dd0_75);
not \U$14100 ( \14353 , \14071 );
or \U$14101 ( \14354 , \14352 , \14353 );
not \U$14102 ( \14355 , \9801 );
nand \U$14103 ( \14356 , \14355 , \12735 );
nand \U$14104 ( \14357 , \14354 , \14356 );
not \U$14105 ( \14358 , \12741 );
and \U$14106 ( \14359 , \14357 , \14358 );
not \U$14107 ( \14360 , \14357 );
and \U$14108 ( \14361 , \14360 , \12746 );
nor \U$14109 ( \14362 , \14359 , \14361 );
not \U$14110 ( \14363 , RIbe29fb0_79);
not \U$14111 ( \14364 , \12707 );
or \U$14112 ( \14365 , \14363 , \14364 );
nand \U$14113 ( \14366 , RIbe29e48_76, \13728 );
nand \U$14114 ( \14367 , \14365 , \14366 );
and \U$14115 ( \14368 , \14367 , \13068 );
not \U$14116 ( \14369 , \14367 );
and \U$14117 ( \14370 , \14369 , \12723 );
nor \U$14118 ( \14371 , \14368 , \14370 );
xor \U$14119 ( \14372 , \14362 , \14371 );
not \U$14120 ( \14373 , \12751 );
not \U$14121 ( \14374 , RIbe2a028_80);
not \U$14122 ( \14375 , \14374 );
and \U$14123 ( \14376 , \14373 , \14375 );
and \U$14124 ( \14377 , \13738 , RIbe2acd0_107);
nor \U$14125 ( \14378 , \14376 , \14377 );
and \U$14126 ( \14379 , \14378 , \12770 );
not \U$14127 ( \14380 , \14378 );
and \U$14128 ( \14381 , \14380 , \12927 );
nor \U$14129 ( \14382 , \14379 , \14381 );
xnor \U$14130 ( \14383 , \14372 , \14382 );
xor \U$14131 ( \14384 , \14351 , \14383 );
not \U$14132 ( \14385 , RIbe2b5b8_126);
not \U$14133 ( \14386 , \10936 );
or \U$14134 ( \14387 , \14385 , \14386 );
nand \U$14135 ( \14388 , \12213 , RIbe2a3e8_88);
nand \U$14136 ( \14389 , \14387 , \14388 );
not \U$14137 ( \14390 , \14389 );
not \U$14138 ( \14391 , \12218 );
and \U$14139 ( \14392 , \14390 , \14391 );
and \U$14140 ( \14393 , \14389 , \10940 );
nor \U$14141 ( \14394 , \14392 , \14393 );
and \U$14142 ( \14395 , \12942 , RIbe2a370_87);
not \U$14143 ( \14396 , RIbe2a2f8_86);
not \U$14144 ( \14397 , \12947 );
nor \U$14145 ( \14398 , \14396 , \14397 );
nor \U$14146 ( \14399 , \14395 , \14398 );
and \U$14147 ( \14400 , \14399 , \12956 );
not \U$14148 ( \14401 , \14399 );
and \U$14149 ( \14402 , \14401 , \12195 );
nor \U$14150 ( \14403 , \14400 , \14402 );
xor \U$14151 ( \14404 , \14394 , \14403 );
and \U$14152 ( \14405 , \9909 , RIbe2a988_100);
and \U$14153 ( \14406 , \10921 , RIbe2a910_99);
nor \U$14154 ( \14407 , \14405 , \14406 );
and \U$14155 ( \14408 , \14407 , \8077 );
not \U$14156 ( \14409 , \14407 );
and \U$14157 ( \14410 , \14409 , \13148 );
nor \U$14158 ( \14411 , \14408 , \14410 );
xor \U$14159 ( \14412 , \14404 , \14411 );
xor \U$14160 ( \14413 , \14384 , \14412 );
nand \U$14161 ( \14414 , \13911 , \13917 );
and \U$14162 ( \14415 , \14414 , \13902 );
nor \U$14163 ( \14416 , \13911 , \13917 );
nor \U$14164 ( \14417 , \14415 , \14416 );
not \U$14165 ( \14418 , \14417 );
not \U$14166 ( \14419 , \14418 );
not \U$14167 ( \14420 , \13969 );
not \U$14168 ( \14421 , \13960 );
or \U$14169 ( \14422 , \14420 , \14421 );
nand \U$14170 ( \14423 , \14422 , \13984 );
not \U$14171 ( \14424 , \13960 );
nand \U$14172 ( \14425 , \14424 , \13970 );
nand \U$14173 ( \14426 , \14423 , \14425 );
not \U$14174 ( \14427 , \14426 );
not \U$14175 ( \14428 , \14427 );
or \U$14176 ( \14429 , \14419 , \14428 );
nand \U$14177 ( \14430 , \14426 , \14417 );
nand \U$14178 ( \14431 , \14429 , \14430 );
xor \U$14179 ( \14432 , \14035 , \14045 );
and \U$14180 ( \14433 , \14432 , \14056 );
and \U$14181 ( \14434 , \14035 , \14045 );
or \U$14182 ( \14435 , \14433 , \14434 );
xor \U$14183 ( \14436 , \14431 , \14435 );
and \U$14184 ( \14437 , \14413 , \14436 );
not \U$14185 ( \14438 , \14413 );
not \U$14186 ( \14439 , \14436 );
and \U$14187 ( \14440 , \14438 , \14439 );
nor \U$14188 ( \14441 , \14437 , \14440 );
xor \U$14189 ( \14442 , \14320 , \14441 );
xor \U$14190 ( \14443 , \14226 , \14442 );
not \U$14191 ( \14444 , \14443 );
and \U$14192 ( \14445 , \14172 , \14444 );
and \U$14193 ( \14446 , \14171 , \14443 );
nor \U$14194 ( \14447 , \14445 , \14446 );
not \U$14195 ( \14448 , \14447 );
xnor \U$14196 ( \14449 , \14155 , \14448 );
xor \U$14197 ( \14450 , \14135 , \14449 );
xor \U$14198 ( \14451 , \13758 , \13801 );
xor \U$14199 ( \14452 , \14451 , \13762 );
not \U$14200 ( \14453 , \14452 );
xor \U$14201 ( \14454 , \7501 , \13514 );
xor \U$14202 ( \14455 , \14454 , \13526 );
not \U$14203 ( \14456 , \14455 );
nand \U$14204 ( \14457 , \14453 , \14456 );
not \U$14205 ( \14458 , \13809 );
not \U$14206 ( \14459 , \13816 );
or \U$14207 ( \14460 , \14458 , \14459 );
or \U$14208 ( \14461 , \13816 , \13809 );
nand \U$14209 ( \14462 , \14460 , \14461 );
and \U$14210 ( \14463 , \14462 , \13812 );
not \U$14211 ( \14464 , \14462 );
and \U$14212 ( \14465 , \14464 , \13819 );
nor \U$14213 ( \14466 , \14463 , \14465 );
not \U$14214 ( \14467 , \14466 );
and \U$14215 ( \14468 , \14457 , \14467 );
nor \U$14216 ( \14469 , \14453 , \14456 );
nor \U$14217 ( \14470 , \14468 , \14469 );
not \U$14218 ( \14471 , \6541 );
not \U$14219 ( \14472 , \13192 );
and \U$14220 ( \14473 , \14471 , \14472 );
and \U$14221 ( \14474 , \6537 , RIbe2ab68_104);
nor \U$14222 ( \14475 , \14473 , \14474 );
and \U$14223 ( \14476 , \14475 , \13412 );
not \U$14224 ( \14477 , \14475 );
and \U$14225 ( \14478 , \14477 , \7935 );
nor \U$14226 ( \14479 , \14476 , \14478 );
xor \U$14227 ( \14480 , \13675 , \13663 );
buf \U$14228 ( \14481 , \13652 );
xor \U$14229 ( \14482 , \14480 , \14481 );
xor \U$14230 ( \14483 , \14479 , \14482 );
xor \U$14231 ( \14484 , \13798 , \13785 );
xnor \U$14232 ( \14485 , \14484 , \13775 );
and \U$14233 ( \14486 , \14483 , \14485 );
and \U$14234 ( \14487 , \14479 , \14482 );
or \U$14235 ( \14488 , \14486 , \14487 );
not \U$14236 ( \14489 , \14488 );
and \U$14237 ( \14490 , \12921 , RIbe2a550_91);
not \U$14238 ( \14491 , \13085 );
and \U$14239 ( \14492 , \14491 , RIbe2a988_100);
nor \U$14240 ( \14493 , \14490 , \14492 );
and \U$14241 ( \14494 , \14493 , \12924 );
not \U$14242 ( \14495 , \14493 );
and \U$14243 ( \14496 , \14495 , \12927 );
nor \U$14244 ( \14497 , \14494 , \14496 );
and \U$14245 ( \14498 , \12943 , RIbe2a190_83);
and \U$14246 ( \14499 , \13669 , RIbe2a5c8_92);
nor \U$14247 ( \14500 , \14498 , \14499 );
not \U$14248 ( \14501 , \14500 );
not \U$14249 ( \14502 , \12195 );
or \U$14250 ( \14503 , \14501 , \14502 );
or \U$14251 ( \14504 , \14500 , \12195 );
nand \U$14252 ( \14505 , \14503 , \14504 );
xor \U$14253 ( \14506 , \14497 , \14505 );
not \U$14254 ( \14507 , \12218 );
not \U$14255 ( \14508 , RIbe2a280_85);
not \U$14256 ( \14509 , \13024 );
or \U$14257 ( \14510 , \14508 , \14509 );
buf \U$14258 ( \14511 , \12212 );
nand \U$14259 ( \14512 , \14511 , RIbe2a208_84);
nand \U$14260 ( \14513 , \14510 , \14512 );
not \U$14261 ( \14514 , \14513 );
or \U$14262 ( \14515 , \14507 , \14514 );
or \U$14263 ( \14516 , \14513 , \9903 );
nand \U$14264 ( \14517 , \14515 , \14516 );
and \U$14265 ( \14518 , \14506 , \14517 );
and \U$14266 ( \14519 , \14497 , \14505 );
or \U$14267 ( \14520 , \14518 , \14519 );
not \U$14268 ( \14521 , \14520 );
not \U$14269 ( \14522 , RIbe2a910_99);
not \U$14270 ( \14523 , \12706 );
not \U$14271 ( \14524 , \14523 );
or \U$14272 ( \14525 , \14522 , \14524 );
nand \U$14273 ( \14526 , RIbe2b5b8_126, \13728 );
nand \U$14274 ( \14527 , \14525 , \14526 );
and \U$14275 ( \14528 , \14527 , \12723 );
not \U$14276 ( \14529 , \14527 );
and \U$14277 ( \14530 , \14529 , \12879 );
nor \U$14278 ( \14531 , \14528 , \14530 );
not \U$14279 ( \14532 , RIbe2a3e8_88);
nand \U$14280 ( \14533 , \12728 , \12729 );
not \U$14281 ( \14534 , \14533 );
not \U$14282 ( \14535 , \14534 );
or \U$14283 ( \14536 , \14532 , \14535 );
nand \U$14284 ( \14537 , \12735 , RIbe2a370_87);
nand \U$14285 ( \14538 , \14536 , \14537 );
not \U$14286 ( \14539 , RIbe2abe0_105);
not \U$14287 ( \14540 , RIbe2a7a8_96);
or \U$14288 ( \14541 , \14539 , \14540 );
nand \U$14289 ( \14542 , \14541 , RIbe2ac58_106);
buf \U$14290 ( \14543 , \14542 );
and \U$14291 ( \14544 , \14538 , \14543 );
not \U$14292 ( \14545 , \14538 );
and \U$14293 ( \14546 , \14545 , \14077 );
nor \U$14294 ( \14547 , \14544 , \14546 );
nand \U$14295 ( \14548 , \14531 , \14547 );
not \U$14296 ( \14549 , RIbe2a2f8_86);
and \U$14297 ( \14550 , \12827 , \12828 );
not \U$14298 ( \14551 , \14550 );
or \U$14299 ( \14552 , \14549 , \14551 );
nand \U$14300 ( \14553 , \12834 , RIbe2acd0_107);
nand \U$14301 ( \14554 , \14552 , \14553 );
not \U$14302 ( \14555 , \12863 );
and \U$14303 ( \14556 , \14554 , \14555 );
not \U$14304 ( \14557 , \14554 );
not \U$14305 ( \14558 , \13595 );
and \U$14306 ( \14559 , \14557 , \14558 );
nor \U$14307 ( \14560 , \14556 , \14559 );
and \U$14308 ( \14561 , \14548 , \14560 );
nor \U$14309 ( \14562 , \14531 , \14547 );
nor \U$14310 ( \14563 , \14561 , \14562 );
not \U$14311 ( \14564 , RIbe2a028_80);
not \U$14312 ( \14565 , \13518 );
or \U$14313 ( \14566 , \14564 , \14565 );
nand \U$14314 ( \14567 , \12794 , RIbe29fb0_79);
nand \U$14315 ( \14568 , \14566 , \14567 );
xnor \U$14316 ( \14569 , \14568 , \12893 );
not \U$14317 ( \14570 , RIbe29e48_76);
not \U$14318 ( \14571 , \13690 );
or \U$14319 ( \14572 , \14570 , \14571 );
nand \U$14320 ( \14573 , RIbe29dd0_75, RIbe2ae38_110);
nand \U$14321 ( \14574 , \14572 , \14573 );
xor \U$14322 ( \14575 , \14574 , RIbe2aeb0_111);
not \U$14323 ( \14576 , \14575 );
nand \U$14324 ( \14577 , \14576 , \13412 );
and \U$14325 ( \14578 , \14569 , \14577 );
nor \U$14326 ( \14579 , \14576 , \7546 );
nor \U$14327 ( \14580 , \14578 , \14579 );
nand \U$14328 ( \14581 , \14563 , \14580 );
not \U$14329 ( \14582 , \14581 );
or \U$14330 ( \14583 , \14521 , \14582 );
not \U$14331 ( \14584 , \14580 );
not \U$14332 ( \14585 , \14563 );
nand \U$14333 ( \14586 , \14584 , \14585 );
nand \U$14334 ( \14587 , \14583 , \14586 );
not \U$14335 ( \14588 , \14587 );
nand \U$14336 ( \14589 , \6540 , RIbe2ab68_104);
and \U$14337 ( \14590 , \14589 , \13412 );
not \U$14338 ( \14591 , \14589 );
and \U$14339 ( \14592 , \14591 , \6546 );
nor \U$14340 ( \14593 , \14590 , \14592 );
not \U$14341 ( \14594 , \14593 );
not \U$14342 ( \14595 , \14594 );
not \U$14343 ( \14596 , RIbe2aaf0_103);
not \U$14344 ( \14597 , \7274 );
or \U$14345 ( \14598 , \14596 , \14597 );
nand \U$14346 ( \14599 , RIbe2b630_127, \6596 );
nand \U$14347 ( \14600 , \14598 , \14599 );
not \U$14348 ( \14601 , \14600 );
not \U$14349 ( \14602 , \7949 );
and \U$14350 ( \14603 , \14601 , \14602 );
and \U$14351 ( \14604 , \14600 , \14262 );
nor \U$14352 ( \14605 , \14603 , \14604 );
not \U$14353 ( \14606 , \14605 );
or \U$14354 ( \14607 , \14595 , \14606 );
not \U$14355 ( \14608 , RIbe2b018_114);
not \U$14356 ( \14609 , \7954 );
or \U$14357 ( \14610 , \14608 , \14609 );
nand \U$14358 ( \14611 , \8202 , RIbe2afa0_113);
nand \U$14359 ( \14612 , \14610 , \14611 );
and \U$14360 ( \14613 , \14612 , \7293 );
not \U$14361 ( \14614 , \14612 );
and \U$14362 ( \14615 , \14614 , \6572 );
nor \U$14363 ( \14616 , \14613 , \14615 );
nand \U$14364 ( \14617 , \14607 , \14616 );
not \U$14365 ( \14618 , \14605 );
nand \U$14366 ( \14619 , \14618 , \14593 );
nand \U$14367 ( \14620 , \14617 , \14619 );
not \U$14368 ( \14621 , RIbe2b108_116);
nor \U$14369 ( \14622 , \8274 , \8273 );
not \U$14370 ( \14623 , \14622 );
or \U$14371 ( \14624 , \14621 , \14623 );
nand \U$14372 ( \14625 , RIbe2b090_115, \13038 );
nand \U$14373 ( \14626 , \14624 , \14625 );
and \U$14374 ( \14627 , \14626 , \13649 );
not \U$14375 ( \14628 , \14626 );
and \U$14376 ( \14629 , \14628 , \8077 );
nor \U$14377 ( \14630 , \14627 , \14629 );
not \U$14378 ( \14631 , \14630 );
not \U$14379 ( \14632 , RIbe2b180_117);
and \U$14380 ( \14633 , \7979 , \6939 );
not \U$14381 ( \14634 , \14633 );
or \U$14382 ( \14635 , \14632 , \14634 );
nand \U$14383 ( \14636 , \9891 , RIbe2b270_119);
nand \U$14384 ( \14637 , \14635 , \14636 );
and \U$14385 ( \14638 , \14637 , \7984 );
not \U$14386 ( \14639 , \14637 );
and \U$14387 ( \14640 , \14639 , \6950 );
nor \U$14388 ( \14641 , \14638 , \14640 );
nand \U$14389 ( \14642 , \14631 , \14641 );
not \U$14390 ( \14643 , \8287 );
not \U$14391 ( \14644 , \14643 );
not \U$14392 ( \14645 , RIbe2b1f8_118);
not \U$14393 ( \14646 , \14645 );
and \U$14394 ( \14647 , \14644 , \14646 );
and \U$14395 ( \14648 , \6980 , RIbe2af28_112);
nor \U$14396 ( \14649 , \14647 , \14648 );
not \U$14397 ( \14650 , \6993 );
and \U$14398 ( \14651 , \14649 , \14650 );
not \U$14399 ( \14652 , \14649 );
and \U$14400 ( \14653 , \14652 , \13227 );
nor \U$14401 ( \14654 , \14651 , \14653 );
and \U$14402 ( \14655 , \14642 , \14654 );
nor \U$14403 ( \14656 , \14641 , \14631 );
nor \U$14404 ( \14657 , \14655 , \14656 );
not \U$14405 ( \14658 , RIbe2b630_127);
not \U$14406 ( \14659 , \6592 );
or \U$14407 ( \14660 , \14658 , \14659 );
nand \U$14408 ( \14661 , \6596 , RIbe2b018_114);
nand \U$14409 ( \14662 , \14660 , \14661 );
not \U$14410 ( \14663 , \14662 );
not \U$14411 ( \14664 , \7646 );
and \U$14412 ( \14665 , \14663 , \14664 );
not \U$14413 ( \14666 , \6601 );
and \U$14414 ( \14667 , \14662 , \14666 );
nor \U$14415 ( \14668 , \14665 , \14667 );
nand \U$14416 ( \14669 , \14657 , \14668 );
and \U$14417 ( \14670 , \14620 , \14669 );
nor \U$14418 ( \14671 , \14657 , \14668 );
nor \U$14419 ( \14672 , \14670 , \14671 );
nand \U$14420 ( \14673 , \14588 , \14672 );
not \U$14421 ( \14674 , \14673 );
or \U$14422 ( \14675 , \14489 , \14674 );
not \U$14423 ( \14676 , \14672 );
nand \U$14424 ( \14677 , \14676 , \14587 );
nand \U$14425 ( \14678 , \14675 , \14677 );
xor \U$14426 ( \14679 , \13529 , \13561 );
xor \U$14427 ( \14680 , \14679 , \13601 );
nor \U$14428 ( \14681 , \14678 , \14680 );
or \U$14429 ( \14682 , \14470 , \14681 );
nand \U$14430 ( \14683 , \14678 , \14680 );
nand \U$14431 ( \14684 , \14682 , \14683 );
xor \U$14432 ( \14685 , \13620 , \13622 );
xor \U$14433 ( \14686 , \14685 , \13631 );
xor \U$14434 ( \14687 , \14684 , \14686 );
xor \U$14435 ( \14688 , \13827 , \13829 );
xor \U$14436 ( \14689 , \14688 , \13832 );
xor \U$14437 ( \14690 , \13753 , \13803 );
xor \U$14438 ( \14691 , \14690 , \13821 );
and \U$14439 ( \14692 , \14689 , \14691 );
and \U$14440 ( \14693 , \14687 , \14692 );
and \U$14441 ( \14694 , \14684 , \14686 );
or \U$14442 ( \14695 , \14693 , \14694 );
not \U$14443 ( \14696 , \14695 );
xor \U$14444 ( \14697 , \13640 , \13824 );
xor \U$14445 ( \14698 , \14697 , \13835 );
xor \U$14446 ( \14699 , \13508 , \13604 );
xor \U$14447 ( \14700 , \14699 , \13615 );
nand \U$14448 ( \14701 , \14698 , \14700 );
not \U$14449 ( \14702 , \14701 );
not \U$14450 ( \14703 , \14702 );
or \U$14451 ( \14704 , \14696 , \14703 );
or \U$14452 ( \14705 , \14702 , \14695 );
xor \U$14453 ( \14706 , \13838 , \13850 );
xor \U$14454 ( \14707 , \14706 , \13638 );
nand \U$14455 ( \14708 , \14705 , \14707 );
nand \U$14456 ( \14709 , \14704 , \14708 );
not \U$14457 ( \14710 , \14709 );
xor \U$14458 ( \14711 , \13431 , \13854 );
not \U$14459 ( \14712 , \14132 );
and \U$14460 ( \14713 , \14711 , \14712 );
not \U$14461 ( \14714 , \14711 );
and \U$14462 ( \14715 , \14714 , \14132 );
nor \U$14463 ( \14716 , \14713 , \14715 );
nor \U$14464 ( \14717 , \14710 , \14716 );
and \U$14465 ( \14718 , \14450 , \14717 );
and \U$14466 ( \14719 , \14135 , \14449 );
nor \U$14467 ( \14720 , \14718 , \14719 );
not \U$14468 ( \14721 , \12752 );
not \U$14469 ( \14722 , RIbe29fb0_79);
not \U$14470 ( \14723 , \14722 );
and \U$14471 ( \14724 , \14721 , \14723 );
not \U$14472 ( \14725 , \12763 );
buf \U$14473 ( \14726 , \14725 );
and \U$14474 ( \14727 , \14726 , RIbe2a028_80);
nor \U$14475 ( \14728 , \14724 , \14727 );
and \U$14476 ( \14729 , \14728 , \12770 );
not \U$14477 ( \14730 , \14728 );
and \U$14478 ( \14731 , \14730 , \12927 );
nor \U$14479 ( \14732 , \14729 , \14731 );
not \U$14480 ( \14733 , \14732 );
not \U$14481 ( \14734 , \14733 );
not \U$14482 ( \14735 , RIbe2a2f8_86);
not \U$14483 ( \14736 , \12943 );
or \U$14484 ( \14737 , \14735 , \14736 );
nand \U$14485 ( \14738 , \12947 , RIbe2acd0_107);
nand \U$14486 ( \14739 , \14737 , \14738 );
not \U$14487 ( \14740 , \14739 );
not \U$14488 ( \14741 , \12957 );
and \U$14489 ( \14742 , \14740 , \14741 );
and \U$14490 ( \14743 , \14739 , \12957 );
nor \U$14491 ( \14744 , \14742 , \14743 );
not \U$14492 ( \14745 , \14744 );
not \U$14493 ( \14746 , \14745 );
or \U$14494 ( \14747 , \14734 , \14746 );
nand \U$14495 ( \14748 , \14744 , \14732 );
nand \U$14496 ( \14749 , \14747 , \14748 );
not \U$14497 ( \14750 , RIbe2a3e8_88);
not \U$14498 ( \14751 , \10937 );
not \U$14499 ( \14752 , \14751 );
or \U$14500 ( \14753 , \14750 , \14752 );
nand \U$14501 ( \14754 , \12213 , RIbe2a370_87);
nand \U$14502 ( \14755 , \14753 , \14754 );
buf \U$14503 ( \14756 , \13030 );
not \U$14504 ( \14757 , \14756 );
and \U$14505 ( \14758 , \14755 , \14757 );
not \U$14506 ( \14759 , \14755 );
and \U$14507 ( \14760 , \14759 , \12218 );
nor \U$14508 ( \14761 , \14758 , \14760 );
not \U$14509 ( \14762 , \14761 );
and \U$14510 ( \14763 , \14749 , \14762 );
not \U$14511 ( \14764 , \14749 );
and \U$14512 ( \14765 , \14764 , \14761 );
nor \U$14513 ( \14766 , \14763 , \14765 );
not \U$14514 ( \14767 , \14766 );
not \U$14515 ( \14768 , \14767 );
and \U$14516 ( \14769 , \10915 , RIbe2a910_99);
not \U$14517 ( \14770 , \13038 );
not \U$14518 ( \14771 , \14770 );
and \U$14519 ( \14772 , \14771 , RIbe2b5b8_126);
nor \U$14520 ( \14773 , \14769 , \14772 );
and \U$14521 ( \14774 , \14773 , \13383 );
not \U$14522 ( \14775 , \14773 );
and \U$14523 ( \14776 , \14775 , \13148 );
nor \U$14524 ( \14777 , \14774 , \14776 );
not \U$14525 ( \14778 , \14777 );
not \U$14526 ( \14779 , \14778 );
not \U$14527 ( \14780 , RIbe2a550_91);
not \U$14528 ( \14781 , \7975 );
or \U$14529 ( \14782 , \14780 , \14781 );
nand \U$14530 ( \14783 , \7981 , RIbe2a988_100);
nand \U$14531 ( \14784 , \14782 , \14783 );
and \U$14532 ( \14785 , \14784 , \7984 );
not \U$14533 ( \14786 , \14784 );
and \U$14534 ( \14787 , \14786 , \9896 );
nor \U$14535 ( \14788 , \14785 , \14787 );
not \U$14536 ( \14789 , \14788 );
not \U$14537 ( \14790 , \14789 );
or \U$14538 ( \14791 , \14779 , \14790 );
nand \U$14539 ( \14792 , \14788 , \14777 );
nand \U$14540 ( \14793 , \14791 , \14792 );
not \U$14541 ( \14794 , \7301 );
not \U$14542 ( \14795 , RIbe2a190_83);
not \U$14543 ( \14796 , \7299 );
or \U$14544 ( \14797 , \14795 , \14796 );
nand \U$14545 ( \14798 , \6985 , RIbe2a5c8_92);
nand \U$14546 ( \14799 , \14797 , \14798 );
not \U$14547 ( \14800 , \14799 );
or \U$14548 ( \14801 , \14794 , \14800 );
or \U$14549 ( \14802 , \14799 , \7661 );
nand \U$14550 ( \14803 , \14801 , \14802 );
xor \U$14551 ( \14804 , \14793 , \14803 );
not \U$14552 ( \14805 , \14804 );
not \U$14553 ( \14806 , \14805 );
or \U$14554 ( \14807 , \14768 , \14806 );
nand \U$14555 ( \14808 , \14804 , \14766 );
nand \U$14556 ( \14809 , \14807 , \14808 );
not \U$14557 ( \14810 , RIbe28f48_44);
not \U$14558 ( \14811 , \13590 );
or \U$14559 ( \14812 , \14810 , \14811 );
nand \U$14560 ( \14813 , \13012 , RIbe28ed0_43);
nand \U$14561 ( \14814 , \14812 , \14813 );
not \U$14562 ( \14815 , \13705 );
and \U$14563 ( \14816 , \14814 , \14815 );
not \U$14564 ( \14817 , \14814 );
and \U$14565 ( \14818 , \14817 , \12866 );
nor \U$14566 ( \14819 , \14816 , \14818 );
not \U$14567 ( \14820 , \14819 );
not \U$14568 ( \14821 , RIbe29c68_72);
not \U$14569 ( \14822 , \12847 );
or \U$14570 ( \14823 , \14821 , \14822 );
nand \U$14571 ( \14824 , \13077 , RIbe29bf0_71);
nand \U$14572 ( \14825 , \14823 , \14824 );
and \U$14573 ( \14826 , \14825 , \12742 );
not \U$14574 ( \14827 , \14825 );
and \U$14575 ( \14828 , \14827 , \12852 );
nor \U$14576 ( \14829 , \14826 , \14828 );
not \U$14577 ( \14830 , \14829 );
not \U$14578 ( \14831 , \14830 );
or \U$14579 ( \14832 , \14820 , \14831 );
not \U$14580 ( \14833 , \14819 );
nand \U$14581 ( \14834 , \14833 , \14829 );
nand \U$14582 ( \14835 , \14832 , \14834 );
not \U$14583 ( \14836 , RIbe29e48_76);
not \U$14584 ( \14837 , \13063 );
or \U$14585 ( \14838 , \14836 , \14837 );
nand \U$14586 ( \14839 , \13728 , RIbe29dd0_75);
nand \U$14587 ( \14840 , \14838 , \14839 );
and \U$14588 ( \14841 , \14840 , \12723 );
not \U$14589 ( \14842 , \14840 );
and \U$14590 ( \14843 , \14842 , \12716 );
nor \U$14591 ( \14844 , \14841 , \14843 );
xnor \U$14592 ( \14845 , \14835 , \14844 );
and \U$14593 ( \14846 , \14809 , \14845 );
not \U$14594 ( \14847 , \14809 );
not \U$14595 ( \14848 , \14845 );
and \U$14596 ( \14849 , \14847 , \14848 );
nor \U$14597 ( \14850 , \14846 , \14849 );
xor \U$14598 ( \14851 , \14351 , \14383 );
and \U$14599 ( \14852 , \14851 , \14412 );
and \U$14600 ( \14853 , \14351 , \14383 );
or \U$14601 ( \14854 , \14852 , \14853 );
not \U$14602 ( \14855 , \14854 );
not \U$14603 ( \14856 , RIbe27e68_8);
not \U$14604 ( \14857 , \12811 );
or \U$14605 ( \14858 , \14856 , \14857 );
nand \U$14606 ( \14859 , RIbe28660_25, RIbe2ae38_110);
nand \U$14607 ( \14860 , \14858 , \14859 );
xor \U$14608 ( \14861 , \14860 , RIbe2aeb0_111);
and \U$14609 ( \14862 , \14861 , \4323 );
not \U$14610 ( \14863 , \14861 );
and \U$14611 ( \14864 , \14863 , \4603 );
nor \U$14612 ( \14865 , \14862 , \14864 );
not \U$14613 ( \14866 , \14865 );
not \U$14614 ( \14867 , RIbe27fd0_11);
not \U$14615 ( \14868 , \12887 );
or \U$14616 ( \14869 , \14867 , \14868 );
nand \U$14617 ( \14870 , \12890 , RIbe27f58_10);
nand \U$14618 ( \14871 , \14869 , \14870 );
and \U$14619 ( \14872 , \14871 , \12804 );
not \U$14620 ( \14873 , \14871 );
and \U$14621 ( \14874 , \14873 , \12801 );
nor \U$14622 ( \14875 , \14872 , \14874 );
not \U$14623 ( \14876 , \14875 );
or \U$14624 ( \14877 , \14866 , \14876 );
or \U$14625 ( \14878 , \14875 , \14865 );
nand \U$14626 ( \14879 , \14877 , \14878 );
not \U$14627 ( \14880 , \14879 );
and \U$14628 ( \14881 , \14855 , \14880 );
and \U$14629 ( \14882 , \14854 , \14879 );
nor \U$14630 ( \14883 , \14881 , \14882 );
xnor \U$14631 ( \14884 , \14850 , \14883 );
not \U$14632 ( \14885 , \14137 );
not \U$14633 ( \14886 , \14141 );
or \U$14634 ( \14887 , \14885 , \14886 );
nand \U$14635 ( \14888 , \14887 , \14149 );
not \U$14636 ( \14889 , \14137 );
nand \U$14637 ( \14890 , \14889 , \14142 );
nand \U$14638 ( \14891 , \14888 , \14890 );
xor \U$14639 ( \14892 , \14884 , \14891 );
xor \U$14640 ( \14893 , \14194 , \14225 );
and \U$14641 ( \14894 , \14893 , \14442 );
and \U$14642 ( \14895 , \14194 , \14225 );
or \U$14643 ( \14896 , \14894 , \14895 );
xor \U$14644 ( \14897 , \14892 , \14896 );
not \U$14645 ( \14898 , \14246 );
nand \U$14646 ( \14899 , \14319 , \14898 );
and \U$14647 ( \14900 , \14899 , \14282 );
nor \U$14648 ( \14901 , \14319 , \14898 );
nor \U$14649 ( \14902 , \14900 , \14901 );
not \U$14650 ( \14903 , \14902 );
and \U$14651 ( \14904 , \14176 , \14185 );
nor \U$14652 ( \14905 , \14904 , \14193 );
nor \U$14653 ( \14906 , \14176 , \14185 );
nor \U$14654 ( \14907 , \14905 , \14906 );
not \U$14655 ( \14908 , \14907 );
not \U$14656 ( \14909 , \14427 );
not \U$14657 ( \14910 , \14435 );
or \U$14658 ( \14911 , \14909 , \14910 );
nand \U$14659 ( \14912 , \14911 , \14418 );
or \U$14660 ( \14913 , \14435 , \14427 );
nand \U$14661 ( \14914 , \14912 , \14913 );
not \U$14662 ( \14915 , \14914 );
or \U$14663 ( \14916 , \14908 , \14915 );
or \U$14664 ( \14917 , \14914 , \14907 );
nand \U$14665 ( \14918 , \14916 , \14917 );
not \U$14666 ( \14919 , \14918 );
or \U$14667 ( \14920 , \14903 , \14919 );
or \U$14668 ( \14921 , \14918 , \14902 );
nand \U$14669 ( \14922 , \14920 , \14921 );
not \U$14670 ( \14923 , \14216 );
not \U$14671 ( \14924 , \14208 );
not \U$14672 ( \14925 , \14924 );
or \U$14673 ( \14926 , \14923 , \14925 );
not \U$14674 ( \14927 , \14217 );
not \U$14675 ( \14928 , \14208 );
or \U$14676 ( \14929 , \14927 , \14928 );
nand \U$14677 ( \14930 , \14929 , \14202 );
nand \U$14678 ( \14931 , \14926 , \14930 );
not \U$14679 ( \14932 , \14436 );
not \U$14680 ( \14933 , \14413 );
or \U$14681 ( \14934 , \14932 , \14933 );
nand \U$14682 ( \14935 , \14934 , \14320 );
not \U$14683 ( \14936 , \14413 );
nand \U$14684 ( \14937 , \14936 , \14439 );
nand \U$14685 ( \14938 , \14935 , \14937 );
xor \U$14686 ( \14939 , \14931 , \14938 );
or \U$14687 ( \14940 , \14281 , \14269 );
nand \U$14688 ( \14941 , \14940 , \14256 );
nand \U$14689 ( \14942 , \14269 , \14281 );
nand \U$14690 ( \14943 , \14941 , \14942 );
and \U$14691 ( \14944 , \14245 , \14235 );
xor \U$14692 ( \14945 , \14943 , \14944 );
or \U$14693 ( \14946 , \14304 , \14318 );
nand \U$14694 ( \14947 , \14946 , \14292 );
nand \U$14695 ( \14948 , \14304 , \14318 );
nand \U$14696 ( \14949 , \14947 , \14948 );
xor \U$14697 ( \14950 , \14945 , \14949 );
not \U$14698 ( \14951 , \14326 );
not \U$14699 ( \14952 , \14340 );
or \U$14700 ( \14953 , \14951 , \14952 );
or \U$14701 ( \14954 , \14326 , \14340 );
nand \U$14702 ( \14955 , \14954 , \14350 );
nand \U$14703 ( \14956 , \14953 , \14955 );
or \U$14704 ( \14957 , \14362 , \14371 );
and \U$14705 ( \14958 , \14957 , \14382 );
and \U$14706 ( \14959 , \14362 , \14371 );
nor \U$14707 ( \14960 , \14958 , \14959 );
not \U$14708 ( \14961 , \14960 );
xor \U$14709 ( \14962 , \14956 , \14961 );
not \U$14710 ( \14963 , \14394 );
or \U$14711 ( \14964 , \14963 , \14411 );
nand \U$14712 ( \14965 , \14964 , \14403 );
nand \U$14713 ( \14966 , \14411 , \14963 );
nand \U$14714 ( \14967 , \14965 , \14966 );
xor \U$14715 ( \14968 , \14962 , \14967 );
xor \U$14716 ( \14969 , \14950 , \14968 );
nand \U$14717 ( \14970 , \4809 , RIbe2ab68_104);
and \U$14718 ( \14971 , \14970 , \4323 );
not \U$14719 ( \14972 , \14970 );
and \U$14720 ( \14973 , \14972 , \4603 );
or \U$14721 ( \14974 , \14971 , \14973 );
not \U$14722 ( \14975 , RIbe2b180_117);
not \U$14723 ( \14976 , \6535 );
or \U$14724 ( \14977 , \14975 , \14976 );
nand \U$14725 ( \14978 , \7076 , RIbe2b270_119);
nand \U$14726 ( \14979 , \14977 , \14978 );
and \U$14727 ( \14980 , \14979 , \6546 );
not \U$14728 ( \14981 , \14979 );
and \U$14729 ( \14982 , \14981 , \6888 );
nor \U$14730 ( \14983 , \14980 , \14982 );
not \U$14731 ( \14984 , RIbe2b108_116);
not \U$14732 ( \14985 , \7274 );
or \U$14733 ( \14986 , \14984 , \14985 );
nand \U$14734 ( \14987 , \7278 , RIbe2b090_115);
nand \U$14735 ( \14988 , \14986 , \14987 );
and \U$14736 ( \14989 , \14988 , \6582 );
not \U$14737 ( \14990 , \14988 );
not \U$14738 ( \14991 , \7948 );
and \U$14739 ( \14992 , \14990 , \14991 );
nor \U$14740 ( \14993 , \14989 , \14992 );
xor \U$14741 ( \14994 , \14983 , \14993 );
not \U$14742 ( \14995 , RIbe2a280_85);
not \U$14743 ( \14996 , \13327 );
or \U$14744 ( \14997 , \14995 , \14996 );
not \U$14745 ( \14998 , \13156 );
nand \U$14746 ( \14999 , \14998 , \6963 );
nand \U$14747 ( \15000 , \14997 , \14999 );
and \U$14748 ( \15001 , \15000 , \7293 );
not \U$14749 ( \15002 , \15000 );
and \U$14750 ( \15003 , \15002 , \6572 );
nor \U$14751 ( \15004 , \15001 , \15003 );
xor \U$14752 ( \15005 , \14994 , \15004 );
xor \U$14753 ( \15006 , \14974 , \15005 );
not \U$14754 ( \15007 , RIbe2af28_112);
not \U$14755 ( \15008 , \6139 );
or \U$14756 ( \15009 , \15007 , \15008 );
nand \U$14757 ( \15010 , \7528 , RIbe2b1f8_118);
nand \U$14758 ( \15011 , \15009 , \15010 );
not \U$14759 ( \15012 , \15011 );
not \U$14760 ( \15013 , \5740 );
and \U$14761 ( \15014 , \15012 , \15013 );
and \U$14762 ( \15015 , \15011 , \7535 );
nor \U$14763 ( \15016 , \15014 , \15015 );
not \U$14764 ( \15017 , RIbe2b018_114);
not \U$14765 ( \15018 , \5455 );
or \U$14766 ( \15019 , \15017 , \15018 );
nand \U$14767 ( \15020 , \8247 , RIbe2afa0_113);
nand \U$14768 ( \15021 , \15019 , \15020 );
and \U$14769 ( \15022 , \15021 , \10272 );
not \U$14770 ( \15023 , \15021 );
and \U$14771 ( \15024 , \15023 , \6637 );
nor \U$14772 ( \15025 , \15022 , \15024 );
xor \U$14773 ( \15026 , \15016 , \15025 );
not \U$14774 ( \15027 , RIbe2aaf0_103);
not \U$14775 ( \15028 , \5727 );
or \U$14776 ( \15029 , \15027 , \15028 );
nand \U$14777 ( \15030 , \5052 , RIbe2b630_127);
nand \U$14778 ( \15031 , \15029 , \15030 );
and \U$14779 ( \15032 , \15031 , \4592 );
not \U$14780 ( \15033 , \15031 );
and \U$14781 ( \15034 , \15033 , \4586 );
nor \U$14782 ( \15035 , \15032 , \15034 );
xor \U$14783 ( \15036 , \15026 , \15035 );
xnor \U$14784 ( \15037 , \15006 , \15036 );
xor \U$14785 ( \15038 , \14969 , \15037 );
xor \U$14786 ( \15039 , \14939 , \15038 );
xor \U$14787 ( \15040 , \14922 , \15039 );
xor \U$14788 ( \15041 , \14897 , \15040 );
not \U$14789 ( \15042 , \14167 );
not \U$14790 ( \15043 , \14162 );
not \U$14791 ( \15044 , \15043 );
or \U$14792 ( \15045 , \15042 , \15044 );
nand \U$14793 ( \15046 , \15045 , \14443 );
not \U$14794 ( \15047 , \14167 );
nand \U$14795 ( \15048 , \15047 , \14162 );
nand \U$14796 ( \15049 , \15046 , \15048 );
and \U$14797 ( \15050 , \15041 , \15049 );
and \U$14798 ( \15051 , \14897 , \15040 );
or \U$14799 ( \15052 , \15050 , \15051 );
xor \U$14800 ( \15053 , \14884 , \14891 );
and \U$14801 ( \15054 , \15053 , \14896 );
and \U$14802 ( \15055 , \14884 , \14891 );
or \U$14803 ( \15056 , \15054 , \15055 );
and \U$14804 ( \15057 , \14922 , \15039 );
xor \U$14805 ( \15058 , \15056 , \15057 );
xor \U$14806 ( \15059 , \14931 , \14938 );
and \U$14807 ( \15060 , \15059 , \15038 );
and \U$14808 ( \15061 , \14931 , \14938 );
or \U$14809 ( \15062 , \15060 , \15061 );
not \U$14810 ( \15063 , \14907 );
not \U$14811 ( \15064 , \14902 );
or \U$14812 ( \15065 , \15063 , \15064 );
nand \U$14813 ( \15066 , \15065 , \14914 );
or \U$14814 ( \15067 , \14907 , \14902 );
nand \U$14815 ( \15068 , \15066 , \15067 );
not \U$14816 ( \15069 , \14850 );
not \U$14817 ( \15070 , \14879 );
nand \U$14818 ( \15071 , \15070 , \14854 );
not \U$14819 ( \15072 , \15071 );
or \U$14820 ( \15073 , \15069 , \15072 );
not \U$14821 ( \15074 , \14854 );
nand \U$14822 ( \15075 , \15074 , \14879 );
nand \U$14823 ( \15076 , \15073 , \15075 );
xor \U$14824 ( \15077 , \15068 , \15076 );
xor \U$14825 ( \15078 , \14950 , \14968 );
and \U$14826 ( \15079 , \15078 , \15037 );
and \U$14827 ( \15080 , \14950 , \14968 );
or \U$14828 ( \15081 , \15079 , \15080 );
xor \U$14829 ( \15082 , \15077 , \15081 );
xor \U$14830 ( \15083 , \15062 , \15082 );
not \U$14831 ( \15084 , \14956 );
nand \U$14832 ( \15085 , \15084 , \14960 );
not \U$14833 ( \15086 , \15085 );
not \U$14834 ( \15087 , \14967 );
or \U$14835 ( \15088 , \15086 , \15087 );
nand \U$14836 ( \15089 , \14961 , \14956 );
nand \U$14837 ( \15090 , \15088 , \15089 );
xor \U$14838 ( \15091 , \14943 , \14944 );
and \U$14839 ( \15092 , \15091 , \14949 );
and \U$14840 ( \15093 , \14943 , \14944 );
or \U$14841 ( \15094 , \15092 , \15093 );
xor \U$14842 ( \15095 , \15090 , \15094 );
not \U$14843 ( \15096 , \15036 );
and \U$14844 ( \15097 , \15096 , \14974 );
not \U$14845 ( \15098 , \15005 );
nor \U$14846 ( \15099 , \15097 , \15098 );
nor \U$14847 ( \15100 , \15096 , \14974 );
nor \U$14848 ( \15101 , \15099 , \15100 );
not \U$14849 ( \15102 , \15101 );
and \U$14850 ( \15103 , \15095 , \15102 );
not \U$14851 ( \15104 , \15095 );
and \U$14852 ( \15105 , \15104 , \15101 );
nor \U$14853 ( \15106 , \15103 , \15105 );
nand \U$14854 ( \15107 , \14844 , \14819 );
and \U$14855 ( \15108 , \15107 , \14830 );
nor \U$14856 ( \15109 , \14844 , \14819 );
nor \U$14857 ( \15110 , \15108 , \15109 );
not \U$14858 ( \15111 , \14861 );
nand \U$14859 ( \15112 , \15111 , \4323 );
and \U$14860 ( \15113 , \14875 , \15112 );
nor \U$14861 ( \15114 , \15111 , \4323 );
nor \U$14862 ( \15115 , \15113 , \15114 );
not \U$14863 ( \15116 , \15115 );
not \U$14864 ( \15117 , \14732 );
not \U$14865 ( \15118 , \14761 );
or \U$14866 ( \15119 , \15117 , \15118 );
or \U$14867 ( \15120 , \14761 , \14732 );
nand \U$14868 ( \15121 , \15120 , \14745 );
nand \U$14869 ( \15122 , \15119 , \15121 );
not \U$14870 ( \15123 , \15122 );
or \U$14871 ( \15124 , \15116 , \15123 );
or \U$14872 ( \15125 , \15122 , \15115 );
nand \U$14873 ( \15126 , \15124 , \15125 );
xnor \U$14874 ( \15127 , \15110 , \15126 );
not \U$14875 ( \15128 , \15127 );
xor \U$14876 ( \15129 , \14983 , \14993 );
and \U$14877 ( \15130 , \15129 , \15004 );
and \U$14878 ( \15131 , \14983 , \14993 );
or \U$14879 ( \15132 , \15130 , \15131 );
nand \U$14880 ( \15133 , \14788 , \14778 );
and \U$14881 ( \15134 , \15133 , \14803 );
nor \U$14882 ( \15135 , \14788 , \14778 );
nor \U$14883 ( \15136 , \15134 , \15135 );
and \U$14884 ( \15137 , \15132 , \15136 );
not \U$14885 ( \15138 , \15132 );
not \U$14886 ( \15139 , \15136 );
and \U$14887 ( \15140 , \15138 , \15139 );
or \U$14888 ( \15141 , \15137 , \15140 );
nand \U$14889 ( \15142 , \15035 , \15016 );
and \U$14890 ( \15143 , \15142 , \15025 );
nor \U$14891 ( \15144 , \15035 , \15016 );
nor \U$14892 ( \15145 , \15143 , \15144 );
and \U$14893 ( \15146 , \15141 , \15145 );
not \U$14894 ( \15147 , \15141 );
not \U$14895 ( \15148 , \15145 );
and \U$14896 ( \15149 , \15147 , \15148 );
nor \U$14897 ( \15150 , \15146 , \15149 );
not \U$14898 ( \15151 , \15150 );
or \U$14899 ( \15152 , \15128 , \15151 );
or \U$14900 ( \15153 , \15150 , \15127 );
nand \U$14901 ( \15154 , \15152 , \15153 );
xor \U$14902 ( \15155 , \15106 , \15154 );
or \U$14903 ( \15156 , \14845 , \14804 );
nand \U$14904 ( \15157 , \15156 , \14767 );
nand \U$14905 ( \15158 , \14804 , \14845 );
nand \U$14906 ( \15159 , \15157 , \15158 );
not \U$14907 ( \15160 , RIbe29bf0_71);
not \U$14908 ( \15161 , \12731 );
not \U$14909 ( \15162 , \15161 );
or \U$14910 ( \15163 , \15160 , \15162 );
nand \U$14911 ( \15164 , RIbe28f48_44, \12735 );
nand \U$14912 ( \15165 , \15163 , \15164 );
not \U$14913 ( \15166 , \12746 );
and \U$14914 ( \15167 , \15165 , \15166 );
not \U$14915 ( \15168 , \15165 );
not \U$14916 ( \15169 , \14358 );
and \U$14917 ( \15170 , \15168 , \15169 );
nor \U$14918 ( \15171 , \15167 , \15170 );
not \U$14919 ( \15172 , \15171 );
not \U$14920 ( \15173 , \15172 );
not \U$14921 ( \15174 , RIbe29dd0_75);
not \U$14922 ( \15175 , \12871 );
or \U$14923 ( \15176 , \15174 , \15175 );
nand \U$14924 ( \15177 , \12711 , RIbe29c68_72);
nand \U$14925 ( \15178 , \15176 , \15177 );
and \U$14926 ( \15179 , \15178 , \12723 );
not \U$14927 ( \15180 , \15178 );
and \U$14928 ( \15181 , \15180 , \12716 );
nor \U$14929 ( \15182 , \15179 , \15181 );
not \U$14930 ( \15183 , \15182 );
not \U$14931 ( \15184 , \15183 );
or \U$14932 ( \15185 , \15173 , \15184 );
nand \U$14933 ( \15186 , \15171 , \15182 );
nand \U$14934 ( \15187 , \15185 , \15186 );
not \U$14935 ( \15188 , \12753 );
not \U$14936 ( \15189 , \12380 );
and \U$14937 ( \15190 , \15188 , \15189 );
and \U$14938 ( \15191 , \14726 , RIbe29fb0_79);
nor \U$14939 ( \15192 , \15190 , \15191 );
and \U$14940 ( \15193 , \15192 , \12924 );
not \U$14941 ( \15194 , \15192 );
and \U$14942 ( \15195 , \15194 , \12774 );
nor \U$14943 ( \15196 , \15193 , \15195 );
not \U$14944 ( \15197 , \15196 );
and \U$14945 ( \15198 , \15187 , \15197 );
not \U$14946 ( \15199 , \15187 );
and \U$14947 ( \15200 , \15199 , \15196 );
nor \U$14948 ( \15201 , \15198 , \15200 );
not \U$14949 ( \15202 , \14397 );
not \U$14950 ( \15203 , \14374 );
and \U$14951 ( \15204 , \15202 , \15203 );
buf \U$14952 ( \15205 , \12941 );
and \U$14953 ( \15206 , \15205 , RIbe2acd0_107);
nor \U$14954 ( \15207 , \15204 , \15206 );
and \U$14955 ( \15208 , \15207 , \12956 );
not \U$14956 ( \15209 , \15207 );
and \U$14957 ( \15210 , \15209 , \12195 );
nor \U$14958 ( \15211 , \15208 , \15210 );
not \U$14959 ( \15212 , \15211 );
not \U$14960 ( \15213 , RIbe2a370_87);
not \U$14961 ( \15214 , \10936 );
or \U$14962 ( \15215 , \15213 , \15214 );
nand \U$14963 ( \15216 , \12213 , RIbe2a2f8_86);
nand \U$14964 ( \15217 , \15215 , \15216 );
not \U$14965 ( \15218 , \15217 );
not \U$14966 ( \15219 , \13030 );
and \U$14967 ( \15220 , \15218 , \15219 );
and \U$14968 ( \15221 , \15217 , \13661 );
nor \U$14969 ( \15222 , \15220 , \15221 );
not \U$14970 ( \15223 , \15222 );
or \U$14971 ( \15224 , \15212 , \15223 );
or \U$14972 ( \15225 , \15222 , \15211 );
nand \U$14973 ( \15226 , \15224 , \15225 );
and \U$14974 ( \15227 , \10916 , RIbe2b5b8_126);
not \U$14975 ( \15228 , \13039 );
and \U$14976 ( \15229 , \15228 , RIbe2a3e8_88);
nor \U$14977 ( \15230 , \15227 , \15229 );
and \U$14978 ( \15231 , \15230 , \10926 );
not \U$14979 ( \15232 , \15230 );
not \U$14980 ( \15233 , \7970 );
and \U$14981 ( \15234 , \15232 , \15233 );
nor \U$14982 ( \15235 , \15231 , \15234 );
not \U$14983 ( \15236 , \15235 );
and \U$14984 ( \15237 , \15226 , \15236 );
not \U$14985 ( \15238 , \15226 );
and \U$14986 ( \15239 , \15238 , \15235 );
nor \U$14987 ( \15240 , \15237 , \15239 );
xor \U$14988 ( \15241 , \15201 , \15240 );
not \U$14989 ( \15242 , RIbe28660_25);
not \U$14990 ( \15243 , \13690 );
or \U$14991 ( \15244 , \15242 , \15243 );
nand \U$14992 ( \15245 , RIbe285e8_24, RIbe2ae38_110);
nand \U$14993 ( \15246 , \15244 , \15245 );
xnor \U$14994 ( \15247 , \15246 , RIbe2aeb0_111);
not \U$14995 ( \15248 , RIbe27f58_10);
and \U$14996 ( \15249 , \12782 , \12784 );
buf \U$14997 ( \15250 , \15249 );
not \U$14998 ( \15251 , \15250 );
or \U$14999 ( \15252 , \15248 , \15251 );
nand \U$15000 ( \15253 , RIbe27e68_8, \12890 );
nand \U$15001 ( \15254 , \15252 , \15253 );
xor \U$15002 ( \15255 , \15254 , \12893 );
xor \U$15003 ( \15256 , \15247 , \15255 );
not \U$15004 ( \15257 , RIbe28ed0_43);
not \U$15005 ( \15258 , \13590 );
or \U$15006 ( \15259 , \15257 , \15258 );
nand \U$15007 ( \15260 , \12835 , RIbe27fd0_11);
nand \U$15008 ( \15261 , \15259 , \15260 );
not \U$15009 ( \15262 , \15261 );
not \U$15010 ( \15263 , \13595 );
not \U$15011 ( \15264 , \15263 );
and \U$15012 ( \15265 , \15262 , \15264 );
and \U$15013 ( \15266 , \15261 , \12823 );
nor \U$15014 ( \15267 , \15265 , \15266 );
xor \U$15015 ( \15268 , \15256 , \15267 );
xor \U$15016 ( \15269 , \15241 , \15268 );
xor \U$15017 ( \15270 , \15159 , \15269 );
not \U$15018 ( \15271 , \6888 );
not \U$15019 ( \15272 , RIbe2b270_119);
not \U$15020 ( \15273 , \6535 );
or \U$15021 ( \15274 , \15272 , \15273 );
nand \U$15022 ( \15275 , \10348 , RIbe2b108_116);
nand \U$15023 ( \15276 , \15274 , \15275 );
not \U$15024 ( \15277 , \15276 );
or \U$15025 ( \15278 , \15271 , \15277 );
or \U$15026 ( \15279 , \6548 , \15276 );
nand \U$15027 ( \15280 , \15278 , \15279 );
not \U$15028 ( \15281 , \6602 );
not \U$15029 ( \15282 , RIbe2b090_115);
not \U$15030 ( \15283 , \13238 );
or \U$15031 ( \15284 , \15282 , \15283 );
nand \U$15032 ( \15285 , \6596 , RIbe2a280_85);
nand \U$15033 ( \15286 , \15284 , \15285 );
not \U$15034 ( \15287 , \15286 );
or \U$15035 ( \15288 , \15281 , \15287 );
or \U$15036 ( \15289 , \15286 , \6583 );
nand \U$15037 ( \15290 , \15288 , \15289 );
xor \U$15038 ( \15291 , \15280 , \15290 );
not \U$15039 ( \15292 , \9944 );
not \U$15040 ( \15293 , RIbe2b1f8_118);
not \U$15041 ( \15294 , \6139 );
or \U$15042 ( \15295 , \15293 , \15294 );
nand \U$15043 ( \15296 , \8235 , RIbe2b180_117);
nand \U$15044 ( \15297 , \15295 , \15296 );
not \U$15045 ( \15298 , \15297 );
or \U$15046 ( \15299 , \15292 , \15298 );
or \U$15047 ( \15300 , \15297 , \6624 );
nand \U$15048 ( \15301 , \15299 , \15300 );
xor \U$15049 ( \15302 , \15291 , \15301 );
not \U$15050 ( \15303 , RIbe2b630_127);
not \U$15051 ( \15304 , \6427 );
or \U$15052 ( \15305 , \15303 , \15304 );
nand \U$15053 ( \15306 , RIbe2b018_114, \7056 );
nand \U$15054 ( \15307 , \15305 , \15306 );
and \U$15055 ( \15308 , \15307 , \4586 );
not \U$15056 ( \15309 , \15307 );
and \U$15057 ( \15310 , \15309 , \4592 );
nor \U$15058 ( \15311 , \15308 , \15310 );
not \U$15059 ( \15312 , RIbe2afa0_113);
not \U$15060 ( \15313 , \6629 );
not \U$15061 ( \15314 , \15313 );
or \U$15062 ( \15315 , \15312 , \15314 );
nand \U$15063 ( \15316 , \6634 , RIbe2af28_112);
nand \U$15064 ( \15317 , \15315 , \15316 );
xor \U$15065 ( \15318 , \15317 , \6640 );
and \U$15066 ( \15319 , \15311 , \15318 );
not \U$15067 ( \15320 , \15311 );
not \U$15068 ( \15321 , \15318 );
and \U$15069 ( \15322 , \15320 , \15321 );
nor \U$15070 ( \15323 , \15319 , \15322 );
not \U$15071 ( \15324 , RIbe2ab68_104);
not \U$15072 ( \15325 , \6414 );
or \U$15073 ( \15326 , \15324 , \15325 );
nand \U$15074 ( \15327 , \4600 , RIbe2aaf0_103);
nand \U$15075 ( \15328 , \15326 , \15327 );
and \U$15076 ( \15329 , \15328 , \4326 );
not \U$15077 ( \15330 , \15328 );
and \U$15078 ( \15331 , \15330 , \4323 );
nor \U$15079 ( \15332 , \15329 , \15331 );
xor \U$15080 ( \15333 , \15323 , \15332 );
xor \U$15081 ( \15334 , \15302 , \15333 );
not \U$15082 ( \15335 , RIbe2a5c8_92);
not \U$15083 ( \15336 , \7298 );
or \U$15084 ( \15337 , \15335 , \15336 );
nand \U$15085 ( \15338 , \12251 , RIbe2a550_91);
nand \U$15086 ( \15339 , \15337 , \15338 );
not \U$15087 ( \15340 , \15339 );
not \U$15088 ( \15341 , \6992 );
and \U$15089 ( \15342 , \15340 , \15341 );
and \U$15090 ( \15343 , \15339 , \10902 );
nor \U$15091 ( \15344 , \15342 , \15343 );
not \U$15092 ( \15345 , \15344 );
not \U$15093 ( \15346 , RIbe2a988_100);
not \U$15094 ( \15347 , \10949 );
or \U$15095 ( \15348 , \15346 , \15347 );
nand \U$15096 ( \15349 , \9891 , RIbe2a910_99);
nand \U$15097 ( \15350 , \15348 , \15349 );
and \U$15098 ( \15351 , \15350 , \12234 );
not \U$15099 ( \15352 , \15350 );
and \U$15100 ( \15353 , \15352 , \7984 );
nor \U$15101 ( \15354 , \15351 , \15353 );
not \U$15102 ( \15355 , \15354 );
or \U$15103 ( \15356 , \15345 , \15355 );
or \U$15104 ( \15357 , \15354 , \15344 );
nand \U$15105 ( \15358 , \15356 , \15357 );
not \U$15106 ( \15359 , RIbe2a208_84);
not \U$15107 ( \15360 , \13327 );
or \U$15108 ( \15361 , \15359 , \15360 );
nand \U$15109 ( \15362 , \6963 , RIbe2a190_83);
nand \U$15110 ( \15363 , \15361 , \15362 );
and \U$15111 ( \15364 , \15363 , \7293 );
not \U$15112 ( \15365 , \15363 );
and \U$15113 ( \15366 , \15365 , \6572 );
nor \U$15114 ( \15367 , \15364 , \15366 );
buf \U$15115 ( \15368 , \15367 );
not \U$15116 ( \15369 , \15368 );
and \U$15117 ( \15370 , \15358 , \15369 );
not \U$15118 ( \15371 , \15358 );
and \U$15119 ( \15372 , \15371 , \15368 );
nor \U$15120 ( \15373 , \15370 , \15372 );
xor \U$15121 ( \15374 , \15334 , \15373 );
xor \U$15122 ( \15375 , \15270 , \15374 );
xor \U$15123 ( \15376 , \15155 , \15375 );
xor \U$15124 ( \15377 , \15083 , \15376 );
xor \U$15125 ( \15378 , \15058 , \15377 );
xnor \U$15126 ( \15379 , \15052 , \15378 );
not \U$15127 ( \15380 , \15379 );
xor \U$15128 ( \15381 , \15056 , \15057 );
and \U$15129 ( \15382 , \15381 , \15377 );
and \U$15130 ( \15383 , \15056 , \15057 );
or \U$15131 ( \15384 , \15382 , \15383 );
xor \U$15132 ( \15385 , \15159 , \15269 );
and \U$15133 ( \15386 , \15385 , \15374 );
and \U$15134 ( \15387 , \15159 , \15269 );
or \U$15135 ( \15388 , \15386 , \15387 );
or \U$15136 ( \15389 , \15094 , \15090 );
and \U$15137 ( \15390 , \15102 , \15389 );
and \U$15138 ( \15391 , \15090 , \15094 );
nor \U$15139 ( \15392 , \15390 , \15391 );
not \U$15140 ( \15393 , \15392 );
not \U$15141 ( \15394 , \15150 );
nand \U$15142 ( \15395 , \15394 , \15127 );
not \U$15143 ( \15396 , \15395 );
xor \U$15144 ( \15397 , \15393 , \15396 );
xor \U$15145 ( \15398 , \15388 , \15397 );
xor \U$15146 ( \15399 , \15062 , \15082 );
and \U$15147 ( \15400 , \15399 , \15376 );
and \U$15148 ( \15401 , \15062 , \15082 );
or \U$15149 ( \15402 , \15400 , \15401 );
xor \U$15150 ( \15403 , \15398 , \15402 );
xor \U$15151 ( \15404 , \15106 , \15154 );
and \U$15152 ( \15405 , \15404 , \15375 );
and \U$15153 ( \15406 , \15106 , \15154 );
or \U$15154 ( \15407 , \15405 , \15406 );
xor \U$15155 ( \15408 , \15068 , \15076 );
and \U$15156 ( \15409 , \15408 , \15081 );
and \U$15157 ( \15410 , \15068 , \15076 );
or \U$15158 ( \15411 , \15409 , \15410 );
xor \U$15159 ( \15412 , \15407 , \15411 );
nand \U$15160 ( \15413 , \4027 , RIbe2ab68_104);
and \U$15161 ( \15414 , \15413 , \3471 );
not \U$15162 ( \15415 , \15413 );
and \U$15163 ( \15416 , \15415 , \4821 );
nor \U$15164 ( \15417 , \15414 , \15416 );
not \U$15165 ( \15418 , RIbe2aaf0_103);
not \U$15166 ( \15419 , \4317 );
or \U$15167 ( \15420 , \15418 , \15419 );
nand \U$15168 ( \15421 , \4809 , RIbe2b630_127);
nand \U$15169 ( \15422 , \15420 , \15421 );
not \U$15170 ( \15423 , \15422 );
not \U$15171 ( \15424 , \4323 );
and \U$15172 ( \15425 , \15423 , \15424 );
and \U$15173 ( \15426 , \15422 , \4323 );
nor \U$15174 ( \15427 , \15425 , \15426 );
not \U$15175 ( \15428 , \15427 );
and \U$15176 ( \15429 , \15417 , \15428 );
not \U$15177 ( \15430 , \15417 );
and \U$15178 ( \15431 , \15430 , \15427 );
nor \U$15179 ( \15432 , \15429 , \15431 );
not \U$15180 ( \15433 , \15432 );
not \U$15181 ( \15434 , \4592 );
not \U$15182 ( \15435 , RIbe2b018_114);
not \U$15183 ( \15436 , \6427 );
or \U$15184 ( \15437 , \15435 , \15436 );
nand \U$15185 ( \15438 , \7056 , RIbe2afa0_113);
nand \U$15186 ( \15439 , \15437 , \15438 );
not \U$15187 ( \15440 , \15439 );
or \U$15188 ( \15441 , \15434 , \15440 );
or \U$15189 ( \15442 , \15439 , \4592 );
nand \U$15190 ( \15443 , \15441 , \15442 );
not \U$15191 ( \15444 , \15443 );
not \U$15192 ( \15445 , \15444 );
not \U$15193 ( \15446 , RIbe2b180_117);
not \U$15194 ( \15447 , \6138 );
or \U$15195 ( \15448 , \15446 , \15447 );
nand \U$15196 ( \15449 , \6859 , RIbe2b270_119);
nand \U$15197 ( \15450 , \15448 , \15449 );
and \U$15198 ( \15451 , \15450 , \7535 );
not \U$15199 ( \15452 , \15450 );
and \U$15200 ( \15453 , \15452 , \10969 );
nor \U$15201 ( \15454 , \15451 , \15453 );
not \U$15202 ( \15455 , \15454 );
not \U$15203 ( \15456 , \8252 );
not \U$15204 ( \15457 , RIbe2af28_112);
not \U$15205 ( \15458 , \15313 );
or \U$15206 ( \15459 , \15457 , \15458 );
nand \U$15207 ( \15460 , \7100 , RIbe2b1f8_118);
nand \U$15208 ( \15461 , \15459 , \15460 );
not \U$15209 ( \15462 , \15461 );
or \U$15210 ( \15463 , \15456 , \15462 );
or \U$15211 ( \15464 , \15461 , \6637 );
nand \U$15212 ( \15465 , \15463 , \15464 );
not \U$15213 ( \15466 , \15465 );
or \U$15214 ( \15467 , \15455 , \15466 );
or \U$15215 ( \15468 , \15454 , \15465 );
nand \U$15216 ( \15469 , \15467 , \15468 );
not \U$15217 ( \15470 , \15469 );
or \U$15218 ( \15471 , \15445 , \15470 );
or \U$15219 ( \15472 , \15469 , \15444 );
nand \U$15220 ( \15473 , \15471 , \15472 );
not \U$15221 ( \15474 , \15473 );
and \U$15222 ( \15475 , \15433 , \15474 );
and \U$15223 ( \15476 , \15473 , \15432 );
nor \U$15224 ( \15477 , \15475 , \15476 );
not \U$15225 ( \15478 , \15477 );
or \U$15226 ( \15479 , \15332 , \15311 );
nand \U$15227 ( \15480 , \15479 , \15321 );
nand \U$15228 ( \15481 , \15332 , \15311 );
nand \U$15229 ( \15482 , \15480 , \15481 );
xor \U$15230 ( \15483 , \15280 , \15290 );
and \U$15231 ( \15484 , \15483 , \15301 );
and \U$15232 ( \15485 , \15280 , \15290 );
or \U$15233 ( \15486 , \15484 , \15485 );
xor \U$15234 ( \15487 , \15482 , \15486 );
or \U$15235 ( \15488 , \15367 , \15354 );
not \U$15236 ( \15489 , \15344 );
nand \U$15237 ( \15490 , \15488 , \15489 );
nand \U$15238 ( \15491 , \15367 , \15354 );
nand \U$15239 ( \15492 , \15490 , \15491 );
xor \U$15240 ( \15493 , \15487 , \15492 );
not \U$15241 ( \15494 , \15493 );
or \U$15242 ( \15495 , \15478 , \15494 );
or \U$15243 ( \15496 , \15493 , \15477 );
nand \U$15244 ( \15497 , \15495 , \15496 );
not \U$15245 ( \15498 , \15172 );
not \U$15246 ( \15499 , \15182 );
or \U$15247 ( \15500 , \15498 , \15499 );
nand \U$15248 ( \15501 , \15500 , \15196 );
nand \U$15249 ( \15502 , \15171 , \15183 );
nand \U$15250 ( \15503 , \15501 , \15502 );
not \U$15251 ( \15504 , \15503 );
not \U$15252 ( \15505 , \15222 );
not \U$15253 ( \15506 , \15235 );
or \U$15254 ( \15507 , \15505 , \15506 );
nand \U$15255 ( \15508 , \15507 , \15211 );
not \U$15256 ( \15509 , \15222 );
nand \U$15257 ( \15510 , \15509 , \15236 );
nand \U$15258 ( \15511 , \15508 , \15510 );
not \U$15259 ( \15512 , \15511 );
not \U$15260 ( \15513 , \15512 );
or \U$15261 ( \15514 , \15504 , \15513 );
not \U$15262 ( \15515 , \15503 );
nand \U$15263 ( \15516 , \15515 , \15511 );
nand \U$15264 ( \15517 , \15514 , \15516 );
not \U$15265 ( \15518 , \15517 );
xor \U$15266 ( \15519 , \15247 , \15255 );
and \U$15267 ( \15520 , \15519 , \15267 );
and \U$15268 ( \15521 , \15247 , \15255 );
or \U$15269 ( \15522 , \15520 , \15521 );
not \U$15270 ( \15523 , \15522 );
and \U$15271 ( \15524 , \15518 , \15523 );
and \U$15272 ( \15525 , \15517 , \15522 );
nor \U$15273 ( \15526 , \15524 , \15525 );
xnor \U$15274 ( \15527 , \15497 , \15526 );
not \U$15275 ( \15528 , \15115 );
not \U$15276 ( \15529 , \15110 );
or \U$15277 ( \15530 , \15528 , \15529 );
nand \U$15278 ( \15531 , \15530 , \15122 );
or \U$15279 ( \15532 , \15110 , \15115 );
nand \U$15280 ( \15533 , \15531 , \15532 );
not \U$15281 ( \15534 , \15136 );
not \U$15282 ( \15535 , \15145 );
or \U$15283 ( \15536 , \15534 , \15535 );
nand \U$15284 ( \15537 , \15536 , \15132 );
not \U$15285 ( \15538 , \15145 );
nand \U$15286 ( \15539 , \15538 , \15139 );
nand \U$15287 ( \15540 , \15537 , \15539 );
not \U$15288 ( \15541 , \15540 );
xor \U$15289 ( \15542 , \15533 , \15541 );
nand \U$15290 ( \15543 , \15373 , \15333 );
and \U$15291 ( \15544 , \15543 , \15302 );
nor \U$15292 ( \15545 , \15373 , \15333 );
nor \U$15293 ( \15546 , \15544 , \15545 );
xor \U$15294 ( \15547 , \15542 , \15546 );
not \U$15295 ( \15548 , \15547 );
and \U$15296 ( \15549 , \15527 , \15548 );
not \U$15297 ( \15550 , \15527 );
and \U$15298 ( \15551 , \15550 , \15547 );
nor \U$15299 ( \15552 , \15549 , \15551 );
not \U$15300 ( \15553 , RIbe27fd0_11);
not \U$15301 ( \15554 , \12858 );
or \U$15302 ( \15555 , \15553 , \15554 );
nand \U$15303 ( \15556 , \13012 , RIbe27f58_10);
nand \U$15304 ( \15557 , \15555 , \15556 );
and \U$15305 ( \15558 , \15557 , \13705 );
not \U$15306 ( \15559 , \15557 );
and \U$15307 ( \15560 , \15559 , \12822 );
nor \U$15308 ( \15561 , \15558 , \15560 );
not \U$15309 ( \15562 , RIbe28f48_44);
not \U$15310 ( \15563 , \14071 );
or \U$15311 ( \15564 , \15562 , \15563 );
nand \U$15312 ( \15565 , \12735 , RIbe28ed0_43);
nand \U$15313 ( \15566 , \15564 , \15565 );
and \U$15314 ( \15567 , \15566 , \12742 );
not \U$15315 ( \15568 , \15566 );
and \U$15316 ( \15569 , \15568 , \14358 );
nor \U$15317 ( \15570 , \15567 , \15569 );
xor \U$15318 ( \15571 , \15561 , \15570 );
not \U$15319 ( \15572 , RIbe29c68_72);
not \U$15320 ( \15573 , \12706 );
not \U$15321 ( \15574 , \15573 );
or \U$15322 ( \15575 , \15572 , \15574 );
nand \U$15323 ( \15576 , \12711 , RIbe29bf0_71);
nand \U$15324 ( \15577 , \15575 , \15576 );
and \U$15325 ( \15578 , \15577 , \12723 );
not \U$15326 ( \15579 , \15577 );
and \U$15327 ( \15580 , \15579 , \13068 );
nor \U$15328 ( \15581 , \15578 , \15580 );
xor \U$15329 ( \15582 , \15571 , \15581 );
not \U$15330 ( \15583 , \15582 );
not \U$15331 ( \15584 , \15583 );
not \U$15332 ( \15585 , RIbe285e8_24);
not \U$15333 ( \15586 , \13690 );
or \U$15334 ( \15587 , \15585 , \15586 );
nand \U$15335 ( \15588 , RIbe287c8_28, RIbe2ae38_110);
nand \U$15336 ( \15589 , \15587 , \15588 );
xor \U$15337 ( \15590 , RIbe2aeb0_111, \15589 );
xor \U$15338 ( \15591 , \3471 , \15590 );
not \U$15339 ( \15592 , RIbe27e68_8);
not \U$15340 ( \15593 , \12887 );
or \U$15341 ( \15594 , \15592 , \15593 );
nand \U$15342 ( \15595 , \12890 , RIbe28660_25);
nand \U$15343 ( \15596 , \15594 , \15595 );
and \U$15344 ( \15597 , \15596 , \14103 );
not \U$15345 ( \15598 , \15596 );
and \U$15346 ( \15599 , \15598 , \12801 );
nor \U$15347 ( \15600 , \15597 , \15599 );
xor \U$15348 ( \15601 , \15591 , \15600 );
not \U$15349 ( \15602 , \15601 );
and \U$15350 ( \15603 , \15584 , \15602 );
and \U$15351 ( \15604 , \15583 , \15601 );
nor \U$15352 ( \15605 , \15603 , \15604 );
nand \U$15353 ( \15606 , \15268 , \15201 );
and \U$15354 ( \15607 , \15606 , \15240 );
nor \U$15355 ( \15608 , \15268 , \15201 );
nor \U$15356 ( \15609 , \15607 , \15608 );
xor \U$15357 ( \15610 , \15605 , \15609 );
not \U$15358 ( \15611 , \12753 );
not \U$15359 ( \15612 , RIbe29dd0_75);
not \U$15360 ( \15613 , \15612 );
and \U$15361 ( \15614 , \15611 , \15613 );
not \U$15362 ( \15615 , \12763 );
and \U$15363 ( \15616 , \15615 , RIbe29e48_76);
nor \U$15364 ( \15617 , \15614 , \15616 );
and \U$15365 ( \15618 , \15617 , \12770 );
not \U$15366 ( \15619 , \15617 );
and \U$15367 ( \15620 , \15619 , \12927 );
nor \U$15368 ( \15621 , \15618 , \15620 );
not \U$15369 ( \15622 , \15621 );
not \U$15370 ( \15623 , \15622 );
not \U$15371 ( \15624 , RIbe2a028_80);
not \U$15372 ( \15625 , \12942 );
or \U$15373 ( \15626 , \15624 , \15625 );
not \U$15374 ( \15627 , \12947 );
not \U$15375 ( \15628 , \15627 );
nand \U$15376 ( \15629 , \15628 , RIbe29fb0_79);
nand \U$15377 ( \15630 , \15626 , \15629 );
not \U$15378 ( \15631 , \15630 );
not \U$15379 ( \15632 , \12960 );
and \U$15380 ( \15633 , \15631 , \15632 );
and \U$15381 ( \15634 , \15630 , \12957 );
nor \U$15382 ( \15635 , \15633 , \15634 );
not \U$15383 ( \15636 , \15635 );
not \U$15384 ( \15637 , \15636 );
or \U$15385 ( \15638 , \15623 , \15637 );
nand \U$15386 ( \15639 , \15635 , \15621 );
nand \U$15387 ( \15640 , \15638 , \15639 );
not \U$15388 ( \15641 , RIbe2a2f8_86);
not \U$15389 ( \15642 , \10936 );
or \U$15390 ( \15643 , \15641 , \15642 );
nand \U$15391 ( \15644 , \14511 , RIbe2acd0_107);
nand \U$15392 ( \15645 , \15643 , \15644 );
not \U$15393 ( \15646 , \15645 );
not \U$15394 ( \15647 , \14756 );
and \U$15395 ( \15648 , \15646 , \15647 );
and \U$15396 ( \15649 , \15645 , \13033 );
nor \U$15397 ( \15650 , \15648 , \15649 );
and \U$15398 ( \15651 , \15640 , \15650 );
not \U$15399 ( \15652 , \15640 );
not \U$15400 ( \15653 , \15650 );
and \U$15401 ( \15654 , \15652 , \15653 );
nor \U$15402 ( \15655 , \15651 , \15654 );
not \U$15403 ( \15656 , \15655 );
not \U$15404 ( \15657 , \15656 );
and \U$15405 ( \15658 , \8276 , RIbe2a3e8_88);
and \U$15406 ( \15659 , \9914 , RIbe2a370_87);
nor \U$15407 ( \15660 , \15658 , \15659 );
and \U$15408 ( \15661 , \15660 , \15233 );
not \U$15409 ( \15662 , \15660 );
and \U$15410 ( \15663 , \15662 , \7970 );
nor \U$15411 ( \15664 , \15661 , \15663 );
not \U$15412 ( \15665 , \15664 );
not \U$15413 ( \15666 , \15665 );
not \U$15414 ( \15667 , RIbe2a910_99);
not \U$15415 ( \15668 , \7975 );
or \U$15416 ( \15669 , \15667 , \15668 );
nand \U$15417 ( \15670 , \8269 , RIbe2b5b8_126);
nand \U$15418 ( \15671 , \15669 , \15670 );
and \U$15419 ( \15672 , \15671 , \7984 );
not \U$15420 ( \15673 , \15671 );
and \U$15421 ( \15674 , \15673 , \7988 );
nor \U$15422 ( \15675 , \15672 , \15674 );
not \U$15423 ( \15676 , \15675 );
not \U$15424 ( \15677 , \15676 );
or \U$15425 ( \15678 , \15666 , \15677 );
nand \U$15426 ( \15679 , \15675 , \15664 );
nand \U$15427 ( \15680 , \15678 , \15679 );
not \U$15428 ( \15681 , RIbe2a550_91);
not \U$15429 ( \15682 , \7299 );
or \U$15430 ( \15683 , \15681 , \15682 );
nand \U$15431 ( \15684 , \9875 , RIbe2a988_100);
nand \U$15432 ( \15685 , \15683 , \15684 );
and \U$15433 ( \15686 , \15685 , \6993 );
not \U$15434 ( \15687 , \15685 );
and \U$15435 ( \15688 , \15687 , \10902 );
nor \U$15436 ( \15689 , \15686 , \15688 );
not \U$15437 ( \15690 , \15689 );
and \U$15438 ( \15691 , \15680 , \15690 );
not \U$15439 ( \15692 , \15680 );
and \U$15440 ( \15693 , \15692 , \15689 );
nor \U$15441 ( \15694 , \15691 , \15693 );
not \U$15442 ( \15695 , \15694 );
or \U$15443 ( \15696 , \15657 , \15695 );
not \U$15444 ( \15697 , \15694 );
nand \U$15445 ( \15698 , \15697 , \15655 );
nand \U$15446 ( \15699 , \15696 , \15698 );
not \U$15447 ( \15700 , RIbe2a190_83);
not \U$15448 ( \15701 , \6560 );
or \U$15449 ( \15702 , \15700 , \15701 );
nand \U$15450 ( \15703 , \8202 , RIbe2a5c8_92);
nand \U$15451 ( \15704 , \15702 , \15703 );
and \U$15452 ( \15705 , \15704 , \6569 );
not \U$15453 ( \15706 , \15704 );
and \U$15454 ( \15707 , \15706 , \7293 );
nor \U$15455 ( \15708 , \15705 , \15707 );
not \U$15456 ( \15709 , \15708 );
not \U$15457 ( \15710 , \15709 );
not \U$15458 ( \15711 , RIbe2a280_85);
not \U$15459 ( \15712 , \7941 );
or \U$15460 ( \15713 , \15711 , \15712 );
nand \U$15461 ( \15714 , \7483 , RIbe2a208_84);
nand \U$15462 ( \15715 , \15713 , \15714 );
and \U$15463 ( \15716 , \15715 , \6601 );
not \U$15464 ( \15717 , \15715 );
and \U$15465 ( \15718 , \15717 , \14991 );
nor \U$15466 ( \15719 , \15716 , \15718 );
not \U$15467 ( \15720 , \15719 );
not \U$15468 ( \15721 , \15720 );
or \U$15469 ( \15722 , \15710 , \15721 );
nand \U$15470 ( \15723 , \15708 , \15719 );
nand \U$15471 ( \15724 , \15722 , \15723 );
not \U$15472 ( \15725 , RIbe2b108_116);
not \U$15473 ( \15726 , \6536 );
or \U$15474 ( \15727 , \15725 , \15726 );
nand \U$15475 ( \15728 , \6540 , RIbe2b090_115);
nand \U$15476 ( \15729 , \15727 , \15728 );
not \U$15477 ( \15730 , \6891 );
and \U$15478 ( \15731 , \15729 , \15730 );
not \U$15479 ( \15732 , \15729 );
and \U$15480 ( \15733 , \15732 , \6548 );
nor \U$15481 ( \15734 , \15731 , \15733 );
xnor \U$15482 ( \15735 , \15724 , \15734 );
not \U$15483 ( \15736 , \15735 );
and \U$15484 ( \15737 , \15699 , \15736 );
not \U$15485 ( \15738 , \15699 );
and \U$15486 ( \15739 , \15738 , \15735 );
nor \U$15487 ( \15740 , \15737 , \15739 );
xor \U$15488 ( \15741 , \15610 , \15740 );
not \U$15489 ( \15742 , \15741 );
and \U$15490 ( \15743 , \15552 , \15742 );
not \U$15491 ( \15744 , \15552 );
and \U$15492 ( \15745 , \15744 , \15741 );
nor \U$15493 ( \15746 , \15743 , \15745 );
xor \U$15494 ( \15747 , \15412 , \15746 );
xor \U$15495 ( \15748 , \15403 , \15747 );
xor \U$15496 ( \15749 , \15384 , \15748 );
nand \U$15497 ( \15750 , \14447 , \14150 );
and \U$15498 ( \15751 , \15750 , \14154 );
nor \U$15499 ( \15752 , \14447 , \14150 );
nor \U$15500 ( \15753 , \15751 , \15752 );
not \U$15501 ( \15754 , \15753 );
not \U$15502 ( \15755 , \15754 );
xor \U$15503 ( \15756 , \14897 , \15040 );
xor \U$15504 ( \15757 , \15756 , \15049 );
not \U$15505 ( \15758 , \15757 );
not \U$15506 ( \15759 , \15758 );
or \U$15507 ( \15760 , \15755 , \15759 );
nand \U$15508 ( \15761 , \15757 , \15753 );
nand \U$15509 ( \15762 , \15760 , \15761 );
nand \U$15510 ( \15763 , \15380 , \15749 , \15762 );
nor \U$15511 ( \15764 , \14720 , \15763 );
nand \U$15512 ( \15765 , \15757 , \15754 );
nor \U$15513 ( \15766 , \15379 , \15765 );
nand \U$15514 ( \15767 , \15766 , \15749 );
and \U$15515 ( \15768 , \15378 , \15052 );
nand \U$15516 ( \15769 , \15749 , \15768 );
nand \U$15517 ( \15770 , \15767 , \15769 );
or \U$15518 ( \15771 , \15764 , \15770 );
not \U$15519 ( \15772 , RIbe28660_25);
not \U$15520 ( \15773 , \15249 );
or \U$15521 ( \15774 , \15772 , \15773 );
nand \U$15522 ( \15775 , \12794 , RIbe285e8_24);
nand \U$15523 ( \15776 , \15774 , \15775 );
and \U$15524 ( \15777 , \15776 , \12801 );
not \U$15525 ( \15778 , \15776 );
and \U$15526 ( \15779 , \15778 , \12995 );
nor \U$15527 ( \15780 , \15777 , \15779 );
not \U$15528 ( \15781 , \15780 );
not \U$15529 ( \15782 , RIbe287c8_28);
not \U$15530 ( \15783 , \12811 );
or \U$15531 ( \15784 , \15782 , \15783 );
nand \U$15532 ( \15785 , RIbe28480_21, RIbe2ae38_110);
nand \U$15533 ( \15786 , \15784 , \15785 );
xnor \U$15534 ( \15787 , \15786 , RIbe2aeb0_111);
and \U$15535 ( \15788 , \15781 , \15787 );
not \U$15536 ( \15789 , \15781 );
not \U$15537 ( \15790 , \15787 );
and \U$15538 ( \15791 , \15789 , \15790 );
nor \U$15539 ( \15792 , \15788 , \15791 );
not \U$15540 ( \15793 , RIbe27f58_10);
not \U$15541 ( \15794 , \13590 );
or \U$15542 ( \15795 , \15793 , \15794 );
nand \U$15543 ( \15796 , \13012 , RIbe27e68_8);
nand \U$15544 ( \15797 , \15795 , \15796 );
and \U$15545 ( \15798 , \15797 , \12866 );
not \U$15546 ( \15799 , \15797 );
and \U$15547 ( \15800 , \15799 , \12863 );
nor \U$15548 ( \15801 , \15798 , \15800 );
not \U$15549 ( \15802 , \15801 );
and \U$15550 ( \15803 , \15792 , \15802 );
not \U$15551 ( \15804 , \15792 );
and \U$15552 ( \15805 , \15804 , \15801 );
nor \U$15553 ( \15806 , \15803 , \15805 );
not \U$15554 ( \15807 , \15806 );
nand \U$15555 ( \15808 , \15582 , \15601 );
nand \U$15556 ( \15809 , \15807 , \15808 );
not \U$15557 ( \15810 , \15809 );
not \U$15558 ( \15811 , \15694 );
not \U$15559 ( \15812 , \15735 );
or \U$15560 ( \15813 , \15811 , \15812 );
nand \U$15561 ( \15814 , \15813 , \15656 );
not \U$15562 ( \15815 , \15694 );
nand \U$15563 ( \15816 , \15815 , \15736 );
nand \U$15564 ( \15817 , \15814 , \15816 );
not \U$15565 ( \15818 , \15817 );
or \U$15566 ( \15819 , \15810 , \15818 );
not \U$15567 ( \15820 , \15808 );
nand \U$15568 ( \15821 , \15820 , \15806 );
nand \U$15569 ( \15822 , \15819 , \15821 );
not \U$15570 ( \15823 , \15822 );
nand \U$15571 ( \15824 , \15427 , \15417 );
not \U$15572 ( \15825 , \15824 );
not \U$15573 ( \15826 , \15473 );
or \U$15574 ( \15827 , \15825 , \15826 );
not \U$15575 ( \15828 , \15417 );
nand \U$15576 ( \15829 , \15828 , \15428 );
nand \U$15577 ( \15830 , \15827 , \15829 );
not \U$15578 ( \15831 , \15830 );
not \U$15579 ( \15832 , \15831 );
not \U$15580 ( \15833 , \15522 );
not \U$15581 ( \15834 , \15512 );
or \U$15582 ( \15835 , \15833 , \15834 );
nand \U$15583 ( \15836 , \15835 , \15503 );
not \U$15584 ( \15837 , \15522 );
nand \U$15585 ( \15838 , \15837 , \15511 );
nand \U$15586 ( \15839 , \15836 , \15838 );
not \U$15587 ( \15840 , \15839 );
not \U$15588 ( \15841 , \15840 );
or \U$15589 ( \15842 , \15832 , \15841 );
xor \U$15590 ( \15843 , \15482 , \15486 );
and \U$15591 ( \15844 , \15843 , \15492 );
and \U$15592 ( \15845 , \15482 , \15486 );
or \U$15593 ( \15846 , \15844 , \15845 );
nand \U$15594 ( \15847 , \15842 , \15846 );
nand \U$15595 ( \15848 , \15830 , \15839 );
nand \U$15596 ( \15849 , \15847 , \15848 );
not \U$15597 ( \15850 , \15849 );
not \U$15598 ( \15851 , \15850 );
or \U$15599 ( \15852 , \15823 , \15851 );
not \U$15600 ( \15853 , \15822 );
nand \U$15601 ( \15854 , \15853 , \15849 );
nand \U$15602 ( \15855 , \15852 , \15854 );
not \U$15603 ( \15856 , \15454 );
or \U$15604 ( \15857 , \15856 , \15443 );
nand \U$15605 ( \15858 , \15857 , \15465 );
nand \U$15606 ( \15859 , \15856 , \15443 );
nand \U$15607 ( \15860 , \15858 , \15859 );
not \U$15608 ( \15861 , \15709 );
not \U$15609 ( \15862 , \15719 );
or \U$15610 ( \15863 , \15861 , \15862 );
or \U$15611 ( \15864 , \15719 , \15709 );
nand \U$15612 ( \15865 , \15864 , \15734 );
nand \U$15613 ( \15866 , \15863 , \15865 );
xor \U$15614 ( \15867 , \15860 , \15866 );
or \U$15615 ( \15868 , \15676 , \15664 );
nand \U$15616 ( \15869 , \15868 , \15689 );
nand \U$15617 ( \15870 , \15676 , \15664 );
nand \U$15618 ( \15871 , \15869 , \15870 );
xor \U$15619 ( \15872 , \15867 , \15871 );
not \U$15620 ( \15873 , RIbe2ab68_104);
nor \U$15621 ( \15874 , \3703 , \15873 );
not \U$15622 ( \15875 , \4027 );
nor \U$15623 ( \15876 , \15875 , \13192 );
nor \U$15624 ( \15877 , \15874 , \15876 );
and \U$15625 ( \15878 , \15877 , \3448 );
not \U$15626 ( \15879 , \15877 );
and \U$15627 ( \15880 , \15879 , \3471 );
nor \U$15628 ( \15881 , \15878 , \15880 );
not \U$15629 ( \15882 , RIbe2b1f8_118);
not \U$15630 ( \15883 , \6630 );
or \U$15631 ( \15884 , \15882 , \15883 );
not \U$15632 ( \15885 , \7098 );
nand \U$15633 ( \15886 , \15885 , RIbe2b180_117);
nand \U$15634 ( \15887 , \15884 , \15886 );
and \U$15635 ( \15888 , \15887 , \6118 );
not \U$15636 ( \15889 , \15887 );
and \U$15637 ( \15890 , \15889 , \10272 );
nor \U$15638 ( \15891 , \15888 , \15890 );
not \U$15639 ( \15892 , \15891 );
not \U$15640 ( \15893 , RIbe2afa0_113);
not \U$15641 ( \15894 , \4828 );
not \U$15642 ( \15895 , \15894 );
or \U$15643 ( \15896 , \15893 , \15895 );
nand \U$15644 ( \15897 , \5052 , RIbe2af28_112);
nand \U$15645 ( \15898 , \15896 , \15897 );
and \U$15646 ( \15899 , \15898 , \4586 );
not \U$15647 ( \15900 , \15898 );
and \U$15648 ( \15901 , \15900 , \4592 );
nor \U$15649 ( \15902 , \15899 , \15901 );
not \U$15650 ( \15903 , \15902 );
or \U$15651 ( \15904 , \15892 , \15903 );
or \U$15652 ( \15905 , \15891 , \15902 );
nand \U$15653 ( \15906 , \15904 , \15905 );
not \U$15654 ( \15907 , RIbe2b630_127);
not \U$15655 ( \15908 , \6413 );
or \U$15656 ( \15909 , \15907 , \15908 );
nand \U$15657 ( \15910 , \4808 , RIbe2b018_114);
nand \U$15658 ( \15911 , \15909 , \15910 );
not \U$15659 ( \15912 , \15911 );
not \U$15660 ( \15913 , \4323 );
and \U$15661 ( \15914 , \15912 , \15913 );
and \U$15662 ( \15915 , \15911 , \4323 );
nor \U$15663 ( \15916 , \15914 , \15915 );
xnor \U$15664 ( \15917 , \15906 , \15916 );
xor \U$15665 ( \15918 , \15881 , \15917 );
not \U$15666 ( \15919 , RIbe2b270_119);
not \U$15667 ( \15920 , \8231 );
or \U$15668 ( \15921 , \15919 , \15920 );
nand \U$15669 ( \15922 , \9939 , RIbe2b108_116);
nand \U$15670 ( \15923 , \15921 , \15922 );
and \U$15671 ( \15924 , \15923 , \10972 );
not \U$15672 ( \15925 , \15923 );
and \U$15673 ( \15926 , \15925 , \10969 );
nor \U$15674 ( \15927 , \15924 , \15926 );
not \U$15675 ( \15928 , \15927 );
not \U$15676 ( \15929 , RIbe2b090_115);
not \U$15677 ( \15930 , \6536 );
or \U$15678 ( \15931 , \15929 , \15930 );
nand \U$15679 ( \15932 , \6540 , RIbe2a280_85);
nand \U$15680 ( \15933 , \15931 , \15932 );
not \U$15681 ( \15934 , \15933 );
not \U$15682 ( \15935 , \6891 );
and \U$15683 ( \15936 , \15934 , \15935 );
and \U$15684 ( \15937 , \15933 , \6548 );
nor \U$15685 ( \15938 , \15936 , \15937 );
not \U$15686 ( \15939 , \15938 );
not \U$15687 ( \15940 , \15939 );
not \U$15688 ( \15941 , RIbe2a208_84);
not \U$15689 ( \15942 , \13238 );
or \U$15690 ( \15943 , \15941 , \15942 );
nand \U$15691 ( \15944 , \6596 , RIbe2a190_83);
nand \U$15692 ( \15945 , \15943 , \15944 );
and \U$15693 ( \15946 , \15945 , \6601 );
not \U$15694 ( \15947 , \15945 );
and \U$15695 ( \15948 , \15947 , \10888 );
nor \U$15696 ( \15949 , \15946 , \15948 );
not \U$15697 ( \15950 , \15949 );
not \U$15698 ( \15951 , \15950 );
or \U$15699 ( \15952 , \15940 , \15951 );
nand \U$15700 ( \15953 , \15949 , \15938 );
nand \U$15701 ( \15954 , \15952 , \15953 );
not \U$15702 ( \15955 , \15954 );
or \U$15703 ( \15956 , \15928 , \15955 );
or \U$15704 ( \15957 , \15954 , \15927 );
nand \U$15705 ( \15958 , \15956 , \15957 );
xor \U$15706 ( \15959 , \15918 , \15958 );
xor \U$15707 ( \15960 , \15872 , \15959 );
not \U$15708 ( \15961 , RIbe29bf0_71);
not \U$15709 ( \15962 , \12871 );
or \U$15710 ( \15963 , \15961 , \15962 );
nand \U$15711 ( \15964 , \13728 , RIbe28f48_44);
nand \U$15712 ( \15965 , \15963 , \15964 );
and \U$15713 ( \15966 , \15965 , \12716 );
not \U$15714 ( \15967 , \15965 );
and \U$15715 ( \15968 , \15967 , \12723 );
nor \U$15716 ( \15969 , \15966 , \15968 );
not \U$15717 ( \15970 , RIbe28ed0_43);
not \U$15718 ( \15971 , \14071 );
or \U$15719 ( \15972 , \15970 , \15971 );
nand \U$15720 ( \15973 , \14074 , RIbe27fd0_11);
nand \U$15721 ( \15974 , \15972 , \15973 );
and \U$15722 ( \15975 , \15974 , \12742 );
not \U$15723 ( \15976 , \15974 );
and \U$15724 ( \15977 , \15976 , \14358 );
nor \U$15725 ( \15978 , \15975 , \15977 );
and \U$15726 ( \15979 , \15969 , \15978 );
not \U$15727 ( \15980 , \15969 );
not \U$15728 ( \15981 , \15978 );
and \U$15729 ( \15982 , \15980 , \15981 );
or \U$15730 ( \15983 , \15979 , \15982 );
not \U$15731 ( \15984 , \12751 );
not \U$15732 ( \15985 , \9801 );
and \U$15733 ( \15986 , \15984 , \15985 );
and \U$15734 ( \15987 , \14726 , RIbe29dd0_75);
nor \U$15735 ( \15988 , \15986 , \15987 );
and \U$15736 ( \15989 , \15988 , \12924 );
not \U$15737 ( \15990 , \15988 );
and \U$15738 ( \15991 , \15990 , \12927 );
nor \U$15739 ( \15992 , \15989 , \15991 );
xor \U$15740 ( \15993 , \15983 , \15992 );
not \U$15741 ( \15994 , RIbe2a988_100);
not \U$15742 ( \15995 , \7299 );
or \U$15743 ( \15996 , \15994 , \15995 );
nand \U$15744 ( \15997 , \8287 , RIbe2a910_99);
nand \U$15745 ( \15998 , \15996 , \15997 );
and \U$15746 ( \15999 , \15998 , \13227 );
not \U$15747 ( \16000 , \15998 );
and \U$15748 ( \16001 , \16000 , \6992 );
nor \U$15749 ( \16002 , \15999 , \16001 );
not \U$15750 ( \16003 , RIbe2b5b8_126);
not \U$15751 ( \16004 , \10949 );
or \U$15752 ( \16005 , \16003 , \16004 );
nand \U$15753 ( \16006 , \10952 , RIbe2a3e8_88);
nand \U$15754 ( \16007 , \16005 , \16006 );
and \U$15755 ( \16008 , \16007 , \6949 );
not \U$15756 ( \16009 , \16007 );
not \U$15757 ( \16010 , \7984 );
and \U$15758 ( \16011 , \16009 , \16010 );
nor \U$15759 ( \16012 , \16008 , \16011 );
and \U$15760 ( \16013 , \16002 , \16012 );
not \U$15761 ( \16014 , \16002 );
not \U$15762 ( \16015 , \16012 );
and \U$15763 ( \16016 , \16014 , \16015 );
or \U$15764 ( \16017 , \16013 , \16016 );
not \U$15765 ( \16018 , RIbe2a5c8_92);
not \U$15766 ( \16019 , \6560 );
or \U$15767 ( \16020 , \16018 , \16019 );
nand \U$15768 ( \16021 , \6963 , RIbe2a550_91);
nand \U$15769 ( \16022 , \16020 , \16021 );
and \U$15770 ( \16023 , \16022 , \6569 );
not \U$15771 ( \16024 , \16022 );
and \U$15772 ( \16025 , \16024 , \7293 );
nor \U$15773 ( \16026 , \16023 , \16025 );
not \U$15774 ( \16027 , \16026 );
and \U$15775 ( \16028 , \16017 , \16027 );
not \U$15776 ( \16029 , \16017 );
and \U$15777 ( \16030 , \16029 , \16026 );
nor \U$15778 ( \16031 , \16028 , \16030 );
xor \U$15779 ( \16032 , \15993 , \16031 );
not \U$15780 ( \16033 , \13669 );
not \U$15781 ( \16034 , \16033 );
not \U$15782 ( \16035 , \12380 );
and \U$15783 ( \16036 , \16034 , \16035 );
and \U$15784 ( \16037 , \15205 , RIbe29fb0_79);
nor \U$15785 ( \16038 , \16036 , \16037 );
and \U$15786 ( \16039 , \16038 , \12956 );
not \U$15787 ( \16040 , \16038 );
and \U$15788 ( \16041 , \16040 , \12195 );
nor \U$15789 ( \16042 , \16039 , \16041 );
not \U$15790 ( \16043 , RIbe2acd0_107);
not \U$15791 ( \16044 , \13024 );
or \U$15792 ( \16045 , \16043 , \16044 );
nand \U$15793 ( \16046 , \12212 , RIbe2a028_80);
nand \U$15794 ( \16047 , \16045 , \16046 );
not \U$15795 ( \16048 , \16047 );
not \U$15796 ( \16049 , \10943 );
and \U$15797 ( \16050 , \16048 , \16049 );
and \U$15798 ( \16051 , \16047 , \13033 );
nor \U$15799 ( \16052 , \16050 , \16051 );
xor \U$15800 ( \16053 , \16042 , \16052 );
and \U$15801 ( \16054 , \10916 , RIbe2a370_87);
and \U$15802 ( \16055 , \9914 , RIbe2a2f8_86);
nor \U$15803 ( \16056 , \16054 , \16055 );
and \U$15804 ( \16057 , \16056 , \7970 );
not \U$15805 ( \16058 , \16056 );
buf \U$15806 ( \16059 , \15233 );
and \U$15807 ( \16060 , \16058 , \16059 );
nor \U$15808 ( \16061 , \16057 , \16060 );
xor \U$15809 ( \16062 , \16053 , \16061 );
xor \U$15810 ( \16063 , \16032 , \16062 );
and \U$15811 ( \16064 , \15960 , \16063 );
and \U$15812 ( \16065 , \15872 , \15959 );
or \U$15813 ( \16066 , \16064 , \16065 );
xnor \U$15814 ( \16067 , \15855 , \16066 );
not \U$15815 ( \16068 , \16067 );
not \U$15816 ( \16069 , \15533 );
and \U$15817 ( \16070 , \16069 , \15541 );
nor \U$15818 ( \16071 , \16070 , \15546 );
nor \U$15819 ( \16072 , \15541 , \16069 );
nor \U$15820 ( \16073 , \16071 , \16072 );
nand \U$15821 ( \16074 , \15609 , \15605 );
and \U$15822 ( \16075 , \15740 , \16074 );
nor \U$15823 ( \16076 , \15609 , \15605 );
nor \U$15824 ( \16077 , \16075 , \16076 );
xor \U$15825 ( \16078 , \16073 , \16077 );
and \U$15826 ( \16079 , \15477 , \15526 );
not \U$15827 ( \16080 , \15493 );
nor \U$15828 ( \16081 , \16079 , \16080 );
nor \U$15829 ( \16082 , \15526 , \15477 );
nor \U$15830 ( \16083 , \16081 , \16082 );
xor \U$15831 ( \16084 , \16078 , \16083 );
not \U$15832 ( \16085 , \16084 );
xor \U$15833 ( \16086 , \15872 , \15959 );
xor \U$15834 ( \16087 , \16086 , \16063 );
not \U$15835 ( \16088 , \16087 );
not \U$15836 ( \16089 , \15817 );
xor \U$15837 ( \16090 , \15808 , \15806 );
not \U$15838 ( \16091 , \16090 );
or \U$15839 ( \16092 , \16089 , \16091 );
or \U$15840 ( \16093 , \15817 , \16090 );
nand \U$15841 ( \16094 , \16092 , \16093 );
not \U$15842 ( \16095 , \16094 );
not \U$15843 ( \16096 , \15653 );
not \U$15844 ( \16097 , \15621 );
or \U$15845 ( \16098 , \16096 , \16097 );
not \U$15846 ( \16099 , \15622 );
not \U$15847 ( \16100 , \15650 );
or \U$15848 ( \16101 , \16099 , \16100 );
nand \U$15849 ( \16102 , \16101 , \15636 );
nand \U$15850 ( \16103 , \16098 , \16102 );
nand \U$15851 ( \16104 , \15570 , \15581 );
and \U$15852 ( \16105 , \16104 , \15561 );
nor \U$15853 ( \16106 , \15570 , \15581 );
nor \U$15854 ( \16107 , \16105 , \16106 );
not \U$15855 ( \16108 , \16107 );
and \U$15856 ( \16109 , \16103 , \16108 );
not \U$15857 ( \16110 , \16103 );
and \U$15858 ( \16111 , \16110 , \16107 );
nor \U$15859 ( \16112 , \16109 , \16111 );
not \U$15860 ( \16113 , \15590 );
nand \U$15861 ( \16114 , \16113 , \4821 );
and \U$15862 ( \16115 , \16114 , \15600 );
and \U$15863 ( \16116 , \3471 , \15590 );
nor \U$15864 ( \16117 , \16115 , \16116 );
not \U$15865 ( \16118 , \16117 );
and \U$15866 ( \16119 , \16112 , \16118 );
not \U$15867 ( \16120 , \16112 );
and \U$15868 ( \16121 , \16120 , \16117 );
or \U$15869 ( \16122 , \16119 , \16121 );
not \U$15870 ( \16123 , \16122 );
and \U$15871 ( \16124 , \16095 , \16123 );
and \U$15872 ( \16125 , \16094 , \16122 );
nor \U$15873 ( \16126 , \16124 , \16125 );
not \U$15874 ( \16127 , \16126 );
or \U$15875 ( \16128 , \16088 , \16127 );
or \U$15876 ( \16129 , \16126 , \16087 );
nand \U$15877 ( \16130 , \16128 , \16129 );
nand \U$15878 ( \16131 , \16085 , \16130 );
not \U$15879 ( \16132 , \16131 );
or \U$15880 ( \16133 , \16068 , \16132 );
not \U$15881 ( \16134 , \15846 );
not \U$15882 ( \16135 , \15840 );
or \U$15883 ( \16136 , \16134 , \16135 );
or \U$15884 ( \16137 , \15840 , \15846 );
nand \U$15885 ( \16138 , \16136 , \16137 );
and \U$15886 ( \16139 , \16138 , \15830 );
not \U$15887 ( \16140 , \16138 );
and \U$15888 ( \16141 , \16140 , \15831 );
nor \U$15889 ( \16142 , \16139 , \16141 );
not \U$15890 ( \16143 , \15396 );
not \U$15891 ( \16144 , \15393 );
or \U$15892 ( \16145 , \16143 , \16144 );
nand \U$15893 ( \16146 , \15392 , \15395 );
nand \U$15894 ( \16147 , \15388 , \16146 );
nand \U$15895 ( \16148 , \16145 , \16147 );
xor \U$15896 ( \16149 , \16142 , \16148 );
not \U$15897 ( \16150 , \15547 );
not \U$15898 ( \16151 , \15527 );
or \U$15899 ( \16152 , \16150 , \16151 );
or \U$15900 ( \16153 , \15527 , \15547 );
nand \U$15901 ( \16154 , \16153 , \15741 );
nand \U$15902 ( \16155 , \16152 , \16154 );
and \U$15903 ( \16156 , \16149 , \16155 );
and \U$15904 ( \16157 , \16142 , \16148 );
or \U$15905 ( \16158 , \16156 , \16157 );
nand \U$15906 ( \16159 , \16133 , \16158 );
or \U$15907 ( \16160 , \16131 , \16067 );
nand \U$15908 ( \16161 , \16159 , \16160 );
not \U$15909 ( \16162 , \16161 );
not \U$15910 ( \16163 , \16108 );
not \U$15911 ( \16164 , \16118 );
or \U$15912 ( \16165 , \16163 , \16164 );
not \U$15913 ( \16166 , \16117 );
not \U$15914 ( \16167 , \16107 );
or \U$15915 ( \16168 , \16166 , \16167 );
nand \U$15916 ( \16169 , \16168 , \16103 );
nand \U$15917 ( \16170 , \16165 , \16169 );
xor \U$15918 ( \16171 , \15860 , \15866 );
and \U$15919 ( \16172 , \16171 , \15871 );
and \U$15920 ( \16173 , \15860 , \15866 );
or \U$15921 ( \16174 , \16172 , \16173 );
xor \U$15922 ( \16175 , \16170 , \16174 );
xor \U$15923 ( \16176 , \15881 , \15917 );
and \U$15924 ( \16177 , \16176 , \15958 );
and \U$15925 ( \16178 , \15881 , \15917 );
or \U$15926 ( \16179 , \16177 , \16178 );
xor \U$15927 ( \16180 , \16175 , \16179 );
nand \U$15928 ( \16181 , \15891 , \15916 );
and \U$15929 ( \16182 , \16181 , \15902 );
nor \U$15930 ( \16183 , \15916 , \15891 );
nor \U$15931 ( \16184 , \16182 , \16183 );
not \U$15932 ( \16185 , \16184 );
not \U$15933 ( \16186 , \16185 );
not \U$15934 ( \16187 , \16015 );
not \U$15935 ( \16188 , \16027 );
or \U$15936 ( \16189 , \16187 , \16188 );
not \U$15937 ( \16190 , \16026 );
not \U$15938 ( \16191 , \16012 );
or \U$15939 ( \16192 , \16190 , \16191 );
nand \U$15940 ( \16193 , \16192 , \16002 );
nand \U$15941 ( \16194 , \16189 , \16193 );
not \U$15942 ( \16195 , \16194 );
not \U$15943 ( \16196 , \16195 );
or \U$15944 ( \16197 , \16186 , \16196 );
nand \U$15945 ( \16198 , \16194 , \16184 );
nand \U$15946 ( \16199 , \16197 , \16198 );
not \U$15947 ( \16200 , \16199 );
not \U$15948 ( \16201 , \15927 );
not \U$15949 ( \16202 , \15950 );
or \U$15950 ( \16203 , \16201 , \16202 );
nand \U$15951 ( \16204 , \16203 , \15939 );
not \U$15952 ( \16205 , \15927 );
nand \U$15953 ( \16206 , \16205 , \15949 );
nand \U$15954 ( \16207 , \16204 , \16206 );
not \U$15955 ( \16208 , \16207 );
not \U$15956 ( \16209 , \16208 );
and \U$15957 ( \16210 , \16200 , \16209 );
and \U$15958 ( \16211 , \16199 , \16208 );
nor \U$15959 ( \16212 , \16210 , \16211 );
nand \U$15960 ( \16213 , \15780 , \15787 );
not \U$15961 ( \16214 , \16213 );
not \U$15962 ( \16215 , \15801 );
or \U$15963 ( \16216 , \16214 , \16215 );
nand \U$15964 ( \16217 , \15781 , \15790 );
nand \U$15965 ( \16218 , \16216 , \16217 );
not \U$15966 ( \16219 , \15981 );
not \U$15967 ( \16220 , \15969 );
or \U$15968 ( \16221 , \16219 , \16220 );
or \U$15969 ( \16222 , \15969 , \15981 );
nand \U$15970 ( \16223 , \16222 , \15992 );
nand \U$15971 ( \16224 , \16221 , \16223 );
xor \U$15972 ( \16225 , \16218 , \16224 );
nand \U$15973 ( \16226 , \16061 , \16052 );
and \U$15974 ( \16227 , \16226 , \16042 );
nor \U$15975 ( \16228 , \16061 , \16052 );
nor \U$15976 ( \16229 , \16227 , \16228 );
xnor \U$15977 ( \16230 , \16225 , \16229 );
xor \U$15978 ( \16231 , \16212 , \16230 );
not \U$15979 ( \16232 , RIbe2b180_117);
not \U$15980 ( \16233 , \5455 );
or \U$15981 ( \16234 , \16232 , \16233 );
nand \U$15982 ( \16235 , \15885 , RIbe2b270_119);
nand \U$15983 ( \16236 , \16234 , \16235 );
and \U$15984 ( \16237 , \16236 , \6117 );
not \U$15985 ( \16238 , \16236 );
and \U$15986 ( \16239 , \16238 , \6637 );
nor \U$15987 ( \16240 , \16237 , \16239 );
not \U$15988 ( \16241 , RIbe2b108_116);
not \U$15989 ( \16242 , \8231 );
or \U$15990 ( \16243 , \16241 , \16242 );
nand \U$15991 ( \16244 , \6859 , RIbe2b090_115);
nand \U$15992 ( \16245 , \16243 , \16244 );
and \U$15993 ( \16246 , \16245 , \6623 );
not \U$15994 ( \16247 , \16245 );
and \U$15995 ( \16248 , \16247 , \6624 );
nor \U$15996 ( \16249 , \16246 , \16248 );
xor \U$15997 ( \16250 , \16240 , \16249 );
not \U$15998 ( \16251 , RIbe2af28_112);
not \U$15999 ( \16252 , \6427 );
or \U$16000 ( \16253 , \16251 , \16252 );
nand \U$16001 ( \16254 , \7056 , RIbe2b1f8_118);
nand \U$16002 ( \16255 , \16253 , \16254 );
and \U$16003 ( \16256 , \16255 , \4586 );
not \U$16004 ( \16257 , \16255 );
and \U$16005 ( \16258 , \16257 , \4592 );
nor \U$16006 ( \16259 , \16256 , \16258 );
xor \U$16007 ( \16260 , \16250 , \16259 );
not \U$16008 ( \16261 , \3290 );
nand \U$16009 ( \16262 , \3457 , RIbe2ab68_104);
not \U$16010 ( \16263 , \16262 );
or \U$16011 ( \16264 , \16261 , \16263 );
or \U$16012 ( \16265 , \4346 , \16262 );
nand \U$16013 ( \16266 , \16264 , \16265 );
not \U$16014 ( \16267 , RIbe2b018_114);
not \U$16015 ( \16268 , \4317 );
or \U$16016 ( \16269 , \16267 , \16268 );
nand \U$16017 ( \16270 , \6418 , RIbe2afa0_113);
nand \U$16018 ( \16271 , \16269 , \16270 );
not \U$16019 ( \16272 , \16271 );
not \U$16020 ( \16273 , \4323 );
and \U$16021 ( \16274 , \16272 , \16273 );
and \U$16022 ( \16275 , \16271 , \4323 );
nor \U$16023 ( \16276 , \16274 , \16275 );
xor \U$16024 ( \16277 , \16266 , \16276 );
not \U$16025 ( \16278 , RIbe2aaf0_103);
not \U$16026 ( \16279 , \6783 );
or \U$16027 ( \16280 , \16278 , \16279 );
nand \U$16028 ( \16281 , \4027 , RIbe2b630_127);
nand \U$16029 ( \16282 , \16280 , \16281 );
not \U$16030 ( \16283 , \16282 );
not \U$16031 ( \16284 , \3448 );
and \U$16032 ( \16285 , \16283 , \16284 );
and \U$16033 ( \16286 , \16282 , \3448 );
nor \U$16034 ( \16287 , \16285 , \16286 );
xnor \U$16035 ( \16288 , \16277 , \16287 );
xor \U$16036 ( \16289 , \16260 , \16288 );
not \U$16037 ( \16290 , RIbe2a550_91);
not \U$16038 ( \16291 , \7954 );
or \U$16039 ( \16292 , \16290 , \16291 );
nand \U$16040 ( \16293 , \7958 , RIbe2a988_100);
nand \U$16041 ( \16294 , \16292 , \16293 );
and \U$16042 ( \16295 , \16294 , \7293 );
not \U$16043 ( \16296 , \16294 );
and \U$16044 ( \16297 , \16296 , \6572 );
nor \U$16045 ( \16298 , \16295 , \16297 );
not \U$16046 ( \16299 , RIbe2a190_83);
not \U$16047 ( \16300 , \6592 );
or \U$16048 ( \16301 , \16299 , \16300 );
nand \U$16049 ( \16302 , \7278 , RIbe2a5c8_92);
nand \U$16050 ( \16303 , \16301 , \16302 );
and \U$16051 ( \16304 , \16303 , \6601 );
not \U$16052 ( \16305 , \16303 );
and \U$16053 ( \16306 , \16305 , \7949 );
nor \U$16054 ( \16307 , \16304 , \16306 );
xor \U$16055 ( \16308 , \16298 , \16307 );
not \U$16056 ( \16309 , RIbe2a280_85);
not \U$16057 ( \16310 , \6537 );
or \U$16058 ( \16311 , \16309 , \16310 );
nand \U$16059 ( \16312 , \6540 , RIbe2a208_84);
nand \U$16060 ( \16313 , \16311 , \16312 );
and \U$16061 ( \16314 , \16313 , \6546 );
not \U$16062 ( \16315 , \16313 );
and \U$16063 ( \16316 , \16315 , \6891 );
nor \U$16064 ( \16317 , \16314 , \16316 );
xor \U$16065 ( \16318 , \16308 , \16317 );
and \U$16066 ( \16319 , \16289 , \16318 );
not \U$16067 ( \16320 , \16289 );
not \U$16068 ( \16321 , \16318 );
and \U$16069 ( \16322 , \16320 , \16321 );
nor \U$16070 ( \16323 , \16319 , \16322 );
not \U$16071 ( \16324 , \16323 );
xnor \U$16072 ( \16325 , \16231 , \16324 );
xor \U$16073 ( \16326 , \16180 , \16325 );
not \U$16074 ( \16327 , RIbe285e8_24);
not \U$16075 ( \16328 , \13518 );
or \U$16076 ( \16329 , \16327 , \16328 );
nand \U$16077 ( \16330 , \12794 , RIbe287c8_28);
nand \U$16078 ( \16331 , \16329 , \16330 );
and \U$16079 ( \16332 , \16331 , \12801 );
not \U$16080 ( \16333 , \16331 );
not \U$16081 ( \16334 , \12893 );
and \U$16082 ( \16335 , \16333 , \16334 );
nor \U$16083 ( \16336 , \16332 , \16335 );
not \U$16084 ( \16337 , \16336 );
not \U$16085 ( \16338 , RIbe28480_21);
not \U$16086 ( \16339 , \13003 );
or \U$16087 ( \16340 , \16338 , \16339 );
nand \U$16088 ( \16341 , RIbe28408_20, RIbe2ae38_110);
nand \U$16089 ( \16342 , \16340 , \16341 );
xor \U$16090 ( \16343 , RIbe2aeb0_111, \16342 );
and \U$16091 ( \16344 , \16343 , \4346 );
not \U$16092 ( \16345 , \16343 );
and \U$16093 ( \16346 , \16345 , \2887 );
nor \U$16094 ( \16347 , \16344 , \16346 );
not \U$16095 ( \16348 , \16347 );
or \U$16096 ( \16349 , \16337 , \16348 );
or \U$16097 ( \16350 , \16347 , \16336 );
nand \U$16098 ( \16351 , \16349 , \16350 );
xor \U$16099 ( \16352 , \15993 , \16031 );
and \U$16100 ( \16353 , \16352 , \16062 );
and \U$16101 ( \16354 , \15993 , \16031 );
or \U$16102 ( \16355 , \16353 , \16354 );
xor \U$16103 ( \16356 , \16351 , \16355 );
not \U$16104 ( \16357 , RIbe27e68_8);
not \U$16105 ( \16358 , \12831 );
or \U$16106 ( \16359 , \16357 , \16358 );
nand \U$16107 ( \16360 , \12834 , RIbe28660_25);
nand \U$16108 ( \16361 , \16359 , \16360 );
not \U$16109 ( \16362 , \16361 );
not \U$16110 ( \16363 , RIbe2a730_95);
not \U$16111 ( \16364 , RIbe2b450_123);
or \U$16112 ( \16365 , \16363 , \16364 );
nand \U$16113 ( \16366 , \16365 , RIbe2a7a8_96);
not \U$16114 ( \16367 , \16366 );
and \U$16115 ( \16368 , \16362 , \16367 );
and \U$16116 ( \16369 , \16361 , \15263 );
nor \U$16117 ( \16370 , \16368 , \16369 );
not \U$16118 ( \16371 , RIbe27fd0_11);
not \U$16119 ( \16372 , \12732 );
or \U$16120 ( \16373 , \16371 , \16372 );
nand \U$16121 ( \16374 , \13077 , RIbe27f58_10);
nand \U$16122 ( \16375 , \16373 , \16374 );
and \U$16123 ( \16376 , \16375 , \13570 );
not \U$16124 ( \16377 , \16375 );
and \U$16125 ( \16378 , \16377 , \12746 );
nor \U$16126 ( \16379 , \16376 , \16378 );
xnor \U$16127 ( \16380 , \16370 , \16379 );
not \U$16128 ( \16381 , RIbe28f48_44);
not \U$16129 ( \16382 , \15573 );
not \U$16130 ( \16383 , \16382 );
not \U$16131 ( \16384 , \16383 );
or \U$16132 ( \16385 , \16381 , \16384 );
nand \U$16133 ( \16386 , \12711 , RIbe28ed0_43);
nand \U$16134 ( \16387 , \16385 , \16386 );
and \U$16135 ( \16388 , \16387 , \12723 );
not \U$16136 ( \16389 , \16387 );
and \U$16137 ( \16390 , \16389 , \13068 );
nor \U$16138 ( \16391 , \16388 , \16390 );
xnor \U$16139 ( \16392 , \16380 , \16391 );
and \U$16140 ( \16393 , \12942 , RIbe29e48_76);
not \U$16141 ( \16394 , RIbe29dd0_75);
nor \U$16142 ( \16395 , \16394 , \14397 );
nor \U$16143 ( \16396 , \16393 , \16395 );
and \U$16144 ( \16397 , \16396 , \12960 );
not \U$16145 ( \16398 , \16396 );
and \U$16146 ( \16399 , \16398 , \12195 );
nor \U$16147 ( \16400 , \16397 , \16399 );
not \U$16148 ( \16401 , RIbe29c68_72);
not \U$16149 ( \16402 , \12920 );
or \U$16150 ( \16403 , \16401 , \16402 );
nand \U$16151 ( \16404 , \14491 , RIbe29bf0_71);
nand \U$16152 ( \16405 , \16403 , \16404 );
not \U$16153 ( \16406 , \16405 );
not \U$16154 ( \16407 , \12924 );
and \U$16155 ( \16408 , \16406 , \16407 );
and \U$16156 ( \16409 , \16405 , \12769 );
nor \U$16157 ( \16410 , \16408 , \16409 );
and \U$16158 ( \16411 , \16400 , \16410 );
not \U$16159 ( \16412 , \16400 );
not \U$16160 ( \16413 , \16410 );
and \U$16161 ( \16414 , \16412 , \16413 );
nor \U$16162 ( \16415 , \16411 , \16414 );
not \U$16163 ( \16416 , RIbe2a028_80);
not \U$16164 ( \16417 , \10936 );
or \U$16165 ( \16418 , \16416 , \16417 );
nand \U$16166 ( \16419 , \12971 , RIbe29fb0_79);
nand \U$16167 ( \16420 , \16418 , \16419 );
not \U$16168 ( \16421 , \16420 );
not \U$16169 ( \16422 , \10943 );
and \U$16170 ( \16423 , \16421 , \16422 );
and \U$16171 ( \16424 , \16420 , \10940 );
nor \U$16172 ( \16425 , \16423 , \16424 );
and \U$16173 ( \16426 , \16415 , \16425 );
not \U$16174 ( \16427 , \16415 );
not \U$16175 ( \16428 , \16425 );
and \U$16176 ( \16429 , \16427 , \16428 );
nor \U$16177 ( \16430 , \16426 , \16429 );
not \U$16178 ( \16431 , \13477 );
and \U$16179 ( \16432 , \16431 , RIbe2a2f8_86);
and \U$16180 ( \16433 , \13038 , RIbe2acd0_107);
nor \U$16181 ( \16434 , \16432 , \16433 );
and \U$16182 ( \16435 , \16434 , \8077 );
not \U$16183 ( \16436 , \16434 );
not \U$16184 ( \16437 , \8077 );
and \U$16185 ( \16438 , \16436 , \16437 );
nor \U$16186 ( \16439 , \16435 , \16438 );
not \U$16187 ( \16440 , RIbe2a3e8_88);
not \U$16188 ( \16441 , \10949 );
or \U$16189 ( \16442 , \16440 , \16441 );
nand \U$16190 ( \16443 , \9891 , RIbe2a370_87);
nand \U$16191 ( \16444 , \16442 , \16443 );
and \U$16192 ( \16445 , \16444 , \7984 );
not \U$16193 ( \16446 , \16444 );
and \U$16194 ( \16447 , \16446 , \16010 );
nor \U$16195 ( \16448 , \16445 , \16447 );
xnor \U$16196 ( \16449 , \16439 , \16448 );
not \U$16197 ( \16450 , RIbe2a910_99);
not \U$16198 ( \16451 , \6980 );
or \U$16199 ( \16452 , \16450 , \16451 );
nand \U$16200 ( \16453 , \9875 , RIbe2b5b8_126);
nand \U$16201 ( \16454 , \16452 , \16453 );
and \U$16202 ( \16455 , \16454 , \13167 );
not \U$16203 ( \16456 , \16454 );
and \U$16204 ( \16457 , \16456 , \6992 );
nor \U$16205 ( \16458 , \16455 , \16457 );
and \U$16206 ( \16459 , \16449 , \16458 );
not \U$16207 ( \16460 , \16449 );
not \U$16208 ( \16461 , \16458 );
and \U$16209 ( \16462 , \16460 , \16461 );
nor \U$16210 ( \16463 , \16459 , \16462 );
xor \U$16211 ( \16464 , \16430 , \16463 );
xor \U$16212 ( \16465 , \16392 , \16464 );
xor \U$16213 ( \16466 , \16356 , \16465 );
xor \U$16214 ( \16467 , \16326 , \16466 );
not \U$16215 ( \16468 , \16094 );
nand \U$16216 ( \16469 , \16468 , \16122 );
and \U$16217 ( \16470 , \16087 , \16469 );
nor \U$16218 ( \16471 , \16468 , \16122 );
nor \U$16219 ( \16472 , \16470 , \16471 );
xor \U$16220 ( \16473 , \16073 , \16077 );
and \U$16221 ( \16474 , \16473 , \16083 );
and \U$16222 ( \16475 , \16073 , \16077 );
or \U$16223 ( \16476 , \16474 , \16475 );
nand \U$16224 ( \16477 , \16472 , \16476 );
and \U$16225 ( \16478 , \16467 , \16477 );
nor \U$16226 ( \16479 , \16472 , \16476 );
nor \U$16227 ( \16480 , \16478 , \16479 );
not \U$16228 ( \16481 , \16212 );
not \U$16229 ( \16482 , \16481 );
not \U$16230 ( \16483 , \16324 );
or \U$16231 ( \16484 , \16482 , \16483 );
not \U$16232 ( \16485 , \16212 );
not \U$16233 ( \16486 , \16323 );
or \U$16234 ( \16487 , \16485 , \16486 );
nand \U$16235 ( \16488 , \16487 , \16230 );
nand \U$16236 ( \16489 , \16484 , \16488 );
not \U$16237 ( \16490 , \16489 );
xor \U$16238 ( \16491 , \16170 , \16174 );
and \U$16239 ( \16492 , \16491 , \16179 );
and \U$16240 ( \16493 , \16170 , \16174 );
or \U$16241 ( \16494 , \16492 , \16493 );
not \U$16242 ( \16495 , \16494 );
not \U$16243 ( \16496 , \16495 );
and \U$16244 ( \16497 , \16490 , \16496 );
and \U$16245 ( \16498 , \16489 , \16495 );
nor \U$16246 ( \16499 , \16497 , \16498 );
xor \U$16247 ( \16500 , \16351 , \16355 );
and \U$16248 ( \16501 , \16500 , \16465 );
and \U$16249 ( \16502 , \16351 , \16355 );
or \U$16250 ( \16503 , \16501 , \16502 );
xnor \U$16251 ( \16504 , \16499 , \16503 );
nor \U$16252 ( \16505 , \16480 , \16504 );
not \U$16253 ( \16506 , \16505 );
nand \U$16254 ( \16507 , \16480 , \16504 );
nand \U$16255 ( \16508 , \16506 , \16507 );
not \U$16256 ( \16509 , \15849 );
not \U$16257 ( \16510 , \15822 );
or \U$16258 ( \16511 , \16509 , \16510 );
not \U$16259 ( \16512 , \15850 );
not \U$16260 ( \16513 , \15853 );
or \U$16261 ( \16514 , \16512 , \16513 );
nand \U$16262 ( \16515 , \16514 , \16066 );
nand \U$16263 ( \16516 , \16511 , \16515 );
xor \U$16264 ( \16517 , \16180 , \16325 );
and \U$16265 ( \16518 , \16517 , \16466 );
and \U$16266 ( \16519 , \16180 , \16325 );
or \U$16267 ( \16520 , \16518 , \16519 );
xor \U$16268 ( \16521 , \16516 , \16520 );
not \U$16269 ( \16522 , \16218 );
not \U$16270 ( \16523 , \16522 );
not \U$16271 ( \16524 , \16229 );
or \U$16272 ( \16525 , \16523 , \16524 );
nand \U$16273 ( \16526 , \16525 , \16224 );
not \U$16274 ( \16527 , \16229 );
nand \U$16275 ( \16528 , \16527 , \16218 );
nand \U$16276 ( \16529 , \16526 , \16528 );
not \U$16277 ( \16530 , \16194 );
not \U$16278 ( \16531 , \16185 );
or \U$16279 ( \16532 , \16530 , \16531 );
not \U$16280 ( \16533 , \16184 );
not \U$16281 ( \16534 , \16195 );
or \U$16282 ( \16535 , \16533 , \16534 );
nand \U$16283 ( \16536 , \16535 , \16207 );
nand \U$16284 ( \16537 , \16532 , \16536 );
not \U$16285 ( \16538 , \16537 );
xor \U$16286 ( \16539 , \16529 , \16538 );
buf \U$16287 ( \16540 , \16260 );
nor \U$16288 ( \16541 , \16318 , \16540 );
or \U$16289 ( \16542 , \16541 , \16288 );
nand \U$16290 ( \16543 , \16318 , \16540 );
nand \U$16291 ( \16544 , \16542 , \16543 );
xor \U$16292 ( \16545 , \16539 , \16544 );
not \U$16293 ( \16546 , \16545 );
not \U$16294 ( \16547 , \16546 );
not \U$16295 ( \16548 , \16266 );
not \U$16296 ( \16549 , \16548 );
not \U$16297 ( \16550 , \16287 );
or \U$16298 ( \16551 , \16549 , \16550 );
not \U$16299 ( \16552 , \16276 );
nand \U$16300 ( \16553 , \16551 , \16552 );
not \U$16301 ( \16554 , \16287 );
nand \U$16302 ( \16555 , \16554 , \16266 );
nand \U$16303 ( \16556 , \16553 , \16555 );
not \U$16304 ( \16557 , RIbe2ab68_104);
not \U$16305 ( \16558 , \3284 );
or \U$16306 ( \16559 , \16557 , \16558 );
nand \U$16307 ( \16560 , \3458 , RIbe2aaf0_103);
nand \U$16308 ( \16561 , \16559 , \16560 );
and \U$16309 ( \16562 , \16561 , \2887 );
not \U$16310 ( \16563 , \16561 );
and \U$16311 ( \16564 , \16563 , \3290 );
nor \U$16312 ( \16565 , \16562 , \16564 );
not \U$16313 ( \16566 , \16565 );
not \U$16314 ( \16567 , RIbe2b630_127);
not \U$16315 ( \16568 , \4021 );
or \U$16316 ( \16569 , \16567 , \16568 );
nand \U$16317 ( \16570 , \7438 , RIbe2b018_114);
nand \U$16318 ( \16571 , \16569 , \16570 );
and \U$16319 ( \16572 , \16571 , \3471 );
not \U$16320 ( \16573 , \16571 );
and \U$16321 ( \16574 , \16573 , \3698 );
nor \U$16322 ( \16575 , \16572 , \16574 );
not \U$16323 ( \16576 , \16575 );
or \U$16324 ( \16577 , \16566 , \16576 );
or \U$16325 ( \16578 , \16565 , \16575 );
nand \U$16326 ( \16579 , \16577 , \16578 );
xor \U$16327 ( \16580 , \16556 , \16579 );
not \U$16328 ( \16581 , \16580 );
not \U$16329 ( \16582 , \16581 );
nor \U$16330 ( \16583 , \16343 , \3290 );
or \U$16331 ( \16584 , \16336 , \16583 );
nand \U$16332 ( \16585 , \16343 , \3290 );
nand \U$16333 ( \16586 , \16584 , \16585 );
not \U$16334 ( \16587 , \16586 );
not \U$16335 ( \16588 , \16400 );
nand \U$16336 ( \16589 , \16425 , \16410 );
not \U$16337 ( \16590 , \16589 );
or \U$16338 ( \16591 , \16588 , \16590 );
nand \U$16339 ( \16592 , \16428 , \16413 );
nand \U$16340 ( \16593 , \16591 , \16592 );
not \U$16341 ( \16594 , \16593 );
not \U$16342 ( \16595 , \16594 );
or \U$16343 ( \16596 , \16587 , \16595 );
not \U$16344 ( \16597 , \16586 );
nand \U$16345 ( \16598 , \16597 , \16593 );
nand \U$16346 ( \16599 , \16596 , \16598 );
nand \U$16347 ( \16600 , \16391 , \16370 );
and \U$16348 ( \16601 , \16600 , \16379 );
nor \U$16349 ( \16602 , \16391 , \16370 );
nor \U$16350 ( \16603 , \16601 , \16602 );
and \U$16351 ( \16604 , \16599 , \16603 );
not \U$16352 ( \16605 , \16599 );
not \U$16353 ( \16606 , \16603 );
and \U$16354 ( \16607 , \16605 , \16606 );
nor \U$16355 ( \16608 , \16604 , \16607 );
not \U$16356 ( \16609 , \16608 );
not \U$16357 ( \16610 , \16609 );
or \U$16358 ( \16611 , \16582 , \16610 );
nand \U$16359 ( \16612 , \16608 , \16580 );
nand \U$16360 ( \16613 , \16611 , \16612 );
not \U$16361 ( \16614 , \16439 );
not \U$16362 ( \16615 , \16448 );
not \U$16363 ( \16616 , \16615 );
or \U$16364 ( \16617 , \16614 , \16616 );
or \U$16365 ( \16618 , \16439 , \16615 );
nand \U$16366 ( \16619 , \16618 , \16458 );
nand \U$16367 ( \16620 , \16617 , \16619 );
xor \U$16368 ( \16621 , \16240 , \16249 );
and \U$16369 ( \16622 , \16621 , \16259 );
and \U$16370 ( \16623 , \16240 , \16249 );
or \U$16371 ( \16624 , \16622 , \16623 );
xor \U$16372 ( \16625 , \16620 , \16624 );
or \U$16373 ( \16626 , \16307 , \16298 );
and \U$16374 ( \16627 , \16626 , \16317 );
and \U$16375 ( \16628 , \16298 , \16307 );
nor \U$16376 ( \16629 , \16627 , \16628 );
xnor \U$16377 ( \16630 , \16625 , \16629 );
xnor \U$16378 ( \16631 , \16613 , \16630 );
not \U$16379 ( \16632 , \16631 );
or \U$16380 ( \16633 , \16547 , \16632 );
not \U$16381 ( \16634 , \16631 );
nand \U$16382 ( \16635 , \16634 , \16545 );
nand \U$16383 ( \16636 , \16633 , \16635 );
not \U$16384 ( \16637 , RIbe2a208_84);
not \U$16385 ( \16638 , \6535 );
or \U$16386 ( \16639 , \16637 , \16638 );
nand \U$16387 ( \16640 , \10348 , RIbe2a190_83);
nand \U$16388 ( \16641 , \16639 , \16640 );
not \U$16389 ( \16642 , \16641 );
not \U$16390 ( \16643 , \7546 );
and \U$16391 ( \16644 , \16642 , \16643 );
and \U$16392 ( \16645 , \16641 , \6551 );
nor \U$16393 ( \16646 , \16644 , \16645 );
not \U$16394 ( \16647 , \16646 );
not \U$16395 ( \16648 , \16647 );
not \U$16396 ( \16649 , RIbe2a5c8_92);
not \U$16397 ( \16650 , \7941 );
or \U$16398 ( \16651 , \16649 , \16650 );
nand \U$16399 ( \16652 , \13436 , RIbe2a550_91);
nand \U$16400 ( \16653 , \16651 , \16652 );
and \U$16401 ( \16654 , \16653 , \7948 );
not \U$16402 ( \16655 , \16653 );
and \U$16403 ( \16656 , \16655 , \14262 );
nor \U$16404 ( \16657 , \16654 , \16656 );
not \U$16405 ( \16658 , \16657 );
not \U$16406 ( \16659 , \16658 );
or \U$16407 ( \16660 , \16648 , \16659 );
nand \U$16408 ( \16661 , \16657 , \16646 );
nand \U$16409 ( \16662 , \16660 , \16661 );
not \U$16410 ( \16663 , RIbe2b090_115);
not \U$16411 ( \16664 , \6139 );
or \U$16412 ( \16665 , \16663 , \16664 );
nand \U$16413 ( \16666 , \7528 , RIbe2a280_85);
nand \U$16414 ( \16667 , \16665 , \16666 );
and \U$16415 ( \16668 , \16667 , \7534 );
not \U$16416 ( \16669 , \16667 );
and \U$16417 ( \16670 , \16669 , \5740 );
nor \U$16418 ( \16671 , \16668 , \16670 );
xnor \U$16419 ( \16672 , \16662 , \16671 );
not \U$16420 ( \16673 , RIbe2a370_87);
not \U$16421 ( \16674 , \7974 );
or \U$16422 ( \16675 , \16673 , \16674 );
nand \U$16423 ( \16676 , \7981 , RIbe2a2f8_86);
nand \U$16424 ( \16677 , \16675 , \16676 );
and \U$16425 ( \16678 , \16677 , \14299 );
not \U$16426 ( \16679 , \16677 );
and \U$16427 ( \16680 , \16679 , \6948 );
nor \U$16428 ( \16681 , \16678 , \16680 );
not \U$16429 ( \16682 , \16681 );
not \U$16430 ( \16683 , RIbe2b5b8_126);
not \U$16431 ( \16684 , \6980 );
or \U$16432 ( \16685 , \16683 , \16684 );
nand \U$16433 ( \16686 , \9875 , RIbe2a3e8_88);
nand \U$16434 ( \16687 , \16685 , \16686 );
not \U$16435 ( \16688 , \16687 );
not \U$16436 ( \16689 , \7301 );
and \U$16437 ( \16690 , \16688 , \16689 );
and \U$16438 ( \16691 , \16687 , \6992 );
nor \U$16439 ( \16692 , \16690 , \16691 );
not \U$16440 ( \16693 , \16692 );
or \U$16441 ( \16694 , \16682 , \16693 );
or \U$16442 ( \16695 , \16681 , \16692 );
nand \U$16443 ( \16696 , \16694 , \16695 );
not \U$16444 ( \16697 , RIbe2a988_100);
not \U$16445 ( \16698 , \6958 );
or \U$16446 ( \16699 , \16697 , \16698 );
nand \U$16447 ( \16700 , \7653 , RIbe2a910_99);
nand \U$16448 ( \16701 , \16699 , \16700 );
and \U$16449 ( \16702 , \16701 , \7293 );
not \U$16450 ( \16703 , \16701 );
and \U$16451 ( \16704 , \16703 , \6569 );
nor \U$16452 ( \16705 , \16702 , \16704 );
xnor \U$16453 ( \16706 , \16696 , \16705 );
xor \U$16454 ( \16707 , \16672 , \16706 );
not \U$16455 ( \16708 , RIbe2b1f8_118);
not \U$16456 ( \16709 , \4829 );
or \U$16457 ( \16710 , \16708 , \16709 );
nand \U$16458 ( \16711 , \5052 , RIbe2b180_117);
nand \U$16459 ( \16712 , \16710 , \16711 );
and \U$16460 ( \16713 , \16712 , \4592 );
not \U$16461 ( \16714 , \16712 );
and \U$16462 ( \16715 , \16714 , \4586 );
nor \U$16463 ( \16716 , \16713 , \16715 );
not \U$16464 ( \16717 , \16716 );
not \U$16465 ( \16718 , RIbe2b270_119);
not \U$16466 ( \16719 , \6630 );
or \U$16467 ( \16720 , \16718 , \16719 );
nand \U$16468 ( \16721 , \14239 , RIbe2b108_116);
nand \U$16469 ( \16722 , \16720 , \16721 );
not \U$16470 ( \16723 , \16722 );
not \U$16471 ( \16724 , \5754 );
and \U$16472 ( \16725 , \16723 , \16724 );
and \U$16473 ( \16726 , \16722 , \5754 );
nor \U$16474 ( \16727 , \16725 , \16726 );
not \U$16475 ( \16728 , \16727 );
not \U$16476 ( \16729 , \16728 );
or \U$16477 ( \16730 , \16717 , \16729 );
not \U$16478 ( \16731 , \16716 );
nand \U$16479 ( \16732 , \16727 , \16731 );
nand \U$16480 ( \16733 , \16730 , \16732 );
not \U$16481 ( \16734 , RIbe2afa0_113);
not \U$16482 ( \16735 , \5058 );
or \U$16483 ( \16736 , \16734 , \16735 );
nand \U$16484 ( \16737 , \7858 , RIbe2af28_112);
nand \U$16485 ( \16738 , \16736 , \16737 );
xor \U$16486 ( \16739 , \16738 , \4323 );
and \U$16487 ( \16740 , \16733 , \16739 );
not \U$16488 ( \16741 , \16733 );
not \U$16489 ( \16742 , \16739 );
and \U$16490 ( \16743 , \16741 , \16742 );
nor \U$16491 ( \16744 , \16740 , \16743 );
xor \U$16492 ( \16745 , \16707 , \16744 );
not \U$16493 ( \16746 , \16745 );
not \U$16494 ( \16747 , RIbe27f58_10);
not \U$16495 ( \16748 , \14534 );
or \U$16496 ( \16749 , \16747 , \16748 );
nand \U$16497 ( \16750 , RIbe27e68_8, \12735 );
nand \U$16498 ( \16751 , \16749 , \16750 );
and \U$16499 ( \16752 , \16751 , \14543 );
not \U$16500 ( \16753 , \16751 );
not \U$16501 ( \16754 , \14542 );
and \U$16502 ( \16755 , \16753 , \16754 );
nor \U$16503 ( \16756 , \16752 , \16755 );
not \U$16504 ( \16757 , \16756 );
not \U$16505 ( \16758 , RIbe28ed0_43);
and \U$16506 ( \16759 , \12703 , \12704 );
not \U$16507 ( \16760 , \16759 );
or \U$16508 ( \16761 , \16758 , \16760 );
nand \U$16509 ( \16762 , \13727 , RIbe27fd0_11);
nand \U$16510 ( \16763 , \16761 , \16762 );
and \U$16511 ( \16764 , \16763 , \12716 );
not \U$16512 ( \16765 , \16763 );
and \U$16513 ( \16766 , \16765 , \12723 );
nor \U$16514 ( \16767 , \16764 , \16766 );
not \U$16515 ( \16768 , \16767 );
or \U$16516 ( \16769 , \16757 , \16768 );
not \U$16517 ( \16770 , \16756 );
not \U$16518 ( \16771 , \16767 );
nand \U$16519 ( \16772 , \16770 , \16771 );
nand \U$16520 ( \16773 , \16769 , \16772 );
not \U$16521 ( \16774 , \12753 );
not \U$16522 ( \16775 , \7775 );
and \U$16523 ( \16776 , \16774 , \16775 );
and \U$16524 ( \16777 , \12765 , RIbe29bf0_71);
nor \U$16525 ( \16778 , \16776 , \16777 );
and \U$16526 ( \16779 , \16778 , \12769 );
not \U$16527 ( \16780 , \16778 );
and \U$16528 ( \16781 , \16780 , \12774 );
nor \U$16529 ( \16782 , \16779 , \16781 );
xnor \U$16530 ( \16783 , \16773 , \16782 );
not \U$16531 ( \16784 , RIbe28408_20);
not \U$16532 ( \16785 , \13690 );
or \U$16533 ( \16786 , \16784 , \16785 );
nand \U$16534 ( \16787 , RIbe28390_19, RIbe2ae38_110);
nand \U$16535 ( \16788 , \16786 , \16787 );
xor \U$16536 ( \16789 , \16788 , RIbe2aeb0_111);
not \U$16537 ( \16790 , RIbe287c8_28);
not \U$16538 ( \16791 , \12786 );
or \U$16539 ( \16792 , \16790 , \16791 );
nand \U$16540 ( \16793 , \12794 , RIbe28480_21);
nand \U$16541 ( \16794 , \16792 , \16793 );
and \U$16542 ( \16795 , \16794 , \14336 );
not \U$16543 ( \16796 , \16794 );
and \U$16544 ( \16797 , \16796 , \14335 );
nor \U$16545 ( \16798 , \16795 , \16797 );
xor \U$16546 ( \16799 , \16789 , \16798 );
not \U$16547 ( \16800 , RIbe28660_25);
not \U$16548 ( \16801 , \12831 );
or \U$16549 ( \16802 , \16800 , \16801 );
nand \U$16550 ( \16803 , \13012 , RIbe285e8_24);
nand \U$16551 ( \16804 , \16802 , \16803 );
and \U$16552 ( \16805 , \16804 , \13705 );
not \U$16553 ( \16806 , \16804 );
and \U$16554 ( \16807 , \16806 , \12823 );
nor \U$16555 ( \16808 , \16805 , \16807 );
xnor \U$16556 ( \16809 , \16799 , \16808 );
xor \U$16557 ( \16810 , \16783 , \16809 );
not \U$16558 ( \16811 , RIbe29fb0_79);
not \U$16559 ( \16812 , \10936 );
or \U$16560 ( \16813 , \16811 , \16812 );
nand \U$16561 ( \16814 , \14511 , RIbe29e48_76);
nand \U$16562 ( \16815 , \16813 , \16814 );
xor \U$16563 ( \16816 , \16815 , \10943 );
not \U$16564 ( \16817 , RIbe29dd0_75);
not \U$16565 ( \16818 , \15205 );
or \U$16566 ( \16819 , \16817 , \16818 );
nand \U$16567 ( \16820 , \13669 , RIbe29c68_72);
nand \U$16568 ( \16821 , \16819 , \16820 );
not \U$16569 ( \16822 , \16821 );
not \U$16570 ( \16823 , \12960 );
and \U$16571 ( \16824 , \16822 , \16823 );
and \U$16572 ( \16825 , \16821 , \12957 );
nor \U$16573 ( \16826 , \16824 , \16825 );
xor \U$16574 ( \16827 , \16816 , \16826 );
not \U$16575 ( \16828 , RIbe2acd0_107);
not \U$16576 ( \16829 , \10916 );
or \U$16577 ( \16830 , \16828 , \16829 );
nand \U$16578 ( \16831 , \15228 , RIbe2a028_80);
nand \U$16579 ( \16832 , \16830 , \16831 );
not \U$16580 ( \16833 , \16832 );
not \U$16581 ( \16834 , \13650 );
and \U$16582 ( \16835 , \16833 , \16834 );
and \U$16583 ( \16836 , \16832 , \7971 );
nor \U$16584 ( \16837 , \16835 , \16836 );
xor \U$16585 ( \16838 , \16827 , \16837 );
xor \U$16586 ( \16839 , \16810 , \16838 );
or \U$16587 ( \16840 , \16463 , \16392 );
nand \U$16588 ( \16841 , \16840 , \16430 );
nand \U$16589 ( \16842 , \16463 , \16392 );
nand \U$16590 ( \16843 , \16841 , \16842 );
xnor \U$16591 ( \16844 , \16839 , \16843 );
not \U$16592 ( \16845 , \16844 );
or \U$16593 ( \16846 , \16746 , \16845 );
or \U$16594 ( \16847 , \16844 , \16745 );
nand \U$16595 ( \16848 , \16846 , \16847 );
and \U$16596 ( \16849 , \16636 , \16848 );
not \U$16597 ( \16850 , \16636 );
not \U$16598 ( \16851 , \16848 );
and \U$16599 ( \16852 , \16850 , \16851 );
nor \U$16600 ( \16853 , \16849 , \16852 );
xnor \U$16601 ( \16854 , \16521 , \16853 );
xor \U$16602 ( \16855 , \16508 , \16854 );
not \U$16603 ( \16856 , \16855 );
or \U$16604 ( \16857 , \16162 , \16856 );
or \U$16605 ( \16858 , \16855 , \16161 );
nand \U$16606 ( \16859 , \16857 , \16858 );
xor \U$16607 ( \16860 , \16067 , \16131 );
xnor \U$16608 ( \16861 , \16860 , \16158 );
not \U$16609 ( \16862 , \16861 );
xnor \U$16610 ( \16863 , \16472 , \16476 );
not \U$16611 ( \16864 , \16863 );
not \U$16612 ( \16865 , \16467 );
or \U$16613 ( \16866 , \16864 , \16865 );
or \U$16614 ( \16867 , \16863 , \16467 );
nand \U$16615 ( \16868 , \16866 , \16867 );
nand \U$16616 ( \16869 , \16862 , \16868 );
xor \U$16617 ( \16870 , \16859 , \16869 );
xor \U$16618 ( \16871 , \15407 , \15411 );
and \U$16619 ( \16872 , \16871 , \15746 );
and \U$16620 ( \16873 , \15407 , \15411 );
or \U$16621 ( \16874 , \16872 , \16873 );
not \U$16622 ( \16875 , \16874 );
not \U$16623 ( \16876 , \16130 );
not \U$16624 ( \16877 , \16084 );
and \U$16625 ( \16878 , \16876 , \16877 );
and \U$16626 ( \16879 , \16084 , \16130 );
nor \U$16627 ( \16880 , \16878 , \16879 );
not \U$16628 ( \16881 , \16880 );
not \U$16629 ( \16882 , \16881 );
xor \U$16630 ( \16883 , \16142 , \16148 );
xor \U$16631 ( \16884 , \16883 , \16155 );
not \U$16632 ( \16885 , \16884 );
nand \U$16633 ( \16886 , \16882 , \16885 );
not \U$16634 ( \16887 , \16886 );
or \U$16635 ( \16888 , \16875 , \16887 );
not \U$16636 ( \16889 , \16885 );
nand \U$16637 ( \16890 , \16889 , \16881 );
nand \U$16638 ( \16891 , \16888 , \16890 );
not \U$16639 ( \16892 , \16891 );
not \U$16640 ( \16893 , \16868 );
not \U$16641 ( \16894 , \16861 );
or \U$16642 ( \16895 , \16893 , \16894 );
or \U$16643 ( \16896 , \16868 , \16861 );
nand \U$16644 ( \16897 , \16895 , \16896 );
not \U$16645 ( \16898 , \16897 );
not \U$16646 ( \16899 , \16898 );
or \U$16647 ( \16900 , \16892 , \16899 );
not \U$16648 ( \16901 , \16891 );
nand \U$16649 ( \16902 , \16901 , \16897 );
nand \U$16650 ( \16903 , \16900 , \16902 );
and \U$16651 ( \16904 , \16884 , \16880 );
not \U$16652 ( \16905 , \16884 );
and \U$16653 ( \16906 , \16905 , \16881 );
nor \U$16654 ( \16907 , \16904 , \16906 );
xor \U$16655 ( \16908 , \16907 , \16874 );
not \U$16656 ( \16909 , \16908 );
not \U$16657 ( \16910 , \16909 );
xor \U$16658 ( \16911 , \15398 , \15402 );
and \U$16659 ( \16912 , \16911 , \15747 );
and \U$16660 ( \16913 , \15398 , \15402 );
or \U$16661 ( \16914 , \16912 , \16913 );
not \U$16662 ( \16915 , \16914 );
not \U$16663 ( \16916 , \16915 );
or \U$16664 ( \16917 , \16910 , \16916 );
nand \U$16665 ( \16918 , \16908 , \16914 );
nand \U$16666 ( \16919 , \16917 , \16918 );
nand \U$16667 ( \16920 , \16903 , \16919 );
nor \U$16668 ( \16921 , \16870 , \16920 );
nand \U$16669 ( \16922 , \15771 , \16921 );
not \U$16670 ( \16923 , \16903 );
and \U$16671 ( \16924 , \15384 , \15748 );
not \U$16672 ( \16925 , \16924 );
not \U$16673 ( \16926 , \16919 );
or \U$16674 ( \16927 , \16925 , \16926 );
not \U$16675 ( \16928 , \16908 );
buf \U$16676 ( \16929 , \16914 );
nand \U$16677 ( \16930 , \16928 , \16929 );
nand \U$16678 ( \16931 , \16927 , \16930 );
not \U$16679 ( \16932 , \16931 );
or \U$16680 ( \16933 , \16923 , \16932 );
nand \U$16681 ( \16934 , \16897 , \16891 );
nand \U$16682 ( \16935 , \16933 , \16934 );
not \U$16683 ( \16936 , \16870 );
nand \U$16684 ( \16937 , \16935 , \16936 );
not \U$16685 ( \16938 , \16869 );
nand \U$16686 ( \16939 , \16938 , \16859 );
nand \U$16687 ( \16940 , \16922 , \16937 , \16939 );
not \U$16688 ( \16941 , \16940 );
xnor \U$16689 ( \16942 , \14678 , \14680 );
not \U$16690 ( \16943 , \14470 );
and \U$16691 ( \16944 , \16942 , \16943 );
not \U$16692 ( \16945 , \16942 );
and \U$16693 ( \16946 , \16945 , \14470 );
nor \U$16694 ( \16947 , \16944 , \16946 );
not \U$16695 ( \16948 , \16947 );
not \U$16696 ( \16949 , \16948 );
not \U$16697 ( \16950 , RIbe2acd0_107);
not \U$16698 ( \16951 , \12786 );
or \U$16699 ( \16952 , \16950 , \16951 );
nand \U$16700 ( \16953 , RIbe2a028_80, \12890 );
nand \U$16701 ( \16954 , \16952 , \16953 );
and \U$16702 ( \16955 , \16954 , \12998 );
not \U$16703 ( \16956 , \16954 );
and \U$16704 ( \16957 , \16956 , \16334 );
nor \U$16705 ( \16958 , \16955 , \16957 );
not \U$16706 ( \16959 , RIbe29fb0_79);
not \U$16707 ( \16960 , \13004 );
or \U$16708 ( \16961 , \16959 , \16960 );
nand \U$16709 ( \16962 , RIbe29e48_76, RIbe2ae38_110);
nand \U$16710 ( \16963 , \16961 , \16962 );
not \U$16711 ( \16964 , RIbe2aeb0_111);
xor \U$16712 ( \16965 , \16963 , \16964 );
nand \U$16713 ( \16966 , \16958 , \16965 );
not \U$16714 ( \16967 , \12823 );
not \U$16715 ( \16968 , RIbe2a370_87);
not \U$16716 ( \16969 , \13010 );
or \U$16717 ( \16970 , \16968 , \16969 );
nand \U$16718 ( \16971 , \12835 , RIbe2a2f8_86);
nand \U$16719 ( \16972 , \16970 , \16971 );
not \U$16720 ( \16973 , \16972 );
or \U$16721 ( \16974 , \16967 , \16973 );
or \U$16722 ( \16975 , \16972 , \12823 );
nand \U$16723 ( \16976 , \16974 , \16975 );
and \U$16724 ( \16977 , \16966 , \16976 );
nor \U$16725 ( \16978 , \16958 , \16965 );
nor \U$16726 ( \16979 , \16977 , \16978 );
not \U$16727 ( \16980 , \16979 );
not \U$16728 ( \16981 , \16980 );
not \U$16729 ( \16982 , RIbe2b090_115);
not \U$16730 ( \16983 , \13024 );
or \U$16731 ( \16984 , \16982 , \16983 );
nand \U$16732 ( \16985 , \12212 , RIbe2a280_85);
nand \U$16733 ( \16986 , \16984 , \16985 );
and \U$16734 ( \16987 , \16986 , \13030 );
not \U$16735 ( \16988 , \16986 );
and \U$16736 ( \16989 , \16988 , \9904 );
nor \U$16737 ( \16990 , \16987 , \16989 );
and \U$16738 ( \16991 , \8278 , RIbe2b270_119);
and \U$16739 ( \16992 , \13380 , RIbe2b108_116);
nor \U$16740 ( \16993 , \16991 , \16992 );
not \U$16741 ( \16994 , \8077 );
and \U$16742 ( \16995 , \16993 , \16994 );
not \U$16743 ( \16996 , \16993 );
and \U$16744 ( \16997 , \16996 , \8077 );
nor \U$16745 ( \16998 , \16995 , \16997 );
and \U$16746 ( \16999 , \16990 , \16998 );
not \U$16747 ( \17000 , RIbe2a208_84);
not \U$16748 ( \17001 , \13049 );
or \U$16749 ( \17002 , \17000 , \17001 );
nand \U$16750 ( \17003 , \12947 , RIbe2a190_83);
nand \U$16751 ( \17004 , \17002 , \17003 );
buf \U$16752 ( \17005 , \12956 );
and \U$16753 ( \17006 , \17004 , \17005 );
not \U$16754 ( \17007 , \17004 );
and \U$16755 ( \17008 , \17007 , \12195 );
nor \U$16756 ( \17009 , \17006 , \17008 );
nor \U$16757 ( \17010 , \16999 , \17009 );
nor \U$16758 ( \17011 , \16998 , \16990 );
nor \U$16759 ( \17012 , \17010 , \17011 );
not \U$16760 ( \17013 , \17012 );
not \U$16761 ( \17014 , \17013 );
or \U$16762 ( \17015 , \16981 , \17014 );
not \U$16763 ( \17016 , \16979 );
not \U$16764 ( \17017 , \17012 );
or \U$16765 ( \17018 , \17016 , \17017 );
not \U$16766 ( \17019 , RIbe2b5b8_126);
not \U$16767 ( \17020 , \12732 );
or \U$16768 ( \17021 , \17019 , \17020 );
nand \U$16769 ( \17022 , \13077 , RIbe2a3e8_88);
nand \U$16770 ( \17023 , \17021 , \17022 );
and \U$16771 ( \17024 , \17023 , \12746 );
not \U$16772 ( \17025 , \17023 );
and \U$16773 ( \17026 , \17025 , \14077 );
nor \U$16774 ( \17027 , \17024 , \17026 );
not \U$16775 ( \17028 , RIbe2a988_100);
not \U$16776 ( \17029 , \14523 );
or \U$16777 ( \17030 , \17028 , \17029 );
nand \U$16778 ( \17031 , \13728 , RIbe2a910_99);
nand \U$16779 ( \17032 , \17030 , \17031 );
and \U$16780 ( \17033 , \17032 , \13583 );
not \U$16781 ( \17034 , \17032 );
and \U$16782 ( \17035 , \17034 , \12879 );
nor \U$16783 ( \17036 , \17033 , \17035 );
nand \U$16784 ( \17037 , \17027 , \17036 );
not \U$16785 ( \17038 , RIbe2a5c8_92);
not \U$16786 ( \17039 , \13738 );
not \U$16787 ( \17040 , \17039 );
not \U$16788 ( \17041 , \17040 );
or \U$16789 ( \17042 , \17038 , \17041 );
not \U$16790 ( \17043 , \12753 );
nand \U$16791 ( \17044 , \17043 , RIbe2a550_91);
nand \U$16792 ( \17045 , \17042 , \17044 );
xnor \U$16793 ( \17046 , \17045 , \12924 );
and \U$16794 ( \17047 , \17037 , \17046 );
nor \U$16795 ( \17048 , \17027 , \17036 );
nor \U$16796 ( \17049 , \17047 , \17048 );
not \U$16797 ( \17050 , \17049 );
nand \U$16798 ( \17051 , \17018 , \17050 );
nand \U$16799 ( \17052 , \17015 , \17051 );
and \U$16800 ( \17053 , \6547 , \14576 );
not \U$16801 ( \17054 , \6547 );
and \U$16802 ( \17055 , \17054 , \14575 );
nor \U$16803 ( \17056 , \17053 , \17055 );
not \U$16804 ( \17057 , \17056 );
not \U$16805 ( \17058 , \14569 );
or \U$16806 ( \17059 , \17057 , \17058 );
or \U$16807 ( \17060 , \17056 , \14569 );
nand \U$16808 ( \17061 , \17059 , \17060 );
xor \U$16809 ( \17062 , \14560 , \14547 );
xor \U$16810 ( \17063 , \17062 , \14531 );
xor \U$16811 ( \17064 , \17061 , \17063 );
xor \U$16812 ( \17065 , \14497 , \14505 );
xor \U$16813 ( \17066 , \17065 , \14517 );
and \U$16814 ( \17067 , \17064 , \17066 );
and \U$16815 ( \17068 , \17061 , \17063 );
or \U$16816 ( \17069 , \17067 , \17068 );
xor \U$16817 ( \17070 , \17052 , \17069 );
xor \U$16818 ( \17071 , \14641 , \14630 );
xnor \U$16819 ( \17072 , \17071 , \14654 );
not \U$16820 ( \17073 , \13167 );
and \U$16821 ( \17074 , \7298 , RIbe2afa0_113);
and \U$16822 ( \17075 , \13792 , RIbe2af28_112);
nor \U$16823 ( \17076 , \17074 , \17075 );
not \U$16824 ( \17077 , \17076 );
or \U$16825 ( \17078 , \17073 , \17077 );
or \U$16826 ( \17079 , \17076 , \7304 );
nand \U$16827 ( \17080 , \17078 , \17079 );
not \U$16828 ( \17081 , RIbe2b630_127);
not \U$16829 ( \17082 , \7954 );
or \U$16830 ( \17083 , \17081 , \17082 );
nand \U$16831 ( \17084 , RIbe2b018_114, \6963 );
nand \U$16832 ( \17085 , \17083 , \17084 );
and \U$16833 ( \17086 , \17085 , \7293 );
not \U$16834 ( \17087 , \17085 );
and \U$16835 ( \17088 , \17087 , \6572 );
nor \U$16836 ( \17089 , \17086 , \17088 );
xor \U$16837 ( \17090 , \17080 , \17089 );
not \U$16838 ( \17091 , RIbe2b1f8_118);
not \U$16839 ( \17092 , \10949 );
or \U$16840 ( \17093 , \17091 , \17092 );
nand \U$16841 ( \17094 , \8269 , RIbe2b180_117);
nand \U$16842 ( \17095 , \17093 , \17094 );
and \U$16843 ( \17096 , \17095 , \14299 );
not \U$16844 ( \17097 , \17095 );
and \U$16845 ( \17098 , \17097 , \7989 );
nor \U$16846 ( \17099 , \17096 , \17098 );
and \U$16847 ( \17100 , \17090 , \17099 );
and \U$16848 ( \17101 , \17080 , \17089 );
or \U$16849 ( \17102 , \17100 , \17101 );
xor \U$16850 ( \17103 , \17072 , \17102 );
xor \U$16851 ( \17104 , \14605 , \14616 );
xnor \U$16852 ( \17105 , \17104 , \14593 );
and \U$16853 ( \17106 , \17103 , \17105 );
and \U$16854 ( \17107 , \17072 , \17102 );
or \U$16855 ( \17108 , \17106 , \17107 );
and \U$16856 ( \17109 , \17070 , \17108 );
and \U$16857 ( \17110 , \17052 , \17069 );
or \U$16858 ( \17111 , \17109 , \17110 );
not \U$16859 ( \17112 , \17111 );
xnor \U$16860 ( \17113 , \13678 , \13748 );
not \U$16861 ( \17114 , \17113 );
not \U$16862 ( \17115 , \13711 );
and \U$16863 ( \17116 , \17114 , \17115 );
and \U$16864 ( \17117 , \13711 , \17113 );
nor \U$16865 ( \17118 , \17116 , \17117 );
and \U$16866 ( \17119 , \17112 , \17118 );
not \U$16867 ( \17120 , \13745 );
not \U$16868 ( \17121 , \13734 );
or \U$16869 ( \17122 , \17120 , \17121 );
nand \U$16870 ( \17123 , \13746 , \13722 );
nand \U$16871 ( \17124 , \17122 , \17123 );
and \U$16872 ( \17125 , \17124 , \13743 );
not \U$16873 ( \17126 , \17124 );
not \U$16874 ( \17127 , \13743 );
and \U$16875 ( \17128 , \17126 , \17127 );
nor \U$16876 ( \17129 , \17125 , \17128 );
not \U$16877 ( \17130 , \17129 );
xor \U$16878 ( \17131 , \13688 , \13695 );
xnor \U$16879 ( \17132 , \17131 , \13708 );
nand \U$16880 ( \17133 , \17130 , \17132 );
not \U$16881 ( \17134 , \17133 );
xor \U$16882 ( \17135 , \14479 , \14482 );
xor \U$16883 ( \17136 , \17135 , \14485 );
not \U$16884 ( \17137 , \17136 );
or \U$16885 ( \17138 , \17134 , \17137 );
not \U$16886 ( \17139 , \17132 );
nand \U$16887 ( \17140 , \17139 , \17129 );
nand \U$16888 ( \17141 , \17138 , \17140 );
not \U$16889 ( \17142 , \17141 );
nor \U$16890 ( \17143 , \17119 , \17142 );
nor \U$16891 ( \17144 , \17112 , \17118 );
nor \U$16892 ( \17145 , \17143 , \17144 );
not \U$16893 ( \17146 , \17145 );
or \U$16894 ( \17147 , \16949 , \17146 );
not \U$16895 ( \17148 , \17145 );
nand \U$16896 ( \17149 , \17148 , \16947 );
nand \U$16897 ( \17150 , \17147 , \17149 );
xnor \U$16898 ( \17151 , \14689 , \14691 );
not \U$16899 ( \17152 , \17151 );
and \U$16900 ( \17153 , \17150 , \17152 );
not \U$16901 ( \17154 , \17150 );
and \U$16902 ( \17155 , \17154 , \17151 );
nor \U$16903 ( \17156 , \17153 , \17155 );
not \U$16904 ( \17157 , \14488 );
not \U$16905 ( \17158 , \14587 );
not \U$16906 ( \17159 , \14672 );
or \U$16907 ( \17160 , \17158 , \17159 );
or \U$16908 ( \17161 , \14672 , \14587 );
nand \U$16909 ( \17162 , \17160 , \17161 );
not \U$16910 ( \17163 , \17162 );
not \U$16911 ( \17164 , \17163 );
or \U$16912 ( \17165 , \17157 , \17164 );
not \U$16913 ( \17166 , \14488 );
nand \U$16914 ( \17167 , \17166 , \17162 );
nand \U$16915 ( \17168 , \17165 , \17167 );
not \U$16916 ( \17169 , \17168 );
not \U$16917 ( \17170 , \17118 );
not \U$16918 ( \17171 , \17170 );
not \U$16919 ( \17172 , \17142 );
or \U$16920 ( \17173 , \17171 , \17172 );
nand \U$16921 ( \17174 , \17141 , \17118 );
nand \U$16922 ( \17175 , \17173 , \17174 );
xor \U$16923 ( \17176 , \17175 , \17112 );
nor \U$16924 ( \17177 , \17169 , \17176 );
not \U$16925 ( \17178 , \17177 );
xor \U$16926 ( \17179 , \14455 , \14452 );
xnor \U$16927 ( \17180 , \17179 , \14466 );
not \U$16928 ( \17181 , \14620 );
buf \U$16929 ( \17182 , \14657 );
not \U$16930 ( \17183 , \17182 );
and \U$16931 ( \17184 , \17181 , \17183 );
and \U$16932 ( \17185 , \14620 , \17182 );
nor \U$16933 ( \17186 , \17184 , \17185 );
xor \U$16934 ( \17187 , \17186 , \14668 );
not \U$16935 ( \17188 , RIbe2ab68_104);
not \U$16936 ( \17189 , \6592 );
or \U$16937 ( \17190 , \17188 , \17189 );
nand \U$16938 ( \17191 , \6596 , RIbe2aaf0_103);
nand \U$16939 ( \17192 , \17190 , \17191 );
not \U$16940 ( \17193 , \17192 );
not \U$16941 ( \17194 , \14666 );
and \U$16942 ( \17195 , \17193 , \17194 );
and \U$16943 ( \17196 , \17192 , \6583 );
nor \U$16944 ( \17197 , \17195 , \17196 );
not \U$16945 ( \17198 , \17197 );
not \U$16946 ( \17199 , RIbe2aaf0_103);
not \U$16947 ( \17200 , \6958 );
or \U$16948 ( \17201 , \17199 , \17200 );
nand \U$16949 ( \17202 , \7653 , RIbe2b630_127);
nand \U$16950 ( \17203 , \17201 , \17202 );
and \U$16951 ( \17204 , \17203 , \7293 );
not \U$16952 ( \17205 , \17203 );
and \U$16953 ( \17206 , \17205 , \6572 );
nor \U$16954 ( \17207 , \17204 , \17206 );
nand \U$16955 ( \17208 , \13436 , RIbe2ab68_104);
and \U$16956 ( \17209 , \17208 , \6601 );
not \U$16957 ( \17210 , \17208 );
and \U$16958 ( \17211 , \17210 , \8957 );
or \U$16959 ( \17212 , \17209 , \17211 );
nand \U$16960 ( \17213 , \17207 , \17212 );
not \U$16961 ( \17214 , \17213 );
or \U$16962 ( \17215 , \17198 , \17214 );
not \U$16963 ( \17216 , RIbe2af28_112);
not \U$16964 ( \17217 , \10949 );
or \U$16965 ( \17218 , \17216 , \17217 );
nand \U$16966 ( \17219 , RIbe2b1f8_118, \9891 );
nand \U$16967 ( \17220 , \17218 , \17219 );
and \U$16968 ( \17221 , \17220 , \7984 );
not \U$16969 ( \17222 , \17220 );
and \U$16970 ( \17223 , \17222 , \9896 );
nor \U$16971 ( \17224 , \17221 , \17223 );
not \U$16972 ( \17225 , \17224 );
buf \U$16973 ( \17226 , \17225 );
and \U$16974 ( \17227 , \9909 , RIbe2b180_117);
not \U$16975 ( \17228 , \13379 );
and \U$16976 ( \17229 , \17228 , RIbe2b270_119);
nor \U$16977 ( \17230 , \17227 , \17229 );
and \U$16978 ( \17231 , \17230 , \8077 );
not \U$16979 ( \17232 , \17230 );
and \U$16980 ( \17233 , \17232 , \13649 );
nor \U$16981 ( \17234 , \17231 , \17233 );
not \U$16982 ( \17235 , \17234 );
not \U$16983 ( \17236 , \17235 );
or \U$16984 ( \17237 , \17226 , \17236 );
and \U$16985 ( \17238 , \7299 , RIbe2b018_114);
and \U$16986 ( \17239 , \6985 , RIbe2afa0_113);
nor \U$16987 ( \17240 , \17238 , \17239 );
and \U$16988 ( \17241 , \17240 , \7660 );
not \U$16989 ( \17242 , \17240 );
and \U$16990 ( \17243 , \17242 , \7301 );
nor \U$16991 ( \17244 , \17241 , \17243 );
not \U$16992 ( \17245 , \17244 );
nand \U$16993 ( \17246 , \17237 , \17245 );
nand \U$16994 ( \17247 , \17226 , \17236 );
nand \U$16995 ( \17248 , \17246 , \17247 );
nand \U$16996 ( \17249 , \17215 , \17248 );
not \U$16997 ( \17250 , \17197 );
nand \U$16998 ( \17251 , \17250 , \17207 , \17212 );
nand \U$16999 ( \17252 , \17249 , \17251 );
not \U$17000 ( \17253 , \17252 );
not \U$17001 ( \17254 , RIbe2a3e8_88);
not \U$17002 ( \17255 , \13590 );
or \U$17003 ( \17256 , \17254 , \17255 );
nand \U$17004 ( \17257 , RIbe2a370_87, \12835 );
nand \U$17005 ( \17258 , \17256 , \17257 );
and \U$17006 ( \17259 , \17258 , \15263 );
not \U$17007 ( \17260 , \17258 );
and \U$17008 ( \17261 , \17260 , \12866 );
nor \U$17009 ( \17262 , \17259 , \17261 );
not \U$17010 ( \17263 , \17262 );
not \U$17011 ( \17264 , \17263 );
not \U$17012 ( \17265 , RIbe2a550_91);
not \U$17013 ( \17266 , \16383 );
or \U$17014 ( \17267 , \17265 , \17266 );
nand \U$17015 ( \17268 , \12711 , RIbe2a988_100);
nand \U$17016 ( \17269 , \17267 , \17268 );
and \U$17017 ( \17270 , \17269 , \13583 );
not \U$17018 ( \17271 , \17269 );
and \U$17019 ( \17272 , \17271 , \12879 );
nor \U$17020 ( \17273 , \17270 , \17272 );
not \U$17021 ( \17274 , \17273 );
not \U$17022 ( \17275 , \17274 );
or \U$17023 ( \17276 , \17264 , \17275 );
nand \U$17024 ( \17277 , \17273 , \17262 );
not \U$17025 ( \17278 , RIbe2a910_99);
not \U$17026 ( \17279 , \12732 );
or \U$17027 ( \17280 , \17278 , \17279 );
nand \U$17028 ( \17281 , \13077 , RIbe2b5b8_126);
nand \U$17029 ( \17282 , \17280 , \17281 );
and \U$17030 ( \17283 , \17282 , \12746 );
not \U$17031 ( \17284 , \17282 );
and \U$17032 ( \17285 , \17284 , \13570 );
nor \U$17033 ( \17286 , \17283 , \17285 );
not \U$17034 ( \17287 , \17286 );
nand \U$17035 ( \17288 , \17277 , \17287 );
nand \U$17036 ( \17289 , \17276 , \17288 );
not \U$17037 ( \17290 , RIbe2b108_116);
not \U$17038 ( \17291 , \10936 );
or \U$17039 ( \17292 , \17290 , \17291 );
nand \U$17040 ( \17293 , \14511 , RIbe2b090_115);
nand \U$17041 ( \17294 , \17292 , \17293 );
and \U$17042 ( \17295 , \17294 , \9903 );
not \U$17043 ( \17296 , \17294 );
not \U$17044 ( \17297 , \13030 );
and \U$17045 ( \17298 , \17296 , \17297 );
nor \U$17046 ( \17299 , \17295 , \17298 );
and \U$17047 ( \17300 , \12765 , RIbe2a190_83);
and \U$17048 ( \17301 , \14491 , RIbe2a5c8_92);
nor \U$17049 ( \17302 , \17300 , \17301 );
and \U$17050 ( \17303 , \17302 , \12774 );
not \U$17051 ( \17304 , \17302 );
and \U$17052 ( \17305 , \17304 , \14000 );
nor \U$17053 ( \17306 , \17303 , \17305 );
and \U$17054 ( \17307 , \17299 , \17306 );
and \U$17055 ( \17308 , \12943 , RIbe2a280_85);
and \U$17056 ( \17309 , \15628 , RIbe2a208_84);
nor \U$17057 ( \17310 , \17308 , \17309 );
not \U$17058 ( \17311 , \17310 );
not \U$17059 ( \17312 , \12195 );
and \U$17060 ( \17313 , \17311 , \17312 );
and \U$17061 ( \17314 , \17310 , \12195 );
nor \U$17062 ( \17315 , \17313 , \17314 );
nor \U$17063 ( \17316 , \17307 , \17315 );
nor \U$17064 ( \17317 , \17299 , \17306 );
nor \U$17065 ( \17318 , \17316 , \17317 );
not \U$17066 ( \17319 , RIbe2a2f8_86);
not \U$17067 ( \17320 , \12787 );
or \U$17068 ( \17321 , \17319 , \17320 );
nand \U$17069 ( \17322 , \12890 , RIbe2acd0_107);
nand \U$17070 ( \17323 , \17321 , \17322 );
and \U$17071 ( \17324 , \17323 , \14103 );
not \U$17072 ( \17325 , \17323 );
and \U$17073 ( \17326 , \17325 , \12801 );
nor \U$17074 ( \17327 , \17324 , \17326 );
not \U$17075 ( \17328 , RIbe2a028_80);
not \U$17076 ( \17329 , \13003 );
or \U$17077 ( \17330 , \17328 , \17329 );
nand \U$17078 ( \17331 , RIbe29fb0_79, RIbe2ae38_110);
nand \U$17079 ( \17332 , \17330 , \17331 );
xor \U$17080 ( \17333 , \17332 , RIbe2aeb0_111);
not \U$17081 ( \17334 , \17333 );
nand \U$17082 ( \17335 , \17334 , \8957 );
and \U$17083 ( \17336 , \17327 , \17335 );
nor \U$17084 ( \17337 , \17334 , \14666 );
nor \U$17085 ( \17338 , \17336 , \17337 );
nand \U$17086 ( \17339 , \17318 , \17338 );
and \U$17087 ( \17340 , \17289 , \17339 );
nor \U$17088 ( \17341 , \17318 , \17338 );
nor \U$17089 ( \17342 , \17340 , \17341 );
nand \U$17090 ( \17343 , \17253 , \17342 );
not \U$17091 ( \17344 , \17343 );
xor \U$17092 ( \17345 , \17009 , \16990 );
and \U$17093 ( \17346 , \17345 , \16998 );
not \U$17094 ( \17347 , \17345 );
not \U$17095 ( \17348 , \16998 );
and \U$17096 ( \17349 , \17347 , \17348 );
nor \U$17097 ( \17350 , \17346 , \17349 );
not \U$17098 ( \17351 , \17350 );
xor \U$17099 ( \17352 , \17036 , \17027 );
xor \U$17100 ( \17353 , \17352 , \17046 );
or \U$17101 ( \17354 , \17351 , \17353 );
xor \U$17102 ( \17355 , \17080 , \17089 );
xor \U$17103 ( \17356 , \17355 , \17099 );
nand \U$17104 ( \17357 , \17354 , \17356 );
nand \U$17105 ( \17358 , \17351 , \17353 );
nand \U$17106 ( \17359 , \17357 , \17358 );
not \U$17107 ( \17360 , \17359 );
or \U$17108 ( \17361 , \17344 , \17360 );
not \U$17109 ( \17362 , \17342 );
nand \U$17110 ( \17363 , \17362 , \17252 );
nand \U$17111 ( \17364 , \17361 , \17363 );
xor \U$17112 ( \17365 , \17187 , \17364 );
xor \U$17113 ( \17366 , \17061 , \17063 );
xor \U$17114 ( \17367 , \17366 , \17066 );
not \U$17115 ( \17368 , \17050 );
not \U$17116 ( \17369 , \17012 );
or \U$17117 ( \17370 , \17368 , \17369 );
nand \U$17118 ( \17371 , \17013 , \17049 );
nand \U$17119 ( \17372 , \17370 , \17371 );
and \U$17120 ( \17373 , \17372 , \16980 );
not \U$17121 ( \17374 , \17372 );
and \U$17122 ( \17375 , \17374 , \16979 );
nor \U$17123 ( \17376 , \17373 , \17375 );
or \U$17124 ( \17377 , \17367 , \17376 );
xor \U$17125 ( \17378 , \17072 , \17102 );
xor \U$17126 ( \17379 , \17378 , \17105 );
nand \U$17127 ( \17380 , \17377 , \17379 );
nand \U$17128 ( \17381 , \17367 , \17376 );
nand \U$17129 ( \17382 , \17380 , \17381 );
and \U$17130 ( \17383 , \17365 , \17382 );
and \U$17131 ( \17384 , \17187 , \17364 );
or \U$17132 ( \17385 , \17383 , \17384 );
xor \U$17133 ( \17386 , \17180 , \17385 );
not \U$17134 ( \17387 , \14585 );
not \U$17135 ( \17388 , \14520 );
not \U$17136 ( \17389 , \14580 );
and \U$17137 ( \17390 , \17388 , \17389 );
and \U$17138 ( \17391 , \14520 , \14580 );
nor \U$17139 ( \17392 , \17390 , \17391 );
not \U$17140 ( \17393 , \17392 );
or \U$17141 ( \17394 , \17387 , \17393 );
or \U$17142 ( \17395 , \17392 , \14585 );
nand \U$17143 ( \17396 , \17394 , \17395 );
xor \U$17144 ( \17397 , \17129 , \17132 );
not \U$17145 ( \17398 , \17397 );
not \U$17146 ( \17399 , \17136 );
or \U$17147 ( \17400 , \17398 , \17399 );
or \U$17148 ( \17401 , \17136 , \17397 );
nand \U$17149 ( \17402 , \17400 , \17401 );
xor \U$17150 ( \17403 , \17396 , \17402 );
xor \U$17151 ( \17404 , \17052 , \17069 );
xor \U$17152 ( \17405 , \17404 , \17108 );
and \U$17153 ( \17406 , \17403 , \17405 );
and \U$17154 ( \17407 , \17396 , \17402 );
or \U$17155 ( \17408 , \17406 , \17407 );
and \U$17156 ( \17409 , \17386 , \17408 );
and \U$17157 ( \17410 , \17180 , \17385 );
or \U$17158 ( \17411 , \17409 , \17410 );
not \U$17159 ( \17412 , \17411 );
nand \U$17160 ( \17413 , \17178 , \17412 );
and \U$17161 ( \17414 , \17156 , \17413 );
and \U$17162 ( \17415 , \17411 , \17177 );
nor \U$17163 ( \17416 , \17414 , \17415 );
not \U$17164 ( \17417 , \17416 );
not \U$17165 ( \17418 , \17417 );
not \U$17166 ( \17419 , \14700 );
not \U$17167 ( \17420 , \14698 );
not \U$17168 ( \17421 , \17420 );
or \U$17169 ( \17422 , \17419 , \17421 );
not \U$17170 ( \17423 , \14700 );
nand \U$17171 ( \17424 , \17423 , \14698 );
nand \U$17172 ( \17425 , \17422 , \17424 );
not \U$17173 ( \17426 , \17151 );
not \U$17174 ( \17427 , \17145 );
or \U$17175 ( \17428 , \17426 , \17427 );
not \U$17176 ( \17429 , \16947 );
nand \U$17177 ( \17430 , \17428 , \17429 );
nand \U$17178 ( \17431 , \17152 , \17148 );
nand \U$17179 ( \17432 , \17430 , \17431 );
xor \U$17180 ( \17433 , \17425 , \17432 );
xor \U$17181 ( \17434 , \14684 , \14686 );
xor \U$17182 ( \17435 , \17434 , \14692 );
xor \U$17183 ( \17436 , \17433 , \17435 );
not \U$17184 ( \17437 , \17436 );
not \U$17185 ( \17438 , \17437 );
or \U$17186 ( \17439 , \17418 , \17438 );
nand \U$17187 ( \17440 , \17436 , \17416 );
nand \U$17188 ( \17441 , \17439 , \17440 );
xor \U$17189 ( \17442 , \17168 , \17112 );
xnor \U$17190 ( \17443 , \17442 , \17175 );
xor \U$17191 ( \17444 , \17180 , \17385 );
xor \U$17192 ( \17445 , \17444 , \17408 );
xor \U$17193 ( \17446 , \17443 , \17445 );
xor \U$17194 ( \17447 , \17187 , \17364 );
xor \U$17195 ( \17448 , \17447 , \17382 );
xor \U$17196 ( \17449 , \17376 , \17379 );
xnor \U$17197 ( \17450 , \17449 , \17367 );
xor \U$17198 ( \17451 , \16965 , \16958 );
xnor \U$17199 ( \17452 , \17451 , \16976 );
xor \U$17200 ( \17453 , \17197 , \17213 );
xnor \U$17201 ( \17454 , \17453 , \17248 );
xor \U$17202 ( \17455 , \17452 , \17454 );
and \U$17203 ( \17456 , \17356 , \17350 );
not \U$17204 ( \17457 , \17356 );
and \U$17205 ( \17458 , \17457 , \17351 );
or \U$17206 ( \17459 , \17456 , \17458 );
xnor \U$17207 ( \17460 , \17459 , \17353 );
and \U$17208 ( \17461 , \17455 , \17460 );
and \U$17209 ( \17462 , \17452 , \17454 );
or \U$17210 ( \17463 , \17461 , \17462 );
not \U$17211 ( \17464 , \17463 );
xor \U$17212 ( \17465 , \17212 , \17207 );
not \U$17213 ( \17466 , \17465 );
not \U$17214 ( \17467 , \17466 );
not \U$17215 ( \17468 , \17235 );
not \U$17216 ( \17469 , \17225 );
or \U$17217 ( \17470 , \17468 , \17469 );
nand \U$17218 ( \17471 , \17224 , \17234 );
nand \U$17219 ( \17472 , \17470 , \17471 );
and \U$17220 ( \17473 , \17472 , \17244 );
not \U$17221 ( \17474 , \17472 );
and \U$17222 ( \17475 , \17474 , \17245 );
nor \U$17223 ( \17476 , \17473 , \17475 );
not \U$17224 ( \17477 , \17476 );
or \U$17225 ( \17478 , \17467 , \17477 );
not \U$17226 ( \17479 , \13227 );
and \U$17227 ( \17480 , \7299 , RIbe2b630_127);
and \U$17228 ( \17481 , \10898 , RIbe2b018_114);
nor \U$17229 ( \17482 , \17480 , \17481 );
not \U$17230 ( \17483 , \17482 );
or \U$17231 ( \17484 , \17479 , \17483 );
or \U$17232 ( \17485 , \17482 , \13167 );
nand \U$17233 ( \17486 , \17484 , \17485 );
not \U$17234 ( \17487 , RIbe2ab68_104);
not \U$17235 ( \17488 , \6561 );
or \U$17236 ( \17489 , \17487 , \17488 );
nand \U$17237 ( \17490 , \6963 , RIbe2aaf0_103);
nand \U$17238 ( \17491 , \17489 , \17490 );
and \U$17239 ( \17492 , \17491 , \7293 );
not \U$17240 ( \17493 , \17491 );
and \U$17241 ( \17494 , \17493 , \6572 );
nor \U$17242 ( \17495 , \17492 , \17494 );
xor \U$17243 ( \17496 , \17486 , \17495 );
not \U$17244 ( \17497 , RIbe2afa0_113);
not \U$17245 ( \17498 , \10949 );
or \U$17246 ( \17499 , \17497 , \17498 );
nand \U$17247 ( \17500 , \10952 , RIbe2af28_112);
nand \U$17248 ( \17501 , \17499 , \17500 );
and \U$17249 ( \17502 , \17501 , \7988 );
not \U$17250 ( \17503 , \17501 );
and \U$17251 ( \17504 , \17503 , \7984 );
nor \U$17252 ( \17505 , \17502 , \17504 );
and \U$17253 ( \17506 , \17496 , \17505 );
and \U$17254 ( \17507 , \17486 , \17495 );
or \U$17255 ( \17508 , \17506 , \17507 );
nand \U$17256 ( \17509 , \17478 , \17508 );
not \U$17257 ( \17510 , \17476 );
nand \U$17258 ( \17511 , \17510 , \17465 );
nand \U$17259 ( \17512 , \17509 , \17511 );
not \U$17260 ( \17513 , RIbe2acd0_107);
not \U$17261 ( \17514 , \13004 );
or \U$17262 ( \17515 , \17513 , \17514 );
nand \U$17263 ( \17516 , RIbe2a028_80, RIbe2ae38_110);
nand \U$17264 ( \17517 , \17515 , \17516 );
xnor \U$17265 ( \17518 , \17517 , RIbe2aeb0_111);
not \U$17266 ( \17519 , \17518 );
not \U$17267 ( \17520 , RIbe2a370_87);
not \U$17268 ( \17521 , \13518 );
or \U$17269 ( \17522 , \17520 , \17521 );
nand \U$17270 ( \17523 , RIbe2a2f8_86, \12890 );
nand \U$17271 ( \17524 , \17522 , \17523 );
and \U$17272 ( \17525 , \17524 , \14103 );
not \U$17273 ( \17526 , \17524 );
and \U$17274 ( \17527 , \17526 , \12893 );
or \U$17275 ( \17528 , \17525 , \17527 );
not \U$17276 ( \17529 , \17528 );
or \U$17277 ( \17530 , \17519 , \17529 );
not \U$17278 ( \17531 , \12823 );
not \U$17279 ( \17532 , RIbe2b5b8_126);
not \U$17280 ( \17533 , \13590 );
or \U$17281 ( \17534 , \17532 , \17533 );
nand \U$17282 ( \17535 , \13012 , RIbe2a3e8_88);
nand \U$17283 ( \17536 , \17534 , \17535 );
not \U$17284 ( \17537 , \17536 );
or \U$17285 ( \17538 , \17531 , \17537 );
or \U$17286 ( \17539 , \17536 , \12863 );
nand \U$17287 ( \17540 , \17538 , \17539 );
nand \U$17288 ( \17541 , \17530 , \17540 );
not \U$17289 ( \17542 , \17528 );
not \U$17290 ( \17543 , \17518 );
nand \U$17291 ( \17544 , \17542 , \17543 );
nand \U$17292 ( \17545 , \17541 , \17544 );
and \U$17293 ( \17546 , \10916 , RIbe2b1f8_118);
buf \U$17294 ( \17547 , \13038 );
and \U$17295 ( \17548 , \17547 , RIbe2b180_117);
nor \U$17296 ( \17549 , \17546 , \17548 );
and \U$17297 ( \17550 , \17549 , \7970 );
not \U$17298 ( \17551 , \17549 );
and \U$17299 ( \17552 , \17551 , \10912 );
nor \U$17300 ( \17553 , \17550 , \17552 );
not \U$17301 ( \17554 , \17553 );
not \U$17302 ( \17555 , \12219 );
not \U$17303 ( \17556 , RIbe2b270_119);
not \U$17304 ( \17557 , \10936 );
or \U$17305 ( \17558 , \17556 , \17557 );
nand \U$17306 ( \17559 , \12971 , RIbe2b108_116);
nand \U$17307 ( \17560 , \17558 , \17559 );
not \U$17308 ( \17561 , \17560 );
and \U$17309 ( \17562 , \17555 , \17561 );
and \U$17310 ( \17563 , \17560 , \13030 );
nor \U$17311 ( \17564 , \17562 , \17563 );
not \U$17312 ( \17565 , \17564 );
or \U$17313 ( \17566 , \17554 , \17565 );
and \U$17314 ( \17567 , \12943 , RIbe2b090_115);
and \U$17315 ( \17568 , \13669 , RIbe2a280_85);
nor \U$17316 ( \17569 , \17567 , \17568 );
and \U$17317 ( \17570 , \17569 , \12956 );
not \U$17318 ( \17571 , \17569 );
and \U$17319 ( \17572 , \17571 , \12195 );
nor \U$17320 ( \17573 , \17570 , \17572 );
nand \U$17321 ( \17574 , \17566 , \17573 );
not \U$17322 ( \17575 , \17564 );
not \U$17323 ( \17576 , \17553 );
nand \U$17324 ( \17577 , \17575 , \17576 );
nand \U$17325 ( \17578 , \17574 , \17577 );
xor \U$17326 ( \17579 , \17545 , \17578 );
not \U$17327 ( \17580 , \12927 );
and \U$17328 ( \17581 , \17040 , RIbe2a208_84);
nor \U$17329 ( \17582 , \12753 , \14285 );
nor \U$17330 ( \17583 , \17581 , \17582 );
not \U$17331 ( \17584 , \17583 );
or \U$17332 ( \17585 , \17580 , \17584 );
or \U$17333 ( \17586 , \17583 , \12774 );
nand \U$17334 ( \17587 , \17585 , \17586 );
not \U$17335 ( \17588 , RIbe2a5c8_92);
not \U$17336 ( \17589 , \16383 );
or \U$17337 ( \17590 , \17588 , \17589 );
nand \U$17338 ( \17591 , \12711 , RIbe2a550_91);
nand \U$17339 ( \17592 , \17590 , \17591 );
and \U$17340 ( \17593 , \17592 , \13068 );
not \U$17341 ( \17594 , \17592 );
and \U$17342 ( \17595 , \17594 , \13583 );
nor \U$17343 ( \17596 , \17593 , \17595 );
xor \U$17344 ( \17597 , \17587 , \17596 );
not \U$17345 ( \17598 , RIbe2a988_100);
not \U$17346 ( \17599 , \12847 );
or \U$17347 ( \17600 , \17598 , \17599 );
nand \U$17348 ( \17601 , \14074 , RIbe2a910_99);
nand \U$17349 ( \17602 , \17600 , \17601 );
and \U$17350 ( \17603 , \17602 , \14077 );
not \U$17351 ( \17604 , \17602 );
and \U$17352 ( \17605 , \17604 , \12746 );
nor \U$17353 ( \17606 , \17603 , \17605 );
and \U$17354 ( \17607 , \17597 , \17606 );
and \U$17355 ( \17608 , \17587 , \17596 );
or \U$17356 ( \17609 , \17607 , \17608 );
and \U$17357 ( \17610 , \17579 , \17609 );
and \U$17358 ( \17611 , \17545 , \17578 );
or \U$17359 ( \17612 , \17610 , \17611 );
xor \U$17360 ( \17613 , \17512 , \17612 );
and \U$17361 ( \17614 , \17333 , \7948 );
not \U$17362 ( \17615 , \17333 );
and \U$17363 ( \17616 , \17615 , \7646 );
or \U$17364 ( \17617 , \17614 , \17616 );
not \U$17365 ( \17618 , \17617 );
not \U$17366 ( \17619 , \17327 );
or \U$17367 ( \17620 , \17618 , \17619 );
or \U$17368 ( \17621 , \17327 , \17617 );
nand \U$17369 ( \17622 , \17620 , \17621 );
xor \U$17370 ( \17623 , \17299 , \17315 );
xnor \U$17371 ( \17624 , \17623 , \17306 );
xor \U$17372 ( \17625 , \17622 , \17624 );
not \U$17373 ( \17626 , \17262 );
not \U$17374 ( \17627 , \17287 );
or \U$17375 ( \17628 , \17626 , \17627 );
nand \U$17376 ( \17629 , \17286 , \17263 );
nand \U$17377 ( \17630 , \17628 , \17629 );
and \U$17378 ( \17631 , \17630 , \17274 );
not \U$17379 ( \17632 , \17630 );
and \U$17380 ( \17633 , \17632 , \17273 );
nor \U$17381 ( \17634 , \17631 , \17633 );
and \U$17382 ( \17635 , \17625 , \17634 );
and \U$17383 ( \17636 , \17622 , \17624 );
or \U$17384 ( \17637 , \17635 , \17636 );
and \U$17385 ( \17638 , \17613 , \17637 );
and \U$17386 ( \17639 , \17512 , \17612 );
or \U$17387 ( \17640 , \17638 , \17639 );
nor \U$17388 ( \17641 , \17464 , \17640 );
or \U$17389 ( \17642 , \17450 , \17641 );
nand \U$17390 ( \17643 , \17464 , \17640 );
nand \U$17391 ( \17644 , \17642 , \17643 );
xor \U$17392 ( \17645 , \17448 , \17644 );
xor \U$17393 ( \17646 , \17396 , \17402 );
xor \U$17394 ( \17647 , \17646 , \17405 );
and \U$17395 ( \17648 , \17645 , \17647 );
and \U$17396 ( \17649 , \17448 , \17644 );
or \U$17397 ( \17650 , \17648 , \17649 );
and \U$17398 ( \17651 , \17446 , \17650 );
and \U$17399 ( \17652 , \17443 , \17445 );
or \U$17400 ( \17653 , \17651 , \17652 );
xor \U$17401 ( \17654 , \17411 , \17177 );
xor \U$17402 ( \17655 , \17654 , \17156 );
xor \U$17403 ( \17656 , \17653 , \17655 );
nand \U$17404 ( \17657 , \17441 , \17656 );
not \U$17405 ( \17658 , \17657 );
not \U$17406 ( \17659 , \17359 );
not \U$17407 ( \17660 , \17362 );
not \U$17408 ( \17661 , \17253 );
and \U$17409 ( \17662 , \17660 , \17661 );
and \U$17410 ( \17663 , \17253 , \17362 );
nor \U$17411 ( \17664 , \17662 , \17663 );
not \U$17412 ( \17665 , \17664 );
or \U$17413 ( \17666 , \17659 , \17665 );
or \U$17414 ( \17667 , \17664 , \17359 );
nand \U$17415 ( \17668 , \17666 , \17667 );
not \U$17416 ( \17669 , \17289 );
xnor \U$17417 ( \17670 , \17318 , \17338 );
not \U$17418 ( \17671 , \17670 );
or \U$17419 ( \17672 , \17669 , \17671 );
or \U$17420 ( \17673 , \17670 , \17289 );
nand \U$17421 ( \17674 , \17672 , \17673 );
not \U$17422 ( \17675 , \17543 );
not \U$17423 ( \17676 , \17528 );
or \U$17424 ( \17677 , \17675 , \17676 );
nand \U$17425 ( \17678 , \17542 , \17518 );
nand \U$17426 ( \17679 , \17677 , \17678 );
xnor \U$17427 ( \17680 , \17679 , \17540 );
not \U$17428 ( \17681 , \17680 );
xor \U$17429 ( \17682 , \17587 , \17596 );
xor \U$17430 ( \17683 , \17682 , \17606 );
nand \U$17431 ( \17684 , \17681 , \17683 );
not \U$17432 ( \17685 , \17684 );
not \U$17433 ( \17686 , \17685 );
not \U$17434 ( \17687 , RIbe2a2f8_86);
not \U$17435 ( \17688 , \13004 );
or \U$17436 ( \17689 , \17687 , \17688 );
nand \U$17437 ( \17690 , RIbe2acd0_107, RIbe2ae38_110);
nand \U$17438 ( \17691 , \17689 , \17690 );
xnor \U$17439 ( \17692 , \17691 , RIbe2aeb0_111);
xor \U$17440 ( \17693 , \6569 , \17692 );
not \U$17441 ( \17694 , RIbe2a3e8_88);
not \U$17442 ( \17695 , \12787 );
or \U$17443 ( \17696 , \17694 , \17695 );
nand \U$17444 ( \17697 , \12890 , RIbe2a370_87);
nand \U$17445 ( \17698 , \17696 , \17697 );
xor \U$17446 ( \17699 , \17698 , \12800 );
and \U$17447 ( \17700 , \17693 , \17699 );
and \U$17448 ( \17701 , \6569 , \17692 );
or \U$17449 ( \17702 , \17700 , \17701 );
not \U$17450 ( \17703 , RIbe2b180_117);
not \U$17451 ( \17704 , \10936 );
or \U$17452 ( \17705 , \17703 , \17704 );
nand \U$17453 ( \17706 , \12213 , RIbe2b270_119);
nand \U$17454 ( \17707 , \17705 , \17706 );
and \U$17455 ( \17708 , \17707 , \9903 );
not \U$17456 ( \17709 , \17707 );
and \U$17457 ( \17710 , \17709 , \14757 );
nor \U$17458 ( \17711 , \17708 , \17710 );
not \U$17459 ( \17712 , RIbe2a280_85);
not \U$17460 ( \17713 , \12921 );
or \U$17461 ( \17714 , \17712 , \17713 );
not \U$17462 ( \17715 , \12752 );
nand \U$17463 ( \17716 , \17715 , RIbe2a208_84);
nand \U$17464 ( \17717 , \17714 , \17716 );
not \U$17465 ( \17718 , \17717 );
not \U$17466 ( \17719 , \12924 );
and \U$17467 ( \17720 , \17718 , \17719 );
and \U$17468 ( \17721 , \17717 , \12924 );
nor \U$17469 ( \17722 , \17720 , \17721 );
and \U$17470 ( \17723 , \17711 , \17722 );
not \U$17471 ( \17724 , RIbe2b108_116);
not \U$17472 ( \17725 , \12942 );
or \U$17473 ( \17726 , \17724 , \17725 );
nand \U$17474 ( \17727 , \13669 , RIbe2b090_115);
nand \U$17475 ( \17728 , \17726 , \17727 );
and \U$17476 ( \17729 , \17728 , \12195 );
not \U$17477 ( \17730 , \17728 );
and \U$17478 ( \17731 , \17730 , \12957 );
nor \U$17479 ( \17732 , \17729 , \17731 );
not \U$17480 ( \17733 , \17732 );
nor \U$17481 ( \17734 , \17723 , \17733 );
nor \U$17482 ( \17735 , \17711 , \17722 );
nor \U$17483 ( \17736 , \17734 , \17735 );
xor \U$17484 ( \17737 , \17702 , \17736 );
not \U$17485 ( \17738 , \16382 );
not \U$17486 ( \17739 , \14285 );
and \U$17487 ( \17740 , \17738 , \17739 );
not \U$17488 ( \17741 , \12711 );
not \U$17489 ( \17742 , RIbe2a5c8_92);
nor \U$17490 ( \17743 , \17741 , \17742 );
nor \U$17491 ( \17744 , \17740 , \17743 );
and \U$17492 ( \17745 , \17744 , \12716 );
not \U$17493 ( \17746 , \17744 );
and \U$17494 ( \17747 , \17746 , \12723 );
nor \U$17495 ( \17748 , \17745 , \17747 );
not \U$17496 ( \17749 , \17748 );
not \U$17497 ( \17750 , RIbe2a550_91);
not \U$17498 ( \17751 , \12732 );
or \U$17499 ( \17752 , \17750 , \17751 );
nand \U$17500 ( \17753 , \13077 , RIbe2a988_100);
nand \U$17501 ( \17754 , \17752 , \17753 );
and \U$17502 ( \17755 , \17754 , \12746 );
not \U$17503 ( \17756 , \17754 );
and \U$17504 ( \17757 , \17756 , \13570 );
nor \U$17505 ( \17758 , \17755 , \17757 );
not \U$17506 ( \17759 , \17758 );
and \U$17507 ( \17760 , \17749 , \17759 );
and \U$17508 ( \17761 , \17748 , \17758 );
not \U$17509 ( \17762 , RIbe2a910_99);
not \U$17510 ( \17763 , \13010 );
or \U$17511 ( \17764 , \17762 , \17763 );
nand \U$17512 ( \17765 , \12835 , RIbe2b5b8_126);
nand \U$17513 ( \17766 , \17764 , \17765 );
and \U$17514 ( \17767 , \17766 , \13595 );
not \U$17515 ( \17768 , \17766 );
and \U$17516 ( \17769 , \17768 , \12863 );
nor \U$17517 ( \17770 , \17767 , \17769 );
not \U$17518 ( \17771 , \17770 );
nor \U$17519 ( \17772 , \17761 , \17771 );
nor \U$17520 ( \17773 , \17760 , \17772 );
and \U$17521 ( \17774 , \17737 , \17773 );
and \U$17522 ( \17775 , \17702 , \17736 );
or \U$17523 ( \17776 , \17774 , \17775 );
not \U$17524 ( \17777 , \17776 );
not \U$17525 ( \17778 , \17777 );
or \U$17526 ( \17779 , \17686 , \17778 );
nand \U$17527 ( \17780 , \17776 , \17684 );
and \U$17528 ( \17781 , \13036 , RIbe2af28_112);
and \U$17529 ( \17782 , \9914 , RIbe2b1f8_118);
nor \U$17530 ( \17783 , \17781 , \17782 );
and \U$17531 ( \17784 , \17783 , \8077 );
not \U$17532 ( \17785 , \17783 );
and \U$17533 ( \17786 , \17785 , \13649 );
nor \U$17534 ( \17787 , \17784 , \17786 );
not \U$17535 ( \17788 , \17787 );
not \U$17536 ( \17789 , \17788 );
not \U$17537 ( \17790 , RIbe2b018_114);
not \U$17538 ( \17791 , \10949 );
or \U$17539 ( \17792 , \17790 , \17791 );
nand \U$17540 ( \17793 , \8269 , RIbe2afa0_113);
nand \U$17541 ( \17794 , \17792 , \17793 );
and \U$17542 ( \17795 , \17794 , \7984 );
not \U$17543 ( \17796 , \17794 );
and \U$17544 ( \17797 , \17796 , \7985 );
nor \U$17545 ( \17798 , \17795 , \17797 );
not \U$17546 ( \17799 , \17798 );
or \U$17547 ( \17800 , \17789 , \17799 );
not \U$17548 ( \17801 , \10897 );
not \U$17549 ( \17802 , RIbe2b630_127);
not \U$17550 ( \17803 , \17802 );
and \U$17551 ( \17804 , \17801 , \17803 );
and \U$17552 ( \17805 , \6980 , RIbe2aaf0_103);
nor \U$17553 ( \17806 , \17804 , \17805 );
and \U$17554 ( \17807 , \17806 , \13353 );
not \U$17555 ( \17808 , \17806 );
and \U$17556 ( \17809 , \17808 , \6992 );
or \U$17557 ( \17810 , \17807 , \17809 );
nand \U$17558 ( \17811 , \17800 , \17810 );
not \U$17559 ( \17812 , \17798 );
nand \U$17560 ( \17813 , \17812 , \17787 );
nand \U$17561 ( \17814 , \17811 , \17813 );
xor \U$17562 ( \17815 , \17486 , \17495 );
xor \U$17563 ( \17816 , \17815 , \17505 );
xor \U$17564 ( \17817 , \17814 , \17816 );
and \U$17565 ( \17818 , \17573 , \17564 );
not \U$17566 ( \17819 , \17573 );
and \U$17567 ( \17820 , \17819 , \17575 );
or \U$17568 ( \17821 , \17818 , \17820 );
and \U$17569 ( \17822 , \17821 , \17576 );
not \U$17570 ( \17823 , \17821 );
and \U$17571 ( \17824 , \17823 , \17553 );
nor \U$17572 ( \17825 , \17822 , \17824 );
and \U$17573 ( \17826 , \17817 , \17825 );
and \U$17574 ( \17827 , \17814 , \17816 );
or \U$17575 ( \17828 , \17826 , \17827 );
nand \U$17576 ( \17829 , \17780 , \17828 );
nand \U$17577 ( \17830 , \17779 , \17829 );
xor \U$17578 ( \17831 , \17674 , \17830 );
not \U$17579 ( \17832 , \17508 );
not \U$17580 ( \17833 , \17832 );
not \U$17581 ( \17834 , \17465 );
not \U$17582 ( \17835 , \17476 );
or \U$17583 ( \17836 , \17834 , \17835 );
or \U$17584 ( \17837 , \17465 , \17476 );
nand \U$17585 ( \17838 , \17836 , \17837 );
not \U$17586 ( \17839 , \17838 );
or \U$17587 ( \17840 , \17833 , \17839 );
or \U$17588 ( \17841 , \17838 , \17832 );
nand \U$17589 ( \17842 , \17840 , \17841 );
xor \U$17590 ( \17843 , \17545 , \17578 );
xor \U$17591 ( \17844 , \17843 , \17609 );
xor \U$17592 ( \17845 , \17842 , \17844 );
xor \U$17593 ( \17846 , \17622 , \17624 );
xor \U$17594 ( \17847 , \17846 , \17634 );
and \U$17595 ( \17848 , \17845 , \17847 );
and \U$17596 ( \17849 , \17842 , \17844 );
or \U$17597 ( \17850 , \17848 , \17849 );
and \U$17598 ( \17851 , \17831 , \17850 );
and \U$17599 ( \17852 , \17674 , \17830 );
or \U$17600 ( \17853 , \17851 , \17852 );
xor \U$17601 ( \17854 , \17668 , \17853 );
xor \U$17602 ( \17855 , \17512 , \17612 );
xor \U$17603 ( \17856 , \17855 , \17637 );
not \U$17604 ( \17857 , \17856 );
xor \U$17605 ( \17858 , \17452 , \17454 );
xor \U$17606 ( \17859 , \17858 , \17460 );
nor \U$17607 ( \17860 , \17857 , \17859 );
and \U$17608 ( \17861 , \17854 , \17860 );
and \U$17609 ( \17862 , \17668 , \17853 );
or \U$17610 ( \17863 , \17861 , \17862 );
xor \U$17611 ( \17864 , \17448 , \17644 );
xor \U$17612 ( \17865 , \17864 , \17647 );
and \U$17613 ( \17866 , \17863 , \17865 );
xor \U$17614 ( \17867 , \17443 , \17445 );
xor \U$17615 ( \17868 , \17867 , \17650 );
and \U$17616 ( \17869 , \17866 , \17868 );
and \U$17617 ( \17870 , \17658 , \17869 );
and \U$17618 ( \17871 , \17653 , \17655 );
not \U$17619 ( \17872 , \17871 );
not \U$17620 ( \17873 , \17441 );
or \U$17621 ( \17874 , \17872 , \17873 );
nand \U$17622 ( \17875 , \17436 , \17417 );
nand \U$17623 ( \17876 , \17874 , \17875 );
nor \U$17624 ( \17877 , \17870 , \17876 );
not \U$17625 ( \17878 , \17859 );
not \U$17626 ( \17879 , \17856 );
and \U$17627 ( \17880 , \17878 , \17879 );
and \U$17628 ( \17881 , \17859 , \17856 );
nor \U$17629 ( \17882 , \17880 , \17881 );
not \U$17630 ( \17883 , \17882 );
not \U$17631 ( \17884 , \17883 );
xor \U$17632 ( \17885 , \17674 , \17830 );
xor \U$17633 ( \17886 , \17885 , \17850 );
not \U$17634 ( \17887 , \17886 );
or \U$17635 ( \17888 , \17884 , \17887 );
or \U$17636 ( \17889 , \17886 , \17883 );
not \U$17637 ( \17890 , \17771 );
not \U$17638 ( \17891 , \17758 );
not \U$17639 ( \17892 , \17891 );
or \U$17640 ( \17893 , \17890 , \17892 );
nand \U$17641 ( \17894 , \17758 , \17770 );
nand \U$17642 ( \17895 , \17893 , \17894 );
not \U$17643 ( \17896 , \17748 );
and \U$17644 ( \17897 , \17895 , \17896 );
not \U$17645 ( \17898 , \17895 );
and \U$17646 ( \17899 , \17898 , \17748 );
nor \U$17647 ( \17900 , \17897 , \17899 );
not \U$17648 ( \17901 , \17900 );
xor \U$17649 ( \17902 , \6569 , \17692 );
xor \U$17650 ( \17903 , \17902 , \17699 );
nor \U$17651 ( \17904 , \17901 , \17903 );
not \U$17652 ( \17905 , RIbe2aeb0_111);
not \U$17653 ( \17906 , RIbe2a370_87);
nor \U$17654 ( \17907 , \17906 , \12810 );
and \U$17655 ( \17908 , RIbe2a2f8_86, RIbe2ae38_110);
nor \U$17656 ( \17909 , \17907 , \17908 );
not \U$17657 ( \17910 , \17909 );
or \U$17658 ( \17911 , \17905 , \17910 );
or \U$17659 ( \17912 , \17909 , RIbe2aeb0_111);
nand \U$17660 ( \17913 , \17911 , \17912 );
not \U$17661 ( \17914 , \17913 );
not \U$17662 ( \17915 , RIbe2b5b8_126);
not \U$17663 ( \17916 , \12787 );
or \U$17664 ( \17917 , \17915 , \17916 );
nand \U$17665 ( \17918 , RIbe2a3e8_88, \12890 );
nand \U$17666 ( \17919 , \17917 , \17918 );
and \U$17667 ( \17920 , \17919 , \12893 );
not \U$17668 ( \17921 , \17919 );
and \U$17669 ( \17922 , \17921 , \16334 );
nor \U$17670 ( \17923 , \17920 , \17922 );
nand \U$17671 ( \17924 , \17914 , \17923 );
not \U$17672 ( \17925 , \12863 );
not \U$17673 ( \17926 , RIbe2a988_100);
not \U$17674 ( \17927 , \13010 );
or \U$17675 ( \17928 , \17926 , \17927 );
nand \U$17676 ( \17929 , \13012 , RIbe2a910_99);
nand \U$17677 ( \17930 , \17928 , \17929 );
not \U$17678 ( \17931 , \17930 );
or \U$17679 ( \17932 , \17925 , \17931 );
or \U$17680 ( \17933 , \17930 , \12823 );
nand \U$17681 ( \17934 , \17932 , \17933 );
and \U$17682 ( \17935 , \17924 , \17934 );
not \U$17683 ( \17936 , \17913 );
nor \U$17684 ( \17937 , \17936 , \17923 );
nor \U$17685 ( \17938 , \17935 , \17937 );
not \U$17686 ( \17939 , \17938 );
not \U$17687 ( \17940 , \17939 );
not \U$17688 ( \17941 , RIbe2b1f8_118);
not \U$17689 ( \17942 , \14751 );
or \U$17690 ( \17943 , \17941 , \17942 );
nand \U$17691 ( \17944 , \12971 , RIbe2b180_117);
nand \U$17692 ( \17945 , \17943 , \17944 );
and \U$17693 ( \17946 , \17945 , \10944 );
not \U$17694 ( \17947 , \17945 );
and \U$17695 ( \17948 , \17947 , \12218 );
nor \U$17696 ( \17949 , \17946 , \17948 );
not \U$17697 ( \17950 , \17949 );
and \U$17698 ( \17951 , \13036 , RIbe2afa0_113);
and \U$17699 ( \17952 , \13040 , RIbe2af28_112);
nor \U$17700 ( \17953 , \17951 , \17952 );
and \U$17701 ( \17954 , \17953 , \7970 );
not \U$17702 ( \17955 , \17953 );
and \U$17703 ( \17956 , \17955 , \8077 );
nor \U$17704 ( \17957 , \17954 , \17956 );
not \U$17705 ( \17958 , \17957 );
not \U$17706 ( \17959 , \17958 );
or \U$17707 ( \17960 , \17950 , \17959 );
not \U$17708 ( \17961 , \17949 );
not \U$17709 ( \17962 , \17961 );
not \U$17710 ( \17963 , \17957 );
or \U$17711 ( \17964 , \17962 , \17963 );
and \U$17712 ( \17965 , \12943 , RIbe2b270_119);
not \U$17713 ( \17966 , RIbe2b108_116);
nor \U$17714 ( \17967 , \17966 , \16033 );
nor \U$17715 ( \17968 , \17965 , \17967 );
and \U$17716 ( \17969 , \17968 , \12195 );
not \U$17717 ( \17970 , \17968 );
and \U$17718 ( \17971 , \17970 , \12960 );
nor \U$17719 ( \17972 , \17969 , \17971 );
not \U$17720 ( \17973 , \17972 );
nand \U$17721 ( \17974 , \17964 , \17973 );
nand \U$17722 ( \17975 , \17960 , \17974 );
not \U$17723 ( \17976 , \17975 );
or \U$17724 ( \17977 , \17940 , \17976 );
not \U$17725 ( \17978 , RIbe2a5c8_92);
not \U$17726 ( \17979 , \12732 );
or \U$17727 ( \17980 , \17978 , \17979 );
nand \U$17728 ( \17981 , \12735 , RIbe2a550_91);
nand \U$17729 ( \17982 , \17980 , \17981 );
and \U$17730 ( \17983 , \17982 , \12743 );
not \U$17731 ( \17984 , \17982 );
and \U$17732 ( \17985 , \17984 , \12742 );
nor \U$17733 ( \17986 , \17983 , \17985 );
not \U$17734 ( \17987 , RIbe2a208_84);
not \U$17735 ( \17988 , \12871 );
or \U$17736 ( \17989 , \17987 , \17988 );
nand \U$17737 ( \17990 , \13728 , RIbe2a190_83);
nand \U$17738 ( \17991 , \17989 , \17990 );
and \U$17739 ( \17992 , \17991 , \12716 );
not \U$17740 ( \17993 , \17991 );
and \U$17741 ( \17994 , \17993 , \12723 );
nor \U$17742 ( \17995 , \17992 , \17994 );
or \U$17743 ( \17996 , \17986 , \17995 );
not \U$17744 ( \17997 , \13087 );
not \U$17745 ( \17998 , RIbe2a280_85);
not \U$17746 ( \17999 , \17998 );
and \U$17747 ( \18000 , \17997 , \17999 );
and \U$17748 ( \18001 , \12765 , RIbe2b090_115);
nor \U$17749 ( \18002 , \18000 , \18001 );
and \U$17750 ( \18003 , \18002 , \12770 );
not \U$17751 ( \18004 , \18002 );
and \U$17752 ( \18005 , \18004 , \12927 );
nor \U$17753 ( \18006 , \18003 , \18005 );
and \U$17754 ( \18007 , \17996 , \18006 );
and \U$17755 ( \18008 , \17995 , \17986 );
nor \U$17756 ( \18009 , \18007 , \18008 );
not \U$17757 ( \18010 , \18009 );
not \U$17758 ( \18011 , \17975 );
nand \U$17759 ( \18012 , \18011 , \17938 );
nand \U$17760 ( \18013 , \18010 , \18012 );
nand \U$17761 ( \18014 , \17977 , \18013 );
xor \U$17762 ( \18015 , \17904 , \18014 );
nand \U$17763 ( \18016 , \7653 , RIbe2ab68_104);
and \U$17764 ( \18017 , \18016 , \6569 );
not \U$17765 ( \18018 , \18016 );
and \U$17766 ( \18019 , \18018 , \7293 );
nor \U$17767 ( \18020 , \18017 , \18019 );
not \U$17768 ( \18021 , \18020 );
not \U$17769 ( \18022 , \17788 );
not \U$17770 ( \18023 , \17812 );
or \U$17771 ( \18024 , \18022 , \18023 );
nand \U$17772 ( \18025 , \17798 , \17787 );
nand \U$17773 ( \18026 , \18024 , \18025 );
not \U$17774 ( \18027 , \17810 );
and \U$17775 ( \18028 , \18026 , \18027 );
not \U$17776 ( \18029 , \18026 );
and \U$17777 ( \18030 , \18029 , \17810 );
nor \U$17778 ( \18031 , \18028 , \18030 );
not \U$17779 ( \18032 , \18031 );
not \U$17780 ( \18033 , \18032 );
or \U$17781 ( \18034 , \18021 , \18033 );
not \U$17782 ( \18035 , \18020 );
nand \U$17783 ( \18036 , \18035 , \18031 );
not \U$17784 ( \18037 , \17711 );
and \U$17785 ( \18038 , \17722 , \17732 );
not \U$17786 ( \18039 , \17722 );
and \U$17787 ( \18040 , \18039 , \17733 );
or \U$17788 ( \18041 , \18038 , \18040 );
not \U$17789 ( \18042 , \18041 );
or \U$17790 ( \18043 , \18037 , \18042 );
or \U$17791 ( \18044 , \18041 , \17711 );
nand \U$17792 ( \18045 , \18043 , \18044 );
nand \U$17793 ( \18046 , \18036 , \18045 );
nand \U$17794 ( \18047 , \18034 , \18046 );
and \U$17795 ( \18048 , \18015 , \18047 );
and \U$17796 ( \18049 , \17904 , \18014 );
or \U$17797 ( \18050 , \18048 , \18049 );
not \U$17798 ( \18051 , \18050 );
not \U$17799 ( \18052 , \17681 );
not \U$17800 ( \18053 , \17683 );
not \U$17801 ( \18054 , \18053 );
or \U$17802 ( \18055 , \18052 , \18054 );
nand \U$17803 ( \18056 , \17683 , \17680 );
nand \U$17804 ( \18057 , \18055 , \18056 );
not \U$17805 ( \18058 , \18057 );
xor \U$17806 ( \18059 , \17702 , \17736 );
xor \U$17807 ( \18060 , \18059 , \17773 );
not \U$17808 ( \18061 , \18060 );
not \U$17809 ( \18062 , \18061 );
or \U$17810 ( \18063 , \18058 , \18062 );
xor \U$17811 ( \18064 , \17814 , \17816 );
xor \U$17812 ( \18065 , \18064 , \17825 );
not \U$17813 ( \18066 , \18057 );
nand \U$17814 ( \18067 , \18066 , \18060 );
nand \U$17815 ( \18068 , \18065 , \18067 );
nand \U$17816 ( \18069 , \18063 , \18068 );
not \U$17817 ( \18070 , \18069 );
or \U$17818 ( \18071 , \18051 , \18070 );
or \U$17819 ( \18072 , \18069 , \18050 );
xor \U$17820 ( \18073 , \17842 , \17844 );
xor \U$17821 ( \18074 , \18073 , \17847 );
nand \U$17822 ( \18075 , \18072 , \18074 );
nand \U$17823 ( \18076 , \18071 , \18075 );
nand \U$17824 ( \18077 , \17889 , \18076 );
nand \U$17825 ( \18078 , \17888 , \18077 );
xor \U$17826 ( \18079 , \17668 , \17853 );
xor \U$17827 ( \18080 , \18079 , \17860 );
xor \U$17828 ( \18081 , \17463 , \17640 );
xnor \U$17829 ( \18082 , \18081 , \17450 );
not \U$17830 ( \18083 , \18082 );
and \U$17831 ( \18084 , \18080 , \18083 );
not \U$17832 ( \18085 , \18080 );
and \U$17833 ( \18086 , \18085 , \18082 );
nor \U$17834 ( \18087 , \18084 , \18086 );
and \U$17835 ( \18088 , \18078 , \18087 );
not \U$17836 ( \18089 , \18088 );
not \U$17837 ( \18090 , \18080 );
nor \U$17838 ( \18091 , \18090 , \18082 );
not \U$17839 ( \18092 , \18091 );
xor \U$17840 ( \18093 , \17863 , \17865 );
not \U$17841 ( \18094 , \18093 );
not \U$17842 ( \18095 , \18094 );
or \U$17843 ( \18096 , \18092 , \18095 );
not \U$17844 ( \18097 , \18091 );
nand \U$17845 ( \18098 , \18097 , \18093 );
nand \U$17846 ( \18099 , \18096 , \18098 );
not \U$17847 ( \18100 , \18099 );
or \U$17848 ( \18101 , \18089 , \18100 );
nand \U$17849 ( \18102 , \18093 , \18091 );
nand \U$17850 ( \18103 , \18101 , \18102 );
xor \U$17851 ( \18104 , \17866 , \17868 );
nand \U$17852 ( \18105 , \17658 , \18103 , \18104 );
nand \U$17853 ( \18106 , \17877 , \18105 );
and \U$17854 ( \18107 , \14695 , \14701 );
not \U$17855 ( \18108 , \14695 );
and \U$17856 ( \18109 , \18108 , \14702 );
or \U$17857 ( \18110 , \18107 , \18109 );
not \U$17858 ( \18111 , \14707 );
and \U$17859 ( \18112 , \18110 , \18111 );
not \U$17860 ( \18113 , \18110 );
and \U$17861 ( \18114 , \18113 , \14707 );
nor \U$17862 ( \18115 , \18112 , \18114 );
not \U$17863 ( \18116 , \18115 );
not \U$17864 ( \18117 , \18116 );
xor \U$17865 ( \18118 , \17425 , \17432 );
and \U$17866 ( \18119 , \18118 , \17435 );
and \U$17867 ( \18120 , \17425 , \17432 );
or \U$17868 ( \18121 , \18119 , \18120 );
not \U$17869 ( \18122 , \18121 );
not \U$17870 ( \18123 , \18122 );
or \U$17871 ( \18124 , \18117 , \18123 );
nand \U$17872 ( \18125 , \18115 , \18121 );
nand \U$17873 ( \18126 , \18124 , \18125 );
buf \U$17874 ( \18127 , \18126 );
nand \U$17875 ( \18128 , \18106 , \18127 );
xor \U$17876 ( \18129 , \17904 , \18014 );
xor \U$17877 ( \18130 , \18129 , \18047 );
not \U$17878 ( \18131 , RIbe2a910_99);
not \U$17879 ( \18132 , \12887 );
or \U$17880 ( \18133 , \18131 , \18132 );
nand \U$17881 ( \18134 , \12890 , RIbe2b5b8_126);
nand \U$17882 ( \18135 , \18133 , \18134 );
xor \U$17883 ( \18136 , \12801 , \18135 );
not \U$17884 ( \18137 , \18136 );
not \U$17885 ( \18138 , RIbe2a3e8_88);
not \U$17886 ( \18139 , \12811 );
or \U$17887 ( \18140 , \18138 , \18139 );
nand \U$17888 ( \18141 , RIbe2a370_87, RIbe2ae38_110);
nand \U$17889 ( \18142 , \18140 , \18141 );
xor \U$17890 ( \18143 , RIbe2aeb0_111, \18142 );
nor \U$17891 ( \18144 , \18143 , \13167 );
not \U$17892 ( \18145 , \18144 );
and \U$17893 ( \18146 , \18137 , \18145 );
and \U$17894 ( \18147 , \13167 , \18143 );
nor \U$17895 ( \18148 , \18146 , \18147 );
not \U$17896 ( \18149 , \18148 );
not \U$17897 ( \18150 , \18149 );
not \U$17898 ( \18151 , RIbe2af28_112);
not \U$17899 ( \18152 , \10936 );
or \U$17900 ( \18153 , \18151 , \18152 );
nand \U$17901 ( \18154 , \12971 , RIbe2b1f8_118);
nand \U$17902 ( \18155 , \18153 , \18154 );
and \U$17903 ( \18156 , \18155 , \10940 );
not \U$17904 ( \18157 , \18155 );
and \U$17905 ( \18158 , \18157 , \9902 );
nor \U$17906 ( \18159 , \18156 , \18158 );
and \U$17907 ( \18160 , \13092 , RIbe2b108_116);
not \U$17908 ( \18161 , RIbe2b090_115);
nor \U$17909 ( \18162 , \18161 , \12752 );
nor \U$17910 ( \18163 , \18160 , \18162 );
and \U$17911 ( \18164 , \18163 , \12927 );
not \U$17912 ( \18165 , \18163 );
and \U$17913 ( \18166 , \18165 , \12770 );
nor \U$17914 ( \18167 , \18164 , \18166 );
nand \U$17915 ( \18168 , \18159 , \18167 );
not \U$17916 ( \18169 , \14397 );
not \U$17917 ( \18170 , \13109 );
and \U$17918 ( \18171 , \18169 , \18170 );
and \U$17919 ( \18172 , \12943 , RIbe2b180_117);
nor \U$17920 ( \18173 , \18171 , \18172 );
not \U$17921 ( \18174 , \18173 );
not \U$17922 ( \18175 , \12195 );
and \U$17923 ( \18176 , \18174 , \18175 );
and \U$17924 ( \18177 , \18173 , \12195 );
nor \U$17925 ( \18178 , \18176 , \18177 );
not \U$17926 ( \18179 , \18178 );
and \U$17927 ( \18180 , \18168 , \18179 );
nor \U$17928 ( \18181 , \18159 , \18167 );
nor \U$17929 ( \18182 , \18180 , \18181 );
not \U$17930 ( \18183 , \18182 );
not \U$17931 ( \18184 , \18183 );
or \U$17932 ( \18185 , \18150 , \18184 );
not \U$17933 ( \18186 , \18148 );
not \U$17934 ( \18187 , \18182 );
or \U$17935 ( \18188 , \18186 , \18187 );
not \U$17936 ( \18189 , RIbe2a550_91);
not \U$17937 ( \18190 , \13010 );
or \U$17938 ( \18191 , \18189 , \18190 );
not \U$17939 ( \18192 , \13552 );
nand \U$17940 ( \18193 , \18192 , \12834 );
nand \U$17941 ( \18194 , \18191 , \18193 );
and \U$17942 ( \18195 , \18194 , \14555 );
not \U$17943 ( \18196 , \18194 );
and \U$17944 ( \18197 , \18196 , \12863 );
nor \U$17945 ( \18198 , \18195 , \18197 );
not \U$17946 ( \18199 , RIbe2a190_83);
not \U$17947 ( \18200 , \13074 );
or \U$17948 ( \18201 , \18199 , \18200 );
not \U$17949 ( \18202 , \17742 );
nand \U$17950 ( \18203 , \18202 , \14074 );
nand \U$17951 ( \18204 , \18201 , \18203 );
and \U$17952 ( \18205 , \18204 , \12743 );
not \U$17953 ( \18206 , \18204 );
and \U$17954 ( \18207 , \18206 , \12742 );
nor \U$17955 ( \18208 , \18205 , \18207 );
xor \U$17956 ( \18209 , \18198 , \18208 );
not \U$17957 ( \18210 , RIbe2a280_85);
not \U$17958 ( \18211 , \14523 );
or \U$17959 ( \18212 , \18210 , \18211 );
nand \U$17960 ( \18213 , \13728 , RIbe2a208_84);
nand \U$17961 ( \18214 , \18212 , \18213 );
and \U$17962 ( \18215 , \18214 , \12879 );
not \U$17963 ( \18216 , \18214 );
and \U$17964 ( \18217 , \18216 , \12723 );
nor \U$17965 ( \18218 , \18215 , \18217 );
and \U$17966 ( \18219 , \18209 , \18218 );
and \U$17967 ( \18220 , \18198 , \18208 );
or \U$17968 ( \18221 , \18219 , \18220 );
nand \U$17969 ( \18222 , \18188 , \18221 );
nand \U$17970 ( \18223 , \18185 , \18222 );
not \U$17971 ( \18224 , \18223 );
not \U$17972 ( \18225 , RIbe2b630_127);
not \U$17973 ( \18226 , \10949 );
or \U$17974 ( \18227 , \18225 , \18226 );
nand \U$17975 ( \18228 , \10952 , RIbe2b018_114);
nand \U$17976 ( \18229 , \18227 , \18228 );
and \U$17977 ( \18230 , \18229 , \7988 );
not \U$17978 ( \18231 , \18229 );
and \U$17979 ( \18232 , \18231 , \7984 );
nor \U$17980 ( \18233 , \18230 , \18232 );
not \U$17981 ( \18234 , \18233 );
not \U$17982 ( \18235 , \14643 );
not \U$17983 ( \18236 , \13192 );
and \U$17984 ( \18237 , \18235 , \18236 );
and \U$17985 ( \18238 , \6980 , RIbe2ab68_104);
nor \U$17986 ( \18239 , \18237 , \18238 );
and \U$17987 ( \18240 , \18239 , \7661 );
not \U$17988 ( \18241 , \18239 );
and \U$17989 ( \18242 , \18241 , \13353 );
nor \U$17990 ( \18243 , \18240 , \18242 );
not \U$17991 ( \18244 , \18243 );
and \U$17992 ( \18245 , \18234 , \18244 );
not \U$17993 ( \18246 , RIbe2aaf0_103);
not \U$17994 ( \18247 , \10949 );
or \U$17995 ( \18248 , \18246 , \18247 );
nand \U$17996 ( \18249 , \7981 , RIbe2b630_127);
nand \U$17997 ( \18250 , \18248 , \18249 );
and \U$17998 ( \18251 , \18250 , \6948 );
not \U$17999 ( \18252 , \18250 );
and \U$18000 ( \18253 , \18252 , \6950 );
or \U$18001 ( \18254 , \18251 , \18253 );
not \U$18002 ( \18255 , \18254 );
nand \U$18003 ( \18256 , \12251 , RIbe2ab68_104);
and \U$18004 ( \18257 , \18256 , \6992 );
not \U$18005 ( \18258 , \18256 );
and \U$18006 ( \18259 , \18258 , \6993 );
nor \U$18007 ( \18260 , \18257 , \18259 );
not \U$18008 ( \18261 , \18260 );
nand \U$18009 ( \18262 , \18255 , \18261 );
and \U$18010 ( \18263 , \13478 , RIbe2b018_114);
and \U$18011 ( \18264 , \13040 , RIbe2afa0_113);
nor \U$18012 ( \18265 , \18263 , \18264 );
and \U$18013 ( \18266 , \18265 , \8077 );
not \U$18014 ( \18267 , \18265 );
and \U$18015 ( \18268 , \18267 , \13649 );
nor \U$18016 ( \18269 , \18266 , \18268 );
and \U$18017 ( \18270 , \18262 , \18269 );
nor \U$18018 ( \18271 , \18255 , \18261 );
nor \U$18019 ( \18272 , \18270 , \18271 );
nor \U$18020 ( \18273 , \18245 , \18272 );
and \U$18021 ( \18274 , \18243 , \18233 );
nor \U$18022 ( \18275 , \18273 , \18274 );
not \U$18023 ( \18276 , \18275 );
and \U$18024 ( \18277 , \18224 , \18276 );
and \U$18025 ( \18278 , \18223 , \18275 );
nor \U$18026 ( \18279 , \18277 , \18278 );
xor \U$18027 ( \18280 , \17995 , \17986 );
xor \U$18028 ( \18281 , \18280 , \18006 );
not \U$18029 ( \18282 , \18281 );
not \U$18030 ( \18283 , \17934 );
xor \U$18031 ( \18284 , \17913 , \17923 );
not \U$18032 ( \18285 , \18284 );
or \U$18033 ( \18286 , \18283 , \18285 );
or \U$18034 ( \18287 , \18284 , \17934 );
nand \U$18035 ( \18288 , \18286 , \18287 );
not \U$18036 ( \18289 , \18288 );
or \U$18037 ( \18290 , \18282 , \18289 );
or \U$18038 ( \18291 , \18288 , \18281 );
not \U$18039 ( \18292 , \17961 );
not \U$18040 ( \18293 , \17973 );
or \U$18041 ( \18294 , \18292 , \18293 );
nand \U$18042 ( \18295 , \17972 , \17949 );
nand \U$18043 ( \18296 , \18294 , \18295 );
and \U$18044 ( \18297 , \18296 , \17958 );
not \U$18045 ( \18298 , \18296 );
and \U$18046 ( \18299 , \18298 , \17957 );
nor \U$18047 ( \18300 , \18297 , \18299 );
nand \U$18048 ( \18301 , \18291 , \18300 );
nand \U$18049 ( \18302 , \18290 , \18301 );
xnor \U$18050 ( \18303 , \18279 , \18302 );
not \U$18051 ( \18304 , \8077 );
not \U$18052 ( \18305 , RIbe2b630_127);
not \U$18053 ( \18306 , \9909 );
or \U$18054 ( \18307 , \18305 , \18306 );
nand \U$18055 ( \18308 , \17547 , RIbe2b018_114);
nand \U$18056 ( \18309 , \18307 , \18308 );
not \U$18057 ( \18310 , \18309 );
or \U$18058 ( \18311 , \18304 , \18310 );
or \U$18059 ( \18312 , \18309 , \16059 );
nand \U$18060 ( \18313 , \18311 , \18312 );
not \U$18061 ( \18314 , \18313 );
not \U$18062 ( \18315 , RIbe2afa0_113);
not \U$18063 ( \18316 , \10936 );
or \U$18064 ( \18317 , \18315 , \18316 );
nand \U$18065 ( \18318 , \14511 , RIbe2af28_112);
nand \U$18066 ( \18319 , \18317 , \18318 );
and \U$18067 ( \18320 , \18319 , \17297 );
not \U$18068 ( \18321 , \18319 );
and \U$18069 ( \18322 , \18321 , \14756 );
nor \U$18070 ( \18323 , \18320 , \18322 );
not \U$18071 ( \18324 , \18323 );
or \U$18072 ( \18325 , \18314 , \18324 );
or \U$18073 ( \18326 , \18313 , \18323 );
not \U$18074 ( \18327 , RIbe2b1f8_118);
not \U$18075 ( \18328 , \13049 );
or \U$18076 ( \18329 , \18327 , \18328 );
nand \U$18077 ( \18330 , \12948 , RIbe2b180_117);
nand \U$18078 ( \18331 , \18329 , \18330 );
and \U$18079 ( \18332 , \18331 , \12195 );
not \U$18080 ( \18333 , \18331 );
and \U$18081 ( \18334 , \18333 , \12960 );
nor \U$18082 ( \18335 , \18332 , \18334 );
nand \U$18083 ( \18336 , \18326 , \18335 );
nand \U$18084 ( \18337 , \18325 , \18336 );
not \U$18085 ( \18338 , RIbe2b5b8_126);
not \U$18086 ( \18339 , \13004 );
or \U$18087 ( \18340 , \18338 , \18339 );
nand \U$18088 ( \18341 , RIbe2a3e8_88, RIbe2ae38_110);
nand \U$18089 ( \18342 , \18340 , \18341 );
xnor \U$18090 ( \18343 , \18342 , RIbe2aeb0_111);
not \U$18091 ( \18344 , \18343 );
not \U$18092 ( \18345 , \18344 );
not \U$18093 ( \18346 , RIbe2a988_100);
not \U$18094 ( \18347 , \15249 );
or \U$18095 ( \18348 , \18346 , \18347 );
nand \U$18096 ( \18349 , \12794 , RIbe2a910_99);
nand \U$18097 ( \18350 , \18348 , \18349 );
and \U$18098 ( \18351 , \18350 , \16334 );
not \U$18099 ( \18352 , \18350 );
and \U$18100 ( \18353 , \18352 , \12801 );
nor \U$18101 ( \18354 , \18351 , \18353 );
not \U$18102 ( \18355 , \18354 );
or \U$18103 ( \18356 , \18345 , \18355 );
not \U$18104 ( \18357 , RIbe2a5c8_92);
not \U$18105 ( \18358 , \12831 );
or \U$18106 ( \18359 , \18357 , \18358 );
nand \U$18107 ( \18360 , \13012 , RIbe2a550_91);
nand \U$18108 ( \18361 , \18359 , \18360 );
and \U$18109 ( \18362 , \18361 , \12823 );
not \U$18110 ( \18363 , \18361 );
not \U$18111 ( \18364 , \14558 );
and \U$18112 ( \18365 , \18363 , \18364 );
nor \U$18113 ( \18366 , \18362 , \18365 );
not \U$18114 ( \18367 , \18366 );
not \U$18115 ( \18368 , \18354 );
nand \U$18116 ( \18369 , \18368 , \18343 );
nand \U$18117 ( \18370 , \18367 , \18369 );
nand \U$18118 ( \18371 , \18356 , \18370 );
nand \U$18119 ( \18372 , \18337 , \18371 );
or \U$18120 ( \18373 , \18337 , \18371 );
not \U$18121 ( \18374 , RIbe2b090_115);
not \U$18122 ( \18375 , \16383 );
or \U$18123 ( \18376 , \18374 , \18375 );
nand \U$18124 ( \18377 , \13728 , RIbe2a280_85);
nand \U$18125 ( \18378 , \18376 , \18377 );
and \U$18126 ( \18379 , \18378 , \12723 );
not \U$18127 ( \18380 , \18378 );
and \U$18128 ( \18381 , \18380 , \12879 );
nor \U$18129 ( \18382 , \18379 , \18381 );
not \U$18130 ( \18383 , RIbe2a208_84);
not \U$18131 ( \18384 , \12847 );
or \U$18132 ( \18385 , \18383 , \18384 );
nand \U$18133 ( \18386 , \13077 , RIbe2a190_83);
nand \U$18134 ( \18387 , \18385 , \18386 );
and \U$18135 ( \18388 , \18387 , \12746 );
not \U$18136 ( \18389 , \18387 );
and \U$18137 ( \18390 , \18389 , \12743 );
nor \U$18138 ( \18391 , \18388 , \18390 );
and \U$18139 ( \18392 , \18382 , \18391 );
not \U$18140 ( \18393 , RIbe2b270_119);
not \U$18141 ( \18394 , \17040 );
or \U$18142 ( \18395 , \18393 , \18394 );
not \U$18143 ( \18396 , \12753 );
nand \U$18144 ( \18397 , \18396 , RIbe2b108_116);
nand \U$18145 ( \18398 , \18395 , \18397 );
not \U$18146 ( \18399 , \18398 );
not \U$18147 ( \18400 , \12924 );
and \U$18148 ( \18401 , \18399 , \18400 );
and \U$18149 ( \18402 , \18398 , \12769 );
nor \U$18150 ( \18403 , \18401 , \18402 );
nor \U$18151 ( \18404 , \18392 , \18403 );
nor \U$18152 ( \18405 , \18382 , \18391 );
nor \U$18153 ( \18406 , \18404 , \18405 );
not \U$18154 ( \18407 , \18406 );
nand \U$18155 ( \18408 , \18373 , \18407 );
nand \U$18156 ( \18409 , \18372 , \18408 );
xor \U$18157 ( \18410 , \18198 , \18208 );
xor \U$18158 ( \18411 , \18410 , \18218 );
xor \U$18159 ( \18412 , \18260 , \18254 );
xor \U$18160 ( \18413 , \18412 , \18269 );
xor \U$18161 ( \18414 , \18411 , \18413 );
not \U$18162 ( \18415 , \18167 );
not \U$18163 ( \18416 , \18179 );
or \U$18164 ( \18417 , \18415 , \18416 );
not \U$18165 ( \18418 , \18167 );
nand \U$18166 ( \18419 , \18418 , \18178 );
nand \U$18167 ( \18420 , \18417 , \18419 );
xnor \U$18168 ( \18421 , \18420 , \18159 );
and \U$18169 ( \18422 , \18414 , \18421 );
and \U$18170 ( \18423 , \18411 , \18413 );
or \U$18171 ( \18424 , \18422 , \18423 );
xor \U$18172 ( \18425 , \18409 , \18424 );
xor \U$18173 ( \18426 , \18281 , \18300 );
and \U$18174 ( \18427 , \18426 , \18288 );
not \U$18175 ( \18428 , \18426 );
not \U$18176 ( \18429 , \18288 );
and \U$18177 ( \18430 , \18428 , \18429 );
nor \U$18178 ( \18431 , \18427 , \18430 );
and \U$18179 ( \18432 , \18425 , \18431 );
and \U$18180 ( \18433 , \18409 , \18424 );
or \U$18181 ( \18434 , \18432 , \18433 );
xor \U$18182 ( \18435 , \18303 , \18434 );
not \U$18183 ( \18436 , \17903 );
not \U$18184 ( \18437 , \18436 );
not \U$18185 ( \18438 , \17901 );
or \U$18186 ( \18439 , \18437 , \18438 );
nand \U$18187 ( \18440 , \17900 , \17903 );
nand \U$18188 ( \18441 , \18439 , \18440 );
xor \U$18189 ( \18442 , \18020 , \17711 );
xnor \U$18190 ( \18443 , \18442 , \18041 );
and \U$18191 ( \18444 , \18443 , \18031 );
not \U$18192 ( \18445 , \18443 );
and \U$18193 ( \18446 , \18445 , \18032 );
nor \U$18194 ( \18447 , \18444 , \18446 );
xor \U$18195 ( \18448 , \18441 , \18447 );
xnor \U$18196 ( \18449 , \17975 , \18009 );
and \U$18197 ( \18450 , \18449 , \17938 );
not \U$18198 ( \18451 , \18449 );
and \U$18199 ( \18452 , \18451 , \17939 );
nor \U$18200 ( \18453 , \18450 , \18452 );
xor \U$18201 ( \18454 , \18448 , \18453 );
and \U$18202 ( \18455 , \18435 , \18454 );
and \U$18203 ( \18456 , \18303 , \18434 );
or \U$18204 ( \18457 , \18455 , \18456 );
xor \U$18205 ( \18458 , \18130 , \18457 );
xor \U$18206 ( \18459 , \18057 , \18061 );
xor \U$18207 ( \18460 , \18459 , \18065 );
not \U$18208 ( \18461 , \18460 );
not \U$18209 ( \18462 , \18441 );
not \U$18210 ( \18463 , \18453 );
not \U$18211 ( \18464 , \18463 );
or \U$18212 ( \18465 , \18462 , \18464 );
not \U$18213 ( \18466 , \18447 );
not \U$18214 ( \18467 , \18441 );
nand \U$18215 ( \18468 , \18467 , \18453 );
nand \U$18216 ( \18469 , \18466 , \18468 );
nand \U$18217 ( \18470 , \18465 , \18469 );
not \U$18218 ( \18471 , \18470 );
not \U$18219 ( \18472 , \18275 );
not \U$18220 ( \18473 , \18223 );
not \U$18221 ( \18474 , \18473 );
or \U$18222 ( \18475 , \18472 , \18474 );
nand \U$18223 ( \18476 , \18475 , \18302 );
not \U$18224 ( \18477 , \18275 );
nand \U$18225 ( \18478 , \18477 , \18223 );
and \U$18226 ( \18479 , \18476 , \18478 );
not \U$18227 ( \18480 , \18479 );
and \U$18228 ( \18481 , \18471 , \18480 );
and \U$18229 ( \18482 , \18470 , \18479 );
nor \U$18230 ( \18483 , \18481 , \18482 );
not \U$18231 ( \18484 , \18483 );
or \U$18232 ( \18485 , \18461 , \18484 );
or \U$18233 ( \18486 , \18483 , \18460 );
nand \U$18234 ( \18487 , \18485 , \18486 );
and \U$18235 ( \18488 , \18458 , \18487 );
and \U$18236 ( \18489 , \18130 , \18457 );
or \U$18237 ( \18490 , \18488 , \18489 );
not \U$18238 ( \18491 , \18490 );
not \U$18239 ( \18492 , \18491 );
not \U$18240 ( \18493 , \17685 );
not \U$18241 ( \18494 , \17777 );
or \U$18242 ( \18495 , \18493 , \18494 );
or \U$18243 ( \18496 , \17777 , \17685 );
nand \U$18244 ( \18497 , \18495 , \18496 );
xor \U$18245 ( \18498 , \17828 , \18497 );
xor \U$18246 ( \18499 , \18050 , \18069 );
xnor \U$18247 ( \18500 , \18499 , \18074 );
xor \U$18248 ( \18501 , \18498 , \18500 );
not \U$18249 ( \18502 , \18470 );
nand \U$18250 ( \18503 , \18502 , \18479 );
and \U$18251 ( \18504 , \18460 , \18503 );
not \U$18252 ( \18505 , \18479 );
and \U$18253 ( \18506 , \18470 , \18505 );
nor \U$18254 ( \18507 , \18504 , \18506 );
xor \U$18255 ( \18508 , \18501 , \18507 );
not \U$18256 ( \18509 , \18508 );
not \U$18257 ( \18510 , \18509 );
or \U$18258 ( \18511 , \18492 , \18510 );
nand \U$18259 ( \18512 , \18508 , \18490 );
nand \U$18260 ( \18513 , \18511 , \18512 );
xor \U$18261 ( \18514 , \18498 , \18500 );
and \U$18262 ( \18515 , \18514 , \18507 );
and \U$18263 ( \18516 , \18498 , \18500 );
or \U$18264 ( \18517 , \18515 , \18516 );
xor \U$18265 ( \18518 , \17882 , \17886 );
xor \U$18266 ( \18519 , \18518 , \18076 );
xor \U$18267 ( \18520 , \18517 , \18519 );
not \U$18268 ( \18521 , \18272 );
xor \U$18269 ( \18522 , \18243 , \18233 );
not \U$18270 ( \18523 , \18522 );
or \U$18271 ( \18524 , \18521 , \18523 );
or \U$18272 ( \18525 , \18522 , \18272 );
nand \U$18273 ( \18526 , \18524 , \18525 );
xor \U$18274 ( \18527 , \18411 , \18413 );
xor \U$18275 ( \18528 , \18527 , \18421 );
not \U$18276 ( \18529 , \18337 );
not \U$18277 ( \18530 , \18529 );
not \U$18278 ( \18531 , \18407 );
or \U$18279 ( \18532 , \18530 , \18531 );
nand \U$18280 ( \18533 , \18406 , \18337 );
nand \U$18281 ( \18534 , \18532 , \18533 );
xnor \U$18282 ( \18535 , \18534 , \18371 );
not \U$18283 ( \18536 , \18535 );
and \U$18284 ( \18537 , \18528 , \18536 );
xor \U$18285 ( \18538 , \18526 , \18537 );
xor \U$18286 ( \18539 , \13167 , \18143 );
not \U$18287 ( \18540 , \18539 );
not \U$18288 ( \18541 , \18136 );
or \U$18289 ( \18542 , \18540 , \18541 );
or \U$18290 ( \18543 , \18136 , \18539 );
nand \U$18291 ( \18544 , \18542 , \18543 );
not \U$18292 ( \18545 , \18544 );
not \U$18293 ( \18546 , RIbe2a550_91);
not \U$18294 ( \18547 , \13518 );
or \U$18295 ( \18548 , \18546 , \18547 );
nand \U$18296 ( \18549 , \12890 , RIbe2a988_100);
nand \U$18297 ( \18550 , \18548 , \18549 );
and \U$18298 ( \18551 , \18550 , \12804 );
not \U$18299 ( \18552 , \18550 );
and \U$18300 ( \18553 , \18552 , \12893 );
nor \U$18301 ( \18554 , \18551 , \18553 );
not \U$18302 ( \18555 , \18554 );
not \U$18303 ( \18556 , RIbe2a910_99);
not \U$18304 ( \18557 , \13004 );
or \U$18305 ( \18558 , \18556 , \18557 );
nand \U$18306 ( \18559 , RIbe2b5b8_126, RIbe2ae38_110);
nand \U$18307 ( \18560 , \18558 , \18559 );
xnor \U$18308 ( \18561 , \18560 , RIbe2aeb0_111);
nand \U$18309 ( \18562 , \18561 , \7984 );
not \U$18310 ( \18563 , \18562 );
or \U$18311 ( \18564 , \18555 , \18563 );
not \U$18312 ( \18565 , \18561 );
nand \U$18313 ( \18566 , \18565 , \8480 );
nand \U$18314 ( \18567 , \18564 , \18566 );
not \U$18315 ( \18568 , \18567 );
not \U$18316 ( \18569 , RIbe2b018_114);
not \U$18317 ( \18570 , \10936 );
or \U$18318 ( \18571 , \18569 , \18570 );
nand \U$18319 ( \18572 , \14511 , RIbe2afa0_113);
nand \U$18320 ( \18573 , \18571 , \18572 );
not \U$18321 ( \18574 , \18573 );
not \U$18322 ( \18575 , \14756 );
and \U$18323 ( \18576 , \18574 , \18575 );
and \U$18324 ( \18577 , \18573 , \12219 );
nor \U$18325 ( \18578 , \18576 , \18577 );
not \U$18326 ( \18579 , \12753 );
not \U$18327 ( \18580 , \13109 );
and \U$18328 ( \18581 , \18579 , \18580 );
and \U$18329 ( \18582 , \13738 , RIbe2b180_117);
nor \U$18330 ( \18583 , \18581 , \18582 );
and \U$18331 ( \18584 , \18583 , \12927 );
not \U$18332 ( \18585 , \18583 );
and \U$18333 ( \18586 , \18585 , \12924 );
nor \U$18334 ( \18587 , \18584 , \18586 );
and \U$18335 ( \18588 , \18578 , \18587 );
not \U$18336 ( \18589 , RIbe2af28_112);
not \U$18337 ( \18590 , \15205 );
or \U$18338 ( \18591 , \18589 , \18590 );
nand \U$18339 ( \18592 , \12948 , RIbe2b1f8_118);
nand \U$18340 ( \18593 , \18591 , \18592 );
not \U$18341 ( \18594 , \18593 );
not \U$18342 ( \18595 , \12957 );
and \U$18343 ( \18596 , \18594 , \18595 );
and \U$18344 ( \18597 , \18593 , \12956 );
nor \U$18345 ( \18598 , \18596 , \18597 );
nor \U$18346 ( \18599 , \18588 , \18598 );
nor \U$18347 ( \18600 , \18578 , \18587 );
nor \U$18348 ( \18601 , \18599 , \18600 );
not \U$18349 ( \18602 , \18601 );
not \U$18350 ( \18603 , \18602 );
or \U$18351 ( \18604 , \18568 , \18603 );
or \U$18352 ( \18605 , \18602 , \18567 );
not \U$18353 ( \18606 , RIbe2a190_83);
buf \U$18354 ( \18607 , \12830 );
not \U$18355 ( \18608 , \18607 );
not \U$18356 ( \18609 , \18608 );
or \U$18357 ( \18610 , \18606 , \18609 );
nand \U$18358 ( \18611 , \12835 , RIbe2a5c8_92);
nand \U$18359 ( \18612 , \18610 , \18611 );
and \U$18360 ( \18613 , \18612 , \18364 );
not \U$18361 ( \18614 , \18612 );
and \U$18362 ( \18615 , \18614 , \15263 );
nor \U$18363 ( \18616 , \18613 , \18615 );
not \U$18364 ( \18617 , \18616 );
not \U$18365 ( \18618 , \13583 );
not \U$18366 ( \18619 , RIbe2b108_116);
not \U$18367 ( \18620 , \15573 );
or \U$18368 ( \18621 , \18619 , \18620 );
nand \U$18369 ( \18622 , \12711 , RIbe2b090_115);
nand \U$18370 ( \18623 , \18621 , \18622 );
not \U$18371 ( \18624 , \18623 );
or \U$18372 ( \18625 , \18618 , \18624 );
or \U$18373 ( \18626 , \18623 , \13583 );
nand \U$18374 ( \18627 , \18625 , \18626 );
not \U$18375 ( \18628 , \18627 );
or \U$18376 ( \18629 , \18617 , \18628 );
or \U$18377 ( \18630 , \18627 , \18616 );
not \U$18378 ( \18631 , \12742 );
not \U$18379 ( \18632 , RIbe2a280_85);
not \U$18380 ( \18633 , \14071 );
or \U$18381 ( \18634 , \18632 , \18633 );
nand \U$18382 ( \18635 , \14074 , RIbe2a208_84);
nand \U$18383 ( \18636 , \18634 , \18635 );
not \U$18384 ( \18637 , \18636 );
or \U$18385 ( \18638 , \18631 , \18637 );
or \U$18386 ( \18639 , \18636 , \12742 );
nand \U$18387 ( \18640 , \18638 , \18639 );
nand \U$18388 ( \18641 , \18630 , \18640 );
nand \U$18389 ( \18642 , \18629 , \18641 );
nand \U$18390 ( \18643 , \18605 , \18642 );
nand \U$18391 ( \18644 , \18604 , \18643 );
not \U$18392 ( \18645 , \18644 );
or \U$18393 ( \18646 , \18545 , \18645 );
or \U$18394 ( \18647 , \18644 , \18544 );
xor \U$18395 ( \18648 , \18382 , \18391 );
xnor \U$18396 ( \18649 , \18648 , \18403 );
and \U$18397 ( \18650 , \10949 , RIbe2ab68_104);
and \U$18398 ( \18651 , \10952 , RIbe2aaf0_103);
nor \U$18399 ( \18652 , \18650 , \18651 );
and \U$18400 ( \18653 , \18652 , \8480 );
not \U$18401 ( \18654 , \18652 );
and \U$18402 ( \18655 , \18654 , \6949 );
nor \U$18403 ( \18656 , \18653 , \18655 );
not \U$18404 ( \18657 , \18656 );
or \U$18405 ( \18658 , \18649 , \18657 );
not \U$18406 ( \18659 , \18313 );
xor \U$18407 ( \18660 , \18335 , \18323 );
not \U$18408 ( \18661 , \18660 );
not \U$18409 ( \18662 , \18661 );
or \U$18410 ( \18663 , \18659 , \18662 );
not \U$18411 ( \18664 , \18313 );
nand \U$18412 ( \18665 , \18664 , \18660 );
nand \U$18413 ( \18666 , \18663 , \18665 );
nand \U$18414 ( \18667 , \18658 , \18666 );
nand \U$18415 ( \18668 , \18649 , \18657 );
nand \U$18416 ( \18669 , \18667 , \18668 );
nand \U$18417 ( \18670 , \18647 , \18669 );
nand \U$18418 ( \18671 , \18646 , \18670 );
and \U$18419 ( \18672 , \18538 , \18671 );
and \U$18420 ( \18673 , \18526 , \18537 );
or \U$18421 ( \18674 , \18672 , \18673 );
or \U$18422 ( \18675 , \18183 , \18148 );
or \U$18423 ( \18676 , \18182 , \18149 );
nand \U$18424 ( \18677 , \18675 , \18676 );
xor \U$18425 ( \18678 , \18221 , \18677 );
xor \U$18426 ( \18679 , \18409 , \18424 );
xor \U$18427 ( \18680 , \18679 , \18431 );
and \U$18428 ( \18681 , \18678 , \18680 );
xor \U$18429 ( \18682 , \18674 , \18681 );
xor \U$18430 ( \18683 , \18303 , \18434 );
xor \U$18431 ( \18684 , \18683 , \18454 );
and \U$18432 ( \18685 , \18682 , \18684 );
and \U$18433 ( \18686 , \18674 , \18681 );
or \U$18434 ( \18687 , \18685 , \18686 );
xor \U$18435 ( \18688 , \18130 , \18457 );
xor \U$18436 ( \18689 , \18688 , \18487 );
xor \U$18437 ( \18690 , \18687 , \18689 );
and \U$18438 ( \18691 , \18354 , \18343 );
not \U$18439 ( \18692 , \18354 );
and \U$18440 ( \18693 , \18692 , \18344 );
nor \U$18441 ( \18694 , \18691 , \18693 );
xnor \U$18442 ( \18695 , \18694 , \18366 );
not \U$18443 ( \18696 , \18695 );
not \U$18444 ( \18697 , RIbe2a988_100);
not \U$18445 ( \18698 , \13690 );
or \U$18446 ( \18699 , \18697 , \18698 );
nand \U$18447 ( \18700 , RIbe2a910_99, RIbe2ae38_110);
nand \U$18448 ( \18701 , \18699 , \18700 );
xnor \U$18449 ( \18702 , \18701 , RIbe2aeb0_111);
not \U$18450 ( \18703 , RIbe2a5c8_92);
not \U$18451 ( \18704 , \12786 );
or \U$18452 ( \18705 , \18703 , \18704 );
nand \U$18453 ( \18706 , \12794 , RIbe2a550_91);
nand \U$18454 ( \18707 , \18705 , \18706 );
xor \U$18455 ( \18708 , \18707 , \12893 );
xor \U$18456 ( \18709 , \18702 , \18708 );
not \U$18457 ( \18710 , RIbe2a208_84);
not \U$18458 ( \18711 , \12831 );
or \U$18459 ( \18712 , \18710 , \18711 );
nand \U$18460 ( \18713 , \12835 , RIbe2a190_83);
nand \U$18461 ( \18714 , \18712 , \18713 );
and \U$18462 ( \18715 , \18714 , \13595 );
not \U$18463 ( \18716 , \18714 );
and \U$18464 ( \18717 , \18716 , \12823 );
or \U$18465 ( \18718 , \18715 , \18717 );
and \U$18466 ( \18719 , \18709 , \18718 );
and \U$18467 ( \18720 , \18702 , \18708 );
or \U$18468 ( \18721 , \18719 , \18720 );
not \U$18469 ( \18722 , \18721 );
not \U$18470 ( \18723 , \18722 );
and \U$18471 ( \18724 , \10916 , RIbe2ab68_104);
and \U$18472 ( \18725 , \10921 , RIbe2aaf0_103);
nor \U$18473 ( \18726 , \18724 , \18725 );
and \U$18474 ( \18727 , \18726 , \10926 );
not \U$18475 ( \18728 , \18726 );
and \U$18476 ( \18729 , \18728 , \8077 );
nor \U$18477 ( \18730 , \18727 , \18729 );
not \U$18478 ( \18731 , RIbe2b630_127);
not \U$18479 ( \18732 , \10936 );
or \U$18480 ( \18733 , \18731 , \18732 );
nand \U$18481 ( \18734 , \14511 , RIbe2b018_114);
nand \U$18482 ( \18735 , \18733 , \18734 );
and \U$18483 ( \18736 , \18735 , \9903 );
not \U$18484 ( \18737 , \18735 );
and \U$18485 ( \18738 , \18737 , \9902 );
nor \U$18486 ( \18739 , \18736 , \18738 );
nand \U$18487 ( \18740 , \18730 , \18739 );
not \U$18488 ( \18741 , \17005 );
not \U$18489 ( \18742 , RIbe2afa0_113);
not \U$18490 ( \18743 , \12943 );
or \U$18491 ( \18744 , \18742 , \18743 );
nand \U$18492 ( \18745 , \15628 , RIbe2af28_112);
nand \U$18493 ( \18746 , \18744 , \18745 );
not \U$18494 ( \18747 , \18746 );
or \U$18495 ( \18748 , \18741 , \18747 );
or \U$18496 ( \18749 , \18746 , \12960 );
nand \U$18497 ( \18750 , \18748 , \18749 );
buf \U$18498 ( \18751 , \18750 );
and \U$18499 ( \18752 , \18740 , \18751 );
nor \U$18500 ( \18753 , \18730 , \18739 );
nor \U$18501 ( \18754 , \18752 , \18753 );
not \U$18502 ( \18755 , \18754 );
not \U$18503 ( \18756 , \18755 );
or \U$18504 ( \18757 , \18723 , \18756 );
not \U$18505 ( \18758 , \18721 );
not \U$18506 ( \18759 , \18754 );
or \U$18507 ( \18760 , \18758 , \18759 );
not \U$18508 ( \18761 , RIbe2b270_119);
not \U$18509 ( \18762 , \12871 );
or \U$18510 ( \18763 , \18761 , \18762 );
nand \U$18511 ( \18764 , \12711 , RIbe2b108_116);
nand \U$18512 ( \18765 , \18763 , \18764 );
not \U$18513 ( \18766 , \18765 );
not \U$18514 ( \18767 , \12723 );
and \U$18515 ( \18768 , \18766 , \18767 );
and \U$18516 ( \18769 , \18765 , \12723 );
nor \U$18517 ( \18770 , \18768 , \18769 );
not \U$18518 ( \18771 , \18770 );
not \U$18519 ( \18772 , RIbe2b090_115);
not \U$18520 ( \18773 , \13074 );
or \U$18521 ( \18774 , \18772 , \18773 );
nand \U$18522 ( \18775 , \12735 , RIbe2a280_85);
nand \U$18523 ( \18776 , \18774 , \18775 );
and \U$18524 ( \18777 , \18776 , \14358 );
not \U$18525 ( \18778 , \18776 );
and \U$18526 ( \18779 , \18778 , \12746 );
nor \U$18527 ( \18780 , \18777 , \18779 );
or \U$18528 ( \18781 , \18771 , \18780 );
and \U$18529 ( \18782 , \17040 , RIbe2b1f8_118);
nor \U$18530 ( \18783 , \13087 , \14248 );
nor \U$18531 ( \18784 , \18782 , \18783 );
and \U$18532 ( \18785 , \18784 , \12770 );
not \U$18533 ( \18786 , \18784 );
and \U$18534 ( \18787 , \18786 , \12927 );
nor \U$18535 ( \18788 , \18785 , \18787 );
nand \U$18536 ( \18789 , \18781 , \18788 );
nand \U$18537 ( \18790 , \18780 , \18771 );
nand \U$18538 ( \18791 , \18789 , \18790 );
nand \U$18539 ( \18792 , \18760 , \18791 );
nand \U$18540 ( \18793 , \18757 , \18792 );
not \U$18541 ( \18794 , \18793 );
not \U$18542 ( \18795 , \18794 );
or \U$18543 ( \18796 , \18696 , \18795 );
not \U$18544 ( \18797 , \15233 );
not \U$18545 ( \18798 , \18797 );
and \U$18546 ( \18799 , \10916 , RIbe2aaf0_103);
and \U$18547 ( \18800 , \9914 , RIbe2b630_127);
nor \U$18548 ( \18801 , \18799 , \18800 );
not \U$18549 ( \18802 , \18801 );
or \U$18550 ( \18803 , \18798 , \18802 );
or \U$18551 ( \18804 , \18801 , \16994 );
nand \U$18552 ( \18805 , \18803 , \18804 );
not \U$18553 ( \18806 , \18805 );
nand \U$18554 ( \18807 , \10952 , RIbe2ab68_104);
and \U$18555 ( \18808 , \18807 , \14299 );
not \U$18556 ( \18809 , \18807 );
and \U$18557 ( \18810 , \18809 , \7989 );
nor \U$18558 ( \18811 , \18808 , \18810 );
nand \U$18559 ( \18812 , \18806 , \18811 );
not \U$18560 ( \18813 , \18812 );
xor \U$18561 ( \18814 , \18598 , \18587 );
xnor \U$18562 ( \18815 , \18814 , \18578 );
not \U$18563 ( \18816 , \18815 );
or \U$18564 ( \18817 , \18813 , \18816 );
not \U$18565 ( \18818 , \18811 );
nand \U$18566 ( \18819 , \18818 , \18805 );
nand \U$18567 ( \18820 , \18817 , \18819 );
nand \U$18568 ( \18821 , \18796 , \18820 );
not \U$18569 ( \18822 , \18695 );
nand \U$18570 ( \18823 , \18822 , \18793 );
nand \U$18571 ( \18824 , \18821 , \18823 );
not \U$18572 ( \18825 , \18824 );
not \U$18573 ( \18826 , \18536 );
not \U$18574 ( \18827 , \18528 );
not \U$18575 ( \18828 , \18827 );
or \U$18576 ( \18829 , \18826 , \18828 );
nand \U$18577 ( \18830 , \18528 , \18535 );
nand \U$18578 ( \18831 , \18829 , \18830 );
not \U$18579 ( \18832 , \18831 );
or \U$18580 ( \18833 , \18825 , \18832 );
or \U$18581 ( \18834 , \18824 , \18831 );
xor \U$18582 ( \18835 , \18544 , \18644 );
xnor \U$18583 ( \18836 , \18835 , \18669 );
not \U$18584 ( \18837 , \18836 );
nand \U$18585 ( \18838 , \18834 , \18837 );
nand \U$18586 ( \18839 , \18833 , \18838 );
xor \U$18587 ( \18840 , \18678 , \18680 );
xor \U$18588 ( \18841 , \18839 , \18840 );
xor \U$18589 ( \18842 , \18526 , \18537 );
xor \U$18590 ( \18843 , \18842 , \18671 );
and \U$18591 ( \18844 , \18841 , \18843 );
and \U$18592 ( \18845 , \18839 , \18840 );
or \U$18593 ( \18846 , \18844 , \18845 );
xor \U$18594 ( \18847 , \18674 , \18681 );
xor \U$18595 ( \18848 , \18847 , \18684 );
xor \U$18596 ( \18849 , \18846 , \18848 );
and \U$18597 ( \18850 , \18513 , \18520 , \18690 , \18849 );
not \U$18598 ( \18851 , \18850 );
xnor \U$18599 ( \18852 , \18770 , \18780 );
xnor \U$18600 ( \18853 , \18852 , \18788 );
not \U$18601 ( \18854 , \18853 );
xnor \U$18602 ( \18855 , \18750 , \18739 );
buf \U$18603 ( \18856 , \18730 );
xor \U$18604 ( \18857 , \18855 , \18856 );
not \U$18605 ( \18858 , \18857 );
not \U$18606 ( \18859 , \18858 );
or \U$18607 ( \18860 , \18854 , \18859 );
not \U$18608 ( \18861 , \18853 );
nand \U$18609 ( \18862 , \18861 , \18857 );
nand \U$18610 ( \18863 , \18860 , \18862 );
xor \U$18611 ( \18864 , \18702 , \18708 );
xor \U$18612 ( \18865 , \18864 , \18718 );
xnor \U$18613 ( \18866 , \18863 , \18865 );
not \U$18614 ( \18867 , \18866 );
not \U$18615 ( \18868 , RIbe2a280_85);
not \U$18616 ( \18869 , \12831 );
or \U$18617 ( \18870 , \18868 , \18869 );
nand \U$18618 ( \18871 , \12835 , RIbe2a208_84);
nand \U$18619 ( \18872 , \18870 , \18871 );
and \U$18620 ( \18873 , \18872 , \12823 );
not \U$18621 ( \18874 , \18872 );
and \U$18622 ( \18875 , \18874 , \14555 );
nor \U$18623 ( \18876 , \18873 , \18875 );
not \U$18624 ( \18877 , RIbe2b180_117);
not \U$18625 ( \18878 , \12871 );
or \U$18626 ( \18879 , \18877 , \18878 );
nand \U$18627 ( \18880 , \13728 , RIbe2b270_119);
nand \U$18628 ( \18881 , \18879 , \18880 );
not \U$18629 ( \18882 , \18881 );
not \U$18630 ( \18883 , \12723 );
and \U$18631 ( \18884 , \18882 , \18883 );
and \U$18632 ( \18885 , \12723 , \18881 );
nor \U$18633 ( \18886 , \18884 , \18885 );
xor \U$18634 ( \18887 , \18876 , \18886 );
not \U$18635 ( \18888 , RIbe2b108_116);
not \U$18636 ( \18889 , \14071 );
or \U$18637 ( \18890 , \18888 , \18889 );
nand \U$18638 ( \18891 , \13077 , RIbe2b090_115);
nand \U$18639 ( \18892 , \18890 , \18891 );
and \U$18640 ( \18893 , \18892 , \12746 );
not \U$18641 ( \18894 , \18892 );
and \U$18642 ( \18895 , \18894 , \12852 );
nor \U$18643 ( \18896 , \18893 , \18895 );
xor \U$18644 ( \18897 , \18887 , \18896 );
nand \U$18645 ( \18898 , \17547 , RIbe2ab68_104);
and \U$18646 ( \18899 , \18898 , \16994 );
not \U$18647 ( \18900 , \18898 );
and \U$18648 ( \18901 , \18900 , \15233 );
nor \U$18649 ( \18902 , \18899 , \18901 );
and \U$18650 ( \18903 , \18897 , \18902 );
not \U$18651 ( \18904 , RIbe2b018_114);
not \U$18652 ( \18905 , \15205 );
or \U$18653 ( \18906 , \18904 , \18905 );
nand \U$18654 ( \18907 , \13669 , RIbe2afa0_113);
nand \U$18655 ( \18908 , \18906 , \18907 );
not \U$18656 ( \18909 , \18908 );
not \U$18657 ( \18910 , \12960 );
and \U$18658 ( \18911 , \18909 , \18910 );
and \U$18659 ( \18912 , \18908 , \12956 );
nor \U$18660 ( \18913 , \18911 , \18912 );
not \U$18661 ( \18914 , \12751 );
not \U$18662 ( \18915 , \14645 );
and \U$18663 ( \18916 , \18914 , \18915 );
and \U$18664 ( \18917 , \14726 , RIbe2af28_112);
nor \U$18665 ( \18918 , \18916 , \18917 );
and \U$18666 ( \18919 , \18918 , \12924 );
not \U$18667 ( \18920 , \18918 );
and \U$18668 ( \18921 , \18920 , \12774 );
nor \U$18669 ( \18922 , \18919 , \18921 );
and \U$18670 ( \18923 , \18913 , \18922 );
not \U$18671 ( \18924 , \18913 );
not \U$18672 ( \18925 , \18922 );
and \U$18673 ( \18926 , \18924 , \18925 );
or \U$18674 ( \18927 , \18923 , \18926 );
not \U$18675 ( \18928 , RIbe2aaf0_103);
not \U$18676 ( \18929 , \10936 );
or \U$18677 ( \18930 , \18928 , \18929 );
nand \U$18678 ( \18931 , \12213 , RIbe2b630_127);
nand \U$18679 ( \18932 , \18930 , \18931 );
not \U$18680 ( \18933 , \18932 );
not \U$18681 ( \18934 , \13030 );
and \U$18682 ( \18935 , \18933 , \18934 );
and \U$18683 ( \18936 , \18932 , \9903 );
nor \U$18684 ( \18937 , \18935 , \18936 );
xor \U$18685 ( \18938 , \18927 , \18937 );
nor \U$18686 ( \18939 , \18903 , \18938 );
nor \U$18687 ( \18940 , \18897 , \18902 );
nor \U$18688 ( \18941 , \18939 , \18940 );
not \U$18689 ( \18942 , \18941 );
not \U$18690 ( \18943 , RIbe2ab68_104);
not \U$18691 ( \18944 , \10936 );
or \U$18692 ( \18945 , \18943 , \18944 );
nand \U$18693 ( \18946 , \12971 , RIbe2aaf0_103);
nand \U$18694 ( \18947 , \18945 , \18946 );
and \U$18695 ( \18948 , \18947 , \9902 );
not \U$18696 ( \18949 , \18947 );
and \U$18697 ( \18950 , \18949 , \12219 );
nor \U$18698 ( \18951 , \18948 , \18950 );
not \U$18699 ( \18952 , \12960 );
not \U$18700 ( \18953 , RIbe2b630_127);
not \U$18701 ( \18954 , \12943 );
or \U$18702 ( \18955 , \18953 , \18954 );
nand \U$18703 ( \18956 , \12948 , RIbe2b018_114);
nand \U$18704 ( \18957 , \18955 , \18956 );
not \U$18705 ( \18958 , \18957 );
or \U$18706 ( \18959 , \18952 , \18958 );
or \U$18707 ( \18960 , \18957 , \12956 );
nand \U$18708 ( \18961 , \18959 , \18960 );
nand \U$18709 ( \18962 , \18951 , \18961 );
not \U$18710 ( \18963 , \18962 );
not \U$18711 ( \18964 , RIbe2a5c8_92);
not \U$18712 ( \18965 , \12811 );
or \U$18713 ( \18966 , \18964 , \18965 );
nand \U$18714 ( \18967 , RIbe2a550_91, RIbe2ae38_110);
nand \U$18715 ( \18968 , \18966 , \18967 );
xnor \U$18716 ( \18969 , \18968 , RIbe2aeb0_111);
not \U$18717 ( \18970 , RIbe2a208_84);
not \U$18718 ( \18971 , \15249 );
or \U$18719 ( \18972 , \18970 , \18971 );
nand \U$18720 ( \18973 , \12890 , RIbe2a190_83);
nand \U$18721 ( \18974 , \18972 , \18973 );
xor \U$18722 ( \18975 , \18974 , \12893 );
xor \U$18723 ( \18976 , \18969 , \18975 );
not \U$18724 ( \18977 , RIbe2b090_115);
not \U$18725 ( \18978 , \13010 );
or \U$18726 ( \18979 , \18977 , \18978 );
nand \U$18727 ( \18980 , \12835 , RIbe2a280_85);
nand \U$18728 ( \18981 , \18979 , \18980 );
and \U$18729 ( \18982 , \18981 , \15263 );
not \U$18730 ( \18983 , \18981 );
and \U$18731 ( \18984 , \18983 , \18364 );
nor \U$18732 ( \18985 , \18982 , \18984 );
and \U$18733 ( \18986 , \18976 , \18985 );
and \U$18734 ( \18987 , \18969 , \18975 );
or \U$18735 ( \18988 , \18986 , \18987 );
not \U$18736 ( \18989 , \18988 );
or \U$18737 ( \18990 , \18963 , \18989 );
not \U$18738 ( \18991 , RIbe2b270_119);
not \U$18739 ( \18992 , \14071 );
or \U$18740 ( \18993 , \18991 , \18992 );
nand \U$18741 ( \18994 , \14074 , RIbe2b108_116);
nand \U$18742 ( \18995 , \18993 , \18994 );
and \U$18743 ( \18996 , \18995 , \12742 );
not \U$18744 ( \18997 , \18995 );
and \U$18745 ( \18998 , \18997 , \15166 );
nor \U$18746 ( \18999 , \18996 , \18998 );
not \U$18747 ( \19000 , \18999 );
not \U$18748 ( \19001 , \19000 );
not \U$18749 ( \19002 , RIbe2b1f8_118);
not \U$18750 ( \19003 , \13063 );
or \U$18751 ( \19004 , \19002 , \19003 );
nand \U$18752 ( \19005 , \13728 , RIbe2b180_117);
nand \U$18753 ( \19006 , \19004 , \19005 );
and \U$18754 ( \19007 , \19006 , \12723 );
not \U$18755 ( \19008 , \19006 );
and \U$18756 ( \19009 , \19008 , \12716 );
nor \U$18757 ( \19010 , \19007 , \19009 );
not \U$18758 ( \19011 , \19010 );
not \U$18759 ( \19012 , \19011 );
or \U$18760 ( \19013 , \19001 , \19012 );
and \U$18761 ( \19014 , \12765 , RIbe2afa0_113);
not \U$18762 ( \19015 , RIbe2af28_112);
nor \U$18763 ( \19016 , \19015 , \13087 );
nor \U$18764 ( \19017 , \19014 , \19016 );
and \U$18765 ( \19018 , \19017 , \12774 );
not \U$18766 ( \19019 , \19017 );
and \U$18767 ( \19020 , \19019 , \12924 );
nor \U$18768 ( \19021 , \19018 , \19020 );
not \U$18769 ( \19022 , \19021 );
nand \U$18770 ( \19023 , \18999 , \19010 );
nand \U$18771 ( \19024 , \19022 , \19023 );
nand \U$18772 ( \19025 , \19013 , \19024 );
nand \U$18773 ( \19026 , \18990 , \19025 );
or \U$18774 ( \19027 , \18962 , \18988 );
nand \U$18775 ( \19028 , \19026 , \19027 );
not \U$18776 ( \19029 , \19028 );
and \U$18777 ( \19030 , \18942 , \19029 );
and \U$18778 ( \19031 , \18941 , \19028 );
nor \U$18779 ( \19032 , \19030 , \19031 );
not \U$18780 ( \19033 , \19032 );
or \U$18781 ( \19034 , \18867 , \19033 );
or \U$18782 ( \19035 , \18866 , \19032 );
nand \U$18783 ( \19036 , \19034 , \19035 );
xor \U$18784 ( \19037 , \18876 , \18886 );
and \U$18785 ( \19038 , \19037 , \18896 );
and \U$18786 ( \19039 , \18876 , \18886 );
or \U$18787 ( \19040 , \19038 , \19039 );
not \U$18788 ( \19041 , \19040 );
and \U$18789 ( \19042 , \18937 , \18925 );
nor \U$18790 ( \19043 , \19042 , \18913 );
nor \U$18791 ( \19044 , \18925 , \18937 );
nor \U$18792 ( \19045 , \19043 , \19044 );
not \U$18793 ( \19046 , RIbe2a190_83);
not \U$18794 ( \19047 , \13518 );
or \U$18795 ( \19048 , \19046 , \19047 );
nand \U$18796 ( \19049 , \12890 , RIbe2a5c8_92);
nand \U$18797 ( \19050 , \19048 , \19049 );
and \U$18798 ( \19051 , \19050 , \12893 );
not \U$18799 ( \19052 , \19050 );
and \U$18800 ( \19053 , \19052 , \12995 );
nor \U$18801 ( \19054 , \19051 , \19053 );
not \U$18802 ( \19055 , RIbe2a550_91);
not \U$18803 ( \19056 , \12811 );
or \U$18804 ( \19057 , \19055 , \19056 );
nand \U$18805 ( \19058 , RIbe2a988_100, RIbe2ae38_110);
nand \U$18806 ( \19059 , \19057 , \19058 );
xor \U$18807 ( \19060 , \19059 , RIbe2aeb0_111);
nor \U$18808 ( \19061 , \19060 , \7970 );
nor \U$18809 ( \19062 , \19054 , \19061 );
and \U$18810 ( \19063 , \19060 , \16994 );
nor \U$18811 ( \19064 , \19062 , \19063 );
and \U$18812 ( \19065 , \19045 , \19064 );
not \U$18813 ( \19066 , \19045 );
not \U$18814 ( \19067 , \19064 );
and \U$18815 ( \19068 , \19066 , \19067 );
nor \U$18816 ( \19069 , \19065 , \19068 );
not \U$18817 ( \19070 , \19069 );
or \U$18818 ( \19071 , \19041 , \19070 );
or \U$18819 ( \19072 , \19069 , \19040 );
nand \U$18820 ( \19073 , \19071 , \19072 );
and \U$18821 ( \19074 , \19060 , \7971 );
not \U$18822 ( \19075 , \19060 );
and \U$18823 ( \19076 , \19075 , \7970 );
nor \U$18824 ( \19077 , \19074 , \19076 );
not \U$18825 ( \19078 , \19077 );
not \U$18826 ( \19079 , \19054 );
not \U$18827 ( \19080 , \19079 );
or \U$18828 ( \19081 , \19078 , \19080 );
or \U$18829 ( \19082 , \19079 , \19077 );
nand \U$18830 ( \19083 , \19081 , \19082 );
not \U$18831 ( \19084 , RIbe2af28_112);
not \U$18832 ( \19085 , \15573 );
or \U$18833 ( \19086 , \19084 , \19085 );
nand \U$18834 ( \19087 , \12711 , RIbe2b1f8_118);
nand \U$18835 ( \19088 , \19086 , \19087 );
and \U$18836 ( \19089 , \19088 , \12723 );
not \U$18837 ( \19090 , \19088 );
and \U$18838 ( \19091 , \19090 , \12716 );
nor \U$18839 ( \19092 , \19089 , \19091 );
not \U$18840 ( \19093 , RIbe2b108_116);
not \U$18841 ( \19094 , \12831 );
or \U$18842 ( \19095 , \19093 , \19094 );
nand \U$18843 ( \19096 , \13012 , RIbe2b090_115);
nand \U$18844 ( \19097 , \19095 , \19096 );
and \U$18845 ( \19098 , \19097 , \12863 );
not \U$18846 ( \19099 , \19097 );
and \U$18847 ( \19100 , \19099 , \12866 );
nor \U$18848 ( \19101 , \19098 , \19100 );
and \U$18849 ( \19102 , \19092 , \19101 );
not \U$18850 ( \19103 , RIbe2b180_117);
not \U$18851 ( \19104 , \12732 );
or \U$18852 ( \19105 , \19103 , \19104 );
nand \U$18853 ( \19106 , \14074 , RIbe2b270_119);
nand \U$18854 ( \19107 , \19105 , \19106 );
and \U$18855 ( \19108 , \19107 , \14077 );
not \U$18856 ( \19109 , \19107 );
and \U$18857 ( \19110 , \19109 , \12746 );
nor \U$18858 ( \19111 , \19108 , \19110 );
not \U$18859 ( \19112 , \19111 );
nor \U$18860 ( \19113 , \19102 , \19112 );
nor \U$18861 ( \19114 , \19092 , \19101 );
nor \U$18862 ( \19115 , \19113 , \19114 );
not \U$18863 ( \19116 , RIbe2a190_83);
not \U$18864 ( \19117 , \12811 );
or \U$18865 ( \19118 , \19116 , \19117 );
nand \U$18866 ( \19119 , RIbe2a5c8_92, RIbe2ae38_110);
nand \U$18867 ( \19120 , \19118 , \19119 );
xnor \U$18868 ( \19121 , \19120 , RIbe2aeb0_111);
xor \U$18869 ( \19122 , \9903 , \19121 );
not \U$18870 ( \19123 , RIbe2a280_85);
not \U$18871 ( \19124 , \12887 );
or \U$18872 ( \19125 , \19123 , \19124 );
nand \U$18873 ( \19126 , \12890 , RIbe2a208_84);
nand \U$18874 ( \19127 , \19125 , \19126 );
xor \U$18875 ( \19128 , \19127 , \12893 );
and \U$18876 ( \19129 , \19122 , \19128 );
and \U$18877 ( \19130 , \9903 , \19121 );
or \U$18878 ( \19131 , \19129 , \19130 );
nand \U$18879 ( \19132 , \19115 , \19131 );
not \U$18880 ( \19133 , \19132 );
nand \U$18881 ( \19134 , \14511 , RIbe2ab68_104);
not \U$18882 ( \19135 , \19134 );
not \U$18883 ( \19136 , \10940 );
not \U$18884 ( \19137 , \19136 );
or \U$18885 ( \19138 , \19135 , \19137 );
not \U$18886 ( \19139 , \13033 );
or \U$18887 ( \19140 , \19134 , \19139 );
nand \U$18888 ( \19141 , \19138 , \19140 );
not \U$18889 ( \19142 , \12770 );
not \U$18890 ( \19143 , RIbe2b018_114);
not \U$18891 ( \19144 , \17040 );
or \U$18892 ( \19145 , \19143 , \19144 );
not \U$18893 ( \19146 , \12752 );
nand \U$18894 ( \19147 , \19146 , RIbe2afa0_113);
nand \U$18895 ( \19148 , \19145 , \19147 );
not \U$18896 ( \19149 , \19148 );
or \U$18897 ( \19150 , \19142 , \19149 );
or \U$18898 ( \19151 , \19148 , \12769 );
nand \U$18899 ( \19152 , \19150 , \19151 );
xor \U$18900 ( \19153 , \19141 , \19152 );
and \U$18901 ( \19154 , \12948 , RIbe2b630_127);
and \U$18902 ( \19155 , \12943 , RIbe2aaf0_103);
nor \U$18903 ( \19156 , \19154 , \19155 );
and \U$18904 ( \19157 , \19156 , \12195 );
not \U$18905 ( \19158 , \19156 );
and \U$18906 ( \19159 , \19158 , \12956 );
or \U$18907 ( \19160 , \19157 , \19159 );
and \U$18908 ( \19161 , \19153 , \19160 );
and \U$18909 ( \19162 , \19141 , \19152 );
or \U$18910 ( \19163 , \19161 , \19162 );
not \U$18911 ( \19164 , \19163 );
or \U$18912 ( \19165 , \19133 , \19164 );
not \U$18913 ( \19166 , \19131 );
not \U$18914 ( \19167 , \19115 );
nand \U$18915 ( \19168 , \19166 , \19167 );
nand \U$18916 ( \19169 , \19165 , \19168 );
xor \U$18917 ( \19170 , \19083 , \19169 );
xor \U$18918 ( \19171 , \18969 , \18975 );
xor \U$18919 ( \19172 , \19171 , \18985 );
xnor \U$18920 ( \19173 , \18951 , \18961 );
nand \U$18921 ( \19174 , \19172 , \19173 );
not \U$18922 ( \19175 , \19021 );
nand \U$18923 ( \19176 , \19000 , \19010 );
nand \U$18924 ( \19177 , \18999 , \19011 );
nand \U$18925 ( \19178 , \19176 , \19177 );
not \U$18926 ( \19179 , \19178 );
or \U$18927 ( \19180 , \19175 , \19179 );
or \U$18928 ( \19181 , \19178 , \19021 );
nand \U$18929 ( \19182 , \19180 , \19181 );
nand \U$18930 ( \19183 , \19174 , \19182 );
or \U$18931 ( \19184 , \19172 , \19173 );
nand \U$18932 ( \19185 , \19183 , \19184 );
and \U$18933 ( \19186 , \19170 , \19185 );
and \U$18934 ( \19187 , \19083 , \19169 );
or \U$18935 ( \19188 , \19186 , \19187 );
xor \U$18936 ( \19189 , \19073 , \19188 );
xor \U$18937 ( \19190 , \18962 , \18988 );
xor \U$18938 ( \19191 , \19190 , \19025 );
not \U$18939 ( \19192 , \18938 );
xor \U$18940 ( \19193 , \18897 , \18902 );
not \U$18941 ( \19194 , \19193 );
or \U$18942 ( \19195 , \19192 , \19194 );
or \U$18943 ( \19196 , \19193 , \18938 );
nand \U$18944 ( \19197 , \19195 , \19196 );
and \U$18945 ( \19198 , \19191 , \19197 );
xor \U$18946 ( \19199 , \19189 , \19198 );
xor \U$18947 ( \19200 , \19036 , \19199 );
xor \U$18948 ( \19201 , \19191 , \19197 );
not \U$18949 ( \19202 , \19201 );
xor \U$18950 ( \19203 , \19173 , \19172 );
xnor \U$18951 ( \19204 , \19203 , \19182 );
xor \U$18952 ( \19205 , \9903 , \19121 );
xor \U$18953 ( \19206 , \19205 , \19128 );
not \U$18954 ( \19207 , \19206 );
and \U$18955 ( \19208 , \19101 , \19111 );
not \U$18956 ( \19209 , \19101 );
and \U$18957 ( \19210 , \19209 , \19112 );
or \U$18958 ( \19211 , \19208 , \19210 );
xnor \U$18959 ( \19212 , \19211 , \19092 );
nand \U$18960 ( \19213 , \19207 , \19212 );
nand \U$18961 ( \19214 , \19204 , \19213 );
not \U$18962 ( \19215 , \19214 );
not \U$18963 ( \19216 , RIbe2a208_84);
not \U$18964 ( \19217 , \13004 );
or \U$18965 ( \19218 , \19216 , \19217 );
nand \U$18966 ( \19219 , RIbe2a190_83, RIbe2ae38_110);
nand \U$18967 ( \19220 , \19218 , \19219 );
xnor \U$18968 ( \19221 , \19220 , RIbe2aeb0_111);
not \U$18969 ( \19222 , \19221 );
not \U$18970 ( \19223 , RIbe2b090_115);
not \U$18971 ( \19224 , \12887 );
or \U$18972 ( \19225 , \19223 , \19224 );
nand \U$18973 ( \19226 , \12890 , RIbe2a280_85);
nand \U$18974 ( \19227 , \19225 , \19226 );
and \U$18975 ( \19228 , \19227 , \12998 );
not \U$18976 ( \19229 , \19227 );
and \U$18977 ( \19230 , \19229 , \16334 );
nor \U$18978 ( \19231 , \19228 , \19230 );
not \U$18979 ( \19232 , \19231 );
or \U$18980 ( \19233 , \19222 , \19232 );
not \U$18981 ( \19234 , \15263 );
not \U$18982 ( \19235 , RIbe2b270_119);
not \U$18983 ( \19236 , \12831 );
or \U$18984 ( \19237 , \19235 , \19236 );
nand \U$18985 ( \19238 , \12835 , RIbe2b108_116);
nand \U$18986 ( \19239 , \19237 , \19238 );
not \U$18987 ( \19240 , \19239 );
or \U$18988 ( \19241 , \19234 , \19240 );
or \U$18989 ( \19242 , \19239 , \13706 );
nand \U$18990 ( \19243 , \19241 , \19242 );
nand \U$18991 ( \19244 , \19233 , \19243 );
not \U$18992 ( \19245 , \19221 );
not \U$18993 ( \19246 , \19231 );
nand \U$18994 ( \19247 , \19245 , \19246 );
nand \U$18995 ( \19248 , \19244 , \19247 );
not \U$18996 ( \19249 , RIbe2b1f8_118);
not \U$18997 ( \19250 , \14071 );
or \U$18998 ( \19251 , \19249 , \19250 );
nand \U$18999 ( \19252 , \14074 , RIbe2b180_117);
nand \U$19000 ( \19253 , \19251 , \19252 );
not \U$19001 ( \19254 , \19253 );
not \U$19002 ( \19255 , \12746 );
and \U$19003 ( \19256 , \19254 , \19255 );
and \U$19004 ( \19257 , \19253 , \12741 );
nor \U$19005 ( \19258 , \19256 , \19257 );
not \U$19006 ( \19259 , \19258 );
not \U$19007 ( \19260 , \19259 );
not \U$19008 ( \19261 , RIbe2afa0_113);
not \U$19009 ( \19262 , \12706 );
not \U$19010 ( \19263 , \19262 );
or \U$19011 ( \19264 , \19261 , \19263 );
nand \U$19012 ( \19265 , \13728 , RIbe2af28_112);
nand \U$19013 ( \19266 , \19264 , \19265 );
and \U$19014 ( \19267 , \19266 , \12723 );
not \U$19015 ( \19268 , \19266 );
and \U$19016 ( \19269 , \19268 , \12879 );
nor \U$19017 ( \19270 , \19267 , \19269 );
not \U$19018 ( \19271 , \19270 );
not \U$19019 ( \19272 , \19271 );
or \U$19020 ( \19273 , \19260 , \19272 );
not \U$19021 ( \19274 , \19258 );
not \U$19022 ( \19275 , \19270 );
or \U$19023 ( \19276 , \19274 , \19275 );
and \U$19024 ( \19277 , \17040 , RIbe2b630_127);
and \U$19025 ( \19278 , \13086 , RIbe2b018_114);
nor \U$19026 ( \19279 , \19277 , \19278 );
and \U$19027 ( \19280 , \19279 , \12924 );
not \U$19028 ( \19281 , \19279 );
and \U$19029 ( \19282 , \19281 , \12927 );
nor \U$19030 ( \19283 , \19280 , \19282 );
nand \U$19031 ( \19284 , \19276 , \19283 );
nand \U$19032 ( \19285 , \19273 , \19284 );
xor \U$19033 ( \19286 , \19248 , \19285 );
xor \U$19034 ( \19287 , \19141 , \19152 );
xor \U$19035 ( \19288 , \19287 , \19160 );
and \U$19036 ( \19289 , \19286 , \19288 );
and \U$19037 ( \19290 , \19248 , \19285 );
or \U$19038 ( \19291 , \19289 , \19290 );
not \U$19039 ( \19292 , \19291 );
or \U$19040 ( \19293 , \19215 , \19292 );
or \U$19041 ( \19294 , \19204 , \19213 );
nand \U$19042 ( \19295 , \19293 , \19294 );
not \U$19043 ( \19296 , \19295 );
or \U$19044 ( \19297 , \19202 , \19296 );
or \U$19045 ( \19298 , \19295 , \19201 );
xor \U$19046 ( \19299 , \19083 , \19169 );
xor \U$19047 ( \19300 , \19299 , \19185 );
nand \U$19048 ( \19301 , \19298 , \19300 );
nand \U$19049 ( \19302 , \19297 , \19301 );
nand \U$19050 ( \19303 , \19200 , \19302 );
not \U$19051 ( \19304 , \19303 );
and \U$19052 ( \19305 , \19036 , \19199 );
buf \U$19053 ( \19306 , \19305 );
not \U$19054 ( \19307 , \19306 );
xor \U$19055 ( \19308 , \19073 , \19188 );
and \U$19056 ( \19309 , \19308 , \19198 );
and \U$19057 ( \19310 , \19073 , \19188 );
or \U$19058 ( \19311 , \19309 , \19310 );
nand \U$19059 ( \19312 , \18853 , \18865 );
and \U$19060 ( \19313 , \19312 , \18858 );
nor \U$19061 ( \19314 , \18853 , \18865 );
nor \U$19062 ( \19315 , \19313 , \19314 );
xor \U$19063 ( \19316 , \18616 , \18640 );
xor \U$19064 ( \19317 , \19316 , \18627 );
not \U$19065 ( \19318 , \19064 );
not \U$19066 ( \19319 , \19040 );
or \U$19067 ( \19320 , \19318 , \19319 );
not \U$19068 ( \19321 , \19045 );
nand \U$19069 ( \19322 , \19320 , \19321 );
not \U$19070 ( \19323 , \19040 );
nand \U$19071 ( \19324 , \19323 , \19067 );
nand \U$19072 ( \19325 , \19322 , \19324 );
xor \U$19073 ( \19326 , \19317 , \19325 );
xnor \U$19074 ( \19327 , \19315 , \19326 );
not \U$19075 ( \19328 , \19028 );
nand \U$19076 ( \19329 , \19328 , \18941 );
and \U$19077 ( \19330 , \18866 , \19329 );
not \U$19078 ( \19331 , \19028 );
nor \U$19079 ( \19332 , \19331 , \18941 );
nor \U$19080 ( \19333 , \19330 , \19332 );
xnor \U$19081 ( \19334 , \19327 , \19333 );
not \U$19082 ( \19335 , \18554 );
and \U$19083 ( \19336 , \18565 , \6949 );
not \U$19084 ( \19337 , \18565 );
and \U$19085 ( \19338 , \19337 , \7988 );
nor \U$19086 ( \19339 , \19336 , \19338 );
not \U$19087 ( \19340 , \19339 );
and \U$19088 ( \19341 , \19335 , \19340 );
and \U$19089 ( \19342 , \18554 , \19339 );
nor \U$19090 ( \19343 , \19341 , \19342 );
not \U$19091 ( \19344 , \18815 );
not \U$19092 ( \19345 , \18805 );
not \U$19093 ( \19346 , \18811 );
and \U$19094 ( \19347 , \19345 , \19346 );
and \U$19095 ( \19348 , \18805 , \18811 );
nor \U$19096 ( \19349 , \19347 , \19348 );
not \U$19097 ( \19350 , \19349 );
and \U$19098 ( \19351 , \19344 , \19350 );
and \U$19099 ( \19352 , \18815 , \19349 );
nor \U$19100 ( \19353 , \19351 , \19352 );
xor \U$19101 ( \19354 , \19343 , \19353 );
and \U$19102 ( \19355 , \18791 , \18755 );
not \U$19103 ( \19356 , \18791 );
and \U$19104 ( \19357 , \19356 , \18754 );
nor \U$19105 ( \19358 , \19355 , \19357 );
and \U$19106 ( \19359 , \19358 , \18721 );
not \U$19107 ( \19360 , \19358 );
and \U$19108 ( \19361 , \19360 , \18722 );
nor \U$19109 ( \19362 , \19359 , \19361 );
xor \U$19110 ( \19363 , \19354 , \19362 );
not \U$19111 ( \19364 , \19363 );
and \U$19112 ( \19365 , \19334 , \19364 );
not \U$19113 ( \19366 , \19334 );
and \U$19114 ( \19367 , \19366 , \19363 );
nor \U$19115 ( \19368 , \19365 , \19367 );
xor \U$19116 ( \19369 , \19311 , \19368 );
not \U$19117 ( \19370 , \19369 );
not \U$19118 ( \19371 , \19370 );
or \U$19119 ( \19372 , \19307 , \19371 );
not \U$19120 ( \19373 , \19305 );
nand \U$19121 ( \19374 , \19373 , \19369 );
nand \U$19122 ( \19375 , \19372 , \19374 );
nand \U$19123 ( \19376 , \19304 , \19375 );
nand \U$19124 ( \19377 , \19369 , \19306 );
nand \U$19125 ( \19378 , \19376 , \19377 );
not \U$19126 ( \19379 , \19378 );
xor \U$19127 ( \19380 , \18839 , \18840 );
xor \U$19128 ( \19381 , \19380 , \18843 );
not \U$19129 ( \19382 , \19381 );
xor \U$19130 ( \19383 , \18601 , \18567 );
xor \U$19131 ( \19384 , \19383 , \18642 );
not \U$19132 ( \19385 , \19384 );
not \U$19133 ( \19386 , \18820 );
not \U$19134 ( \19387 , \18695 );
and \U$19135 ( \19388 , \19386 , \19387 );
and \U$19136 ( \19389 , \18820 , \18695 );
nor \U$19137 ( \19390 , \19388 , \19389 );
and \U$19138 ( \19391 , \19390 , \18794 );
not \U$19139 ( \19392 , \19390 );
and \U$19140 ( \19393 , \19392 , \18793 );
nor \U$19141 ( \19394 , \19391 , \19393 );
nand \U$19142 ( \19395 , \19385 , \19394 );
xor \U$19143 ( \19396 , \18656 , \18666 );
xor \U$19144 ( \19397 , \19396 , \18649 );
not \U$19145 ( \19398 , \19317 );
not \U$19146 ( \19399 , \19325 );
and \U$19147 ( \19400 , \19398 , \19399 );
nor \U$19148 ( \19401 , \19400 , \19315 );
and \U$19149 ( \19402 , \19317 , \19325 );
nor \U$19150 ( \19403 , \19401 , \19402 );
xor \U$19151 ( \19404 , \19397 , \19403 );
xor \U$19152 ( \19405 , \19343 , \19353 );
and \U$19153 ( \19406 , \19405 , \19362 );
and \U$19154 ( \19407 , \19343 , \19353 );
or \U$19155 ( \19408 , \19406 , \19407 );
and \U$19156 ( \19409 , \19404 , \19408 );
and \U$19157 ( \19410 , \19397 , \19403 );
or \U$19158 ( \19411 , \19409 , \19410 );
xor \U$19159 ( \19412 , \19395 , \19411 );
xor \U$19160 ( \19413 , \18824 , \18831 );
xor \U$19161 ( \19414 , \19413 , \18836 );
and \U$19162 ( \19415 , \19412 , \19414 );
and \U$19163 ( \19416 , \19395 , \19411 );
or \U$19164 ( \19417 , \19415 , \19416 );
not \U$19165 ( \19418 , \19417 );
and \U$19166 ( \19419 , \19382 , \19418 );
and \U$19167 ( \19420 , \19381 , \19417 );
nor \U$19168 ( \19421 , \19419 , \19420 );
not \U$19169 ( \19422 , \19421 );
xor \U$19170 ( \19423 , \19397 , \19403 );
xor \U$19171 ( \19424 , \19423 , \19408 );
not \U$19172 ( \19425 , \19424 );
not \U$19173 ( \19426 , \19425 );
not \U$19174 ( \19427 , \19333 );
not \U$19175 ( \19428 , \19363 );
or \U$19176 ( \19429 , \19427 , \19428 );
nand \U$19177 ( \19430 , \19429 , \19327 );
not \U$19178 ( \19431 , \19333 );
nand \U$19179 ( \19432 , \19431 , \19364 );
nand \U$19180 ( \19433 , \19430 , \19432 );
not \U$19181 ( \19434 , \19433 );
not \U$19182 ( \19435 , \19434 );
or \U$19183 ( \19436 , \19426 , \19435 );
nand \U$19184 ( \19437 , \19433 , \19424 );
nand \U$19185 ( \19438 , \19436 , \19437 );
not \U$19186 ( \19439 , \19438 );
xor \U$19187 ( \19440 , \18793 , \19384 );
xnor \U$19188 ( \19441 , \19440 , \19390 );
not \U$19189 ( \19442 , \19441 );
and \U$19190 ( \19443 , \19439 , \19442 );
and \U$19191 ( \19444 , \19438 , \19441 );
nor \U$19192 ( \19445 , \19443 , \19444 );
not \U$19193 ( \19446 , \19445 );
and \U$19194 ( \19447 , \19311 , \19368 );
not \U$19195 ( \19448 , \19447 );
or \U$19196 ( \19449 , \19446 , \19448 );
or \U$19197 ( \19450 , \19445 , \19447 );
nand \U$19198 ( \19451 , \19449 , \19450 );
xor \U$19199 ( \19452 , \19395 , \19411 );
xor \U$19200 ( \19453 , \19452 , \19414 );
not \U$19201 ( \19454 , \19453 );
not \U$19202 ( \19455 , \19454 );
not \U$19203 ( \19456 , \19441 );
not \U$19204 ( \19457 , \19434 );
or \U$19205 ( \19458 , \19456 , \19457 );
nand \U$19206 ( \19459 , \19458 , \19425 );
not \U$19207 ( \19460 , \19441 );
nand \U$19208 ( \19461 , \19460 , \19433 );
nand \U$19209 ( \19462 , \19459 , \19461 );
not \U$19210 ( \19463 , \19462 );
not \U$19211 ( \19464 , \19463 );
or \U$19212 ( \19465 , \19455 , \19464 );
nand \U$19213 ( \19466 , \19462 , \19453 );
nand \U$19214 ( \19467 , \19465 , \19466 );
and \U$19215 ( \19468 , \19422 , \19451 , \19467 );
not \U$19216 ( \19469 , \19468 );
or \U$19217 ( \19470 , \19379 , \19469 );
not \U$19218 ( \19471 , \19445 );
nand \U$19219 ( \19472 , \19471 , \19447 );
nor \U$19220 ( \19473 , \19421 , \19472 );
and \U$19221 ( \19474 , \19467 , \19473 );
nand \U$19222 ( \19475 , \19454 , \19462 );
or \U$19223 ( \19476 , \19421 , \19475 );
not \U$19224 ( \19477 , \19381 );
or \U$19225 ( \19478 , \19477 , \19417 );
nand \U$19226 ( \19479 , \19476 , \19478 );
nor \U$19227 ( \19480 , \19474 , \19479 );
nand \U$19228 ( \19481 , \19470 , \19480 );
not \U$19229 ( \19482 , \19481 );
or \U$19230 ( \19483 , \18851 , \19482 );
not \U$19231 ( \19484 , \18517 );
not \U$19232 ( \19485 , \18519 );
and \U$19233 ( \19486 , \19484 , \19485 );
and \U$19234 ( \19487 , \18846 , \18848 );
and \U$19235 ( \19488 , \18690 , \19487 );
and \U$19236 ( \19489 , \18687 , \18689 );
nor \U$19237 ( \19490 , \19488 , \19489 );
not \U$19238 ( \19491 , \18513 );
or \U$19239 ( \19492 , \19490 , \19491 );
not \U$19240 ( \19493 , \18491 );
nand \U$19241 ( \19494 , \19493 , \18509 );
nand \U$19242 ( \19495 , \19492 , \19494 );
and \U$19243 ( \19496 , \19495 , \18520 );
nor \U$19244 ( \19497 , \19486 , \19496 );
nand \U$19245 ( \19498 , \19483 , \19497 );
nand \U$19246 ( \19499 , \18099 , \18104 );
nor \U$19247 ( \19500 , \19499 , \17657 );
xor \U$19248 ( \19501 , \18078 , \18087 );
and \U$19249 ( \19502 , \18126 , \19501 );
nand \U$19250 ( \19503 , \19498 , \19500 , \19502 );
nand \U$19251 ( \19504 , \18116 , \18121 );
nand \U$19252 ( \19505 , \18128 , \19503 , \19504 );
not \U$19253 ( \19506 , \16920 );
not \U$19254 ( \19507 , \15763 );
not \U$19255 ( \19508 , \16870 );
xor \U$19256 ( \19509 , \14709 , \14716 );
not \U$19257 ( \19510 , \14450 );
nor \U$19258 ( \19511 , \19509 , \19510 );
and \U$19259 ( \19512 , \19506 , \19507 , \19508 , \19511 );
nand \U$19260 ( \19513 , \19505 , \19512 );
not \U$19261 ( \19514 , \19421 );
and \U$19262 ( \19515 , \19514 , \19451 , \19467 , \19375 );
xor \U$19263 ( \19516 , \19200 , \19302 );
and \U$19264 ( \19517 , \19515 , \18850 , \19516 );
not \U$19265 ( \19518 , \12195 );
and \U$19266 ( \19519 , \13049 , RIbe2ab68_104);
and \U$19267 ( \19520 , \13669 , RIbe2aaf0_103);
nor \U$19268 ( \19521 , \19519 , \19520 );
not \U$19269 ( \19522 , \19521 );
or \U$19270 ( \19523 , \19518 , \19522 );
or \U$19271 ( \19524 , \19521 , \12195 );
nand \U$19272 ( \19525 , \19523 , \19524 );
not \U$19273 ( \19526 , \19525 );
not \U$19274 ( \19527 , RIbe2a280_85);
nor \U$19275 ( \19528 , \19527 , \12810 );
and \U$19276 ( \19529 , RIbe2a208_84, RIbe2ae38_110);
nor \U$19277 ( \19530 , \19528 , \19529 );
xnor \U$19278 ( \19531 , \19530 , RIbe2aeb0_111);
not \U$19279 ( \19532 , \19531 );
nand \U$19280 ( \19533 , \19532 , \12956 );
not \U$19281 ( \19534 , \19533 );
not \U$19282 ( \19535 , \12893 );
not \U$19283 ( \19536 , RIbe2b108_116);
not \U$19284 ( \19537 , \15250 );
or \U$19285 ( \19538 , \19536 , \19537 );
nand \U$19286 ( \19539 , \12890 , RIbe2b090_115);
nand \U$19287 ( \19540 , \19538 , \19539 );
not \U$19288 ( \19541 , \19540 );
or \U$19289 ( \19542 , \19535 , \19541 );
or \U$19290 ( \19543 , \19540 , \12801 );
nand \U$19291 ( \19544 , \19542 , \19543 );
not \U$19292 ( \19545 , \19544 );
or \U$19293 ( \19546 , \19534 , \19545 );
nand \U$19294 ( \19547 , \19531 , \12195 );
nand \U$19295 ( \19548 , \19546 , \19547 );
not \U$19296 ( \19549 , \19548 );
or \U$19297 ( \19550 , \19526 , \19549 );
not \U$19298 ( \19551 , RIbe2b180_117);
not \U$19299 ( \19552 , \13010 );
or \U$19300 ( \19553 , \19551 , \19552 );
nand \U$19301 ( \19554 , \13012 , RIbe2b270_119);
nand \U$19302 ( \19555 , \19553 , \19554 );
and \U$19303 ( \19556 , \19555 , \13595 );
not \U$19304 ( \19557 , \19555 );
and \U$19305 ( \19558 , \19557 , \12823 );
nor \U$19306 ( \19559 , \19556 , \19558 );
not \U$19307 ( \19560 , \19559 );
not \U$19308 ( \19561 , RIbe2b018_114);
not \U$19309 ( \19562 , \13063 );
or \U$19310 ( \19563 , \19561 , \19562 );
nand \U$19311 ( \19564 , \13728 , RIbe2afa0_113);
nand \U$19312 ( \19565 , \19563 , \19564 );
and \U$19313 ( \19566 , \19565 , \13068 );
not \U$19314 ( \19567 , \19565 );
and \U$19315 ( \19568 , \19567 , \12723 );
nor \U$19316 ( \19569 , \19566 , \19568 );
not \U$19317 ( \19570 , \19569 );
or \U$19318 ( \19571 , \19560 , \19570 );
or \U$19319 ( \19572 , \19569 , \19559 );
not \U$19320 ( \19573 , RIbe2af28_112);
not \U$19321 ( \19574 , \14071 );
or \U$19322 ( \19575 , \19573 , \19574 );
nand \U$19323 ( \19576 , RIbe2b1f8_118, \14074 );
nand \U$19324 ( \19577 , \19575 , \19576 );
and \U$19325 ( \19578 , \19577 , \12746 );
not \U$19326 ( \19579 , \19577 );
and \U$19327 ( \19580 , \19579 , \12743 );
nor \U$19328 ( \19581 , \19578 , \19580 );
not \U$19329 ( \19582 , \19581 );
nand \U$19330 ( \19583 , \19572 , \19582 );
nand \U$19331 ( \19584 , \19571 , \19583 );
not \U$19332 ( \19585 , \19525 );
not \U$19333 ( \19586 , \19548 );
nand \U$19334 ( \19587 , \19585 , \19586 );
nand \U$19335 ( \19588 , \19584 , \19587 );
nand \U$19336 ( \19589 , \19550 , \19588 );
not \U$19337 ( \19590 , \19206 );
not \U$19338 ( \19591 , \19212 );
or \U$19339 ( \19592 , \19590 , \19591 );
or \U$19340 ( \19593 , \19212 , \19206 );
nand \U$19341 ( \19594 , \19592 , \19593 );
xor \U$19342 ( \19595 , \19589 , \19594 );
xor \U$19343 ( \19596 , \19248 , \19285 );
xor \U$19344 ( \19597 , \19596 , \19288 );
and \U$19345 ( \19598 , \19595 , \19597 );
and \U$19346 ( \19599 , \19589 , \19594 );
or \U$19347 ( \19600 , \19598 , \19599 );
not \U$19348 ( \19601 , \19600 );
not \U$19349 ( \19602 , \19131 );
not \U$19350 ( \19603 , \19163 );
and \U$19351 ( \19604 , \19602 , \19603 );
and \U$19352 ( \19605 , \19131 , \19163 );
nor \U$19353 ( \19606 , \19604 , \19605 );
xor \U$19354 ( \19607 , \19606 , \19167 );
or \U$19355 ( \19608 , \19601 , \19607 );
not \U$19356 ( \19609 , \19607 );
not \U$19357 ( \19610 , \19601 );
or \U$19358 ( \19611 , \19609 , \19610 );
xor \U$19359 ( \19612 , \19213 , \19291 );
xnor \U$19360 ( \19613 , \19612 , \19204 );
not \U$19361 ( \19614 , \19613 );
nand \U$19362 ( \19615 , \19611 , \19614 );
nand \U$19363 ( \19616 , \19608 , \19615 );
xnor \U$19364 ( \19617 , \19295 , \19201 );
not \U$19365 ( \19618 , \19617 );
not \U$19366 ( \19619 , \19300 );
and \U$19367 ( \19620 , \19618 , \19619 );
and \U$19368 ( \19621 , \19617 , \19300 );
nor \U$19369 ( \19622 , \19620 , \19621 );
xnor \U$19370 ( \19623 , \19616 , \19622 );
not \U$19371 ( \19624 , \19623 );
not \U$19372 ( \19625 , RIbe2af28_112);
not \U$19373 ( \19626 , \12858 );
or \U$19374 ( \19627 , \19625 , \19626 );
nand \U$19375 ( \19628 , \12834 , RIbe2b1f8_118);
nand \U$19376 ( \19629 , \19627 , \19628 );
and \U$19377 ( \19630 , \19629 , \14815 );
not \U$19378 ( \19631 , \19629 );
and \U$19379 ( \19632 , \19631 , \13595 );
nor \U$19380 ( \19633 , \19630 , \19632 );
not \U$19381 ( \19634 , RIbe2aaf0_103);
not \U$19382 ( \19635 , \14523 );
or \U$19383 ( \19636 , \19634 , \19635 );
nand \U$19384 ( \19637 , \13728 , RIbe2b630_127);
nand \U$19385 ( \19638 , \19636 , \19637 );
and \U$19386 ( \19639 , \19638 , \13583 );
not \U$19387 ( \19640 , \19638 );
and \U$19388 ( \19641 , \19640 , \13068 );
nor \U$19389 ( \19642 , \19639 , \19641 );
nand \U$19390 ( \19643 , \19633 , \19642 );
not \U$19391 ( \19644 , RIbe2b018_114);
not \U$19392 ( \19645 , \12847 );
or \U$19393 ( \19646 , \19644 , \19645 );
nand \U$19394 ( \19647 , \12735 , RIbe2afa0_113);
nand \U$19395 ( \19648 , \19646 , \19647 );
and \U$19396 ( \19649 , \19648 , \12852 );
not \U$19397 ( \19650 , \19648 );
and \U$19398 ( \19651 , \19650 , \12746 );
nor \U$19399 ( \19652 , \19649 , \19651 );
nand \U$19400 ( \19653 , \19643 , \19652 );
or \U$19401 ( \19654 , \19633 , \19642 );
and \U$19402 ( \19655 , \19653 , \19654 );
not \U$19403 ( \19656 , RIbe2b108_116);
not \U$19404 ( \19657 , \13690 );
or \U$19405 ( \19658 , \19656 , \19657 );
nand \U$19406 ( \19659 , RIbe2b090_115, RIbe2ae38_110);
nand \U$19407 ( \19660 , \19658 , \19659 );
xnor \U$19408 ( \19661 , \19660 , RIbe2aeb0_111);
xor \U$19409 ( \19662 , \12924 , \19661 );
not \U$19410 ( \19663 , RIbe2b180_117);
not \U$19411 ( \19664 , \13518 );
or \U$19412 ( \19665 , \19663 , \19664 );
nand \U$19413 ( \19666 , \12890 , RIbe2b270_119);
nand \U$19414 ( \19667 , \19665 , \19666 );
and \U$19415 ( \19668 , \19667 , \12998 );
not \U$19416 ( \19669 , \19667 );
and \U$19417 ( \19670 , \19669 , \16334 );
nor \U$19418 ( \19671 , \19668 , \19670 );
and \U$19419 ( \19672 , \19662 , \19671 );
and \U$19420 ( \19673 , \12924 , \19661 );
or \U$19421 ( \19674 , \19672 , \19673 );
nand \U$19422 ( \19675 , \19655 , \19674 );
not \U$19423 ( \19676 , \12723 );
not \U$19424 ( \19677 , RIbe2b630_127);
not \U$19425 ( \19678 , \12707 );
or \U$19426 ( \19679 , \19677 , \19678 );
nand \U$19427 ( \19680 , \12711 , RIbe2b018_114);
nand \U$19428 ( \19681 , \19679 , \19680 );
not \U$19429 ( \19682 , \19681 );
or \U$19430 ( \19683 , \19676 , \19682 );
or \U$19431 ( \19684 , \19681 , \12723 );
nand \U$19432 ( \19685 , \19683 , \19684 );
not \U$19433 ( \19686 , RIbe2afa0_113);
not \U$19434 ( \19687 , \12847 );
or \U$19435 ( \19688 , \19686 , \19687 );
nand \U$19436 ( \19689 , \13077 , RIbe2af28_112);
nand \U$19437 ( \19690 , \19688 , \19689 );
and \U$19438 ( \19691 , \19690 , \12852 );
not \U$19439 ( \19692 , \19690 );
and \U$19440 ( \19693 , \19692 , \12742 );
nor \U$19441 ( \19694 , \19691 , \19693 );
xor \U$19442 ( \19695 , \19685 , \19694 );
not \U$19443 ( \19696 , \12751 );
not \U$19444 ( \19697 , \13192 );
and \U$19445 ( \19698 , \19696 , \19697 );
and \U$19446 ( \19699 , \15615 , RIbe2ab68_104);
nor \U$19447 ( \19700 , \19698 , \19699 );
and \U$19448 ( \19701 , \19700 , \12924 );
not \U$19449 ( \19702 , \19700 );
and \U$19450 ( \19703 , \19702 , \12774 );
nor \U$19451 ( \19704 , \19701 , \19703 );
xor \U$19452 ( \19705 , \19695 , \19704 );
and \U$19453 ( \19706 , \19675 , \19705 );
nor \U$19454 ( \19707 , \19655 , \19674 );
nor \U$19455 ( \19708 , \19706 , \19707 );
not \U$19456 ( \19709 , \19708 );
not \U$19457 ( \19710 , \19709 );
nand \U$19458 ( \19711 , \13669 , RIbe2ab68_104);
and \U$19459 ( \19712 , \19711 , \12195 );
not \U$19460 ( \19713 , \19711 );
and \U$19461 ( \19714 , \19713 , \12960 );
nor \U$19462 ( \19715 , \19712 , \19714 );
not \U$19463 ( \19716 , \19715 );
nor \U$19464 ( \19717 , \19531 , \17005 );
not \U$19465 ( \19718 , \19717 );
nand \U$19466 ( \19719 , \19531 , \12960 );
nand \U$19467 ( \19720 , \19718 , \19719 );
xor \U$19468 ( \19721 , \19720 , \19544 );
not \U$19469 ( \19722 , \19721 );
or \U$19470 ( \19723 , \19716 , \19722 );
or \U$19471 ( \19724 , \19721 , \19715 );
nand \U$19472 ( \19725 , \19723 , \19724 );
not \U$19473 ( \19726 , \19725 );
not \U$19474 ( \19727 , \19559 );
not \U$19475 ( \19728 , \19727 );
not \U$19476 ( \19729 , \19582 );
or \U$19477 ( \19730 , \19728 , \19729 );
nand \U$19478 ( \19731 , \19581 , \19559 );
nand \U$19479 ( \19732 , \19730 , \19731 );
not \U$19480 ( \19733 , \19569 );
and \U$19481 ( \19734 , \19732 , \19733 );
not \U$19482 ( \19735 , \19732 );
and \U$19483 ( \19736 , \19735 , \19569 );
nor \U$19484 ( \19737 , \19734 , \19736 );
not \U$19485 ( \19738 , \19737 );
and \U$19486 ( \19739 , \19726 , \19738 );
and \U$19487 ( \19740 , \19737 , \19725 );
nor \U$19488 ( \19741 , \19739 , \19740 );
not \U$19489 ( \19742 , \19741 );
not \U$19490 ( \19743 , \19742 );
or \U$19491 ( \19744 , \19710 , \19743 );
not \U$19492 ( \19745 , \19741 );
not \U$19493 ( \19746 , \19708 );
or \U$19494 ( \19747 , \19745 , \19746 );
and \U$19495 ( \19748 , \13738 , RIbe2aaf0_103);
not \U$19496 ( \19749 , \12751 );
and \U$19497 ( \19750 , \19749 , RIbe2b630_127);
nor \U$19498 ( \19751 , \19748 , \19750 );
and \U$19499 ( \19752 , \19751 , \12924 );
not \U$19500 ( \19753 , \19751 );
and \U$19501 ( \19754 , \19753 , \12927 );
nor \U$19502 ( \19755 , \19752 , \19754 );
xor \U$19503 ( \19756 , \19685 , \19694 );
and \U$19504 ( \19757 , \19756 , \19704 );
and \U$19505 ( \19758 , \19685 , \19694 );
or \U$19506 ( \19759 , \19757 , \19758 );
xor \U$19507 ( \19760 , \19755 , \19759 );
not \U$19508 ( \19761 , RIbe2b090_115);
not \U$19509 ( \19762 , \13004 );
or \U$19510 ( \19763 , \19761 , \19762 );
nand \U$19511 ( \19764 , RIbe2a280_85, RIbe2ae38_110);
nand \U$19512 ( \19765 , \19763 , \19764 );
xor \U$19513 ( \19766 , \19765 , RIbe2aeb0_111);
not \U$19514 ( \19767 , \12801 );
not \U$19515 ( \19768 , RIbe2b270_119);
not \U$19516 ( \19769 , \12887 );
or \U$19517 ( \19770 , \19768 , \19769 );
nand \U$19518 ( \19771 , \12890 , RIbe2b108_116);
nand \U$19519 ( \19772 , \19770 , \19771 );
not \U$19520 ( \19773 , \19772 );
or \U$19521 ( \19774 , \19767 , \19773 );
or \U$19522 ( \19775 , \19772 , \12801 );
nand \U$19523 ( \19776 , \19774 , \19775 );
xor \U$19524 ( \19777 , \19766 , \19776 );
not \U$19525 ( \19778 , RIbe2b1f8_118);
nor \U$19526 ( \19779 , \19778 , \18607 );
not \U$19527 ( \19780 , \13012 );
nor \U$19528 ( \19781 , \19780 , \14248 );
nor \U$19529 ( \19782 , \19779 , \19781 );
not \U$19530 ( \19783 , \13705 );
and \U$19531 ( \19784 , \19782 , \19783 );
not \U$19532 ( \19785 , \19782 );
and \U$19533 ( \19786 , \19785 , \13705 );
nor \U$19534 ( \19787 , \19784 , \19786 );
and \U$19535 ( \19788 , \19777 , \19787 );
and \U$19536 ( \19789 , \19766 , \19776 );
or \U$19537 ( \19790 , \19788 , \19789 );
xor \U$19538 ( \19791 , \19760 , \19790 );
nand \U$19539 ( \19792 , \19747 , \19791 );
nand \U$19540 ( \19793 , \19744 , \19792 );
not \U$19541 ( \19794 , \19793 );
not \U$19542 ( \19795 , \19525 );
not \U$19543 ( \19796 , \19586 );
or \U$19544 ( \19797 , \19795 , \19796 );
or \U$19545 ( \19798 , \19586 , \19525 );
nand \U$19546 ( \19799 , \19797 , \19798 );
xnor \U$19547 ( \19800 , \19584 , \19799 );
and \U$19548 ( \19801 , \19221 , \19231 );
not \U$19549 ( \19802 , \19221 );
and \U$19550 ( \19803 , \19802 , \19246 );
nor \U$19551 ( \19804 , \19801 , \19803 );
xor \U$19552 ( \19805 , \19243 , \19804 );
nand \U$19553 ( \19806 , \19800 , \19805 );
not \U$19554 ( \19807 , \19806 );
nor \U$19555 ( \19808 , \19800 , \19805 );
nor \U$19556 ( \19809 , \19807 , \19808 );
not \U$19557 ( \19810 , \19809 );
or \U$19558 ( \19811 , \19794 , \19810 );
or \U$19559 ( \19812 , \19793 , \19809 );
nand \U$19560 ( \19813 , \19811 , \19812 );
not \U$19561 ( \19814 , \19813 );
not \U$19562 ( \19815 , \19259 );
not \U$19563 ( \19816 , \19270 );
or \U$19564 ( \19817 , \19815 , \19816 );
nand \U$19565 ( \19818 , \19258 , \19271 );
nand \U$19566 ( \19819 , \19817 , \19818 );
xor \U$19567 ( \19820 , \19819 , \19283 );
not \U$19568 ( \19821 , \19715 );
not \U$19569 ( \19822 , \19821 );
not \U$19570 ( \19823 , \19721 );
or \U$19571 ( \19824 , \19822 , \19823 );
not \U$19572 ( \19825 , \19737 );
or \U$19573 ( \19826 , \19721 , \19821 );
nand \U$19574 ( \19827 , \19825 , \19826 );
nand \U$19575 ( \19828 , \19824 , \19827 );
xor \U$19576 ( \19829 , \19820 , \19828 );
xor \U$19577 ( \19830 , \19755 , \19759 );
and \U$19578 ( \19831 , \19830 , \19790 );
and \U$19579 ( \19832 , \19755 , \19759 );
or \U$19580 ( \19833 , \19831 , \19832 );
xor \U$19581 ( \19834 , \19829 , \19833 );
not \U$19582 ( \19835 , \19834 );
not \U$19583 ( \19836 , \19835 );
and \U$19584 ( \19837 , \19814 , \19836 );
and \U$19585 ( \19838 , \19813 , \19835 );
nor \U$19586 ( \19839 , \19837 , \19838 );
not \U$19587 ( \19840 , \19839 );
xor \U$19588 ( \19841 , \19766 , \19776 );
xor \U$19589 ( \19842 , \19841 , \19787 );
nand \U$19590 ( \19843 , \19749 , RIbe2ab68_104);
and \U$19591 ( \19844 , \19843 , \12924 );
not \U$19592 ( \19845 , \19843 );
and \U$19593 ( \19846 , \19845 , \12927 );
nor \U$19594 ( \19847 , \19844 , \19846 );
not \U$19595 ( \19848 , RIbe2b270_119);
not \U$19596 ( \19849 , \12811 );
or \U$19597 ( \19850 , \19848 , \19849 );
nand \U$19598 ( \19851 , RIbe2b108_116, RIbe2ae38_110);
nand \U$19599 ( \19852 , \19850 , \19851 );
xor \U$19600 ( \19853 , \19852 , RIbe2aeb0_111);
not \U$19601 ( \19854 , RIbe2b1f8_118);
not \U$19602 ( \19855 , \13518 );
or \U$19603 ( \19856 , \19854 , \19855 );
not \U$19604 ( \19857 , \14248 );
nand \U$19605 ( \19858 , \19857 , \12794 );
nand \U$19606 ( \19859 , \19856 , \19858 );
and \U$19607 ( \19860 , \19859 , \16334 );
not \U$19608 ( \19861 , \19859 );
and \U$19609 ( \19862 , \19861 , \12893 );
nor \U$19610 ( \19863 , \19860 , \19862 );
xor \U$19611 ( \19864 , \19853 , \19863 );
not \U$19612 ( \19865 , RIbe2afa0_113);
not \U$19613 ( \19866 , \12831 );
or \U$19614 ( \19867 , \19865 , \19866 );
nand \U$19615 ( \19868 , \13012 , RIbe2af28_112);
nand \U$19616 ( \19869 , \19867 , \19868 );
and \U$19617 ( \19870 , \19869 , \14555 );
not \U$19618 ( \19871 , \19869 );
and \U$19619 ( \19872 , \19871 , \12863 );
nor \U$19620 ( \19873 , \19870 , \19872 );
and \U$19621 ( \19874 , \19864 , \19873 );
and \U$19622 ( \19875 , \19853 , \19863 );
or \U$19623 ( \19876 , \19874 , \19875 );
xor \U$19624 ( \19877 , \19847 , \19876 );
not \U$19625 ( \19878 , \19642 );
not \U$19626 ( \19879 , \19633 );
not \U$19627 ( \19880 , \19652 );
or \U$19628 ( \19881 , \19879 , \19880 );
or \U$19629 ( \19882 , \19652 , \19633 );
nand \U$19630 ( \19883 , \19881 , \19882 );
not \U$19631 ( \19884 , \19883 );
or \U$19632 ( \19885 , \19878 , \19884 );
or \U$19633 ( \19886 , \19642 , \19883 );
nand \U$19634 ( \19887 , \19885 , \19886 );
and \U$19635 ( \19888 , \19877 , \19887 );
and \U$19636 ( \19889 , \19847 , \19876 );
or \U$19637 ( \19890 , \19888 , \19889 );
xor \U$19638 ( \19891 , \19842 , \19890 );
xor \U$19639 ( \19892 , \19674 , \19655 );
xor \U$19640 ( \19893 , \19892 , \19705 );
and \U$19641 ( \19894 , \19891 , \19893 );
and \U$19642 ( \19895 , \19842 , \19890 );
or \U$19643 ( \19896 , \19894 , \19895 );
and \U$19644 ( \19897 , \19742 , \19708 );
not \U$19645 ( \19898 , \19742 );
and \U$19646 ( \19899 , \19898 , \19709 );
nor \U$19647 ( \19900 , \19897 , \19899 );
not \U$19648 ( \19901 , \19791 );
and \U$19649 ( \19902 , \19900 , \19901 );
not \U$19650 ( \19903 , \19900 );
and \U$19651 ( \19904 , \19903 , \19791 );
nor \U$19652 ( \19905 , \19902 , \19904 );
and \U$19653 ( \19906 , \19896 , \19905 );
not \U$19654 ( \19907 , \19906 );
and \U$19655 ( \19908 , \19840 , \19907 );
and \U$19656 ( \19909 , \19839 , \19906 );
nor \U$19657 ( \19910 , \19908 , \19909 );
not \U$19658 ( \19911 , \19910 );
not \U$19659 ( \19912 , \16382 );
not \U$19660 ( \19913 , \15873 );
and \U$19661 ( \19914 , \19912 , \19913 );
nor \U$19662 ( \19915 , \17741 , \13192 );
nor \U$19663 ( \19916 , \19914 , \19915 );
and \U$19664 ( \19917 , \19916 , \13068 );
not \U$19665 ( \19918 , \19916 );
and \U$19666 ( \19919 , \19918 , \13583 );
nor \U$19667 ( \19920 , \19917 , \19919 );
not \U$19668 ( \19921 , \19920 );
xor \U$19669 ( \19922 , \19853 , \19863 );
xor \U$19670 ( \19923 , \19922 , \19873 );
nand \U$19671 ( \19924 , \19921 , \19923 );
xor \U$19672 ( \19925 , \12924 , \19661 );
xor \U$19673 ( \19926 , \19925 , \19671 );
xor \U$19674 ( \19927 , \19924 , \19926 );
not \U$19675 ( \19928 , RIbe2b180_117);
not \U$19676 ( \19929 , \13003 );
or \U$19677 ( \19930 , \19928 , \19929 );
nand \U$19678 ( \19931 , RIbe2b270_119, RIbe2ae38_110);
nand \U$19679 ( \19932 , \19930 , \19931 );
xor \U$19680 ( \19933 , \19932 , RIbe2aeb0_111);
not \U$19681 ( \19934 , \19933 );
nand \U$19682 ( \19935 , \19934 , \13583 );
not \U$19683 ( \19936 , \19935 );
not \U$19684 ( \19937 , RIbe2af28_112);
not \U$19685 ( \19938 , \13518 );
or \U$19686 ( \19939 , \19937 , \19938 );
nand \U$19687 ( \19940 , \12890 , RIbe2b1f8_118);
nand \U$19688 ( \19941 , \19939 , \19940 );
and \U$19689 ( \19942 , \19941 , \12804 );
not \U$19690 ( \19943 , \19941 );
and \U$19691 ( \19944 , \19943 , \12998 );
nor \U$19692 ( \19945 , \19942 , \19944 );
not \U$19693 ( \19946 , \19945 );
or \U$19694 ( \19947 , \19936 , \19946 );
nand \U$19695 ( \19948 , \19933 , \13068 );
nand \U$19696 ( \19949 , \19947 , \19948 );
not \U$19697 ( \19950 , \19949 );
not \U$19698 ( \19951 , \19950 );
and \U$19699 ( \19952 , \14074 , RIbe2b018_114);
and \U$19700 ( \19953 , \12847 , RIbe2b630_127);
nor \U$19701 ( \19954 , \19952 , \19953 );
and \U$19702 ( \19955 , \19954 , \12743 );
not \U$19703 ( \19956 , \19954 );
and \U$19704 ( \19957 , \19956 , \12742 );
nor \U$19705 ( \19958 , \19955 , \19957 );
not \U$19706 ( \19959 , \19958 );
and \U$19707 ( \19960 , \19951 , \19959 );
nand \U$19708 ( \19961 , \12711 , RIbe2ab68_104);
and \U$19709 ( \19962 , \19961 , \12723 );
not \U$19710 ( \19963 , \19961 );
and \U$19711 ( \19964 , \19963 , \13068 );
nor \U$19712 ( \19965 , \19962 , \19964 );
not \U$19713 ( \19966 , RIbe2aaf0_103);
not \U$19714 ( \19967 , \12847 );
or \U$19715 ( \19968 , \19966 , \19967 );
nand \U$19716 ( \19969 , \14074 , RIbe2b630_127);
nand \U$19717 ( \19970 , \19968 , \19969 );
and \U$19718 ( \19971 , \19970 , \12743 );
not \U$19719 ( \19972 , \19970 );
and \U$19720 ( \19973 , \19972 , \12742 );
nor \U$19721 ( \19974 , \19971 , \19973 );
xor \U$19722 ( \19975 , \19965 , \19974 );
not \U$19723 ( \19976 , RIbe2b018_114);
nor \U$19724 ( \19977 , \19976 , \12830 );
not \U$19725 ( \19978 , RIbe2afa0_113);
not \U$19726 ( \19979 , \12835 );
nor \U$19727 ( \19980 , \19978 , \19979 );
nor \U$19728 ( \19981 , \19977 , \19980 );
and \U$19729 ( \19982 , \19981 , \15263 );
not \U$19730 ( \19983 , \19981 );
and \U$19731 ( \19984 , \19983 , \13595 );
nor \U$19732 ( \19985 , \19982 , \19984 );
and \U$19733 ( \19986 , \19975 , \19985 );
and \U$19734 ( \19987 , \19965 , \19974 );
or \U$19735 ( \19988 , \19986 , \19987 );
nand \U$19736 ( \19989 , \19950 , \19958 );
and \U$19737 ( \19990 , \19988 , \19989 );
nor \U$19738 ( \19991 , \19960 , \19990 );
and \U$19739 ( \19992 , \19927 , \19991 );
and \U$19740 ( \19993 , \19924 , \19926 );
or \U$19741 ( \19994 , \19992 , \19993 );
not \U$19742 ( \19995 , \19994 );
xor \U$19743 ( \19996 , \19842 , \19890 );
xor \U$19744 ( \19997 , \19996 , \19893 );
nand \U$19745 ( \19998 , \19995 , \19997 );
not \U$19746 ( \19999 , \19998 );
not \U$19747 ( \20000 , \19999 );
xor \U$19748 ( \20001 , \19896 , \19905 );
not \U$19749 ( \20002 , \20001 );
not \U$19750 ( \20003 , \20002 );
or \U$19751 ( \20004 , \20000 , \20003 );
nand \U$19752 ( \20005 , \20001 , \19998 );
nand \U$19753 ( \20006 , \20004 , \20005 );
xor \U$19754 ( \20007 , \19847 , \19876 );
xor \U$19755 ( \20008 , \20007 , \19887 );
not \U$19756 ( \20009 , \20008 );
xor \U$19757 ( \20010 , \19924 , \19926 );
xor \U$19758 ( \20011 , \20010 , \19991 );
nor \U$19759 ( \20012 , \20009 , \20011 );
not \U$19760 ( \20013 , \19994 );
not \U$19761 ( \20014 , \19997 );
or \U$19762 ( \20015 , \20013 , \20014 );
or \U$19763 ( \20016 , \19997 , \19994 );
nand \U$19764 ( \20017 , \20015 , \20016 );
xor \U$19765 ( \20018 , \20012 , \20017 );
and \U$19766 ( \20019 , \19911 , \20006 , \20018 );
xor \U$19767 ( \20020 , \19607 , \19600 );
xnor \U$19768 ( \20021 , \20020 , \19613 );
xor \U$19769 ( \20022 , \19820 , \19828 );
and \U$19770 ( \20023 , \20022 , \19833 );
and \U$19771 ( \20024 , \19820 , \19828 );
or \U$19772 ( \20025 , \20023 , \20024 );
not \U$19773 ( \20026 , \19805 );
nor \U$19774 ( \20027 , \20026 , \19800 );
or \U$19775 ( \20028 , \20025 , \20027 );
xor \U$19776 ( \20029 , \19589 , \19594 );
xor \U$19777 ( \20030 , \20029 , \19597 );
and \U$19778 ( \20031 , \20028 , \20030 );
and \U$19779 ( \20032 , \20025 , \20027 );
nor \U$19780 ( \20033 , \20031 , \20032 );
xor \U$19781 ( \20034 , \20021 , \20033 );
not \U$19782 ( \20035 , \19793 );
or \U$19783 ( \20036 , \20035 , \19809 );
not \U$19784 ( \20037 , \19809 );
not \U$19785 ( \20038 , \20035 );
or \U$19786 ( \20039 , \20037 , \20038 );
nand \U$19787 ( \20040 , \20039 , \19834 );
nand \U$19788 ( \20041 , \20036 , \20040 );
not \U$19789 ( \20042 , \20041 );
xor \U$19790 ( \20043 , \20025 , \20027 );
xor \U$19791 ( \20044 , \20043 , \20030 );
not \U$19792 ( \20045 , \20044 );
not \U$19793 ( \20046 , \20045 );
or \U$19794 ( \20047 , \20042 , \20046 );
not \U$19795 ( \20048 , \20041 );
nand \U$19796 ( \20049 , \20048 , \20044 );
nand \U$19797 ( \20050 , \20047 , \20049 );
and \U$19798 ( \20051 , \20019 , \20034 , \20050 );
not \U$19799 ( \20052 , \20051 );
not \U$19800 ( \20053 , \20008 );
not \U$19801 ( \20054 , \20011 );
or \U$19802 ( \20055 , \20053 , \20054 );
or \U$19803 ( \20056 , \20011 , \20008 );
nand \U$19804 ( \20057 , \20055 , \20056 );
not \U$19805 ( \20058 , \20057 );
and \U$19806 ( \20059 , \13068 , \19934 );
not \U$19807 ( \20060 , \13068 );
and \U$19808 ( \20061 , \20060 , \19933 );
nor \U$19809 ( \20062 , \20059 , \20061 );
not \U$19810 ( \20063 , \20062 );
not \U$19811 ( \20064 , \19945 );
or \U$19812 ( \20065 , \20063 , \20064 );
or \U$19813 ( \20066 , \20062 , \19945 );
nand \U$19814 ( \20067 , \20065 , \20066 );
not \U$19815 ( \20068 , RIbe2b1f8_118);
not \U$19816 ( \20069 , \13004 );
or \U$19817 ( \20070 , \20068 , \20069 );
nand \U$19818 ( \20071 , RIbe2b180_117, RIbe2ae38_110);
nand \U$19819 ( \20072 , \20070 , \20071 );
xor \U$19820 ( \20073 , \20072 , RIbe2aeb0_111);
not \U$19821 ( \20074 , RIbe2afa0_113);
not \U$19822 ( \20075 , \13518 );
or \U$19823 ( \20076 , \20074 , \20075 );
nand \U$19824 ( \20077 , \12890 , RIbe2af28_112);
nand \U$19825 ( \20078 , \20076 , \20077 );
and \U$19826 ( \20079 , \20078 , \14103 );
not \U$19827 ( \20080 , \20078 );
and \U$19828 ( \20081 , \20080 , \12893 );
nor \U$19829 ( \20082 , \20079 , \20081 );
xor \U$19830 ( \20083 , \20073 , \20082 );
not \U$19831 ( \20084 , RIbe2b630_127);
nor \U$19832 ( \20085 , \20084 , \12830 );
not \U$19833 ( \20086 , RIbe2b018_114);
nor \U$19834 ( \20087 , \20086 , \19979 );
nor \U$19835 ( \20088 , \20085 , \20087 );
and \U$19836 ( \20089 , \20088 , \19783 );
not \U$19837 ( \20090 , \20088 );
and \U$19838 ( \20091 , \20090 , \13595 );
nor \U$19839 ( \20092 , \20089 , \20091 );
and \U$19840 ( \20093 , \20083 , \20092 );
and \U$19841 ( \20094 , \20073 , \20082 );
or \U$19842 ( \20095 , \20093 , \20094 );
xor \U$19843 ( \20096 , \20067 , \20095 );
xor \U$19844 ( \20097 , \19965 , \19974 );
xor \U$19845 ( \20098 , \20097 , \19985 );
and \U$19846 ( \20099 , \20096 , \20098 );
and \U$19847 ( \20100 , \20067 , \20095 );
or \U$19848 ( \20101 , \20099 , \20100 );
not \U$19849 ( \20102 , \19920 );
not \U$19850 ( \20103 , \19923 );
or \U$19851 ( \20104 , \20102 , \20103 );
or \U$19852 ( \20105 , \19923 , \19920 );
nand \U$19853 ( \20106 , \20104 , \20105 );
xor \U$19854 ( \20107 , \20101 , \20106 );
not \U$19855 ( \20108 , \19988 );
not \U$19856 ( \20109 , \19958 );
not \U$19857 ( \20110 , \19949 );
and \U$19858 ( \20111 , \20109 , \20110 );
and \U$19859 ( \20112 , \19949 , \19958 );
nor \U$19860 ( \20113 , \20111 , \20112 );
not \U$19861 ( \20114 , \20113 );
or \U$19862 ( \20115 , \20108 , \20114 );
or \U$19863 ( \20116 , \20113 , \19988 );
nand \U$19864 ( \20117 , \20115 , \20116 );
and \U$19865 ( \20118 , \20107 , \20117 );
and \U$19866 ( \20119 , \20101 , \20106 );
or \U$19867 ( \20120 , \20118 , \20119 );
not \U$19868 ( \20121 , \20120 );
or \U$19869 ( \20122 , \20058 , \20121 );
and \U$19870 ( \20123 , \12847 , RIbe2ab68_104);
and \U$19871 ( \20124 , \14074 , RIbe2aaf0_103);
nor \U$19872 ( \20125 , \20123 , \20124 );
and \U$19873 ( \20126 , \20125 , \12742 );
not \U$19874 ( \20127 , \20125 );
and \U$19875 ( \20128 , \20127 , \12743 );
nor \U$19876 ( \20129 , \20126 , \20128 );
not \U$19877 ( \20130 , RIbe2aaf0_103);
not \U$19878 ( \20131 , \13010 );
or \U$19879 ( \20132 , \20130 , \20131 );
nand \U$19880 ( \20133 , \12835 , RIbe2b630_127);
nand \U$19881 ( \20134 , \20132 , \20133 );
and \U$19882 ( \20135 , \20134 , \14555 );
not \U$19883 ( \20136 , \20134 );
and \U$19884 ( \20137 , \20136 , \14558 );
nor \U$19885 ( \20138 , \20135 , \20137 );
nand \U$19886 ( \20139 , \14074 , RIbe2ab68_104);
and \U$19887 ( \20140 , \20139 , \12746 );
not \U$19888 ( \20141 , \20139 );
and \U$19889 ( \20142 , \20141 , \14358 );
nor \U$19890 ( \20143 , \20140 , \20142 );
and \U$19891 ( \20144 , \20138 , \20143 );
xor \U$19892 ( \20145 , \20129 , \20144 );
not \U$19893 ( \20146 , \12743 );
not \U$19894 ( \20147 , RIbe2af28_112);
not \U$19895 ( \20148 , \12811 );
or \U$19896 ( \20149 , \20147 , \20148 );
nand \U$19897 ( \20150 , RIbe2b1f8_118, RIbe2ae38_110);
nand \U$19898 ( \20151 , \20149 , \20150 );
xor \U$19899 ( \20152 , \20151 , RIbe2aeb0_111);
not \U$19900 ( \20153 , \20152 );
or \U$19901 ( \20154 , \20146 , \20153 );
or \U$19902 ( \20155 , \20152 , \12743 );
not \U$19903 ( \20156 , RIbe2b018_114);
not \U$19904 ( \20157 , \12887 );
or \U$19905 ( \20158 , \20156 , \20157 );
nand \U$19906 ( \20159 , \12890 , RIbe2afa0_113);
nand \U$19907 ( \20160 , \20158 , \20159 );
xnor \U$19908 ( \20161 , \20160 , \12801 );
nand \U$19909 ( \20162 , \20155 , \20161 );
nand \U$19910 ( \20163 , \20154 , \20162 );
and \U$19911 ( \20164 , \20145 , \20163 );
and \U$19912 ( \20165 , \20129 , \20144 );
or \U$19913 ( \20166 , \20164 , \20165 );
xor \U$19914 ( \20167 , \20067 , \20095 );
xor \U$19915 ( \20168 , \20167 , \20098 );
and \U$19916 ( \20169 , \20166 , \20168 );
not \U$19917 ( \20170 , \20169 );
xor \U$19918 ( \20171 , \20101 , \20106 );
xor \U$19919 ( \20172 , \20171 , \20117 );
not \U$19920 ( \20173 , \20172 );
or \U$19921 ( \20174 , \20170 , \20173 );
not \U$19922 ( \20175 , RIbe2b018_114);
not \U$19923 ( \20176 , \13004 );
or \U$19924 ( \20177 , \20175 , \20176 );
nand \U$19925 ( \20178 , RIbe2afa0_113, RIbe2ae38_110);
nand \U$19926 ( \20179 , \20177 , \20178 );
xor \U$19927 ( \20180 , \20179 , RIbe2aeb0_111);
xor \U$19928 ( \20181 , \13595 , \20180 );
and \U$19929 ( \20182 , \12890 , RIbe2b630_127);
and \U$19930 ( \20183 , \12787 , RIbe2aaf0_103);
nor \U$19931 ( \20184 , \20182 , \20183 );
and \U$19932 ( \20185 , \20184 , \12801 );
not \U$19933 ( \20186 , \20184 );
and \U$19934 ( \20187 , \20186 , \14103 );
nor \U$19935 ( \20188 , \20185 , \20187 );
and \U$19936 ( \20189 , \20181 , \20188 );
and \U$19937 ( \20190 , \13595 , \20180 );
or \U$19938 ( \20191 , \20189 , \20190 );
not \U$19939 ( \20192 , RIbe2afa0_113);
not \U$19940 ( \20193 , \13004 );
or \U$19941 ( \20194 , \20192 , \20193 );
nand \U$19942 ( \20195 , RIbe2af28_112, RIbe2ae38_110);
nand \U$19943 ( \20196 , \20194 , \20195 );
xor \U$19944 ( \20197 , RIbe2aeb0_111, \20196 );
not \U$19945 ( \20198 , \12863 );
not \U$19946 ( \20199 , RIbe2ab68_104);
not \U$19947 ( \20200 , \13010 );
or \U$19948 ( \20201 , \20199 , \20200 );
nand \U$19949 ( \20202 , \12835 , RIbe2aaf0_103);
nand \U$19950 ( \20203 , \20201 , \20202 );
not \U$19951 ( \20204 , \20203 );
or \U$19952 ( \20205 , \20198 , \20204 );
or \U$19953 ( \20206 , \20203 , \13706 );
nand \U$19954 ( \20207 , \20205 , \20206 );
xor \U$19955 ( \20208 , \20197 , \20207 );
not \U$19956 ( \20209 , \12998 );
not \U$19957 ( \20210 , RIbe2b630_127);
not \U$19958 ( \20211 , \15250 );
or \U$19959 ( \20212 , \20210 , \20211 );
nand \U$19960 ( \20213 , \12794 , RIbe2b018_114);
nand \U$19961 ( \20214 , \20212 , \20213 );
not \U$19962 ( \20215 , \20214 );
or \U$19963 ( \20216 , \20209 , \20215 );
or \U$19964 ( \20217 , \20214 , \12893 );
nand \U$19965 ( \20218 , \20216 , \20217 );
xor \U$19966 ( \20219 , \20208 , \20218 );
and \U$19967 ( \20220 , \20191 , \20219 );
not \U$19968 ( \20221 , \20220 );
xor \U$19969 ( \20222 , \20143 , \20138 );
xor \U$19970 ( \20223 , \20197 , \20207 );
and \U$19971 ( \20224 , \20223 , \20218 );
and \U$19972 ( \20225 , \20197 , \20207 );
or \U$19973 ( \20226 , \20224 , \20225 );
xor \U$19974 ( \20227 , \20222 , \20226 );
xor \U$19975 ( \20228 , \12743 , \20152 );
xnor \U$19976 ( \20229 , \20228 , \20161 );
not \U$19977 ( \20230 , \20229 );
xor \U$19978 ( \20231 , \20227 , \20230 );
not \U$19979 ( \20232 , \20231 );
or \U$19980 ( \20233 , \20221 , \20232 );
nand \U$19981 ( \20234 , \13012 , RIbe2ab68_104);
and \U$19982 ( \20235 , \20234 , \19783 );
not \U$19983 ( \20236 , \20234 );
and \U$19984 ( \20237 , \20236 , \13705 );
nor \U$19985 ( \20238 , \20235 , \20237 );
xor \U$19986 ( \20239 , \13595 , \20180 );
xor \U$19987 ( \20240 , \20239 , \20188 );
and \U$19988 ( \20241 , \20238 , \20240 );
not \U$19989 ( \20242 , \20241 );
xor \U$19990 ( \20243 , \20191 , \20219 );
not \U$19991 ( \20244 , \20243 );
or \U$19992 ( \20245 , \20242 , \20244 );
not \U$19993 ( \20246 , RIbe2aaf0_103);
not \U$19994 ( \20247 , \13690 );
or \U$19995 ( \20248 , \20246 , \20247 );
nand \U$19996 ( \20249 , RIbe2b630_127, RIbe2ae38_110);
nand \U$19997 ( \20250 , \20248 , \20249 );
xnor \U$19998 ( \20251 , \20250 , RIbe2aeb0_111);
and \U$19999 ( \20252 , \20251 , \12801 );
not \U$20000 ( \20253 , \20251 );
and \U$20001 ( \20254 , \20253 , \14103 );
nor \U$20002 ( \20255 , \20252 , \20254 );
not \U$20003 ( \20256 , \20255 );
nand \U$20004 ( \20257 , \12890 , RIbe2ab68_104);
and \U$20005 ( \20258 , \20257 , \12801 );
not \U$20006 ( \20259 , \20257 );
and \U$20007 ( \20260 , \20259 , \14103 );
or \U$20008 ( \20261 , \20258 , \20260 );
or \U$20009 ( \20262 , \20256 , \20261 );
not \U$20010 ( \20263 , \20261 );
not \U$20011 ( \20264 , \20255 );
or \U$20012 ( \20265 , \20263 , \20264 );
or \U$20013 ( \20266 , \20255 , \20261 );
nand \U$20014 ( \20267 , \20265 , \20266 );
and \U$20015 ( \20268 , \12811 , RIbe2ab68_104);
and \U$20016 ( \20269 , RIbe2aaf0_103, RIbe2ae38_110);
nor \U$20017 ( \20270 , \20268 , \20269 );
xnor \U$20018 ( \20271 , \20270 , RIbe2aeb0_111);
not \U$20019 ( \20272 , RIbe2aeb0_111);
nand \U$20020 ( \20273 , RIbe2ae38_110, RIbe2ab68_104);
not \U$20021 ( \20274 , \20273 );
not \U$20022 ( \20275 , RIbe2aeb0_111);
and \U$20023 ( \20276 , \20274 , \20275 );
and \U$20024 ( \20277 , \20273 , RIbe2aeb0_111);
nor \U$20025 ( \20278 , \20276 , \20277 );
nor \U$20026 ( \20279 , \20272 , \20278 );
nand \U$20027 ( \20280 , \20267 , \20271 , \20279 );
nand \U$20028 ( \20281 , \20262 , \20280 );
not \U$20029 ( \20282 , \20281 );
or \U$20030 ( \20283 , \20251 , \12998 );
not \U$20031 ( \20284 , \20283 );
and \U$20032 ( \20285 , \12811 , RIbe2b630_127);
and \U$20033 ( \20286 , RIbe2b018_114, RIbe2ae38_110);
nor \U$20034 ( \20287 , \20285 , \20286 );
xnor \U$20035 ( \20288 , \20287 , RIbe2aeb0_111);
not \U$20036 ( \20289 , RIbe2ab68_104);
not \U$20037 ( \20290 , \13518 );
or \U$20038 ( \20291 , \20289 , \20290 );
nand \U$20039 ( \20292 , \12890 , RIbe2aaf0_103);
nand \U$20040 ( \20293 , \20291 , \20292 );
and \U$20041 ( \20294 , \20293 , \12995 );
not \U$20042 ( \20295 , \20293 );
and \U$20043 ( \20296 , \20295 , \12998 );
nor \U$20044 ( \20297 , \20294 , \20296 );
xor \U$20045 ( \20298 , \20288 , \20297 );
not \U$20046 ( \20299 , \20298 );
or \U$20047 ( \20300 , \20284 , \20299 );
or \U$20048 ( \20301 , \20298 , \20283 );
nand \U$20049 ( \20302 , \20300 , \20301 );
not \U$20050 ( \20303 , \20302 );
or \U$20051 ( \20304 , \20282 , \20303 );
not \U$20052 ( \20305 , \20298 );
or \U$20053 ( \20306 , \20305 , \20283 );
nand \U$20054 ( \20307 , \20304 , \20306 );
not \U$20055 ( \20308 , \20307 );
xor \U$20056 ( \20309 , \20238 , \20240 );
and \U$20057 ( \20310 , \20288 , \20297 );
and \U$20058 ( \20311 , \20309 , \20310 );
not \U$20059 ( \20312 , \20309 );
not \U$20060 ( \20313 , \20310 );
and \U$20061 ( \20314 , \20312 , \20313 );
nor \U$20062 ( \20315 , \20311 , \20314 );
not \U$20063 ( \20316 , \20315 );
or \U$20064 ( \20317 , \20308 , \20316 );
nand \U$20065 ( \20318 , \20310 , \20309 );
nand \U$20066 ( \20319 , \20317 , \20318 );
xor \U$20067 ( \20320 , \20241 , \20243 );
nand \U$20068 ( \20321 , \20319 , \20320 );
nand \U$20069 ( \20322 , \20245 , \20321 );
xor \U$20070 ( \20323 , \20231 , \20220 );
nand \U$20071 ( \20324 , \20322 , \20323 );
nand \U$20072 ( \20325 , \20233 , \20324 );
not \U$20073 ( \20326 , \20325 );
xor \U$20074 ( \20327 , \20166 , \20168 );
not \U$20075 ( \20328 , \20327 );
xor \U$20076 ( \20329 , \20129 , \20144 );
xor \U$20077 ( \20330 , \20329 , \20163 );
xor \U$20078 ( \20331 , \20073 , \20082 );
xor \U$20079 ( \20332 , \20331 , \20092 );
nand \U$20080 ( \20333 , \20330 , \20332 );
not \U$20081 ( \20334 , \20333 );
and \U$20082 ( \20335 , \20328 , \20334 );
and \U$20083 ( \20336 , \20327 , \20333 );
nor \U$20084 ( \20337 , \20335 , \20336 );
not \U$20085 ( \20338 , \20332 );
nor \U$20086 ( \20339 , \20338 , \20330 );
not \U$20087 ( \20340 , \20339 );
not \U$20088 ( \20341 , \20332 );
nand \U$20089 ( \20342 , \20341 , \20330 );
nand \U$20090 ( \20343 , \20340 , \20342 );
not \U$20091 ( \20344 , \20343 );
xor \U$20092 ( \20345 , \20222 , \20226 );
not \U$20093 ( \20346 , \20229 );
and \U$20094 ( \20347 , \20345 , \20346 );
and \U$20095 ( \20348 , \20222 , \20226 );
or \U$20096 ( \20349 , \20347 , \20348 );
not \U$20097 ( \20350 , \20349 );
not \U$20098 ( \20351 , \20350 );
and \U$20099 ( \20352 , \20344 , \20351 );
and \U$20100 ( \20353 , \20343 , \20350 );
nor \U$20101 ( \20354 , \20352 , \20353 );
nor \U$20102 ( \20355 , \20337 , \20354 );
not \U$20103 ( \20356 , \20355 );
or \U$20104 ( \20357 , \20326 , \20356 );
not \U$20105 ( \20358 , \20337 );
not \U$20106 ( \20359 , \20343 );
nor \U$20107 ( \20360 , \20359 , \20350 );
and \U$20108 ( \20361 , \20358 , \20360 );
not \U$20109 ( \20362 , \20333 );
and \U$20110 ( \20363 , \20327 , \20362 );
nor \U$20111 ( \20364 , \20361 , \20363 );
nand \U$20112 ( \20365 , \20357 , \20364 );
xor \U$20113 ( \20366 , \20172 , \20169 );
nand \U$20114 ( \20367 , \20365 , \20366 );
nand \U$20115 ( \20368 , \20174 , \20367 );
xor \U$20116 ( \20369 , \20120 , \20057 );
nand \U$20117 ( \20370 , \20368 , \20369 );
nand \U$20118 ( \20371 , \20122 , \20370 );
not \U$20119 ( \20372 , \20371 );
or \U$20120 ( \20373 , \20052 , \20372 );
not \U$20121 ( \20374 , \20021 );
not \U$20122 ( \20375 , \20033 );
and \U$20123 ( \20376 , \20374 , \20375 );
not \U$20124 ( \20377 , \20050 );
not \U$20125 ( \20378 , \20002 );
not \U$20126 ( \20379 , \19999 );
not \U$20127 ( \20380 , \20379 );
and \U$20128 ( \20381 , \20378 , \20380 );
and \U$20129 ( \20382 , \20012 , \20017 );
and \U$20130 ( \20383 , \20006 , \20382 );
nor \U$20131 ( \20384 , \20381 , \20383 );
or \U$20132 ( \20385 , \20384 , \19910 );
not \U$20133 ( \20386 , \19839 );
nand \U$20134 ( \20387 , \20386 , \19906 );
nand \U$20135 ( \20388 , \20385 , \20387 );
not \U$20136 ( \20389 , \20388 );
or \U$20137 ( \20390 , \20377 , \20389 );
nand \U$20138 ( \20391 , \20044 , \20041 );
nand \U$20139 ( \20392 , \20390 , \20391 );
and \U$20140 ( \20393 , \20392 , \20034 );
nor \U$20141 ( \20394 , \20376 , \20393 );
nand \U$20142 ( \20395 , \20373 , \20394 );
not \U$20143 ( \20396 , \20395 );
or \U$20144 ( \20397 , \19624 , \20396 );
not \U$20145 ( \20398 , \19622 );
nand \U$20146 ( \20399 , \20398 , \19616 );
nand \U$20147 ( \20400 , \20397 , \20399 );
and \U$20148 ( \20401 , \19500 , \19517 , \20400 , \19502 );
nand \U$20149 ( \20402 , \19512 , \20401 );
nand \U$20150 ( \20403 , \16941 , \19513 , \20402 );
not \U$20151 ( \20404 , \14622 );
not \U$20152 ( \20405 , \20404 );
and \U$20153 ( \20406 , \20405 , RIbe27fd0_11);
and \U$20154 ( \20407 , \10919 , RIbe27f58_10);
nor \U$20155 ( \20408 , \20406 , \20407 );
and \U$20156 ( \20409 , \20408 , \8077 );
not \U$20157 ( \20410 , \20408 );
and \U$20158 ( \20411 , \20410 , \7970 );
nor \U$20159 ( \20412 , \20409 , \20411 );
buf \U$20160 ( \20413 , \20412 );
not \U$20161 ( \20414 , RIbe28f48_44);
not \U$20162 ( \20415 , \14633 );
or \U$20163 ( \20416 , \20414 , \20415 );
nand \U$20164 ( \20417 , RIbe28ed0_43, \13158 );
nand \U$20165 ( \20418 , \20416 , \20417 );
and \U$20166 ( \20419 , \20418 , \6949 );
not \U$20167 ( \20420 , \20418 );
and \U$20168 ( \20421 , \20420 , \7988 );
nor \U$20169 ( \20422 , \20419 , \20421 );
not \U$20170 ( \20423 , \20422 );
or \U$20171 ( \20424 , \20413 , \20423 );
not \U$20172 ( \20425 , RIbe29c68_72);
not \U$20173 ( \20426 , \6980 );
or \U$20174 ( \20427 , \20425 , \20426 );
nand \U$20175 ( \20428 , \13224 , RIbe29bf0_71);
nand \U$20176 ( \20429 , \20427 , \20428 );
and \U$20177 ( \20430 , \20429 , \7304 );
not \U$20178 ( \20431 , \20429 );
and \U$20179 ( \20432 , \20431 , \7301 );
nor \U$20180 ( \20433 , \20430 , \20432 );
nand \U$20181 ( \20434 , \20424 , \20433 );
nand \U$20182 ( \20435 , \20423 , \20413 );
nand \U$20183 ( \20436 , \20434 , \20435 );
not \U$20184 ( \20437 , \20436 );
not \U$20185 ( \20438 , \20437 );
not \U$20186 ( \20439 , \7098 );
nand \U$20187 ( \20440 , \5453 , RIbe2a910_99);
or \U$20188 ( \20441 , \20439 , \20440 );
not \U$20189 ( \20442 , \7098 );
nand \U$20190 ( \20443 , \20442 , RIbe2b5b8_126);
nand \U$20191 ( \20444 , \20441 , \20443 );
and \U$20192 ( \20445 , \20444 , \6637 );
not \U$20193 ( \20446 , \20444 );
and \U$20194 ( \20447 , \20446 , \6907 );
nor \U$20195 ( \20448 , \20445 , \20447 );
not \U$20196 ( \20449 , RIbe2a3e8_88);
not \U$20197 ( \20450 , \6138 );
or \U$20198 ( \20451 , \20449 , \20450 );
nand \U$20199 ( \20452 , RIbe2a370_87, \8235 );
nand \U$20200 ( \20453 , \20451 , \20452 );
not \U$20201 ( \20454 , \20453 );
not \U$20202 ( \20455 , \5740 );
and \U$20203 ( \20456 , \20454 , \20455 );
and \U$20204 ( \20457 , \20453 , \9944 );
nor \U$20205 ( \20458 , \20456 , \20457 );
xor \U$20206 ( \20459 , \20448 , \20458 );
not \U$20207 ( \20460 , RIbe2a550_91);
not \U$20208 ( \20461 , \15894 );
or \U$20209 ( \20462 , \20460 , \20461 );
nand \U$20210 ( \20463 , \5731 , RIbe2a988_100);
nand \U$20211 ( \20464 , \20462 , \20463 );
not \U$20212 ( \20465 , \4945 );
and \U$20213 ( \20466 , \20464 , \20465 );
not \U$20214 ( \20467 , \20464 );
and \U$20215 ( \20468 , \20467 , \4586 );
nor \U$20216 ( \20469 , \20466 , \20468 );
and \U$20217 ( \20470 , \20459 , \20469 );
and \U$20218 ( \20471 , \20448 , \20458 );
or \U$20219 ( \20472 , \20470 , \20471 );
not \U$20220 ( \20473 , \20472 );
or \U$20221 ( \20474 , \20438 , \20473 );
not \U$20222 ( \20475 , RIbe29e48_76);
not \U$20223 ( \20476 , \6560 );
or \U$20224 ( \20477 , \20475 , \20476 );
nand \U$20225 ( \20478 , \6963 , RIbe29dd0_75);
nand \U$20226 ( \20479 , \20477 , \20478 );
and \U$20227 ( \20480 , \20479 , \7293 );
not \U$20228 ( \20481 , \20479 );
and \U$20229 ( \20482 , \20481 , \6572 );
nor \U$20230 ( \20483 , \20480 , \20482 );
not \U$20231 ( \20484 , \20483 );
not \U$20232 ( \20485 , RIbe2a028_80);
nand \U$20233 ( \20486 , \6587 , \6588 );
not \U$20234 ( \20487 , \20486 );
not \U$20235 ( \20488 , \20487 );
or \U$20236 ( \20489 , \20485 , \20488 );
nand \U$20237 ( \20490 , \7278 , RIbe29fb0_79);
nand \U$20238 ( \20491 , \20489 , \20490 );
and \U$20239 ( \20492 , \20491 , \14991 );
not \U$20240 ( \20493 , \20491 );
and \U$20241 ( \20494 , \20493 , \6601 );
nor \U$20242 ( \20495 , \20492 , \20494 );
nand \U$20243 ( \20496 , \20484 , \20495 );
not \U$20244 ( \20497 , \13412 );
not \U$20245 ( \20498 , RIbe2a2f8_86);
not \U$20246 ( \20499 , \6535 );
or \U$20247 ( \20500 , \20498 , \20499 );
nand \U$20248 ( \20501 , \10348 , RIbe2acd0_107);
nand \U$20249 ( \20502 , \20500 , \20501 );
not \U$20250 ( \20503 , \20502 );
or \U$20251 ( \20504 , \20497 , \20503 );
or \U$20252 ( \20505 , \6548 , \20502 );
nand \U$20253 ( \20506 , \20504 , \20505 );
and \U$20254 ( \20507 , \20496 , \20506 );
nor \U$20255 ( \20508 , \20484 , \20495 );
nor \U$20256 ( \20509 , \20507 , \20508 );
not \U$20257 ( \20510 , \20509 );
nand \U$20258 ( \20511 , \20474 , \20510 );
not \U$20259 ( \20512 , \20472 );
nand \U$20260 ( \20513 , \20512 , \20436 );
nand \U$20261 ( \20514 , \20511 , \20513 );
not \U$20262 ( \20515 , \13085 );
not \U$20263 ( \20516 , RIbe28408_20);
not \U$20264 ( \20517 , \20516 );
and \U$20265 ( \20518 , \20515 , \20517 );
or \U$20266 ( \20519 , RIbe2b540_125, \12758 );
nand \U$20267 ( \20520 , \20519 , \12761 );
and \U$20268 ( \20521 , \20520 , RIbe28480_21);
nor \U$20269 ( \20522 , \20518 , \20521 );
and \U$20270 ( \20523 , \20522 , \12769 );
not \U$20271 ( \20524 , \20522 );
and \U$20272 ( \20525 , \20524 , \12773 );
or \U$20273 ( \20526 , \20523 , \20525 );
not \U$20274 ( \20527 , \20526 );
not \U$20275 ( \20528 , \12218 );
not \U$20276 ( \20529 , RIbe27e68_8);
and \U$20277 ( \20530 , \10932 , \10934 , \10930 );
not \U$20278 ( \20531 , \20530 );
or \U$20279 ( \20532 , \20529 , \20531 );
nand \U$20280 ( \20533 , \12212 , RIbe28660_25);
nand \U$20281 ( \20534 , \20532 , \20533 );
not \U$20282 ( \20535 , \20534 );
and \U$20283 ( \20536 , \20528 , \20535 );
and \U$20284 ( \20537 , \20534 , \13033 );
nor \U$20285 ( \20538 , \20536 , \20537 );
not \U$20286 ( \20539 , \20538 );
or \U$20287 ( \20540 , \20527 , \20539 );
not \U$20288 ( \20541 , \12956 );
not \U$20289 ( \20542 , RIbe285e8_24);
not \U$20290 ( \20543 , \12941 );
or \U$20291 ( \20544 , \20542 , \20543 );
nand \U$20292 ( \20545 , \12947 , RIbe287c8_28);
nand \U$20293 ( \20546 , \20544 , \20545 );
not \U$20294 ( \20547 , \20546 );
or \U$20295 ( \20548 , \20541 , \20547 );
or \U$20296 ( \20549 , \20546 , \12956 );
nand \U$20297 ( \20550 , \20548 , \20549 );
nand \U$20298 ( \20551 , \20540 , \20550 );
or \U$20299 ( \20552 , \20526 , \20538 );
nand \U$20300 ( \20553 , \20551 , \20552 );
not \U$20301 ( \20554 , RIbe28228_16);
not \U$20302 ( \20555 , \13002 );
or \U$20303 ( \20556 , \20554 , \20555 );
nand \U$20304 ( \20557 , RIbe281b0_15, RIbe2ae38_110);
nand \U$20305 ( \20558 , \20556 , \20557 );
xor \U$20306 ( \20559 , RIbe2aeb0_111, \20558 );
not \U$20307 ( \20560 , \20559 );
nand \U$20308 ( \20561 , \20560 , \1153 );
not \U$20309 ( \20562 , \20561 );
not \U$20310 ( \20563 , RIbe28930_31);
not \U$20311 ( \20564 , \12786 );
or \U$20312 ( \20565 , \20563 , \20564 );
nand \U$20313 ( \20566 , \12794 , RIbe29560_57);
nand \U$20314 ( \20567 , \20565 , \20566 );
and \U$20315 ( \20568 , \20567 , \14336 );
not \U$20316 ( \20569 , \20567 );
and \U$20317 ( \20570 , \20569 , \14335 );
nor \U$20318 ( \20571 , \20568 , \20570 );
not \U$20319 ( \20572 , \20571 );
or \U$20320 ( \20573 , \20562 , \20572 );
nand \U$20321 ( \20574 , \20559 , \1469 );
nand \U$20322 ( \20575 , \20573 , \20574 );
or \U$20323 ( \20576 , \20553 , \20575 );
not \U$20324 ( \20577 , RIbe28390_19);
not \U$20325 ( \20578 , \13063 );
or \U$20326 ( \20579 , \20577 , \20578 );
nand \U$20327 ( \20580 , \13728 , RIbe28b10_35);
nand \U$20328 ( \20581 , \20579 , \20580 );
and \U$20329 ( \20582 , \20581 , \12879 );
not \U$20330 ( \20583 , \20581 );
and \U$20331 ( \20584 , \20583 , \12723 );
nor \U$20332 ( \20585 , \20582 , \20584 );
not \U$20333 ( \20586 , RIbe28b88_36);
not \U$20334 ( \20587 , \14534 );
or \U$20335 ( \20588 , \20586 , \20587 );
nand \U$20336 ( \20589 , \12735 , RIbe29290_51);
nand \U$20337 ( \20590 , \20588 , \20589 );
and \U$20338 ( \20591 , \20590 , \14543 );
not \U$20339 ( \20592 , \20590 );
and \U$20340 ( \20593 , \20592 , \16754 );
nor \U$20341 ( \20594 , \20591 , \20593 );
not \U$20342 ( \20595 , \20594 );
or \U$20343 ( \20596 , \20585 , \20595 );
not \U$20344 ( \20597 , RIbe28a20_33);
not \U$20345 ( \20598 , \14550 );
or \U$20346 ( \20599 , \20597 , \20598 );
nand \U$20347 ( \20600 , \12834 , RIbe289a8_32);
nand \U$20348 ( \20601 , \20599 , \20600 );
not \U$20349 ( \20602 , \16366 );
and \U$20350 ( \20603 , \20601 , \20602 );
not \U$20351 ( \20604 , \20601 );
and \U$20352 ( \20605 , \20604 , \16366 );
nor \U$20353 ( \20606 , \20603 , \20605 );
nand \U$20354 ( \20607 , \20596 , \20606 );
nand \U$20355 ( \20608 , \20585 , \20595 );
nand \U$20356 ( \20609 , \20607 , \20608 );
nand \U$20357 ( \20610 , \20576 , \20609 );
nand \U$20358 ( \20611 , \20553 , \20575 );
nand \U$20359 ( \20612 , \20610 , \20611 );
or \U$20360 ( \20613 , \20514 , \20612 );
not \U$20361 ( \20614 , RIbe2ab68_104);
not \U$20362 ( \20615 , \1143 );
or \U$20363 ( \20616 , \20614 , \20615 );
nand \U$20364 ( \20617 , \1147 , RIbe2aaf0_103);
nand \U$20365 ( \20618 , \20616 , \20617 );
and \U$20366 ( \20619 , \20618 , \7899 );
not \U$20367 ( \20620 , \20618 );
and \U$20368 ( \20621 , \20620 , \1157 );
nor \U$20369 ( \20622 , \20619 , \20621 );
not \U$20370 ( \20623 , RIbe2a280_85);
not \U$20371 ( \20624 , \3701 );
nor \U$20372 ( \20625 , \20624 , \4024 );
not \U$20373 ( \20626 , \20625 );
or \U$20374 ( \20627 , \20623 , \20626 );
nand \U$20375 ( \20628 , \6787 , RIbe2a208_84);
nand \U$20376 ( \20629 , \20627 , \20628 );
xor \U$20377 ( \20630 , \20629 , \3448 );
not \U$20378 ( \20631 , \20630 );
not \U$20379 ( \20632 , RIbe2b108_116);
not \U$20380 ( \20633 , \3451 );
or \U$20381 ( \20634 , \20632 , \20633 );
nand \U$20382 ( \20635 , \6800 , RIbe2b090_115);
nand \U$20383 ( \20636 , \20634 , \20635 );
xor \U$20384 ( \20637 , \20636 , \2887 );
not \U$20385 ( \20638 , \20637 );
or \U$20386 ( \20639 , \20631 , \20638 );
not \U$20387 ( \20640 , RIbe2a190_83);
not \U$20388 ( \20641 , \6413 );
or \U$20389 ( \20642 , \20640 , \20641 );
nand \U$20390 ( \20643 , \4808 , RIbe2a5c8_92);
nand \U$20391 ( \20644 , \20642 , \20643 );
and \U$20392 ( \20645 , \20644 , \4007 );
not \U$20393 ( \20646 , \20644 );
and \U$20394 ( \20647 , \20646 , \4323 );
nor \U$20395 ( \20648 , \20645 , \20647 );
nand \U$20396 ( \20649 , \20639 , \20648 );
or \U$20397 ( \20650 , \20630 , \20637 );
nand \U$20398 ( \20651 , \20649 , \20650 );
xor \U$20399 ( \20652 , \20622 , \20651 );
not \U$20400 ( \20653 , RIbe2b180_117);
not \U$20401 ( \20654 , \10010 );
or \U$20402 ( \20655 , \20653 , \20654 );
nand \U$20403 ( \20656 , \4284 , RIbe2b270_119);
nand \U$20404 ( \20657 , \20655 , \20656 );
and \U$20405 ( \20658 , \20657 , \3481 );
not \U$20406 ( \20659 , \20657 );
and \U$20407 ( \20660 , \20659 , \2576 );
nor \U$20408 ( \20661 , \20658 , \20660 );
and \U$20409 ( \20662 , \6380 , RIbe2b018_114);
not \U$20410 ( \20663 , \6382 );
buf \U$20411 ( \20664 , \20663 );
and \U$20412 ( \20665 , \20664 , RIbe2afa0_113);
nor \U$20413 ( \20666 , \20662 , \20665 );
and \U$20414 ( \20667 , \20666 , \1448 );
not \U$20415 ( \20668 , \20666 );
and \U$20416 ( \20669 , \20668 , \1132 );
nor \U$20417 ( \20670 , \20667 , \20669 );
or \U$20418 ( \20671 , \20661 , \20670 );
not \U$20419 ( \20672 , RIbe2af28_112);
or \U$20420 ( \20673 , \1266 , RIbe29740_61);
nand \U$20421 ( \20674 , \20673 , \1269 );
not \U$20422 ( \20675 , \20674 );
or \U$20423 ( \20676 , \20672 , \20675 );
nand \U$20424 ( \20677 , \2384 , RIbe2b1f8_118);
nand \U$20425 ( \20678 , \20676 , \20677 );
not \U$20426 ( \20679 , \20678 );
not \U$20427 ( \20680 , \3516 );
and \U$20428 ( \20681 , \20679 , \20680 );
and \U$20429 ( \20682 , \20678 , \1076 );
nor \U$20430 ( \20683 , \20681 , \20682 );
not \U$20431 ( \20684 , \20683 );
nand \U$20432 ( \20685 , \20671 , \20684 );
nand \U$20433 ( \20686 , \20670 , \20661 );
nand \U$20434 ( \20687 , \20685 , \20686 );
and \U$20435 ( \20688 , \20652 , \20687 );
and \U$20436 ( \20689 , \20622 , \20651 );
or \U$20437 ( \20690 , \20688 , \20689 );
nand \U$20438 ( \20691 , \20613 , \20690 );
nand \U$20439 ( \20692 , \20514 , \20612 );
nand \U$20440 ( \20693 , \20691 , \20692 );
not \U$20441 ( \20694 , RIbe281b0_15);
not \U$20442 ( \20695 , \13690 );
or \U$20443 ( \20696 , \20694 , \20695 );
nand \U$20444 ( \20697 , RIbe280c0_13, RIbe2ae38_110);
nand \U$20445 ( \20698 , \20696 , \20697 );
xnor \U$20446 ( \20699 , \20698 , RIbe2aeb0_111);
not \U$20447 ( \20700 , RIbe29560_57);
not \U$20448 ( \20701 , \15249 );
or \U$20449 ( \20702 , \20700 , \20701 );
nand \U$20450 ( \20703 , \12794 , RIbe28228_16);
nand \U$20451 ( \20704 , \20702 , \20703 );
xor \U$20452 ( \20705 , \20704 , \14335 );
xor \U$20453 ( \20706 , \20699 , \20705 );
not \U$20454 ( \20707 , RIbe289a8_32);
not \U$20455 ( \20708 , \13590 );
or \U$20456 ( \20709 , \20707 , \20708 );
nand \U$20457 ( \20710 , \13012 , RIbe28930_31);
nand \U$20458 ( \20711 , \20709 , \20710 );
xor \U$20459 ( \20712 , \20711 , \12863 );
xor \U$20460 ( \20713 , \20706 , \20712 );
not \U$20461 ( \20714 , \20713 );
not \U$20462 ( \20715 , RIbe28b10_35);
not \U$20463 ( \20716 , \16759 );
or \U$20464 ( \20717 , \20715 , \20716 );
nand \U$20465 ( \20718 , \12710 , RIbe28b88_36);
nand \U$20466 ( \20719 , \20717 , \20718 );
and \U$20467 ( \20720 , \20719 , \13583 );
not \U$20468 ( \20721 , \20719 );
and \U$20469 ( \20722 , \20721 , \12716 );
nor \U$20470 ( \20723 , \20720 , \20722 );
not \U$20471 ( \20724 , \20723 );
not \U$20472 ( \20725 , RIbe29290_51);
not \U$20473 ( \20726 , \14534 );
or \U$20474 ( \20727 , \20725 , \20726 );
nand \U$20475 ( \20728 , \12735 , RIbe28a20_33);
nand \U$20476 ( \20729 , \20727 , \20728 );
and \U$20477 ( \20730 , \20729 , \14543 );
not \U$20478 ( \20731 , \20729 );
and \U$20479 ( \20732 , \20731 , \14358 );
nor \U$20480 ( \20733 , \20730 , \20732 );
not \U$20481 ( \20734 , \20733 );
not \U$20482 ( \20735 , \20734 );
or \U$20483 ( \20736 , \20724 , \20735 );
or \U$20484 ( \20737 , \20723 , \20734 );
nand \U$20485 ( \20738 , \20736 , \20737 );
not \U$20486 ( \20739 , \12769 );
not \U$20487 ( \20740 , RIbe28408_20);
not \U$20488 ( \20741 , \13738 );
or \U$20489 ( \20742 , \20740 , \20741 );
not \U$20490 ( \20743 , \12752 );
nand \U$20491 ( \20744 , \20743 , RIbe28390_19);
nand \U$20492 ( \20745 , \20742 , \20744 );
not \U$20493 ( \20746 , \20745 );
or \U$20494 ( \20747 , \20739 , \20746 );
or \U$20495 ( \20748 , \20745 , \12770 );
nand \U$20496 ( \20749 , \20747 , \20748 );
xor \U$20497 ( \20750 , \20738 , \20749 );
nand \U$20498 ( \20751 , \20714 , \20750 );
not \U$20499 ( \20752 , \20751 );
not \U$20500 ( \20753 , RIbe2b090_115);
not \U$20501 ( \20754 , \3451 );
or \U$20502 ( \20755 , \20753 , \20754 );
nand \U$20503 ( \20756 , \3457 , RIbe2a280_85);
nand \U$20504 ( \20757 , \20755 , \20756 );
and \U$20505 ( \20758 , \20757 , \2887 );
not \U$20506 ( \20759 , \20757 );
and \U$20507 ( \20760 , \20759 , \4346 );
nor \U$20508 ( \20761 , \20758 , \20760 );
not \U$20509 ( \20762 , \20761 );
not \U$20510 ( \20763 , RIbe2a208_84);
not \U$20511 ( \20764 , \3703 );
not \U$20512 ( \20765 , \20764 );
or \U$20513 ( \20766 , \20763 , \20765 );
not \U$20514 ( \20767 , \6786 );
nand \U$20515 ( \20768 , \20767 , RIbe2a190_83);
nand \U$20516 ( \20769 , \20766 , \20768 );
and \U$20517 ( \20770 , \20769 , \3471 );
not \U$20518 ( \20771 , \20769 );
and \U$20519 ( \20772 , \20771 , \3698 );
nor \U$20520 ( \20773 , \20770 , \20772 );
not \U$20521 ( \20774 , \20773 );
or \U$20522 ( \20775 , \20762 , \20774 );
or \U$20523 ( \20776 , \20761 , \20773 );
nand \U$20524 ( \20777 , \20775 , \20776 );
not \U$20525 ( \20778 , RIbe2b270_119);
not \U$20526 ( \20779 , \8342 );
or \U$20527 ( \20780 , \20778 , \20779 );
nand \U$20528 ( \20781 , \4284 , RIbe2b108_116);
nand \U$20529 ( \20782 , \20780 , \20781 );
not \U$20530 ( \20783 , \20782 );
not \U$20531 ( \20784 , \2379 );
and \U$20532 ( \20785 , \20783 , \20784 );
and \U$20533 ( \20786 , \20782 , \3275 );
nor \U$20534 ( \20787 , \20785 , \20786 );
and \U$20535 ( \20788 , \20777 , \20787 );
not \U$20536 ( \20789 , \20777 );
not \U$20537 ( \20790 , \20787 );
and \U$20538 ( \20791 , \20789 , \20790 );
nor \U$20539 ( \20792 , \20788 , \20791 );
not \U$20540 ( \20793 , \20792 );
not \U$20541 ( \20794 , \20793 );
not \U$20542 ( \20795 , RIbe2b5b8_126);
and \U$20543 ( \20796 , \5747 , \5453 );
not \U$20544 ( \20797 , \20796 );
or \U$20545 ( \20798 , \20795 , \20797 );
nand \U$20546 ( \20799 , \6633 , RIbe2a3e8_88);
nand \U$20547 ( \20800 , \20798 , \20799 );
not \U$20548 ( \20801 , \6640 );
and \U$20549 ( \20802 , \20800 , \20801 );
not \U$20550 ( \20803 , \20800 );
and \U$20551 ( \20804 , \20803 , \5457 );
nor \U$20552 ( \20805 , \20802 , \20804 );
not \U$20553 ( \20806 , \20805 );
not \U$20554 ( \20807 , \20806 );
not \U$20555 ( \20808 , RIbe2a988_100);
and \U$20556 ( \20809 , \5051 , \4826 );
not \U$20557 ( \20810 , \20809 );
or \U$20558 ( \20811 , \20808 , \20810 );
nand \U$20559 ( \20812 , \7056 , RIbe2a910_99);
nand \U$20560 ( \20813 , \20811 , \20812 );
and \U$20561 ( \20814 , \20813 , \4946 );
not \U$20562 ( \20815 , \20813 );
and \U$20563 ( \20816 , \20815 , \4586 );
nor \U$20564 ( \20817 , \20814 , \20816 );
not \U$20565 ( \20818 , \20817 );
not \U$20566 ( \20819 , \20818 );
or \U$20567 ( \20820 , \20807 , \20819 );
nand \U$20568 ( \20821 , \20817 , \20805 );
nand \U$20569 ( \20822 , \20820 , \20821 );
not \U$20570 ( \20823 , RIbe2a5c8_92);
not \U$20571 ( \20824 , \6413 );
or \U$20572 ( \20825 , \20823 , \20824 );
nand \U$20573 ( \20826 , \4808 , RIbe2a550_91);
nand \U$20574 ( \20827 , \20825 , \20826 );
and \U$20575 ( \20828 , \20827 , \4326 );
not \U$20576 ( \20829 , \20827 );
and \U$20577 ( \20830 , \20829 , \7865 );
nor \U$20578 ( \20831 , \20828 , \20830 );
xor \U$20579 ( \20832 , \20822 , \20831 );
not \U$20580 ( \20833 , \20832 );
or \U$20581 ( \20834 , \20794 , \20833 );
not \U$20582 ( \20835 , \1076 );
not \U$20583 ( \20836 , RIbe2b1f8_118);
not \U$20584 ( \20837 , \20674 );
or \U$20585 ( \20838 , \20836 , \20837 );
nand \U$20586 ( \20839 , \2384 , RIbe2b180_117);
nand \U$20587 ( \20840 , \20838 , \20839 );
not \U$20588 ( \20841 , \20840 );
and \U$20589 ( \20842 , \20835 , \20841 );
and \U$20590 ( \20843 , \20840 , \7038 );
nor \U$20591 ( \20844 , \20842 , \20843 );
not \U$20592 ( \20845 , \20844 );
not \U$20593 ( \20846 , RIbe2afa0_113);
not \U$20594 ( \20847 , \1111 );
or \U$20595 ( \20848 , \20846 , \20847 );
not \U$20596 ( \20849 , \6382 );
nand \U$20597 ( \20850 , RIbe2af28_112, \20849 );
nand \U$20598 ( \20851 , \20848 , \20850 );
and \U$20599 ( \20852 , \20851 , \1131 );
not \U$20600 ( \20853 , \20851 );
and \U$20601 ( \20854 , \20853 , \1123 );
nor \U$20602 ( \20855 , \20852 , \20854 );
not \U$20603 ( \20856 , \20855 );
or \U$20604 ( \20857 , \20845 , \20856 );
or \U$20605 ( \20858 , \20844 , \20855 );
nand \U$20606 ( \20859 , \20857 , \20858 );
not \U$20607 ( \20860 , RIbe2b630_127);
not \U$20608 ( \20861 , \1632 );
or \U$20609 ( \20862 , \20860 , \20861 );
nand \U$20610 ( \20863 , RIbe2b018_114, \1454 );
nand \U$20611 ( \20864 , \20862 , \20863 );
and \U$20612 ( \20865 , \20864 , \2418 );
not \U$20613 ( \20866 , \20864 );
and \U$20614 ( \20867 , \20866 , \1309 );
nor \U$20615 ( \20868 , \20865 , \20867 );
and \U$20616 ( \20869 , \20859 , \20868 );
not \U$20617 ( \20870 , \20859 );
not \U$20618 ( \20871 , \20868 );
and \U$20619 ( \20872 , \20870 , \20871 );
nor \U$20620 ( \20873 , \20869 , \20872 );
not \U$20621 ( \20874 , \20873 );
not \U$20622 ( \20875 , \20832 );
nand \U$20623 ( \20876 , \20875 , \20792 );
nand \U$20624 ( \20877 , \20874 , \20876 );
nand \U$20625 ( \20878 , \20834 , \20877 );
nor \U$20626 ( \20879 , \20752 , \20878 );
not \U$20627 ( \20880 , RIbe28ed0_43);
not \U$20628 ( \20881 , \7974 );
or \U$20629 ( \20882 , \20880 , \20881 );
nand \U$20630 ( \20883 , \13339 , RIbe27fd0_11);
nand \U$20631 ( \20884 , \20882 , \20883 );
and \U$20632 ( \20885 , \20884 , \14299 );
not \U$20633 ( \20886 , \20884 );
and \U$20634 ( \20887 , \20886 , \6948 );
nor \U$20635 ( \20888 , \20885 , \20887 );
and \U$20636 ( \20889 , \6980 , RIbe29bf0_71);
and \U$20637 ( \20890 , \13792 , RIbe28f48_44);
nor \U$20638 ( \20891 , \20889 , \20890 );
and \U$20639 ( \20892 , \20891 , \13227 );
not \U$20640 ( \20893 , \20891 );
and \U$20641 ( \20894 , \20893 , \6992 );
nor \U$20642 ( \20895 , \20892 , \20894 );
and \U$20643 ( \20896 , \20888 , \20895 );
not \U$20644 ( \20897 , \20888 );
not \U$20645 ( \20898 , \20895 );
and \U$20646 ( \20899 , \20897 , \20898 );
or \U$20647 ( \20900 , \20896 , \20899 );
not \U$20648 ( \20901 , RIbe29dd0_75);
not \U$20649 ( \20902 , \8199 );
or \U$20650 ( \20903 , \20901 , \20902 );
nand \U$20651 ( \20904 , \8202 , RIbe29c68_72);
nand \U$20652 ( \20905 , \20903 , \20904 );
and \U$20653 ( \20906 , \20905 , \7293 );
not \U$20654 ( \20907 , \20905 );
and \U$20655 ( \20908 , \20907 , \6572 );
nor \U$20656 ( \20909 , \20906 , \20908 );
xor \U$20657 ( \20910 , \20900 , \20909 );
not \U$20658 ( \20911 , \12957 );
not \U$20659 ( \20912 , RIbe287c8_28);
not \U$20660 ( \20913 , \12942 );
or \U$20661 ( \20914 , \20912 , \20913 );
nand \U$20662 ( \20915 , \12947 , RIbe28480_21);
nand \U$20663 ( \20916 , \20914 , \20915 );
not \U$20664 ( \20917 , \20916 );
or \U$20665 ( \20918 , \20911 , \20917 );
or \U$20666 ( \20919 , \20916 , \12957 );
nand \U$20667 ( \20920 , \20918 , \20919 );
not \U$20668 ( \20921 , \20920 );
not \U$20669 ( \20922 , RIbe28660_25);
not \U$20670 ( \20923 , \13024 );
or \U$20671 ( \20924 , \20922 , \20923 );
nand \U$20672 ( \20925 , \12212 , RIbe285e8_24);
nand \U$20673 ( \20926 , \20924 , \20925 );
not \U$20674 ( \20927 , \20926 );
not \U$20675 ( \20928 , \13033 );
and \U$20676 ( \20929 , \20927 , \20928 );
and \U$20677 ( \20930 , \20926 , \13661 );
nor \U$20678 ( \20931 , \20929 , \20930 );
not \U$20679 ( \20932 , \20931 );
or \U$20680 ( \20933 , \20921 , \20932 );
or \U$20681 ( \20934 , \20931 , \20920 );
nand \U$20682 ( \20935 , \20933 , \20934 );
and \U$20683 ( \20936 , \8276 , RIbe27f58_10);
and \U$20684 ( \20937 , \13038 , RIbe27e68_8);
nor \U$20685 ( \20938 , \20936 , \20937 );
and \U$20686 ( \20939 , \20938 , \16437 );
not \U$20687 ( \20940 , \20938 );
and \U$20688 ( \20941 , \20940 , \12202 );
nor \U$20689 ( \20942 , \20939 , \20941 );
not \U$20690 ( \20943 , \20942 );
buf \U$20691 ( \20944 , \20943 );
and \U$20692 ( \20945 , \20935 , \20944 );
not \U$20693 ( \20946 , \20935 );
not \U$20694 ( \20947 , \20944 );
and \U$20695 ( \20948 , \20946 , \20947 );
nor \U$20696 ( \20949 , \20945 , \20948 );
or \U$20697 ( \20950 , \20910 , \20949 );
and \U$20698 ( \20951 , \6535 , RIbe2acd0_107);
and \U$20699 ( \20952 , \6884 , RIbe2a028_80);
nor \U$20700 ( \20953 , \20951 , \20952 );
and \U$20701 ( \20954 , \20953 , \13412 );
not \U$20702 ( \20955 , \20953 );
and \U$20703 ( \20956 , \20955 , \15730 );
nor \U$20704 ( \20957 , \20954 , \20956 );
not \U$20705 ( \20958 , RIbe29fb0_79);
not \U$20706 ( \20959 , \6591 );
or \U$20707 ( \20960 , \20958 , \20959 );
nand \U$20708 ( \20961 , \13436 , RIbe29e48_76);
nand \U$20709 ( \20962 , \20960 , \20961 );
and \U$20710 ( \20963 , \20962 , \6582 );
not \U$20711 ( \20964 , \20962 );
and \U$20712 ( \20965 , \20964 , \7949 );
nor \U$20713 ( \20966 , \20963 , \20965 );
xor \U$20714 ( \20967 , \20957 , \20966 );
not \U$20715 ( \20968 , \5740 );
not \U$20716 ( \20969 , RIbe2a370_87);
not \U$20717 ( \20970 , \12268 );
or \U$20718 ( \20971 , \20969 , \20970 );
nand \U$20719 ( \20972 , \8235 , RIbe2a2f8_86);
nand \U$20720 ( \20973 , \20971 , \20972 );
not \U$20721 ( \20974 , \20973 );
or \U$20722 ( \20975 , \20968 , \20974 );
or \U$20723 ( \20976 , \20973 , \9944 );
nand \U$20724 ( \20977 , \20975 , \20976 );
xor \U$20725 ( \20978 , \20967 , \20977 );
and \U$20726 ( \20979 , \20950 , \20978 );
and \U$20727 ( \20980 , \20910 , \20949 );
nor \U$20728 ( \20981 , \20979 , \20980 );
or \U$20729 ( \20982 , \20879 , \20981 );
not \U$20730 ( \20983 , \20751 );
nand \U$20731 ( \20984 , \20878 , \20983 );
nand \U$20732 ( \20985 , \20982 , \20984 );
xor \U$20733 ( \20986 , \20693 , \20985 );
not \U$20734 ( \20987 , \12998 );
not \U$20735 ( \20988 , RIbe28228_16);
not \U$20736 ( \20989 , \12787 );
or \U$20737 ( \20990 , \20988 , \20989 );
nand \U$20738 ( \20991 , \12794 , RIbe281b0_15);
nand \U$20739 ( \20992 , \20990 , \20991 );
not \U$20740 ( \20993 , \20992 );
or \U$20741 ( \20994 , \20987 , \20993 );
or \U$20742 ( \20995 , \20992 , \12893 );
nand \U$20743 ( \20996 , \20994 , \20995 );
not \U$20744 ( \20997 , RIbe280c0_13);
not \U$20745 ( \20998 , \12811 );
or \U$20746 ( \20999 , \20997 , \20998 );
nand \U$20747 ( \21000 , RIbe29830_63, RIbe2ae38_110);
nand \U$20748 ( \21001 , \20999 , \21000 );
xnor \U$20749 ( \21002 , \21001 , RIbe2aeb0_111);
not \U$20750 ( \21003 , \21002 );
xor \U$20751 ( \21004 , \1011 , \21003 );
xor \U$20752 ( \21005 , \20996 , \21004 );
not \U$20753 ( \21006 , RIbe28a20_33);
not \U$20754 ( \21007 , \14534 );
or \U$20755 ( \21008 , \21006 , \21007 );
nand \U$20756 ( \21009 , \12735 , RIbe289a8_32);
nand \U$20757 ( \21010 , \21008 , \21009 );
and \U$20758 ( \21011 , \21010 , \14543 );
not \U$20759 ( \21012 , \21010 );
not \U$20760 ( \21013 , \14543 );
and \U$20761 ( \21014 , \21012 , \21013 );
nor \U$20762 ( \21015 , \21011 , \21014 );
not \U$20763 ( \21016 , RIbe28930_31);
not \U$20764 ( \21017 , \12858 );
or \U$20765 ( \21018 , \21016 , \21017 );
nand \U$20766 ( \21019 , \12834 , RIbe29560_57);
nand \U$20767 ( \21020 , \21018 , \21019 );
xnor \U$20768 ( \21021 , \21020 , \16366 );
xor \U$20769 ( \21022 , \21015 , \21021 );
not \U$20770 ( \21023 , RIbe28b88_36);
not \U$20771 ( \21024 , \16759 );
or \U$20772 ( \21025 , \21023 , \21024 );
nand \U$20773 ( \21026 , \13728 , RIbe29290_51);
nand \U$20774 ( \21027 , \21025 , \21026 );
and \U$20775 ( \21028 , \21027 , \12723 );
not \U$20776 ( \21029 , \21027 );
and \U$20777 ( \21030 , \21029 , \12879 );
nor \U$20778 ( \21031 , \21028 , \21030 );
xnor \U$20779 ( \21032 , \21022 , \21031 );
and \U$20780 ( \21033 , \21005 , \21032 );
not \U$20781 ( \21034 , \21005 );
not \U$20782 ( \21035 , \21032 );
and \U$20783 ( \21036 , \21034 , \21035 );
or \U$20784 ( \21037 , \21033 , \21036 );
not \U$20785 ( \21038 , \21037 );
not \U$20786 ( \21039 , RIbe2a550_91);
and \U$20787 ( \21040 , \4313 , \4314 );
not \U$20788 ( \21041 , \21040 );
or \U$20789 ( \21042 , \21039 , \21041 );
not \U$20790 ( \21043 , \4598 );
nand \U$20791 ( \21044 , \21043 , RIbe2a988_100);
nand \U$20792 ( \21045 , \21042 , \21044 );
and \U$20793 ( \21046 , \21045 , \4326 );
not \U$20794 ( \21047 , \21045 );
and \U$20795 ( \21048 , \21047 , \4323 );
nor \U$20796 ( \21049 , \21046 , \21048 );
not \U$20797 ( \21050 , \21049 );
not \U$20798 ( \21051 , RIbe2a190_83);
not \U$20799 ( \21052 , \20625 );
or \U$20800 ( \21053 , \21051 , \21052 );
nand \U$20801 ( \21054 , \6787 , RIbe2a5c8_92);
nand \U$20802 ( \21055 , \21053 , \21054 );
not \U$20803 ( \21056 , \21055 );
not \U$20804 ( \21057 , \3698 );
and \U$20805 ( \21058 , \21056 , \21057 );
and \U$20806 ( \21059 , \21055 , \3448 );
nor \U$20807 ( \21060 , \21058 , \21059 );
not \U$20808 ( \21061 , \21060 );
or \U$20809 ( \21062 , \21050 , \21061 );
or \U$20810 ( \21063 , \21049 , \21060 );
nand \U$20811 ( \21064 , \21062 , \21063 );
not \U$20812 ( \21065 , RIbe2a280_85);
not \U$20813 ( \21066 , \3451 );
or \U$20814 ( \21067 , \21065 , \21066 );
nand \U$20815 ( \21068 , \3457 , RIbe2a208_84);
nand \U$20816 ( \21069 , \21067 , \21068 );
and \U$20817 ( \21070 , \21069 , \2887 );
not \U$20818 ( \21071 , \21069 );
and \U$20819 ( \21072 , \21071 , \4346 );
nor \U$20820 ( \21073 , \21070 , \21072 );
not \U$20821 ( \21074 , \21073 );
and \U$20822 ( \21075 , \21064 , \21074 );
not \U$20823 ( \21076 , \21064 );
and \U$20824 ( \21077 , \21076 , \21073 );
nor \U$20825 ( \21078 , \21075 , \21077 );
not \U$20826 ( \21079 , \21078 );
not \U$20827 ( \21080 , RIbe2a2f8_86);
and \U$20828 ( \21081 , \6614 , \6134 );
not \U$20829 ( \21082 , \21081 );
or \U$20830 ( \21083 , \21080 , \21082 );
not \U$20831 ( \21084 , \6615 );
nand \U$20832 ( \21085 , \21084 , RIbe2acd0_107);
nand \U$20833 ( \21086 , \21083 , \21085 );
not \U$20834 ( \21087 , RIbe29d58_74);
not \U$20835 ( \21088 , RIbe29ce0_73);
or \U$20836 ( \21089 , \21087 , \21088 );
nand \U$20837 ( \21090 , \21089 , RIbe29b78_70);
and \U$20838 ( \21091 , \21086 , \21090 );
not \U$20839 ( \21092 , \21086 );
not \U$20840 ( \21093 , \21090 );
and \U$20841 ( \21094 , \21092 , \21093 );
nor \U$20842 ( \21095 , \21091 , \21094 );
not \U$20843 ( \21096 , RIbe2a910_99);
not \U$20844 ( \21097 , \4828 );
not \U$20845 ( \21098 , \21097 );
or \U$20846 ( \21099 , \21096 , \21098 );
nand \U$20847 ( \21100 , \7056 , RIbe2b5b8_126);
nand \U$20848 ( \21101 , \21099 , \21100 );
not \U$20849 ( \21102 , \21101 );
not \U$20850 ( \21103 , \4946 );
and \U$20851 ( \21104 , \21102 , \21103 );
and \U$20852 ( \21105 , \21101 , \4592 );
nor \U$20853 ( \21106 , \21104 , \21105 );
xor \U$20854 ( \21107 , \21095 , \21106 );
not \U$20855 ( \21108 , RIbe2a3e8_88);
not \U$20856 ( \21109 , \6630 );
or \U$20857 ( \21110 , \21108 , \21109 );
nand \U$20858 ( \21111 , \20439 , RIbe2a370_87);
nand \U$20859 ( \21112 , \21110 , \21111 );
not \U$20860 ( \21113 , \21112 );
not \U$20861 ( \21114 , \5754 );
and \U$20862 ( \21115 , \21113 , \21114 );
and \U$20863 ( \21116 , \21112 , \5754 );
nor \U$20864 ( \21117 , \21115 , \21116 );
xor \U$20865 ( \21118 , \21107 , \21117 );
not \U$20866 ( \21119 , \21118 );
or \U$20867 ( \21120 , \21079 , \21119 );
or \U$20868 ( \21121 , \21118 , \21078 );
nand \U$20869 ( \21122 , \21120 , \21121 );
not \U$20870 ( \21123 , \2385 );
not \U$20871 ( \21124 , \13109 );
and \U$20872 ( \21125 , \21123 , \21124 );
and \U$20873 ( \21126 , \8833 , RIbe2b180_117);
nor \U$20874 ( \21127 , \21125 , \21126 );
and \U$20875 ( \21128 , \21127 , \1277 );
not \U$20876 ( \21129 , \21127 );
and \U$20877 ( \21130 , \21129 , \1076 );
nor \U$20878 ( \21131 , \21128 , \21130 );
not \U$20879 ( \21132 , RIbe2b108_116);
not \U$20880 ( \21133 , \7007 );
or \U$20881 ( \21134 , \21132 , \21133 );
nand \U$20882 ( \21135 , \3267 , RIbe2b090_115);
nand \U$20883 ( \21136 , \21134 , \21135 );
and \U$20884 ( \21137 , \21136 , \7457 );
not \U$20885 ( \21138 , \21136 );
and \U$20886 ( \21139 , \21138 , \2379 );
nor \U$20887 ( \21140 , \21137 , \21139 );
and \U$20888 ( \21141 , \21131 , \21140 );
not \U$20889 ( \21142 , \21131 );
not \U$20890 ( \21143 , \21140 );
and \U$20891 ( \21144 , \21142 , \21143 );
or \U$20892 ( \21145 , \21141 , \21144 );
and \U$20893 ( \21146 , \10759 , RIbe2af28_112);
and \U$20894 ( \21147 , \10761 , RIbe2b1f8_118);
nor \U$20895 ( \21148 , \21146 , \21147 );
and \U$20896 ( \21149 , \21148 , \1132 );
not \U$20897 ( \21150 , \21148 );
and \U$20898 ( \21151 , \21150 , \2563 );
nor \U$20899 ( \21152 , \21149 , \21151 );
xnor \U$20900 ( \21153 , \21145 , \21152 );
not \U$20901 ( \21154 , \21153 );
and \U$20902 ( \21155 , \21122 , \21154 );
not \U$20903 ( \21156 , \21122 );
and \U$20904 ( \21157 , \21156 , \21153 );
nor \U$20905 ( \21158 , \21155 , \21157 );
nand \U$20906 ( \21159 , \21038 , \21158 );
not \U$20907 ( \21160 , \21159 );
not \U$20908 ( \21161 , \12751 );
not \U$20909 ( \21162 , RIbe28b10_35);
not \U$20910 ( \21163 , \21162 );
and \U$20911 ( \21164 , \21161 , \21163 );
and \U$20912 ( \21165 , \20520 , RIbe28390_19);
nor \U$20913 ( \21166 , \21164 , \21165 );
and \U$20914 ( \21167 , \21166 , \12774 );
not \U$20915 ( \21168 , \21166 );
and \U$20916 ( \21169 , \21168 , \12769 );
nor \U$20917 ( \21170 , \21167 , \21169 );
not \U$20918 ( \21171 , \12956 );
not \U$20919 ( \21172 , RIbe28480_21);
not \U$20920 ( \21173 , \12942 );
or \U$20921 ( \21174 , \21172 , \21173 );
nand \U$20922 ( \21175 , \12947 , RIbe28408_20);
nand \U$20923 ( \21176 , \21174 , \21175 );
not \U$20924 ( \21177 , \21176 );
or \U$20925 ( \21178 , \21171 , \21177 );
or \U$20926 ( \21179 , \21176 , \17005 );
nand \U$20927 ( \21180 , \21178 , \21179 );
xor \U$20928 ( \21181 , \21170 , \21180 );
not \U$20929 ( \21182 , RIbe285e8_24);
not \U$20930 ( \21183 , \20530 );
or \U$20931 ( \21184 , \21182 , \21183 );
nand \U$20932 ( \21185 , \12212 , RIbe287c8_28);
nand \U$20933 ( \21186 , \21184 , \21185 );
not \U$20934 ( \21187 , \21186 );
not \U$20935 ( \21188 , \13661 );
and \U$20936 ( \21189 , \21187 , \21188 );
and \U$20937 ( \21190 , \10940 , \21186 );
nor \U$20938 ( \21191 , \21189 , \21190 );
buf \U$20939 ( \21192 , \21191 );
xnor \U$20940 ( \21193 , \21181 , \21192 );
not \U$20941 ( \21194 , \21193 );
not \U$20942 ( \21195 , \21194 );
not \U$20943 ( \21196 , \20404 );
and \U$20944 ( \21197 , \21196 , RIbe27e68_8);
and \U$20945 ( \21198 , \10919 , RIbe28660_25);
nor \U$20946 ( \21199 , \21197 , \21198 );
and \U$20947 ( \21200 , \21199 , \7969 );
not \U$20948 ( \21201 , \21199 );
and \U$20949 ( \21202 , \21201 , \7970 );
nor \U$20950 ( \21203 , \21200 , \21202 );
not \U$20951 ( \21204 , RIbe27fd0_11);
not \U$20952 ( \21205 , \14633 );
or \U$20953 ( \21206 , \21204 , \21205 );
nand \U$20954 ( \21207 , \8269 , RIbe27f58_10);
nand \U$20955 ( \21208 , \21206 , \21207 );
and \U$20956 ( \21209 , \21208 , \6949 );
not \U$20957 ( \21210 , \21208 );
and \U$20958 ( \21211 , \21210 , \14299 );
nor \U$20959 ( \21212 , \21209 , \21211 );
xor \U$20960 ( \21213 , \21203 , \21212 );
not \U$20961 ( \21214 , \6992 );
not \U$20962 ( \21215 , RIbe28f48_44);
not \U$20963 ( \21216 , \6980 );
or \U$20964 ( \21217 , \21215 , \21216 );
nand \U$20965 ( \21218 , \6985 , RIbe28ed0_43);
nand \U$20966 ( \21219 , \21217 , \21218 );
not \U$20967 ( \21220 , \21219 );
or \U$20968 ( \21221 , \21214 , \21220 );
or \U$20969 ( \21222 , \21219 , \10902 );
nand \U$20970 ( \21223 , \21221 , \21222 );
not \U$20971 ( \21224 , \21223 );
xor \U$20972 ( \21225 , \21213 , \21224 );
not \U$20973 ( \21226 , \21225 );
not \U$20974 ( \21227 , \21226 );
or \U$20975 ( \21228 , \21195 , \21227 );
nand \U$20976 ( \21229 , \21225 , \21193 );
nand \U$20977 ( \21230 , \21228 , \21229 );
not \U$20978 ( \21231 , RIbe29e48_76);
not \U$20979 ( \21232 , \6591 );
or \U$20980 ( \21233 , \21231 , \21232 );
nand \U$20981 ( \21234 , \13436 , RIbe29dd0_75);
nand \U$20982 ( \21235 , \21233 , \21234 );
and \U$20983 ( \21236 , \21235 , \6601 );
not \U$20984 ( \21237 , \21235 );
not \U$20985 ( \21238 , \7948 );
and \U$20986 ( \21239 , \21237 , \21238 );
nor \U$20987 ( \21240 , \21236 , \21239 );
not \U$20988 ( \21241 , RIbe29c68_72);
not \U$20989 ( \21242 , \6560 );
or \U$20990 ( \21243 , \21241 , \21242 );
nand \U$20991 ( \21244 , \7958 , RIbe29bf0_71);
nand \U$20992 ( \21245 , \21243 , \21244 );
and \U$20993 ( \21246 , \21245 , \7293 );
not \U$20994 ( \21247 , \21245 );
and \U$20995 ( \21248 , \21247 , \6569 );
nor \U$20996 ( \21249 , \21246 , \21248 );
xor \U$20997 ( \21250 , \21240 , \21249 );
not \U$20998 ( \21251 , RIbe2a028_80);
not \U$20999 ( \21252 , \6535 );
or \U$21000 ( \21253 , \21251 , \21252 );
nand \U$21001 ( \21254 , \10348 , RIbe29fb0_79);
nand \U$21002 ( \21255 , \21253 , \21254 );
and \U$21003 ( \21256 , \21255 , \6552 );
not \U$21004 ( \21257 , \21255 );
and \U$21005 ( \21258 , \21257 , \7546 );
nor \U$21006 ( \21259 , \21256 , \21258 );
not \U$21007 ( \21260 , \21259 );
and \U$21008 ( \21261 , \21250 , \21260 );
not \U$21009 ( \21262 , \21250 );
and \U$21010 ( \21263 , \21262 , \21259 );
nor \U$21011 ( \21264 , \21261 , \21263 );
not \U$21012 ( \21265 , \21264 );
and \U$21013 ( \21266 , \21230 , \21265 );
not \U$21014 ( \21267 , \21230 );
and \U$21015 ( \21268 , \21267 , \21264 );
nor \U$21016 ( \21269 , \21266 , \21268 );
not \U$21017 ( \21270 , \21269 );
or \U$21018 ( \21271 , \21160 , \21270 );
not \U$21019 ( \21272 , \21158 );
nand \U$21020 ( \21273 , \21272 , \21037 );
nand \U$21021 ( \21274 , \21271 , \21273 );
and \U$21022 ( \21275 , \20986 , \21274 );
and \U$21023 ( \21276 , \20693 , \20985 );
or \U$21024 ( \21277 , \21275 , \21276 );
not \U$21025 ( \21278 , \21277 );
not \U$21026 ( \21279 , \20942 );
not \U$21027 ( \21280 , \20931 );
or \U$21028 ( \21281 , \21279 , \21280 );
nand \U$21029 ( \21282 , \21281 , \20920 );
not \U$21030 ( \21283 , \20931 );
nand \U$21031 ( \21284 , \21283 , \20943 );
nand \U$21032 ( \21285 , \21282 , \21284 );
not \U$21033 ( \21286 , \21285 );
not \U$21034 ( \21287 , \21286 );
nand \U$21035 ( \21288 , \20733 , \20723 );
and \U$21036 ( \21289 , \21288 , \20749 );
nor \U$21037 ( \21290 , \20733 , \20723 );
nor \U$21038 ( \21291 , \21289 , \21290 );
not \U$21039 ( \21292 , \21291 );
not \U$21040 ( \21293 , \21292 );
or \U$21041 ( \21294 , \21287 , \21293 );
nand \U$21042 ( \21295 , \21291 , \21285 );
nand \U$21043 ( \21296 , \21294 , \21295 );
not \U$21044 ( \21297 , \21296 );
xor \U$21045 ( \21298 , \20699 , \20705 );
and \U$21046 ( \21299 , \21298 , \20712 );
and \U$21047 ( \21300 , \20699 , \20705 );
or \U$21048 ( \21301 , \21299 , \21300 );
not \U$21049 ( \21302 , \21301 );
and \U$21050 ( \21303 , \21297 , \21302 );
and \U$21051 ( \21304 , \21296 , \21301 );
nor \U$21052 ( \21305 , \21303 , \21304 );
not \U$21053 ( \21306 , \20966 );
not \U$21054 ( \21307 , \20977 );
or \U$21055 ( \21308 , \21306 , \21307 );
or \U$21056 ( \21309 , \20966 , \20977 );
nand \U$21057 ( \21310 , \21309 , \20957 );
nand \U$21058 ( \21311 , \21308 , \21310 );
not \U$21059 ( \21312 , \20805 );
not \U$21060 ( \21313 , \20831 );
or \U$21061 ( \21314 , \21312 , \21313 );
or \U$21062 ( \21315 , \20831 , \20805 );
nand \U$21063 ( \21316 , \21315 , \20818 );
nand \U$21064 ( \21317 , \21314 , \21316 );
xor \U$21065 ( \21318 , \21311 , \21317 );
or \U$21066 ( \21319 , \20909 , \20888 );
nand \U$21067 ( \21320 , \21319 , \20898 );
nand \U$21068 ( \21321 , \20888 , \20909 );
nand \U$21069 ( \21322 , \21320 , \21321 );
xor \U$21070 ( \21323 , \21318 , \21322 );
not \U$21071 ( \21324 , \21323 );
nand \U$21072 ( \21325 , \21305 , \21324 );
not \U$21073 ( \21326 , \20855 );
and \U$21074 ( \21327 , \21326 , \20868 );
nor \U$21075 ( \21328 , \21327 , \20844 );
nor \U$21076 ( \21329 , \20868 , \21326 );
nor \U$21077 ( \21330 , \21328 , \21329 );
nand \U$21078 ( \21331 , \20761 , \20787 );
and \U$21079 ( \21332 , \21331 , \20773 );
nor \U$21080 ( \21333 , \20761 , \20787 );
nor \U$21081 ( \21334 , \21332 , \21333 );
xor \U$21082 ( \21335 , \21330 , \21334 );
nand \U$21083 ( \21336 , \1202 , RIbe2ab68_104);
and \U$21084 ( \21337 , \21336 , \1813 );
not \U$21085 ( \21338 , \21336 );
and \U$21086 ( \21339 , \21338 , \1010 );
nor \U$21087 ( \21340 , \21337 , \21339 );
not \U$21088 ( \21341 , RIbe2aaf0_103);
not \U$21089 ( \21342 , \1138 );
nand \U$21090 ( \21343 , \21342 , \1140 );
not \U$21091 ( \21344 , \21343 );
not \U$21092 ( \21345 , \21344 );
or \U$21093 ( \21346 , \21341 , \21345 );
nand \U$21094 ( \21347 , RIbe2b630_127, \1146 );
nand \U$21095 ( \21348 , \21346 , \21347 );
and \U$21096 ( \21349 , \21348 , \1154 );
not \U$21097 ( \21350 , \21348 );
and \U$21098 ( \21351 , \21350 , \8327 );
nor \U$21099 ( \21352 , \21349 , \21351 );
xor \U$21100 ( \21353 , \21340 , \21352 );
not \U$21101 ( \21354 , \2418 );
not \U$21102 ( \21355 , RIbe2b018_114);
not \U$21103 ( \21356 , \1632 );
or \U$21104 ( \21357 , \21355 , \21356 );
nand \U$21105 ( \21358 , \4730 , RIbe2afa0_113);
nand \U$21106 ( \21359 , \21357 , \21358 );
not \U$21107 ( \21360 , \21359 );
or \U$21108 ( \21361 , \21354 , \21360 );
or \U$21109 ( \21362 , \21359 , \4251 );
nand \U$21110 ( \21363 , \21361 , \21362 );
xnor \U$21111 ( \21364 , \21353 , \21363 );
xor \U$21112 ( \21365 , \21335 , \21364 );
not \U$21113 ( \21366 , \21365 );
and \U$21114 ( \21367 , \21325 , \21366 );
nor \U$21115 ( \21368 , \21305 , \21324 );
nor \U$21116 ( \21369 , \21367 , \21368 );
not \U$21117 ( \21370 , \21369 );
not \U$21118 ( \21371 , \21170 );
not \U$21119 ( \21372 , \21191 );
or \U$21120 ( \21373 , \21371 , \21372 );
nand \U$21121 ( \21374 , \21373 , \21180 );
or \U$21122 ( \21375 , \21170 , \21191 );
nand \U$21123 ( \21376 , \21374 , \21375 );
not \U$21124 ( \21377 , \21376 );
not \U$21125 ( \21378 , \21377 );
nand \U$21126 ( \21379 , \21015 , \21031 );
and \U$21127 ( \21380 , \21379 , \21021 );
nor \U$21128 ( \21381 , \21031 , \21015 );
nor \U$21129 ( \21382 , \21380 , \21381 );
not \U$21130 ( \21383 , \21382 );
not \U$21131 ( \21384 , \21383 );
or \U$21132 ( \21385 , \21378 , \21384 );
nand \U$21133 ( \21386 , \21382 , \21376 );
nand \U$21134 ( \21387 , \21385 , \21386 );
nand \U$21135 ( \21388 , \21002 , \1813 );
and \U$21136 ( \21389 , \20996 , \21388 );
nor \U$21137 ( \21390 , \21002 , \1813 );
nor \U$21138 ( \21391 , \21389 , \21390 );
and \U$21139 ( \21392 , \21387 , \21391 );
not \U$21140 ( \21393 , \21387 );
not \U$21141 ( \21394 , \21391 );
and \U$21142 ( \21395 , \21393 , \21394 );
nor \U$21143 ( \21396 , \21392 , \21395 );
not \U$21144 ( \21397 , \21340 );
not \U$21145 ( \21398 , \21352 );
nand \U$21146 ( \21399 , \21397 , \21398 );
and \U$21147 ( \21400 , \21399 , \21363 );
not \U$21148 ( \21401 , \21340 );
nor \U$21149 ( \21402 , \21401 , \21398 );
nor \U$21150 ( \21403 , \21400 , \21402 );
not \U$21151 ( \21404 , \21403 );
not \U$21152 ( \21405 , \21404 );
not \U$21153 ( \21406 , \21060 );
not \U$21154 ( \21407 , \21073 );
or \U$21155 ( \21408 , \21406 , \21407 );
nand \U$21156 ( \21409 , \21408 , \21049 );
not \U$21157 ( \21410 , \21060 );
nand \U$21158 ( \21411 , \21410 , \21074 );
nand \U$21159 ( \21412 , \21409 , \21411 );
not \U$21160 ( \21413 , \21412 );
not \U$21161 ( \21414 , \21413 );
or \U$21162 ( \21415 , \21405 , \21414 );
nand \U$21163 ( \21416 , \21403 , \21412 );
nand \U$21164 ( \21417 , \21415 , \21416 );
not \U$21165 ( \21418 , \21417 );
and \U$21166 ( \21419 , \21143 , \21152 );
nor \U$21167 ( \21420 , \21419 , \21131 );
nor \U$21168 ( \21421 , \21143 , \21152 );
nor \U$21169 ( \21422 , \21420 , \21421 );
not \U$21170 ( \21423 , \21422 );
and \U$21171 ( \21424 , \21418 , \21423 );
and \U$21172 ( \21425 , \21417 , \21422 );
nor \U$21173 ( \21426 , \21424 , \21425 );
xor \U$21174 ( \21427 , \21396 , \21426 );
xor \U$21175 ( \21428 , \21095 , \21106 );
and \U$21176 ( \21429 , \21428 , \21117 );
and \U$21177 ( \21430 , \21095 , \21106 );
or \U$21178 ( \21431 , \21429 , \21430 );
not \U$21179 ( \21432 , \21249 );
not \U$21180 ( \21433 , \21240 );
or \U$21181 ( \21434 , \21432 , \21433 );
or \U$21182 ( \21435 , \21240 , \21249 );
nand \U$21183 ( \21436 , \21435 , \21259 );
nand \U$21184 ( \21437 , \21434 , \21436 );
not \U$21185 ( \21438 , \21437 );
not \U$21186 ( \21439 , \21438 );
not \U$21187 ( \21440 , \21203 );
nand \U$21188 ( \21441 , \21440 , \21212 );
and \U$21189 ( \21442 , \21441 , \21223 );
nor \U$21190 ( \21443 , \21440 , \21212 );
nor \U$21191 ( \21444 , \21442 , \21443 );
not \U$21192 ( \21445 , \21444 );
not \U$21193 ( \21446 , \21445 );
or \U$21194 ( \21447 , \21439 , \21446 );
nand \U$21195 ( \21448 , \21444 , \21437 );
nand \U$21196 ( \21449 , \21447 , \21448 );
xor \U$21197 ( \21450 , \21431 , \21449 );
xor \U$21198 ( \21451 , \21427 , \21450 );
not \U$21199 ( \21452 , \21451 );
or \U$21200 ( \21453 , \21370 , \21452 );
not \U$21201 ( \21454 , RIbe2ab68_104);
not \U$21202 ( \21455 , \1806 );
or \U$21203 ( \21456 , \21454 , \21455 );
nand \U$21204 ( \21457 , \7905 , RIbe2aaf0_103);
nand \U$21205 ( \21458 , \21456 , \21457 );
and \U$21206 ( \21459 , \21458 , \1011 );
not \U$21207 ( \21460 , \21458 );
and \U$21208 ( \21461 , \21460 , \1608 );
nor \U$21209 ( \21462 , \21459 , \21461 );
not \U$21210 ( \21463 , RIbe2b630_127);
not \U$21211 ( \21464 , \21344 );
or \U$21212 ( \21465 , \21463 , \21464 );
nand \U$21213 ( \21466 , \1146 , RIbe2b018_114);
nand \U$21214 ( \21467 , \21465 , \21466 );
and \U$21215 ( \21468 , \21467 , \3994 );
not \U$21216 ( \21469 , \21467 );
and \U$21217 ( \21470 , \21469 , \7899 );
nor \U$21218 ( \21471 , \21468 , \21470 );
and \U$21219 ( \21472 , \21462 , \21471 );
not \U$21220 ( \21473 , \21462 );
not \U$21221 ( \21474 , \21471 );
and \U$21222 ( \21475 , \21473 , \21474 );
or \U$21223 ( \21476 , \21472 , \21475 );
not \U$21224 ( \21477 , RIbe2a208_84);
and \U$21225 ( \21478 , \3280 , \3281 );
not \U$21226 ( \21479 , \21478 );
or \U$21227 ( \21480 , \21477 , \21479 );
nand \U$21228 ( \21481 , \3456 , RIbe2a190_83);
nand \U$21229 ( \21482 , \21480 , \21481 );
not \U$21230 ( \21483 , \21482 );
not \U$21231 ( \21484 , \2887 );
or \U$21232 ( \21485 , \21483 , \21484 );
or \U$21233 ( \21486 , \21482 , \2887 );
nand \U$21234 ( \21487 , \21485 , \21486 );
not \U$21235 ( \21488 , RIbe2a5c8_92);
not \U$21236 ( \21489 , \20625 );
or \U$21237 ( \21490 , \21488 , \21489 );
not \U$21238 ( \21491 , RIbe2a550_91);
not \U$21239 ( \21492 , \21491 );
nand \U$21240 ( \21493 , \21492 , \4332 );
nand \U$21241 ( \21494 , \21490 , \21493 );
and \U$21242 ( \21495 , \21494 , \3471 );
not \U$21243 ( \21496 , \21494 );
and \U$21244 ( \21497 , \21496 , \3448 );
nor \U$21245 ( \21498 , \21495 , \21497 );
xor \U$21246 ( \21499 , \21487 , \21498 );
not \U$21247 ( \21500 , RIbe2b090_115);
not \U$21248 ( \21501 , \10010 );
or \U$21249 ( \21502 , \21500 , \21501 );
nand \U$21250 ( \21503 , \4284 , RIbe2a280_85);
nand \U$21251 ( \21504 , \21502 , \21503 );
and \U$21252 ( \21505 , \21504 , \3272 );
not \U$21253 ( \21506 , \21504 );
and \U$21254 ( \21507 , \21506 , \2379 );
nor \U$21255 ( \21508 , \21505 , \21507 );
xor \U$21256 ( \21509 , \21499 , \21508 );
xor \U$21257 ( \21510 , \21476 , \21509 );
not \U$21258 ( \21511 , \4064 );
not \U$21259 ( \21512 , RIbe2b108_116);
not \U$21260 ( \21513 , \21512 );
and \U$21261 ( \21514 , \21511 , \21513 );
and \U$21262 ( \21515 , \20674 , RIbe2b270_119);
nor \U$21263 ( \21516 , \21514 , \21515 );
and \U$21264 ( \21517 , \21516 , \1276 );
not \U$21265 ( \21518 , \21516 );
and \U$21266 ( \21519 , \21518 , \1076 );
nor \U$21267 ( \21520 , \21517 , \21519 );
not \U$21268 ( \21521 , RIbe2b1f8_118);
not \U$21269 ( \21522 , \1111 );
or \U$21270 ( \21523 , \21521 , \21522 );
nand \U$21271 ( \21524 , \20663 , RIbe2b180_117);
nand \U$21272 ( \21525 , \21523 , \21524 );
and \U$21273 ( \21526 , \21525 , \6831 );
not \U$21274 ( \21527 , \21525 );
and \U$21275 ( \21528 , \21527 , \1131 );
nor \U$21276 ( \21529 , \21526 , \21528 );
xor \U$21277 ( \21530 , \21520 , \21529 );
not \U$21278 ( \21531 , RIbe2afa0_113);
not \U$21279 ( \21532 , \1632 );
or \U$21280 ( \21533 , \21531 , \21532 );
nand \U$21281 ( \21534 , \1454 , RIbe2af28_112);
nand \U$21282 ( \21535 , \21533 , \21534 );
and \U$21283 ( \21536 , \21535 , \5125 );
not \U$21284 ( \21537 , \21535 );
and \U$21285 ( \21538 , \21537 , \1309 );
nor \U$21286 ( \21539 , \21536 , \21538 );
xnor \U$21287 ( \21540 , \21530 , \21539 );
xnor \U$21288 ( \21541 , \21510 , \21540 );
not \U$21289 ( \21542 , \10888 );
not \U$21290 ( \21543 , RIbe29dd0_75);
not \U$21291 ( \21544 , \20487 );
or \U$21292 ( \21545 , \21543 , \21544 );
nand \U$21293 ( \21546 , \7277 , RIbe29c68_72);
nand \U$21294 ( \21547 , \21545 , \21546 );
not \U$21295 ( \21548 , \21547 );
and \U$21296 ( \21549 , \21542 , \21548 );
and \U$21297 ( \21550 , \21547 , \7488 );
nor \U$21298 ( \21551 , \21549 , \21550 );
not \U$21299 ( \21552 , \21551 );
not \U$21300 ( \21553 , RIbe29fb0_79);
not \U$21301 ( \21554 , \6535 );
or \U$21302 ( \21555 , \21553 , \21554 );
nand \U$21303 ( \21556 , RIbe29e48_76, \7075 );
nand \U$21304 ( \21557 , \21555 , \21556 );
and \U$21305 ( \21558 , \21557 , \6546 );
not \U$21306 ( \21559 , \21557 );
and \U$21307 ( \21560 , \21559 , \6888 );
nor \U$21308 ( \21561 , \21558 , \21560 );
not \U$21309 ( \21562 , \21561 );
or \U$21310 ( \21563 , \21552 , \21562 );
or \U$21311 ( \21564 , \21561 , \21551 );
nand \U$21312 ( \21565 , \21563 , \21564 );
not \U$21313 ( \21566 , RIbe2acd0_107);
not \U$21314 ( \21567 , \13894 );
or \U$21315 ( \21568 , \21566 , \21567 );
nand \U$21316 ( \21569 , \6859 , RIbe2a028_80);
nand \U$21317 ( \21570 , \21568 , \21569 );
and \U$21318 ( \21571 , \21570 , \9944 );
not \U$21319 ( \21572 , \21570 );
and \U$21320 ( \21573 , \21572 , \6623 );
nor \U$21321 ( \21574 , \21571 , \21573 );
and \U$21322 ( \21575 , \21565 , \21574 );
not \U$21323 ( \21576 , \21565 );
not \U$21324 ( \21577 , \21574 );
and \U$21325 ( \21578 , \21576 , \21577 );
nor \U$21326 ( \21579 , \21575 , \21578 );
not \U$21327 ( \21580 , \21579 );
not \U$21328 ( \21581 , \8004 );
not \U$21329 ( \21582 , RIbe28ed0_43);
not \U$21330 ( \21583 , \7298 );
or \U$21331 ( \21584 , \21582 , \21583 );
nand \U$21332 ( \21585 , \13224 , RIbe27fd0_11);
nand \U$21333 ( \21586 , \21584 , \21585 );
not \U$21334 ( \21587 , \21586 );
or \U$21335 ( \21588 , \21581 , \21587 );
or \U$21336 ( \21589 , \21586 , \8004 );
nand \U$21337 ( \21590 , \21588 , \21589 );
not \U$21338 ( \21591 , \21590 );
not \U$21339 ( \21592 , RIbe27f58_10);
not \U$21340 ( \21593 , \14633 );
or \U$21341 ( \21594 , \21592 , \21593 );
nand \U$21342 ( \21595 , \8269 , RIbe27e68_8);
nand \U$21343 ( \21596 , \21594 , \21595 );
and \U$21344 ( \21597 , \21596 , \7984 );
not \U$21345 ( \21598 , \21596 );
and \U$21346 ( \21599 , \21598 , \7988 );
nor \U$21347 ( \21600 , \21597 , \21599 );
not \U$21348 ( \21601 , \21600 );
or \U$21349 ( \21602 , \21591 , \21601 );
or \U$21350 ( \21603 , \21600 , \21590 );
nand \U$21351 ( \21604 , \21602 , \21603 );
not \U$21352 ( \21605 , RIbe29bf0_71);
not \U$21353 ( \21606 , \6961 );
nand \U$21354 ( \21607 , \21606 , \6557 );
not \U$21355 ( \21608 , \21607 );
not \U$21356 ( \21609 , \21608 );
or \U$21357 ( \21610 , \21605 , \21609 );
nand \U$21358 ( \21611 , \7958 , RIbe28f48_44);
nand \U$21359 ( \21612 , \21610 , \21611 );
xor \U$21360 ( \21613 , \21612 , \6569 );
and \U$21361 ( \21614 , \21604 , \21613 );
not \U$21362 ( \21615 , \21604 );
not \U$21363 ( \21616 , \21613 );
and \U$21364 ( \21617 , \21615 , \21616 );
nor \U$21365 ( \21618 , \21614 , \21617 );
not \U$21366 ( \21619 , \21618 );
not \U$21367 ( \21620 , \21619 );
or \U$21368 ( \21621 , \21580 , \21620 );
not \U$21369 ( \21622 , \21579 );
nand \U$21370 ( \21623 , \21618 , \21622 );
nand \U$21371 ( \21624 , \21621 , \21623 );
not \U$21372 ( \21625 , RIbe2b5b8_126);
not \U$21373 ( \21626 , \20809 );
or \U$21374 ( \21627 , \21625 , \21626 );
nand \U$21375 ( \21628 , RIbe2a3e8_88, \7056 );
nand \U$21376 ( \21629 , \21627 , \21628 );
and \U$21377 ( \21630 , \21629 , \20465 );
not \U$21378 ( \21631 , \21629 );
and \U$21379 ( \21632 , \21631 , \4586 );
nor \U$21380 ( \21633 , \21630 , \21632 );
not \U$21381 ( \21634 , RIbe2a370_87);
not \U$21382 ( \21635 , \15313 );
or \U$21383 ( \21636 , \21634 , \21635 );
nand \U$21384 ( \21637 , \8246 , RIbe2a2f8_86);
nand \U$21385 ( \21638 , \21636 , \21637 );
not \U$21386 ( \21639 , \21638 );
not \U$21387 ( \21640 , \8252 );
and \U$21388 ( \21641 , \21639 , \21640 );
and \U$21389 ( \21642 , \21638 , \5046 );
nor \U$21390 ( \21643 , \21641 , \21642 );
xor \U$21391 ( \21644 , \21633 , \21643 );
not \U$21392 ( \21645 , RIbe2a988_100);
not \U$21393 ( \21646 , \4804 );
or \U$21394 ( \21647 , \21645 , \21646 );
nand \U$21395 ( \21648 , \4599 , RIbe2a910_99);
nand \U$21396 ( \21649 , \21647 , \21648 );
and \U$21397 ( \21650 , \21649 , \4323 );
not \U$21398 ( \21651 , \21649 );
and \U$21399 ( \21652 , \21651 , \4326 );
nor \U$21400 ( \21653 , \21650 , \21652 );
xor \U$21401 ( \21654 , \21644 , \21653 );
not \U$21402 ( \21655 , \21654 );
xor \U$21403 ( \21656 , \21624 , \21655 );
or \U$21404 ( \21657 , \21541 , \21656 );
nand \U$21405 ( \21658 , \21656 , \21541 );
nand \U$21406 ( \21659 , \21657 , \21658 );
not \U$21407 ( \21660 , RIbe29830_63);
not \U$21408 ( \21661 , \13690 );
or \U$21409 ( \21662 , \21660 , \21661 );
nand \U$21410 ( \21663 , RIbe296c8_60, RIbe2ae38_110);
nand \U$21411 ( \21664 , \21662 , \21663 );
xor \U$21412 ( \21665 , \21664 , RIbe2aeb0_111);
not \U$21413 ( \21666 , RIbe281b0_15);
not \U$21414 ( \21667 , \12786 );
or \U$21415 ( \21668 , \21666 , \21667 );
nand \U$21416 ( \21669 , \12794 , RIbe280c0_13);
nand \U$21417 ( \21670 , \21668 , \21669 );
and \U$21418 ( \21671 , \21670 , \14336 );
not \U$21419 ( \21672 , \21670 );
and \U$21420 ( \21673 , \21672 , \14335 );
nor \U$21421 ( \21674 , \21671 , \21673 );
xor \U$21422 ( \21675 , \21665 , \21674 );
not \U$21423 ( \21676 , RIbe29560_57);
not \U$21424 ( \21677 , \13010 );
or \U$21425 ( \21678 , \21676 , \21677 );
not \U$21426 ( \21679 , \12827 );
nand \U$21427 ( \21680 , \21679 , RIbe28228_16);
nand \U$21428 ( \21681 , \21678 , \21680 );
and \U$21429 ( \21682 , \21681 , \13595 );
not \U$21430 ( \21683 , \21681 );
and \U$21431 ( \21684 , \21683 , \12823 );
nor \U$21432 ( \21685 , \21682 , \21684 );
xor \U$21433 ( \21686 , \21675 , \21685 );
not \U$21434 ( \21687 , RIbe289a8_32);
not \U$21435 ( \21688 , \13074 );
or \U$21436 ( \21689 , \21687 , \21688 );
nand \U$21437 ( \21690 , RIbe28930_31, \12735 );
nand \U$21438 ( \21691 , \21689 , \21690 );
and \U$21439 ( \21692 , \21691 , \12741 );
not \U$21440 ( \21693 , \21691 );
and \U$21441 ( \21694 , \21693 , \15166 );
nor \U$21442 ( \21695 , \21692 , \21694 );
not \U$21443 ( \21696 , RIbe29290_51);
not \U$21444 ( \21697 , \12707 );
or \U$21445 ( \21698 , \21696 , \21697 );
nand \U$21446 ( \21699 , \13728 , RIbe28a20_33);
nand \U$21447 ( \21700 , \21698 , \21699 );
xor \U$21448 ( \21701 , \21700 , \12723 );
xor \U$21449 ( \21702 , \21695 , \21701 );
not \U$21450 ( \21703 , \12752 );
not \U$21451 ( \21704 , RIbe28b88_36);
not \U$21452 ( \21705 , \21704 );
and \U$21453 ( \21706 , \21703 , \21705 );
and \U$21454 ( \21707 , \12921 , RIbe28b10_35);
nor \U$21455 ( \21708 , \21706 , \21707 );
and \U$21456 ( \21709 , \21708 , \12927 );
not \U$21457 ( \21710 , \21708 );
and \U$21458 ( \21711 , \21710 , \12769 );
nor \U$21459 ( \21712 , \21709 , \21711 );
xor \U$21460 ( \21713 , \21702 , \21712 );
not \U$21461 ( \21714 , \21713 );
xor \U$21462 ( \21715 , \21686 , \21714 );
not \U$21463 ( \21716 , RIbe287c8_28);
not \U$21464 ( \21717 , \10936 );
or \U$21465 ( \21718 , \21716 , \21717 );
nand \U$21466 ( \21719 , \12213 , RIbe28480_21);
nand \U$21467 ( \21720 , \21718 , \21719 );
and \U$21468 ( \21721 , \21720 , \9902 );
not \U$21469 ( \21722 , \21720 );
and \U$21470 ( \21723 , \21722 , \9903 );
nor \U$21471 ( \21724 , \21721 , \21723 );
not \U$21472 ( \21725 , \21724 );
not \U$21473 ( \21726 , \21725 );
and \U$21474 ( \21727 , \13049 , RIbe28408_20);
and \U$21475 ( \21728 , \13669 , RIbe28390_19);
nor \U$21476 ( \21729 , \21727 , \21728 );
and \U$21477 ( \21730 , \21729 , \12195 );
not \U$21478 ( \21731 , \21729 );
and \U$21479 ( \21732 , \21731 , \12956 );
nor \U$21480 ( \21733 , \21730 , \21732 );
not \U$21481 ( \21734 , \21733 );
not \U$21482 ( \21735 , \21734 );
or \U$21483 ( \21736 , \21726 , \21735 );
nand \U$21484 ( \21737 , \21733 , \21724 );
nand \U$21485 ( \21738 , \21736 , \21737 );
and \U$21486 ( \21739 , \13478 , RIbe28660_25);
and \U$21487 ( \21740 , \13040 , RIbe285e8_24);
nor \U$21488 ( \21741 , \21739 , \21740 );
and \U$21489 ( \21742 , \21741 , \8077 );
not \U$21490 ( \21743 , \21741 );
and \U$21491 ( \21744 , \21743 , \13384 );
nor \U$21492 ( \21745 , \21742 , \21744 );
xor \U$21493 ( \21746 , \21738 , \21745 );
xnor \U$21494 ( \21747 , \21715 , \21746 );
not \U$21495 ( \21748 , \21747 );
and \U$21496 ( \21749 , \21659 , \21748 );
not \U$21497 ( \21750 , \21659 );
and \U$21498 ( \21751 , \21750 , \21747 );
nor \U$21499 ( \21752 , \21749 , \21751 );
nand \U$21500 ( \21753 , \21453 , \21752 );
not \U$21501 ( \21754 , \21451 );
not \U$21502 ( \21755 , \21369 );
nand \U$21503 ( \21756 , \21754 , \21755 );
nand \U$21504 ( \21757 , \21753 , \21756 );
not \U$21505 ( \21758 , \21757 );
not \U$21506 ( \21759 , \21758 );
or \U$21507 ( \21760 , \21278 , \21759 );
not \U$21508 ( \21761 , \21277 );
nand \U$21509 ( \21762 , \21761 , \21757 );
nand \U$21510 ( \21763 , \21760 , \21762 );
not \U$21511 ( \21764 , \21391 );
not \U$21512 ( \21765 , \21377 );
or \U$21513 ( \21766 , \21764 , \21765 );
nand \U$21514 ( \21767 , \21766 , \21383 );
not \U$21515 ( \21768 , \21377 );
nand \U$21516 ( \21769 , \21768 , \21394 );
nand \U$21517 ( \21770 , \21767 , \21769 );
not \U$21518 ( \21771 , \21770 );
not \U$21519 ( \21772 , \21431 );
not \U$21520 ( \21773 , \21438 );
or \U$21521 ( \21774 , \21772 , \21773 );
nand \U$21522 ( \21775 , \21774 , \21445 );
not \U$21523 ( \21776 , \21431 );
nand \U$21524 ( \21777 , \21776 , \21437 );
nand \U$21525 ( \21778 , \21775 , \21777 );
not \U$21526 ( \21779 , \21778 );
not \U$21527 ( \21780 , \21779 );
or \U$21528 ( \21781 , \21771 , \21780 );
not \U$21529 ( \21782 , \21770 );
nand \U$21530 ( \21783 , \21778 , \21782 );
nand \U$21531 ( \21784 , \21781 , \21783 );
not \U$21532 ( \21785 , \21412 );
not \U$21533 ( \21786 , \21422 );
not \U$21534 ( \21787 , \21786 );
or \U$21535 ( \21788 , \21785 , \21787 );
not \U$21536 ( \21789 , \21413 );
not \U$21537 ( \21790 , \21422 );
or \U$21538 ( \21791 , \21789 , \21790 );
nand \U$21539 ( \21792 , \21791 , \21404 );
nand \U$21540 ( \21793 , \21788 , \21792 );
xor \U$21541 ( \21794 , \21784 , \21793 );
not \U$21542 ( \21795 , \21794 );
or \U$21543 ( \21796 , \21509 , \21476 );
nand \U$21544 ( \21797 , \21796 , \21540 );
nand \U$21545 ( \21798 , \21509 , \21476 );
nand \U$21546 ( \21799 , \21797 , \21798 );
not \U$21547 ( \21800 , \21799 );
not \U$21548 ( \21801 , \21622 );
not \U$21549 ( \21802 , \21655 );
or \U$21550 ( \21803 , \21801 , \21802 );
not \U$21551 ( \21804 , \21654 );
not \U$21552 ( \21805 , \21579 );
or \U$21553 ( \21806 , \21804 , \21805 );
nand \U$21554 ( \21807 , \21806 , \21619 );
nand \U$21555 ( \21808 , \21803 , \21807 );
not \U$21556 ( \21809 , \21808 );
not \U$21557 ( \21810 , \21809 );
or \U$21558 ( \21811 , \21800 , \21810 );
or \U$21559 ( \21812 , \21799 , \21809 );
nand \U$21560 ( \21813 , \21811 , \21812 );
not \U$21561 ( \21814 , \21686 );
not \U$21562 ( \21815 , \21814 );
not \U$21563 ( \21816 , \21713 );
or \U$21564 ( \21817 , \21815 , \21816 );
nand \U$21565 ( \21818 , \21817 , \21746 );
nand \U$21566 ( \21819 , \21714 , \21686 );
nand \U$21567 ( \21820 , \21818 , \21819 );
not \U$21568 ( \21821 , \21820 );
and \U$21569 ( \21822 , \21813 , \21821 );
not \U$21570 ( \21823 , \21813 );
and \U$21571 ( \21824 , \21823 , \21820 );
nor \U$21572 ( \21825 , \21822 , \21824 );
not \U$21573 ( \21826 , \21825 );
or \U$21574 ( \21827 , \21795 , \21826 );
or \U$21575 ( \21828 , \21825 , \21794 );
nand \U$21576 ( \21829 , \21827 , \21828 );
not \U$21577 ( \21830 , RIbe280c0_13);
not \U$21578 ( \21831 , \15249 );
or \U$21579 ( \21832 , \21830 , \21831 );
nand \U$21580 ( \21833 , \12794 , RIbe29830_63);
nand \U$21581 ( \21834 , \21832 , \21833 );
and \U$21582 ( \21835 , \21834 , \12995 );
not \U$21583 ( \21836 , \21834 );
and \U$21584 ( \21837 , \21836 , \12801 );
nor \U$21585 ( \21838 , \21835 , \21837 );
not \U$21586 ( \21839 , RIbe296c8_60);
not \U$21587 ( \21840 , \12811 );
or \U$21588 ( \21841 , \21839 , \21840 );
nand \U$21589 ( \21842 , RIbe29650_59, RIbe2ae38_110);
nand \U$21590 ( \21843 , \21841 , \21842 );
xnor \U$21591 ( \21844 , \21843 , RIbe2aeb0_111);
not \U$21592 ( \21845 , \21844 );
and \U$21593 ( \21846 , \21845 , \564 );
not \U$21594 ( \21847 , \21845 );
and \U$21595 ( \21848 , \21847 , \1621 );
nor \U$21596 ( \21849 , \21846 , \21848 );
xor \U$21597 ( \21850 , \21838 , \21849 );
and \U$21598 ( \21851 , \21196 , RIbe285e8_24);
and \U$21599 ( \21852 , \9913 , RIbe287c8_28);
nor \U$21600 ( \21853 , \21851 , \21852 );
and \U$21601 ( \21854 , \21853 , \13383 );
not \U$21602 ( \21855 , \21853 );
and \U$21603 ( \21856 , \21855 , \16994 );
nor \U$21604 ( \21857 , \21854 , \21856 );
not \U$21605 ( \21858 , RIbe27e68_8);
not \U$21606 ( \21859 , \7974 );
or \U$21607 ( \21860 , \21858 , \21859 );
nand \U$21608 ( \21861 , \9891 , RIbe28660_25);
nand \U$21609 ( \21862 , \21860 , \21861 );
not \U$21610 ( \21863 , \21862 );
not \U$21611 ( \21864 , \7984 );
and \U$21612 ( \21865 , \21863 , \21864 );
and \U$21613 ( \21866 , \21862 , \6948 );
nor \U$21614 ( \21867 , \21865 , \21866 );
and \U$21615 ( \21868 , \21857 , \21867 );
not \U$21616 ( \21869 , \21857 );
not \U$21617 ( \21870 , \21867 );
and \U$21618 ( \21871 , \21869 , \21870 );
or \U$21619 ( \21872 , \21868 , \21871 );
and \U$21620 ( \21873 , \6980 , RIbe27fd0_11);
and \U$21621 ( \21874 , \10898 , RIbe27f58_10);
nor \U$21622 ( \21875 , \21873 , \21874 );
and \U$21623 ( \21876 , \21875 , \6992 );
not \U$21624 ( \21877 , \21875 );
and \U$21625 ( \21878 , \21877 , \13227 );
nor \U$21626 ( \21879 , \21876 , \21878 );
and \U$21627 ( \21880 , \21872 , \21879 );
not \U$21628 ( \21881 , \21872 );
not \U$21629 ( \21882 , \21879 );
and \U$21630 ( \21883 , \21881 , \21882 );
nor \U$21631 ( \21884 , \21880 , \21883 );
buf \U$21632 ( \21885 , \21884 );
xor \U$21633 ( \21886 , \21850 , \21885 );
not \U$21634 ( \21887 , \13085 );
not \U$21635 ( \21888 , \5423 );
and \U$21636 ( \21889 , \21887 , \21888 );
and \U$21637 ( \21890 , \12764 , RIbe28b88_36);
nor \U$21638 ( \21891 , \21889 , \21890 );
and \U$21639 ( \21892 , \21891 , \12774 );
not \U$21640 ( \21893 , \21891 );
and \U$21641 ( \21894 , \21893 , \12924 );
nor \U$21642 ( \21895 , \21892 , \21894 );
not \U$21643 ( \21896 , RIbe28390_19);
not \U$21644 ( \21897 , \12942 );
or \U$21645 ( \21898 , \21896 , \21897 );
nand \U$21646 ( \21899 , \15628 , RIbe28b10_35);
nand \U$21647 ( \21900 , \21898 , \21899 );
not \U$21648 ( \21901 , \21900 );
not \U$21649 ( \21902 , \12957 );
and \U$21650 ( \21903 , \21901 , \21902 );
and \U$21651 ( \21904 , \21900 , \17005 );
nor \U$21652 ( \21905 , \21903 , \21904 );
xor \U$21653 ( \21906 , \21895 , \21905 );
not \U$21654 ( \21907 , RIbe28480_21);
not \U$21655 ( \21908 , \13024 );
or \U$21656 ( \21909 , \21907 , \21908 );
nand \U$21657 ( \21910 , \14511 , RIbe28408_20);
nand \U$21658 ( \21911 , \21909 , \21910 );
not \U$21659 ( \21912 , \21911 );
not \U$21660 ( \21913 , \13033 );
and \U$21661 ( \21914 , \21912 , \21913 );
and \U$21662 ( \21915 , \21911 , \10943 );
nor \U$21663 ( \21916 , \21914 , \21915 );
xnor \U$21664 ( \21917 , \21906 , \21916 );
not \U$21665 ( \21918 , RIbe28228_16);
not \U$21666 ( \21919 , \14550 );
or \U$21667 ( \21920 , \21918 , \21919 );
not \U$21668 ( \21921 , \3663 );
nand \U$21669 ( \21922 , \21921 , \13012 );
nand \U$21670 ( \21923 , \21920 , \21922 );
and \U$21671 ( \21924 , \21923 , \20602 );
not \U$21672 ( \21925 , \21923 );
and \U$21673 ( \21926 , \21925 , \16366 );
nor \U$21674 ( \21927 , \21924 , \21926 );
not \U$21675 ( \21928 , \21927 );
not \U$21676 ( \21929 , \21928 );
not \U$21677 ( \21930 , RIbe28930_31);
not \U$21678 ( \21931 , \14534 );
or \U$21679 ( \21932 , \21930 , \21931 );
nand \U$21680 ( \21933 , \12735 , RIbe29560_57);
nand \U$21681 ( \21934 , \21932 , \21933 );
and \U$21682 ( \21935 , \21934 , \14543 );
not \U$21683 ( \21936 , \21934 );
and \U$21684 ( \21937 , \21936 , \21013 );
nor \U$21685 ( \21938 , \21935 , \21937 );
not \U$21686 ( \21939 , \21938 );
not \U$21687 ( \21940 , \21939 );
or \U$21688 ( \21941 , \21929 , \21940 );
nand \U$21689 ( \21942 , \21938 , \21927 );
nand \U$21690 ( \21943 , \21941 , \21942 );
not \U$21691 ( \21944 , RIbe28a20_33);
not \U$21692 ( \21945 , \19262 );
or \U$21693 ( \21946 , \21944 , \21945 );
nand \U$21694 ( \21947 , \12710 , RIbe289a8_32);
nand \U$21695 ( \21948 , \21946 , \21947 );
xor \U$21696 ( \21949 , \21948 , \12723 );
xnor \U$21697 ( \21950 , \21943 , \21949 );
xor \U$21698 ( \21951 , \21917 , \21950 );
xnor \U$21699 ( \21952 , \21886 , \21951 );
not \U$21700 ( \21953 , RIbe2a550_91);
not \U$21701 ( \21954 , \20625 );
or \U$21702 ( \21955 , \21953 , \21954 );
nand \U$21703 ( \21956 , \6787 , RIbe2a988_100);
nand \U$21704 ( \21957 , \21955 , \21956 );
and \U$21705 ( \21958 , \21957 , \3471 );
not \U$21706 ( \21959 , \21957 );
and \U$21707 ( \21960 , \21959 , \3698 );
nor \U$21708 ( \21961 , \21958 , \21960 );
not \U$21709 ( \21962 , \21961 );
not \U$21710 ( \21963 , \21962 );
not \U$21711 ( \21964 , RIbe2a910_99);
not \U$21712 ( \21965 , \4595 );
or \U$21713 ( \21966 , \21964 , \21965 );
nand \U$21714 ( \21967 , \7858 , RIbe2b5b8_126);
nand \U$21715 ( \21968 , \21966 , \21967 );
and \U$21716 ( \21969 , \21968 , \7865 );
not \U$21717 ( \21970 , \21968 );
and \U$21718 ( \21971 , \21970 , \4007 );
nor \U$21719 ( \21972 , \21969 , \21971 );
not \U$21720 ( \21973 , \21972 );
not \U$21721 ( \21974 , \21973 );
or \U$21722 ( \21975 , \21963 , \21974 );
nand \U$21723 ( \21976 , \21961 , \21972 );
nand \U$21724 ( \21977 , \21975 , \21976 );
not \U$21725 ( \21978 , RIbe2a190_83);
not \U$21726 ( \21979 , \6797 );
or \U$21727 ( \21980 , \21978 , \21979 );
nand \U$21728 ( \21981 , \6800 , RIbe2a5c8_92);
nand \U$21729 ( \21982 , \21980 , \21981 );
and \U$21730 ( \21983 , \21982 , \2887 );
not \U$21731 ( \21984 , \21982 );
and \U$21732 ( \21985 , \21984 , \3290 );
nor \U$21733 ( \21986 , \21983 , \21985 );
and \U$21734 ( \21987 , \21977 , \21986 );
not \U$21735 ( \21988 , \21977 );
not \U$21736 ( \21989 , \21986 );
and \U$21737 ( \21990 , \21988 , \21989 );
nor \U$21738 ( \21991 , \21987 , \21990 );
not \U$21739 ( \21992 , \21090 );
not \U$21740 ( \21993 , RIbe2a028_80);
not \U$21741 ( \21994 , \21081 );
or \U$21742 ( \21995 , \21993 , \21994 );
nand \U$21743 ( \21996 , \8235 , RIbe29fb0_79);
nand \U$21744 ( \21997 , \21995 , \21996 );
not \U$21745 ( \21998 , \21997 );
or \U$21746 ( \21999 , \21992 , \21998 );
or \U$21747 ( \22000 , \5740 , \21997 );
nand \U$21748 ( \22001 , \21999 , \22000 );
not \U$21749 ( \22002 , RIbe2a2f8_86);
not \U$21750 ( \22003 , \15313 );
or \U$21751 ( \22004 , \22002 , \22003 );
nand \U$21752 ( \22005 , \15885 , RIbe2acd0_107);
nand \U$21753 ( \22006 , \22004 , \22005 );
not \U$21754 ( \22007 , \5754 );
and \U$21755 ( \22008 , \22006 , \22007 );
not \U$21756 ( \22009 , \22006 );
and \U$21757 ( \22010 , \22009 , \6640 );
nor \U$21758 ( \22011 , \22008 , \22010 );
xor \U$21759 ( \22012 , \22001 , \22011 );
not \U$21760 ( \22013 , RIbe2a3e8_88);
not \U$21761 ( \22014 , \6427 );
or \U$21762 ( \22015 , \22013 , \22014 );
nand \U$21763 ( \22016 , \7056 , RIbe2a370_87);
nand \U$21764 ( \22017 , \22015 , \22016 );
and \U$21765 ( \22018 , \22017 , \4586 );
not \U$21766 ( \22019 , \22017 );
and \U$21767 ( \22020 , \22019 , \4592 );
nor \U$21768 ( \22021 , \22018 , \22020 );
xor \U$21769 ( \22022 , \22012 , \22021 );
xor \U$21770 ( \22023 , \21991 , \22022 );
not \U$21771 ( \22024 , RIbe29c68_72);
not \U$21772 ( \22025 , \7941 );
or \U$21773 ( \22026 , \22024 , \22025 );
nand \U$21774 ( \22027 , \6596 , RIbe29bf0_71);
nand \U$21775 ( \22028 , \22026 , \22027 );
and \U$21776 ( \22029 , \22028 , \6601 );
not \U$21777 ( \22030 , \22028 );
and \U$21778 ( \22031 , \22030 , \6602 );
nor \U$21779 ( \22032 , \22029 , \22031 );
not \U$21780 ( \22033 , RIbe28f48_44);
not \U$21781 ( \22034 , \7954 );
or \U$21782 ( \22035 , \22033 , \22034 );
nand \U$21783 ( \22036 , \7958 , RIbe28ed0_43);
nand \U$21784 ( \22037 , \22035 , \22036 );
and \U$21785 ( \22038 , \22037 , \6572 );
not \U$21786 ( \22039 , \22037 );
and \U$21787 ( \22040 , \22039 , \7293 );
nor \U$21788 ( \22041 , \22038 , \22040 );
and \U$21789 ( \22042 , \22032 , \22041 );
not \U$21790 ( \22043 , \22032 );
not \U$21791 ( \22044 , \22041 );
and \U$21792 ( \22045 , \22043 , \22044 );
nor \U$21793 ( \22046 , \22042 , \22045 );
not \U$21794 ( \22047 , RIbe29e48_76);
not \U$21795 ( \22048 , \6536 );
or \U$21796 ( \22049 , \22047 , \22048 );
nand \U$21797 ( \22050 , \7076 , RIbe29dd0_75);
nand \U$21798 ( \22051 , \22049 , \22050 );
and \U$21799 ( \22052 , \22051 , \7935 );
not \U$21800 ( \22053 , \22051 );
and \U$21801 ( \22054 , \22053 , \6891 );
nor \U$21802 ( \22055 , \22052 , \22054 );
xor \U$21803 ( \22056 , \22046 , \22055 );
xnor \U$21804 ( \22057 , \22023 , \22056 );
xnor \U$21805 ( \22058 , \21952 , \22057 );
and \U$21806 ( \22059 , \21829 , \22058 );
not \U$21807 ( \22060 , \21829 );
not \U$21808 ( \22061 , \22058 );
and \U$21809 ( \22062 , \22060 , \22061 );
nor \U$21810 ( \22063 , \22059 , \22062 );
and \U$21811 ( \22064 , \21763 , \22063 );
not \U$21812 ( \22065 , \21763 );
not \U$21813 ( \22066 , \22063 );
and \U$21814 ( \22067 , \22065 , \22066 );
nor \U$21815 ( \22068 , \22064 , \22067 );
not \U$21816 ( \22069 , \22068 );
not \U$21817 ( \22070 , \22069 );
not \U$21818 ( \22071 , \22070 );
not \U$21819 ( \22072 , \21747 );
not \U$21820 ( \22073 , \21656 );
not \U$21821 ( \22074 , \22073 );
or \U$21822 ( \22075 , \22072 , \22074 );
not \U$21823 ( \22076 , \21541 );
nand \U$21824 ( \22077 , \22075 , \22076 );
not \U$21825 ( \22078 , \22073 );
nand \U$21826 ( \22079 , \22078 , \21748 );
nand \U$21827 ( \22080 , \22077 , \22079 );
not \U$21828 ( \22081 , \21301 );
not \U$21829 ( \22082 , \21286 );
or \U$21830 ( \22083 , \22081 , \22082 );
nand \U$21831 ( \22084 , \22083 , \21292 );
or \U$21832 ( \22085 , \21286 , \21301 );
nand \U$21833 ( \22086 , \22084 , \22085 );
xor \U$21834 ( \22087 , \21311 , \21317 );
and \U$21835 ( \22088 , \22087 , \21322 );
and \U$21836 ( \22089 , \21311 , \21317 );
or \U$21837 ( \22090 , \22088 , \22089 );
nor \U$21838 ( \22091 , \22086 , \22090 );
xor \U$21839 ( \22092 , \21330 , \21334 );
and \U$21840 ( \22093 , \22092 , \21364 );
and \U$21841 ( \22094 , \21330 , \21334 );
or \U$21842 ( \22095 , \22093 , \22094 );
or \U$21843 ( \22096 , \22091 , \22095 );
nand \U$21844 ( \22097 , \22086 , \22090 );
nand \U$21845 ( \22098 , \22096 , \22097 );
not \U$21846 ( \22099 , \22098 );
not \U$21847 ( \22100 , \21078 );
not \U$21848 ( \22101 , \22100 );
not \U$21849 ( \22102 , \21118 );
or \U$21850 ( \22103 , \22101 , \22102 );
nand \U$21851 ( \22104 , \22103 , \21153 );
or \U$21852 ( \22105 , \21118 , \22100 );
and \U$21853 ( \22106 , \22104 , \22105 );
nand \U$21854 ( \22107 , \21035 , \21005 );
and \U$21855 ( \22108 , \22106 , \22107 );
and \U$21856 ( \22109 , \21226 , \21264 );
nor \U$21857 ( \22110 , \22109 , \21193 );
nor \U$21858 ( \22111 , \21226 , \21264 );
nor \U$21859 ( \22112 , \22110 , \22111 );
nor \U$21860 ( \22113 , \22108 , \22112 );
nor \U$21861 ( \22114 , \22106 , \22107 );
nor \U$21862 ( \22115 , \22113 , \22114 );
not \U$21863 ( \22116 , \22115 );
or \U$21864 ( \22117 , \22099 , \22116 );
or \U$21865 ( \22118 , \22115 , \22098 );
nand \U$21866 ( \22119 , \22117 , \22118 );
not \U$21867 ( \22120 , \22119 );
and \U$21868 ( \22121 , \22080 , \22120 );
not \U$21869 ( \22122 , \22080 );
and \U$21870 ( \22123 , \22122 , \22119 );
or \U$21871 ( \22124 , \22121 , \22123 );
not \U$21872 ( \22125 , \22124 );
or \U$21873 ( \22126 , \22071 , \22125 );
not \U$21874 ( \22127 , \21613 );
not \U$21875 ( \22128 , \21600 );
or \U$21876 ( \22129 , \22127 , \22128 );
nand \U$21877 ( \22130 , \22129 , \21590 );
not \U$21878 ( \22131 , \21600 );
nand \U$21879 ( \22132 , \22131 , \21616 );
nand \U$21880 ( \22133 , \22130 , \22132 );
not \U$21881 ( \22134 , \22133 );
not \U$21882 ( \22135 , \22134 );
nand \U$21883 ( \22136 , \21574 , \21551 );
and \U$21884 ( \22137 , \22136 , \21561 );
nor \U$21885 ( \22138 , \21574 , \21551 );
nor \U$21886 ( \22139 , \22137 , \22138 );
not \U$21887 ( \22140 , \22139 );
not \U$21888 ( \22141 , \22140 );
or \U$21889 ( \22142 , \22135 , \22141 );
nand \U$21890 ( \22143 , \22139 , \22133 );
nand \U$21891 ( \22144 , \22142 , \22143 );
xor \U$21892 ( \22145 , \21633 , \21643 );
and \U$21893 ( \22146 , \22145 , \21653 );
and \U$21894 ( \22147 , \21633 , \21643 );
or \U$21895 ( \22148 , \22146 , \22147 );
not \U$21896 ( \22149 , \22148 );
and \U$21897 ( \22150 , \22144 , \22149 );
not \U$21898 ( \22151 , \22144 );
and \U$21899 ( \22152 , \22151 , \22148 );
nor \U$21900 ( \22153 , \22150 , \22152 );
not \U$21901 ( \22154 , \22153 );
nand \U$21902 ( \22155 , \21529 , \21539 );
not \U$21903 ( \22156 , \21520 );
and \U$21904 ( \22157 , \22155 , \22156 );
nor \U$21905 ( \22158 , \21529 , \21539 );
nor \U$21906 ( \22159 , \22157 , \22158 );
xor \U$21907 ( \22160 , \21487 , \21498 );
and \U$21908 ( \22161 , \22160 , \21508 );
and \U$21909 ( \22162 , \21487 , \21498 );
or \U$21910 ( \22163 , \22161 , \22162 );
xor \U$21911 ( \22164 , \22159 , \22163 );
nand \U$21912 ( \22165 , \21474 , \21462 );
xnor \U$21913 ( \22166 , \22164 , \22165 );
not \U$21914 ( \22167 , \22166 );
or \U$21915 ( \22168 , \22154 , \22167 );
or \U$21916 ( \22169 , \22153 , \22166 );
nand \U$21917 ( \22170 , \22168 , \22169 );
nand \U$21918 ( \22171 , \1179 , RIbe2ab68_104);
and \U$21919 ( \22172 , \22171 , \1621 );
not \U$21920 ( \22173 , \22171 );
and \U$21921 ( \22174 , \22173 , \564 );
or \U$21922 ( \22175 , \22172 , \22174 );
not \U$21923 ( \22176 , RIbe2af28_112);
not \U$21924 ( \22177 , \1631 );
or \U$21925 ( \22178 , \22176 , \22177 );
nand \U$21926 ( \22179 , \1098 , RIbe2b1f8_118);
nand \U$21927 ( \22180 , \22178 , \22179 );
and \U$21928 ( \22181 , \22180 , \1309 );
not \U$21929 ( \22182 , \22180 );
and \U$21930 ( \22183 , \22182 , \2418 );
nor \U$21931 ( \22184 , \22181 , \22183 );
not \U$21932 ( \22185 , RIbe2b018_114);
not \U$21933 ( \22186 , \21344 );
or \U$21934 ( \22187 , \22185 , \22186 );
nand \U$21935 ( \22188 , \1146 , RIbe2afa0_113);
nand \U$21936 ( \22189 , \22187 , \22188 );
and \U$21937 ( \22190 , \22189 , \1153 );
not \U$21938 ( \22191 , \22189 );
and \U$21939 ( \22192 , \22191 , \7899 );
nor \U$21940 ( \22193 , \22190 , \22192 );
xor \U$21941 ( \22194 , \22184 , \22193 );
not \U$21942 ( \22195 , RIbe2aaf0_103);
not \U$21943 ( \22196 , \2424 );
or \U$21944 ( \22197 , \22195 , \22196 );
nand \U$21945 ( \22198 , \7905 , RIbe2b630_127);
nand \U$21946 ( \22199 , \22197 , \22198 );
and \U$21947 ( \22200 , \22199 , \1813 );
not \U$21948 ( \22201 , \22199 );
and \U$21949 ( \22202 , \22201 , \1010 );
nor \U$21950 ( \22203 , \22200 , \22202 );
not \U$21951 ( \22204 , \22203 );
xor \U$21952 ( \22205 , \22194 , \22204 );
xor \U$21953 ( \22206 , \22175 , \22205 );
not \U$21954 ( \22207 , RIbe2b108_116);
not \U$21955 ( \22208 , \20674 );
or \U$21956 ( \22209 , \22207 , \22208 );
nand \U$21957 ( \22210 , \2384 , RIbe2b090_115);
nand \U$21958 ( \22211 , \22209 , \22210 );
not \U$21959 ( \22212 , \22211 );
not \U$21960 ( \22213 , \3516 );
and \U$21961 ( \22214 , \22212 , \22213 );
and \U$21962 ( \22215 , \22211 , \1075 );
nor \U$21963 ( \22216 , \22214 , \22215 );
not \U$21964 ( \22217 , \22216 );
not \U$21965 ( \22218 , RIbe2a280_85);
not \U$21966 ( \22219 , \4050 );
or \U$21967 ( \22220 , \22218 , \22219 );
nand \U$21968 ( \22221 , \2900 , RIbe2a208_84);
nand \U$21969 ( \22222 , \22220 , \22221 );
and \U$21970 ( \22223 , \22222 , \4058 );
not \U$21971 ( \22224 , \22222 );
and \U$21972 ( \22225 , \22224 , \3275 );
nor \U$21973 ( \22226 , \22223 , \22225 );
not \U$21974 ( \22227 , \22226 );
or \U$21975 ( \22228 , \22217 , \22227 );
or \U$21976 ( \22229 , \22216 , \22226 );
nand \U$21977 ( \22230 , \22228 , \22229 );
and \U$21978 ( \22231 , \1113 , RIbe2b180_117);
and \U$21979 ( \22232 , \20664 , RIbe2b270_119);
nor \U$21980 ( \22233 , \22231 , \22232 );
and \U$21981 ( \22234 , \22233 , \1132 );
not \U$21982 ( \22235 , \22233 );
and \U$21983 ( \22236 , \22235 , \1448 );
nor \U$21984 ( \22237 , \22234 , \22236 );
xnor \U$21985 ( \22238 , \22230 , \22237 );
xor \U$21986 ( \22239 , \22206 , \22238 );
xnor \U$21987 ( \22240 , \22170 , \22239 );
not \U$21988 ( \22241 , \22240 );
xor \U$21989 ( \22242 , \21396 , \21426 );
and \U$21990 ( \22243 , \22242 , \21450 );
and \U$21991 ( \22244 , \21396 , \21426 );
or \U$21992 ( \22245 , \22243 , \22244 );
xor \U$21993 ( \22246 , \21695 , \21701 );
and \U$21994 ( \22247 , \22246 , \21712 );
and \U$21995 ( \22248 , \21695 , \21701 );
or \U$21996 ( \22249 , \22247 , \22248 );
not \U$21997 ( \22250 , \21745 );
not \U$21998 ( \22251 , \21724 );
or \U$21999 ( \22252 , \22250 , \22251 );
or \U$22000 ( \22253 , \21724 , \21745 );
nand \U$22001 ( \22254 , \22253 , \21734 );
nand \U$22002 ( \22255 , \22252 , \22254 );
xor \U$22003 ( \22256 , \22249 , \22255 );
or \U$22004 ( \22257 , \21674 , \21665 );
and \U$22005 ( \22258 , \21685 , \22257 );
and \U$22006 ( \22259 , \21665 , \21674 );
nor \U$22007 ( \22260 , \22258 , \22259 );
xnor \U$22008 ( \22261 , \22256 , \22260 );
xnor \U$22009 ( \22262 , \22245 , \22261 );
not \U$22010 ( \22263 , \22262 );
or \U$22011 ( \22264 , \22241 , \22263 );
or \U$22012 ( \22265 , \22262 , \22240 );
nand \U$22013 ( \22266 , \22264 , \22265 );
not \U$22014 ( \22267 , \22266 );
xor \U$22015 ( \22268 , \1153 , \20559 );
xnor \U$22016 ( \22269 , \22268 , \20571 );
not \U$22017 ( \22270 , \22269 );
not \U$22018 ( \22271 , \20526 );
not \U$22019 ( \22272 , \20550 );
or \U$22020 ( \22273 , \22271 , \22272 );
or \U$22021 ( \22274 , \20526 , \20550 );
nand \U$22022 ( \22275 , \22273 , \22274 );
not \U$22023 ( \22276 , \22275 );
not \U$22024 ( \22277 , \20538 );
and \U$22025 ( \22278 , \22276 , \22277 );
and \U$22026 ( \22279 , \22275 , \20538 );
nor \U$22027 ( \22280 , \22278 , \22279 );
nand \U$22028 ( \22281 , \22270 , \22280 );
and \U$22029 ( \22282 , \20606 , \20594 );
not \U$22030 ( \22283 , \20606 );
and \U$22031 ( \22284 , \22283 , \20595 );
or \U$22032 ( \22285 , \22282 , \22284 );
xor \U$22033 ( \22286 , \22285 , \20585 );
and \U$22034 ( \22287 , \22281 , \22286 );
not \U$22035 ( \22288 , \22269 );
nor \U$22036 ( \22289 , \22288 , \22280 );
nor \U$22037 ( \22290 , \22287 , \22289 );
buf \U$22038 ( \22291 , \22290 );
not \U$22039 ( \22292 , \22291 );
xor \U$22040 ( \22293 , \20448 , \20458 );
xor \U$22041 ( \22294 , \22293 , \20469 );
not \U$22042 ( \22295 , \22294 );
and \U$22043 ( \22296 , \20412 , \20422 );
not \U$22044 ( \22297 , \20412 );
and \U$22045 ( \22298 , \22297 , \20423 );
or \U$22046 ( \22299 , \22296 , \22298 );
not \U$22047 ( \22300 , \20433 );
and \U$22048 ( \22301 , \22299 , \22300 );
not \U$22049 ( \22302 , \22299 );
and \U$22050 ( \22303 , \22302 , \20433 );
nor \U$22051 ( \22304 , \22301 , \22303 );
not \U$22052 ( \22305 , \22304 );
or \U$22053 ( \22306 , \22295 , \22305 );
xor \U$22054 ( \22307 , \20495 , \20483 );
xnor \U$22055 ( \22308 , \22307 , \20506 );
nand \U$22056 ( \22309 , \22306 , \22308 );
not \U$22057 ( \22310 , \22304 );
not \U$22058 ( \22311 , \22294 );
nand \U$22059 ( \22312 , \22310 , \22311 );
nand \U$22060 ( \22313 , \22309 , \22312 );
nand \U$22061 ( \22314 , \22292 , \22313 );
not \U$22062 ( \22315 , RIbe29fb0_79);
not \U$22063 ( \22316 , \8199 );
or \U$22064 ( \22317 , \22315 , \22316 );
nand \U$22065 ( \22318 , \7958 , RIbe29e48_76);
nand \U$22066 ( \22319 , \22317 , \22318 );
xor \U$22067 ( \22320 , \22319 , \6572 );
not \U$22068 ( \22321 , \22320 );
not \U$22069 ( \22322 , \22321 );
not \U$22070 ( \22323 , RIbe29bf0_71);
not \U$22071 ( \22324 , \6942 );
or \U$22072 ( \22325 , \22323 , \22324 );
nand \U$22073 ( \22326 , RIbe28f48_44, \13158 );
nand \U$22074 ( \22327 , \22325 , \22326 );
and \U$22075 ( \22328 , \22327 , \16010 );
not \U$22076 ( \22329 , \22327 );
and \U$22077 ( \22330 , \22329 , \6948 );
nor \U$22078 ( \22331 , \22328 , \22330 );
not \U$22079 ( \22332 , \22331 );
or \U$22080 ( \22333 , \22322 , \22332 );
not \U$22081 ( \22334 , \22331 );
not \U$22082 ( \22335 , \22334 );
not \U$22083 ( \22336 , \22320 );
or \U$22084 ( \22337 , \22335 , \22336 );
not \U$22085 ( \22338 , RIbe29dd0_75);
not \U$22086 ( \22339 , \7298 );
or \U$22087 ( \22340 , \22338 , \22339 );
nand \U$22088 ( \22341 , \13792 , RIbe29c68_72);
nand \U$22089 ( \22342 , \22340 , \22341 );
not \U$22090 ( \22343 , \22342 );
not \U$22091 ( \22344 , \6992 );
and \U$22092 ( \22345 , \22343 , \22344 );
and \U$22093 ( \22346 , \22342 , \6992 );
nor \U$22094 ( \22347 , \22345 , \22346 );
not \U$22095 ( \22348 , \22347 );
nand \U$22096 ( \22349 , \22337 , \22348 );
nand \U$22097 ( \22350 , \22333 , \22349 );
not \U$22098 ( \22351 , RIbe2a208_84);
not \U$22099 ( \22352 , \4317 );
or \U$22100 ( \22353 , \22351 , \22352 );
not \U$22101 ( \22354 , \14285 );
nand \U$22102 ( \22355 , \22354 , \7858 );
nand \U$22103 ( \22356 , \22353 , \22355 );
and \U$22104 ( \22357 , \22356 , \7865 );
not \U$22105 ( \22358 , \22356 );
and \U$22106 ( \22359 , \22358 , \4603 );
nor \U$22107 ( \22360 , \22357 , \22359 );
not \U$22108 ( \22361 , \22360 );
not \U$22109 ( \22362 , RIbe2a988_100);
not \U$22110 ( \22363 , \15313 );
or \U$22111 ( \22364 , \22362 , \22363 );
nand \U$22112 ( \22365 , \5749 , RIbe2a910_99);
nand \U$22113 ( \22366 , \22364 , \22365 );
not \U$22114 ( \22367 , \22366 );
not \U$22115 ( \22368 , \5046 );
and \U$22116 ( \22369 , \22367 , \22368 );
and \U$22117 ( \22370 , \22366 , \10984 );
nor \U$22118 ( \22371 , \22369 , \22370 );
not \U$22119 ( \22372 , \22371 );
or \U$22120 ( \22373 , \22361 , \22372 );
not \U$22121 ( \22374 , RIbe2a5c8_92);
not \U$22122 ( \22375 , \21097 );
or \U$22123 ( \22376 , \22374 , \22375 );
buf \U$22124 ( \22377 , \5051 );
not \U$22125 ( \22378 , \22377 );
nand \U$22126 ( \22379 , \22378 , RIbe2a550_91);
nand \U$22127 ( \22380 , \22376 , \22379 );
and \U$22128 ( \22381 , \22380 , \4586 );
not \U$22129 ( \22382 , \22380 );
and \U$22130 ( \22383 , \22382 , \4592 );
nor \U$22131 ( \22384 , \22381 , \22383 );
nand \U$22132 ( \22385 , \22373 , \22384 );
or \U$22133 ( \22386 , \22371 , \22360 );
and \U$22134 ( \22387 , \22385 , \22386 );
not \U$22135 ( \22388 , RIbe2b5b8_126);
not \U$22136 ( \22389 , \6138 );
or \U$22137 ( \22390 , \22388 , \22389 );
nand \U$22138 ( \22391 , RIbe2a3e8_88, \6616 );
nand \U$22139 ( \22392 , \22390 , \22391 );
and \U$22140 ( \22393 , \22392 , \9944 );
not \U$22141 ( \22394 , \22392 );
and \U$22142 ( \22395 , \22394 , \10969 );
nor \U$22143 ( \22396 , \22393 , \22395 );
nand \U$22144 ( \22397 , \6588 , RIbe2acd0_107);
or \U$22145 ( \22398 , \22397 , \6595 );
nand \U$22146 ( \22399 , \7277 , RIbe2a028_80);
nand \U$22147 ( \22400 , \22398 , \22399 );
not \U$22148 ( \22401 , \22400 );
not \U$22149 ( \22402 , \7271 );
and \U$22150 ( \22403 , \22401 , \22402 );
and \U$22151 ( \22404 , \22400 , \9868 );
nor \U$22152 ( \22405 , \22403 , \22404 );
nand \U$22153 ( \22406 , \22396 , \22405 );
not \U$22154 ( \22407 , RIbe2a370_87);
not \U$22155 ( \22408 , \6535 );
or \U$22156 ( \22409 , \22407 , \22408 );
nand \U$22157 ( \22410 , RIbe2a2f8_86, \6540 );
nand \U$22158 ( \22411 , \22409 , \22410 );
and \U$22159 ( \22412 , \22411 , \6546 );
not \U$22160 ( \22413 , \22411 );
and \U$22161 ( \22414 , \22413 , \6891 );
nor \U$22162 ( \22415 , \22412 , \22414 );
and \U$22163 ( \22416 , \22406 , \22415 );
nor \U$22164 ( \22417 , \22396 , \22405 );
nor \U$22165 ( \22418 , \22416 , \22417 );
nand \U$22166 ( \22419 , \22387 , \22418 );
and \U$22167 ( \22420 , \22350 , \22419 );
nor \U$22168 ( \22421 , \22387 , \22418 );
nor \U$22169 ( \22422 , \22420 , \22421 );
not \U$22170 ( \22423 , RIbe2aaf0_103);
not \U$22171 ( \22424 , \1633 );
or \U$22172 ( \22425 , \22423 , \22424 );
nand \U$22173 ( \22426 , \1099 , RIbe2b630_127);
nand \U$22174 ( \22427 , \22425 , \22426 );
and \U$22175 ( \22428 , \22427 , \4251 );
not \U$22176 ( \22429 , \22427 );
and \U$22177 ( \22430 , \22429 , \1309 );
nor \U$22178 ( \22431 , \22428 , \22430 );
not \U$22179 ( \22432 , \22431 );
not \U$22180 ( \22433 , RIbe2b630_127);
not \U$22181 ( \22434 , \1112 );
or \U$22182 ( \22435 , \22433 , \22434 );
nand \U$22183 ( \22436 , RIbe2b018_114, \20849 );
nand \U$22184 ( \22437 , \22435 , \22436 );
not \U$22185 ( \22438 , \22437 );
not \U$22186 ( \22439 , \1123 );
and \U$22187 ( \22440 , \22438 , \22439 );
and \U$22188 ( \22441 , \22437 , \1123 );
nor \U$22189 ( \22442 , \22440 , \22441 );
not \U$22190 ( \22443 , RIbe2ab68_104);
not \U$22191 ( \22444 , \8868 );
or \U$22192 ( \22445 , \22443 , \22444 );
not \U$22193 ( \22446 , \13192 );
nand \U$22194 ( \22447 , \22446 , \1454 );
nand \U$22195 ( \22448 , \22445 , \22447 );
and \U$22196 ( \22449 , \22448 , \1082 );
not \U$22197 ( \22450 , \22448 );
and \U$22198 ( \22451 , \22450 , \1309 );
nor \U$22199 ( \22452 , \22449 , \22451 );
nand \U$22200 ( \22453 , \22442 , \22452 );
not \U$22201 ( \22454 , \4064 );
not \U$22202 ( \22455 , RIbe2af28_112);
not \U$22203 ( \22456 , \22455 );
and \U$22204 ( \22457 , \22454 , \22456 );
and \U$22205 ( \22458 , \2390 , RIbe2afa0_113);
nor \U$22206 ( \22459 , \22457 , \22458 );
and \U$22207 ( \22460 , \22459 , \1076 );
not \U$22208 ( \22461 , \22459 );
and \U$22209 ( \22462 , \22461 , \9083 );
nor \U$22210 ( \22463 , \22460 , \22462 );
and \U$22211 ( \22464 , \22453 , \22463 );
nor \U$22212 ( \22465 , \22442 , \22452 );
nor \U$22213 ( \22466 , \22464 , \22465 );
not \U$22214 ( \22467 , \22466 );
or \U$22215 ( \22468 , \22432 , \22467 );
nand \U$22216 ( \22469 , \3701 , RIbe2b090_115);
or \U$22217 ( \22470 , \22469 , \20767 );
nand \U$22218 ( \22471 , RIbe2a280_85, \6787 );
nand \U$22219 ( \22472 , \22470 , \22471 );
xor \U$22220 ( \22473 , \22472 , \3448 );
not \U$22221 ( \22474 , \22473 );
not \U$22222 ( \22475 , RIbe2b1f8_118);
not \U$22223 ( \22476 , \7827 );
or \U$22224 ( \22477 , \22475 , \22476 );
nand \U$22225 ( \22478 , \3267 , RIbe2b180_117);
nand \U$22226 ( \22479 , \22477 , \22478 );
and \U$22227 ( \22480 , \22479 , \4783 );
not \U$22228 ( \22481 , \22479 );
and \U$22229 ( \22482 , \22481 , \4287 );
nor \U$22230 ( \22483 , \22480 , \22482 );
not \U$22231 ( \22484 , \22483 );
or \U$22232 ( \22485 , \22474 , \22484 );
not \U$22233 ( \22486 , \2887 );
and \U$22234 ( \22487 , \3456 , RIbe2b108_116);
not \U$22235 ( \22488 , \3456 );
and \U$22236 ( \22489 , \3281 , RIbe2b270_119);
and \U$22237 ( \22490 , \22488 , \22489 );
or \U$22238 ( \22491 , \22487 , \22490 );
not \U$22239 ( \22492 , \22491 );
or \U$22240 ( \22493 , \22486 , \22492 );
or \U$22241 ( \22494 , \22491 , \2887 );
nand \U$22242 ( \22495 , \22493 , \22494 );
nand \U$22243 ( \22496 , \22485 , \22495 );
or \U$22244 ( \22497 , \22483 , \22473 );
nand \U$22245 ( \22498 , \22496 , \22497 );
nand \U$22246 ( \22499 , \22468 , \22498 );
not \U$22247 ( \22500 , \22466 );
not \U$22248 ( \22501 , \22431 );
nand \U$22249 ( \22502 , \22500 , \22501 );
and \U$22250 ( \22503 , \22499 , \22502 );
nand \U$22251 ( \22504 , \22422 , \22503 );
not \U$22252 ( \22505 , \12218 );
not \U$22253 ( \22506 , RIbe27f58_10);
not \U$22254 ( \22507 , \20530 );
or \U$22255 ( \22508 , \22506 , \22507 );
nand \U$22256 ( \22509 , \12212 , RIbe27e68_8);
nand \U$22257 ( \22510 , \22508 , \22509 );
not \U$22258 ( \22511 , \22510 );
and \U$22259 ( \22512 , \22505 , \22511 );
and \U$22260 ( \22513 , \22510 , \13661 );
nor \U$22261 ( \22514 , \22512 , \22513 );
not \U$22262 ( \22515 , RIbe28660_25);
not \U$22263 ( \22516 , \12942 );
or \U$22264 ( \22517 , \22515 , \22516 );
nand \U$22265 ( \22518 , \12947 , RIbe285e8_24);
nand \U$22266 ( \22519 , \22517 , \22518 );
not \U$22267 ( \22520 , \22519 );
not \U$22268 ( \22521 , \17005 );
and \U$22269 ( \22522 , \22520 , \22521 );
and \U$22270 ( \22523 , \22519 , \12957 );
nor \U$22271 ( \22524 , \22522 , \22523 );
xor \U$22272 ( \22525 , \22514 , \22524 );
and \U$22273 ( \22526 , \9909 , RIbe28ed0_43);
and \U$22274 ( \22527 , \13643 , RIbe27fd0_11);
nor \U$22275 ( \22528 , \22526 , \22527 );
and \U$22276 ( \22529 , \22528 , \16437 );
not \U$22277 ( \22530 , \22528 );
and \U$22278 ( \22531 , \22530 , \8077 );
nor \U$22279 ( \22532 , \22529 , \22531 );
and \U$22280 ( \22533 , \22525 , \22532 );
and \U$22281 ( \22534 , \22514 , \22524 );
or \U$22282 ( \22535 , \22533 , \22534 );
not \U$22283 ( \22536 , \22535 );
not \U$22284 ( \22537 , RIbe29560_57);
not \U$22285 ( \22538 , \13004 );
or \U$22286 ( \22539 , \22537 , \22538 );
nand \U$22287 ( \22540 , RIbe28228_16, RIbe2ae38_110);
nand \U$22288 ( \22541 , \22539 , \22540 );
not \U$22289 ( \22542 , RIbe2aeb0_111);
xor \U$22290 ( \22543 , \22541 , \22542 );
not \U$22291 ( \22544 , \22543 );
not \U$22292 ( \22545 , RIbe289a8_32);
not \U$22293 ( \22546 , \12887 );
or \U$22294 ( \22547 , \22545 , \22546 );
nand \U$22295 ( \22548 , \12890 , RIbe28930_31);
nand \U$22296 ( \22549 , \22547 , \22548 );
not \U$22297 ( \22550 , \22549 );
not \U$22298 ( \22551 , \12801 );
and \U$22299 ( \22552 , \22550 , \22551 );
and \U$22300 ( \22553 , \22549 , \12893 );
nor \U$22301 ( \22554 , \22552 , \22553 );
not \U$22302 ( \22555 , \22554 );
or \U$22303 ( \22556 , \22544 , \22555 );
not \U$22304 ( \22557 , \14558 );
not \U$22305 ( \22558 , RIbe29290_51);
not \U$22306 ( \22559 , \18608 );
or \U$22307 ( \22560 , \22558 , \22559 );
nand \U$22308 ( \22561 , \12835 , RIbe28a20_33);
nand \U$22309 ( \22562 , \22560 , \22561 );
not \U$22310 ( \22563 , \22562 );
or \U$22311 ( \22564 , \22557 , \22563 );
or \U$22312 ( \22565 , \22562 , \13706 );
nand \U$22313 ( \22566 , \22564 , \22565 );
nand \U$22314 ( \22567 , \22556 , \22566 );
not \U$22315 ( \22568 , \22554 );
not \U$22316 ( \22569 , \22543 );
nand \U$22317 ( \22570 , \22568 , \22569 );
nand \U$22318 ( \22571 , \22567 , \22570 );
nor \U$22319 ( \22572 , \22536 , \22571 );
not \U$22320 ( \22573 , RIbe28b10_35);
not \U$22321 ( \22574 , \13074 );
or \U$22322 ( \22575 , \22573 , \22574 );
nand \U$22323 ( \22576 , \12735 , RIbe28b88_36);
nand \U$22324 ( \22577 , \22575 , \22576 );
and \U$22325 ( \22578 , \22577 , \21013 );
not \U$22326 ( \22579 , \22577 );
and \U$22327 ( \22580 , \22579 , \14543 );
nor \U$22328 ( \22581 , \22578 , \22580 );
not \U$22329 ( \22582 , \22581 );
not \U$22330 ( \22583 , RIbe28408_20);
not \U$22331 ( \22584 , \12707 );
or \U$22332 ( \22585 , \22583 , \22584 );
nand \U$22333 ( \22586 , \12710 , RIbe28390_19);
nand \U$22334 ( \22587 , \22585 , \22586 );
xor \U$22335 ( \22588 , \22587 , \12723 );
nand \U$22336 ( \22589 , \22582 , \22588 );
not \U$22337 ( \22590 , \14000 );
not \U$22338 ( \22591 , RIbe287c8_28);
not \U$22339 ( \22592 , \13738 );
or \U$22340 ( \22593 , \22591 , \22592 );
not \U$22341 ( \22594 , \12752 );
nand \U$22342 ( \22595 , \22594 , RIbe28480_21);
nand \U$22343 ( \22596 , \22593 , \22595 );
not \U$22344 ( \22597 , \22596 );
or \U$22345 ( \22598 , \22590 , \22597 );
or \U$22346 ( \22599 , \22596 , \12770 );
nand \U$22347 ( \22600 , \22598 , \22599 );
and \U$22348 ( \22601 , \22589 , \22600 );
nor \U$22349 ( \22602 , \22582 , \22588 );
nor \U$22350 ( \22603 , \22601 , \22602 );
or \U$22351 ( \22604 , \22572 , \22603 );
nand \U$22352 ( \22605 , \22536 , \22571 );
nand \U$22353 ( \22606 , \22604 , \22605 );
and \U$22354 ( \22607 , \22504 , \22606 );
nor \U$22355 ( \22608 , \22422 , \22503 );
nor \U$22356 ( \22609 , \22607 , \22608 );
nand \U$22357 ( \22610 , \1147 , RIbe2ab68_104);
and \U$22358 ( \22611 , \22610 , \1154 );
not \U$22359 ( \22612 , \22610 );
and \U$22360 ( \22613 , \22612 , \1157 );
or \U$22361 ( \22614 , \22611 , \22613 );
not \U$22362 ( \22615 , \22614 );
not \U$22363 ( \22616 , \20630 );
not \U$22364 ( \22617 , \20648 );
or \U$22365 ( \22618 , \22616 , \22617 );
or \U$22366 ( \22619 , \20648 , \20630 );
nand \U$22367 ( \22620 , \22618 , \22619 );
nor \U$22368 ( \22621 , \22620 , \20637 );
not \U$22369 ( \22622 , \22621 );
nand \U$22370 ( \22623 , \22620 , \20637 );
nand \U$22371 ( \22624 , \22622 , \22623 );
not \U$22372 ( \22625 , \22624 );
or \U$22373 ( \22626 , \22615 , \22625 );
not \U$22374 ( \22627 , \22621 );
not \U$22375 ( \22628 , \22614 );
nand \U$22376 ( \22629 , \22627 , \22623 , \22628 );
xor \U$22377 ( \22630 , \20683 , \20661 );
xnor \U$22378 ( \22631 , \22630 , \20670 );
nand \U$22379 ( \22632 , \22629 , \22631 );
nand \U$22380 ( \22633 , \22626 , \22632 );
nand \U$22381 ( \22634 , \22309 , \22290 , \22312 );
nand \U$22382 ( \22635 , \22633 , \22634 );
nand \U$22383 ( \22636 , \22314 , \22609 , \22635 );
not \U$22384 ( \22637 , \22636 );
not \U$22385 ( \22638 , \20713 );
not \U$22386 ( \22639 , \20750 );
or \U$22387 ( \22640 , \22638 , \22639 );
or \U$22388 ( \22641 , \20750 , \20713 );
nand \U$22389 ( \22642 , \22640 , \22641 );
not \U$22390 ( \22643 , \22642 );
and \U$22391 ( \22644 , \20873 , \20832 );
not \U$22392 ( \22645 , \20873 );
not \U$22393 ( \22646 , \20832 );
and \U$22394 ( \22647 , \22645 , \22646 );
nor \U$22395 ( \22648 , \22644 , \22647 );
not \U$22396 ( \22649 , \22648 );
not \U$22397 ( \22650 , \20793 );
and \U$22398 ( \22651 , \22649 , \22650 );
and \U$22399 ( \22652 , \22648 , \20793 );
nor \U$22400 ( \22653 , \22651 , \22652 );
nand \U$22401 ( \22654 , \22643 , \22653 );
not \U$22402 ( \22655 , \22654 );
xor \U$22403 ( \22656 , \20910 , \20949 );
xor \U$22404 ( \22657 , \20978 , \22656 );
not \U$22405 ( \22658 , \22657 );
or \U$22406 ( \22659 , \22655 , \22658 );
not \U$22407 ( \22660 , \22653 );
nand \U$22408 ( \22661 , \22660 , \22642 );
nand \U$22409 ( \22662 , \22659 , \22661 );
not \U$22410 ( \22663 , \22662 );
or \U$22411 ( \22664 , \22637 , \22663 );
not \U$22412 ( \22665 , \22609 );
nand \U$22413 ( \22666 , \22314 , \22635 );
nand \U$22414 ( \22667 , \22665 , \22666 );
nand \U$22415 ( \22668 , \22664 , \22667 );
not \U$22416 ( \22669 , \22668 );
xor \U$22417 ( \22670 , \22107 , \22112 );
xnor \U$22418 ( \22671 , \22670 , \22106 );
not \U$22419 ( \22672 , \22671 );
nand \U$22420 ( \22673 , \22669 , \22672 );
not \U$22421 ( \22674 , \20437 );
not \U$22422 ( \22675 , \20510 );
or \U$22423 ( \22676 , \22674 , \22675 );
nand \U$22424 ( \22677 , \20509 , \20436 );
nand \U$22425 ( \22678 , \22676 , \22677 );
not \U$22426 ( \22679 , \22678 );
not \U$22427 ( \22680 , \20472 );
and \U$22428 ( \22681 , \22679 , \22680 );
and \U$22429 ( \22682 , \20472 , \22678 );
nor \U$22430 ( \22683 , \22681 , \22682 );
not \U$22431 ( \22684 , \22683 );
not \U$22432 ( \22685 , \22684 );
xor \U$22433 ( \22686 , \20575 , \20553 );
xnor \U$22434 ( \22687 , \22686 , \20609 );
not \U$22435 ( \22688 , \22687 );
not \U$22436 ( \22689 , \22688 );
or \U$22437 ( \22690 , \22685 , \22689 );
not \U$22438 ( \22691 , \22687 );
not \U$22439 ( \22692 , \22683 );
or \U$22440 ( \22693 , \22691 , \22692 );
xor \U$22441 ( \22694 , \20622 , \20651 );
xor \U$22442 ( \22695 , \22694 , \20687 );
nand \U$22443 ( \22696 , \22693 , \22695 );
nand \U$22444 ( \22697 , \22690 , \22696 );
not \U$22445 ( \22698 , \22697 );
or \U$22446 ( \22699 , \21365 , \21323 );
nand \U$22447 ( \22700 , \21365 , \21323 );
nand \U$22448 ( \22701 , \22699 , \22700 );
xor \U$22449 ( \22702 , \22701 , \21305 );
or \U$22450 ( \22703 , \22698 , \22702 );
not \U$22451 ( \22704 , \22698 );
not \U$22452 ( \22705 , \22702 );
or \U$22453 ( \22706 , \22704 , \22705 );
xor \U$22454 ( \22707 , \21037 , \21272 );
xor \U$22455 ( \22708 , \22707 , \21269 );
nand \U$22456 ( \22709 , \22706 , \22708 );
nand \U$22457 ( \22710 , \22703 , \22709 );
and \U$22458 ( \22711 , \22673 , \22710 );
and \U$22459 ( \22712 , \22668 , \22671 );
nor \U$22460 ( \22713 , \22711 , \22712 );
nand \U$22461 ( \22714 , \22267 , \22713 );
not \U$22462 ( \22715 , \22714 );
xor \U$22463 ( \22716 , \21451 , \21755 );
xnor \U$22464 ( \22717 , \22716 , \21752 );
not \U$22465 ( \22718 , \22717 );
xor \U$22466 ( \22719 , \20693 , \20985 );
xor \U$22467 ( \22720 , \22719 , \21274 );
not \U$22468 ( \22721 , \22720 );
xor \U$22469 ( \22722 , \22095 , \22090 );
xor \U$22470 ( \22723 , \22722 , \22086 );
nand \U$22471 ( \22724 , \22721 , \22723 );
not \U$22472 ( \22725 , \22724 );
or \U$22473 ( \22726 , \22718 , \22725 );
not \U$22474 ( \22727 , \22723 );
nand \U$22475 ( \22728 , \22727 , \22720 );
nand \U$22476 ( \22729 , \22726 , \22728 );
not \U$22477 ( \22730 , \22729 );
or \U$22478 ( \22731 , \22715 , \22730 );
not \U$22479 ( \22732 , \22713 );
nand \U$22480 ( \22733 , \22732 , \22266 );
nand \U$22481 ( \22734 , \22731 , \22733 );
not \U$22482 ( \22735 , \22734 );
nand \U$22483 ( \22736 , \22126 , \22735 );
not \U$22484 ( \22737 , \22736 );
not \U$22485 ( \22738 , \22098 );
nand \U$22486 ( \22739 , \22115 , \22738 );
and \U$22487 ( \22740 , \22080 , \22739 );
nor \U$22488 ( \22741 , \22115 , \22738 );
nor \U$22489 ( \22742 , \22740 , \22741 );
nand \U$22490 ( \22743 , \22245 , \22261 );
and \U$22491 ( \22744 , \22240 , \22743 );
nor \U$22492 ( \22745 , \22245 , \22261 );
nor \U$22493 ( \22746 , \22744 , \22745 );
xor \U$22494 ( \22747 , \22742 , \22746 );
not \U$22495 ( \22748 , \21794 );
nand \U$22496 ( \22749 , \21825 , \22748 );
and \U$22497 ( \22750 , \22058 , \22749 );
nor \U$22498 ( \22751 , \21825 , \22748 );
nor \U$22499 ( \22752 , \22750 , \22751 );
xor \U$22500 ( \22753 , \22747 , \22752 );
nand \U$22501 ( \22754 , \22249 , \22260 );
and \U$22502 ( \22755 , \22754 , \22255 );
nor \U$22503 ( \22756 , \22249 , \22260 );
nor \U$22504 ( \22757 , \22755 , \22756 );
not \U$22505 ( \22758 , \22757 );
not \U$22506 ( \22759 , \22165 );
not \U$22507 ( \22760 , \22159 );
or \U$22508 ( \22761 , \22759 , \22760 );
nand \U$22509 ( \22762 , \22761 , \22163 );
or \U$22510 ( \22763 , \22159 , \22165 );
nand \U$22511 ( \22764 , \22762 , \22763 );
not \U$22512 ( \22765 , \22764 );
not \U$22513 ( \22766 , \22133 );
not \U$22514 ( \22767 , \22149 );
or \U$22515 ( \22768 , \22766 , \22767 );
not \U$22516 ( \22769 , \22148 );
not \U$22517 ( \22770 , \22134 );
or \U$22518 ( \22771 , \22769 , \22770 );
nand \U$22519 ( \22772 , \22771 , \22140 );
nand \U$22520 ( \22773 , \22768 , \22772 );
not \U$22521 ( \22774 , \22773 );
not \U$22522 ( \22775 , \22774 );
or \U$22523 ( \22776 , \22765 , \22775 );
or \U$22524 ( \22777 , \22774 , \22764 );
nand \U$22525 ( \22778 , \22776 , \22777 );
not \U$22526 ( \22779 , \22778 );
or \U$22527 ( \22780 , \22758 , \22779 );
or \U$22528 ( \22781 , \22778 , \22757 );
nand \U$22529 ( \22782 , \22780 , \22781 );
not \U$22530 ( \22783 , \22782 );
not \U$22531 ( \22784 , \22175 );
nand \U$22532 ( \22785 , \22784 , \22205 );
not \U$22533 ( \22786 , \22785 );
not \U$22534 ( \22787 , \22238 );
or \U$22535 ( \22788 , \22786 , \22787 );
not \U$22536 ( \22789 , \22205 );
nand \U$22537 ( \22790 , \22789 , \22175 );
nand \U$22538 ( \22791 , \22788 , \22790 );
not \U$22539 ( \22792 , \22791 );
not \U$22540 ( \22793 , \21950 );
not \U$22541 ( \22794 , \21884 );
or \U$22542 ( \22795 , \22793 , \22794 );
or \U$22543 ( \22796 , \21950 , \21884 );
nand \U$22544 ( \22797 , \22796 , \21917 );
nand \U$22545 ( \22798 , \22795 , \22797 );
not \U$22546 ( \22799 , \22798 );
not \U$22547 ( \22800 , \22799 );
or \U$22548 ( \22801 , \22792 , \22800 );
not \U$22549 ( \22802 , \22791 );
nand \U$22550 ( \22803 , \22802 , \22798 );
nand \U$22551 ( \22804 , \22801 , \22803 );
not \U$22552 ( \22805 , \22804 );
not \U$22553 ( \22806 , \21991 );
not \U$22554 ( \22807 , \22806 );
nand \U$22555 ( \22808 , \22056 , \22807 );
and \U$22556 ( \22809 , \22808 , \22022 );
nor \U$22557 ( \22810 , \22056 , \22807 );
nor \U$22558 ( \22811 , \22809 , \22810 );
buf \U$22559 ( \22812 , \22811 );
not \U$22560 ( \22813 , \22812 );
and \U$22561 ( \22814 , \22805 , \22813 );
and \U$22562 ( \22815 , \22804 , \22812 );
nor \U$22563 ( \22816 , \22814 , \22815 );
not \U$22564 ( \22817 , \22816 );
and \U$22565 ( \22818 , \22783 , \22817 );
and \U$22566 ( \22819 , \22782 , \22816 );
nor \U$22567 ( \22820 , \22818 , \22819 );
nand \U$22568 ( \22821 , \21818 , \21797 );
not \U$22569 ( \22822 , \21686 );
not \U$22570 ( \22823 , \21714 );
or \U$22571 ( \22824 , \22822 , \22823 );
nand \U$22572 ( \22825 , \22824 , \21798 );
nor \U$22573 ( \22826 , \22821 , \22825 );
not \U$22574 ( \22827 , \22826 );
not \U$22575 ( \22828 , \21809 );
and \U$22576 ( \22829 , \22827 , \22828 );
and \U$22577 ( \22830 , \21799 , \21820 );
nor \U$22578 ( \22831 , \22829 , \22830 );
not \U$22579 ( \22832 , \21782 );
not \U$22580 ( \22833 , \21779 );
or \U$22581 ( \22834 , \22832 , \22833 );
nand \U$22582 ( \22835 , \22834 , \21793 );
not \U$22583 ( \22836 , \21779 );
nand \U$22584 ( \22837 , \22836 , \21770 );
and \U$22585 ( \22838 , \22835 , \22837 );
xor \U$22586 ( \22839 , \22831 , \22838 );
nand \U$22587 ( \22840 , \22057 , \21850 );
xor \U$22588 ( \22841 , \21951 , \21885 );
and \U$22589 ( \22842 , \22840 , \22841 );
nor \U$22590 ( \22843 , \22057 , \21850 );
nor \U$22591 ( \22844 , \22842 , \22843 );
xor \U$22592 ( \22845 , \22839 , \22844 );
xor \U$22593 ( \22846 , \22820 , \22845 );
nand \U$22594 ( \22847 , \22239 , \22166 );
and \U$22595 ( \22848 , \22847 , \22153 );
nor \U$22596 ( \22849 , \22239 , \22166 );
nor \U$22597 ( \22850 , \22848 , \22849 );
not \U$22598 ( \22851 , \21838 );
nand \U$22599 ( \22852 , \21844 , \1618 );
not \U$22600 ( \22853 , \22852 );
or \U$22601 ( \22854 , \22851 , \22853 );
nand \U$22602 ( \22855 , \21845 , \3959 );
nand \U$22603 ( \22856 , \22854 , \22855 );
and \U$22604 ( \22857 , \21916 , \21895 );
nor \U$22605 ( \22858 , \22857 , \21905 );
nor \U$22606 ( \22859 , \21916 , \21895 );
nor \U$22607 ( \22860 , \22858 , \22859 );
xor \U$22608 ( \22861 , \22856 , \22860 );
and \U$22609 ( \22862 , \21949 , \21938 );
nor \U$22610 ( \22863 , \22862 , \21928 );
nor \U$22611 ( \22864 , \21949 , \21938 );
nor \U$22612 ( \22865 , \22863 , \22864 );
xnor \U$22613 ( \22866 , \22861 , \22865 );
or \U$22614 ( \22867 , \21870 , \21857 );
nand \U$22615 ( \22868 , \22867 , \21879 );
nand \U$22616 ( \22869 , \21870 , \21857 );
nand \U$22617 ( \22870 , \22868 , \22869 );
xor \U$22618 ( \22871 , \22001 , \22011 );
and \U$22619 ( \22872 , \22871 , \22021 );
and \U$22620 ( \22873 , \22001 , \22011 );
or \U$22621 ( \22874 , \22872 , \22873 );
xor \U$22622 ( \22875 , \22870 , \22874 );
buf \U$22623 ( \22876 , \22032 );
or \U$22624 ( \22877 , \22876 , \22044 );
nand \U$22625 ( \22878 , \22877 , \22055 );
nand \U$22626 ( \22879 , \22876 , \22044 );
nand \U$22627 ( \22880 , \22878 , \22879 );
xor \U$22628 ( \22881 , \22875 , \22880 );
xnor \U$22629 ( \22882 , \22866 , \22881 );
nand \U$22630 ( \22883 , \22203 , \22193 );
not \U$22631 ( \22884 , \22883 );
not \U$22632 ( \22885 , \22184 );
or \U$22633 ( \22886 , \22884 , \22885 );
not \U$22634 ( \22887 , \22193 );
nand \U$22635 ( \22888 , \22887 , \22204 );
nand \U$22636 ( \22889 , \22886 , \22888 );
not \U$22637 ( \22890 , \22889 );
not \U$22638 ( \22891 , \21962 );
not \U$22639 ( \22892 , \21986 );
or \U$22640 ( \22893 , \22891 , \22892 );
nand \U$22641 ( \22894 , \22893 , \21973 );
nand \U$22642 ( \22895 , \21989 , \21961 );
nand \U$22643 ( \22896 , \22894 , \22895 );
not \U$22644 ( \22897 , \22896 );
not \U$22645 ( \22898 , \22897 );
or \U$22646 ( \22899 , \22890 , \22898 );
not \U$22647 ( \22900 , \22889 );
nand \U$22648 ( \22901 , \22900 , \22896 );
nand \U$22649 ( \22902 , \22899 , \22901 );
not \U$22650 ( \22903 , \22902 );
not \U$22651 ( \22904 , \22226 );
and \U$22652 ( \22905 , \22904 , \22237 );
nor \U$22653 ( \22906 , \22905 , \22216 );
nor \U$22654 ( \22907 , \22904 , \22237 );
nor \U$22655 ( \22908 , \22906 , \22907 );
not \U$22656 ( \22909 , \22908 );
and \U$22657 ( \22910 , \22903 , \22909 );
and \U$22658 ( \22911 , \22902 , \22908 );
nor \U$22659 ( \22912 , \22910 , \22911 );
and \U$22660 ( \22913 , \22882 , \22912 );
not \U$22661 ( \22914 , \22882 );
not \U$22662 ( \22915 , \22912 );
and \U$22663 ( \22916 , \22914 , \22915 );
nor \U$22664 ( \22917 , \22913 , \22916 );
xor \U$22665 ( \22918 , \22850 , \22917 );
not \U$22666 ( \22919 , RIbe289a8_32);
not \U$22667 ( \22920 , \16759 );
or \U$22668 ( \22921 , \22919 , \22920 );
nand \U$22669 ( \22922 , \12710 , RIbe28930_31);
nand \U$22670 ( \22923 , \22921 , \22922 );
xor \U$22671 ( \22924 , \22923 , \12723 );
not \U$22672 ( \22925 , RIbe29560_57);
not \U$22673 ( \22926 , \14534 );
or \U$22674 ( \22927 , \22925 , \22926 );
nand \U$22675 ( \22928 , \12735 , RIbe28228_16);
nand \U$22676 ( \22929 , \22927 , \22928 );
not \U$22677 ( \22930 , \22929 );
not \U$22678 ( \22931 , \14542 );
and \U$22679 ( \22932 , \22930 , \22931 );
and \U$22680 ( \22933 , \22929 , \14543 );
nor \U$22681 ( \22934 , \22932 , \22933 );
xor \U$22682 ( \22935 , \22924 , \22934 );
not \U$22683 ( \22936 , \12752 );
not \U$22684 ( \22937 , \5177 );
and \U$22685 ( \22938 , \22936 , \22937 );
and \U$22686 ( \22939 , \15615 , RIbe29290_51);
nor \U$22687 ( \22940 , \22938 , \22939 );
and \U$22688 ( \22941 , \22940 , \12927 );
not \U$22689 ( \22942 , \22940 );
and \U$22690 ( \22943 , \22942 , \12924 );
nor \U$22691 ( \22944 , \22941 , \22943 );
xor \U$22692 ( \22945 , \22935 , \22944 );
not \U$22693 ( \22946 , \22945 );
and \U$22694 ( \22947 , \20405 , RIbe287c8_28);
and \U$22695 ( \22948 , \10919 , RIbe28480_21);
nor \U$22696 ( \22949 , \22947 , \22948 );
and \U$22697 ( \22950 , \22949 , \8077 );
not \U$22698 ( \22951 , \22949 );
and \U$22699 ( \22952 , \22951 , \7970 );
nor \U$22700 ( \22953 , \22950 , \22952 );
not \U$22701 ( \22954 , RIbe28b10_35);
not \U$22702 ( \22955 , \12942 );
or \U$22703 ( \22956 , \22954 , \22955 );
nand \U$22704 ( \22957 , \12948 , RIbe28b88_36);
nand \U$22705 ( \22958 , \22956 , \22957 );
and \U$22706 ( \22959 , \22958 , \12195 );
not \U$22707 ( \22960 , \22958 );
and \U$22708 ( \22961 , \22960 , \12957 );
nor \U$22709 ( \22962 , \22959 , \22961 );
xor \U$22710 ( \22963 , \22953 , \22962 );
not \U$22711 ( \22964 , RIbe28408_20);
not \U$22712 ( \22965 , \13024 );
or \U$22713 ( \22966 , \22964 , \22965 );
nand \U$22714 ( \22967 , \12212 , RIbe28390_19);
nand \U$22715 ( \22968 , \22966 , \22967 );
and \U$22716 ( \22969 , \22968 , \9902 );
not \U$22717 ( \22970 , \22968 );
and \U$22718 ( \22971 , \22970 , \13030 );
nor \U$22719 ( \22972 , \22969 , \22971 );
xor \U$22720 ( \22973 , \22963 , \22972 );
not \U$22721 ( \22974 , \22973 );
or \U$22722 ( \22975 , \22946 , \22974 );
or \U$22723 ( \22976 , \22973 , \22945 );
nand \U$22724 ( \22977 , \22975 , \22976 );
not \U$22725 ( \22978 , RIbe29650_59);
not \U$22726 ( \22979 , \12811 );
or \U$22727 ( \22980 , \22978 , \22979 );
nand \U$22728 ( \22981 , RIbe29038_46, RIbe2ae38_110);
nand \U$22729 ( \22982 , \22980 , \22981 );
xnor \U$22730 ( \22983 , \22982 , RIbe2aeb0_111);
not \U$22731 ( \22984 , \22983 );
not \U$22732 ( \22985 , \22984 );
not \U$22733 ( \22986 , RIbe29830_63);
not \U$22734 ( \22987 , \12786 );
or \U$22735 ( \22988 , \22986 , \22987 );
nand \U$22736 ( \22989 , RIbe296c8_60, \12794 );
nand \U$22737 ( \22990 , \22988 , \22989 );
and \U$22738 ( \22991 , \22990 , \12801 );
not \U$22739 ( \22992 , \22990 );
and \U$22740 ( \22993 , \22992 , \16334 );
nor \U$22741 ( \22994 , \22991 , \22993 );
not \U$22742 ( \22995 , \22994 );
or \U$22743 ( \22996 , \22985 , \22995 );
not \U$22744 ( \22997 , \22994 );
nand \U$22745 ( \22998 , \22997 , \22983 );
nand \U$22746 ( \22999 , \22996 , \22998 );
not \U$22747 ( \23000 , RIbe281b0_15);
not \U$22748 ( \23001 , \13010 );
or \U$22749 ( \23002 , \23000 , \23001 );
nand \U$22750 ( \23003 , \21679 , RIbe280c0_13);
nand \U$22751 ( \23004 , \23002 , \23003 );
and \U$22752 ( \23005 , \23004 , \14555 );
not \U$22753 ( \23006 , \23004 );
and \U$22754 ( \23007 , \23006 , \14558 );
nor \U$22755 ( \23008 , \23005 , \23007 );
xor \U$22756 ( \23009 , \22999 , \23008 );
not \U$22757 ( \23010 , \23009 );
and \U$22758 ( \23011 , \22977 , \23010 );
not \U$22759 ( \23012 , \22977 );
and \U$22760 ( \23013 , \23012 , \23009 );
nor \U$22761 ( \23014 , \23011 , \23013 );
and \U$22762 ( \23015 , \6980 , RIbe27f58_10);
not \U$22763 ( \23016 , RIbe27e68_8);
nor \U$22764 ( \23017 , \23016 , \6984 );
nor \U$22765 ( \23018 , \23015 , \23017 );
xor \U$22766 ( \23019 , \23018 , \8004 );
not \U$22767 ( \23020 , \23019 );
not \U$22768 ( \23021 , RIbe28660_25);
not \U$22769 ( \23022 , \14633 );
or \U$22770 ( \23023 , \23021 , \23022 );
nand \U$22771 ( \23024 , \13339 , RIbe285e8_24);
nand \U$22772 ( \23025 , \23023 , \23024 );
and \U$22773 ( \23026 , \23025 , \6948 );
not \U$22774 ( \23027 , \23025 );
and \U$22775 ( \23028 , \23027 , \9896 );
nor \U$22776 ( \23029 , \23026 , \23028 );
not \U$22777 ( \23030 , \23029 );
or \U$22778 ( \23031 , \23020 , \23030 );
or \U$22779 ( \23032 , \23029 , \23019 );
nand \U$22780 ( \23033 , \23031 , \23032 );
not \U$22781 ( \23034 , RIbe28ed0_43);
not \U$22782 ( \23035 , \6958 );
or \U$22783 ( \23036 , \23034 , \23035 );
nand \U$22784 ( \23037 , \6962 , RIbe27fd0_11);
nand \U$22785 ( \23038 , \23036 , \23037 );
not \U$22786 ( \23039 , \23038 );
not \U$22787 ( \23040 , \6572 );
and \U$22788 ( \23041 , \23039 , \23040 );
and \U$22789 ( \23042 , \23038 , \6569 );
nor \U$22790 ( \23043 , \23041 , \23042 );
not \U$22791 ( \23044 , \23043 );
and \U$22792 ( \23045 , \23033 , \23044 );
not \U$22793 ( \23046 , \23033 );
and \U$22794 ( \23047 , \23046 , \23043 );
nor \U$22795 ( \23048 , \23045 , \23047 );
not \U$22796 ( \23049 , RIbe29dd0_75);
not \U$22797 ( \23050 , \6535 );
or \U$22798 ( \23051 , \23049 , \23050 );
nand \U$22799 ( \23052 , \6540 , RIbe29c68_72);
nand \U$22800 ( \23053 , \23051 , \23052 );
and \U$22801 ( \23054 , \23053 , \6552 );
not \U$22802 ( \23055 , \23053 );
and \U$22803 ( \23056 , \23055 , \6891 );
nor \U$22804 ( \23057 , \23054 , \23056 );
not \U$22805 ( \23058 , RIbe29fb0_79);
not \U$22806 ( \23059 , \6138 );
or \U$22807 ( \23060 , \23058 , \23059 );
nand \U$22808 ( \23061 , \9939 , RIbe29e48_76);
nand \U$22809 ( \23062 , \23060 , \23061 );
and \U$22810 ( \23063 , \23062 , \6623 );
not \U$22811 ( \23064 , \23062 );
and \U$22812 ( \23065 , \23064 , \10972 );
nor \U$22813 ( \23066 , \23063 , \23065 );
xor \U$22814 ( \23067 , \23057 , \23066 );
not \U$22815 ( \23068 , RIbe29bf0_71);
not \U$22816 ( \23069 , \6868 );
or \U$22817 ( \23070 , \23068 , \23069 );
nand \U$22818 ( \23071 , \13436 , RIbe28f48_44);
nand \U$22819 ( \23072 , \23070 , \23071 );
and \U$22820 ( \23073 , \23072 , \6601 );
not \U$22821 ( \23074 , \23072 );
and \U$22822 ( \23075 , \23074 , \7271 );
nor \U$22823 ( \23076 , \23073 , \23075 );
xor \U$22824 ( \23077 , \23067 , \23076 );
xor \U$22825 ( \23078 , \23048 , \23077 );
not \U$22826 ( \23079 , RIbe2a370_87);
not \U$22827 ( \23080 , \4829 );
or \U$22828 ( \23081 , \23079 , \23080 );
nand \U$22829 ( \23082 , \5052 , RIbe2a2f8_86);
nand \U$22830 ( \23083 , \23081 , \23082 );
and \U$22831 ( \23084 , \23083 , \4586 );
not \U$22832 ( \23085 , \23083 );
and \U$22833 ( \23086 , \23085 , \4946 );
nor \U$22834 ( \23087 , \23084 , \23086 );
not \U$22835 ( \23088 , \23087 );
not \U$22836 ( \23089 , \23088 );
not \U$22837 ( \23090 , RIbe2acd0_107);
not \U$22838 ( \23091 , \5455 );
or \U$22839 ( \23092 , \23090 , \23091 );
nand \U$22840 ( \23093 , \6634 , RIbe2a028_80);
nand \U$22841 ( \23094 , \23092 , \23093 );
not \U$22842 ( \23095 , \23094 );
not \U$22843 ( \23096 , \5754 );
and \U$22844 ( \23097 , \23095 , \23096 );
and \U$22845 ( \23098 , \23094 , \6641 );
nor \U$22846 ( \23099 , \23097 , \23098 );
not \U$22847 ( \23100 , \23099 );
not \U$22848 ( \23101 , \23100 );
or \U$22849 ( \23102 , \23089 , \23101 );
nand \U$22850 ( \23103 , \23099 , \23087 );
nand \U$22851 ( \23104 , \23102 , \23103 );
not \U$22852 ( \23105 , RIbe2b5b8_126);
not \U$22853 ( \23106 , \6413 );
or \U$22854 ( \23107 , \23105 , \23106 );
nand \U$22855 ( \23108 , \4808 , RIbe2a3e8_88);
nand \U$22856 ( \23109 , \23107 , \23108 );
not \U$22857 ( \23110 , \23109 );
not \U$22858 ( \23111 , \4323 );
and \U$22859 ( \23112 , \23110 , \23111 );
and \U$22860 ( \23113 , \23109 , \7865 );
nor \U$22861 ( \23114 , \23112 , \23113 );
not \U$22862 ( \23115 , \23114 );
and \U$22863 ( \23116 , \23104 , \23115 );
not \U$22864 ( \23117 , \23104 );
and \U$22865 ( \23118 , \23117 , \23114 );
nor \U$22866 ( \23119 , \23116 , \23118 );
xor \U$22867 ( \23120 , \23078 , \23119 );
or \U$22868 ( \23121 , \23014 , \23120 );
nand \U$22869 ( \23122 , \23014 , \23120 );
nand \U$22870 ( \23123 , \23121 , \23122 );
and \U$22871 ( \23124 , \2583 , RIbe2b090_115);
and \U$22872 ( \23125 , \2384 , RIbe2a280_85);
nor \U$22873 ( \23126 , \23124 , \23125 );
and \U$22874 ( \23127 , \23126 , \1274 );
not \U$22875 ( \23128 , \23126 );
and \U$22876 ( \23129 , \23128 , \1076 );
nor \U$22877 ( \23130 , \23127 , \23129 );
and \U$22878 ( \23131 , \2554 , RIbe2b270_119);
and \U$22879 ( \23132 , \5467 , RIbe2b108_116);
nor \U$22880 ( \23133 , \23131 , \23132 );
and \U$22881 ( \23134 , \23133 , \1131 );
not \U$22882 ( \23135 , \23133 );
and \U$22883 ( \23136 , \23135 , \6831 );
nor \U$22884 ( \23137 , \23134 , \23136 );
and \U$22885 ( \23138 , \23130 , \23137 );
not \U$22886 ( \23139 , \23130 );
not \U$22887 ( \23140 , \23137 );
and \U$22888 ( \23141 , \23139 , \23140 );
nor \U$22889 ( \23142 , \23138 , \23141 );
not \U$22890 ( \23143 , RIbe2b1f8_118);
not \U$22891 ( \23144 , \1298 );
or \U$22892 ( \23145 , \23143 , \23144 );
nand \U$22893 ( \23146 , \1454 , RIbe2b180_117);
nand \U$22894 ( \23147 , \23145 , \23146 );
not \U$22895 ( \23148 , \23147 );
not \U$22896 ( \23149 , \1458 );
and \U$22897 ( \23150 , \23148 , \23149 );
and \U$22898 ( \23151 , \23147 , \1458 );
nor \U$22899 ( \23152 , \23150 , \23151 );
not \U$22900 ( \23153 , \23152 );
xor \U$22901 ( \23154 , \23142 , \23153 );
not \U$22902 ( \23155 , RIbe2a5c8_92);
not \U$22903 ( \23156 , \3451 );
or \U$22904 ( \23157 , \23155 , \23156 );
nand \U$22905 ( \23158 , \6800 , RIbe2a550_91);
nand \U$22906 ( \23159 , \23157 , \23158 );
and \U$22907 ( \23160 , \23159 , \2887 );
not \U$22908 ( \23161 , \23159 );
and \U$22909 ( \23162 , \23161 , \4346 );
nor \U$22910 ( \23163 , \23160 , \23162 );
not \U$22911 ( \23164 , RIbe2a988_100);
not \U$22912 ( \23165 , \20764 );
or \U$22913 ( \23166 , \23164 , \23165 );
nand \U$22914 ( \23167 , \8368 , RIbe2a910_99);
nand \U$22915 ( \23168 , \23166 , \23167 );
and \U$22916 ( \23169 , \23168 , \3471 );
not \U$22917 ( \23170 , \23168 );
and \U$22918 ( \23171 , \23170 , \3448 );
nor \U$22919 ( \23172 , \23169 , \23171 );
xor \U$22920 ( \23173 , \23163 , \23172 );
not \U$22921 ( \23174 , RIbe2a208_84);
not \U$22922 ( \23175 , \7827 );
or \U$22923 ( \23176 , \23174 , \23175 );
nand \U$22924 ( \23177 , \4284 , RIbe2a190_83);
nand \U$22925 ( \23178 , \23176 , \23177 );
not \U$22926 ( \23179 , \23178 );
not \U$22927 ( \23180 , \3275 );
and \U$22928 ( \23181 , \23179 , \23180 );
and \U$22929 ( \23182 , \23178 , \2379 );
nor \U$22930 ( \23183 , \23181 , \23182 );
xor \U$22931 ( \23184 , \23173 , \23183 );
xor \U$22932 ( \23185 , \23154 , \23184 );
not \U$22933 ( \23186 , RIbe2ab68_104);
not \U$22934 ( \23187 , \7363 );
or \U$22935 ( \23188 , \23186 , \23187 );
nand \U$22936 ( \23189 , \740 , RIbe2aaf0_103);
nand \U$22937 ( \23190 , \23188 , \23189 );
and \U$22938 ( \23191 , \23190 , \3959 );
not \U$22939 ( \23192 , \23190 );
and \U$22940 ( \23193 , \23192 , \564 );
nor \U$22941 ( \23194 , \23191 , \23193 );
not \U$22942 ( \23195 , RIbe2afa0_113);
not \U$22943 ( \23196 , \2597 );
or \U$22944 ( \23197 , \23195 , \23196 );
nand \U$22945 ( \23198 , \1147 , RIbe2af28_112);
nand \U$22946 ( \23199 , \23197 , \23198 );
not \U$22947 ( \23200 , \23199 );
not \U$22948 ( \23201 , \4742 );
and \U$22949 ( \23202 , \23200 , \23201 );
and \U$22950 ( \23203 , \23199 , \1153 );
nor \U$22951 ( \23204 , \23202 , \23203 );
xor \U$22952 ( \23205 , \23194 , \23204 );
and \U$22953 ( \23206 , \5973 , RIbe2b630_127);
and \U$22954 ( \23207 , \1203 , RIbe2b018_114);
nor \U$22955 ( \23208 , \23206 , \23207 );
and \U$22956 ( \23209 , \23208 , \1011 );
not \U$22957 ( \23210 , \23208 );
and \U$22958 ( \23211 , \23210 , \1813 );
nor \U$22959 ( \23212 , \23209 , \23211 );
xor \U$22960 ( \23213 , \23205 , \23212 );
xor \U$22961 ( \23214 , \23185 , \23213 );
not \U$22962 ( \23215 , \23214 );
and \U$22963 ( \23216 , \23123 , \23215 );
not \U$22964 ( \23217 , \23123 );
and \U$22965 ( \23218 , \23217 , \23214 );
nor \U$22966 ( \23219 , \23216 , \23218 );
xor \U$22967 ( \23220 , \22918 , \23219 );
xor \U$22968 ( \23221 , \22846 , \23220 );
xor \U$22969 ( \23222 , \22753 , \23221 );
nand \U$22970 ( \23223 , \22066 , \21761 );
and \U$22971 ( \23224 , \23223 , \21757 );
nor \U$22972 ( \23225 , \22066 , \21761 );
nor \U$22973 ( \23226 , \23224 , \23225 );
xor \U$22974 ( \23227 , \23222 , \23226 );
not \U$22975 ( \23228 , \23227 );
not \U$22976 ( \23229 , \23228 );
or \U$22977 ( \23230 , \22737 , \23229 );
nand \U$22978 ( \23231 , \22070 , \22734 , \22124 );
nand \U$22979 ( \23232 , \23230 , \23231 );
not \U$22980 ( \23233 , \22816 );
nand \U$22981 ( \23234 , \23233 , \22782 );
xor \U$22982 ( \23235 , \22831 , \22838 );
and \U$22983 ( \23236 , \23235 , \22844 );
and \U$22984 ( \23237 , \22831 , \22838 );
or \U$22985 ( \23238 , \23236 , \23237 );
xor \U$22986 ( \23239 , \23234 , \23238 );
xor \U$22987 ( \23240 , \22850 , \22917 );
and \U$22988 ( \23241 , \23240 , \23219 );
and \U$22989 ( \23242 , \22850 , \22917 );
or \U$22990 ( \23243 , \23241 , \23242 );
xor \U$22991 ( \23244 , \23239 , \23243 );
xor \U$22992 ( \23245 , \22753 , \23221 );
and \U$22993 ( \23246 , \23245 , \23226 );
and \U$22994 ( \23247 , \22753 , \23221 );
or \U$22995 ( \23248 , \23246 , \23247 );
xor \U$22996 ( \23249 , \23244 , \23248 );
xor \U$22997 ( \23250 , \22742 , \22746 );
and \U$22998 ( \23251 , \23250 , \22752 );
and \U$22999 ( \23252 , \22742 , \22746 );
or \U$23000 ( \23253 , \23251 , \23252 );
xor \U$23001 ( \23254 , \22820 , \22845 );
and \U$23002 ( \23255 , \23254 , \23220 );
and \U$23003 ( \23256 , \22820 , \22845 );
or \U$23004 ( \23257 , \23255 , \23256 );
xor \U$23005 ( \23258 , \23253 , \23257 );
not \U$23006 ( \23259 , \22799 );
not \U$23007 ( \23260 , \22811 );
or \U$23008 ( \23261 , \23259 , \23260 );
nand \U$23009 ( \23262 , \23261 , \22791 );
not \U$23010 ( \23263 , \22811 );
nand \U$23011 ( \23264 , \23263 , \22798 );
nand \U$23012 ( \23265 , \23262 , \23264 );
not \U$23013 ( \23266 , \23265 );
not \U$23014 ( \23267 , \22774 );
not \U$23015 ( \23268 , \22757 );
or \U$23016 ( \23269 , \23267 , \23268 );
nand \U$23017 ( \23270 , \23269 , \22764 );
not \U$23018 ( \23271 , \22757 );
nand \U$23019 ( \23272 , \23271 , \22773 );
nand \U$23020 ( \23273 , \23270 , \23272 );
not \U$23021 ( \23274 , \23273 );
not \U$23022 ( \23275 , \23274 );
and \U$23023 ( \23276 , \23266 , \23275 );
and \U$23024 ( \23277 , \23265 , \23274 );
nor \U$23025 ( \23278 , \23276 , \23277 );
not \U$23026 ( \23279 , \23014 );
not \U$23027 ( \23280 , \23279 );
not \U$23028 ( \23281 , \23120 );
or \U$23029 ( \23282 , \23280 , \23281 );
or \U$23030 ( \23283 , \23279 , \23120 );
nand \U$23031 ( \23284 , \23283 , \23214 );
nand \U$23032 ( \23285 , \23282 , \23284 );
xor \U$23033 ( \23286 , \23278 , \23285 );
not \U$23034 ( \23287 , \23286 );
not \U$23035 ( \23288 , \22866 );
not \U$23036 ( \23289 , \22912 );
or \U$23037 ( \23290 , \23288 , \23289 );
nand \U$23038 ( \23291 , \23290 , \22881 );
not \U$23039 ( \23292 , \22866 );
nand \U$23040 ( \23293 , \23292 , \22915 );
nand \U$23041 ( \23294 , \23291 , \23293 );
not \U$23042 ( \23295 , \22983 );
not \U$23043 ( \23296 , \22994 );
or \U$23044 ( \23297 , \23295 , \23296 );
nand \U$23045 ( \23298 , \23297 , \23008 );
nand \U$23046 ( \23299 , \22984 , \22997 );
nand \U$23047 ( \23300 , \23298 , \23299 );
xor \U$23048 ( \23301 , \22924 , \22934 );
and \U$23049 ( \23302 , \23301 , \22944 );
and \U$23050 ( \23303 , \22924 , \22934 );
or \U$23051 ( \23304 , \23302 , \23303 );
not \U$23052 ( \23305 , \23304 );
xor \U$23053 ( \23306 , \23300 , \23305 );
xor \U$23054 ( \23307 , \22953 , \22962 );
and \U$23055 ( \23308 , \23307 , \22972 );
and \U$23056 ( \23309 , \22953 , \22962 );
or \U$23057 ( \23310 , \23308 , \23309 );
xor \U$23058 ( \23311 , \23306 , \23310 );
not \U$23059 ( \23312 , \23029 );
not \U$23060 ( \23313 , \23043 );
or \U$23061 ( \23314 , \23312 , \23313 );
nand \U$23062 ( \23315 , \23314 , \23019 );
not \U$23063 ( \23316 , \23029 );
nand \U$23064 ( \23317 , \23316 , \23044 );
nand \U$23065 ( \23318 , \23315 , \23317 );
not \U$23066 ( \23319 , \23115 );
not \U$23067 ( \23320 , \23087 );
or \U$23068 ( \23321 , \23319 , \23320 );
not \U$23069 ( \23322 , \23088 );
not \U$23070 ( \23323 , \23114 );
or \U$23071 ( \23324 , \23322 , \23323 );
nand \U$23072 ( \23325 , \23324 , \23100 );
nand \U$23073 ( \23326 , \23321 , \23325 );
xor \U$23074 ( \23327 , \23318 , \23326 );
xor \U$23075 ( \23328 , \23057 , \23066 );
and \U$23076 ( \23329 , \23328 , \23076 );
and \U$23077 ( \23330 , \23057 , \23066 );
or \U$23078 ( \23331 , \23329 , \23330 );
xor \U$23079 ( \23332 , \23327 , \23331 );
xor \U$23080 ( \23333 , \23311 , \23332 );
xor \U$23081 ( \23334 , \23294 , \23333 );
not \U$23082 ( \23335 , \1813 );
not \U$23083 ( \23336 , RIbe2b018_114);
not \U$23084 ( \23337 , \998 );
nand \U$23085 ( \23338 , \23337 , \1000 );
not \U$23086 ( \23339 , \23338 );
not \U$23087 ( \23340 , \23339 );
or \U$23088 ( \23341 , \23336 , \23340 );
nand \U$23089 ( \23342 , RIbe2afa0_113, \1202 );
nand \U$23090 ( \23343 , \23341 , \23342 );
not \U$23091 ( \23344 , \23343 );
and \U$23092 ( \23345 , \23335 , \23344 );
and \U$23093 ( \23346 , \23343 , \1813 );
nor \U$23094 ( \23347 , \23345 , \23346 );
not \U$23095 ( \23348 , RIbe2af28_112);
not \U$23096 ( \23349 , \21344 );
or \U$23097 ( \23350 , \23348 , \23349 );
nand \U$23098 ( \23351 , RIbe2b1f8_118, \1146 );
nand \U$23099 ( \23352 , \23350 , \23351 );
and \U$23100 ( \23353 , \23352 , \1153 );
not \U$23101 ( \23354 , \23352 );
and \U$23102 ( \23355 , \23354 , \7899 );
nor \U$23103 ( \23356 , \23353 , \23355 );
xor \U$23104 ( \23357 , \23347 , \23356 );
not \U$23105 ( \23358 , \1082 );
not \U$23106 ( \23359 , RIbe2b180_117);
not \U$23107 ( \23360 , \8868 );
or \U$23108 ( \23361 , \23359 , \23360 );
nand \U$23109 ( \23362 , \4730 , RIbe2b270_119);
nand \U$23110 ( \23363 , \23361 , \23362 );
not \U$23111 ( \23364 , \23363 );
or \U$23112 ( \23365 , \23358 , \23364 );
or \U$23113 ( \23366 , \23363 , \1458 );
nand \U$23114 ( \23367 , \23365 , \23366 );
xor \U$23115 ( \23368 , \23357 , \23367 );
nand \U$23116 ( \23369 , \553 , RIbe2ab68_104);
and \U$23117 ( \23370 , \23369 , \424 );
not \U$23118 ( \23371 , \23369 );
and \U$23119 ( \23372 , \23371 , \1330 );
or \U$23120 ( \23373 , \23370 , \23372 );
not \U$23121 ( \23374 , \23373 );
not \U$23122 ( \23375 , RIbe2aaf0_103);
not \U$23123 ( \23376 , \2531 );
or \U$23124 ( \23377 , \23375 , \23376 );
nand \U$23125 ( \23378 , \1179 , RIbe2b630_127);
nand \U$23126 ( \23379 , \23377 , \23378 );
and \U$23127 ( \23380 , \23379 , \3959 );
not \U$23128 ( \23381 , \23379 );
and \U$23129 ( \23382 , \23381 , \1618 );
nor \U$23130 ( \23383 , \23380 , \23382 );
not \U$23131 ( \23384 , \23383 );
or \U$23132 ( \23385 , \23374 , \23384 );
or \U$23133 ( \23386 , \23383 , \23373 );
nand \U$23134 ( \23387 , \23385 , \23386 );
xor \U$23135 ( \23388 , \23368 , \23387 );
not \U$23136 ( \23389 , \23388 );
not \U$23137 ( \23390 , \23389 );
not \U$23138 ( \23391 , \23130 );
nand \U$23139 ( \23392 , \23152 , \23137 );
nand \U$23140 ( \23393 , \23391 , \23392 );
nand \U$23141 ( \23394 , \23140 , \23153 );
nand \U$23142 ( \23395 , \23393 , \23394 );
nand \U$23143 ( \23396 , \23163 , \23183 );
and \U$23144 ( \23397 , \23396 , \23172 );
nor \U$23145 ( \23398 , \23163 , \23183 );
nor \U$23146 ( \23399 , \23397 , \23398 );
xor \U$23147 ( \23400 , \23395 , \23399 );
nand \U$23148 ( \23401 , \23204 , \23212 );
and \U$23149 ( \23402 , \23401 , \23194 );
nor \U$23150 ( \23403 , \23204 , \23212 );
nor \U$23151 ( \23404 , \23402 , \23403 );
xnor \U$23152 ( \23405 , \23400 , \23404 );
not \U$23153 ( \23406 , \23405 );
not \U$23154 ( \23407 , \23406 );
or \U$23155 ( \23408 , \23390 , \23407 );
nand \U$23156 ( \23409 , \23405 , \23388 );
nand \U$23157 ( \23410 , \23408 , \23409 );
not \U$23158 ( \23411 , RIbe2a910_99);
not \U$23159 ( \23412 , \20764 );
or \U$23160 ( \23413 , \23411 , \23412 );
nand \U$23161 ( \23414 , \6787 , RIbe2b5b8_126);
nand \U$23162 ( \23415 , \23413 , \23414 );
and \U$23163 ( \23416 , \23415 , \3471 );
not \U$23164 ( \23417 , \23415 );
and \U$23165 ( \23418 , \23417 , \3698 );
nor \U$23166 ( \23419 , \23416 , \23418 );
not \U$23167 ( \23420 , \23419 );
not \U$23168 ( \23421 , RIbe2a3e8_88);
not \U$23169 ( \23422 , \21040 );
or \U$23170 ( \23423 , \23421 , \23422 );
nand \U$23171 ( \23424 , \7858 , RIbe2a370_87);
nand \U$23172 ( \23425 , \23423 , \23424 );
and \U$23173 ( \23426 , \23425 , \4323 );
not \U$23174 ( \23427 , \23425 );
and \U$23175 ( \23428 , \23427 , \4326 );
nor \U$23176 ( \23429 , \23426 , \23428 );
not \U$23177 ( \23430 , \23429 );
or \U$23178 ( \23431 , \23420 , \23430 );
or \U$23179 ( \23432 , \23419 , \23429 );
nand \U$23180 ( \23433 , \23431 , \23432 );
not \U$23181 ( \23434 , RIbe2a550_91);
not \U$23182 ( \23435 , \6797 );
or \U$23183 ( \23436 , \23434 , \23435 );
nand \U$23184 ( \23437 , \6800 , RIbe2a988_100);
nand \U$23185 ( \23438 , \23436 , \23437 );
and \U$23186 ( \23439 , \23438 , \2887 );
not \U$23187 ( \23440 , \23438 );
and \U$23188 ( \23441 , \23440 , \3290 );
nor \U$23189 ( \23442 , \23439 , \23441 );
not \U$23190 ( \23443 , \23442 );
and \U$23191 ( \23444 , \23433 , \23443 );
not \U$23192 ( \23445 , \23433 );
and \U$23193 ( \23446 , \23445 , \23442 );
nor \U$23194 ( \23447 , \23444 , \23446 );
not \U$23195 ( \23448 , \23447 );
not \U$23196 ( \23449 , RIbe2a028_80);
not \U$23197 ( \23450 , \15313 );
or \U$23198 ( \23451 , \23449 , \23450 );
nand \U$23199 ( \23452 , \20439 , RIbe29fb0_79);
nand \U$23200 ( \23453 , \23451 , \23452 );
and \U$23201 ( \23454 , \23453 , \8253 );
not \U$23202 ( \23455 , \23453 );
and \U$23203 ( \23456 , \23455 , \5046 );
nor \U$23204 ( \23457 , \23454 , \23456 );
not \U$23205 ( \23458 , RIbe29e48_76);
not \U$23206 ( \23459 , \6856 );
or \U$23207 ( \23460 , \23458 , \23459 );
nand \U$23208 ( \23461 , \21084 , RIbe29dd0_75);
nand \U$23209 ( \23462 , \23460 , \23461 );
and \U$23210 ( \23463 , \23462 , \21093 );
not \U$23211 ( \23464 , \23462 );
and \U$23212 ( \23465 , \23464 , \21090 );
or \U$23213 ( \23466 , \23463 , \23465 );
xor \U$23214 ( \23467 , \23457 , \23466 );
not \U$23215 ( \23468 , RIbe2a2f8_86);
not \U$23216 ( \23469 , \21097 );
or \U$23217 ( \23470 , \23468 , \23469 );
nand \U$23218 ( \23471 , \5052 , RIbe2acd0_107);
nand \U$23219 ( \23472 , \23470 , \23471 );
and \U$23220 ( \23473 , \23472 , \4592 );
not \U$23221 ( \23474 , \23472 );
and \U$23222 ( \23475 , \23474 , \4586 );
nor \U$23223 ( \23476 , \23473 , \23475 );
not \U$23224 ( \23477 , \23476 );
xor \U$23225 ( \23478 , \23467 , \23477 );
not \U$23226 ( \23479 , \23478 );
or \U$23227 ( \23480 , \23448 , \23479 );
or \U$23228 ( \23481 , \23478 , \23447 );
nand \U$23229 ( \23482 , \23480 , \23481 );
not \U$23230 ( \23483 , RIbe2a190_83);
not \U$23231 ( \23484 , \10010 );
or \U$23232 ( \23485 , \23483 , \23484 );
nand \U$23233 ( \23486 , \2901 , RIbe2a5c8_92);
nand \U$23234 ( \23487 , \23485 , \23486 );
not \U$23235 ( \23488 , \23487 );
not \U$23236 ( \23489 , \2379 );
and \U$23237 ( \23490 , \23488 , \23489 );
and \U$23238 ( \23491 , \23487 , \2576 );
nor \U$23239 ( \23492 , \23490 , \23491 );
not \U$23240 ( \23493 , \23492 );
not \U$23241 ( \23494 , \3516 );
not \U$23242 ( \23495 , RIbe2a280_85);
not \U$23243 ( \23496 , \2583 );
or \U$23244 ( \23497 , \23495 , \23496 );
nand \U$23245 ( \23498 , \2384 , RIbe2a208_84);
nand \U$23246 ( \23499 , \23497 , \23498 );
not \U$23247 ( \23500 , \23499 );
or \U$23248 ( \23501 , \23494 , \23500 );
or \U$23249 ( \23502 , \23499 , \7038 );
nand \U$23250 ( \23503 , \23501 , \23502 );
not \U$23251 ( \23504 , \23503 );
or \U$23252 ( \23505 , \23493 , \23504 );
or \U$23253 ( \23506 , \23503 , \23492 );
nand \U$23254 ( \23507 , \23505 , \23506 );
not \U$23255 ( \23508 , RIbe2b108_116);
not \U$23256 ( \23509 , \1284 );
not \U$23257 ( \23510 , \23509 );
or \U$23258 ( \23511 , \23508 , \23510 );
nand \U$23259 ( \23512 , \20849 , RIbe2b090_115);
nand \U$23260 ( \23513 , \23511 , \23512 );
not \U$23261 ( \23514 , \23513 );
not \U$23262 ( \23515 , \2563 );
and \U$23263 ( \23516 , \23514 , \23515 );
and \U$23264 ( \23517 , \23513 , \1448 );
nor \U$23265 ( \23518 , \23516 , \23517 );
buf \U$23266 ( \23519 , \23518 );
xnor \U$23267 ( \23520 , \23507 , \23519 );
not \U$23268 ( \23521 , \23520 );
and \U$23269 ( \23522 , \23482 , \23521 );
not \U$23270 ( \23523 , \23482 );
and \U$23271 ( \23524 , \23523 , \23520 );
nor \U$23272 ( \23525 , \23522 , \23524 );
not \U$23273 ( \23526 , \23525 );
and \U$23274 ( \23527 , \23410 , \23526 );
not \U$23275 ( \23528 , \23410 );
and \U$23276 ( \23529 , \23528 , \23525 );
nor \U$23277 ( \23530 , \23527 , \23529 );
xor \U$23278 ( \23531 , \23334 , \23530 );
not \U$23279 ( \23532 , \23531 );
or \U$23280 ( \23533 , \23287 , \23532 );
not \U$23281 ( \23534 , \23531 );
not \U$23282 ( \23535 , \23286 );
nand \U$23283 ( \23536 , \23534 , \23535 );
nand \U$23284 ( \23537 , \23533 , \23536 );
not \U$23285 ( \23538 , RIbe28f48_44);
not \U$23286 ( \23539 , \6868 );
or \U$23287 ( \23540 , \23538 , \23539 );
nand \U$23288 ( \23541 , \7278 , RIbe28ed0_43);
nand \U$23289 ( \23542 , \23540 , \23541 );
and \U$23290 ( \23543 , \23542 , \6582 );
not \U$23291 ( \23544 , \23542 );
and \U$23292 ( \23545 , \23544 , \6583 );
nor \U$23293 ( \23546 , \23543 , \23545 );
not \U$23294 ( \23547 , RIbe27fd0_11);
not \U$23295 ( \23548 , \21608 );
or \U$23296 ( \23549 , \23547 , \23548 );
nand \U$23297 ( \23550 , \7958 , RIbe27f58_10);
nand \U$23298 ( \23551 , \23549 , \23550 );
and \U$23299 ( \23552 , \23551 , \7293 );
not \U$23300 ( \23553 , \23551 );
and \U$23301 ( \23554 , \23553 , \6572 );
nor \U$23302 ( \23555 , \23552 , \23554 );
xor \U$23303 ( \23556 , \23546 , \23555 );
not \U$23304 ( \23557 , RIbe29c68_72);
not \U$23305 ( \23558 , \6536 );
or \U$23306 ( \23559 , \23557 , \23558 );
nand \U$23307 ( \23560 , \6540 , RIbe29bf0_71);
nand \U$23308 ( \23561 , \23559 , \23560 );
and \U$23309 ( \23562 , \23561 , \15730 );
not \U$23310 ( \23563 , \23561 );
and \U$23311 ( \23564 , \23563 , \13412 );
nor \U$23312 ( \23565 , \23562 , \23564 );
not \U$23313 ( \23566 , \23565 );
and \U$23314 ( \23567 , \23556 , \23566 );
not \U$23315 ( \23568 , \23556 );
and \U$23316 ( \23569 , \23568 , \23565 );
nor \U$23317 ( \23570 , \23567 , \23569 );
not \U$23318 ( \23571 , \23570 );
not \U$23319 ( \23572 , \13085 );
not \U$23320 ( \23573 , \3421 );
and \U$23321 ( \23574 , \23572 , \23573 );
and \U$23322 ( \23575 , \12764 , RIbe28a20_33);
nor \U$23323 ( \23576 , \23574 , \23575 );
and \U$23324 ( \23577 , \23576 , \12774 );
not \U$23325 ( \23578 , \23576 );
and \U$23326 ( \23579 , \23578 , \14000 );
nor \U$23327 ( \23580 , \23577 , \23579 );
not \U$23328 ( \23581 , \23580 );
not \U$23329 ( \23582 , RIbe28b88_36);
not \U$23330 ( \23583 , \12942 );
or \U$23331 ( \23584 , \23582 , \23583 );
nand \U$23332 ( \23585 , \12947 , RIbe29290_51);
nand \U$23333 ( \23586 , \23584 , \23585 );
and \U$23334 ( \23587 , \23586 , \12195 );
not \U$23335 ( \23588 , \23586 );
and \U$23336 ( \23589 , \23588 , \12960 );
nor \U$23337 ( \23590 , \23587 , \23589 );
not \U$23338 ( \23591 , \23590 );
or \U$23339 ( \23592 , \23581 , \23591 );
or \U$23340 ( \23593 , \23590 , \23580 );
nand \U$23341 ( \23594 , \23592 , \23593 );
not \U$23342 ( \23595 , RIbe28390_19);
not \U$23343 ( \23596 , \10936 );
or \U$23344 ( \23597 , \23595 , \23596 );
nand \U$23345 ( \23598 , \12971 , RIbe28b10_35);
nand \U$23346 ( \23599 , \23597 , \23598 );
and \U$23347 ( \23600 , \23599 , \10940 );
not \U$23348 ( \23601 , \23599 );
and \U$23349 ( \23602 , \23601 , \9901 );
nor \U$23350 ( \23603 , \23600 , \23602 );
buf \U$23351 ( \23604 , \23603 );
and \U$23352 ( \23605 , \23594 , \23604 );
not \U$23353 ( \23606 , \23594 );
not \U$23354 ( \23607 , \23604 );
and \U$23355 ( \23608 , \23606 , \23607 );
nor \U$23356 ( \23609 , \23605 , \23608 );
not \U$23357 ( \23610 , \23609 );
not \U$23358 ( \23611 , \23610 );
or \U$23359 ( \23612 , \23571 , \23611 );
not \U$23360 ( \23613 , \23570 );
nand \U$23361 ( \23614 , \23609 , \23613 );
nand \U$23362 ( \23615 , \23612 , \23614 );
not \U$23363 ( \23616 , RIbe28480_21);
not \U$23364 ( \23617 , \14622 );
or \U$23365 ( \23618 , \23616 , \23617 );
nand \U$23366 ( \23619 , \13038 , RIbe28408_20);
nand \U$23367 ( \23620 , \23618 , \23619 );
xor \U$23368 ( \23621 , \23620 , \8077 );
not \U$23369 ( \23622 , \23621 );
not \U$23370 ( \23623 , RIbe285e8_24);
not \U$23371 ( \23624 , \14633 );
or \U$23372 ( \23625 , \23623 , \23624 );
nand \U$23373 ( \23626 , \9891 , RIbe287c8_28);
nand \U$23374 ( \23627 , \23625 , \23626 );
and \U$23375 ( \23628 , \23627 , \14299 );
not \U$23376 ( \23629 , \23627 );
and \U$23377 ( \23630 , \23629 , \6949 );
nor \U$23378 ( \23631 , \23628 , \23630 );
not \U$23379 ( \23632 , \23631 );
or \U$23380 ( \23633 , \23622 , \23632 );
or \U$23381 ( \23634 , \23621 , \23631 );
nand \U$23382 ( \23635 , \23633 , \23634 );
not \U$23383 ( \23636 , RIbe27e68_8);
not \U$23384 ( \23637 , \7298 );
or \U$23385 ( \23638 , \23636 , \23637 );
nand \U$23386 ( \23639 , \9875 , RIbe28660_25);
nand \U$23387 ( \23640 , \23638 , \23639 );
and \U$23388 ( \23641 , \23640 , \7660 );
not \U$23389 ( \23642 , \23640 );
and \U$23390 ( \23643 , \23642 , \6992 );
nor \U$23391 ( \23644 , \23641 , \23643 );
not \U$23392 ( \23645 , \23644 );
and \U$23393 ( \23646 , \23635 , \23645 );
not \U$23394 ( \23647 , \23635 );
and \U$23395 ( \23648 , \23647 , \23644 );
nor \U$23396 ( \23649 , \23646 , \23648 );
xnor \U$23397 ( \23650 , \23615 , \23649 );
not \U$23398 ( \23651 , \23650 );
not \U$23399 ( \23652 , RIbe29038_46);
not \U$23400 ( \23653 , \13003 );
or \U$23401 ( \23654 , \23652 , \23653 );
nand \U$23402 ( \23655 , RIbe28fc0_45, RIbe2ae38_110);
nand \U$23403 ( \23656 , \23654 , \23655 );
xnor \U$23404 ( \23657 , \23656 , RIbe2aeb0_111);
and \U$23405 ( \23658 , \23657 , \1764 );
not \U$23406 ( \23659 , \23657 );
and \U$23407 ( \23660 , \23659 , \1245 );
nor \U$23408 ( \23661 , \23658 , \23660 );
not \U$23409 ( \23662 , \12893 );
not \U$23410 ( \23663 , RIbe296c8_60);
not \U$23411 ( \23664 , \15249 );
or \U$23412 ( \23665 , \23663 , \23664 );
nand \U$23413 ( \23666 , \12794 , RIbe29650_59);
nand \U$23414 ( \23667 , \23665 , \23666 );
not \U$23415 ( \23668 , \23667 );
or \U$23416 ( \23669 , \23662 , \23668 );
or \U$23417 ( \23670 , \23667 , \12998 );
nand \U$23418 ( \23671 , \23669 , \23670 );
xor \U$23419 ( \23672 , \23661 , \23671 );
not \U$23420 ( \23673 , RIbe280c0_13);
not \U$23421 ( \23674 , \13590 );
or \U$23422 ( \23675 , \23673 , \23674 );
nand \U$23423 ( \23676 , \13012 , RIbe29830_63);
nand \U$23424 ( \23677 , \23675 , \23676 );
and \U$23425 ( \23678 , \23677 , \12866 );
not \U$23426 ( \23679 , \23677 );
and \U$23427 ( \23680 , \23679 , \14558 );
nor \U$23428 ( \23681 , \23678 , \23680 );
not \U$23429 ( \23682 , RIbe28228_16);
not \U$23430 ( \23683 , \13074 );
or \U$23431 ( \23684 , \23682 , \23683 );
nand \U$23432 ( \23685 , \13077 , RIbe281b0_15);
nand \U$23433 ( \23686 , \23684 , \23685 );
and \U$23434 ( \23687 , \23686 , \12746 );
not \U$23435 ( \23688 , \23686 );
and \U$23436 ( \23689 , \23688 , \14077 );
nor \U$23437 ( \23690 , \23687 , \23689 );
and \U$23438 ( \23691 , \23681 , \23690 );
not \U$23439 ( \23692 , \23681 );
not \U$23440 ( \23693 , \23690 );
and \U$23441 ( \23694 , \23692 , \23693 );
or \U$23442 ( \23695 , \23691 , \23694 );
not \U$23443 ( \23696 , RIbe28930_31);
not \U$23444 ( \23697 , \19262 );
or \U$23445 ( \23698 , \23696 , \23697 );
nand \U$23446 ( \23699 , \12711 , RIbe29560_57);
nand \U$23447 ( \23700 , \23698 , \23699 );
not \U$23448 ( \23701 , \23700 );
not \U$23449 ( \23702 , \12723 );
and \U$23450 ( \23703 , \23701 , \23702 );
and \U$23451 ( \23704 , \23700 , \12723 );
nor \U$23452 ( \23705 , \23703 , \23704 );
and \U$23453 ( \23706 , \23695 , \23705 );
not \U$23454 ( \23707 , \23695 );
not \U$23455 ( \23708 , \23705 );
and \U$23456 ( \23709 , \23707 , \23708 );
nor \U$23457 ( \23710 , \23706 , \23709 );
and \U$23458 ( \23711 , \23672 , \23710 );
not \U$23459 ( \23712 , \23672 );
not \U$23460 ( \23713 , \23710 );
and \U$23461 ( \23714 , \23712 , \23713 );
nor \U$23462 ( \23715 , \23711 , \23714 );
not \U$23463 ( \23716 , \23715 );
and \U$23464 ( \23717 , \23651 , \23716 );
and \U$23465 ( \23718 , \23650 , \23715 );
nor \U$23466 ( \23719 , \23717 , \23718 );
not \U$23467 ( \23720 , \23719 );
not \U$23468 ( \23721 , \22856 );
not \U$23469 ( \23722 , \22865 );
not \U$23470 ( \23723 , \23722 );
or \U$23471 ( \23724 , \23721 , \23723 );
not \U$23472 ( \23725 , \22856 );
not \U$23473 ( \23726 , \23725 );
not \U$23474 ( \23727 , \22865 );
or \U$23475 ( \23728 , \23726 , \23727 );
not \U$23476 ( \23729 , \22860 );
nand \U$23477 ( \23730 , \23728 , \23729 );
nand \U$23478 ( \23731 , \23724 , \23730 );
not \U$23479 ( \23732 , \23731 );
xor \U$23480 ( \23733 , \22870 , \22874 );
and \U$23481 ( \23734 , \23733 , \22880 );
and \U$23482 ( \23735 , \22870 , \22874 );
or \U$23483 ( \23736 , \23734 , \23735 );
not \U$23484 ( \23737 , \23736 );
not \U$23485 ( \23738 , \23737 );
or \U$23486 ( \23739 , \23732 , \23738 );
or \U$23487 ( \23740 , \23731 , \23737 );
nand \U$23488 ( \23741 , \23739 , \23740 );
not \U$23489 ( \23742 , \22897 );
not \U$23490 ( \23743 , \22908 );
or \U$23491 ( \23744 , \23742 , \23743 );
nand \U$23492 ( \23745 , \23744 , \22889 );
not \U$23493 ( \23746 , \22908 );
nand \U$23494 ( \23747 , \23746 , \22896 );
nand \U$23495 ( \23748 , \23745 , \23747 );
not \U$23496 ( \23749 , \23748 );
and \U$23497 ( \23750 , \23741 , \23749 );
not \U$23498 ( \23751 , \23741 );
and \U$23499 ( \23752 , \23751 , \23748 );
nor \U$23500 ( \23753 , \23750 , \23752 );
not \U$23501 ( \23754 , \23753 );
not \U$23502 ( \23755 , \23754 );
or \U$23503 ( \23756 , \23720 , \23755 );
not \U$23504 ( \23757 , \23719 );
nand \U$23505 ( \23758 , \23757 , \23753 );
nand \U$23506 ( \23759 , \23756 , \23758 );
xor \U$23507 ( \23760 , \23048 , \23077 );
and \U$23508 ( \23761 , \23760 , \23119 );
and \U$23509 ( \23762 , \23048 , \23077 );
or \U$23510 ( \23763 , \23761 , \23762 );
not \U$23511 ( \23764 , \23009 );
not \U$23512 ( \23765 , \22945 );
not \U$23513 ( \23766 , \23765 );
or \U$23514 ( \23767 , \23764 , \23766 );
or \U$23515 ( \23768 , \23765 , \23009 );
nand \U$23516 ( \23769 , \23768 , \22973 );
nand \U$23517 ( \23770 , \23767 , \23769 );
and \U$23518 ( \23771 , \23763 , \23770 );
not \U$23519 ( \23772 , \23763 );
not \U$23520 ( \23773 , \23770 );
and \U$23521 ( \23774 , \23772 , \23773 );
nor \U$23522 ( \23775 , \23771 , \23774 );
not \U$23523 ( \23776 , \23775 );
or \U$23524 ( \23777 , \23184 , \23154 );
and \U$23525 ( \23778 , \23777 , \23213 );
and \U$23526 ( \23779 , \23154 , \23184 );
nor \U$23527 ( \23780 , \23778 , \23779 );
not \U$23528 ( \23781 , \23780 );
and \U$23529 ( \23782 , \23776 , \23781 );
and \U$23530 ( \23783 , \23775 , \23780 );
nor \U$23531 ( \23784 , \23782 , \23783 );
not \U$23532 ( \23785 , \23784 );
and \U$23533 ( \23786 , \23759 , \23785 );
not \U$23534 ( \23787 , \23759 );
and \U$23535 ( \23788 , \23787 , \23784 );
nor \U$23536 ( \23789 , \23786 , \23788 );
not \U$23537 ( \23790 , \23789 );
and \U$23538 ( \23791 , \23537 , \23790 );
not \U$23539 ( \23792 , \23537 );
and \U$23540 ( \23793 , \23792 , \23789 );
nor \U$23541 ( \23794 , \23791 , \23793 );
xor \U$23542 ( \23795 , \23258 , \23794 );
xnor \U$23543 ( \23796 , \23249 , \23795 );
xor \U$23544 ( \23797 , \23232 , \23796 );
not \U$23545 ( \23798 , \22672 );
not \U$23546 ( \23799 , \22668 );
or \U$23547 ( \23800 , \23798 , \23799 );
or \U$23548 ( \23801 , \22668 , \22672 );
nand \U$23549 ( \23802 , \23800 , \23801 );
xor \U$23550 ( \23803 , \22710 , \23802 );
not \U$23551 ( \23804 , RIbe2a988_100);
not \U$23552 ( \23805 , \12268 );
or \U$23553 ( \23806 , \23804 , \23805 );
nand \U$23554 ( \23807 , \8235 , RIbe2a910_99);
nand \U$23555 ( \23808 , \23806 , \23807 );
and \U$23556 ( \23809 , \23808 , \9944 );
not \U$23557 ( \23810 , \23808 );
and \U$23558 ( \23811 , \23810 , \7534 );
nor \U$23559 ( \23812 , \23809 , \23811 );
not \U$23560 ( \23813 , \23812 );
not \U$23561 ( \23814 , \23813 );
not \U$23562 ( \23815 , RIbe2a370_87);
not \U$23563 ( \23816 , \20487 );
or \U$23564 ( \23817 , \23815 , \23816 );
nand \U$23565 ( \23818 , \7483 , RIbe2a2f8_86);
nand \U$23566 ( \23819 , \23817 , \23818 );
and \U$23567 ( \23820 , \23819 , \14666 );
not \U$23568 ( \23821 , \23819 );
and \U$23569 ( \23822 , \23821 , \6582 );
nor \U$23570 ( \23823 , \23820 , \23822 );
not \U$23571 ( \23824 , \23823 );
not \U$23572 ( \23825 , \23824 );
or \U$23573 ( \23826 , \23814 , \23825 );
not \U$23574 ( \23827 , \23823 );
not \U$23575 ( \23828 , \23812 );
or \U$23576 ( \23829 , \23827 , \23828 );
not \U$23577 ( \23830 , \6891 );
not \U$23578 ( \23831 , RIbe2b5b8_126);
not \U$23579 ( \23832 , \6535 );
or \U$23580 ( \23833 , \23831 , \23832 );
nand \U$23581 ( \23834 , \6540 , RIbe2a3e8_88);
nand \U$23582 ( \23835 , \23833 , \23834 );
not \U$23583 ( \23836 , \23835 );
or \U$23584 ( \23837 , \23830 , \23836 );
or \U$23585 ( \23838 , \23835 , \6888 );
nand \U$23586 ( \23839 , \23837 , \23838 );
nand \U$23587 ( \23840 , \23829 , \23839 );
nand \U$23588 ( \23841 , \23826 , \23840 );
not \U$23589 ( \23842 , RIbe2a5c8_92);
not \U$23590 ( \23843 , \6630 );
or \U$23591 ( \23844 , \23842 , \23843 );
nand \U$23592 ( \23845 , \15885 , RIbe2a550_91);
nand \U$23593 ( \23846 , \23844 , \23845 );
and \U$23594 ( \23847 , \23846 , \6640 );
not \U$23595 ( \23848 , \23846 );
and \U$23596 ( \23849 , \23848 , \10272 );
nor \U$23597 ( \23850 , \23847 , \23849 );
not \U$23598 ( \23851 , \23850 );
not \U$23599 ( \23852 , \23851 );
not \U$23600 ( \23853 , RIbe2b090_115);
not \U$23601 ( \23854 , \4595 );
or \U$23602 ( \23855 , \23853 , \23854 );
nand \U$23603 ( \23856 , \7858 , RIbe2a280_85);
nand \U$23604 ( \23857 , \23855 , \23856 );
and \U$23605 ( \23858 , \23857 , \4323 );
not \U$23606 ( \23859 , \23857 );
and \U$23607 ( \23860 , \23859 , \4326 );
nor \U$23608 ( \23861 , \23858 , \23860 );
not \U$23609 ( \23862 , \23861 );
not \U$23610 ( \23863 , \23862 );
or \U$23611 ( \23864 , \23852 , \23863 );
and \U$23612 ( \23865 , \4826 , RIbe2a208_84);
or \U$23613 ( \23866 , \5052 , \23865 );
not \U$23614 ( \23867 , RIbe2a190_83);
nand \U$23615 ( \23868 , \23867 , \22378 );
nand \U$23616 ( \23869 , \23866 , \23868 );
not \U$23617 ( \23870 , \23869 );
not \U$23618 ( \23871 , \4586 );
and \U$23619 ( \23872 , \23870 , \23871 );
and \U$23620 ( \23873 , \23869 , \4586 );
nor \U$23621 ( \23874 , \23872 , \23873 );
not \U$23622 ( \23875 , \23874 );
nand \U$23623 ( \23876 , \23861 , \23850 );
nand \U$23624 ( \23877 , \23875 , \23876 );
nand \U$23625 ( \23878 , \23864 , \23877 );
or \U$23626 ( \23879 , \23841 , \23878 );
not \U$23627 ( \23880 , RIbe2acd0_107);
not \U$23628 ( \23881 , \8199 );
or \U$23629 ( \23882 , \23880 , \23881 );
nand \U$23630 ( \23883 , \6963 , RIbe2a028_80);
nand \U$23631 ( \23884 , \23882 , \23883 );
and \U$23632 ( \23885 , \23884 , \7293 );
not \U$23633 ( \23886 , \23884 );
and \U$23634 ( \23887 , \23886 , \6572 );
nor \U$23635 ( \23888 , \23885 , \23887 );
not \U$23636 ( \23889 , \23888 );
nand \U$23637 ( \23890 , \7981 , RIbe29c68_72);
nand \U$23638 ( \23891 , \6939 , RIbe2a0a0_81, RIbe2b360_121, RIbe29dd0_75);
nor \U$23639 ( \23892 , RIbe2a0a0_81, RIbe2b360_121);
nand \U$23640 ( \23893 , \6939 , \23892 , RIbe29dd0_75);
nand \U$23641 ( \23894 , \23890 , \23891 , \23893 );
and \U$23642 ( \23895 , \23894 , \16010 );
not \U$23643 ( \23896 , \23894 );
and \U$23644 ( \23897 , \23896 , \7984 );
nor \U$23645 ( \23898 , \23895 , \23897 );
not \U$23646 ( \23899 , \23898 );
or \U$23647 ( \23900 , \23889 , \23899 );
or \U$23648 ( \23901 , \23888 , \23898 );
and \U$23649 ( \23902 , \7298 , RIbe29fb0_79);
and \U$23650 ( \23903 , \6983 , RIbe29e48_76);
nor \U$23651 ( \23904 , \23902 , \23903 );
and \U$23652 ( \23905 , \23904 , \6992 );
not \U$23653 ( \23906 , \23904 );
and \U$23654 ( \23907 , \23906 , \7660 );
nor \U$23655 ( \23908 , \23905 , \23907 );
nand \U$23656 ( \23909 , \23901 , \23908 );
nand \U$23657 ( \23910 , \23900 , \23909 );
nand \U$23658 ( \23911 , \23879 , \23910 );
nand \U$23659 ( \23912 , \23841 , \23878 );
nand \U$23660 ( \23913 , \23911 , \23912 );
not \U$23661 ( \23914 , \23913 );
not \U$23662 ( \23915 , RIbe29290_51);
not \U$23663 ( \23916 , \12786 );
or \U$23664 ( \23917 , \23915 , \23916 );
nand \U$23665 ( \23918 , \12794 , RIbe28a20_33);
nand \U$23666 ( \23919 , \23917 , \23918 );
and \U$23667 ( \23920 , \23919 , \14335 );
not \U$23668 ( \23921 , \23919 );
and \U$23669 ( \23922 , \23921 , \14336 );
nor \U$23670 ( \23923 , \23920 , \23922 );
not \U$23671 ( \23924 , RIbe289a8_32);
not \U$23672 ( \23925 , \13690 );
or \U$23673 ( \23926 , \23924 , \23925 );
nand \U$23674 ( \23927 , RIbe28930_31, RIbe2ae38_110);
nand \U$23675 ( \23928 , \23926 , \23927 );
xnor \U$23676 ( \23929 , \23928 , RIbe2aeb0_111);
nand \U$23677 ( \23930 , \23923 , \23929 );
not \U$23678 ( \23931 , \12863 );
not \U$23679 ( \23932 , RIbe28b10_35);
not \U$23680 ( \23933 , \12858 );
or \U$23681 ( \23934 , \23932 , \23933 );
nand \U$23682 ( \23935 , \13012 , RIbe28b88_36);
nand \U$23683 ( \23936 , \23934 , \23935 );
not \U$23684 ( \23937 , \23936 );
or \U$23685 ( \23938 , \23931 , \23937 );
or \U$23686 ( \23939 , \23936 , \12823 );
nand \U$23687 ( \23940 , \23938 , \23939 );
and \U$23688 ( \23941 , \23930 , \23940 );
nor \U$23689 ( \23942 , \23923 , \23929 );
nor \U$23690 ( \23943 , \23941 , \23942 );
not \U$23691 ( \23944 , \23943 );
not \U$23692 ( \23945 , RIbe28408_20);
not \U$23693 ( \23946 , \14534 );
or \U$23694 ( \23947 , \23945 , \23946 );
nand \U$23695 ( \23948 , \12735 , RIbe28390_19);
nand \U$23696 ( \23949 , \23947 , \23948 );
and \U$23697 ( \23950 , \23949 , \14542 );
not \U$23698 ( \23951 , \23949 );
and \U$23699 ( \23952 , \23951 , \16754 );
nor \U$23700 ( \23953 , \23950 , \23952 );
not \U$23701 ( \23954 , RIbe287c8_28);
not \U$23702 ( \23955 , \16759 );
or \U$23703 ( \23956 , \23954 , \23955 );
nand \U$23704 ( \23957 , \12710 , RIbe28480_21);
nand \U$23705 ( \23958 , \23956 , \23957 );
and \U$23706 ( \23959 , \23958 , \12723 );
not \U$23707 ( \23960 , \23958 );
and \U$23708 ( \23961 , \23960 , \12879 );
nor \U$23709 ( \23962 , \23959 , \23961 );
nand \U$23710 ( \23963 , \23953 , \23962 );
not \U$23711 ( \23964 , \12770 );
not \U$23712 ( \23965 , RIbe28660_25);
not \U$23713 ( \23966 , \12921 );
or \U$23714 ( \23967 , \23965 , \23966 );
nand \U$23715 ( \23968 , \17715 , RIbe285e8_24);
nand \U$23716 ( \23969 , \23967 , \23968 );
not \U$23717 ( \23970 , \23969 );
or \U$23718 ( \23971 , \23964 , \23970 );
or \U$23719 ( \23972 , \23969 , \12924 );
nand \U$23720 ( \23973 , \23971 , \23972 );
and \U$23721 ( \23974 , \23963 , \23973 );
nor \U$23722 ( \23975 , \23953 , \23962 );
nor \U$23723 ( \23976 , \23974 , \23975 );
not \U$23724 ( \23977 , \23976 );
or \U$23725 ( \23978 , \23944 , \23977 );
not \U$23726 ( \23979 , RIbe28ed0_43);
not \U$23727 ( \23980 , \20530 );
or \U$23728 ( \23981 , \23979 , \23980 );
nand \U$23729 ( \23982 , RIbe27fd0_11, \12212 );
nand \U$23730 ( \23983 , \23981 , \23982 );
and \U$23731 ( \23984 , \23983 , \19139 );
not \U$23732 ( \23985 , \23983 );
and \U$23733 ( \23986 , \23985 , \10943 );
nor \U$23734 ( \23987 , \23984 , \23986 );
not \U$23735 ( \23988 , RIbe27f58_10);
not \U$23736 ( \23989 , \12942 );
or \U$23737 ( \23990 , \23988 , \23989 );
nand \U$23738 ( \23991 , \12948 , RIbe27e68_8);
nand \U$23739 ( \23992 , \23990 , \23991 );
and \U$23740 ( \23993 , \23992 , \12195 );
not \U$23741 ( \23994 , \23992 );
and \U$23742 ( \23995 , \23994 , \12956 );
nor \U$23743 ( \23996 , \23993 , \23995 );
xor \U$23744 ( \23997 , \23987 , \23996 );
and \U$23745 ( \23998 , \13478 , RIbe29bf0_71);
and \U$23746 ( \23999 , \13038 , RIbe28f48_44);
nor \U$23747 ( \24000 , \23998 , \23999 );
and \U$23748 ( \24001 , \24000 , \10912 );
not \U$23749 ( \24002 , \24000 );
and \U$23750 ( \24003 , \24002 , \7970 );
nor \U$23751 ( \24004 , \24001 , \24003 );
and \U$23752 ( \24005 , \23997 , \24004 );
and \U$23753 ( \24006 , \23987 , \23996 );
or \U$23754 ( \24007 , \24005 , \24006 );
nand \U$23755 ( \24008 , \23978 , \24007 );
not \U$23756 ( \24009 , \23976 );
not \U$23757 ( \24010 , \23943 );
nand \U$23758 ( \24011 , \24009 , \24010 );
nand \U$23759 ( \24012 , \24008 , \24011 );
not \U$23760 ( \24013 , \24012 );
and \U$23761 ( \24014 , \23914 , \24013 );
nand \U$23762 ( \24015 , \1099 , RIbe2ab68_104);
and \U$23763 ( \24016 , \24015 , \1309 );
not \U$23764 ( \24017 , \24015 );
and \U$23765 ( \24018 , \24017 , \4251 );
nor \U$23766 ( \24019 , \24016 , \24018 );
not \U$23767 ( \24020 , RIbe2afa0_113);
not \U$23768 ( \24021 , \8342 );
or \U$23769 ( \24022 , \24020 , \24021 );
nand \U$23770 ( \24023 , \2901 , RIbe2af28_112);
nand \U$23771 ( \24024 , \24022 , \24023 );
not \U$23772 ( \24025 , \24024 );
not \U$23773 ( \24026 , \2576 );
and \U$23774 ( \24027 , \24025 , \24026 );
and \U$23775 ( \24028 , \24024 , \4059 );
nor \U$23776 ( \24029 , \24027 , \24028 );
not \U$23777 ( \24030 , RIbe2b270_119);
not \U$23778 ( \24031 , \7880 );
or \U$23779 ( \24032 , \24030 , \24031 );
nand \U$23780 ( \24033 , \6787 , RIbe2b108_116);
nand \U$23781 ( \24034 , \24032 , \24033 );
and \U$23782 ( \24035 , \24034 , \3448 );
not \U$23783 ( \24036 , \24034 );
and \U$23784 ( \24037 , \24036 , \3471 );
nor \U$23785 ( \24038 , \24035 , \24037 );
and \U$23786 ( \24039 , \24029 , \24038 );
not \U$23787 ( \24040 , RIbe2b1f8_118);
not \U$23788 ( \24041 , \3685 );
or \U$23789 ( \24042 , \24040 , \24041 );
nand \U$23790 ( \24043 , \3689 , RIbe2b180_117);
nand \U$23791 ( \24044 , \24042 , \24043 );
and \U$23792 ( \24045 , \24044 , \2887 );
not \U$23793 ( \24046 , \24044 );
and \U$23794 ( \24047 , \24046 , \3290 );
nor \U$23795 ( \24048 , \24045 , \24047 );
nor \U$23796 ( \24049 , \24039 , \24048 );
nor \U$23797 ( \24050 , \24029 , \24038 );
nor \U$23798 ( \24051 , \24049 , \24050 );
xor \U$23799 ( \24052 , \24019 , \24051 );
and \U$23800 ( \24053 , \1112 , RIbe2aaf0_103);
and \U$23801 ( \24054 , \20663 , RIbe2b630_127);
nor \U$23802 ( \24055 , \24053 , \24054 );
and \U$23803 ( \24056 , \24055 , \1132 );
not \U$23804 ( \24057 , \24055 );
and \U$23805 ( \24058 , \24057 , \1448 );
nor \U$23806 ( \24059 , \24056 , \24058 );
and \U$23807 ( \24060 , \1272 , RIbe2b018_114);
and \U$23808 ( \24061 , \2384 , RIbe2afa0_113);
nor \U$23809 ( \24062 , \24060 , \24061 );
not \U$23810 ( \24063 , \1275 );
xor \U$23811 ( \24064 , \24062 , \24063 );
xor \U$23812 ( \24065 , \24059 , \24064 );
not \U$23813 ( \24066 , RIbe2af28_112);
not \U$23814 ( \24067 , \8342 );
or \U$23815 ( \24068 , \24066 , \24067 );
nand \U$23816 ( \24069 , \3267 , RIbe2b1f8_118);
nand \U$23817 ( \24070 , \24068 , \24069 );
and \U$23818 ( \24071 , \24070 , \3275 );
not \U$23819 ( \24072 , \24070 );
and \U$23820 ( \24073 , \24072 , \4058 );
nor \U$23821 ( \24074 , \24071 , \24073 );
xor \U$23822 ( \24075 , \24065 , \24074 );
and \U$23823 ( \24076 , \24052 , \24075 );
and \U$23824 ( \24077 , \24019 , \24051 );
or \U$23825 ( \24078 , \24076 , \24077 );
nor \U$23826 ( \24079 , \24014 , \24078 );
and \U$23827 ( \24080 , \24012 , \23913 );
nor \U$23828 ( \24081 , \24079 , \24080 );
and \U$23829 ( \24082 , \22554 , \22543 );
not \U$23830 ( \24083 , \22554 );
and \U$23831 ( \24084 , \24083 , \22569 );
nor \U$23832 ( \24085 , \24082 , \24084 );
xnor \U$23833 ( \24086 , \24085 , \22566 );
nand \U$23834 ( \24087 , \6557 , RIbe2a028_80);
or \U$23835 ( \24088 , \6961 , \24087 );
nand \U$23836 ( \24089 , RIbe29fb0_79, \7957 );
nand \U$23837 ( \24090 , \24088 , \24089 );
and \U$23838 ( \24091 , \24090 , \7293 );
not \U$23839 ( \24092 , \24090 );
and \U$23840 ( \24093 , \24092 , \6572 );
nor \U$23841 ( \24094 , \24091 , \24093 );
and \U$23842 ( \24095 , \7277 , RIbe2acd0_107);
not \U$23843 ( \24096 , \7277 );
and \U$23844 ( \24097 , \6588 , RIbe2a2f8_86);
and \U$23845 ( \24098 , \24096 , \24097 );
or \U$23846 ( \24099 , \24095 , \24098 );
and \U$23847 ( \24100 , \24099 , \6582 );
not \U$23848 ( \24101 , \24099 );
and \U$23849 ( \24102 , \24101 , \6873 );
nor \U$23850 ( \24103 , \24100 , \24102 );
xor \U$23851 ( \24104 , \24094 , \24103 );
not \U$23852 ( \24105 , RIbe2a3e8_88);
not \U$23853 ( \24106 , \6535 );
or \U$23854 ( \24107 , \24105 , \24106 );
nand \U$23855 ( \24108 , \6884 , RIbe2a370_87);
nand \U$23856 ( \24109 , \24107 , \24108 );
not \U$23857 ( \24110 , \24109 );
not \U$23858 ( \24111 , \6891 );
and \U$23859 ( \24112 , \24110 , \24111 );
and \U$23860 ( \24113 , \24109 , \6551 );
nor \U$23861 ( \24114 , \24112 , \24113 );
not \U$23862 ( \24115 , \24114 );
and \U$23863 ( \24116 , \24104 , \24115 );
not \U$23864 ( \24117 , \24104 );
and \U$23865 ( \24118 , \24117 , \24114 );
nor \U$23866 ( \24119 , \24116 , \24118 );
not \U$23867 ( \24120 , RIbe2a190_83);
not \U$23868 ( \24121 , \21097 );
or \U$23869 ( \24122 , \24120 , \24121 );
nand \U$23870 ( \24123 , \7056 , RIbe2a5c8_92);
nand \U$23871 ( \24124 , \24122 , \24123 );
xor \U$23872 ( \24125 , \24124 , \4592 );
not \U$23873 ( \24126 , \24125 );
nand \U$23874 ( \24127 , \5748 , RIbe2a988_100);
not \U$23875 ( \24128 , \24127 );
nor \U$23876 ( \24129 , \5044 , \5453 );
not \U$23877 ( \24130 , \24129 );
or \U$23878 ( \24131 , \24128 , \24130 );
nand \U$23879 ( \24132 , \6634 , \24127 , \5460 );
nand \U$23880 ( \24133 , \24131 , \24132 );
or \U$23881 ( \24134 , \24127 , \5045 );
nand \U$23882 ( \24135 , \5453 , RIbe2a550_91);
or \U$23883 ( \24136 , \5749 , \24135 , \5460 );
nand \U$23884 ( \24137 , \24127 , \5460 , \21491 );
nand \U$23885 ( \24138 , \24134 , \24136 , \24137 );
nor \U$23886 ( \24139 , \24133 , \24138 );
and \U$23887 ( \24140 , \8234 , RIbe2b5b8_126);
not \U$23888 ( \24141 , \8234 );
and \U$23889 ( \24142 , \6134 , RIbe2a910_99);
and \U$23890 ( \24143 , \24141 , \24142 );
or \U$23891 ( \24144 , \24140 , \24143 );
and \U$23892 ( \24145 , \24144 , \21090 );
not \U$23893 ( \24146 , \24144 );
and \U$23894 ( \24147 , \24146 , \21093 );
nor \U$23895 ( \24148 , \24145 , \24147 );
and \U$23896 ( \24149 , \24139 , \24148 );
not \U$23897 ( \24150 , \24139 );
not \U$23898 ( \24151 , \24148 );
and \U$23899 ( \24152 , \24150 , \24151 );
nor \U$23900 ( \24153 , \24149 , \24152 );
not \U$23901 ( \24154 , \24153 );
or \U$23902 ( \24155 , \24126 , \24154 );
or \U$23903 ( \24156 , \24125 , \24153 );
nand \U$23904 ( \24157 , \24155 , \24156 );
xor \U$23905 ( \24158 , \24119 , \24157 );
and \U$23906 ( \24159 , \4314 , RIbe2a280_85);
not \U$23907 ( \24160 , \24159 );
not \U$23908 ( \24161 , \4807 );
or \U$23909 ( \24162 , \24160 , \24161 );
not \U$23910 ( \24163 , \13156 );
nand \U$23911 ( \24164 , \24163 , \21043 );
nand \U$23912 ( \24165 , \24162 , \24164 );
and \U$23913 ( \24166 , \24165 , \4326 );
not \U$23914 ( \24167 , \24165 );
and \U$23915 ( \24168 , \24167 , \7865 );
nor \U$23916 ( \24169 , \24166 , \24168 );
not \U$23917 ( \24170 , RIbe2b108_116);
not \U$23918 ( \24171 , \20764 );
or \U$23919 ( \24172 , \24170 , \24171 );
nand \U$23920 ( \24173 , \20767 , RIbe2b090_115);
nand \U$23921 ( \24174 , \24172 , \24173 );
not \U$23922 ( \24175 , \24174 );
not \U$23923 ( \24176 , \3698 );
and \U$23924 ( \24177 , \24175 , \24176 );
and \U$23925 ( \24178 , \24174 , \3448 );
nor \U$23926 ( \24179 , \24177 , \24178 );
xor \U$23927 ( \24180 , \24169 , \24179 );
not \U$23928 ( \24181 , RIbe2b180_117);
not \U$23929 ( \24182 , \3451 );
or \U$23930 ( \24183 , \24181 , \24182 );
nand \U$23931 ( \24184 , \4011 , RIbe2b270_119);
nand \U$23932 ( \24185 , \24183 , \24184 );
and \U$23933 ( \24186 , \24185 , \3290 );
not \U$23934 ( \24187 , \24185 );
and \U$23935 ( \24188 , \24187 , \3461 );
nor \U$23936 ( \24189 , \24186 , \24188 );
xnor \U$23937 ( \24190 , \24180 , \24189 );
and \U$23938 ( \24191 , \24158 , \24190 );
and \U$23939 ( \24192 , \24119 , \24157 );
or \U$23940 ( \24193 , \24191 , \24192 );
not \U$23941 ( \24194 , \24193 );
xor \U$23942 ( \24195 , \24086 , \24194 );
and \U$23943 ( \24196 , \20405 , RIbe28f48_44);
and \U$23944 ( \24197 , \10919 , RIbe28ed0_43);
nor \U$23945 ( \24198 , \24196 , \24197 );
and \U$23946 ( \24199 , \24198 , \7970 );
not \U$23947 ( \24200 , \24198 );
and \U$23948 ( \24201 , \24200 , \8077 );
nor \U$23949 ( \24202 , \24199 , \24201 );
not \U$23950 ( \24203 , RIbe29c68_72);
not \U$23951 ( \24204 , \7974 );
or \U$23952 ( \24205 , \24203 , \24204 );
nand \U$23953 ( \24206 , \8269 , RIbe29bf0_71);
nand \U$23954 ( \24207 , \24205 , \24206 );
not \U$23955 ( \24208 , \24207 );
not \U$23956 ( \24209 , \7984 );
and \U$23957 ( \24210 , \24208 , \24209 );
and \U$23958 ( \24211 , \24207 , \6949 );
nor \U$23959 ( \24212 , \24210 , \24211 );
xor \U$23960 ( \24213 , \24202 , \24212 );
not \U$23961 ( \24214 , RIbe29e48_76);
not \U$23962 ( \24215 , \7298 );
or \U$23963 ( \24216 , \24214 , \24215 );
nand \U$23964 ( \24217 , \13792 , RIbe29dd0_75);
nand \U$23965 ( \24218 , \24216 , \24217 );
not \U$23966 ( \24219 , \24218 );
not \U$23967 ( \24220 , \7301 );
and \U$23968 ( \24221 , \24219 , \24220 );
and \U$23969 ( \24222 , \24218 , \6992 );
nor \U$23970 ( \24223 , \24221 , \24222 );
xor \U$23971 ( \24224 , \24213 , \24223 );
not \U$23972 ( \24225 , RIbe28b88_36);
not \U$23973 ( \24226 , \14550 );
or \U$23974 ( \24227 , \24225 , \24226 );
nand \U$23975 ( \24228 , \12834 , RIbe29290_51);
nand \U$23976 ( \24229 , \24227 , \24228 );
not \U$23977 ( \24230 , \24229 );
not \U$23978 ( \24231 , \16366 );
and \U$23979 ( \24232 , \24230 , \24231 );
and \U$23980 ( \24233 , \24229 , \16366 );
nor \U$23981 ( \24234 , \24232 , \24233 );
not \U$23982 ( \24235 , \24234 );
not \U$23983 ( \24236 , RIbe28390_19);
not \U$23984 ( \24237 , \15161 );
or \U$23985 ( \24238 , \24236 , \24237 );
nand \U$23986 ( \24239 , \12735 , RIbe28b10_35);
nand \U$23987 ( \24240 , \24238 , \24239 );
and \U$23988 ( \24241 , \24240 , \15166 );
not \U$23989 ( \24242 , \24240 );
and \U$23990 ( \24243 , \24242 , \12742 );
nor \U$23991 ( \24244 , \24241 , \24243 );
not \U$23992 ( \24245 , \24244 );
or \U$23993 ( \24246 , \24235 , \24245 );
or \U$23994 ( \24247 , \24244 , \24234 );
nand \U$23995 ( \24248 , \24246 , \24247 );
not \U$23996 ( \24249 , RIbe28480_21);
not \U$23997 ( \24250 , \19262 );
or \U$23998 ( \24251 , \24249 , \24250 );
nand \U$23999 ( \24252 , \12710 , RIbe28408_20);
nand \U$24000 ( \24253 , \24251 , \24252 );
xor \U$24001 ( \24254 , \24253 , \12723 );
and \U$24002 ( \24255 , \24248 , \24254 );
not \U$24003 ( \24256 , \24248 );
not \U$24004 ( \24257 , \24254 );
and \U$24005 ( \24258 , \24256 , \24257 );
nor \U$24006 ( \24259 , \24255 , \24258 );
nand \U$24007 ( \24260 , \24224 , \24259 );
not \U$24008 ( \24261 , \12774 );
not \U$24009 ( \24262 , \13087 );
not \U$24010 ( \24263 , \10854 );
and \U$24011 ( \24264 , \24262 , \24263 );
and \U$24012 ( \24265 , \12764 , RIbe285e8_24);
nor \U$24013 ( \24266 , \24264 , \24265 );
not \U$24014 ( \24267 , \24266 );
or \U$24015 ( \24268 , \24261 , \24267 );
or \U$24016 ( \24269 , \24266 , \12927 );
nand \U$24017 ( \24270 , \24268 , \24269 );
not \U$24018 ( \24271 , RIbe27e68_8);
not \U$24019 ( \24272 , \12943 );
or \U$24020 ( \24273 , \24271 , \24272 );
nand \U$24021 ( \24274 , \12948 , RIbe28660_25);
nand \U$24022 ( \24275 , \24273 , \24274 );
and \U$24023 ( \24276 , \24275 , \12195 );
not \U$24024 ( \24277 , \24275 );
and \U$24025 ( \24278 , \24277 , \17005 );
nor \U$24026 ( \24279 , \24276 , \24278 );
xor \U$24027 ( \24280 , \24270 , \24279 );
not \U$24028 ( \24281 , RIbe27fd0_11);
not \U$24029 ( \24282 , \10936 );
or \U$24030 ( \24283 , \24281 , \24282 );
nand \U$24031 ( \24284 , \12212 , RIbe27f58_10);
nand \U$24032 ( \24285 , \24283 , \24284 );
and \U$24033 ( \24286 , \24285 , \9902 );
not \U$24034 ( \24287 , \24285 );
and \U$24035 ( \24288 , \24287 , \13033 );
nor \U$24036 ( \24289 , \24286 , \24288 );
xor \U$24037 ( \24290 , \24280 , \24289 );
and \U$24038 ( \24291 , \24260 , \24290 );
nor \U$24039 ( \24292 , \24224 , \24259 );
nor \U$24040 ( \24293 , \24291 , \24292 );
and \U$24041 ( \24294 , \24195 , \24293 );
and \U$24042 ( \24295 , \24086 , \24194 );
or \U$24043 ( \24296 , \24294 , \24295 );
xor \U$24044 ( \24297 , \24081 , \24296 );
xor \U$24045 ( \24298 , \24059 , \24064 );
and \U$24046 ( \24299 , \24298 , \24074 );
and \U$24047 ( \24300 , \24059 , \24064 );
or \U$24048 ( \24301 , \24299 , \24300 );
xor \U$24049 ( \24302 , \22463 , \22442 );
xnor \U$24050 ( \24303 , \24302 , \22452 );
xor \U$24051 ( \24304 , \24301 , \24303 );
not \U$24052 ( \24305 , \24189 );
not \U$24053 ( \24306 , \24169 );
and \U$24054 ( \24307 , \24305 , \24306 );
nor \U$24055 ( \24308 , \24307 , \24179 );
nor \U$24056 ( \24309 , \24305 , \24306 );
nor \U$24057 ( \24310 , \24308 , \24309 );
xor \U$24058 ( \24311 , \24304 , \24310 );
not \U$24059 ( \24312 , \22473 );
not \U$24060 ( \24313 , \22495 );
or \U$24061 ( \24314 , \24312 , \24313 );
or \U$24062 ( \24315 , \22473 , \22495 );
nand \U$24063 ( \24316 , \24314 , \24315 );
not \U$24064 ( \24317 , \24316 );
not \U$24065 ( \24318 , \22483 );
and \U$24066 ( \24319 , \24317 , \24318 );
and \U$24067 ( \24320 , \24316 , \22483 );
nor \U$24068 ( \24321 , \24319 , \24320 );
not \U$24069 ( \24322 , \24321 );
not \U$24070 ( \24323 , \22415 );
not \U$24071 ( \24324 , \22405 );
or \U$24072 ( \24325 , \24323 , \24324 );
or \U$24073 ( \24326 , \22415 , \22405 );
nand \U$24074 ( \24327 , \24325 , \24326 );
not \U$24075 ( \24328 , \22396 );
and \U$24076 ( \24329 , \24327 , \24328 );
not \U$24077 ( \24330 , \24327 );
and \U$24078 ( \24331 , \24330 , \22396 );
nor \U$24079 ( \24332 , \24329 , \24331 );
not \U$24080 ( \24333 , \24332 );
or \U$24081 ( \24334 , \24322 , \24333 );
or \U$24082 ( \24335 , \24321 , \24332 );
nand \U$24083 ( \24336 , \24334 , \24335 );
xor \U$24084 ( \24337 , \22371 , \22384 );
xnor \U$24085 ( \24338 , \24337 , \22360 );
not \U$24086 ( \24339 , \24338 );
and \U$24087 ( \24340 , \24336 , \24339 );
not \U$24088 ( \24341 , \24336 );
and \U$24089 ( \24342 , \24341 , \24338 );
nor \U$24090 ( \24343 , \24340 , \24342 );
not \U$24091 ( \24344 , \24343 );
and \U$24092 ( \24345 , \24311 , \24344 );
not \U$24093 ( \24346 , \22348 );
not \U$24094 ( \24347 , \22334 );
or \U$24095 ( \24348 , \24346 , \24347 );
nand \U$24096 ( \24349 , \22331 , \22347 );
nand \U$24097 ( \24350 , \24348 , \24349 );
and \U$24098 ( \24351 , \24350 , \22320 );
not \U$24099 ( \24352 , \24350 );
and \U$24100 ( \24353 , \24352 , \22321 );
nor \U$24101 ( \24354 , \24351 , \24353 );
not \U$24102 ( \24355 , \24354 );
not \U$24103 ( \24356 , \24355 );
xor \U$24104 ( \24357 , \22514 , \22524 );
xor \U$24105 ( \24358 , \24357 , \22532 );
not \U$24106 ( \24359 , \24358 );
or \U$24107 ( \24360 , \24356 , \24359 );
not \U$24108 ( \24361 , \24358 );
nand \U$24109 ( \24362 , \24354 , \24361 );
nand \U$24110 ( \24363 , \24360 , \24362 );
not \U$24111 ( \24364 , \22588 );
not \U$24112 ( \24365 , \22581 );
or \U$24113 ( \24366 , \24364 , \24365 );
or \U$24114 ( \24367 , \22588 , \22581 );
nand \U$24115 ( \24368 , \24366 , \24367 );
not \U$24116 ( \24369 , \22600 );
and \U$24117 ( \24370 , \24368 , \24369 );
not \U$24118 ( \24371 , \24368 );
and \U$24119 ( \24372 , \24371 , \22600 );
nor \U$24120 ( \24373 , \24370 , \24372 );
and \U$24121 ( \24374 , \24363 , \24373 );
not \U$24122 ( \24375 , \24363 );
not \U$24123 ( \24376 , \24373 );
and \U$24124 ( \24377 , \24375 , \24376 );
nor \U$24125 ( \24378 , \24374 , \24377 );
nor \U$24126 ( \24379 , \24345 , \24378 );
nor \U$24127 ( \24380 , \24311 , \24344 );
nor \U$24128 ( \24381 , \24379 , \24380 );
and \U$24129 ( \24382 , \24297 , \24381 );
and \U$24130 ( \24383 , \24081 , \24296 );
or \U$24131 ( \24384 , \24382 , \24383 );
not \U$24132 ( \24385 , \24384 );
not \U$24133 ( \24386 , \24385 );
or \U$24134 ( \24387 , \24103 , \24094 );
and \U$24135 ( \24388 , \24115 , \24387 );
and \U$24136 ( \24389 , \24094 , \24103 );
nor \U$24137 ( \24390 , \24388 , \24389 );
not \U$24138 ( \24391 , \24390 );
xor \U$24139 ( \24392 , \24202 , \24212 );
and \U$24140 ( \24393 , \24392 , \24223 );
and \U$24141 ( \24394 , \24202 , \24212 );
or \U$24142 ( \24395 , \24393 , \24394 );
not \U$24143 ( \24396 , \24395 );
or \U$24144 ( \24397 , \24391 , \24396 );
not \U$24145 ( \24398 , \24125 );
not \U$24146 ( \24399 , \24148 );
or \U$24147 ( \24400 , \24398 , \24399 );
not \U$24148 ( \24401 , \24139 );
nand \U$24149 ( \24402 , \24400 , \24401 );
not \U$24150 ( \24403 , \24125 );
nand \U$24151 ( \24404 , \24403 , \24151 );
nand \U$24152 ( \24405 , \24402 , \24404 );
nand \U$24153 ( \24406 , \24397 , \24405 );
not \U$24154 ( \24407 , \24390 );
not \U$24155 ( \24408 , \24395 );
nand \U$24156 ( \24409 , \24407 , \24408 );
nand \U$24157 ( \24410 , \24406 , \24409 );
not \U$24158 ( \24411 , RIbe28a20_33);
not \U$24159 ( \24412 , \12887 );
or \U$24160 ( \24413 , \24411 , \24412 );
nand \U$24161 ( \24414 , \12794 , RIbe289a8_32);
nand \U$24162 ( \24415 , \24413 , \24414 );
xor \U$24163 ( \24416 , \24415 , \12801 );
not \U$24164 ( \24417 , RIbe28930_31);
not \U$24165 ( \24418 , \13003 );
or \U$24166 ( \24419 , \24417 , \24418 );
nand \U$24167 ( \24420 , RIbe29560_57, RIbe2ae38_110);
nand \U$24168 ( \24421 , \24419 , \24420 );
xor \U$24169 ( \24422 , \24421 , RIbe2aeb0_111);
nor \U$24170 ( \24423 , \24422 , \1309 );
or \U$24171 ( \24424 , \24416 , \24423 );
nand \U$24172 ( \24425 , \24422 , \1309 );
nand \U$24173 ( \24426 , \24424 , \24425 );
not \U$24174 ( \24427 , \24234 );
not \U$24175 ( \24428 , \24254 );
or \U$24176 ( \24429 , \24427 , \24428 );
nand \U$24177 ( \24430 , \24429 , \24244 );
not \U$24178 ( \24431 , \24234 );
nand \U$24179 ( \24432 , \24431 , \24257 );
nand \U$24180 ( \24433 , \24430 , \24432 );
xor \U$24181 ( \24434 , \24426 , \24433 );
xor \U$24182 ( \24435 , \24270 , \24279 );
and \U$24183 ( \24436 , \24435 , \24289 );
and \U$24184 ( \24437 , \24270 , \24279 );
or \U$24185 ( \24438 , \24436 , \24437 );
and \U$24186 ( \24439 , \24434 , \24438 );
and \U$24187 ( \24440 , \24426 , \24433 );
or \U$24188 ( \24441 , \24439 , \24440 );
xor \U$24189 ( \24442 , \24410 , \24441 );
xor \U$24190 ( \24443 , \24301 , \24303 );
and \U$24191 ( \24444 , \24443 , \24310 );
and \U$24192 ( \24445 , \24301 , \24303 );
or \U$24193 ( \24446 , \24444 , \24445 );
xor \U$24194 ( \24447 , \24442 , \24446 );
not \U$24195 ( \24448 , \24447 );
nand \U$24196 ( \24449 , \24338 , \24321 );
buf \U$24197 ( \24450 , \24332 );
and \U$24198 ( \24451 , \24449 , \24450 );
nor \U$24199 ( \24452 , \24338 , \24321 );
nor \U$24200 ( \24453 , \24451 , \24452 );
not \U$24201 ( \24454 , \24453 );
not \U$24202 ( \24455 , \24358 );
not \U$24203 ( \24456 , \24373 );
or \U$24204 ( \24457 , \24455 , \24456 );
nand \U$24205 ( \24458 , \24457 , \24355 );
nand \U$24206 ( \24459 , \24376 , \24361 );
nand \U$24207 ( \24460 , \24458 , \24459 );
not \U$24208 ( \24461 , \24460 );
or \U$24209 ( \24462 , \24454 , \24461 );
not \U$24210 ( \24463 , \24460 );
not \U$24211 ( \24464 , \24453 );
nand \U$24212 ( \24465 , \24463 , \24464 );
nand \U$24213 ( \24466 , \24462 , \24465 );
not \U$24214 ( \24467 , \22280 );
xor \U$24215 ( \24468 , \22269 , \24467 );
xnor \U$24216 ( \24469 , \24468 , \22286 );
not \U$24217 ( \24470 , \24469 );
and \U$24218 ( \24471 , \24466 , \24470 );
not \U$24219 ( \24472 , \24466 );
and \U$24220 ( \24473 , \24472 , \24469 );
nor \U$24221 ( \24474 , \24471 , \24473 );
nand \U$24222 ( \24475 , \24448 , \24474 );
not \U$24223 ( \24476 , \24475 );
not \U$24224 ( \24477 , \24476 );
or \U$24225 ( \24478 , \24386 , \24477 );
not \U$24226 ( \24479 , \24384 );
not \U$24227 ( \24480 , \24475 );
or \U$24228 ( \24481 , \24479 , \24480 );
not \U$24229 ( \24482 , \22536 );
not \U$24230 ( \24483 , \22603 );
or \U$24231 ( \24484 , \24482 , \24483 );
or \U$24232 ( \24485 , \22603 , \22536 );
nand \U$24233 ( \24486 , \24484 , \24485 );
xnor \U$24234 ( \24487 , \24486 , \22571 );
xor \U$24235 ( \24488 , \22387 , \22418 );
xor \U$24236 ( \24489 , \24488 , \22350 );
not \U$24237 ( \24490 , \24489 );
nand \U$24238 ( \24491 , \24487 , \24490 );
not \U$24239 ( \24492 , \24491 );
not \U$24240 ( \24493 , \22304 );
not \U$24241 ( \24494 , \22308 );
or \U$24242 ( \24495 , \24493 , \24494 );
or \U$24243 ( \24496 , \22308 , \22304 );
nand \U$24244 ( \24497 , \24495 , \24496 );
and \U$24245 ( \24498 , \24497 , \22311 );
not \U$24246 ( \24499 , \24497 );
and \U$24247 ( \24500 , \24499 , \22294 );
nor \U$24248 ( \24501 , \24498 , \24500 );
xor \U$24249 ( \24502 , \22501 , \22500 );
xor \U$24250 ( \24503 , \24502 , \22498 );
xor \U$24251 ( \24504 , \22614 , \20637 );
xnor \U$24252 ( \24505 , \24504 , \22620 );
xor \U$24253 ( \24506 , \24505 , \22631 );
xor \U$24254 ( \24507 , \24503 , \24506 );
xor \U$24255 ( \24508 , \24501 , \24507 );
not \U$24256 ( \24509 , \24508 );
or \U$24257 ( \24510 , \24492 , \24509 );
not \U$24258 ( \24511 , \24487 );
nand \U$24259 ( \24512 , \24511 , \24489 );
nand \U$24260 ( \24513 , \24510 , \24512 );
nand \U$24261 ( \24514 , \24481 , \24513 );
nand \U$24262 ( \24515 , \24478 , \24514 );
xor \U$24263 ( \24516 , \20690 , \20612 );
xor \U$24264 ( \24517 , \20514 , \24516 );
not \U$24265 ( \24518 , \22609 );
not \U$24266 ( \24519 , \22666 );
and \U$24267 ( \24520 , \24518 , \24519 );
and \U$24268 ( \24521 , \22666 , \22609 );
nor \U$24269 ( \24522 , \24520 , \24521 );
not \U$24270 ( \24523 , \24522 );
not \U$24271 ( \24524 , \22662 );
and \U$24272 ( \24525 , \24523 , \24524 );
and \U$24273 ( \24526 , \24522 , \22662 );
nor \U$24274 ( \24527 , \24525 , \24526 );
xor \U$24275 ( \24528 , \24517 , \24527 );
not \U$24276 ( \24529 , \22708 );
not \U$24277 ( \24530 , \24529 );
not \U$24278 ( \24531 , \22702 );
not \U$24279 ( \24532 , \22697 );
or \U$24280 ( \24533 , \24531 , \24532 );
or \U$24281 ( \24534 , \22702 , \22697 );
nand \U$24282 ( \24535 , \24533 , \24534 );
not \U$24283 ( \24536 , \24535 );
or \U$24284 ( \24537 , \24530 , \24536 );
or \U$24285 ( \24538 , \24535 , \24529 );
nand \U$24286 ( \24539 , \24537 , \24538 );
xnor \U$24287 ( \24540 , \24528 , \24539 );
xor \U$24288 ( \24541 , \24515 , \24540 );
not \U$24289 ( \24542 , \22606 );
buf \U$24290 ( \24543 , \22422 );
not \U$24291 ( \24544 , \24543 );
not \U$24292 ( \24545 , \22503 );
not \U$24293 ( \24546 , \24545 );
and \U$24294 ( \24547 , \24544 , \24546 );
and \U$24295 ( \24548 , \24543 , \24545 );
nor \U$24296 ( \24549 , \24547 , \24548 );
not \U$24297 ( \24550 , \24549 );
or \U$24298 ( \24551 , \24542 , \24550 );
or \U$24299 ( \24552 , \24549 , \22606 );
nand \U$24300 ( \24553 , \24551 , \24552 );
nor \U$24301 ( \24554 , \24441 , \24410 );
or \U$24302 ( \24555 , \24446 , \24554 );
nand \U$24303 ( \24556 , \24441 , \24410 );
nand \U$24304 ( \24557 , \24555 , \24556 );
not \U$24305 ( \24558 , \24464 );
not \U$24306 ( \24559 , \24470 );
or \U$24307 ( \24560 , \24558 , \24559 );
not \U$24308 ( \24561 , \24469 );
not \U$24309 ( \24562 , \24453 );
or \U$24310 ( \24563 , \24561 , \24562 );
nand \U$24311 ( \24564 , \24563 , \24460 );
nand \U$24312 ( \24565 , \24560 , \24564 );
xor \U$24313 ( \24566 , \24557 , \24565 );
or \U$24314 ( \24567 , \24506 , \24501 );
nand \U$24315 ( \24568 , \24567 , \24503 );
nand \U$24316 ( \24569 , \24501 , \24506 );
nand \U$24317 ( \24570 , \24568 , \24569 );
xor \U$24318 ( \24571 , \24566 , \24570 );
xor \U$24319 ( \24572 , \24553 , \24571 );
not \U$24320 ( \24573 , \22633 );
not \U$24321 ( \24574 , \22291 );
and \U$24322 ( \24575 , \24573 , \24574 );
and \U$24323 ( \24576 , \22633 , \22291 );
nor \U$24324 ( \24577 , \24575 , \24576 );
xor \U$24325 ( \24578 , \24577 , \22313 );
not \U$24326 ( \24579 , \22695 );
not \U$24327 ( \24580 , \24579 );
not \U$24328 ( \24581 , \22688 );
or \U$24329 ( \24582 , \24580 , \24581 );
nand \U$24330 ( \24583 , \22687 , \22695 );
nand \U$24331 ( \24584 , \24582 , \24583 );
and \U$24332 ( \24585 , \24584 , \22684 );
not \U$24333 ( \24586 , \24584 );
and \U$24334 ( \24587 , \24586 , \22683 );
nor \U$24335 ( \24588 , \24585 , \24587 );
xor \U$24336 ( \24589 , \24578 , \24588 );
xor \U$24337 ( \24590 , \22642 , \22653 );
xnor \U$24338 ( \24591 , \24590 , \22657 );
xnor \U$24339 ( \24592 , \24589 , \24591 );
and \U$24340 ( \24593 , \24572 , \24592 );
and \U$24341 ( \24594 , \24553 , \24571 );
or \U$24342 ( \24595 , \24593 , \24594 );
and \U$24343 ( \24596 , \24541 , \24595 );
and \U$24344 ( \24597 , \24515 , \24540 );
or \U$24345 ( \24598 , \24596 , \24597 );
xor \U$24346 ( \24599 , \23803 , \24598 );
xor \U$24347 ( \24600 , \24557 , \24565 );
and \U$24348 ( \24601 , \24600 , \24570 );
and \U$24349 ( \24602 , \24557 , \24565 );
or \U$24350 ( \24603 , \24601 , \24602 );
not \U$24351 ( \24604 , \20981 );
not \U$24352 ( \24605 , \20751 );
and \U$24353 ( \24606 , \24604 , \24605 );
and \U$24354 ( \24607 , \20981 , \20751 );
nor \U$24355 ( \24608 , \24606 , \24607 );
xor \U$24356 ( \24609 , \24608 , \20878 );
nor \U$24357 ( \24610 , \24603 , \24609 );
not \U$24358 ( \24611 , \24588 );
buf \U$24359 ( \24612 , \24578 );
nand \U$24360 ( \24613 , \24611 , \24612 );
and \U$24361 ( \24614 , \24613 , \24591 );
nor \U$24362 ( \24615 , \24611 , \24612 );
nor \U$24363 ( \24616 , \24614 , \24615 );
or \U$24364 ( \24617 , \24610 , \24616 );
nand \U$24365 ( \24618 , \24603 , \24609 );
nand \U$24366 ( \24619 , \24617 , \24618 );
not \U$24367 ( \24620 , \24517 );
nand \U$24368 ( \24621 , \24620 , \24527 );
not \U$24369 ( \24622 , \24621 );
not \U$24370 ( \24623 , \24539 );
or \U$24371 ( \24624 , \24622 , \24623 );
not \U$24372 ( \24625 , \24527 );
nand \U$24373 ( \24626 , \24625 , \24517 );
nand \U$24374 ( \24627 , \24624 , \24626 );
xor \U$24375 ( \24628 , \24619 , \24627 );
xor \U$24376 ( \24629 , \22723 , \22720 );
xnor \U$24377 ( \24630 , \24629 , \22717 );
xor \U$24378 ( \24631 , \24628 , \24630 );
and \U$24379 ( \24632 , \24599 , \24631 );
and \U$24380 ( \24633 , \23803 , \24598 );
or \U$24381 ( \24634 , \24632 , \24633 );
xor \U$24382 ( \24635 , \22266 , \22732 );
xnor \U$24383 ( \24636 , \24635 , \22729 );
not \U$24384 ( \24637 , \24636 );
xor \U$24385 ( \24638 , \24619 , \24627 );
and \U$24386 ( \24639 , \24638 , \24630 );
and \U$24387 ( \24640 , \24619 , \24627 );
or \U$24388 ( \24641 , \24639 , \24640 );
not \U$24389 ( \24642 , \24641 );
and \U$24390 ( \24643 , \22124 , \22069 );
not \U$24391 ( \24644 , \22124 );
and \U$24392 ( \24645 , \24644 , \22068 );
nor \U$24393 ( \24646 , \24643 , \24645 );
not \U$24394 ( \24647 , \24646 );
or \U$24395 ( \24648 , \24642 , \24647 );
not \U$24396 ( \24649 , \24641 );
not \U$24397 ( \24650 , \24646 );
nand \U$24398 ( \24651 , \24649 , \24650 );
nand \U$24399 ( \24652 , \24648 , \24651 );
not \U$24400 ( \24653 , \24652 );
or \U$24401 ( \24654 , \24637 , \24653 );
or \U$24402 ( \24655 , \24652 , \24636 );
nand \U$24403 ( \24656 , \24654 , \24655 );
xor \U$24404 ( \24657 , \24634 , \24656 );
and \U$24405 ( \24658 , \23797 , \24657 );
not \U$24406 ( \24659 , \24636 );
not \U$24407 ( \24660 , \24646 );
or \U$24408 ( \24661 , \24659 , \24660 );
nand \U$24409 ( \24662 , \24661 , \24641 );
not \U$24410 ( \24663 , \24636 );
nand \U$24411 ( \24664 , \24663 , \24650 );
and \U$24412 ( \24665 , \24662 , \24664 );
not \U$24413 ( \24666 , \24665 );
not \U$24414 ( \24667 , \23227 );
not \U$24415 ( \24668 , \22734 );
nand \U$24416 ( \24669 , \22068 , \22124 );
not \U$24417 ( \24670 , \24669 );
or \U$24418 ( \24671 , \24668 , \24670 );
or \U$24419 ( \24672 , \24669 , \22734 );
nand \U$24420 ( \24673 , \24671 , \24672 );
not \U$24421 ( \24674 , \24673 );
or \U$24422 ( \24675 , \24667 , \24674 );
not \U$24423 ( \24676 , \24673 );
nand \U$24424 ( \24677 , \24676 , \23228 );
nand \U$24425 ( \24678 , \24675 , \24677 );
not \U$24426 ( \24679 , \24678 );
or \U$24427 ( \24680 , \24666 , \24679 );
or \U$24428 ( \24681 , \24678 , \24665 );
nand \U$24429 ( \24682 , \24680 , \24681 );
xor \U$24430 ( \24683 , \23803 , \24598 );
xor \U$24431 ( \24684 , \24683 , \24631 );
xor \U$24432 ( \24685 , \24086 , \24194 );
xor \U$24433 ( \24686 , \24685 , \24293 );
not \U$24434 ( \24687 , \24686 );
not \U$24435 ( \24688 , \24078 );
xor \U$24436 ( \24689 , \24012 , \23913 );
not \U$24437 ( \24690 , \24689 );
or \U$24438 ( \24691 , \24688 , \24690 );
or \U$24439 ( \24692 , \24689 , \24078 );
nand \U$24440 ( \24693 , \24691 , \24692 );
nand \U$24441 ( \24694 , \24687 , \24693 );
not \U$24442 ( \24695 , \24694 );
not \U$24443 ( \24696 , \24695 );
not \U$24444 ( \24697 , \2385 );
not \U$24445 ( \24698 , RIbe2b018_114);
not \U$24446 ( \24699 , \24698 );
and \U$24447 ( \24700 , \24697 , \24699 );
and \U$24448 ( \24701 , \8833 , RIbe2b630_127);
nor \U$24449 ( \24702 , \24700 , \24701 );
and \U$24450 ( \24703 , \24702 , \1076 );
not \U$24451 ( \24704 , \24702 );
and \U$24452 ( \24705 , \24704 , \9083 );
nor \U$24453 ( \24706 , \24703 , \24705 );
not \U$24454 ( \24707 , \24706 );
not \U$24455 ( \24708 , \24707 );
not \U$24456 ( \24709 , RIbe2b108_116);
not \U$24457 ( \24710 , \6414 );
or \U$24458 ( \24711 , \24709 , \24710 );
nand \U$24459 ( \24712 , \4600 , RIbe2b090_115);
nand \U$24460 ( \24713 , \24711 , \24712 );
and \U$24461 ( \24714 , \24713 , \4603 );
not \U$24462 ( \24715 , \24713 );
and \U$24463 ( \24716 , \24715 , \4323 );
nor \U$24464 ( \24717 , \24714 , \24716 );
not \U$24465 ( \24718 , RIbe2b180_117);
not \U$24466 ( \24719 , \7880 );
or \U$24467 ( \24720 , \24718 , \24719 );
nand \U$24468 ( \24721 , \6787 , RIbe2b270_119);
nand \U$24469 ( \24722 , \24720 , \24721 );
and \U$24470 ( \24723 , \24722 , \3448 );
not \U$24471 ( \24724 , \24722 );
and \U$24472 ( \24725 , \24724 , \3471 );
nor \U$24473 ( \24726 , \24723 , \24725 );
not \U$24474 ( \24727 , RIbe2af28_112);
not \U$24475 ( \24728 , \6797 );
or \U$24476 ( \24729 , \24727 , \24728 );
nand \U$24477 ( \24730 , RIbe2b1f8_118, \6800 );
nand \U$24478 ( \24731 , \24729 , \24730 );
and \U$24479 ( \24732 , \24731 , \4346 );
not \U$24480 ( \24733 , \24731 );
and \U$24481 ( \24734 , \24733 , \2887 );
nor \U$24482 ( \24735 , \24732 , \24734 );
not \U$24483 ( \24736 , \24735 );
nand \U$24484 ( \24737 , \24726 , \24736 );
and \U$24485 ( \24738 , \24717 , \24737 );
nor \U$24486 ( \24739 , \24726 , \24736 );
nor \U$24487 ( \24740 , \24738 , \24739 );
not \U$24488 ( \24741 , \24740 );
or \U$24489 ( \24742 , \24708 , \24741 );
nand \U$24490 ( \24743 , \5467 , RIbe2ab68_104);
and \U$24491 ( \24744 , \24743 , \2563 );
not \U$24492 ( \24745 , \24743 );
and \U$24493 ( \24746 , \24745 , \1131 );
nor \U$24494 ( \24747 , \24744 , \24746 );
not \U$24495 ( \24748 , \24747 );
not \U$24496 ( \24749 , RIbe2b018_114);
not \U$24497 ( \24750 , \10010 );
or \U$24498 ( \24751 , \24749 , \24750 );
nand \U$24499 ( \24752 , RIbe2afa0_113, \2901 );
nand \U$24500 ( \24753 , \24751 , \24752 );
xor \U$24501 ( \24754 , \24753 , \2379 );
nand \U$24502 ( \24755 , \24748 , \24754 );
not \U$24503 ( \24756 , \24755 );
not \U$24504 ( \24757 , \2889 );
not \U$24505 ( \24758 , \17802 );
and \U$24506 ( \24759 , \24757 , \24758 );
and \U$24507 ( \24760 , \2583 , RIbe2aaf0_103);
nor \U$24508 ( \24761 , \24759 , \24760 );
and \U$24509 ( \24762 , \24761 , \1076 );
not \U$24510 ( \24763 , \24761 );
and \U$24511 ( \24764 , \24763 , \1277 );
nor \U$24512 ( \24765 , \24762 , \24764 );
not \U$24513 ( \24766 , \24765 );
or \U$24514 ( \24767 , \24756 , \24766 );
not \U$24515 ( \24768 , \24754 );
nand \U$24516 ( \24769 , \24768 , \24747 );
nand \U$24517 ( \24770 , \24767 , \24769 );
nand \U$24518 ( \24771 , \24742 , \24770 );
not \U$24519 ( \24772 , \24740 );
nand \U$24520 ( \24773 , \24772 , \24706 );
and \U$24521 ( \24774 , \24771 , \24773 );
not \U$24522 ( \24775 , \24774 );
not \U$24523 ( \24776 , RIbe2a280_85);
not \U$24524 ( \24777 , \20809 );
or \U$24525 ( \24778 , \24776 , \24777 );
nand \U$24526 ( \24779 , \7056 , RIbe2a208_84);
nand \U$24527 ( \24780 , \24778 , \24779 );
and \U$24528 ( \24781 , \24780 , \4592 );
not \U$24529 ( \24782 , \24780 );
and \U$24530 ( \24783 , \24782 , \4586 );
nor \U$24531 ( \24784 , \24781 , \24783 );
not \U$24532 ( \24785 , RIbe2a190_83);
not \U$24533 ( \24786 , \20796 );
or \U$24534 ( \24787 , \24785 , \24786 );
nand \U$24535 ( \24788 , \5749 , RIbe2a5c8_92);
nand \U$24536 ( \24789 , \24787 , \24788 );
and \U$24537 ( \24790 , \24789 , \10984 );
not \U$24538 ( \24791 , \24789 );
and \U$24539 ( \24792 , \24791 , \8253 );
nor \U$24540 ( \24793 , \24790 , \24792 );
nand \U$24541 ( \24794 , \24784 , \24793 );
not \U$24542 ( \24795 , RIbe2a550_91);
not \U$24543 ( \24796 , \21081 );
or \U$24544 ( \24797 , \24795 , \24796 );
nand \U$24545 ( \24798 , \21084 , RIbe2a988_100);
nand \U$24546 ( \24799 , \24797 , \24798 );
xnor \U$24547 ( \24800 , \24799 , \21090 );
and \U$24548 ( \24801 , \24794 , \24800 );
nor \U$24549 ( \24802 , \24793 , \24784 );
nor \U$24550 ( \24803 , \24801 , \24802 );
not \U$24551 ( \24804 , \24803 );
not \U$24552 ( \24805 , RIbe29e48_76);
not \U$24553 ( \24806 , \7974 );
or \U$24554 ( \24807 , \24805 , \24806 );
nand \U$24555 ( \24808 , \7981 , RIbe29dd0_75);
nand \U$24556 ( \24809 , \24807 , \24808 );
xnor \U$24557 ( \24810 , \24809 , \7984 );
and \U$24558 ( \24811 , \20405 , RIbe29c68_72);
and \U$24559 ( \24812 , \10919 , RIbe29bf0_71);
nor \U$24560 ( \24813 , \24811 , \24812 );
and \U$24561 ( \24814 , \24813 , \8077 );
not \U$24562 ( \24815 , \24813 );
and \U$24563 ( \24816 , \24815 , \7970 );
nor \U$24564 ( \24817 , \24814 , \24816 );
or \U$24565 ( \24818 , \24810 , \24817 );
and \U$24566 ( \24819 , \7299 , RIbe2a028_80);
not \U$24567 ( \24820 , RIbe29fb0_79);
nor \U$24568 ( \24821 , \24820 , \10897 );
nor \U$24569 ( \24822 , \24819 , \24821 );
and \U$24570 ( \24823 , \24822 , \14650 );
not \U$24571 ( \24824 , \24822 );
and \U$24572 ( \24825 , \24824 , \7660 );
nor \U$24573 ( \24826 , \24823 , \24825 );
and \U$24574 ( \24827 , \24818 , \24826 );
and \U$24575 ( \24828 , \24810 , \24817 );
nor \U$24576 ( \24829 , \24827 , \24828 );
not \U$24577 ( \24830 , \24829 );
or \U$24578 ( \24831 , \24804 , \24830 );
not \U$24579 ( \24832 , RIbe2a2f8_86);
not \U$24580 ( \24833 , \21608 );
or \U$24581 ( \24834 , \24832 , \24833 );
nand \U$24582 ( \24835 , RIbe2acd0_107, \6962 );
nand \U$24583 ( \24836 , \24834 , \24835 );
and \U$24584 ( \24837 , \24836 , \7293 );
not \U$24585 ( \24838 , \24836 );
and \U$24586 ( \24839 , \24838 , \6572 );
nor \U$24587 ( \24840 , \24837 , \24839 );
not \U$24588 ( \24841 , \24840 );
not \U$24589 ( \24842 , RIbe2a3e8_88);
not \U$24590 ( \24843 , \20487 );
or \U$24591 ( \24844 , \24842 , \24843 );
nand \U$24592 ( \24845 , RIbe2a370_87, \6595 );
nand \U$24593 ( \24846 , \24844 , \24845 );
and \U$24594 ( \24847 , \24846 , \6873 );
not \U$24595 ( \24848 , \24846 );
and \U$24596 ( \24849 , \24848 , \6601 );
nor \U$24597 ( \24850 , \24847 , \24849 );
not \U$24598 ( \24851 , \24850 );
not \U$24599 ( \24852 , \24851 );
or \U$24600 ( \24853 , \24841 , \24852 );
not \U$24601 ( \24854 , \24840 );
not \U$24602 ( \24855 , \24854 );
not \U$24603 ( \24856 , \24850 );
or \U$24604 ( \24857 , \24855 , \24856 );
not \U$24605 ( \24858 , RIbe2a910_99);
not \U$24606 ( \24859 , \6880 );
or \U$24607 ( \24860 , \24858 , \24859 );
nand \U$24608 ( \24861 , \7076 , RIbe2b5b8_126);
nand \U$24609 ( \24862 , \24860 , \24861 );
and \U$24610 ( \24863 , \24862 , \6546 );
not \U$24611 ( \24864 , \24862 );
and \U$24612 ( \24865 , \24864 , \9933 );
nor \U$24613 ( \24866 , \24863 , \24865 );
nand \U$24614 ( \24867 , \24857 , \24866 );
nand \U$24615 ( \24868 , \24853 , \24867 );
nand \U$24616 ( \24869 , \24831 , \24868 );
not \U$24617 ( \24870 , \24829 );
not \U$24618 ( \24871 , \24803 );
nand \U$24619 ( \24872 , \24870 , \24871 );
nand \U$24620 ( \24873 , \24869 , \24872 );
not \U$24621 ( \24874 , \24873 );
not \U$24622 ( \24875 , \24874 );
or \U$24623 ( \24876 , \24775 , \24875 );
not \U$24624 ( \24877 , RIbe28b88_36);
not \U$24625 ( \24878 , \15249 );
or \U$24626 ( \24879 , \24877 , \24878 );
nand \U$24627 ( \24880 , \12794 , RIbe29290_51);
nand \U$24628 ( \24881 , \24879 , \24880 );
and \U$24629 ( \24882 , \24881 , \14336 );
not \U$24630 ( \24883 , \24881 );
and \U$24631 ( \24884 , \24883 , \14335 );
nor \U$24632 ( \24885 , \24882 , \24884 );
not \U$24633 ( \24886 , \24885 );
not \U$24634 ( \24887 , RIbe28a20_33);
not \U$24635 ( \24888 , \13002 );
or \U$24636 ( \24889 , \24887 , \24888 );
nand \U$24637 ( \24890 , RIbe289a8_32, RIbe2ae38_110);
nand \U$24638 ( \24891 , \24889 , \24890 );
xor \U$24639 ( \24892 , \24891 , RIbe2aeb0_111);
not \U$24640 ( \24893 , \24892 );
nand \U$24641 ( \24894 , \24893 , \2563 );
not \U$24642 ( \24895 , \24894 );
or \U$24643 ( \24896 , \24886 , \24895 );
nand \U$24644 ( \24897 , \24892 , \1132 );
nand \U$24645 ( \24898 , \24896 , \24897 );
not \U$24646 ( \24899 , \24898 );
and \U$24647 ( \24900 , \14725 , RIbe27e68_8);
and \U$24648 ( \24901 , \13086 , RIbe28660_25);
nor \U$24649 ( \24902 , \24900 , \24901 );
and \U$24650 ( \24903 , \24902 , \12770 );
not \U$24651 ( \24904 , \24902 );
and \U$24652 ( \24905 , \24904 , \12927 );
nor \U$24653 ( \24906 , \24903 , \24905 );
not \U$24654 ( \24907 , \24906 );
not \U$24655 ( \24908 , RIbe28f48_44);
not \U$24656 ( \24909 , \10936 );
or \U$24657 ( \24910 , \24908 , \24909 );
nand \U$24658 ( \24911 , \12971 , RIbe28ed0_43);
nand \U$24659 ( \24912 , \24910 , \24911 );
and \U$24660 ( \24913 , \24912 , \9902 );
not \U$24661 ( \24914 , \24912 );
and \U$24662 ( \24915 , \24914 , \12218 );
nor \U$24663 ( \24916 , \24913 , \24915 );
not \U$24664 ( \24917 , \24916 );
or \U$24665 ( \24918 , \24907 , \24917 );
or \U$24666 ( \24919 , \24916 , \24906 );
and \U$24667 ( \24920 , \15205 , RIbe27fd0_11);
and \U$24668 ( \24921 , \12947 , RIbe27f58_10);
nor \U$24669 ( \24922 , \24920 , \24921 );
not \U$24670 ( \24923 , \24922 );
not \U$24671 ( \24924 , \12195 );
and \U$24672 ( \24925 , \24923 , \24924 );
and \U$24673 ( \24926 , \24922 , \12195 );
nor \U$24674 ( \24927 , \24925 , \24926 );
not \U$24675 ( \24928 , \24927 );
nand \U$24676 ( \24929 , \24919 , \24928 );
nand \U$24677 ( \24930 , \24918 , \24929 );
not \U$24678 ( \24931 , \24930 );
or \U$24679 ( \24932 , \24899 , \24931 );
not \U$24680 ( \24933 , \24898 );
not \U$24681 ( \24934 , \24930 );
nand \U$24682 ( \24935 , \24933 , \24934 );
not \U$24683 ( \24936 , RIbe285e8_24);
not \U$24684 ( \24937 , \19262 );
or \U$24685 ( \24938 , \24936 , \24937 );
nand \U$24686 ( \24939 , \12711 , RIbe287c8_28);
nand \U$24687 ( \24940 , \24938 , \24939 );
and \U$24688 ( \24941 , \24940 , \13068 );
not \U$24689 ( \24942 , \24940 );
and \U$24690 ( \24943 , \24942 , \12723 );
nor \U$24691 ( \24944 , \24941 , \24943 );
not \U$24692 ( \24945 , RIbe28480_21);
not \U$24693 ( \24946 , \15161 );
or \U$24694 ( \24947 , \24945 , \24946 );
nand \U$24695 ( \24948 , \12735 , RIbe28408_20);
nand \U$24696 ( \24949 , \24947 , \24948 );
and \U$24697 ( \24950 , \24949 , \12746 );
not \U$24698 ( \24951 , \24949 );
and \U$24699 ( \24952 , \24951 , \14358 );
nor \U$24700 ( \24953 , \24950 , \24952 );
not \U$24701 ( \24954 , \24953 );
or \U$24702 ( \24955 , \24944 , \24954 );
not \U$24703 ( \24956 , RIbe28390_19);
not \U$24704 ( \24957 , \14550 );
or \U$24705 ( \24958 , \24956 , \24957 );
nand \U$24706 ( \24959 , \13012 , RIbe28b10_35);
nand \U$24707 ( \24960 , \24958 , \24959 );
and \U$24708 ( \24961 , \24960 , \13595 );
not \U$24709 ( \24962 , \24960 );
and \U$24710 ( \24963 , \24962 , \12863 );
nor \U$24711 ( \24964 , \24961 , \24963 );
nand \U$24712 ( \24965 , \24955 , \24964 );
nand \U$24713 ( \24966 , \24944 , \24954 );
nand \U$24714 ( \24967 , \24965 , \24966 );
nand \U$24715 ( \24968 , \24935 , \24967 );
nand \U$24716 ( \24969 , \24932 , \24968 );
nand \U$24717 ( \24970 , \24876 , \24969 );
not \U$24718 ( \24971 , \24774 );
nand \U$24719 ( \24972 , \24971 , \24873 );
nand \U$24720 ( \24973 , \24970 , \24972 );
and \U$24721 ( \24974 , \24422 , \1082 );
not \U$24722 ( \24975 , \24422 );
and \U$24723 ( \24976 , \24975 , \1309 );
or \U$24724 ( \24977 , \24974 , \24976 );
xnor \U$24725 ( \24978 , \24977 , \24416 );
not \U$24726 ( \24979 , \24978 );
and \U$24727 ( \24980 , \1286 , RIbe2ab68_104);
and \U$24728 ( \24981 , \1117 , RIbe2aaf0_103);
nor \U$24729 ( \24982 , \24980 , \24981 );
and \U$24730 ( \24983 , \24982 , \1131 );
not \U$24731 ( \24984 , \24982 );
and \U$24732 ( \24985 , \24984 , \1448 );
nor \U$24733 ( \24986 , \24983 , \24985 );
not \U$24734 ( \24987 , \24986 );
xor \U$24735 ( \24988 , \24038 , \24048 );
and \U$24736 ( \24989 , \24988 , \24029 );
not \U$24737 ( \24990 , \24988 );
not \U$24738 ( \24991 , \24029 );
and \U$24739 ( \24992 , \24990 , \24991 );
nor \U$24740 ( \24993 , \24989 , \24992 );
not \U$24741 ( \24994 , \24993 );
or \U$24742 ( \24995 , \24987 , \24994 );
not \U$24743 ( \24996 , \23874 );
not \U$24744 ( \24997 , \23851 );
or \U$24745 ( \24998 , \24996 , \24997 );
or \U$24746 ( \24999 , \23851 , \23874 );
nand \U$24747 ( \25000 , \24998 , \24999 );
and \U$24748 ( \25001 , \25000 , \23862 );
not \U$24749 ( \25002 , \25000 );
and \U$24750 ( \25003 , \25002 , \23861 );
nor \U$24751 ( \25004 , \25001 , \25003 );
nand \U$24752 ( \25005 , \24995 , \25004 );
not \U$24753 ( \25006 , \24986 );
not \U$24754 ( \25007 , \24993 );
nand \U$24755 ( \25008 , \25006 , \25007 );
nand \U$24756 ( \25009 , \24979 , \25005 , \25008 );
not \U$24757 ( \25010 , \25009 );
xor \U$24758 ( \25011 , \23987 , \23996 );
xor \U$24759 ( \25012 , \25011 , \24004 );
not \U$24760 ( \25013 , \23812 );
not \U$24761 ( \25014 , \23839 );
not \U$24762 ( \25015 , \23823 );
or \U$24763 ( \25016 , \25014 , \25015 );
or \U$24764 ( \25017 , \23823 , \23839 );
nand \U$24765 ( \25018 , \25016 , \25017 );
not \U$24766 ( \25019 , \25018 );
or \U$24767 ( \25020 , \25013 , \25019 );
or \U$24768 ( \25021 , \25018 , \23812 );
nand \U$24769 ( \25022 , \25020 , \25021 );
xor \U$24770 ( \25023 , \25012 , \25022 );
xor \U$24771 ( \25024 , \23894 , \7984 );
xor \U$24772 ( \25025 , \25024 , \23908 );
xnor \U$24773 ( \25026 , \25025 , \23888 );
and \U$24774 ( \25027 , \25023 , \25026 );
and \U$24775 ( \25028 , \25012 , \25022 );
or \U$24776 ( \25029 , \25027 , \25028 );
not \U$24777 ( \25030 , \25029 );
or \U$24778 ( \25031 , \25010 , \25030 );
nand \U$24779 ( \25032 , \25005 , \25008 );
nand \U$24780 ( \25033 , \25032 , \24978 );
nand \U$24781 ( \25034 , \25031 , \25033 );
xor \U$24782 ( \25035 , \24973 , \25034 );
xor \U$24783 ( \25036 , \24019 , \24051 );
xor \U$24784 ( \25037 , \25036 , \24075 );
not \U$24785 ( \25038 , \25037 );
xor \U$24786 ( \25039 , \24119 , \24157 );
xor \U$24787 ( \25040 , \25039 , \24190 );
not \U$24788 ( \25041 , \25040 );
not \U$24789 ( \25042 , \25041 );
or \U$24790 ( \25043 , \25038 , \25042 );
xor \U$24791 ( \25044 , \24224 , \24290 );
xor \U$24792 ( \25045 , \25044 , \24259 );
nand \U$24793 ( \25046 , \25043 , \25045 );
not \U$24794 ( \25047 , \25037 );
nand \U$24795 ( \25048 , \25040 , \25047 );
nand \U$24796 ( \25049 , \25046 , \25048 );
and \U$24797 ( \25050 , \25035 , \25049 );
and \U$24798 ( \25051 , \24973 , \25034 );
or \U$24799 ( \25052 , \25050 , \25051 );
not \U$24800 ( \25053 , \25052 );
or \U$24801 ( \25054 , \24696 , \25053 );
not \U$24802 ( \25055 , \24694 );
not \U$24803 ( \25056 , \25052 );
not \U$24804 ( \25057 , \25056 );
or \U$24805 ( \25058 , \25055 , \25057 );
xor \U$24806 ( \25059 , \24426 , \24433 );
xor \U$24807 ( \25060 , \25059 , \24438 );
not \U$24808 ( \25061 , \25060 );
not \U$24809 ( \25062 , \24405 );
not \U$24810 ( \25063 , \24390 );
and \U$24811 ( \25064 , \25062 , \25063 );
and \U$24812 ( \25065 , \24405 , \24390 );
nor \U$24813 ( \25066 , \25064 , \25065 );
and \U$24814 ( \25067 , \25066 , \24408 );
not \U$24815 ( \25068 , \25066 );
and \U$24816 ( \25069 , \25068 , \24395 );
nor \U$24817 ( \25070 , \25067 , \25069 );
nand \U$24818 ( \25071 , \25061 , \25070 );
not \U$24819 ( \25072 , \25071 );
not \U$24820 ( \25073 , \24343 );
not \U$24821 ( \25074 , \24378 );
or \U$24822 ( \25075 , \25073 , \25074 );
or \U$24823 ( \25076 , \24378 , \24343 );
nand \U$24824 ( \25077 , \25075 , \25076 );
not \U$24825 ( \25078 , \24311 );
and \U$24826 ( \25079 , \25077 , \25078 );
not \U$24827 ( \25080 , \25077 );
and \U$24828 ( \25081 , \25080 , \24311 );
nor \U$24829 ( \25082 , \25079 , \25081 );
not \U$24830 ( \25083 , \25082 );
or \U$24831 ( \25084 , \25072 , \25083 );
not \U$24832 ( \25085 , \25070 );
nand \U$24833 ( \25086 , \25085 , \25060 );
nand \U$24834 ( \25087 , \25084 , \25086 );
nand \U$24835 ( \25088 , \25058 , \25087 );
nand \U$24836 ( \25089 , \25054 , \25088 );
not \U$24837 ( \25090 , \24490 );
not \U$24838 ( \25091 , \24511 );
or \U$24839 ( \25092 , \25090 , \25091 );
nand \U$24840 ( \25093 , \24487 , \24489 );
nand \U$24841 ( \25094 , \25092 , \25093 );
xor \U$24842 ( \25095 , \24501 , \25094 );
xnor \U$24843 ( \25096 , \25095 , \24507 );
not \U$24844 ( \25097 , \25096 );
not \U$24845 ( \25098 , \25097 );
not \U$24846 ( \25099 , \24447 );
not \U$24847 ( \25100 , \24474 );
or \U$24848 ( \25101 , \25099 , \25100 );
or \U$24849 ( \25102 , \24474 , \24447 );
nand \U$24850 ( \25103 , \25101 , \25102 );
not \U$24851 ( \25104 , \25103 );
or \U$24852 ( \25105 , \25098 , \25104 );
not \U$24853 ( \25106 , \25103 );
not \U$24854 ( \25107 , \25106 );
not \U$24855 ( \25108 , \25096 );
or \U$24856 ( \25109 , \25107 , \25108 );
xor \U$24857 ( \25110 , \24081 , \24296 );
xor \U$24858 ( \25111 , \25110 , \24381 );
not \U$24859 ( \25112 , \25111 );
nand \U$24860 ( \25113 , \25109 , \25112 );
nand \U$24861 ( \25114 , \25105 , \25113 );
xor \U$24862 ( \25115 , \25089 , \25114 );
xor \U$24863 ( \25116 , \24553 , \24571 );
xor \U$24864 ( \25117 , \25116 , \24592 );
and \U$24865 ( \25118 , \25115 , \25117 );
and \U$24866 ( \25119 , \25089 , \25114 );
or \U$24867 ( \25120 , \25118 , \25119 );
not \U$24868 ( \25121 , \25120 );
not \U$24869 ( \25122 , \24609 );
buf \U$24870 ( \25123 , \24603 );
xor \U$24871 ( \25124 , \25122 , \25123 );
xnor \U$24872 ( \25125 , \25124 , \24616 );
nand \U$24873 ( \25126 , \25121 , \25125 );
not \U$24874 ( \25127 , \25126 );
xor \U$24875 ( \25128 , \24515 , \24540 );
xor \U$24876 ( \25129 , \25128 , \24595 );
not \U$24877 ( \25130 , \25129 );
or \U$24878 ( \25131 , \25127 , \25130 );
not \U$24879 ( \25132 , \25125 );
nand \U$24880 ( \25133 , \25132 , \25120 );
nand \U$24881 ( \25134 , \25131 , \25133 );
nand \U$24882 ( \25135 , \24684 , \25134 );
not \U$24883 ( \25136 , \24684 );
not \U$24884 ( \25137 , \25134 );
nand \U$24885 ( \25138 , \25136 , \25137 );
and \U$24886 ( \25139 , \24682 , \25135 , \25138 );
not \U$24887 ( \25140 , \24513 );
not \U$24888 ( \25141 , \25140 );
not \U$24889 ( \25142 , \24384 );
not \U$24890 ( \25143 , \24476 );
or \U$24891 ( \25144 , \25142 , \25143 );
nand \U$24892 ( \25145 , \24475 , \24385 );
nand \U$24893 ( \25146 , \25144 , \25145 );
not \U$24894 ( \25147 , \25146 );
or \U$24895 ( \25148 , \25141 , \25147 );
or \U$24896 ( \25149 , \25146 , \25140 );
nand \U$24897 ( \25150 , \25148 , \25149 );
xnor \U$24898 ( \25151 , \23923 , \23929 );
not \U$24899 ( \25152 , \25151 );
not \U$24900 ( \25153 , \23940 );
and \U$24901 ( \25154 , \25152 , \25153 );
and \U$24902 ( \25155 , \25151 , \23940 );
nor \U$24903 ( \25156 , \25154 , \25155 );
not \U$24904 ( \25157 , \25156 );
xor \U$24905 ( \25158 , \23862 , \24986 );
xnor \U$24906 ( \25159 , \25158 , \25000 );
and \U$24907 ( \25160 , \25159 , \24993 );
not \U$24908 ( \25161 , \25159 );
and \U$24909 ( \25162 , \25161 , \25007 );
nor \U$24910 ( \25163 , \25160 , \25162 );
not \U$24911 ( \25164 , \25163 );
or \U$24912 ( \25165 , \25157 , \25164 );
xor \U$24913 ( \25166 , \25012 , \25022 );
xor \U$24914 ( \25167 , \25166 , \25026 );
nand \U$24915 ( \25168 , \25165 , \25167 );
not \U$24916 ( \25169 , \25156 );
not \U$24917 ( \25170 , \25163 );
nand \U$24918 ( \25171 , \25169 , \25170 );
nand \U$24919 ( \25172 , \25168 , \25171 );
not \U$24920 ( \25173 , \24854 );
not \U$24921 ( \25174 , \24851 );
or \U$24922 ( \25175 , \25173 , \25174 );
nand \U$24923 ( \25176 , \24850 , \24840 );
nand \U$24924 ( \25177 , \25175 , \25176 );
xor \U$24925 ( \25178 , \25177 , \24866 );
not \U$24926 ( \25179 , \25178 );
xor \U$24927 ( \25180 , \24784 , \24800 );
xor \U$24928 ( \25181 , \25180 , \24793 );
not \U$24929 ( \25182 , \25181 );
or \U$24930 ( \25183 , \25179 , \25182 );
or \U$24931 ( \25184 , \25178 , \25181 );
xor \U$24932 ( \25185 , \24810 , \24817 );
xor \U$24933 ( \25186 , \25185 , \24826 );
nand \U$24934 ( \25187 , \25184 , \25186 );
nand \U$24935 ( \25188 , \25183 , \25187 );
not \U$24936 ( \25189 , \23973 );
xnor \U$24937 ( \25190 , \23953 , \23962 );
not \U$24938 ( \25191 , \25190 );
or \U$24939 ( \25192 , \25189 , \25191 );
or \U$24940 ( \25193 , \25190 , \23973 );
nand \U$24941 ( \25194 , \25192 , \25193 );
nor \U$24942 ( \25195 , \25188 , \25194 );
not \U$24943 ( \25196 , \24964 );
not \U$24944 ( \25197 , \25196 );
not \U$24945 ( \25198 , \24954 );
or \U$24946 ( \25199 , \25197 , \25198 );
nand \U$24947 ( \25200 , \24953 , \24964 );
nand \U$24948 ( \25201 , \25199 , \25200 );
buf \U$24949 ( \25202 , \24944 );
not \U$24950 ( \25203 , \25202 );
and \U$24951 ( \25204 , \25201 , \25203 );
not \U$24952 ( \25205 , \25201 );
and \U$24953 ( \25206 , \25205 , \25202 );
nor \U$24954 ( \25207 , \25204 , \25206 );
and \U$24955 ( \25208 , \24892 , \2563 );
not \U$24956 ( \25209 , \24892 );
and \U$24957 ( \25210 , \25209 , \1131 );
nor \U$24958 ( \25211 , \25208 , \25210 );
not \U$24959 ( \25212 , \25211 );
not \U$24960 ( \25213 , \24885 );
or \U$24961 ( \25214 , \25212 , \25213 );
or \U$24962 ( \25215 , \24885 , \25211 );
nand \U$24963 ( \25216 , \25214 , \25215 );
not \U$24964 ( \25217 , \25216 );
and \U$24965 ( \25218 , \25207 , \25217 );
and \U$24966 ( \25219 , \24906 , \24927 );
not \U$24967 ( \25220 , \24906 );
and \U$24968 ( \25221 , \25220 , \24928 );
or \U$24969 ( \25222 , \25219 , \25221 );
buf \U$24970 ( \25223 , \24916 );
not \U$24971 ( \25224 , \25223 );
and \U$24972 ( \25225 , \25222 , \25224 );
not \U$24973 ( \25226 , \25222 );
and \U$24974 ( \25227 , \25226 , \25223 );
nor \U$24975 ( \25228 , \25225 , \25227 );
nor \U$24976 ( \25229 , \25218 , \25228 );
nor \U$24977 ( \25230 , \25207 , \25217 );
nor \U$24978 ( \25231 , \25229 , \25230 );
or \U$24979 ( \25232 , \25195 , \25231 );
nand \U$24980 ( \25233 , \25188 , \25194 );
nand \U$24981 ( \25234 , \25232 , \25233 );
not \U$24982 ( \25235 , \25234 );
not \U$24983 ( \25236 , RIbe2b270_119);
not \U$24984 ( \25237 , \4804 );
or \U$24985 ( \25238 , \25236 , \25237 );
nand \U$24986 ( \25239 , \7858 , RIbe2b108_116);
nand \U$24987 ( \25240 , \25238 , \25239 );
not \U$24988 ( \25241 , \25240 );
not \U$24989 ( \25242 , \7865 );
and \U$24990 ( \25243 , \25241 , \25242 );
and \U$24991 ( \25244 , \25240 , \4323 );
nor \U$24992 ( \25245 , \25243 , \25244 );
not \U$24993 ( \25246 , RIbe2b090_115);
not \U$24994 ( \25247 , \21097 );
or \U$24995 ( \25248 , \25246 , \25247 );
nand \U$24996 ( \25249 , \22378 , RIbe2a280_85);
nand \U$24997 ( \25250 , \25248 , \25249 );
xor \U$24998 ( \25251 , \25250 , \4592 );
nand \U$24999 ( \25252 , \25245 , \25251 );
not \U$25000 ( \25253 , RIbe2a208_84);
not \U$25001 ( \25254 , \6630 );
or \U$25002 ( \25255 , \25253 , \25254 );
nand \U$25003 ( \25256 , \10269 , RIbe2a190_83);
nand \U$25004 ( \25257 , \25255 , \25256 );
not \U$25005 ( \25258 , \8253 );
not \U$25006 ( \25259 , \25258 );
and \U$25007 ( \25260 , \25257 , \25259 );
not \U$25008 ( \25261 , \25257 );
and \U$25009 ( \25262 , \25261 , \6118 );
nor \U$25010 ( \25263 , \25260 , \25262 );
and \U$25011 ( \25264 , \25252 , \25263 );
nor \U$25012 ( \25265 , \25245 , \25251 );
nor \U$25013 ( \25266 , \25264 , \25265 );
not \U$25014 ( \25267 , \25266 );
not \U$25015 ( \25268 , RIbe2a988_100);
not \U$25016 ( \25269 , \6535 );
or \U$25017 ( \25270 , \25268 , \25269 );
nand \U$25018 ( \25271 , \7075 , RIbe2a910_99);
nand \U$25019 ( \25272 , \25270 , \25271 );
not \U$25020 ( \25273 , \25272 );
not \U$25021 ( \25274 , \9933 );
and \U$25022 ( \25275 , \25273 , \25274 );
and \U$25023 ( \25276 , \25272 , \7546 );
nor \U$25024 ( \25277 , \25275 , \25276 );
not \U$25025 ( \25278 , RIbe2a5c8_92);
not \U$25026 ( \25279 , \6138 );
or \U$25027 ( \25280 , \25278 , \25279 );
nand \U$25028 ( \25281 , \7087 , RIbe2a550_91);
nand \U$25029 ( \25282 , \25280 , \25281 );
not \U$25030 ( \25283 , \25282 );
not \U$25031 ( \25284 , \5740 );
and \U$25032 ( \25285 , \25283 , \25284 );
and \U$25033 ( \25286 , \25282 , \6141 );
nor \U$25034 ( \25287 , \25285 , \25286 );
xor \U$25035 ( \25288 , \25277 , \25287 );
not \U$25036 ( \25289 , RIbe2b5b8_126);
not \U$25037 ( \25290 , \7941 );
or \U$25038 ( \25291 , \25289 , \25290 );
nand \U$25039 ( \25292 , \6596 , RIbe2a3e8_88);
nand \U$25040 ( \25293 , \25291 , \25292 );
and \U$25041 ( \25294 , \25293 , \7949 );
not \U$25042 ( \25295 , \25293 );
and \U$25043 ( \25296 , \25295 , \6582 );
nor \U$25044 ( \25297 , \25294 , \25296 );
and \U$25045 ( \25298 , \25288 , \25297 );
and \U$25046 ( \25299 , \25277 , \25287 );
or \U$25047 ( \25300 , \25298 , \25299 );
not \U$25048 ( \25301 , \25300 );
or \U$25049 ( \25302 , \25267 , \25301 );
not \U$25050 ( \25303 , RIbe29fb0_79);
not \U$25051 ( \25304 , \7974 );
or \U$25052 ( \25305 , \25303 , \25304 );
nand \U$25053 ( \25306 , \9891 , RIbe29e48_76);
nand \U$25054 ( \25307 , \25305 , \25306 );
not \U$25055 ( \25308 , \25307 );
not \U$25056 ( \25309 , \6948 );
and \U$25057 ( \25310 , \25308 , \25309 );
and \U$25058 ( \25311 , \25307 , \6948 );
nor \U$25059 ( \25312 , \25310 , \25311 );
not \U$25060 ( \25313 , \25312 );
not \U$25061 ( \25314 , \25313 );
not \U$25062 ( \25315 , RIbe2a370_87);
not \U$25063 ( \25316 , \6958 );
or \U$25064 ( \25317 , \25315 , \25316 );
nand \U$25065 ( \25318 , \7653 , RIbe2a2f8_86);
nand \U$25066 ( \25319 , \25317 , \25318 );
and \U$25067 ( \25320 , \25319 , \6569 );
not \U$25068 ( \25321 , \25319 );
and \U$25069 ( \25322 , \25321 , \7293 );
nor \U$25070 ( \25323 , \25320 , \25322 );
not \U$25071 ( \25324 , \25323 );
not \U$25072 ( \25325 , \25324 );
or \U$25073 ( \25326 , \25314 , \25325 );
not \U$25074 ( \25327 , \25323 );
not \U$25075 ( \25328 , \25312 );
or \U$25076 ( \25329 , \25327 , \25328 );
not \U$25077 ( \25330 , \6992 );
not \U$25078 ( \25331 , RIbe2acd0_107);
not \U$25079 ( \25332 , \6980 );
or \U$25080 ( \25333 , \25331 , \25332 );
nand \U$25081 ( \25334 , \6985 , RIbe2a028_80);
nand \U$25082 ( \25335 , \25333 , \25334 );
not \U$25083 ( \25336 , \25335 );
or \U$25084 ( \25337 , \25330 , \25336 );
or \U$25085 ( \25338 , \25335 , \6992 );
nand \U$25086 ( \25339 , \25337 , \25338 );
nand \U$25087 ( \25340 , \25329 , \25339 );
nand \U$25088 ( \25341 , \25326 , \25340 );
nand \U$25089 ( \25342 , \25302 , \25341 );
not \U$25090 ( \25343 , \25300 );
not \U$25091 ( \25344 , \25266 );
nand \U$25092 ( \25345 , \25343 , \25344 );
nand \U$25093 ( \25346 , \25342 , \25345 );
not \U$25094 ( \25347 , RIbe28b10_35);
not \U$25095 ( \25348 , \13518 );
or \U$25096 ( \25349 , \25347 , \25348 );
nand \U$25097 ( \25350 , \12794 , RIbe28b88_36);
nand \U$25098 ( \25351 , \25349 , \25350 );
and \U$25099 ( \25352 , \25351 , \12801 );
not \U$25100 ( \25353 , \25351 );
and \U$25101 ( \25354 , \25353 , \16334 );
nor \U$25102 ( \25355 , \25352 , \25354 );
not \U$25103 ( \25356 , RIbe29290_51);
not \U$25104 ( \25357 , \12811 );
or \U$25105 ( \25358 , \25356 , \25357 );
nand \U$25106 ( \25359 , RIbe28a20_33, RIbe2ae38_110);
nand \U$25107 ( \25360 , \25358 , \25359 );
xnor \U$25108 ( \25361 , \25360 , RIbe2aeb0_111);
nand \U$25109 ( \25362 , \25355 , \25361 );
not \U$25110 ( \25363 , \12823 );
not \U$25111 ( \25364 , RIbe28408_20);
not \U$25112 ( \25365 , \13590 );
or \U$25113 ( \25366 , \25364 , \25365 );
nand \U$25114 ( \25367 , \21679 , RIbe28390_19);
nand \U$25115 ( \25368 , \25366 , \25367 );
not \U$25116 ( \25369 , \25368 );
or \U$25117 ( \25370 , \25363 , \25369 );
or \U$25118 ( \25371 , \25368 , \15263 );
nand \U$25119 ( \25372 , \25370 , \25371 );
and \U$25120 ( \25373 , \25362 , \25372 );
nor \U$25121 ( \25374 , \25355 , \25361 );
nor \U$25122 ( \25375 , \25373 , \25374 );
not \U$25123 ( \25376 , \25375 );
not \U$25124 ( \25377 , RIbe29bf0_71);
not \U$25125 ( \25378 , \10936 );
or \U$25126 ( \25379 , \25377 , \25378 );
nand \U$25127 ( \25380 , \12971 , RIbe28f48_44);
nand \U$25128 ( \25381 , \25379 , \25380 );
and \U$25129 ( \25382 , \25381 , \19139 );
not \U$25130 ( \25383 , \25381 );
and \U$25131 ( \25384 , \25383 , \13030 );
nor \U$25132 ( \25385 , \25382 , \25384 );
not \U$25133 ( \25386 , \25385 );
and \U$25134 ( \25387 , \16431 , RIbe29dd0_75);
and \U$25135 ( \25388 , \17228 , RIbe29c68_72);
nor \U$25136 ( \25389 , \25387 , \25388 );
and \U$25137 ( \25390 , \25389 , \13384 );
not \U$25138 ( \25391 , \25389 );
and \U$25139 ( \25392 , \25391 , \13383 );
nor \U$25140 ( \25393 , \25390 , \25392 );
nand \U$25141 ( \25394 , \25386 , \25393 );
and \U$25142 ( \25395 , \15205 , RIbe28ed0_43);
and \U$25143 ( \25396 , \12947 , RIbe27fd0_11);
nor \U$25144 ( \25397 , \25395 , \25396 );
and \U$25145 ( \25398 , \25397 , \12195 );
not \U$25146 ( \25399 , \25397 );
and \U$25147 ( \25400 , \25399 , \17005 );
nor \U$25148 ( \25401 , \25398 , \25400 );
not \U$25149 ( \25402 , \25401 );
and \U$25150 ( \25403 , \25394 , \25402 );
nor \U$25151 ( \25404 , \25386 , \25393 );
nor \U$25152 ( \25405 , \25403 , \25404 );
not \U$25153 ( \25406 , \25405 );
or \U$25154 ( \25407 , \25376 , \25406 );
not \U$25155 ( \25408 , RIbe28660_25);
not \U$25156 ( \25409 , \12871 );
or \U$25157 ( \25410 , \25408 , \25409 );
nand \U$25158 ( \25411 , \12711 , RIbe285e8_24);
nand \U$25159 ( \25412 , \25410 , \25411 );
and \U$25160 ( \25413 , \25412 , \12879 );
not \U$25161 ( \25414 , \25412 );
and \U$25162 ( \25415 , \25414 , \12723 );
nor \U$25163 ( \25416 , \25413 , \25415 );
not \U$25164 ( \25417 , \25416 );
not \U$25165 ( \25418 , RIbe287c8_28);
not \U$25166 ( \25419 , \14071 );
or \U$25167 ( \25420 , \25418 , \25419 );
nand \U$25168 ( \25421 , \14074 , RIbe28480_21);
nand \U$25169 ( \25422 , \25420 , \25421 );
and \U$25170 ( \25423 , \25422 , \12746 );
not \U$25171 ( \25424 , \25422 );
and \U$25172 ( \25425 , \25424 , \13570 );
nor \U$25173 ( \25426 , \25423 , \25425 );
not \U$25174 ( \25427 , \25426 );
not \U$25175 ( \25428 , \25427 );
or \U$25176 ( \25429 , \25417 , \25428 );
not \U$25177 ( \25430 , \25426 );
not \U$25178 ( \25431 , \25416 );
not \U$25179 ( \25432 , \25431 );
or \U$25180 ( \25433 , \25430 , \25432 );
not \U$25181 ( \25434 , \12753 );
not \U$25182 ( \25435 , \6347 );
and \U$25183 ( \25436 , \25434 , \25435 );
and \U$25184 ( \25437 , \13738 , RIbe27f58_10);
nor \U$25185 ( \25438 , \25436 , \25437 );
and \U$25186 ( \25439 , \25438 , \12770 );
not \U$25187 ( \25440 , \25438 );
and \U$25188 ( \25441 , \25440 , \12927 );
nor \U$25189 ( \25442 , \25439 , \25441 );
nand \U$25190 ( \25443 , \25433 , \25442 );
nand \U$25191 ( \25444 , \25429 , \25443 );
nand \U$25192 ( \25445 , \25407 , \25444 );
not \U$25193 ( \25446 , \25405 );
not \U$25194 ( \25447 , \25375 );
nand \U$25195 ( \25448 , \25446 , \25447 );
nand \U$25196 ( \25449 , \25445 , \25448 );
nor \U$25197 ( \25450 , \25346 , \25449 );
xor \U$25198 ( \25451 , \24735 , \24726 );
xor \U$25199 ( \25452 , \25451 , \24717 );
not \U$25200 ( \25453 , RIbe2afa0_113);
not \U$25201 ( \25454 , \6797 );
or \U$25202 ( \25455 , \25453 , \25454 );
nand \U$25203 ( \25456 , \3689 , RIbe2af28_112);
nand \U$25204 ( \25457 , \25455 , \25456 );
and \U$25205 ( \25458 , \25457 , \4346 );
not \U$25206 ( \25459 , \25457 );
and \U$25207 ( \25460 , \25459 , \2887 );
nor \U$25208 ( \25461 , \25458 , \25460 );
not \U$25209 ( \25462 , RIbe2b1f8_118);
not \U$25210 ( \25463 , \6783 );
or \U$25211 ( \25464 , \25462 , \25463 );
nand \U$25212 ( \25465 , \8368 , RIbe2b180_117);
nand \U$25213 ( \25466 , \25464 , \25465 );
and \U$25214 ( \25467 , \25466 , \3471 );
not \U$25215 ( \25468 , \25466 );
and \U$25216 ( \25469 , \25468 , \3698 );
nor \U$25217 ( \25470 , \25467 , \25469 );
xor \U$25218 ( \25471 , \25461 , \25470 );
not \U$25219 ( \25472 , RIbe2b630_127);
not \U$25220 ( \25473 , \7827 );
or \U$25221 ( \25474 , \25472 , \25473 );
nand \U$25222 ( \25475 , \4284 , RIbe2b018_114);
nand \U$25223 ( \25476 , \25474 , \25475 );
not \U$25224 ( \25477 , \2576 );
and \U$25225 ( \25478 , \25476 , \25477 );
not \U$25226 ( \25479 , \25476 );
and \U$25227 ( \25480 , \25479 , \4059 );
nor \U$25228 ( \25481 , \25478 , \25480 );
and \U$25229 ( \25482 , \25471 , \25481 );
and \U$25230 ( \25483 , \25461 , \25470 );
or \U$25231 ( \25484 , \25482 , \25483 );
not \U$25232 ( \25485 , \25484 );
nand \U$25233 ( \25486 , \25452 , \25485 );
xor \U$25234 ( \25487 , \24747 , \24754 );
xnor \U$25235 ( \25488 , \25487 , \24765 );
and \U$25236 ( \25489 , \25486 , \25488 );
nor \U$25237 ( \25490 , \25485 , \25452 );
nor \U$25238 ( \25491 , \25489 , \25490 );
or \U$25239 ( \25492 , \25450 , \25491 );
not \U$25240 ( \25493 , \25342 );
not \U$25241 ( \25494 , \25345 );
or \U$25242 ( \25495 , \25493 , \25494 );
nand \U$25243 ( \25496 , \25495 , \25449 );
nand \U$25244 ( \25497 , \25492 , \25496 );
not \U$25245 ( \25498 , \25497 );
nand \U$25246 ( \25499 , \25235 , \25498 );
and \U$25247 ( \25500 , \25172 , \25499 );
and \U$25248 ( \25501 , \25234 , \25497 );
nor \U$25249 ( \25502 , \25500 , \25501 );
buf \U$25250 ( \25503 , \25502 );
xor \U$25251 ( \25504 , \23910 , \23841 );
xnor \U$25252 ( \25505 , \25504 , \23878 );
not \U$25253 ( \25506 , \24007 );
xor \U$25254 ( \25507 , \23976 , \25506 );
and \U$25255 ( \25508 , \25507 , \23943 );
not \U$25256 ( \25509 , \25507 );
and \U$25257 ( \25510 , \25509 , \24010 );
nor \U$25258 ( \25511 , \25508 , \25510 );
nand \U$25259 ( \25512 , \25505 , \25511 );
not \U$25260 ( \25513 , \25512 );
xor \U$25261 ( \25514 , \24898 , \24930 );
xnor \U$25262 ( \25515 , \25514 , \24967 );
not \U$25263 ( \25516 , \25515 );
xor \U$25264 ( \25517 , \24868 , \24871 );
xor \U$25265 ( \25518 , \25517 , \24829 );
not \U$25266 ( \25519 , \25518 );
or \U$25267 ( \25520 , \25516 , \25519 );
xor \U$25268 ( \25521 , \24706 , \24770 );
xnor \U$25269 ( \25522 , \25521 , \24740 );
nand \U$25270 ( \25523 , \25520 , \25522 );
not \U$25271 ( \25524 , \25515 );
not \U$25272 ( \25525 , \25518 );
nand \U$25273 ( \25526 , \25524 , \25525 );
nand \U$25274 ( \25527 , \25523 , \25526 );
not \U$25275 ( \25528 , \25527 );
or \U$25276 ( \25529 , \25513 , \25528 );
not \U$25277 ( \25530 , \25511 );
not \U$25278 ( \25531 , \25505 );
nand \U$25279 ( \25532 , \25530 , \25531 );
nand \U$25280 ( \25533 , \25529 , \25532 );
not \U$25281 ( \25534 , \25533 );
nand \U$25282 ( \25535 , \25503 , \25534 );
not \U$25283 ( \25536 , \25535 );
xor \U$25284 ( \25537 , \24978 , \25029 );
xnor \U$25285 ( \25538 , \25537 , \25032 );
not \U$25286 ( \25539 , \25538 );
not \U$25287 ( \25540 , \25539 );
not \U$25288 ( \25541 , \25047 );
not \U$25289 ( \25542 , \25041 );
or \U$25290 ( \25543 , \25541 , \25542 );
nand \U$25291 ( \25544 , \25040 , \25037 );
nand \U$25292 ( \25545 , \25543 , \25544 );
not \U$25293 ( \25546 , \25045 );
and \U$25294 ( \25547 , \25545 , \25546 );
not \U$25295 ( \25548 , \25545 );
and \U$25296 ( \25549 , \25548 , \25045 );
nor \U$25297 ( \25550 , \25547 , \25549 );
not \U$25298 ( \25551 , \25550 );
not \U$25299 ( \25552 , \25551 );
or \U$25300 ( \25553 , \25540 , \25552 );
not \U$25301 ( \25554 , \25538 );
not \U$25302 ( \25555 , \25550 );
or \U$25303 ( \25556 , \25554 , \25555 );
not \U$25304 ( \25557 , \24874 );
not \U$25305 ( \25558 , \24969 );
or \U$25306 ( \25559 , \25557 , \25558 );
or \U$25307 ( \25560 , \24874 , \24969 );
nand \U$25308 ( \25561 , \25559 , \25560 );
not \U$25309 ( \25562 , \25561 );
buf \U$25310 ( \25563 , \24774 );
not \U$25311 ( \25564 , \25563 );
and \U$25312 ( \25565 , \25562 , \25564 );
and \U$25313 ( \25566 , \25561 , \25563 );
nor \U$25314 ( \25567 , \25565 , \25566 );
not \U$25315 ( \25568 , \25567 );
nand \U$25316 ( \25569 , \25556 , \25568 );
nand \U$25317 ( \25570 , \25553 , \25569 );
not \U$25318 ( \25571 , \25570 );
or \U$25319 ( \25572 , \25536 , \25571 );
or \U$25320 ( \25573 , \25503 , \25534 );
nand \U$25321 ( \25574 , \25572 , \25573 );
not \U$25322 ( \25575 , \25574 );
not \U$25323 ( \25576 , \25575 );
not \U$25324 ( \25577 , \24693 );
not \U$25325 ( \25578 , \24686 );
or \U$25326 ( \25579 , \25577 , \25578 );
or \U$25327 ( \25580 , \24686 , \24693 );
nand \U$25328 ( \25581 , \25579 , \25580 );
xor \U$25329 ( \25582 , \24973 , \25034 );
xor \U$25330 ( \25583 , \25582 , \25049 );
xor \U$25331 ( \25584 , \25581 , \25583 );
not \U$25332 ( \25585 , \25070 );
not \U$25333 ( \25586 , \25060 );
or \U$25334 ( \25587 , \25585 , \25586 );
or \U$25335 ( \25588 , \25060 , \25070 );
nand \U$25336 ( \25589 , \25587 , \25588 );
xor \U$25337 ( \25590 , \24311 , \25589 );
xnor \U$25338 ( \25591 , \25590 , \25077 );
and \U$25339 ( \25592 , \25584 , \25591 );
and \U$25340 ( \25593 , \25581 , \25583 );
or \U$25341 ( \25594 , \25592 , \25593 );
not \U$25342 ( \25595 , \25594 );
not \U$25343 ( \25596 , \25595 );
or \U$25344 ( \25597 , \25576 , \25596 );
not \U$25345 ( \25598 , \25106 );
not \U$25346 ( \25599 , \25111 );
not \U$25347 ( \25600 , \25599 );
or \U$25348 ( \25601 , \25598 , \25600 );
nand \U$25349 ( \25602 , \25103 , \25111 );
nand \U$25350 ( \25603 , \25601 , \25602 );
and \U$25351 ( \25604 , \25603 , \25097 );
not \U$25352 ( \25605 , \25603 );
and \U$25353 ( \25606 , \25605 , \25096 );
nor \U$25354 ( \25607 , \25604 , \25606 );
nand \U$25355 ( \25608 , \25597 , \25607 );
not \U$25356 ( \25609 , \25595 );
nand \U$25357 ( \25610 , \25609 , \25574 );
nand \U$25358 ( \25611 , \25608 , \25610 );
xor \U$25359 ( \25612 , \25150 , \25611 );
xor \U$25360 ( \25613 , \25089 , \25114 );
xor \U$25361 ( \25614 , \25613 , \25117 );
and \U$25362 ( \25615 , \25612 , \25614 );
and \U$25363 ( \25616 , \25150 , \25611 );
or \U$25364 ( \25617 , \25615 , \25616 );
not \U$25365 ( \25618 , \25617 );
xor \U$25366 ( \25619 , \25125 , \25120 );
xor \U$25367 ( \25620 , \25619 , \25129 );
not \U$25368 ( \25621 , \25620 );
or \U$25369 ( \25622 , \25618 , \25621 );
or \U$25370 ( \25623 , \25620 , \25617 );
nand \U$25371 ( \25624 , \25622 , \25623 );
and \U$25372 ( \25625 , \24658 , \25139 , \25624 );
not \U$25373 ( \25626 , \25625 );
not \U$25374 ( \25627 , \16575 );
nand \U$25375 ( \25628 , \25627 , \16565 );
not \U$25376 ( \25629 , \25628 );
not \U$25377 ( \25630 , \16556 );
or \U$25378 ( \25631 , \25629 , \25630 );
not \U$25379 ( \25632 , \16565 );
nand \U$25380 ( \25633 , \25632 , \16575 );
nand \U$25381 ( \25634 , \25631 , \25633 );
not \U$25382 ( \25635 , \25634 );
not \U$25383 ( \25636 , \25635 );
not \U$25384 ( \25637 , \16624 );
not \U$25385 ( \25638 , \16620 );
and \U$25386 ( \25639 , \25637 , \25638 );
nor \U$25387 ( \25640 , \25639 , \16629 );
and \U$25388 ( \25641 , \16620 , \16624 );
nor \U$25389 ( \25642 , \25640 , \25641 );
not \U$25390 ( \25643 , \25642 );
or \U$25391 ( \25644 , \25636 , \25643 );
not \U$25392 ( \25645 , \16586 );
not \U$25393 ( \25646 , \16593 );
or \U$25394 ( \25647 , \25645 , \25646 );
not \U$25395 ( \25648 , \16586 );
nand \U$25396 ( \25649 , \25648 , \16594 );
nand \U$25397 ( \25650 , \16606 , \25649 );
nand \U$25398 ( \25651 , \25647 , \25650 );
nand \U$25399 ( \25652 , \25644 , \25651 );
not \U$25400 ( \25653 , \25642 );
nand \U$25401 ( \25654 , \25653 , \25634 );
nand \U$25402 ( \25655 , \25652 , \25654 );
not \U$25403 ( \25656 , RIbe28390_19);
not \U$25404 ( \25657 , \13690 );
or \U$25405 ( \25658 , \25656 , \25657 );
nand \U$25406 ( \25659 , RIbe28b10_35, RIbe2ae38_110);
nand \U$25407 ( \25660 , \25658 , \25659 );
xnor \U$25408 ( \25661 , \25660 , RIbe2aeb0_111);
not \U$25409 ( \25662 , \25661 );
and \U$25410 ( \25663 , \25662 , \2576 );
not \U$25411 ( \25664 , \25662 );
and \U$25412 ( \25665 , \25664 , \3481 );
nor \U$25413 ( \25666 , \25663 , \25665 );
not \U$25414 ( \25667 , \25666 );
not \U$25415 ( \25668 , RIbe28480_21);
not \U$25416 ( \25669 , \12786 );
or \U$25417 ( \25670 , \25668 , \25669 );
nand \U$25418 ( \25671 , RIbe28408_20, \12890 );
nand \U$25419 ( \25672 , \25670 , \25671 );
and \U$25420 ( \25673 , \25672 , \12801 );
not \U$25421 ( \25674 , \25672 );
and \U$25422 ( \25675 , \25674 , \16334 );
or \U$25423 ( \25676 , \25673 , \25675 );
not \U$25424 ( \25677 , \25676 );
or \U$25425 ( \25678 , \25667 , \25677 );
or \U$25426 ( \25679 , \25666 , \25676 );
nand \U$25427 ( \25680 , \25678 , \25679 );
nand \U$25428 ( \25681 , \3267 , RIbe2ab68_104);
and \U$25429 ( \25682 , \25681 , \2379 );
not \U$25430 ( \25683 , \25681 );
and \U$25431 ( \25684 , \25683 , \7457 );
nor \U$25432 ( \25685 , \25682 , \25684 );
not \U$25433 ( \25686 , RIbe2af28_112);
not \U$25434 ( \25687 , \4317 );
or \U$25435 ( \25688 , \25686 , \25687 );
nand \U$25436 ( \25689 , \7858 , RIbe2b1f8_118);
nand \U$25437 ( \25690 , \25688 , \25689 );
and \U$25438 ( \25691 , \25690 , \4007 );
not \U$25439 ( \25692 , \25690 );
and \U$25440 ( \25693 , \25692 , \7865 );
nor \U$25441 ( \25694 , \25691 , \25693 );
not \U$25442 ( \25695 , \25694 );
not \U$25443 ( \25696 , RIbe2b018_114);
not \U$25444 ( \25697 , \7880 );
or \U$25445 ( \25698 , \25696 , \25697 );
nand \U$25446 ( \25699 , \7438 , RIbe2afa0_113);
nand \U$25447 ( \25700 , \25698 , \25699 );
not \U$25448 ( \25701 , \25700 );
not \U$25449 ( \25702 , \3698 );
and \U$25450 ( \25703 , \25701 , \25702 );
and \U$25451 ( \25704 , \25700 , \3448 );
nor \U$25452 ( \25705 , \25703 , \25704 );
not \U$25453 ( \25706 , \25705 );
or \U$25454 ( \25707 , \25695 , \25706 );
or \U$25455 ( \25708 , \25694 , \25705 );
nand \U$25456 ( \25709 , \25707 , \25708 );
not \U$25457 ( \25710 , RIbe2aaf0_103);
not \U$25458 ( \25711 , \3452 );
or \U$25459 ( \25712 , \25710 , \25711 );
nand \U$25460 ( \25713 , \4011 , RIbe2b630_127);
nand \U$25461 ( \25714 , \25712 , \25713 );
and \U$25462 ( \25715 , \25714 , \3461 );
not \U$25463 ( \25716 , \25714 );
and \U$25464 ( \25717 , \25716 , \3290 );
nor \U$25465 ( \25718 , \25715 , \25717 );
not \U$25466 ( \25719 , \25718 );
and \U$25467 ( \25720 , \25709 , \25719 );
not \U$25468 ( \25721 , \25709 );
and \U$25469 ( \25722 , \25721 , \25718 );
nor \U$25470 ( \25723 , \25720 , \25722 );
xor \U$25471 ( \25724 , \25685 , \25723 );
not \U$25472 ( \25725 , RIbe2b108_116);
not \U$25473 ( \25726 , \5455 );
or \U$25474 ( \25727 , \25725 , \25726 );
nand \U$25475 ( \25728 , \6634 , RIbe2b090_115);
nand \U$25476 ( \25729 , \25727 , \25728 );
and \U$25477 ( \25730 , \25729 , \25258 );
not \U$25478 ( \25731 , \25729 );
and \U$25479 ( \25732 , \25731 , \6117 );
nor \U$25480 ( \25733 , \25730 , \25732 );
not \U$25481 ( \25734 , RIbe2a280_85);
not \U$25482 ( \25735 , \12268 );
or \U$25483 ( \25736 , \25734 , \25735 );
nand \U$25484 ( \25737 , \7087 , RIbe2a208_84);
nand \U$25485 ( \25738 , \25736 , \25737 );
and \U$25486 ( \25739 , \25738 , \7535 );
not \U$25487 ( \25740 , \25738 );
and \U$25488 ( \25741 , \25740 , \10969 );
nor \U$25489 ( \25742 , \25739 , \25741 );
not \U$25490 ( \25743 , \25742 );
and \U$25491 ( \25744 , \25733 , \25743 );
not \U$25492 ( \25745 , \25733 );
and \U$25493 ( \25746 , \25745 , \25742 );
or \U$25494 ( \25747 , \25744 , \25746 );
not \U$25495 ( \25748 , RIbe2b180_117);
not \U$25496 ( \25749 , \15894 );
or \U$25497 ( \25750 , \25748 , \25749 );
nand \U$25498 ( \25751 , \5052 , RIbe2b270_119);
nand \U$25499 ( \25752 , \25750 , \25751 );
not \U$25500 ( \25753 , \25752 );
not \U$25501 ( \25754 , \4592 );
and \U$25502 ( \25755 , \25753 , \25754 );
and \U$25503 ( \25756 , \25752 , \4592 );
nor \U$25504 ( \25757 , \25755 , \25756 );
not \U$25505 ( \25758 , \25757 );
and \U$25506 ( \25759 , \25747 , \25758 );
not \U$25507 ( \25760 , \25747 );
and \U$25508 ( \25761 , \25760 , \25757 );
nor \U$25509 ( \25762 , \25759 , \25761 );
xor \U$25510 ( \25763 , \25724 , \25762 );
xor \U$25511 ( \25764 , \25680 , \25763 );
not \U$25512 ( \25765 , \12752 );
not \U$25513 ( \25766 , \6757 );
and \U$25514 ( \25767 , \25765 , \25766 );
and \U$25515 ( \25768 , \13738 , RIbe28f48_44);
nor \U$25516 ( \25769 , \25767 , \25768 );
and \U$25517 ( \25770 , \25769 , \12927 );
not \U$25518 ( \25771 , \25769 );
and \U$25519 ( \25772 , \25771 , \12924 );
nor \U$25520 ( \25773 , \25770 , \25772 );
not \U$25521 ( \25774 , \25773 );
and \U$25522 ( \25775 , \15205 , RIbe29c68_72);
not \U$25523 ( \25776 , RIbe29bf0_71);
nor \U$25524 ( \25777 , \25776 , \15627 );
nor \U$25525 ( \25778 , \25775 , \25777 );
and \U$25526 ( \25779 , \25778 , \12960 );
not \U$25527 ( \25780 , \25778 );
and \U$25528 ( \25781 , \25780 , \12195 );
nor \U$25529 ( \25782 , \25779 , \25781 );
not \U$25530 ( \25783 , \25782 );
or \U$25531 ( \25784 , \25774 , \25783 );
not \U$25532 ( \25785 , \25782 );
not \U$25533 ( \25786 , \25773 );
nand \U$25534 ( \25787 , \25785 , \25786 );
nand \U$25535 ( \25788 , \25784 , \25787 );
not \U$25536 ( \25789 , RIbe29e48_76);
not \U$25537 ( \25790 , \10936 );
or \U$25538 ( \25791 , \25789 , \25790 );
nand \U$25539 ( \25792 , \12971 , RIbe29dd0_75);
nand \U$25540 ( \25793 , \25791 , \25792 );
and \U$25541 ( \25794 , \25793 , \19136 );
not \U$25542 ( \25795 , \25793 );
and \U$25543 ( \25796 , \25795 , \10940 );
nor \U$25544 ( \25797 , \25794 , \25796 );
not \U$25545 ( \25798 , \25797 );
and \U$25546 ( \25799 , \25788 , \25798 );
not \U$25547 ( \25800 , \25788 );
and \U$25548 ( \25801 , \25800 , \25797 );
nor \U$25549 ( \25802 , \25799 , \25801 );
and \U$25550 ( \25803 , \21196 , RIbe2a028_80);
and \U$25551 ( \25804 , \10919 , RIbe29fb0_79);
nor \U$25552 ( \25805 , \25803 , \25804 );
and \U$25553 ( \25806 , \25805 , \7970 );
not \U$25554 ( \25807 , \25805 );
not \U$25555 ( \25808 , \7970 );
and \U$25556 ( \25809 , \25807 , \25808 );
nor \U$25557 ( \25810 , \25806 , \25809 );
not \U$25558 ( \25811 , \25810 );
not \U$25559 ( \25812 , RIbe2a2f8_86);
not \U$25560 ( \25813 , \14633 );
or \U$25561 ( \25814 , \25812 , \25813 );
nand \U$25562 ( \25815 , \8269 , RIbe2acd0_107);
nand \U$25563 ( \25816 , \25814 , \25815 );
and \U$25564 ( \25817 , \25816 , \8480 );
not \U$25565 ( \25818 , \25816 );
and \U$25566 ( \25819 , \25818 , \7989 );
nor \U$25567 ( \25820 , \25817 , \25819 );
not \U$25568 ( \25821 , \25820 );
or \U$25569 ( \25822 , \25811 , \25821 );
not \U$25570 ( \25823 , \25810 );
not \U$25571 ( \25824 , \25820 );
nand \U$25572 ( \25825 , \25823 , \25824 );
nand \U$25573 ( \25826 , \25822 , \25825 );
not \U$25574 ( \25827 , \6992 );
not \U$25575 ( \25828 , RIbe2a3e8_88);
not \U$25576 ( \25829 , \7298 );
or \U$25577 ( \25830 , \25828 , \25829 );
nand \U$25578 ( \25831 , \8287 , RIbe2a370_87);
nand \U$25579 ( \25832 , \25830 , \25831 );
not \U$25580 ( \25833 , \25832 );
or \U$25581 ( \25834 , \25827 , \25833 );
or \U$25582 ( \25835 , \25832 , \10902 );
nand \U$25583 ( \25836 , \25834 , \25835 );
not \U$25584 ( \25837 , \25836 );
and \U$25585 ( \25838 , \25826 , \25837 );
not \U$25586 ( \25839 , \25826 );
and \U$25587 ( \25840 , \25839 , \25836 );
nor \U$25588 ( \25841 , \25838 , \25840 );
xor \U$25589 ( \25842 , \25802 , \25841 );
not \U$25590 ( \25843 , \6572 );
not \U$25591 ( \25844 , RIbe2a910_99);
not \U$25592 ( \25845 , \6560 );
or \U$25593 ( \25846 , \25844 , \25845 );
nand \U$25594 ( \25847 , \7958 , RIbe2b5b8_126);
nand \U$25595 ( \25848 , \25846 , \25847 );
not \U$25596 ( \25849 , \25848 );
or \U$25597 ( \25850 , \25843 , \25849 );
or \U$25598 ( \25851 , \25848 , \6572 );
nand \U$25599 ( \25852 , \25850 , \25851 );
not \U$25600 ( \25853 , \25852 );
not \U$25601 ( \25854 , RIbe2a550_91);
not \U$25602 ( \25855 , \6591 );
or \U$25603 ( \25856 , \25854 , \25855 );
nand \U$25604 ( \25857 , \7278 , RIbe2a988_100);
nand \U$25605 ( \25858 , \25856 , \25857 );
and \U$25606 ( \25859 , \25858 , \14666 );
not \U$25607 ( \25860 , \25858 );
and \U$25608 ( \25861 , \25860 , \6582 );
nor \U$25609 ( \25862 , \25859 , \25861 );
not \U$25610 ( \25863 , \25862 );
or \U$25611 ( \25864 , \25853 , \25863 );
or \U$25612 ( \25865 , \25862 , \25852 );
nand \U$25613 ( \25866 , \25864 , \25865 );
not \U$25614 ( \25867 , RIbe2a190_83);
not \U$25615 ( \25868 , \6536 );
or \U$25616 ( \25869 , \25867 , \25868 );
nand \U$25617 ( \25870 , \10348 , RIbe2a5c8_92);
nand \U$25618 ( \25871 , \25869 , \25870 );
xor \U$25619 ( \25872 , \25871 , \9933 );
and \U$25620 ( \25873 , \25866 , \25872 );
not \U$25621 ( \25874 , \25866 );
not \U$25622 ( \25875 , \25872 );
and \U$25623 ( \25876 , \25874 , \25875 );
nor \U$25624 ( \25877 , \25873 , \25876 );
not \U$25625 ( \25878 , \25877 );
and \U$25626 ( \25879 , \25842 , \25878 );
not \U$25627 ( \25880 , \25842 );
and \U$25628 ( \25881 , \25880 , \25877 );
nor \U$25629 ( \25882 , \25879 , \25881 );
and \U$25630 ( \25883 , \25764 , \25882 );
and \U$25631 ( \25884 , \25680 , \25763 );
or \U$25632 ( \25885 , \25883 , \25884 );
xor \U$25633 ( \25886 , \25655 , \25885 );
not \U$25634 ( \25887 , RIbe27fd0_11);
not \U$25635 ( \25888 , \19262 );
or \U$25636 ( \25889 , \25887 , \25888 );
nand \U$25637 ( \25890 , \13728 , RIbe27f58_10);
nand \U$25638 ( \25891 , \25889 , \25890 );
and \U$25639 ( \25892 , \25891 , \12879 );
not \U$25640 ( \25893 , \25891 );
and \U$25641 ( \25894 , \25893 , \13583 );
nor \U$25642 ( \25895 , \25892 , \25894 );
not \U$25643 ( \25896 , RIbe27e68_8);
not \U$25644 ( \25897 , \14071 );
or \U$25645 ( \25898 , \25896 , \25897 );
not \U$25646 ( \25899 , RIbe28660_25);
not \U$25647 ( \25900 , \25899 );
nand \U$25648 ( \25901 , \25900 , \14074 );
nand \U$25649 ( \25902 , \25898 , \25901 );
and \U$25650 ( \25903 , \25902 , \12852 );
not \U$25651 ( \25904 , \25902 );
and \U$25652 ( \25905 , \25904 , \12746 );
nor \U$25653 ( \25906 , \25903 , \25905 );
not \U$25654 ( \25907 , RIbe285e8_24);
not \U$25655 ( \25908 , \13590 );
or \U$25656 ( \25909 , \25907 , \25908 );
nand \U$25657 ( \25910 , \13012 , RIbe287c8_28);
nand \U$25658 ( \25911 , \25909 , \25910 );
and \U$25659 ( \25912 , \25911 , \14555 );
not \U$25660 ( \25913 , \25911 );
and \U$25661 ( \25914 , \25913 , \12863 );
nor \U$25662 ( \25915 , \25912 , \25914 );
xor \U$25663 ( \25916 , \25906 , \25915 );
xnor \U$25664 ( \25917 , \25895 , \25916 );
xor \U$25665 ( \25918 , \16783 , \16809 );
and \U$25666 ( \25919 , \25918 , \16838 );
and \U$25667 ( \25920 , \16783 , \16809 );
or \U$25668 ( \25921 , \25919 , \25920 );
xor \U$25669 ( \25922 , \25917 , \25921 );
xor \U$25670 ( \25923 , \16672 , \16706 );
and \U$25671 ( \25924 , \25923 , \16744 );
and \U$25672 ( \25925 , \16672 , \16706 );
or \U$25673 ( \25926 , \25924 , \25925 );
and \U$25674 ( \25927 , \25922 , \25926 );
and \U$25675 ( \25928 , \25917 , \25921 );
or \U$25676 ( \25929 , \25927 , \25928 );
xor \U$25677 ( \25930 , \25886 , \25929 );
xor \U$25678 ( \25931 , \25680 , \25763 );
xor \U$25679 ( \25932 , \25931 , \25882 );
not \U$25680 ( \25933 , \16742 );
not \U$25681 ( \25934 , \16731 );
or \U$25682 ( \25935 , \25933 , \25934 );
not \U$25683 ( \25936 , \16727 );
nand \U$25684 ( \25937 , \16716 , \16739 );
nand \U$25685 ( \25938 , \25936 , \25937 );
nand \U$25686 ( \25939 , \25935 , \25938 );
not \U$25687 ( \25940 , \25939 );
not \U$25688 ( \25941 , \16681 );
not \U$25689 ( \25942 , \16705 );
or \U$25690 ( \25943 , \25941 , \25942 );
or \U$25691 ( \25944 , \16705 , \16681 );
not \U$25692 ( \25945 , \16692 );
nand \U$25693 ( \25946 , \25944 , \25945 );
nand \U$25694 ( \25947 , \25943 , \25946 );
not \U$25695 ( \25948 , \16671 );
not \U$25696 ( \25949 , \16657 );
or \U$25697 ( \25950 , \25948 , \25949 );
or \U$25698 ( \25951 , \16657 , \16671 );
nand \U$25699 ( \25952 , \25951 , \16647 );
nand \U$25700 ( \25953 , \25950 , \25952 );
xnor \U$25701 ( \25954 , \25947 , \25953 );
not \U$25702 ( \25955 , \25954 );
or \U$25703 ( \25956 , \25940 , \25955 );
or \U$25704 ( \25957 , \25954 , \25939 );
nand \U$25705 ( \25958 , \25956 , \25957 );
not \U$25706 ( \25959 , \25958 );
xor \U$25707 ( \25960 , \16816 , \16826 );
and \U$25708 ( \25961 , \25960 , \16837 );
and \U$25709 ( \25962 , \16816 , \16826 );
or \U$25710 ( \25963 , \25961 , \25962 );
not \U$25711 ( \25964 , \25963 );
not \U$25712 ( \25965 , \16771 );
not \U$25713 ( \25966 , \16756 );
or \U$25714 ( \25967 , \25965 , \25966 );
nand \U$25715 ( \25968 , \25967 , \16782 );
not \U$25716 ( \25969 , \16771 );
nand \U$25717 ( \25970 , \25969 , \16770 );
nand \U$25718 ( \25971 , \25968 , \25970 );
not \U$25719 ( \25972 , \25971 );
and \U$25720 ( \25973 , \25964 , \25972 );
and \U$25721 ( \25974 , \25963 , \25971 );
nor \U$25722 ( \25975 , \25973 , \25974 );
not \U$25723 ( \25976 , \16789 );
not \U$25724 ( \25977 , \16798 );
or \U$25725 ( \25978 , \25976 , \25977 );
or \U$25726 ( \25979 , \16798 , \16789 );
nand \U$25727 ( \25980 , \25979 , \16808 );
nand \U$25728 ( \25981 , \25978 , \25980 );
xor \U$25729 ( \25982 , \25975 , \25981 );
not \U$25730 ( \25983 , \25982 );
and \U$25731 ( \25984 , \25959 , \25983 );
and \U$25732 ( \25985 , \25958 , \25982 );
nor \U$25733 ( \25986 , \25984 , \25985 );
xor \U$25734 ( \25987 , \25932 , \25986 );
xor \U$25735 ( \25988 , \25635 , \25651 );
xnor \U$25736 ( \25989 , \25988 , \25642 );
nand \U$25737 ( \25990 , \25987 , \25989 );
not \U$25738 ( \25991 , \16843 );
nand \U$25739 ( \25992 , \16745 , \25991 );
not \U$25740 ( \25993 , \16839 );
and \U$25741 ( \25994 , \25992 , \25993 );
nor \U$25742 ( \25995 , \16745 , \25991 );
nor \U$25743 ( \25996 , \25994 , \25995 );
not \U$25744 ( \25997 , \25996 );
not \U$25745 ( \25998 , \16581 );
not \U$25746 ( \25999 , \16608 );
or \U$25747 ( \26000 , \25998 , \25999 );
nand \U$25748 ( \26001 , \26000 , \16630 );
not \U$25749 ( \26002 , \16581 );
nand \U$25750 ( \26003 , \26002 , \16609 );
nand \U$25751 ( \26004 , \26001 , \26003 );
not \U$25752 ( \26005 , \16529 );
not \U$25753 ( \26006 , \26005 );
not \U$25754 ( \26007 , \16538 );
or \U$25755 ( \26008 , \26006 , \26007 );
nand \U$25756 ( \26009 , \26008 , \16544 );
nand \U$25757 ( \26010 , \16537 , \16529 );
nand \U$25758 ( \26011 , \26009 , \26010 );
xor \U$25759 ( \26012 , \26004 , \26011 );
not \U$25760 ( \26013 , \26012 );
or \U$25761 ( \26014 , \25997 , \26013 );
or \U$25762 ( \26015 , \26012 , \25996 );
nand \U$25763 ( \26016 , \26014 , \26015 );
and \U$25764 ( \26017 , \25990 , \26016 );
nor \U$25765 ( \26018 , \25987 , \25989 );
nor \U$25766 ( \26019 , \26017 , \26018 );
xor \U$25767 ( \26020 , \25930 , \26019 );
nand \U$25768 ( \26021 , \16631 , \16545 );
and \U$25769 ( \26022 , \26021 , \16848 );
nor \U$25770 ( \26023 , \16631 , \16545 );
nor \U$25771 ( \26024 , \26022 , \26023 );
xor \U$25772 ( \26025 , \25917 , \25921 );
xor \U$25773 ( \26026 , \26025 , \25926 );
nand \U$25774 ( \26027 , \26024 , \26026 );
not \U$25775 ( \26028 , \16494 );
not \U$25776 ( \26029 , \16489 );
or \U$25777 ( \26030 , \26028 , \26029 );
or \U$25778 ( \26031 , \16489 , \16494 );
nand \U$25779 ( \26032 , \26031 , \16503 );
nand \U$25780 ( \26033 , \26030 , \26032 );
and \U$25781 ( \26034 , \26027 , \26033 );
nor \U$25782 ( \26035 , \26024 , \26026 );
nor \U$25783 ( \26036 , \26034 , \26035 );
and \U$25784 ( \26037 , \26020 , \26036 );
and \U$25785 ( \26038 , \25930 , \26019 );
or \U$25786 ( \26039 , \26037 , \26038 );
not \U$25787 ( \26040 , \26039 );
not \U$25788 ( \26041 , \25996 );
or \U$25789 ( \26042 , \26011 , \26004 );
and \U$25790 ( \26043 , \26041 , \26042 );
and \U$25791 ( \26044 , \26004 , \26011 );
nor \U$25792 ( \26045 , \26043 , \26044 );
not \U$25793 ( \26046 , \26045 );
not \U$25794 ( \26047 , \26046 );
not \U$25795 ( \26048 , \25958 );
nand \U$25796 ( \26049 , \26048 , \25982 );
and \U$25797 ( \26050 , \25932 , \26049 );
not \U$25798 ( \26051 , \25958 );
nor \U$25799 ( \26052 , \26051 , \25982 );
nor \U$25800 ( \26053 , \26050 , \26052 );
not \U$25801 ( \26054 , \26053 );
not \U$25802 ( \26055 , \26054 );
or \U$25803 ( \26056 , \26047 , \26055 );
nor \U$25804 ( \26057 , \25981 , \25971 );
or \U$25805 ( \26058 , \25963 , \26057 );
nand \U$25806 ( \26059 , \25981 , \25971 );
nand \U$25807 ( \26060 , \26058 , \26059 );
or \U$25808 ( \26061 , \25939 , \25953 );
nand \U$25809 ( \26062 , \26061 , \25947 );
nand \U$25810 ( \26063 , \25953 , \25939 );
nand \U$25811 ( \26064 , \26062 , \26063 );
xor \U$25812 ( \26065 , \26060 , \26064 );
xor \U$25813 ( \26066 , \25685 , \25723 );
and \U$25814 ( \26067 , \26066 , \25762 );
and \U$25815 ( \26068 , \25685 , \25723 );
or \U$25816 ( \26069 , \26067 , \26068 );
xor \U$25817 ( \26070 , \26065 , \26069 );
not \U$25818 ( \26071 , \7546 );
not \U$25819 ( \26072 , RIbe2a5c8_92);
not \U$25820 ( \26073 , \6535 );
or \U$25821 ( \26074 , \26072 , \26073 );
not \U$25822 ( \26075 , \21491 );
nand \U$25823 ( \26076 , \26075 , \6540 );
nand \U$25824 ( \26077 , \26074 , \26076 );
not \U$25825 ( \26078 , \26077 );
or \U$25826 ( \26079 , \26071 , \26078 );
or \U$25827 ( \26080 , \26077 , \13412 );
nand \U$25828 ( \26081 , \26079 , \26080 );
not \U$25829 ( \26082 , \7646 );
not \U$25830 ( \26083 , RIbe2a988_100);
not \U$25831 ( \26084 , \7941 );
or \U$25832 ( \26085 , \26083 , \26084 );
nand \U$25833 ( \26086 , \13436 , RIbe2a910_99);
nand \U$25834 ( \26087 , \26085 , \26086 );
not \U$25835 ( \26088 , \26087 );
or \U$25836 ( \26089 , \26082 , \26088 );
or \U$25837 ( \26090 , \26087 , \14262 );
nand \U$25838 ( \26091 , \26089 , \26090 );
xor \U$25839 ( \26092 , \26081 , \26091 );
not \U$25840 ( \26093 , RIbe2a208_84);
not \U$25841 ( \26094 , \12268 );
or \U$25842 ( \26095 , \26093 , \26094 );
nand \U$25843 ( \26096 , \8235 , RIbe2a190_83);
nand \U$25844 ( \26097 , \26095 , \26096 );
and \U$25845 ( \26098 , \26097 , \6144 );
not \U$25846 ( \26099 , \26097 );
and \U$25847 ( \26100 , \26099 , \6141 );
nor \U$25848 ( \26101 , \26098 , \26100 );
xor \U$25849 ( \26102 , \26092 , \26101 );
and \U$25850 ( \26103 , \16431 , RIbe29fb0_79);
and \U$25851 ( \26104 , \10919 , RIbe29e48_76);
nor \U$25852 ( \26105 , \26103 , \26104 );
and \U$25853 ( \26106 , \26105 , \16437 );
not \U$25854 ( \26107 , \26105 );
and \U$25855 ( \26108 , \26107 , \12202 );
nor \U$25856 ( \26109 , \26106 , \26108 );
not \U$25857 ( \26110 , RIbe29dd0_75);
not \U$25858 ( \26111 , \13024 );
or \U$25859 ( \26112 , \26110 , \26111 );
nand \U$25860 ( \26113 , \12971 , RIbe29c68_72);
nand \U$25861 ( \26114 , \26112 , \26113 );
not \U$25862 ( \26115 , \26114 );
not \U$25863 ( \26116 , \13033 );
and \U$25864 ( \26117 , \26115 , \26116 );
and \U$25865 ( \26118 , \26114 , \10940 );
nor \U$25866 ( \26119 , \26117 , \26118 );
xor \U$25867 ( \26120 , \26109 , \26119 );
not \U$25868 ( \26121 , RIbe29bf0_71);
not \U$25869 ( \26122 , \12942 );
or \U$25870 ( \26123 , \26121 , \26122 );
nand \U$25871 ( \26124 , \12947 , RIbe28f48_44);
nand \U$25872 ( \26125 , \26123 , \26124 );
not \U$25873 ( \26126 , \26125 );
not \U$25874 ( \26127 , \12960 );
and \U$25875 ( \26128 , \26126 , \26127 );
and \U$25876 ( \26129 , \26125 , \12956 );
nor \U$25877 ( \26130 , \26128 , \26129 );
xor \U$25878 ( \26131 , \26120 , \26130 );
xor \U$25879 ( \26132 , \26102 , \26131 );
not \U$25880 ( \26133 , RIbe2a370_87);
not \U$25881 ( \26134 , \7298 );
or \U$25882 ( \26135 , \26133 , \26134 );
nand \U$25883 ( \26136 , \13792 , RIbe2a2f8_86);
nand \U$25884 ( \26137 , \26135 , \26136 );
not \U$25885 ( \26138 , \26137 );
not \U$25886 ( \26139 , \7301 );
and \U$25887 ( \26140 , \26138 , \26139 );
and \U$25888 ( \26141 , \26137 , \7661 );
nor \U$25889 ( \26142 , \26140 , \26141 );
not \U$25890 ( \26143 , RIbe2acd0_107);
not \U$25891 ( \26144 , \6942 );
or \U$25892 ( \26145 , \26143 , \26144 );
not \U$25893 ( \26146 , \14374 );
nand \U$25894 ( \26147 , \26146 , \10952 );
nand \U$25895 ( \26148 , \26145 , \26147 );
xor \U$25896 ( \26149 , \26148 , \14302 );
xor \U$25897 ( \26150 , \26142 , \26149 );
not \U$25898 ( \26151 , RIbe2b5b8_126);
not \U$25899 ( \26152 , \6561 );
or \U$25900 ( \26153 , \26151 , \26152 );
nand \U$25901 ( \26154 , \7958 , RIbe2a3e8_88);
nand \U$25902 ( \26155 , \26153 , \26154 );
not \U$25903 ( \26156 , \26155 );
not \U$25904 ( \26157 , \6572 );
and \U$25905 ( \26158 , \26156 , \26157 );
and \U$25906 ( \26159 , \26155 , \6572 );
nor \U$25907 ( \26160 , \26158 , \26159 );
xor \U$25908 ( \26161 , \26150 , \26160 );
xor \U$25909 ( \26162 , \26132 , \26161 );
and \U$25910 ( \26163 , \25877 , \25841 );
nor \U$25911 ( \26164 , \26163 , \25802 );
nor \U$25912 ( \26165 , \25877 , \25841 );
nor \U$25913 ( \26166 , \26164 , \26165 );
not \U$25914 ( \26167 , \12752 );
not \U$25915 ( \26168 , \7360 );
and \U$25916 ( \26169 , \26167 , \26168 );
and \U$25917 ( \26170 , \13738 , RIbe28ed0_43);
nor \U$25918 ( \26171 , \26169 , \26170 );
not \U$25919 ( \26172 , \13999 );
and \U$25920 ( \26173 , \26171 , \26172 );
not \U$25921 ( \26174 , \26171 );
and \U$25922 ( \26175 , \26174 , \12927 );
nor \U$25923 ( \26176 , \26173 , \26175 );
not \U$25924 ( \26177 , RIbe27f58_10);
not \U$25925 ( \26178 , \19262 );
or \U$25926 ( \26179 , \26177 , \26178 );
nand \U$25927 ( \26180 , \12711 , RIbe27e68_8);
nand \U$25928 ( \26181 , \26179 , \26180 );
and \U$25929 ( \26182 , \26181 , \12716 );
not \U$25930 ( \26183 , \26181 );
and \U$25931 ( \26184 , \26183 , \12723 );
nor \U$25932 ( \26185 , \26182 , \26184 );
xor \U$25933 ( \26186 , \26176 , \26185 );
not \U$25934 ( \26187 , RIbe28660_25);
not \U$25935 ( \26188 , \12847 );
or \U$25936 ( \26189 , \26187 , \26188 );
nand \U$25937 ( \26190 , \14074 , RIbe285e8_24);
nand \U$25938 ( \26191 , \26189 , \26190 );
and \U$25939 ( \26192 , \26191 , \12743 );
not \U$25940 ( \26193 , \26191 );
and \U$25941 ( \26194 , \26193 , \12746 );
nor \U$25942 ( \26195 , \26192 , \26194 );
xor \U$25943 ( \26196 , \26186 , \26195 );
not \U$25944 ( \26197 , RIbe28b10_35);
not \U$25945 ( \26198 , \13003 );
or \U$25946 ( \26199 , \26197 , \26198 );
nand \U$25947 ( \26200 , RIbe28b88_36, RIbe2ae38_110);
nand \U$25948 ( \26201 , \26199 , \26200 );
xnor \U$25949 ( \26202 , \26201 , RIbe2aeb0_111);
not \U$25950 ( \26203 , RIbe28408_20);
not \U$25951 ( \26204 , \15249 );
or \U$25952 ( \26205 , \26203 , \26204 );
nand \U$25953 ( \26206 , \12794 , RIbe28390_19);
nand \U$25954 ( \26207 , \26205 , \26206 );
not \U$25955 ( \26208 , \26207 );
not \U$25956 ( \26209 , \12801 );
and \U$25957 ( \26210 , \26208 , \26209 );
and \U$25958 ( \26211 , \26207 , \12998 );
nor \U$25959 ( \26212 , \26210 , \26211 );
xor \U$25960 ( \26213 , \26202 , \26212 );
not \U$25961 ( \26214 , RIbe287c8_28);
not \U$25962 ( \26215 , \13590 );
or \U$25963 ( \26216 , \26214 , \26215 );
nand \U$25964 ( \26217 , \21679 , RIbe28480_21);
nand \U$25965 ( \26218 , \26216 , \26217 );
not \U$25966 ( \26219 , \26218 );
not \U$25967 ( \26220 , \13706 );
and \U$25968 ( \26221 , \26219 , \26220 );
and \U$25969 ( \26222 , \26218 , \12823 );
nor \U$25970 ( \26223 , \26221 , \26222 );
xor \U$25971 ( \26224 , \26213 , \26223 );
and \U$25972 ( \26225 , \26196 , \26224 );
not \U$25973 ( \26226 , \26196 );
not \U$25974 ( \26227 , \26224 );
and \U$25975 ( \26228 , \26226 , \26227 );
or \U$25976 ( \26229 , \26225 , \26228 );
not \U$25977 ( \26230 , \26229 );
and \U$25978 ( \26231 , \26166 , \26230 );
not \U$25979 ( \26232 , \26166 );
and \U$25980 ( \26233 , \26232 , \26229 );
nor \U$25981 ( \26234 , \26231 , \26233 );
xor \U$25982 ( \26235 , \26162 , \26234 );
xor \U$25983 ( \26236 , \26070 , \26235 );
not \U$25984 ( \26237 , \25676 );
nand \U$25985 ( \26238 , \25661 , \3275 );
not \U$25986 ( \26239 , \26238 );
or \U$25987 ( \26240 , \26237 , \26239 );
nand \U$25988 ( \26241 , \25662 , \7457 );
nand \U$25989 ( \26242 , \26240 , \26241 );
or \U$25990 ( \26243 , \25797 , \25786 );
nand \U$25991 ( \26244 , \26243 , \25782 );
nand \U$25992 ( \26245 , \25797 , \25786 );
nand \U$25993 ( \26246 , \26244 , \26245 );
xor \U$25994 ( \26247 , \26242 , \26246 );
or \U$25995 ( \26248 , \25895 , \25906 );
nand \U$25996 ( \26249 , \26248 , \25915 );
nand \U$25997 ( \26250 , \25906 , \25895 );
nand \U$25998 ( \26251 , \26249 , \26250 );
xor \U$25999 ( \26252 , \26247 , \26251 );
not \U$26000 ( \26253 , \26252 );
nand \U$26001 ( \26254 , \25733 , \25757 );
and \U$26002 ( \26255 , \26254 , \25743 );
nor \U$26003 ( \26256 , \25733 , \25757 );
nor \U$26004 ( \26257 , \26255 , \26256 );
not \U$26005 ( \26258 , \26257 );
not \U$26006 ( \26259 , \26258 );
not \U$26007 ( \26260 , \25810 );
not \U$26008 ( \26261 , \25824 );
or \U$26009 ( \26262 , \26260 , \26261 );
nand \U$26010 ( \26263 , \26262 , \25836 );
nand \U$26011 ( \26264 , \25820 , \25823 );
nand \U$26012 ( \26265 , \26263 , \26264 );
not \U$26013 ( \26266 , \26265 );
not \U$26014 ( \26267 , \26266 );
or \U$26015 ( \26268 , \26259 , \26267 );
nand \U$26016 ( \26269 , \26265 , \26257 );
nand \U$26017 ( \26270 , \26268 , \26269 );
not \U$26018 ( \26271 , \26270 );
not \U$26019 ( \26272 , \25862 );
or \U$26020 ( \26273 , \26272 , \25852 );
nand \U$26021 ( \26274 , \26273 , \25875 );
nand \U$26022 ( \26275 , \26272 , \25852 );
nand \U$26023 ( \26276 , \26274 , \26275 );
not \U$26024 ( \26277 , \26276 );
not \U$26025 ( \26278 , \26277 );
and \U$26026 ( \26279 , \26271 , \26278 );
and \U$26027 ( \26280 , \26270 , \26277 );
nor \U$26028 ( \26281 , \26279 , \26280 );
not \U$26029 ( \26282 , \26281 );
or \U$26030 ( \26283 , \26253 , \26282 );
or \U$26031 ( \26284 , \26281 , \26252 );
nand \U$26032 ( \26285 , \26283 , \26284 );
nand \U$26033 ( \26286 , \25705 , \25718 );
and \U$26034 ( \26287 , \26286 , \25694 );
nor \U$26035 ( \26288 , \25705 , \25718 );
nor \U$26036 ( \26289 , \26287 , \26288 );
not \U$26037 ( \26290 , RIbe2b270_119);
not \U$26038 ( \26291 , \4829 );
or \U$26039 ( \26292 , \26290 , \26291 );
nand \U$26040 ( \26293 , RIbe2b108_116, \5731 );
nand \U$26041 ( \26294 , \26292 , \26293 );
and \U$26042 ( \26295 , \26294 , \4586 );
not \U$26043 ( \26296 , \26294 );
and \U$26044 ( \26297 , \26296 , \4946 );
nor \U$26045 ( \26298 , \26295 , \26297 );
not \U$26046 ( \26299 , RIbe2b090_115);
not \U$26047 ( \26300 , \5455 );
or \U$26048 ( \26301 , \26299 , \26300 );
nand \U$26049 ( \26302 , \7100 , RIbe2a280_85);
nand \U$26050 ( \26303 , \26301 , \26302 );
and \U$26051 ( \26304 , \26303 , \25259 );
not \U$26052 ( \26305 , \26303 );
and \U$26053 ( \26306 , \26305 , \6641 );
nor \U$26054 ( \26307 , \26304 , \26306 );
xor \U$26055 ( \26308 , \26298 , \26307 );
not \U$26056 ( \26309 , RIbe2b1f8_118);
not \U$26057 ( \26310 , \4595 );
or \U$26058 ( \26311 , \26309 , \26310 );
nand \U$26059 ( \26312 , \4600 , RIbe2b180_117);
nand \U$26060 ( \26313 , \26311 , \26312 );
and \U$26061 ( \26314 , \26313 , \4603 );
not \U$26062 ( \26315 , \26313 );
and \U$26063 ( \26316 , \26315 , \7865 );
nor \U$26064 ( \26317 , \26314 , \26316 );
xnor \U$26065 ( \26318 , \26308 , \26317 );
xor \U$26066 ( \26319 , \26289 , \26318 );
not \U$26067 ( \26320 , RIbe2afa0_113);
not \U$26068 ( \26321 , \4021 );
or \U$26069 ( \26322 , \26320 , \26321 );
nand \U$26070 ( \26323 , \4027 , RIbe2af28_112);
nand \U$26071 ( \26324 , \26322 , \26323 );
and \U$26072 ( \26325 , \26324 , \3448 );
not \U$26073 ( \26326 , \26324 );
and \U$26074 ( \26327 , \26326 , \3471 );
nor \U$26075 ( \26328 , \26325 , \26327 );
not \U$26076 ( \26329 , RIbe2b630_127);
not \U$26077 ( \26330 , \3452 );
or \U$26078 ( \26331 , \26329 , \26330 );
nand \U$26079 ( \26332 , \3458 , RIbe2b018_114);
nand \U$26080 ( \26333 , \26331 , \26332 );
and \U$26081 ( \26334 , \26333 , \4346 );
not \U$26082 ( \26335 , \26333 );
and \U$26083 ( \26336 , \26335 , \3461 );
nor \U$26084 ( \26337 , \26334 , \26336 );
xor \U$26085 ( \26338 , \26328 , \26337 );
not \U$26086 ( \26339 , RIbe2ab68_104);
not \U$26087 ( \26340 , \4050 );
or \U$26088 ( \26341 , \26339 , \26340 );
nand \U$26089 ( \26342 , \2901 , RIbe2aaf0_103);
nand \U$26090 ( \26343 , \26341 , \26342 );
and \U$26091 ( \26344 , \26343 , \7457 );
not \U$26092 ( \26345 , \26343 );
and \U$26093 ( \26346 , \26345 , \3275 );
nor \U$26094 ( \26347 , \26344 , \26346 );
xor \U$26095 ( \26348 , \26338 , \26347 );
xor \U$26096 ( \26349 , \26319 , \26348 );
not \U$26097 ( \26350 , \26349 );
and \U$26098 ( \26351 , \26285 , \26350 );
not \U$26099 ( \26352 , \26285 );
and \U$26100 ( \26353 , \26352 , \26349 );
nor \U$26101 ( \26354 , \26351 , \26353 );
xor \U$26102 ( \26355 , \26236 , \26354 );
nand \U$26103 ( \26356 , \26053 , \26045 );
nand \U$26104 ( \26357 , \26355 , \26356 );
nand \U$26105 ( \26358 , \26056 , \26357 );
xor \U$26106 ( \26359 , \26289 , \26318 );
and \U$26107 ( \26360 , \26359 , \26348 );
and \U$26108 ( \26361 , \26289 , \26318 );
or \U$26109 ( \26362 , \26360 , \26361 );
xor \U$26110 ( \26363 , \26242 , \26246 );
and \U$26111 ( \26364 , \26363 , \26251 );
and \U$26112 ( \26365 , \26242 , \26246 );
or \U$26113 ( \26366 , \26364 , \26365 );
not \U$26114 ( \26367 , \26257 );
not \U$26115 ( \26368 , \26266 );
or \U$26116 ( \26369 , \26367 , \26368 );
nand \U$26117 ( \26370 , \26369 , \26276 );
nand \U$26118 ( \26371 , \26265 , \26258 );
nand \U$26119 ( \26372 , \26370 , \26371 );
xor \U$26120 ( \26373 , \26366 , \26372 );
xnor \U$26121 ( \26374 , \26362 , \26373 );
not \U$26122 ( \26375 , \25655 );
not \U$26123 ( \26376 , \26375 );
not \U$26124 ( \26377 , \25929 );
or \U$26125 ( \26378 , \26376 , \26377 );
nand \U$26126 ( \26379 , \26378 , \25885 );
not \U$26127 ( \26380 , \25929 );
nand \U$26128 ( \26381 , \26380 , \25655 );
nand \U$26129 ( \26382 , \26379 , \26381 );
xor \U$26130 ( \26383 , \26374 , \26382 );
xor \U$26131 ( \26384 , \26070 , \26235 );
and \U$26132 ( \26385 , \26384 , \26354 );
and \U$26133 ( \26386 , \26070 , \26235 );
or \U$26134 ( \26387 , \26385 , \26386 );
xor \U$26135 ( \26388 , \26383 , \26387 );
xor \U$26136 ( \26389 , \26358 , \26388 );
xor \U$26137 ( \26390 , \26060 , \26064 );
and \U$26138 ( \26391 , \26390 , \26069 );
and \U$26139 ( \26392 , \26060 , \26064 );
or \U$26140 ( \26393 , \26391 , \26392 );
not \U$26141 ( \26394 , \26230 );
not \U$26142 ( \26395 , \26166 );
or \U$26143 ( \26396 , \26394 , \26395 );
nand \U$26144 ( \26397 , \26396 , \26162 );
not \U$26145 ( \26398 , \26166 );
nand \U$26146 ( \26399 , \26398 , \26229 );
nand \U$26147 ( \26400 , \26397 , \26399 );
xor \U$26148 ( \26401 , \26393 , \26400 );
not \U$26149 ( \26402 , \26252 );
not \U$26150 ( \26403 , \26350 );
or \U$26151 ( \26404 , \26402 , \26403 );
not \U$26152 ( \26405 , \26281 );
not \U$26153 ( \26406 , \26252 );
nand \U$26154 ( \26407 , \26406 , \26349 );
nand \U$26155 ( \26408 , \26405 , \26407 );
nand \U$26156 ( \26409 , \26404 , \26408 );
xor \U$26157 ( \26410 , \26401 , \26409 );
xor \U$26158 ( \26411 , \26202 , \26212 );
and \U$26159 ( \26412 , \26411 , \26223 );
and \U$26160 ( \26413 , \26202 , \26212 );
or \U$26161 ( \26414 , \26412 , \26413 );
xor \U$26162 ( \26415 , \26109 , \26119 );
and \U$26163 ( \26416 , \26415 , \26130 );
and \U$26164 ( \26417 , \26109 , \26119 );
or \U$26165 ( \26418 , \26416 , \26417 );
not \U$26166 ( \26419 , \26418 );
xor \U$26167 ( \26420 , \26414 , \26419 );
xor \U$26168 ( \26421 , \26176 , \26185 );
and \U$26169 ( \26422 , \26421 , \26195 );
and \U$26170 ( \26423 , \26176 , \26185 );
or \U$26171 ( \26424 , \26422 , \26423 );
not \U$26172 ( \26425 , \26424 );
xor \U$26173 ( \26426 , \26420 , \26425 );
not \U$26174 ( \26427 , RIbe28b88_36);
not \U$26175 ( \26428 , \13003 );
or \U$26176 ( \26429 , \26427 , \26428 );
nand \U$26177 ( \26430 , RIbe29290_51, RIbe2ae38_110);
nand \U$26178 ( \26431 , \26429 , \26430 );
xnor \U$26179 ( \26432 , \26431 , RIbe2aeb0_111);
xor \U$26180 ( \26433 , \1076 , \26432 );
not \U$26181 ( \26434 , RIbe28390_19);
not \U$26182 ( \26435 , \12786 );
or \U$26183 ( \26436 , \26434 , \26435 );
nand \U$26184 ( \26437 , \12794 , RIbe28b10_35);
nand \U$26185 ( \26438 , \26436 , \26437 );
and \U$26186 ( \26439 , \26438 , \12801 );
not \U$26187 ( \26440 , \26438 );
and \U$26188 ( \26441 , \26440 , \12804 );
nor \U$26189 ( \26442 , \26439 , \26441 );
xor \U$26190 ( \26443 , \26433 , \26442 );
not \U$26191 ( \26444 , \15263 );
not \U$26192 ( \26445 , RIbe28480_21);
not \U$26193 ( \26446 , \12858 );
or \U$26194 ( \26447 , \26445 , \26446 );
nand \U$26195 ( \26448 , \12835 , RIbe28408_20);
nand \U$26196 ( \26449 , \26447 , \26448 );
not \U$26197 ( \26450 , \26449 );
or \U$26198 ( \26451 , \26444 , \26450 );
or \U$26199 ( \26452 , \26449 , \12863 );
nand \U$26200 ( \26453 , \26451 , \26452 );
not \U$26201 ( \26454 , RIbe285e8_24);
not \U$26202 ( \26455 , \15161 );
or \U$26203 ( \26456 , \26454 , \26455 );
nand \U$26204 ( \26457 , \12735 , RIbe287c8_28);
nand \U$26205 ( \26458 , \26456 , \26457 );
not \U$26206 ( \26459 , \26458 );
not \U$26207 ( \26460 , \12746 );
and \U$26208 ( \26461 , \26459 , \26460 );
and \U$26209 ( \26462 , \26458 , \15169 );
nor \U$26210 ( \26463 , \26461 , \26462 );
xor \U$26211 ( \26464 , \26453 , \26463 );
not \U$26212 ( \26465 , RIbe27e68_8);
not \U$26213 ( \26466 , \14523 );
or \U$26214 ( \26467 , \26465 , \26466 );
nand \U$26215 ( \26468 , \13728 , RIbe28660_25);
nand \U$26216 ( \26469 , \26467 , \26468 );
and \U$26217 ( \26470 , \26469 , \12716 );
not \U$26218 ( \26471 , \26469 );
and \U$26219 ( \26472 , \26471 , \12723 );
nor \U$26220 ( \26473 , \26470 , \26472 );
xor \U$26221 ( \26474 , \26464 , \26473 );
xor \U$26222 ( \26475 , \26443 , \26474 );
not \U$26223 ( \26476 , RIbe27fd0_11);
not \U$26224 ( \26477 , \14725 );
or \U$26225 ( \26478 , \26476 , \26477 );
nand \U$26226 ( \26479 , \13086 , RIbe27f58_10);
nand \U$26227 ( \26480 , \26478 , \26479 );
not \U$26228 ( \26481 , \26480 );
not \U$26229 ( \26482 , \12769 );
and \U$26230 ( \26483 , \26481 , \26482 );
and \U$26231 ( \26484 , \26480 , \12924 );
nor \U$26232 ( \26485 , \26483 , \26484 );
not \U$26233 ( \26486 , RIbe28f48_44);
not \U$26234 ( \26487 , \12943 );
or \U$26235 ( \26488 , \26486 , \26487 );
nand \U$26236 ( \26489 , \13669 , RIbe28ed0_43);
nand \U$26237 ( \26490 , \26488 , \26489 );
and \U$26238 ( \26491 , \26490 , \12195 );
not \U$26239 ( \26492 , \26490 );
and \U$26240 ( \26493 , \26492 , \12960 );
nor \U$26241 ( \26494 , \26491 , \26493 );
xor \U$26242 ( \26495 , \26485 , \26494 );
not \U$26243 ( \26496 , RIbe29c68_72);
not \U$26244 ( \26497 , \10936 );
or \U$26245 ( \26498 , \26496 , \26497 );
nand \U$26246 ( \26499 , \12213 , RIbe29bf0_71);
nand \U$26247 ( \26500 , \26498 , \26499 );
and \U$26248 ( \26501 , \26500 , \9903 );
not \U$26249 ( \26502 , \26500 );
and \U$26250 ( \26503 , \26502 , \19139 );
nor \U$26251 ( \26504 , \26501 , \26503 );
xnor \U$26252 ( \26505 , \26495 , \26504 );
xor \U$26253 ( \26506 , \26475 , \26505 );
xor \U$26254 ( \26507 , \26426 , \26506 );
nand \U$26255 ( \26508 , \26227 , \26196 );
not \U$26256 ( \26509 , \26508 );
not \U$26257 ( \26510 , \26102 );
and \U$26258 ( \26511 , \26161 , \26510 );
nor \U$26259 ( \26512 , \26511 , \26131 );
nor \U$26260 ( \26513 , \26161 , \26510 );
nor \U$26261 ( \26514 , \26512 , \26513 );
not \U$26262 ( \26515 , \26514 );
not \U$26263 ( \26516 , \26515 );
or \U$26264 ( \26517 , \26509 , \26516 );
not \U$26265 ( \26518 , \26508 );
nand \U$26266 ( \26519 , \26514 , \26518 );
nand \U$26267 ( \26520 , \26517 , \26519 );
xnor \U$26268 ( \26521 , \26507 , \26520 );
xor \U$26269 ( \26522 , \26142 , \26149 );
and \U$26270 ( \26523 , \26522 , \26160 );
and \U$26271 ( \26524 , \26142 , \26149 );
or \U$26272 ( \26525 , \26523 , \26524 );
not \U$26273 ( \26526 , \26525 );
or \U$26274 ( \26527 , \26317 , \26298 );
nand \U$26275 ( \26528 , \26527 , \26307 );
nand \U$26276 ( \26529 , \26317 , \26298 );
nand \U$26277 ( \26530 , \26528 , \26529 );
xor \U$26278 ( \26531 , \26081 , \26091 );
and \U$26279 ( \26532 , \26531 , \26101 );
and \U$26280 ( \26533 , \26081 , \26091 );
or \U$26281 ( \26534 , \26532 , \26533 );
xor \U$26282 ( \26535 , \26530 , \26534 );
not \U$26283 ( \26536 , \26535 );
or \U$26284 ( \26537 , \26526 , \26536 );
or \U$26285 ( \26538 , \26535 , \26525 );
nand \U$26286 ( \26539 , \26537 , \26538 );
not \U$26287 ( \26540 , RIbe2af28_112);
not \U$26288 ( \26541 , \7880 );
or \U$26289 ( \26542 , \26540 , \26541 );
nand \U$26290 ( \26543 , \4332 , RIbe2b1f8_118);
nand \U$26291 ( \26544 , \26542 , \26543 );
and \U$26292 ( \26545 , \26544 , \3448 );
not \U$26293 ( \26546 , \26544 );
and \U$26294 ( \26547 , \26546 , \3471 );
nor \U$26295 ( \26548 , \26545 , \26547 );
not \U$26296 ( \26549 , RIbe2b180_117);
not \U$26297 ( \26550 , \5058 );
or \U$26298 ( \26551 , \26549 , \26550 );
nand \U$26299 ( \26552 , \4600 , RIbe2b270_119);
nand \U$26300 ( \26553 , \26551 , \26552 );
and \U$26301 ( \26554 , \26553 , \4326 );
not \U$26302 ( \26555 , \26553 );
and \U$26303 ( \26556 , \26555 , \4323 );
nor \U$26304 ( \26557 , \26554 , \26556 );
and \U$26305 ( \26558 , \26548 , \26557 );
not \U$26306 ( \26559 , \26548 );
not \U$26307 ( \26560 , \26557 );
and \U$26308 ( \26561 , \26559 , \26560 );
or \U$26309 ( \26562 , \26558 , \26561 );
not \U$26310 ( \26563 , RIbe2b018_114);
not \U$26311 ( \26564 , \4764 );
or \U$26312 ( \26565 , \26563 , \26564 );
nand \U$26313 ( \26566 , \4011 , RIbe2afa0_113);
nand \U$26314 ( \26567 , \26565 , \26566 );
and \U$26315 ( \26568 , \26567 , \2887 );
not \U$26316 ( \26569 , \26567 );
and \U$26317 ( \26570 , \26569 , \4346 );
nor \U$26318 ( \26571 , \26568 , \26570 );
xnor \U$26319 ( \26572 , \26562 , \26571 );
not \U$26320 ( \26573 , \26328 );
or \U$26321 ( \26574 , \26573 , \26347 );
nand \U$26322 ( \26575 , \26574 , \26337 );
nand \U$26323 ( \26576 , \26573 , \26347 );
nand \U$26324 ( \26577 , \26575 , \26576 );
not \U$26325 ( \26578 , RIbe2aaf0_103);
not \U$26326 ( \26579 , \2898 );
or \U$26327 ( \26580 , \26578 , \26579 );
nand \U$26328 ( \26581 , \2901 , RIbe2b630_127);
nand \U$26329 ( \26582 , \26580 , \26581 );
and \U$26330 ( \26583 , \26582 , \2573 );
not \U$26331 ( \26584 , \26582 );
and \U$26332 ( \26585 , \26584 , \3275 );
nor \U$26333 ( \26586 , \26583 , \26585 );
not \U$26334 ( \26587 , \4065 );
nand \U$26335 ( \26588 , \26587 , RIbe2ab68_104);
not \U$26336 ( \26589 , \26588 );
not \U$26337 ( \26590 , \1274 );
and \U$26338 ( \26591 , \26589 , \26590 );
and \U$26339 ( \26592 , \26588 , \1277 );
nor \U$26340 ( \26593 , \26591 , \26592 );
and \U$26341 ( \26594 , \26586 , \26593 );
not \U$26342 ( \26595 , \26586 );
not \U$26343 ( \26596 , \26593 );
and \U$26344 ( \26597 , \26595 , \26596 );
or \U$26345 ( \26598 , \26594 , \26597 );
xor \U$26346 ( \26599 , \26577 , \26598 );
xor \U$26347 ( \26600 , \26572 , \26599 );
xor \U$26348 ( \26601 , \26539 , \26600 );
and \U$26349 ( \26602 , \20405 , RIbe29e48_76);
and \U$26350 ( \26603 , \13038 , RIbe29dd0_75);
nor \U$26351 ( \26604 , \26602 , \26603 );
and \U$26352 ( \26605 , \26604 , \25808 );
not \U$26353 ( \26606 , \26604 );
and \U$26354 ( \26607 , \26606 , \7970 );
nor \U$26355 ( \26608 , \26605 , \26607 );
not \U$26356 ( \26609 , RIbe2a028_80);
not \U$26357 ( \26610 , \6942 );
or \U$26358 ( \26611 , \26609 , \26610 );
nand \U$26359 ( \26612 , \7981 , RIbe29fb0_79);
nand \U$26360 ( \26613 , \26611 , \26612 );
not \U$26361 ( \26614 , \26613 );
not \U$26362 ( \26615 , \7984 );
and \U$26363 ( \26616 , \26614 , \26615 );
and \U$26364 ( \26617 , \26613 , \7989 );
nor \U$26365 ( \26618 , \26616 , \26617 );
xor \U$26366 ( \26619 , \26608 , \26618 );
not \U$26367 ( \26620 , RIbe2a2f8_86);
not \U$26368 ( \26621 , \13171 );
or \U$26369 ( \26622 , \26620 , \26621 );
nand \U$26370 ( \26623 , \9875 , RIbe2acd0_107);
nand \U$26371 ( \26624 , \26622 , \26623 );
and \U$26372 ( \26625 , \26624 , \13227 );
not \U$26373 ( \26626 , \26624 );
and \U$26374 ( \26627 , \26626 , \14650 );
nor \U$26375 ( \26628 , \26625 , \26627 );
xor \U$26376 ( \26629 , \26619 , \26628 );
not \U$26377 ( \26630 , \5740 );
not \U$26378 ( \26631 , RIbe2a190_83);
not \U$26379 ( \26632 , \13894 );
or \U$26380 ( \26633 , \26631 , \26632 );
nand \U$26381 ( \26634 , \6616 , RIbe2a5c8_92);
nand \U$26382 ( \26635 , \26633 , \26634 );
not \U$26383 ( \26636 , \26635 );
or \U$26384 ( \26637 , \26630 , \26636 );
or \U$26385 ( \26638 , \26635 , \10972 );
nand \U$26386 ( \26639 , \26637 , \26638 );
not \U$26387 ( \26640 , \26639 );
not \U$26388 ( \26641 , RIbe2a280_85);
not \U$26389 ( \26642 , \15313 );
or \U$26390 ( \26643 , \26641 , \26642 );
nand \U$26391 ( \26644 , \15885 , RIbe2a208_84);
nand \U$26392 ( \26645 , \26643 , \26644 );
not \U$26393 ( \26646 , \26645 );
not \U$26394 ( \26647 , \5046 );
and \U$26395 ( \26648 , \26646 , \26647 );
and \U$26396 ( \26649 , \26645 , \6637 );
nor \U$26397 ( \26650 , \26648 , \26649 );
not \U$26398 ( \26651 , \26650 );
or \U$26399 ( \26652 , \26640 , \26651 );
or \U$26400 ( \26653 , \26650 , \26639 );
nand \U$26401 ( \26654 , \26652 , \26653 );
not \U$26402 ( \26655 , RIbe2b108_116);
not \U$26403 ( \26656 , \5727 );
or \U$26404 ( \26657 , \26655 , \26656 );
nand \U$26405 ( \26658 , \7056 , RIbe2b090_115);
nand \U$26406 ( \26659 , \26657 , \26658 );
and \U$26407 ( \26660 , \26659 , \4946 );
not \U$26408 ( \26661 , \26659 );
and \U$26409 ( \26662 , \26661 , \4586 );
nor \U$26410 ( \26663 , \26660 , \26662 );
not \U$26411 ( \26664 , \26663 );
and \U$26412 ( \26665 , \26654 , \26664 );
not \U$26413 ( \26666 , \26654 );
and \U$26414 ( \26667 , \26666 , \26663 );
nor \U$26415 ( \26668 , \26665 , \26667 );
xor \U$26416 ( \26669 , \26629 , \26668 );
not \U$26417 ( \26670 , RIbe2a910_99);
not \U$26418 ( \26671 , \6591 );
or \U$26419 ( \26672 , \26670 , \26671 );
nand \U$26420 ( \26673 , \7278 , RIbe2b5b8_126);
nand \U$26421 ( \26674 , \26672 , \26673 );
not \U$26422 ( \26675 , \26674 );
not \U$26423 ( \26676 , \8957 );
and \U$26424 ( \26677 , \26675 , \26676 );
and \U$26425 ( \26678 , \26674 , \7488 );
nor \U$26426 ( \26679 , \26677 , \26678 );
not \U$26427 ( \26680 , \26679 );
not \U$26428 ( \26681 , RIbe2a3e8_88);
not \U$26429 ( \26682 , \6958 );
or \U$26430 ( \26683 , \26681 , \26682 );
nand \U$26431 ( \26684 , \8202 , RIbe2a370_87);
nand \U$26432 ( \26685 , \26683 , \26684 );
and \U$26433 ( \26686 , \26685 , \7293 );
not \U$26434 ( \26687 , \26685 );
and \U$26435 ( \26688 , \26687 , \6572 );
nor \U$26436 ( \26689 , \26686 , \26688 );
not \U$26437 ( \26690 , \26689 );
or \U$26438 ( \26691 , \26680 , \26690 );
or \U$26439 ( \26692 , \26679 , \26689 );
nand \U$26440 ( \26693 , \26691 , \26692 );
not \U$26441 ( \26694 , RIbe2a550_91);
not \U$26442 ( \26695 , \6536 );
or \U$26443 ( \26696 , \26694 , \26695 );
nand \U$26444 ( \26697 , \6540 , RIbe2a988_100);
nand \U$26445 ( \26698 , \26696 , \26697 );
and \U$26446 ( \26699 , \26698 , \6546 );
not \U$26447 ( \26700 , \26698 );
and \U$26448 ( \26701 , \26700 , \6891 );
nor \U$26449 ( \26702 , \26699 , \26701 );
not \U$26450 ( \26703 , \26702 );
and \U$26451 ( \26704 , \26693 , \26703 );
not \U$26452 ( \26705 , \26693 );
and \U$26453 ( \26706 , \26705 , \26702 );
nor \U$26454 ( \26707 , \26704 , \26706 );
xor \U$26455 ( \26708 , \26669 , \26707 );
xnor \U$26456 ( \26709 , \26601 , \26708 );
not \U$26457 ( \26710 , \26709 );
and \U$26458 ( \26711 , \26521 , \26710 );
not \U$26459 ( \26712 , \26521 );
and \U$26460 ( \26713 , \26712 , \26709 );
nor \U$26461 ( \26714 , \26711 , \26713 );
xor \U$26462 ( \26715 , \26410 , \26714 );
xor \U$26463 ( \26716 , \26389 , \26715 );
nand \U$26464 ( \26717 , \26040 , \26716 );
not \U$26465 ( \26718 , \26717 );
xor \U$26466 ( \26719 , \26443 , \26474 );
and \U$26467 ( \26720 , \26719 , \26505 );
and \U$26468 ( \26721 , \26443 , \26474 );
or \U$26469 ( \26722 , \26720 , \26721 );
nand \U$26470 ( \26723 , \26629 , \26707 );
and \U$26471 ( \26724 , \26723 , \26668 );
nor \U$26472 ( \26725 , \26629 , \26707 );
nor \U$26473 ( \26726 , \26724 , \26725 );
xor \U$26474 ( \26727 , \26722 , \26726 );
xnor \U$26475 ( \26728 , \25355 , \25361 );
not \U$26476 ( \26729 , \26728 );
not \U$26477 ( \26730 , \25372 );
and \U$26478 ( \26731 , \26729 , \26730 );
and \U$26479 ( \26732 , \26728 , \25372 );
nor \U$26480 ( \26733 , \26731 , \26732 );
xnor \U$26481 ( \26734 , \26727 , \26733 );
xor \U$26482 ( \26735 , \26393 , \26400 );
and \U$26483 ( \26736 , \26735 , \26409 );
and \U$26484 ( \26737 , \26393 , \26400 );
or \U$26485 ( \26738 , \26736 , \26737 );
xor \U$26486 ( \26739 , \26734 , \26738 );
not \U$26487 ( \26740 , \26426 );
not \U$26488 ( \26741 , \26710 );
or \U$26489 ( \26742 , \26740 , \26741 );
not \U$26490 ( \26743 , \26426 );
not \U$26491 ( \26744 , \26743 );
not \U$26492 ( \26745 , \26709 );
or \U$26493 ( \26746 , \26744 , \26745 );
xnor \U$26494 ( \26747 , \26506 , \26520 );
nand \U$26495 ( \26748 , \26746 , \26747 );
nand \U$26496 ( \26749 , \26742 , \26748 );
xor \U$26497 ( \26750 , \26739 , \26749 );
xor \U$26498 ( \26751 , \26358 , \26388 );
and \U$26499 ( \26752 , \26751 , \26715 );
and \U$26500 ( \26753 , \26358 , \26388 );
or \U$26501 ( \26754 , \26752 , \26753 );
xor \U$26502 ( \26755 , \26750 , \26754 );
or \U$26503 ( \26756 , \26577 , \26598 );
and \U$26504 ( \26757 , \26756 , \26572 );
and \U$26505 ( \26758 , \26577 , \26598 );
nor \U$26506 ( \26759 , \26757 , \26758 );
not \U$26507 ( \26760 , \26759 );
or \U$26508 ( \26761 , \26534 , \26530 );
not \U$26509 ( \26762 , \26525 );
and \U$26510 ( \26763 , \26761 , \26762 );
and \U$26511 ( \26764 , \26530 , \26534 );
nor \U$26512 ( \26765 , \26763 , \26764 );
nand \U$26513 ( \26766 , \26418 , \26414 );
and \U$26514 ( \26767 , \26766 , \26424 );
nor \U$26515 ( \26768 , \26418 , \26414 );
nor \U$26516 ( \26769 , \26767 , \26768 );
xor \U$26517 ( \26770 , \26765 , \26769 );
not \U$26518 ( \26771 , \26770 );
or \U$26519 ( \26772 , \26760 , \26771 );
or \U$26520 ( \26773 , \26770 , \26759 );
nand \U$26521 ( \26774 , \26772 , \26773 );
not \U$26522 ( \26775 , \26463 );
or \U$26523 ( \26776 , \26473 , \26775 );
nand \U$26524 ( \26777 , \26776 , \26453 );
nand \U$26525 ( \26778 , \26473 , \26775 );
nand \U$26526 ( \26779 , \26777 , \26778 );
not \U$26527 ( \26780 , \26779 );
nand \U$26528 ( \26781 , \26504 , \26485 );
and \U$26529 ( \26782 , \26781 , \26494 );
nor \U$26530 ( \26783 , \26504 , \26485 );
nor \U$26531 ( \26784 , \26782 , \26783 );
xor \U$26532 ( \26785 , \1076 , \26432 );
and \U$26533 ( \26786 , \26785 , \26442 );
and \U$26534 ( \26787 , \1076 , \26432 );
or \U$26535 ( \26788 , \26786 , \26787 );
not \U$26536 ( \26789 , \26788 );
and \U$26537 ( \26790 , \26784 , \26789 );
not \U$26538 ( \26791 , \26784 );
and \U$26539 ( \26792 , \26791 , \26788 );
nor \U$26540 ( \26793 , \26790 , \26792 );
not \U$26541 ( \26794 , \26793 );
or \U$26542 ( \26795 , \26780 , \26794 );
or \U$26543 ( \26796 , \26793 , \26779 );
nand \U$26544 ( \26797 , \26795 , \26796 );
not \U$26545 ( \26798 , \26679 );
or \U$26546 ( \26799 , \26798 , \26689 );
nand \U$26547 ( \26800 , \26799 , \26702 );
nand \U$26548 ( \26801 , \26689 , \26798 );
nand \U$26549 ( \26802 , \26800 , \26801 );
not \U$26550 ( \26803 , \26664 );
not \U$26551 ( \26804 , \26650 );
not \U$26552 ( \26805 , \26804 );
or \U$26553 ( \26806 , \26803 , \26805 );
not \U$26554 ( \26807 , \26663 );
not \U$26555 ( \26808 , \26650 );
or \U$26556 ( \26809 , \26807 , \26808 );
nand \U$26557 ( \26810 , \26809 , \26639 );
nand \U$26558 ( \26811 , \26806 , \26810 );
xor \U$26559 ( \26812 , \26802 , \26811 );
not \U$26560 ( \26813 , \26608 );
not \U$26561 ( \26814 , \26618 );
not \U$26562 ( \26815 , \26814 );
or \U$26563 ( \26816 , \26813 , \26815 );
not \U$26564 ( \26817 , \26608 );
not \U$26565 ( \26818 , \26817 );
not \U$26566 ( \26819 , \26618 );
or \U$26567 ( \26820 , \26818 , \26819 );
nand \U$26568 ( \26821 , \26820 , \26628 );
nand \U$26569 ( \26822 , \26816 , \26821 );
xor \U$26570 ( \26823 , \26812 , \26822 );
xor \U$26571 ( \26824 , \26797 , \26823 );
not \U$26572 ( \26825 , \2889 );
not \U$26573 ( \26826 , \13192 );
and \U$26574 ( \26827 , \26825 , \26826 );
and \U$26575 ( \26828 , \2583 , RIbe2ab68_104);
nor \U$26576 ( \26829 , \26827 , \26828 );
and \U$26577 ( \26830 , \26829 , \7038 );
not \U$26578 ( \26831 , \26829 );
and \U$26579 ( \26832 , \26831 , \1277 );
nor \U$26580 ( \26833 , \26830 , \26832 );
nand \U$26581 ( \26834 , \26596 , \26586 );
xor \U$26582 ( \26835 , \26833 , \26834 );
and \U$26583 ( \26836 , \26571 , \26548 );
nor \U$26584 ( \26837 , \26836 , \26560 );
nor \U$26585 ( \26838 , \26571 , \26548 );
nor \U$26586 ( \26839 , \26837 , \26838 );
xnor \U$26587 ( \26840 , \26835 , \26839 );
xor \U$26588 ( \26841 , \25461 , \25470 );
xor \U$26589 ( \26842 , \26841 , \25481 );
xor \U$26590 ( \26843 , \25277 , \25287 );
xor \U$26591 ( \26844 , \26843 , \25297 );
xor \U$26592 ( \26845 , \26842 , \26844 );
xor \U$26593 ( \26846 , \25251 , \25263 );
xnor \U$26594 ( \26847 , \26846 , \25245 );
xor \U$26595 ( \26848 , \26845 , \26847 );
xor \U$26596 ( \26849 , \26840 , \26848 );
not \U$26597 ( \26850 , \25402 );
not \U$26598 ( \26851 , \25386 );
or \U$26599 ( \26852 , \26850 , \26851 );
nand \U$26600 ( \26853 , \25401 , \25385 );
nand \U$26601 ( \26854 , \26852 , \26853 );
xor \U$26602 ( \26855 , \26854 , \25393 );
not \U$26603 ( \26856 , \25339 );
not \U$26604 ( \26857 , \25312 );
or \U$26605 ( \26858 , \26856 , \26857 );
or \U$26606 ( \26859 , \25312 , \25339 );
nand \U$26607 ( \26860 , \26858 , \26859 );
xor \U$26608 ( \26861 , \26860 , \25324 );
xor \U$26609 ( \26862 , \26855 , \26861 );
not \U$26610 ( \26863 , \25431 );
not \U$26611 ( \26864 , \25427 );
or \U$26612 ( \26865 , \26863 , \26864 );
nand \U$26613 ( \26866 , \25426 , \25416 );
nand \U$26614 ( \26867 , \26865 , \26866 );
xnor \U$26615 ( \26868 , \26867 , \25442 );
xor \U$26616 ( \26869 , \26862 , \26868 );
xnor \U$26617 ( \26870 , \26849 , \26869 );
xor \U$26618 ( \26871 , \26824 , \26870 );
xor \U$26619 ( \26872 , \26774 , \26871 );
nor \U$26620 ( \26873 , \26372 , \26366 );
or \U$26621 ( \26874 , \26362 , \26873 );
nand \U$26622 ( \26875 , \26372 , \26366 );
nand \U$26623 ( \26876 , \26874 , \26875 );
or \U$26624 ( \26877 , \26539 , \26600 );
and \U$26625 ( \26878 , \26708 , \26877 );
and \U$26626 ( \26879 , \26539 , \26600 );
nor \U$26627 ( \26880 , \26878 , \26879 );
not \U$26628 ( \26881 , \26880 );
xor \U$26629 ( \26882 , \26876 , \26881 );
not \U$26630 ( \26883 , \26508 );
not \U$26631 ( \26884 , \26506 );
or \U$26632 ( \26885 , \26883 , \26884 );
nand \U$26633 ( \26886 , \26885 , \26515 );
not \U$26634 ( \26887 , \26506 );
nand \U$26635 ( \26888 , \26887 , \26518 );
nand \U$26636 ( \26889 , \26886 , \26888 );
xor \U$26637 ( \26890 , \26882 , \26889 );
xor \U$26638 ( \26891 , \26872 , \26890 );
not \U$26639 ( \26892 , \26891 );
nand \U$26640 ( \26893 , \26714 , \26410 );
not \U$26641 ( \26894 , \26893 );
xor \U$26642 ( \26895 , \26374 , \26382 );
and \U$26643 ( \26896 , \26895 , \26387 );
and \U$26644 ( \26897 , \26374 , \26382 );
or \U$26645 ( \26898 , \26896 , \26897 );
not \U$26646 ( \26899 , \26898 );
and \U$26647 ( \26900 , \26894 , \26899 );
and \U$26648 ( \26901 , \26893 , \26898 );
nor \U$26649 ( \26902 , \26900 , \26901 );
not \U$26650 ( \26903 , \26902 );
or \U$26651 ( \26904 , \26892 , \26903 );
or \U$26652 ( \26905 , \26902 , \26891 );
nand \U$26653 ( \26906 , \26904 , \26905 );
xor \U$26654 ( \26907 , \26755 , \26906 );
not \U$26655 ( \26908 , \26907 );
or \U$26656 ( \26909 , \26718 , \26908 );
or \U$26657 ( \26910 , \26907 , \26717 );
nand \U$26658 ( \26911 , \26909 , \26910 );
buf \U$26659 ( \26912 , \26911 );
xor \U$26660 ( \26913 , \26750 , \26754 );
and \U$26661 ( \26914 , \26913 , \26906 );
and \U$26662 ( \26915 , \26750 , \26754 );
or \U$26663 ( \26916 , \26914 , \26915 );
not \U$26664 ( \26917 , \26916 );
and \U$26665 ( \26918 , \26733 , \26726 );
nor \U$26666 ( \26919 , \26918 , \26722 );
nor \U$26667 ( \26920 , \26726 , \26733 );
nor \U$26668 ( \26921 , \26919 , \26920 );
not \U$26669 ( \26922 , \26921 );
and \U$26670 ( \26923 , \26769 , \26759 );
nor \U$26671 ( \26924 , \26923 , \26765 );
nor \U$26672 ( \26925 , \26759 , \26769 );
nor \U$26673 ( \26926 , \26924 , \26925 );
not \U$26674 ( \26927 , \26926 );
and \U$26675 ( \26928 , \26922 , \26927 );
not \U$26676 ( \26929 , \26922 );
and \U$26677 ( \26930 , \26929 , \26926 );
nor \U$26678 ( \26931 , \26928 , \26930 );
not \U$26679 ( \26932 , \26848 );
nand \U$26680 ( \26933 , \26932 , \26840 );
not \U$26681 ( \26934 , \26933 );
not \U$26682 ( \26935 , \26869 );
or \U$26683 ( \26936 , \26934 , \26935 );
not \U$26684 ( \26937 , \26840 );
nand \U$26685 ( \26938 , \26937 , \26848 );
nand \U$26686 ( \26939 , \26936 , \26938 );
xor \U$26687 ( \26940 , \26931 , \26939 );
xor \U$26688 ( \26941 , \26797 , \26823 );
and \U$26689 ( \26942 , \26941 , \26870 );
and \U$26690 ( \26943 , \26797 , \26823 );
or \U$26691 ( \26944 , \26942 , \26943 );
not \U$26692 ( \26945 , \26944 );
xor \U$26693 ( \26946 , \26940 , \26945 );
not \U$26694 ( \26947 , \26822 );
not \U$26695 ( \26948 , \26811 );
or \U$26696 ( \26949 , \26947 , \26948 );
or \U$26697 ( \26950 , \26811 , \26822 );
nand \U$26698 ( \26951 , \26950 , \26802 );
nand \U$26699 ( \26952 , \26949 , \26951 );
not \U$26700 ( \26953 , \26788 );
not \U$26701 ( \26954 , \26784 );
or \U$26702 ( \26955 , \26953 , \26954 );
nand \U$26703 ( \26956 , \26955 , \26779 );
not \U$26704 ( \26957 , \26784 );
nand \U$26705 ( \26958 , \26957 , \26789 );
nand \U$26706 ( \26959 , \26956 , \26958 );
xor \U$26707 ( \26960 , \26952 , \26959 );
not \U$26708 ( \26961 , \26833 );
not \U$26709 ( \26962 , \26834 );
not \U$26710 ( \26963 , \26962 );
or \U$26711 ( \26964 , \26961 , \26963 );
not \U$26712 ( \26965 , \26839 );
not \U$26713 ( \26966 , \26833 );
nand \U$26714 ( \26967 , \26966 , \26834 );
nand \U$26715 ( \26968 , \26965 , \26967 );
nand \U$26716 ( \26969 , \26964 , \26968 );
xor \U$26717 ( \26970 , \26960 , \26969 );
not \U$26718 ( \26971 , \26970 );
not \U$26719 ( \26972 , \26876 );
not \U$26720 ( \26973 , \26881 );
or \U$26721 ( \26974 , \26972 , \26973 );
not \U$26722 ( \26975 , \26876 );
nand \U$26723 ( \26976 , \26975 , \26880 );
nand \U$26724 ( \26977 , \26976 , \26889 );
nand \U$26725 ( \26978 , \26974 , \26977 );
nor \U$26726 ( \26979 , \26971 , \26978 );
not \U$26727 ( \26980 , \26979 );
not \U$26728 ( \26981 , \26970 );
nand \U$26729 ( \26982 , \26981 , \26978 );
nand \U$26730 ( \26983 , \26980 , \26982 );
xnor \U$26731 ( \26984 , \26946 , \26983 );
not \U$26732 ( \26985 , \26984 );
not \U$26733 ( \26986 , \26985 );
xor \U$26734 ( \26987 , \25444 , \25446 );
xor \U$26735 ( \26988 , \25447 , \26987 );
xor \U$26736 ( \26989 , \25216 , \25228 );
xor \U$26737 ( \26990 , \26989 , \25207 );
not \U$26738 ( \26991 , \26990 );
xor \U$26739 ( \26992 , \26988 , \26991 );
not \U$26740 ( \26993 , \26842 );
and \U$26741 ( \26994 , \26847 , \26993 );
nor \U$26742 ( \26995 , \26994 , \26844 );
nor \U$26743 ( \26996 , \26993 , \26847 );
nor \U$26744 ( \26997 , \26995 , \26996 );
not \U$26745 ( \26998 , \26997 );
not \U$26746 ( \26999 , \26998 );
nand \U$26747 ( \27000 , \26855 , \26868 );
and \U$26748 ( \27001 , \27000 , \26861 );
nor \U$26749 ( \27002 , \26855 , \26868 );
nor \U$26750 ( \27003 , \27001 , \27002 );
not \U$26751 ( \27004 , \27003 );
or \U$26752 ( \27005 , \26999 , \27004 );
not \U$26753 ( \27006 , \27003 );
nand \U$26754 ( \27007 , \27006 , \26997 );
nand \U$26755 ( \27008 , \27005 , \27007 );
xor \U$26756 ( \27009 , \26992 , \27008 );
not \U$26757 ( \27010 , \27009 );
and \U$26758 ( \27011 , \25300 , \25344 );
not \U$26759 ( \27012 , \25300 );
and \U$26760 ( \27013 , \27012 , \25266 );
or \U$26761 ( \27014 , \27011 , \27013 );
xnor \U$26762 ( \27015 , \27014 , \25341 );
not \U$26763 ( \27016 , \27015 );
and \U$26764 ( \27017 , \25488 , \25485 );
not \U$26765 ( \27018 , \25488 );
and \U$26766 ( \27019 , \27018 , \25484 );
or \U$26767 ( \27020 , \27017 , \27019 );
xor \U$26768 ( \27021 , \27020 , \25452 );
not \U$26769 ( \27022 , \27021 );
not \U$26770 ( \27023 , \27022 );
or \U$26771 ( \27024 , \27016 , \27023 );
not \U$26772 ( \27025 , \27015 );
nand \U$26773 ( \27026 , \27025 , \27021 );
nand \U$26774 ( \27027 , \27024 , \27026 );
xor \U$26775 ( \27028 , \25181 , \25186 );
not \U$26776 ( \27029 , \25178 );
xor \U$26777 ( \27030 , \27028 , \27029 );
not \U$26778 ( \27031 , \27030 );
and \U$26779 ( \27032 , \27027 , \27031 );
not \U$26780 ( \27033 , \27027 );
and \U$26781 ( \27034 , \27033 , \27030 );
nor \U$26782 ( \27035 , \27032 , \27034 );
not \U$26783 ( \27036 , \27035 );
and \U$26784 ( \27037 , \27010 , \27036 );
and \U$26785 ( \27038 , \27009 , \27035 );
nor \U$26786 ( \27039 , \27037 , \27038 );
not \U$26787 ( \27040 , \27039 );
not \U$26788 ( \27041 , \27040 );
xor \U$26789 ( \27042 , \26734 , \26738 );
and \U$26790 ( \27043 , \27042 , \26749 );
and \U$26791 ( \27044 , \26734 , \26738 );
or \U$26792 ( \27045 , \27043 , \27044 );
not \U$26793 ( \27046 , \27045 );
not \U$26794 ( \27047 , \27046 );
or \U$26795 ( \27048 , \27041 , \27047 );
nand \U$26796 ( \27049 , \27045 , \27039 );
nand \U$26797 ( \27050 , \27048 , \27049 );
xor \U$26798 ( \27051 , \26774 , \26871 );
and \U$26799 ( \27052 , \27051 , \26890 );
and \U$26800 ( \27053 , \26774 , \26871 );
or \U$26801 ( \27054 , \27052 , \27053 );
not \U$26802 ( \27055 , \27054 );
and \U$26803 ( \27056 , \27050 , \27055 );
not \U$26804 ( \27057 , \27050 );
and \U$26805 ( \27058 , \27057 , \27054 );
nor \U$26806 ( \27059 , \27056 , \27058 );
not \U$26807 ( \27060 , \27059 );
not \U$26808 ( \27061 , \27060 );
or \U$26809 ( \27062 , \26986 , \27061 );
nand \U$26810 ( \27063 , \27059 , \26984 );
nand \U$26811 ( \27064 , \27062 , \27063 );
not \U$26812 ( \27065 , \26898 );
nand \U$26813 ( \27066 , \27065 , \26893 );
and \U$26814 ( \27067 , \26891 , \27066 );
not \U$26815 ( \27068 , \26898 );
nor \U$26816 ( \27069 , \27068 , \26893 );
nor \U$26817 ( \27070 , \27067 , \27069 );
and \U$26818 ( \27071 , \27064 , \27070 );
not \U$26819 ( \27072 , \27064 );
not \U$26820 ( \27073 , \27070 );
and \U$26821 ( \27074 , \27072 , \27073 );
nor \U$26822 ( \27075 , \27071 , \27074 );
xor \U$26823 ( \27076 , \26917 , \27075 );
buf \U$26824 ( \27077 , \27076 );
xor \U$26825 ( \27078 , \25930 , \26019 );
xor \U$26826 ( \27079 , \27078 , \26036 );
not \U$26827 ( \27080 , \27079 );
not \U$26828 ( \27081 , \27080 );
xor \U$26829 ( \27082 , \26054 , \26046 );
xor \U$26830 ( \27083 , \26355 , \27082 );
not \U$26831 ( \27084 , \27083 );
or \U$26832 ( \27085 , \27081 , \27084 );
not \U$26833 ( \27086 , \27083 );
not \U$26834 ( \27087 , \27086 );
not \U$26835 ( \27088 , \27079 );
or \U$26836 ( \27089 , \27087 , \27088 );
not \U$26837 ( \27090 , \26026 );
and \U$26838 ( \27091 , \26033 , \27090 );
not \U$26839 ( \27092 , \26033 );
and \U$26840 ( \27093 , \27092 , \26026 );
nor \U$26841 ( \27094 , \27091 , \27093 );
buf \U$26842 ( \27095 , \26024 );
not \U$26843 ( \27096 , \27095 );
and \U$26844 ( \27097 , \27094 , \27096 );
not \U$26845 ( \27098 , \27094 );
and \U$26846 ( \27099 , \27098 , \27095 );
nor \U$26847 ( \27100 , \27097 , \27099 );
not \U$26848 ( \27101 , \16516 );
not \U$26849 ( \27102 , \16853 );
or \U$26850 ( \27103 , \27101 , \27102 );
or \U$26851 ( \27104 , \16516 , \16853 );
nand \U$26852 ( \27105 , \27104 , \16520 );
nand \U$26853 ( \27106 , \27103 , \27105 );
xor \U$26854 ( \27107 , \27100 , \27106 );
xor \U$26855 ( \27108 , \25989 , \25987 );
xor \U$26856 ( \27109 , \27108 , \26016 );
and \U$26857 ( \27110 , \27107 , \27109 );
and \U$26858 ( \27111 , \27100 , \27106 );
or \U$26859 ( \27112 , \27110 , \27111 );
nand \U$26860 ( \27113 , \27089 , \27112 );
nand \U$26861 ( \27114 , \27085 , \27113 );
xnor \U$26862 ( \27115 , \26039 , \26716 );
xor \U$26863 ( \27116 , \27114 , \27115 );
buf \U$26864 ( \27117 , \27116 );
xor \U$26865 ( \27118 , \27100 , \27106 );
xor \U$26866 ( \27119 , \27118 , \27109 );
buf \U$26867 ( \27120 , \16480 );
not \U$26868 ( \27121 , \27120 );
not \U$26869 ( \27122 , \27121 );
not \U$26870 ( \27123 , \16504 );
or \U$26871 ( \27124 , \27122 , \27123 );
not \U$26872 ( \27125 , \16854 );
not \U$26873 ( \27126 , \16504 );
nand \U$26874 ( \27127 , \27126 , \27120 );
nand \U$26875 ( \27128 , \27125 , \27127 );
nand \U$26876 ( \27129 , \27124 , \27128 );
nand \U$26877 ( \27130 , \27119 , \27129 );
not \U$26878 ( \27131 , \27130 );
not \U$26879 ( \27132 , \27086 );
not \U$26880 ( \27133 , \27080 );
or \U$26881 ( \27134 , \27132 , \27133 );
nand \U$26882 ( \27135 , \27079 , \27083 );
nand \U$26883 ( \27136 , \27134 , \27135 );
not \U$26884 ( \27137 , \27112 );
and \U$26885 ( \27138 , \27136 , \27137 );
not \U$26886 ( \27139 , \27136 );
and \U$26887 ( \27140 , \27139 , \27112 );
nor \U$26888 ( \27141 , \27138 , \27140 );
not \U$26889 ( \27142 , \27141 );
not \U$26890 ( \27143 , \27142 );
or \U$26891 ( \27144 , \27131 , \27143 );
not \U$26892 ( \27145 , \27130 );
nand \U$26893 ( \27146 , \27141 , \27145 );
nand \U$26894 ( \27147 , \27144 , \27146 );
not \U$26895 ( \27148 , \16855 );
nand \U$26896 ( \27149 , \27148 , \16161 );
not \U$26897 ( \27150 , \27149 );
xor \U$26898 ( \27151 , \27119 , \27129 );
not \U$26899 ( \27152 , \27151 );
or \U$26900 ( \27153 , \27150 , \27152 );
or \U$26901 ( \27154 , \27149 , \27151 );
nand \U$26902 ( \27155 , \27153 , \27154 );
and \U$26903 ( \27156 , \27147 , \27155 );
nand \U$26904 ( \27157 , \26912 , \27077 , \27117 , \27156 );
nor \U$26905 ( \27158 , \25626 , \27157 );
xor \U$26906 ( \27159 , \25150 , \25611 );
xor \U$26907 ( \27160 , \27159 , \25614 );
and \U$26908 ( \27161 , \25574 , \25594 );
not \U$26909 ( \27162 , \25574 );
and \U$26910 ( \27163 , \27162 , \25595 );
nor \U$26911 ( \27164 , \27161 , \27163 );
not \U$26912 ( \27165 , \25607 );
and \U$26913 ( \27166 , \27164 , \27165 );
not \U$26914 ( \27167 , \27164 );
and \U$26915 ( \27168 , \27167 , \25607 );
nor \U$26916 ( \27169 , \27166 , \27168 );
not \U$26917 ( \27170 , \27169 );
not \U$26918 ( \27171 , \27170 );
not \U$26919 ( \27172 , \24695 );
not \U$26920 ( \27173 , \25056 );
or \U$26921 ( \27174 , \27172 , \27173 );
nand \U$26922 ( \27175 , \24694 , \25052 );
nand \U$26923 ( \27176 , \27174 , \27175 );
not \U$26924 ( \27177 , \25087 );
xor \U$26925 ( \27178 , \27176 , \27177 );
not \U$26926 ( \27179 , \27178 );
not \U$26927 ( \27180 , \27179 );
or \U$26928 ( \27181 , \27171 , \27180 );
not \U$26929 ( \27182 , \27178 );
not \U$26930 ( \27183 , \27169 );
or \U$26931 ( \27184 , \27182 , \27183 );
not \U$26932 ( \27185 , \25502 );
not \U$26933 ( \27186 , \25533 );
and \U$26934 ( \27187 , \27185 , \27186 );
and \U$26935 ( \27188 , \25502 , \25533 );
nor \U$26936 ( \27189 , \27187 , \27188 );
not \U$26937 ( \27190 , \27189 );
not \U$26938 ( \27191 , \25570 );
or \U$26939 ( \27192 , \27190 , \27191 );
or \U$26940 ( \27193 , \25570 , \27189 );
nand \U$26941 ( \27194 , \27192 , \27193 );
xor \U$26942 ( \27195 , \25581 , \25583 );
xor \U$26943 ( \27196 , \27195 , \25591 );
xor \U$26944 ( \27197 , \27194 , \27196 );
nand \U$26945 ( \27198 , \27030 , \27015 );
and \U$26946 ( \27199 , \27198 , \27022 );
nor \U$26947 ( \27200 , \27015 , \27030 );
nor \U$26948 ( \27201 , \27199 , \27200 );
not \U$26949 ( \27202 , \27201 );
not \U$26950 ( \27203 , \27003 );
not \U$26951 ( \27204 , \26997 );
or \U$26952 ( \27205 , \27203 , \27204 );
nand \U$26953 ( \27206 , \27205 , \26990 );
nand \U$26954 ( \27207 , \27006 , \26998 );
not \U$26955 ( \27208 , \26969 );
not \U$26956 ( \27209 , \26952 );
or \U$26957 ( \27210 , \27208 , \27209 );
or \U$26958 ( \27211 , \26952 , \26969 );
nand \U$26959 ( \27212 , \27211 , \26959 );
nand \U$26960 ( \27213 , \27210 , \27212 );
not \U$26961 ( \27214 , \27213 );
nand \U$26962 ( \27215 , \27206 , \27207 , \27214 );
nand \U$26963 ( \27216 , \27202 , \27215 );
nand \U$26964 ( \27217 , \27206 , \27207 );
nand \U$26965 ( \27218 , \27217 , \27213 );
nand \U$26966 ( \27219 , \27216 , \27218 );
xor \U$26967 ( \27220 , \25194 , \25188 );
xnor \U$26968 ( \27221 , \27220 , \25231 );
not \U$26969 ( \27222 , \25522 );
not \U$26970 ( \27223 , \25515 );
or \U$26971 ( \27224 , \27222 , \27223 );
or \U$26972 ( \27225 , \25515 , \25522 );
nand \U$26973 ( \27226 , \27224 , \27225 );
and \U$26974 ( \27227 , \27226 , \25525 );
not \U$26975 ( \27228 , \27226 );
and \U$26976 ( \27229 , \27228 , \25518 );
nor \U$26977 ( \27230 , \27227 , \27229 );
xor \U$26978 ( \27231 , \27221 , \27230 );
xor \U$26979 ( \27232 , \25156 , \25167 );
xnor \U$26980 ( \27233 , \27232 , \25170 );
and \U$26981 ( \27234 , \27231 , \27233 );
and \U$26982 ( \27235 , \27221 , \27230 );
or \U$26983 ( \27236 , \27234 , \27235 );
xor \U$26984 ( \27237 , \27219 , \27236 );
not \U$26985 ( \27238 , \25568 );
not \U$26986 ( \27239 , \25538 );
or \U$26987 ( \27240 , \27238 , \27239 );
nand \U$26988 ( \27241 , \25539 , \25567 );
nand \U$26989 ( \27242 , \27240 , \27241 );
and \U$26990 ( \27243 , \27242 , \25551 );
not \U$26991 ( \27244 , \27242 );
and \U$26992 ( \27245 , \27244 , \25550 );
nor \U$26993 ( \27246 , \27243 , \27245 );
and \U$26994 ( \27247 , \27237 , \27246 );
and \U$26995 ( \27248 , \27219 , \27236 );
or \U$26996 ( \27249 , \27247 , \27248 );
and \U$26997 ( \27250 , \27197 , \27249 );
and \U$26998 ( \27251 , \27194 , \27196 );
or \U$26999 ( \27252 , \27250 , \27251 );
nand \U$27000 ( \27253 , \27184 , \27252 );
nand \U$27001 ( \27254 , \27181 , \27253 );
nand \U$27002 ( \27255 , \27160 , \27254 );
not \U$27003 ( \27256 , \27255 );
nor \U$27004 ( \27257 , \27254 , \27160 );
nor \U$27005 ( \27258 , \27256 , \27257 );
not \U$27006 ( \27259 , \27040 );
not \U$27007 ( \27260 , \27046 );
not \U$27008 ( \27261 , \27260 );
or \U$27009 ( \27262 , \27259 , \27261 );
not \U$27010 ( \27263 , \27039 );
not \U$27011 ( \27264 , \27046 );
or \U$27012 ( \27265 , \27263 , \27264 );
nand \U$27013 ( \27266 , \27265 , \27054 );
nand \U$27014 ( \27267 , \27262 , \27266 );
not \U$27015 ( \27268 , \27267 );
not \U$27016 ( \27269 , \26945 );
not \U$27017 ( \27270 , \26983 );
or \U$27018 ( \27271 , \27269 , \27270 );
or \U$27019 ( \27272 , \26983 , \26945 );
nand \U$27020 ( \27273 , \27271 , \27272 );
nand \U$27021 ( \27274 , \27273 , \26940 );
not \U$27022 ( \27275 , \27274 );
not \U$27023 ( \27276 , \27275 );
or \U$27024 ( \27277 , \27268 , \27276 );
or \U$27025 ( \27278 , \27267 , \27275 );
not \U$27026 ( \27279 , \26970 );
not \U$27027 ( \27280 , \26978 );
or \U$27028 ( \27281 , \27279 , \27280 );
or \U$27029 ( \27282 , \26978 , \26970 );
nand \U$27030 ( \27283 , \27282 , \26944 );
nand \U$27031 ( \27284 , \27281 , \27283 );
xor \U$27032 ( \27285 , \25449 , \25346 );
xor \U$27033 ( \27286 , \27285 , \25491 );
not \U$27034 ( \27287 , \27286 );
not \U$27035 ( \27288 , \27287 );
not \U$27036 ( \27289 , \26926 );
not \U$27037 ( \27290 , \26921 );
or \U$27038 ( \27291 , \27289 , \27290 );
nand \U$27039 ( \27292 , \27291 , \26939 );
nand \U$27040 ( \27293 , \26922 , \26927 );
nand \U$27041 ( \27294 , \27292 , \27293 );
not \U$27042 ( \27295 , \27294 );
not \U$27043 ( \27296 , \27295 );
or \U$27044 ( \27297 , \27288 , \27296 );
nand \U$27045 ( \27298 , \27294 , \27286 );
nand \U$27046 ( \27299 , \27297 , \27298 );
not \U$27047 ( \27300 , \26988 );
not \U$27048 ( \27301 , \26991 );
not \U$27049 ( \27302 , \27008 );
or \U$27050 ( \27303 , \27301 , \27302 );
or \U$27051 ( \27304 , \27008 , \26991 );
nand \U$27052 ( \27305 , \27303 , \27304 );
not \U$27053 ( \27306 , \27305 );
or \U$27054 ( \27307 , \27300 , \27306 );
or \U$27055 ( \27308 , \27305 , \26988 );
nand \U$27056 ( \27309 , \27308 , \27035 );
nand \U$27057 ( \27310 , \27307 , \27309 );
xor \U$27058 ( \27311 , \27299 , \27310 );
xor \U$27059 ( \27312 , \27284 , \27311 );
xor \U$27060 ( \27313 , \27214 , \27217 );
xnor \U$27061 ( \27314 , \27313 , \27201 );
not \U$27062 ( \27315 , \27314 );
xor \U$27063 ( \27316 , \27221 , \27230 );
xor \U$27064 ( \27317 , \27316 , \27233 );
not \U$27065 ( \27318 , \27317 );
or \U$27066 ( \27319 , \27315 , \27318 );
or \U$27067 ( \27320 , \27317 , \27314 );
nand \U$27068 ( \27321 , \27319 , \27320 );
xor \U$27069 ( \27322 , \27312 , \27321 );
nand \U$27070 ( \27323 , \27278 , \27322 );
nand \U$27071 ( \27324 , \27277 , \27323 );
not \U$27072 ( \27325 , \27284 );
not \U$27073 ( \27326 , \27321 );
or \U$27074 ( \27327 , \27325 , \27326 );
or \U$27075 ( \27328 , \27321 , \27284 );
nand \U$27076 ( \27329 , \27328 , \27311 );
nand \U$27077 ( \27330 , \27327 , \27329 );
xnor \U$27078 ( \27331 , \25234 , \25498 );
xor \U$27079 ( \27332 , \25172 , \27331 );
xor \U$27080 ( \27333 , \27219 , \27236 );
xor \U$27081 ( \27334 , \27333 , \27246 );
and \U$27082 ( \27335 , \27332 , \27334 );
not \U$27083 ( \27336 , \27332 );
not \U$27084 ( \27337 , \27334 );
and \U$27085 ( \27338 , \27336 , \27337 );
nor \U$27086 ( \27339 , \27335 , \27338 );
xor \U$27087 ( \27340 , \27330 , \27339 );
xor \U$27088 ( \27341 , \25531 , \25511 );
xnor \U$27089 ( \27342 , \27341 , \25527 );
not \U$27090 ( \27343 , \27314 );
nand \U$27091 ( \27344 , \27343 , \27317 );
xor \U$27092 ( \27345 , \27342 , \27344 );
not \U$27093 ( \27346 , \27294 );
nand \U$27094 ( \27347 , \27346 , \27286 );
nand \U$27095 ( \27348 , \27310 , \27347 );
not \U$27096 ( \27349 , \27346 );
nand \U$27097 ( \27350 , \27349 , \27287 );
nand \U$27098 ( \27351 , \27348 , \27350 );
xnor \U$27099 ( \27352 , \27345 , \27351 );
xor \U$27100 ( \27353 , \27340 , \27352 );
xor \U$27101 ( \27354 , \27324 , \27353 );
xor \U$27102 ( \27355 , \27330 , \27339 );
and \U$27103 ( \27356 , \27355 , \27352 );
and \U$27104 ( \27357 , \27330 , \27339 );
or \U$27105 ( \27358 , \27356 , \27357 );
and \U$27106 ( \27359 , \27334 , \27332 );
not \U$27107 ( \27360 , \27342 );
not \U$27108 ( \27361 , \27351 );
or \U$27109 ( \27362 , \27360 , \27361 );
not \U$27110 ( \27363 , \27348 );
and \U$27111 ( \27364 , \27349 , \27287 );
nor \U$27112 ( \27365 , \27364 , \27342 );
not \U$27113 ( \27366 , \27365 );
or \U$27114 ( \27367 , \27363 , \27366 );
not \U$27115 ( \27368 , \27344 );
nand \U$27116 ( \27369 , \27367 , \27368 );
nand \U$27117 ( \27370 , \27362 , \27369 );
and \U$27118 ( \27371 , \27359 , \27370 );
not \U$27119 ( \27372 , \27359 );
not \U$27120 ( \27373 , \27370 );
and \U$27121 ( \27374 , \27372 , \27373 );
nor \U$27122 ( \27375 , \27371 , \27374 );
not \U$27123 ( \27376 , \27375 );
not \U$27124 ( \27377 , \27376 );
xor \U$27125 ( \27378 , \27194 , \27196 );
xor \U$27126 ( \27379 , \27378 , \27249 );
not \U$27127 ( \27380 , \27379 );
or \U$27128 ( \27381 , \27377 , \27380 );
not \U$27129 ( \27382 , \27379 );
nand \U$27130 ( \27383 , \27382 , \27375 );
nand \U$27131 ( \27384 , \27381 , \27383 );
xor \U$27132 ( \27385 , \27358 , \27384 );
nand \U$27133 ( \27386 , \27258 , \27354 , \27385 );
not \U$27134 ( \27387 , \27386 );
not \U$27135 ( \27388 , \27379 );
not \U$27136 ( \27389 , \27332 );
not \U$27137 ( \27390 , \27337 );
not \U$27138 ( \27391 , \27390 );
or \U$27139 ( \27392 , \27389 , \27391 );
nand \U$27140 ( \27393 , \27392 , \27373 );
not \U$27141 ( \27394 , \27393 );
or \U$27142 ( \27395 , \27388 , \27394 );
nand \U$27143 ( \27396 , \27370 , \27390 , \27332 );
nand \U$27144 ( \27397 , \27395 , \27396 );
not \U$27145 ( \27398 , \27397 );
xor \U$27146 ( \27399 , \27178 , \27252 );
xnor \U$27147 ( \27400 , \27399 , \27169 );
not \U$27148 ( \27401 , \27400 );
not \U$27149 ( \27402 , \27401 );
or \U$27150 ( \27403 , \27398 , \27402 );
not \U$27151 ( \27404 , \27397 );
nand \U$27152 ( \27405 , \27400 , \27404 );
nand \U$27153 ( \27406 , \27403 , \27405 );
not \U$27154 ( \27407 , \27406 );
not \U$27155 ( \27408 , \27322 );
not \U$27156 ( \27409 , \27408 );
not \U$27157 ( \27410 , \27267 );
not \U$27158 ( \27411 , \27410 );
not \U$27159 ( \27412 , \27275 );
or \U$27160 ( \27413 , \27411 , \27412 );
nand \U$27161 ( \27414 , \27267 , \27274 );
nand \U$27162 ( \27415 , \27413 , \27414 );
not \U$27163 ( \27416 , \27415 );
or \U$27164 ( \27417 , \27409 , \27416 );
or \U$27165 ( \27418 , \27415 , \27408 );
nand \U$27166 ( \27419 , \27417 , \27418 );
not \U$27167 ( \27420 , \26984 );
not \U$27168 ( \27421 , \27073 );
or \U$27169 ( \27422 , \27420 , \27421 );
not \U$27170 ( \27423 , \26985 );
not \U$27171 ( \27424 , \27070 );
or \U$27172 ( \27425 , \27423 , \27424 );
not \U$27173 ( \27426 , \27059 );
nand \U$27174 ( \27427 , \27425 , \27426 );
nand \U$27175 ( \27428 , \27422 , \27427 );
xor \U$27176 ( \27429 , \27419 , \27428 );
and \U$27177 ( \27430 , \27387 , \27407 , \27429 );
nand \U$27178 ( \27431 , \20403 , \27158 , \27430 );
not \U$27179 ( \27432 , \27431 );
not \U$27180 ( \27433 , \27075 );
nand \U$27181 ( \27434 , \27433 , \26916 );
not \U$27182 ( \27435 , \27434 );
nand \U$27183 ( \27436 , \27430 , \25625 , \27435 );
not \U$27184 ( \27437 , \25617 );
nor \U$27185 ( \27438 , \27437 , \25620 );
not \U$27186 ( \27439 , \27438 );
xor \U$27187 ( \27440 , \24684 , \25134 );
not \U$27188 ( \27441 , \27440 );
or \U$27189 ( \27442 , \27439 , \27441 );
buf \U$27190 ( \27443 , \25135 );
nand \U$27191 ( \27444 , \27442 , \27443 );
not \U$27192 ( \27445 , \23797 );
not \U$27193 ( \27446 , \27445 );
buf \U$27194 ( \27447 , \24657 );
buf \U$27195 ( \27448 , \24682 );
nand \U$27196 ( \27449 , \27444 , \27446 , \27447 , \27448 );
and \U$27197 ( \27450 , \24634 , \24656 );
not \U$27198 ( \27451 , \27450 );
not \U$27199 ( \27452 , \24682 );
or \U$27200 ( \27453 , \27451 , \27452 );
not \U$27201 ( \27454 , \24665 );
nand \U$27202 ( \27455 , \27454 , \24678 );
nand \U$27203 ( \27456 , \27453 , \27455 );
not \U$27204 ( \27457 , \27445 );
and \U$27205 ( \27458 , \27456 , \27457 );
and \U$27206 ( \27459 , \23232 , \23796 );
nor \U$27207 ( \27460 , \27458 , \27459 );
nand \U$27208 ( \27461 , \27449 , \27460 );
not \U$27209 ( \27462 , \12752 );
not \U$27210 ( \27463 , \3537 );
and \U$27211 ( \27464 , \27462 , \27463 );
and \U$27212 ( \27465 , \14726 , RIbe281b0_15);
nor \U$27213 ( \27466 , \27464 , \27465 );
and \U$27214 ( \27467 , \27466 , \12770 );
not \U$27215 ( \27468 , \27466 );
and \U$27216 ( \27469 , \27468 , \12927 );
nor \U$27217 ( \27470 , \27467 , \27469 );
not \U$27218 ( \27471 , RIbe29830_63);
not \U$27219 ( \27472 , \16383 );
or \U$27220 ( \27473 , \27471 , \27472 );
nand \U$27221 ( \27474 , \13728 , RIbe296c8_60);
nand \U$27222 ( \27475 , \27473 , \27474 );
and \U$27223 ( \27476 , \27475 , \13068 );
not \U$27224 ( \27477 , \27475 );
and \U$27225 ( \27478 , \27477 , \12723 );
nor \U$27226 ( \27479 , \27476 , \27478 );
xor \U$27227 ( \27480 , \27470 , \27479 );
not \U$27228 ( \27481 , RIbe29650_59);
not \U$27229 ( \27482 , \12732 );
or \U$27230 ( \27483 , \27481 , \27482 );
nand \U$27231 ( \27484 , \14074 , RIbe29038_46);
nand \U$27232 ( \27485 , \27483 , \27484 );
and \U$27233 ( \27486 , \27485 , \12743 );
not \U$27234 ( \27487 , \27485 );
and \U$27235 ( \27488 , \27487 , \12742 );
nor \U$27236 ( \27489 , \27486 , \27488 );
and \U$27237 ( \27490 , \27480 , \27489 );
and \U$27238 ( \27491 , \27470 , \27479 );
or \U$27239 ( \27492 , \27490 , \27491 );
and \U$27240 ( \27493 , \8278 , RIbe29290_51);
and \U$27241 ( \27494 , \13643 , RIbe28a20_33);
nor \U$27242 ( \27495 , \27493 , \27494 );
and \U$27243 ( \27496 , \27495 , \8077 );
not \U$27244 ( \27497 , \27495 );
and \U$27245 ( \27498 , \27497 , \7970 );
nor \U$27246 ( \27499 , \27496 , \27498 );
not \U$27247 ( \27500 , RIbe29560_57);
not \U$27248 ( \27501 , \13049 );
or \U$27249 ( \27502 , \27500 , \27501 );
nand \U$27250 ( \27503 , \12948 , RIbe28228_16);
nand \U$27251 ( \27504 , \27502 , \27503 );
and \U$27252 ( \27505 , \27504 , \12195 );
not \U$27253 ( \27506 , \27504 );
and \U$27254 ( \27507 , \27506 , \17005 );
nor \U$27255 ( \27508 , \27505 , \27507 );
xor \U$27256 ( \27509 , \27499 , \27508 );
not \U$27257 ( \27510 , RIbe289a8_32);
not \U$27258 ( \27511 , \10936 );
or \U$27259 ( \27512 , \27510 , \27511 );
nand \U$27260 ( \27513 , \14511 , RIbe28930_31);
nand \U$27261 ( \27514 , \27512 , \27513 );
and \U$27262 ( \27515 , \27514 , \9902 );
not \U$27263 ( \27516 , \27514 );
and \U$27264 ( \27517 , \27516 , \13030 );
nor \U$27265 ( \27518 , \27515 , \27517 );
and \U$27266 ( \27519 , \27509 , \27518 );
and \U$27267 ( \27520 , \27499 , \27508 );
or \U$27268 ( \27521 , \27519 , \27520 );
xor \U$27269 ( \27522 , \27492 , \27521 );
not \U$27270 ( \27523 , RIbe27d00_5);
not \U$27271 ( \27524 , \13003 );
or \U$27272 ( \27525 , \27523 , \27524 );
nand \U$27273 ( \27526 , RIbe27c10_3, RIbe2ae38_110);
nand \U$27274 ( \27527 , \27525 , \27526 );
xor \U$27275 ( \27528 , \27527 , RIbe2aeb0_111);
not \U$27276 ( \27529 , \27528 );
not \U$27277 ( \27530 , RIbe29a88_68);
not \U$27278 ( \27531 , \15249 );
or \U$27279 ( \27532 , \27530 , \27531 );
nand \U$27280 ( \27533 , \12794 , RIbe27d78_6);
nand \U$27281 ( \27534 , \27532 , \27533 );
not \U$27282 ( \27535 , \27534 );
not \U$27283 ( \27536 , \14335 );
and \U$27284 ( \27537 , \27535 , \27536 );
and \U$27285 ( \27538 , \27534 , \12893 );
nor \U$27286 ( \27539 , \27537 , \27538 );
not \U$27287 ( \27540 , \27539 );
not \U$27288 ( \27541 , \27540 );
or \U$27289 ( \27542 , \27529 , \27541 );
not \U$27290 ( \27543 , RIbe28fc0_45);
not \U$27291 ( \27544 , \13590 );
or \U$27292 ( \27545 , \27543 , \27544 );
nand \U$27293 ( \27546 , \12835 , RIbe290b0_47);
nand \U$27294 ( \27547 , \27545 , \27546 );
not \U$27295 ( \27548 , \27547 );
not \U$27296 ( \27549 , \14558 );
and \U$27297 ( \27550 , \27548 , \27549 );
and \U$27298 ( \27551 , \27547 , \12823 );
nor \U$27299 ( \27552 , \27550 , \27551 );
not \U$27300 ( \27553 , \27552 );
not \U$27301 ( \27554 , \27528 );
nand \U$27302 ( \27555 , \27554 , \27539 );
nand \U$27303 ( \27556 , \27553 , \27555 );
nand \U$27304 ( \27557 , \27542 , \27556 );
xor \U$27305 ( \27558 , \27522 , \27557 );
not \U$27306 ( \27559 , RIbe2a3e8_88);
not \U$27307 ( \27560 , \6797 );
or \U$27308 ( \27561 , \27559 , \27560 );
nand \U$27309 ( \27562 , \3457 , RIbe2a370_87);
nand \U$27310 ( \27563 , \27561 , \27562 );
and \U$27311 ( \27564 , \27563 , \2887 );
not \U$27312 ( \27565 , \27563 );
and \U$27313 ( \27566 , \27565 , \3290 );
nor \U$27314 ( \27567 , \27564 , \27566 );
not \U$27315 ( \27568 , RIbe2a028_80);
not \U$27316 ( \27569 , \21040 );
or \U$27317 ( \27570 , \27568 , \27569 );
nand \U$27318 ( \27571 , \4599 , RIbe29fb0_79);
nand \U$27319 ( \27572 , \27570 , \27571 );
not \U$27320 ( \27573 , \27572 );
not \U$27321 ( \27574 , \4323 );
and \U$27322 ( \27575 , \27573 , \27574 );
and \U$27323 ( \27576 , \27572 , \4322 );
nor \U$27324 ( \27577 , \27575 , \27576 );
nand \U$27325 ( \27578 , \27567 , \27577 );
not \U$27326 ( \27579 , RIbe2a2f8_86);
not \U$27327 ( \27580 , \20625 );
or \U$27328 ( \27581 , \27579 , \27580 );
nand \U$27329 ( \27582 , \6787 , RIbe2acd0_107);
nand \U$27330 ( \27583 , \27581 , \27582 );
and \U$27331 ( \27584 , \27583 , \3471 );
not \U$27332 ( \27585 , \27583 );
and \U$27333 ( \27586 , \27585 , \3448 );
nor \U$27334 ( \27587 , \27584 , \27586 );
and \U$27335 ( \27588 , \27578 , \27587 );
nor \U$27336 ( \27589 , \27567 , \27577 );
nor \U$27337 ( \27590 , \27588 , \27589 );
not \U$27338 ( \27591 , \27590 );
not \U$27339 ( \27592 , RIbe2a910_99);
not \U$27340 ( \27593 , \7007 );
or \U$27341 ( \27594 , \27592 , \27593 );
nand \U$27342 ( \27595 , \4284 , RIbe2b5b8_126);
nand \U$27343 ( \27596 , \27594 , \27595 );
and \U$27344 ( \27597 , \27596 , \4059 );
not \U$27345 ( \27598 , \27596 );
and \U$27346 ( \27599 , \27598 , \7457 );
nor \U$27347 ( \27600 , \27597 , \27599 );
not \U$27348 ( \27601 , \1284 );
and \U$27349 ( \27602 , \27601 , RIbe2a190_83);
and \U$27350 ( \27603 , \5467 , RIbe2a5c8_92);
nor \U$27351 ( \27604 , \27602 , \27603 );
and \U$27352 ( \27605 , \27604 , \1131 );
not \U$27353 ( \27606 , \27604 );
and \U$27354 ( \27607 , \27606 , \3491 );
nor \U$27355 ( \27608 , \27605 , \27607 );
nand \U$27356 ( \27609 , \27600 , \27608 );
not \U$27357 ( \27610 , \2385 );
not \U$27358 ( \27611 , \13552 );
and \U$27359 ( \27612 , \27610 , \27611 );
not \U$27360 ( \27613 , \2389 );
buf \U$27361 ( \27614 , \27613 );
and \U$27362 ( \27615 , \27614 , RIbe2a550_91);
nor \U$27363 ( \27616 , \27612 , \27615 );
and \U$27364 ( \27617 , \27616 , \1277 );
not \U$27365 ( \27618 , \27616 );
and \U$27366 ( \27619 , \27618 , \1076 );
nor \U$27367 ( \27620 , \27617 , \27619 );
not \U$27368 ( \27621 , \27620 );
and \U$27369 ( \27622 , \27609 , \27621 );
nor \U$27370 ( \27623 , \27600 , \27608 );
nor \U$27371 ( \27624 , \27622 , \27623 );
not \U$27372 ( \27625 , \27624 );
not \U$27373 ( \27626 , \27625 );
or \U$27374 ( \27627 , \27591 , \27626 );
not \U$27375 ( \27628 , \27590 );
nand \U$27376 ( \27629 , \27628 , \27624 );
nand \U$27377 ( \27630 , \27627 , \27629 );
not \U$27378 ( \27631 , \27630 );
and \U$27379 ( \27632 , \1807 , RIbe2b180_117);
and \U$27380 ( \27633 , \1203 , RIbe2b270_119);
nor \U$27381 ( \27634 , \27632 , \27633 );
and \U$27382 ( \27635 , \27634 , \752 );
not \U$27383 ( \27636 , \27634 );
and \U$27384 ( \27637 , \27636 , \1011 );
nor \U$27385 ( \27638 , \27635 , \27637 );
not \U$27386 ( \27639 , RIbe2b108_116);
not \U$27387 ( \27640 , \4257 );
or \U$27388 ( \27641 , \27639 , \27640 );
nand \U$27389 ( \27642 , \1147 , RIbe2b090_115);
nand \U$27390 ( \27643 , \27641 , \27642 );
and \U$27391 ( \27644 , \27643 , \1153 );
not \U$27392 ( \27645 , \27643 );
and \U$27393 ( \27646 , \27645 , \7899 );
nor \U$27394 ( \27647 , \27644 , \27646 );
not \U$27395 ( \27648 , \27647 );
or \U$27396 ( \27649 , \27638 , \27648 );
not \U$27397 ( \27650 , RIbe2a280_85);
not \U$27398 ( \27651 , \1633 );
or \U$27399 ( \27652 , \27650 , \27651 );
nand \U$27400 ( \27653 , \1455 , RIbe2a208_84);
nand \U$27401 ( \27654 , \27652 , \27653 );
and \U$27402 ( \27655 , \27654 , \1309 );
not \U$27403 ( \27656 , \27654 );
and \U$27404 ( \27657 , \27656 , \1082 );
nor \U$27405 ( \27658 , \27655 , \27657 );
nand \U$27406 ( \27659 , \27649 , \27658 );
nand \U$27407 ( \27660 , \27638 , \27648 );
nand \U$27408 ( \27661 , \27659 , \27660 );
not \U$27409 ( \27662 , \27661 );
not \U$27410 ( \27663 , \27662 );
and \U$27411 ( \27664 , \27631 , \27663 );
and \U$27412 ( \27665 , \27630 , \27662 );
nor \U$27413 ( \27666 , \27664 , \27665 );
not \U$27414 ( \27667 , \27666 );
not \U$27415 ( \27668 , \27667 );
not \U$27416 ( \27669 , RIbe2acd0_107);
not \U$27417 ( \27670 , \20625 );
or \U$27418 ( \27671 , \27669 , \27670 );
nand \U$27419 ( \27672 , \7438 , RIbe2a028_80);
nand \U$27420 ( \27673 , \27671 , \27672 );
and \U$27421 ( \27674 , \27673 , \3471 );
not \U$27422 ( \27675 , \27673 );
and \U$27423 ( \27676 , \27675 , \3698 );
nor \U$27424 ( \27677 , \27674 , \27676 );
not \U$27425 ( \27678 , RIbe2a370_87);
not \U$27426 ( \27679 , \3451 );
or \U$27427 ( \27680 , \27678 , \27679 );
nand \U$27428 ( \27681 , \3457 , RIbe2a2f8_86);
nand \U$27429 ( \27682 , \27680 , \27681 );
and \U$27430 ( \27683 , \27682 , \4346 );
not \U$27431 ( \27684 , \27682 );
and \U$27432 ( \27685 , \27684 , \3461 );
nor \U$27433 ( \27686 , \27683 , \27685 );
xor \U$27434 ( \27687 , \27677 , \27686 );
not \U$27435 ( \27688 , RIbe2b5b8_126);
not \U$27436 ( \27689 , \8342 );
or \U$27437 ( \27690 , \27688 , \27689 );
nand \U$27438 ( \27691 , \4284 , RIbe2a3e8_88);
nand \U$27439 ( \27692 , \27690 , \27691 );
and \U$27440 ( \27693 , \27692 , \3272 );
not \U$27441 ( \27694 , \27692 );
and \U$27442 ( \27695 , \27694 , \4783 );
nor \U$27443 ( \27696 , \27693 , \27695 );
xor \U$27444 ( \27697 , \27687 , \27696 );
not \U$27445 ( \27698 , \27697 );
not \U$27446 ( \27699 , RIbe29bf0_71);
not \U$27447 ( \27700 , \20796 );
or \U$27448 ( \27701 , \27699 , \27700 );
nand \U$27449 ( \27702 , \6633 , RIbe28f48_44);
nand \U$27450 ( \27703 , \27701 , \27702 );
and \U$27451 ( \27704 , \27703 , \5460 );
not \U$27452 ( \27705 , \27703 );
and \U$27453 ( \27706 , \27705 , \5754 );
nor \U$27454 ( \27707 , \27704 , \27706 );
not \U$27455 ( \27708 , \27707 );
not \U$27456 ( \27709 , RIbe29dd0_75);
not \U$27457 ( \27710 , \20809 );
or \U$27458 ( \27711 , \27709 , \27710 );
nand \U$27459 ( \27712 , \5052 , RIbe29c68_72);
nand \U$27460 ( \27713 , \27711 , \27712 );
and \U$27461 ( \27714 , \27713 , \20465 );
not \U$27462 ( \27715 , \27713 );
and \U$27463 ( \27716 , \27715 , \4586 );
nor \U$27464 ( \27717 , \27714 , \27716 );
not \U$27465 ( \27718 , \27717 );
nand \U$27466 ( \27719 , \27708 , \27718 );
nand \U$27467 ( \27720 , \27717 , \27707 );
nand \U$27468 ( \27721 , \27719 , \27720 );
not \U$27469 ( \27722 , RIbe29fb0_79);
not \U$27470 ( \27723 , \4317 );
or \U$27471 ( \27724 , \27722 , \27723 );
nand \U$27472 ( \27725 , \7858 , RIbe29e48_76);
nand \U$27473 ( \27726 , \27724 , \27725 );
xor \U$27474 ( \27727 , \27726 , \4323 );
and \U$27475 ( \27728 , \27721 , \27727 );
not \U$27476 ( \27729 , \27721 );
not \U$27477 ( \27730 , \27727 );
and \U$27478 ( \27731 , \27729 , \27730 );
nor \U$27479 ( \27732 , \27728 , \27731 );
not \U$27480 ( \27733 , \27732 );
or \U$27481 ( \27734 , \27698 , \27733 );
or \U$27482 ( \27735 , \27697 , \27732 );
nand \U$27483 ( \27736 , \27734 , \27735 );
and \U$27484 ( \27737 , \10759 , RIbe2a5c8_92);
and \U$27485 ( \27738 , \5467 , RIbe2a550_91);
nor \U$27486 ( \27739 , \27737 , \27738 );
and \U$27487 ( \27740 , \27739 , \6831 );
not \U$27488 ( \27741 , \27739 );
and \U$27489 ( \27742 , \27741 , \1131 );
nor \U$27490 ( \27743 , \27740 , \27742 );
not \U$27491 ( \27744 , \2889 );
not \U$27492 ( \27745 , RIbe2a910_99);
not \U$27493 ( \27746 , \27745 );
and \U$27494 ( \27747 , \27744 , \27746 );
and \U$27495 ( \27748 , \8833 , RIbe2a988_100);
nor \U$27496 ( \27749 , \27747 , \27748 );
and \U$27497 ( \27750 , \27749 , \24063 );
not \U$27498 ( \27751 , \27749 );
and \U$27499 ( \27752 , \27751 , \1076 );
nor \U$27500 ( \27753 , \27750 , \27752 );
and \U$27501 ( \27754 , \27743 , \27753 );
not \U$27502 ( \27755 , \27743 );
not \U$27503 ( \27756 , \27753 );
and \U$27504 ( \27757 , \27755 , \27756 );
nor \U$27505 ( \27758 , \27754 , \27757 );
not \U$27506 ( \27759 , RIbe2a208_84);
not \U$27507 ( \27760 , \1094 );
or \U$27508 ( \27761 , \27759 , \27760 );
nand \U$27509 ( \27762 , \1455 , RIbe2a190_83);
nand \U$27510 ( \27763 , \27761 , \27762 );
and \U$27511 ( \27764 , \27763 , \1309 );
not \U$27512 ( \27765 , \27763 );
and \U$27513 ( \27766 , \27765 , \5125 );
nor \U$27514 ( \27767 , \27764 , \27766 );
xor \U$27515 ( \27768 , \27758 , \27767 );
not \U$27516 ( \27769 , \27768 );
and \U$27517 ( \27770 , \27736 , \27769 );
not \U$27518 ( \27771 , \27736 );
and \U$27519 ( \27772 , \27771 , \27768 );
nor \U$27520 ( \27773 , \27770 , \27772 );
buf \U$27521 ( \27774 , \27773 );
not \U$27522 ( \27775 , \27774 );
or \U$27523 ( \27776 , \27668 , \27775 );
or \U$27524 ( \27777 , \27774 , \27667 );
not \U$27525 ( \27778 , RIbe2b018_114);
not \U$27526 ( \27779 , \3244 );
or \U$27527 ( \27780 , \27778 , \27779 );
nand \U$27528 ( \27781 , \552 , RIbe2afa0_113);
nand \U$27529 ( \27782 , \27780 , \27781 );
and \U$27530 ( \27783 , \27782 , \3415 );
not \U$27531 ( \27784 , \27782 );
and \U$27532 ( \27785 , \27784 , \424 );
nor \U$27533 ( \27786 , \27783 , \27785 );
not \U$27534 ( \27787 , RIbe2aaf0_103);
not \U$27535 ( \27788 , \383 );
or \U$27536 ( \27789 , \27787 , \27788 );
nand \U$27537 ( \27790 , \429 , RIbe2b630_127);
nand \U$27538 ( \27791 , \27789 , \27790 );
and \U$27539 ( \27792 , \27791 , \306 );
not \U$27540 ( \27793 , \27791 );
and \U$27541 ( \27794 , \27793 , \1547 );
nor \U$27542 ( \27795 , \27792 , \27794 );
or \U$27543 ( \27796 , \27786 , \27795 );
and \U$27544 ( \27797 , \2531 , RIbe2af28_112);
not \U$27545 ( \27798 , RIbe2b1f8_118);
nor \U$27546 ( \27799 , \27798 , \1611 );
nor \U$27547 ( \27800 , \27797 , \27799 );
and \U$27548 ( \27801 , \27800 , \564 );
not \U$27549 ( \27802 , \27800 );
and \U$27550 ( \27803 , \27802 , \1621 );
nor \U$27551 ( \27804 , \27801 , \27803 );
nand \U$27552 ( \27805 , \27796 , \27804 );
nand \U$27553 ( \27806 , \27786 , \27795 );
and \U$27554 ( \27807 , \27805 , \27806 );
not \U$27555 ( \27808 , \27807 );
not \U$27556 ( \27809 , RIbe2b1f8_118);
not \U$27557 ( \27810 , \664 );
or \U$27558 ( \27811 , \27809 , \27810 );
nand \U$27559 ( \27812 , \1179 , RIbe2b180_117);
nand \U$27560 ( \27813 , \27811 , \27812 );
xor \U$27561 ( \27814 , \27813 , \564 );
not \U$27562 ( \27815 , RIbe2b090_115);
not \U$27563 ( \27816 , \4257 );
or \U$27564 ( \27817 , \27815 , \27816 );
nand \U$27565 ( \27818 , \1146 , RIbe2a280_85);
nand \U$27566 ( \27819 , \27817 , \27818 );
and \U$27567 ( \27820 , \27819 , \3993 );
not \U$27568 ( \27821 , \27819 );
and \U$27569 ( \27822 , \27821 , \1157 );
nor \U$27570 ( \27823 , \27820 , \27822 );
xor \U$27571 ( \27824 , \27814 , \27823 );
and \U$27572 ( \27825 , \1807 , RIbe2b270_119);
and \U$27573 ( \27826 , \1203 , RIbe2b108_116);
nor \U$27574 ( \27827 , \27825 , \27826 );
and \U$27575 ( \27828 , \27827 , \750 );
not \U$27576 ( \27829 , \27827 );
and \U$27577 ( \27830 , \27829 , \1011 );
nor \U$27578 ( \27831 , \27828 , \27830 );
xnor \U$27579 ( \27832 , \27824 , \27831 );
not \U$27580 ( \27833 , \27832 );
or \U$27581 ( \27834 , \27808 , \27833 );
or \U$27582 ( \27835 , \27832 , \27807 );
nand \U$27583 ( \27836 , \27834 , \27835 );
not \U$27584 ( \27837 , RIbe2b630_127);
not \U$27585 ( \27838 , \9239 );
or \U$27586 ( \27839 , \27837 , \27838 );
nand \U$27587 ( \27840 , \429 , RIbe2b018_114);
nand \U$27588 ( \27841 , \27839 , \27840 );
and \U$27589 ( \27842 , \27841 , \306 );
not \U$27590 ( \27843 , \27841 );
and \U$27591 ( \27844 , \27843 , \313 );
nor \U$27592 ( \27845 , \27842 , \27844 );
not \U$27593 ( \27846 , \27845 );
not \U$27594 ( \27847 , RIbe2afa0_113);
not \U$27595 ( \27848 , \546 );
or \U$27596 ( \27849 , \27847 , \27848 );
nand \U$27597 ( \27850 , \552 , RIbe2af28_112);
nand \U$27598 ( \27851 , \27849 , \27850 );
not \U$27599 ( \27852 , \27851 );
not \U$27600 ( \27853 , \7124 );
and \U$27601 ( \27854 , \27852 , \27853 );
and \U$27602 ( \27855 , \27851 , \7124 );
nor \U$27603 ( \27856 , \27854 , \27855 );
not \U$27604 ( \27857 , \27856 );
or \U$27605 ( \27858 , \27846 , \27857 );
or \U$27606 ( \27859 , \27856 , \27845 );
nand \U$27607 ( \27860 , \27858 , \27859 );
and \U$27608 ( \27861 , \1528 , RIbe2ab68_104);
and \U$27609 ( \27862 , \1531 , RIbe2aaf0_103);
nor \U$27610 ( \27863 , \27861 , \27862 );
and \U$27611 ( \27864 , \27863 , \293 );
not \U$27612 ( \27865 , \27863 );
and \U$27613 ( \27866 , \27865 , \300 );
nor \U$27614 ( \27867 , \27864 , \27866 );
and \U$27615 ( \27868 , \27860 , \27867 );
not \U$27616 ( \27869 , \27860 );
not \U$27617 ( \27870 , \27867 );
and \U$27618 ( \27871 , \27869 , \27870 );
nor \U$27619 ( \27872 , \27868 , \27871 );
buf \U$27620 ( \27873 , \27872 );
not \U$27621 ( \27874 , \27873 );
and \U$27622 ( \27875 , \27836 , \27874 );
not \U$27623 ( \27876 , \27836 );
and \U$27624 ( \27877 , \27876 , \27873 );
nor \U$27625 ( \27878 , \27875 , \27877 );
nand \U$27626 ( \27879 , \27777 , \27878 );
nand \U$27627 ( \27880 , \27776 , \27879 );
xor \U$27628 ( \27881 , \27558 , \27880 );
or \U$27629 ( \27882 , \27823 , \27831 );
not \U$27630 ( \27883 , \27814 );
nand \U$27631 ( \27884 , \27882 , \27883 );
nand \U$27632 ( \27885 , \27831 , \27823 );
nand \U$27633 ( \27886 , \27884 , \27885 );
xor \U$27634 ( \27887 , \27677 , \27686 );
and \U$27635 ( \27888 , \27887 , \27696 );
and \U$27636 ( \27889 , \27677 , \27686 );
or \U$27637 ( \27890 , \27888 , \27889 );
xor \U$27638 ( \27891 , \27886 , \27890 );
or \U$27639 ( \27892 , \27767 , \27743 );
nand \U$27640 ( \27893 , \27892 , \27756 );
nand \U$27641 ( \27894 , \27767 , \27743 );
nand \U$27642 ( \27895 , \27893 , \27894 );
xor \U$27643 ( \27896 , \27891 , \27895 );
not \U$27644 ( \27897 , RIbe287c8_28);
not \U$27645 ( \27898 , \13327 );
or \U$27646 ( \27899 , \27897 , \27898 );
nand \U$27647 ( \27900 , \8202 , RIbe28480_21);
nand \U$27648 ( \27901 , \27899 , \27900 );
and \U$27649 ( \27902 , \27901 , \7293 );
not \U$27650 ( \27903 , \27901 );
and \U$27651 ( \27904 , \27903 , \6572 );
nor \U$27652 ( \27905 , \27902 , \27904 );
not \U$27653 ( \27906 , RIbe28b10_35);
not \U$27654 ( \27907 , \14633 );
or \U$27655 ( \27908 , \27906 , \27907 );
nand \U$27656 ( \27909 , \8269 , RIbe28b88_36);
nand \U$27657 ( \27910 , \27908 , \27909 );
and \U$27658 ( \27911 , \27910 , \9896 );
not \U$27659 ( \27912 , \27910 );
and \U$27660 ( \27913 , \27912 , \6949 );
nor \U$27661 ( \27914 , \27911 , \27913 );
or \U$27662 ( \27915 , \27905 , \27914 );
not \U$27663 ( \27916 , RIbe28408_20);
not \U$27664 ( \27917 , \6980 );
or \U$27665 ( \27918 , \27916 , \27917 );
nand \U$27666 ( \27919 , \13224 , RIbe28390_19);
nand \U$27667 ( \27920 , \27918 , \27919 );
not \U$27668 ( \27921 , \27920 );
not \U$27669 ( \27922 , \8004 );
and \U$27670 ( \27923 , \27921 , \27922 );
and \U$27671 ( \27924 , \27920 , \7301 );
nor \U$27672 ( \27925 , \27923 , \27924 );
not \U$27673 ( \27926 , \27925 );
nand \U$27674 ( \27927 , \27915 , \27926 );
nand \U$27675 ( \27928 , \27905 , \27914 );
nand \U$27676 ( \27929 , \27927 , \27928 );
not \U$27677 ( \27930 , \27707 );
not \U$27678 ( \27931 , \27730 );
or \U$27679 ( \27932 , \27930 , \27931 );
or \U$27680 ( \27933 , \27730 , \27707 );
nand \U$27681 ( \27934 , \27933 , \27718 );
nand \U$27682 ( \27935 , \27932 , \27934 );
xor \U$27683 ( \27936 , \27929 , \27935 );
not \U$27684 ( \27937 , RIbe28660_25);
not \U$27685 ( \27938 , \6591 );
or \U$27686 ( \27939 , \27937 , \27938 );
nand \U$27687 ( \27940 , \13436 , RIbe285e8_24);
nand \U$27688 ( \27941 , \27939 , \27940 );
and \U$27689 ( \27942 , \27941 , \7948 );
not \U$27690 ( \27943 , \27941 );
and \U$27691 ( \27944 , \27943 , \7949 );
nor \U$27692 ( \27945 , \27942 , \27944 );
not \U$27693 ( \27946 , \6883 );
not \U$27694 ( \27947 , \6347 );
and \U$27695 ( \27948 , \27946 , \27947 );
and \U$27696 ( \27949 , \6535 , RIbe27f58_10);
nor \U$27697 ( \27950 , \27948 , \27949 );
and \U$27698 ( \27951 , \27950 , \6891 );
not \U$27699 ( \27952 , \27950 );
and \U$27700 ( \27953 , \27952 , \7935 );
nor \U$27701 ( \27954 , \27951 , \27953 );
xor \U$27702 ( \27955 , \27945 , \27954 );
not \U$27703 ( \27956 , RIbe28ed0_43);
not \U$27704 ( \27957 , \8231 );
or \U$27705 ( \27958 , \27956 , \27957 );
nand \U$27706 ( \27959 , \6617 , RIbe27fd0_11);
nand \U$27707 ( \27960 , \27958 , \27959 );
and \U$27708 ( \27961 , \27960 , \6620 );
not \U$27709 ( \27962 , \27960 );
and \U$27710 ( \27963 , \27962 , \5740 );
nor \U$27711 ( \27964 , \27961 , \27963 );
and \U$27712 ( \27965 , \27955 , \27964 );
and \U$27713 ( \27966 , \27945 , \27954 );
or \U$27714 ( \27967 , \27965 , \27966 );
xor \U$27715 ( \27968 , \27936 , \27967 );
xor \U$27716 ( \27969 , \27896 , \27968 );
nand \U$27717 ( \27970 , \264 , RIbe2ab68_104);
and \U$27718 ( \27971 , \27970 , \269 );
not \U$27719 ( \27972 , \27970 );
and \U$27720 ( \27973 , \27972 , \1362 );
nor \U$27721 ( \27974 , \27971 , \27973 );
not \U$27722 ( \27975 , \27974 );
and \U$27723 ( \27976 , \283 , RIbe2aaf0_103);
and \U$27724 ( \27977 , \1256 , RIbe2b630_127);
nor \U$27725 ( \27978 , \27976 , \27977 );
and \U$27726 ( \27979 , \27978 , \300 );
not \U$27727 ( \27980 , \27978 );
and \U$27728 ( \27981 , \27980 , \293 );
nor \U$27729 ( \27982 , \27979 , \27981 );
not \U$27730 ( \27983 , \27982 );
or \U$27731 ( \27984 , \27975 , \27983 );
or \U$27732 ( \27985 , \27982 , \27974 );
nand \U$27733 ( \27986 , \27984 , \27985 );
not \U$27734 ( \27987 , \27867 );
not \U$27735 ( \27988 , \27856 );
or \U$27736 ( \27989 , \27987 , \27988 );
nand \U$27737 ( \27990 , \27989 , \27845 );
not \U$27738 ( \27991 , \27856 );
nand \U$27739 ( \27992 , \27991 , \27870 );
nand \U$27740 ( \27993 , \27990 , \27992 );
xor \U$27741 ( \27994 , \27986 , \27993 );
not \U$27742 ( \27995 , \6345 );
not \U$27743 ( \27996 , \13109 );
and \U$27744 ( \27997 , \27995 , \27996 );
and \U$27745 ( \27998 , \1744 , RIbe2b180_117);
nor \U$27746 ( \27999 , \27997 , \27998 );
and \U$27747 ( \28000 , \27999 , \1618 );
not \U$27748 ( \28001 , \27999 );
and \U$27749 ( \28002 , \28001 , \1621 );
nor \U$27750 ( \28003 , \28000 , \28002 );
not \U$27751 ( \28004 , RIbe2af28_112);
not \U$27752 ( \28005 , \546 );
or \U$27753 ( \28006 , \28004 , \28005 );
nand \U$27754 ( \28007 , \552 , RIbe2b1f8_118);
nand \U$27755 ( \28008 , \28006 , \28007 );
not \U$27756 ( \28009 , \28008 );
not \U$27757 ( \28010 , \1333 );
and \U$27758 ( \28011 , \28009 , \28010 );
and \U$27759 ( \28012 , \28008 , \6340 );
nor \U$27760 ( \28013 , \28011 , \28012 );
xor \U$27761 ( \28014 , \28003 , \28013 );
not \U$27762 ( \28015 , RIbe2b018_114);
not \U$27763 ( \28016 , \1337 );
or \U$27764 ( \28017 , \28015 , \28016 );
nand \U$27765 ( \28018 , \429 , RIbe2afa0_113);
nand \U$27766 ( \28019 , \28017 , \28018 );
and \U$27767 ( \28020 , \28019 , \3175 );
not \U$27768 ( \28021 , \28019 );
and \U$27769 ( \28022 , \28021 , \306 );
nor \U$27770 ( \28023 , \28020 , \28022 );
xor \U$27771 ( \28024 , \28014 , \28023 );
xor \U$27772 ( \28025 , \27994 , \28024 );
and \U$27773 ( \28026 , \27969 , \28025 );
not \U$27774 ( \28027 , \27969 );
not \U$27775 ( \28028 , \28025 );
and \U$27776 ( \28029 , \28027 , \28028 );
nor \U$27777 ( \28030 , \28026 , \28029 );
and \U$27778 ( \28031 , \27881 , \28030 );
and \U$27779 ( \28032 , \27558 , \27880 );
or \U$27780 ( \28033 , \28031 , \28032 );
not \U$27781 ( \28034 , \28033 );
not \U$27782 ( \28035 , \28034 );
not \U$27783 ( \28036 , \27624 );
not \U$27784 ( \28037 , \27590 );
or \U$27785 ( \28038 , \28036 , \28037 );
nand \U$27786 ( \28039 , \28038 , \27661 );
not \U$27787 ( \28040 , \27590 );
nand \U$27788 ( \28041 , \28040 , \27625 );
nand \U$27789 ( \28042 , \28039 , \28041 );
not \U$27790 ( \28043 , \28042 );
not \U$27791 ( \28044 , \28043 );
not \U$27792 ( \28045 , RIbe29e48_76);
not \U$27793 ( \28046 , \15894 );
or \U$27794 ( \28047 , \28045 , \28046 );
nand \U$27795 ( \28048 , \22378 , RIbe29dd0_75);
nand \U$27796 ( \28049 , \28047 , \28048 );
and \U$27797 ( \28050 , \28049 , \20465 );
not \U$27798 ( \28051 , \28049 );
and \U$27799 ( \28052 , \28051 , \4586 );
nor \U$27800 ( \28053 , \28050 , \28052 );
not \U$27801 ( \28054 , RIbe28f48_44);
not \U$27802 ( \28055 , \6138 );
or \U$27803 ( \28056 , \28054 , \28055 );
nand \U$27804 ( \28057 , \8235 , RIbe28ed0_43);
nand \U$27805 ( \28058 , \28056 , \28057 );
not \U$27806 ( \28059 , \28058 );
not \U$27807 ( \28060 , \21090 );
and \U$27808 ( \28061 , \28059 , \28060 );
and \U$27809 ( \28062 , \28058 , \9944 );
nor \U$27810 ( \28063 , \28061 , \28062 );
nand \U$27811 ( \28064 , \28053 , \28063 );
not \U$27812 ( \28065 , RIbe29c68_72);
not \U$27813 ( \28066 , \6630 );
or \U$27814 ( \28067 , \28065 , \28066 );
nand \U$27815 ( \28068 , \15885 , RIbe29bf0_71);
nand \U$27816 ( \28069 , \28067 , \28068 );
and \U$27817 ( \28070 , \28069 , \6117 );
not \U$27818 ( \28071 , \28069 );
and \U$27819 ( \28072 , \28071 , \6637 );
nor \U$27820 ( \28073 , \28070 , \28072 );
and \U$27821 ( \28074 , \28064 , \28073 );
nor \U$27822 ( \28075 , \28053 , \28063 );
nor \U$27823 ( \28076 , \28074 , \28075 );
not \U$27824 ( \28077 , RIbe27e68_8);
not \U$27825 ( \28078 , \7274 );
or \U$27826 ( \28079 , \28077 , \28078 );
nand \U$27827 ( \28080 , \7278 , RIbe28660_25);
nand \U$27828 ( \28081 , \28079 , \28080 );
and \U$27829 ( \28082 , \28081 , \14991 );
not \U$27830 ( \28083 , \28081 );
and \U$27831 ( \28084 , \28083 , \7948 );
nor \U$27832 ( \28085 , \28082 , \28084 );
not \U$27833 ( \28086 , RIbe285e8_24);
not \U$27834 ( \28087 , \6958 );
or \U$27835 ( \28088 , \28086 , \28087 );
nand \U$27836 ( \28089 , \8202 , RIbe287c8_28);
nand \U$27837 ( \28090 , \28088 , \28089 );
and \U$27838 ( \28091 , \28090 , \7293 );
not \U$27839 ( \28092 , \28090 );
and \U$27840 ( \28093 , \28092 , \6572 );
nor \U$27841 ( \28094 , \28091 , \28093 );
not \U$27842 ( \28095 , \28094 );
and \U$27843 ( \28096 , \28085 , \28095 );
not \U$27844 ( \28097 , RIbe27fd0_11);
not \U$27845 ( \28098 , \6536 );
or \U$27846 ( \28099 , \28097 , \28098 );
nand \U$27847 ( \28100 , \6540 , RIbe27f58_10);
nand \U$27848 ( \28101 , \28099 , \28100 );
not \U$27849 ( \28102 , \28101 );
not \U$27850 ( \28103 , \6891 );
and \U$27851 ( \28104 , \28102 , \28103 );
and \U$27852 ( \28105 , \28101 , \6548 );
nor \U$27853 ( \28106 , \28104 , \28105 );
nor \U$27854 ( \28107 , \28096 , \28106 );
nor \U$27855 ( \28108 , \28085 , \28095 );
nor \U$27856 ( \28109 , \28107 , \28108 );
and \U$27857 ( \28110 , \28076 , \28109 );
not \U$27858 ( \28111 , RIbe28390_19);
not \U$27859 ( \28112 , \6942 );
or \U$27860 ( \28113 , \28111 , \28112 );
nand \U$27861 ( \28114 , \13339 , RIbe28b10_35);
nand \U$27862 ( \28115 , \28113 , \28114 );
and \U$27863 ( \28116 , \28115 , \7984 );
not \U$27864 ( \28117 , \28115 );
and \U$27865 ( \28118 , \28117 , \7988 );
nor \U$27866 ( \28119 , \28116 , \28118 );
and \U$27867 ( \28120 , \9909 , RIbe28b88_36);
and \U$27868 ( \28121 , \10919 , RIbe29290_51);
nor \U$27869 ( \28122 , \28120 , \28121 );
and \U$27870 ( \28123 , \28122 , \13383 );
not \U$27871 ( \28124 , \28122 );
and \U$27872 ( \28125 , \28124 , \7970 );
nor \U$27873 ( \28126 , \28123 , \28125 );
not \U$27874 ( \28127 , \28126 );
nand \U$27875 ( \28128 , \28119 , \28127 );
not \U$27876 ( \28129 , \7661 );
not \U$27877 ( \28130 , RIbe28480_21);
not \U$27878 ( \28131 , \6980 );
or \U$27879 ( \28132 , \28130 , \28131 );
nand \U$27880 ( \28133 , \8287 , RIbe28408_20);
nand \U$27881 ( \28134 , \28132 , \28133 );
not \U$27882 ( \28135 , \28134 );
or \U$27883 ( \28136 , \28129 , \28135 );
or \U$27884 ( \28137 , \28134 , \7301 );
nand \U$27885 ( \28138 , \28136 , \28137 );
and \U$27886 ( \28139 , \28128 , \28138 );
nor \U$27887 ( \28140 , \28119 , \28127 );
nor \U$27888 ( \28141 , \28139 , \28140 );
nor \U$27889 ( \28142 , \28110 , \28141 );
nor \U$27890 ( \28143 , \28076 , \28109 );
nor \U$27891 ( \28144 , \28142 , \28143 );
not \U$27892 ( \28145 , \28144 );
not \U$27893 ( \28146 , \12801 );
not \U$27894 ( \28147 , RIbe290b0_47);
not \U$27895 ( \28148 , \15249 );
or \U$27896 ( \28149 , \28147 , \28148 );
nand \U$27897 ( \28150 , \12794 , RIbe29a88_68);
nand \U$27898 ( \28151 , \28149 , \28150 );
not \U$27899 ( \28152 , \28151 );
or \U$27900 ( \28153 , \28146 , \28152 );
or \U$27901 ( \28154 , \28151 , \12893 );
nand \U$27902 ( \28155 , \28153 , \28154 );
not \U$27903 ( \28156 , RIbe27d78_6);
not \U$27904 ( \28157 , \12811 );
or \U$27905 ( \28158 , \28156 , \28157 );
nand \U$27906 ( \28159 , RIbe27d00_5, RIbe2ae38_110);
nand \U$27907 ( \28160 , \28158 , \28159 );
xnor \U$27908 ( \28161 , \28160 , RIbe2aeb0_111);
nand \U$27909 ( \28162 , \28161 , \300 );
and \U$27910 ( \28163 , \28155 , \28162 );
nor \U$27911 ( \28164 , \28161 , \300 );
nor \U$27912 ( \28165 , \28163 , \28164 );
not \U$27913 ( \28166 , RIbe29038_46);
not \U$27914 ( \28167 , \14550 );
or \U$27915 ( \28168 , \28166 , \28167 );
nand \U$27916 ( \28169 , \12834 , RIbe28fc0_45);
nand \U$27917 ( \28170 , \28168 , \28169 );
and \U$27918 ( \28171 , \28170 , \16366 );
not \U$27919 ( \28172 , \28170 );
and \U$27920 ( \28173 , \28172 , \20602 );
nor \U$27921 ( \28174 , \28171 , \28173 );
not \U$27922 ( \28175 , RIbe280c0_13);
not \U$27923 ( \28176 , \19262 );
or \U$27924 ( \28177 , \28175 , \28176 );
nand \U$27925 ( \28178 , \12711 , RIbe29830_63);
nand \U$27926 ( \28179 , \28177 , \28178 );
and \U$27927 ( \28180 , \28179 , \12723 );
not \U$27928 ( \28181 , \28179 );
and \U$27929 ( \28182 , \28181 , \12716 );
nor \U$27930 ( \28183 , \28180 , \28182 );
nand \U$27931 ( \28184 , \28174 , \28183 );
not \U$27932 ( \28185 , RIbe296c8_60);
not \U$27933 ( \28186 , \15161 );
or \U$27934 ( \28187 , \28185 , \28186 );
nand \U$27935 ( \28188 , \12735 , RIbe29650_59);
nand \U$27936 ( \28189 , \28187 , \28188 );
and \U$27937 ( \28190 , \28189 , \14077 );
not \U$27938 ( \28191 , \28189 );
and \U$27939 ( \28192 , \28191 , \15169 );
nor \U$27940 ( \28193 , \28190 , \28192 );
and \U$27941 ( \28194 , \28184 , \28193 );
nor \U$27942 ( \28195 , \28183 , \28174 );
nor \U$27943 ( \28196 , \28194 , \28195 );
and \U$27944 ( \28197 , \28165 , \28196 );
not \U$27945 ( \28198 , RIbe28a20_33);
not \U$27946 ( \28199 , \10936 );
or \U$27947 ( \28200 , \28198 , \28199 );
nand \U$27948 ( \28201 , \12213 , RIbe289a8_32);
nand \U$27949 ( \28202 , \28200 , \28201 );
and \U$27950 ( \28203 , \28202 , \10943 );
not \U$27951 ( \28204 , \28202 );
and \U$27952 ( \28205 , \28204 , \19139 );
nor \U$27953 ( \28206 , \28203 , \28205 );
not \U$27954 ( \28207 , \12752 );
not \U$27955 ( \28208 , \3663 );
and \U$27956 ( \28209 , \28207 , \28208 );
and \U$27957 ( \28210 , \13738 , RIbe28228_16);
nor \U$27958 ( \28211 , \28209 , \28210 );
and \U$27959 ( \28212 , \28211 , \12927 );
not \U$27960 ( \28213 , \28211 );
and \U$27961 ( \28214 , \28213 , \12924 );
nor \U$27962 ( \28215 , \28212 , \28214 );
not \U$27963 ( \28216 , \28215 );
not \U$27964 ( \28217 , \28216 );
nand \U$27965 ( \28218 , \28206 , \28217 );
and \U$27966 ( \28219 , \15205 , RIbe28930_31);
not \U$27967 ( \28220 , RIbe29560_57);
nor \U$27968 ( \28221 , \14397 , \28220 );
nor \U$27969 ( \28222 , \28219 , \28221 );
and \U$27970 ( \28223 , \28222 , \12960 );
not \U$27971 ( \28224 , \28222 );
and \U$27972 ( \28225 , \28224 , \12195 );
nor \U$27973 ( \28226 , \28223 , \28225 );
and \U$27974 ( \28227 , \28218 , \28226 );
nor \U$27975 ( \28228 , \28206 , \28217 );
nor \U$27976 ( \28229 , \28227 , \28228 );
nor \U$27977 ( \28230 , \28197 , \28229 );
nor \U$27978 ( \28231 , \28196 , \28165 );
nor \U$27979 ( \28232 , \28230 , \28231 );
not \U$27980 ( \28233 , \28232 );
and \U$27981 ( \28234 , \28145 , \28233 );
not \U$27982 ( \28235 , \28145 );
and \U$27983 ( \28236 , \28235 , \28232 );
nor \U$27984 ( \28237 , \28234 , \28236 );
not \U$27985 ( \28238 , \28237 );
or \U$27986 ( \28239 , \28044 , \28238 );
or \U$27987 ( \28240 , \28237 , \28043 );
nand \U$27988 ( \28241 , \28239 , \28240 );
nand \U$27989 ( \28242 , \27872 , \27807 );
and \U$27990 ( \28243 , \28242 , \27832 );
nor \U$27991 ( \28244 , \27807 , \27872 );
nor \U$27992 ( \28245 , \28243 , \28244 );
xor \U$27993 ( \28246 , \27945 , \27954 );
xor \U$27994 ( \28247 , \28246 , \27964 );
xor \U$27995 ( \28248 , \27925 , \27914 );
xnor \U$27996 ( \28249 , \28248 , \27905 );
xor \U$27997 ( \28250 , \28247 , \28249 );
xor \U$27998 ( \28251 , \27499 , \27508 );
xor \U$27999 ( \28252 , \28251 , \27518 );
and \U$28000 ( \28253 , \28250 , \28252 );
and \U$28001 ( \28254 , \28247 , \28249 );
or \U$28002 ( \28255 , \28253 , \28254 );
not \U$28003 ( \28256 , \27697 );
and \U$28004 ( \28257 , \28256 , \27732 );
nor \U$28005 ( \28258 , \28257 , \27768 );
nor \U$28006 ( \28259 , \27732 , \28256 );
nor \U$28007 ( \28260 , \28258 , \28259 );
not \U$28008 ( \28261 , \28260 );
and \U$28009 ( \28262 , \28255 , \28261 );
not \U$28010 ( \28263 , \28255 );
and \U$28011 ( \28264 , \28263 , \28260 );
nor \U$28012 ( \28265 , \28262 , \28264 );
xnor \U$28013 ( \28266 , \28245 , \28265 );
xor \U$28014 ( \28267 , \28241 , \28266 );
not \U$28015 ( \28268 , \1362 );
not \U$28016 ( \28269 , RIbe27c10_3);
not \U$28017 ( \28270 , \13690 );
or \U$28018 ( \28271 , \28269 , \28270 );
nand \U$28019 ( \28272 , RIbe28e58_42, RIbe2ae38_110);
nand \U$28020 ( \28273 , \28271 , \28272 );
xnor \U$28021 ( \28274 , \28273 , RIbe2aeb0_111);
not \U$28022 ( \28275 , \28274 );
not \U$28023 ( \28276 , \28275 );
or \U$28024 ( \28277 , \28268 , \28276 );
or \U$28025 ( \28278 , \28275 , \270 );
nand \U$28026 ( \28279 , \28277 , \28278 );
not \U$28027 ( \28280 , \28279 );
not \U$28028 ( \28281 , RIbe27d78_6);
not \U$28029 ( \28282 , \12787 );
or \U$28030 ( \28283 , \28281 , \28282 );
nand \U$28031 ( \28284 , \12890 , RIbe27d00_5);
nand \U$28032 ( \28285 , \28283 , \28284 );
and \U$28033 ( \28286 , \28285 , \14103 );
not \U$28034 ( \28287 , \28285 );
and \U$28035 ( \28288 , \28287 , \12893 );
nor \U$28036 ( \28289 , \28286 , \28288 );
not \U$28037 ( \28290 , \28289 );
not \U$28038 ( \28291 , \28290 );
or \U$28039 ( \28292 , \28280 , \28291 );
or \U$28040 ( \28293 , \28279 , \28290 );
nand \U$28041 ( \28294 , \28292 , \28293 );
not \U$28042 ( \28295 , RIbe296c8_60);
not \U$28043 ( \28296 , \14523 );
or \U$28044 ( \28297 , \28295 , \28296 );
nand \U$28045 ( \28298 , \12711 , RIbe29650_59);
nand \U$28046 ( \28299 , \28297 , \28298 );
and \U$28047 ( \28300 , \28299 , \12716 );
not \U$28048 ( \28301 , \28299 );
and \U$28049 ( \28302 , \28301 , \13583 );
nor \U$28050 ( \28303 , \28300 , \28302 );
not \U$28051 ( \28304 , RIbe29038_46);
not \U$28052 ( \28305 , \15161 );
or \U$28053 ( \28306 , \28304 , \28305 );
nand \U$28054 ( \28307 , \12735 , RIbe28fc0_45);
nand \U$28055 ( \28308 , \28306 , \28307 );
and \U$28056 ( \28309 , \28308 , \14358 );
not \U$28057 ( \28310 , \28308 );
and \U$28058 ( \28311 , \28310 , \12742 );
nor \U$28059 ( \28312 , \28309 , \28311 );
not \U$28060 ( \28313 , RIbe290b0_47);
not \U$28061 ( \28314 , \12858 );
or \U$28062 ( \28315 , \28313 , \28314 );
nand \U$28063 ( \28316 , \13012 , RIbe29a88_68);
nand \U$28064 ( \28317 , \28315 , \28316 );
and \U$28065 ( \28318 , \28317 , \12863 );
not \U$28066 ( \28319 , \28317 );
and \U$28067 ( \28320 , \28319 , \18364 );
nor \U$28068 ( \28321 , \28318 , \28320 );
and \U$28069 ( \28322 , \28312 , \28321 );
not \U$28070 ( \28323 , \28312 );
not \U$28071 ( \28324 , \28321 );
and \U$28072 ( \28325 , \28323 , \28324 );
or \U$28073 ( \28326 , \28322 , \28325 );
xor \U$28074 ( \28327 , \28303 , \28326 );
xor \U$28075 ( \28328 , \28294 , \28327 );
not \U$28076 ( \28329 , \12752 );
not \U$28077 ( \28330 , RIbe29830_63);
not \U$28078 ( \28331 , \28330 );
and \U$28079 ( \28332 , \28329 , \28331 );
and \U$28080 ( \28333 , \13738 , RIbe280c0_13);
nor \U$28081 ( \28334 , \28332 , \28333 );
and \U$28082 ( \28335 , \28334 , \26172 );
not \U$28083 ( \28336 , \28334 );
and \U$28084 ( \28337 , \28336 , \12927 );
nor \U$28085 ( \28338 , \28335 , \28337 );
not \U$28086 ( \28339 , RIbe28228_16);
not \U$28087 ( \28340 , \12942 );
or \U$28088 ( \28341 , \28339 , \28340 );
nand \U$28089 ( \28342 , \13669 , RIbe281b0_15);
nand \U$28090 ( \28343 , \28341 , \28342 );
and \U$28091 ( \28344 , \28343 , \12195 );
not \U$28092 ( \28345 , \28343 );
and \U$28093 ( \28346 , \28345 , \17005 );
nor \U$28094 ( \28347 , \28344 , \28346 );
xor \U$28095 ( \28348 , \28338 , \28347 );
not \U$28096 ( \28349 , \10940 );
not \U$28097 ( \28350 , RIbe28930_31);
not \U$28098 ( \28351 , \13024 );
or \U$28099 ( \28352 , \28350 , \28351 );
nand \U$28100 ( \28353 , \14511 , RIbe29560_57);
nand \U$28101 ( \28354 , \28352 , \28353 );
not \U$28102 ( \28355 , \28354 );
or \U$28103 ( \28356 , \28349 , \28355 );
or \U$28104 ( \28357 , \28354 , \13661 );
nand \U$28105 ( \28358 , \28356 , \28357 );
xor \U$28106 ( \28359 , \28348 , \28358 );
xor \U$28107 ( \28360 , \28328 , \28359 );
not \U$28108 ( \28361 , RIbe2b108_116);
not \U$28109 ( \28362 , \6747 );
or \U$28110 ( \28363 , \28361 , \28362 );
nand \U$28111 ( \28364 , \1165 , RIbe2b090_115);
nand \U$28112 ( \28365 , \28363 , \28364 );
and \U$28113 ( \28366 , \28365 , \1011 );
not \U$28114 ( \28367 , \28365 );
and \U$28115 ( \28368 , \28367 , \1608 );
nor \U$28116 ( \28369 , \28366 , \28368 );
not \U$28117 ( \28370 , RIbe2a280_85);
not \U$28118 ( \28371 , \2597 );
or \U$28119 ( \28372 , \28370 , \28371 );
nand \U$28120 ( \28373 , \1147 , RIbe2a208_84);
nand \U$28121 ( \28374 , \28372 , \28373 );
and \U$28122 ( \28375 , \28374 , \7899 );
not \U$28123 ( \28376 , \28374 );
and \U$28124 ( \28377 , \28376 , \1157 );
nor \U$28125 ( \28378 , \28375 , \28377 );
xor \U$28126 ( \28379 , \28369 , \28378 );
not \U$28127 ( \28380 , RIbe2a190_83);
not \U$28128 ( \28381 , \8868 );
or \U$28129 ( \28382 , \28380 , \28381 );
nand \U$28130 ( \28383 , \1455 , RIbe2a5c8_92);
nand \U$28131 ( \28384 , \28382 , \28383 );
and \U$28132 ( \28385 , \28384 , \1309 );
not \U$28133 ( \28386 , \28384 );
and \U$28134 ( \28387 , \28386 , \4251 );
nor \U$28135 ( \28388 , \28385 , \28387 );
xor \U$28136 ( \28389 , \28379 , \28388 );
not \U$28137 ( \28390 , \3448 );
not \U$28138 ( \28391 , RIbe2a028_80);
not \U$28139 ( \28392 , \6783 );
or \U$28140 ( \28393 , \28391 , \28392 );
nand \U$28141 ( \28394 , \8368 , RIbe29fb0_79);
nand \U$28142 ( \28395 , \28393 , \28394 );
not \U$28143 ( \28396 , \28395 );
or \U$28144 ( \28397 , \28390 , \28396 );
or \U$28145 ( \28398 , \28395 , \3698 );
nand \U$28146 ( \28399 , \28397 , \28398 );
not \U$28147 ( \28400 , RIbe29e48_76);
not \U$28148 ( \28401 , \4317 );
or \U$28149 ( \28402 , \28400 , \28401 );
nand \U$28150 ( \28403 , \7858 , RIbe29dd0_75);
nand \U$28151 ( \28404 , \28402 , \28403 );
xor \U$28152 ( \28405 , \28404 , \4323 );
xor \U$28153 ( \28406 , \28399 , \28405 );
not \U$28154 ( \28407 , RIbe2a2f8_86);
not \U$28155 ( \28408 , \3452 );
or \U$28156 ( \28409 , \28407 , \28408 );
nand \U$28157 ( \28410 , \4011 , RIbe2acd0_107);
nand \U$28158 ( \28411 , \28409 , \28410 );
and \U$28159 ( \28412 , \28411 , \3290 );
not \U$28160 ( \28413 , \28411 );
and \U$28161 ( \28414 , \28413 , \3461 );
nor \U$28162 ( \28415 , \28412 , \28414 );
xnor \U$28163 ( \28416 , \28406 , \28415 );
xor \U$28164 ( \28417 , \28389 , \28416 );
and \U$28165 ( \28418 , \2583 , RIbe2a910_99);
not \U$28166 ( \28419 , RIbe2b5b8_126);
nor \U$28167 ( \28420 , \28419 , \2385 );
nor \U$28168 ( \28421 , \28418 , \28420 );
and \U$28169 ( \28422 , \28421 , \1277 );
not \U$28170 ( \28423 , \28421 );
and \U$28171 ( \28424 , \28423 , \3516 );
nor \U$28172 ( \28425 , \28422 , \28424 );
not \U$28173 ( \28426 , RIbe2a3e8_88);
not \U$28174 ( \28427 , \2898 );
or \U$28175 ( \28428 , \28426 , \28427 );
nand \U$28176 ( \28429 , \4284 , RIbe2a370_87);
nand \U$28177 ( \28430 , \28428 , \28429 );
and \U$28178 ( \28431 , \28430 , \4058 );
not \U$28179 ( \28432 , \28430 );
and \U$28180 ( \28433 , \28432 , \2576 );
nor \U$28181 ( \28434 , \28431 , \28433 );
and \U$28182 ( \28435 , \28425 , \28434 );
not \U$28183 ( \28436 , \28425 );
not \U$28184 ( \28437 , \28434 );
and \U$28185 ( \28438 , \28436 , \28437 );
or \U$28186 ( \28439 , \28435 , \28438 );
and \U$28187 ( \28440 , \6380 , RIbe2a550_91);
and \U$28188 ( \28441 , \5467 , RIbe2a988_100);
nor \U$28189 ( \28442 , \28440 , \28441 );
and \U$28190 ( \28443 , \28442 , \1131 );
not \U$28191 ( \28444 , \28442 );
and \U$28192 ( \28445 , \28444 , \3491 );
nor \U$28193 ( \28446 , \28443 , \28445 );
xnor \U$28194 ( \28447 , \28439 , \28446 );
xor \U$28195 ( \28448 , \28417 , \28447 );
xor \U$28196 ( \28449 , \28360 , \28448 );
and \U$28197 ( \28450 , \21196 , RIbe28a20_33);
and \U$28198 ( \28451 , \9913 , RIbe289a8_32);
nor \U$28199 ( \28452 , \28450 , \28451 );
and \U$28200 ( \28453 , \28452 , \7971 );
not \U$28201 ( \28454 , \28452 );
and \U$28202 ( \28455 , \28454 , \7970 );
nor \U$28203 ( \28456 , \28453 , \28455 );
not \U$28204 ( \28457 , RIbe28b88_36);
not \U$28205 ( \28458 , \7974 );
or \U$28206 ( \28459 , \28457 , \28458 );
nand \U$28207 ( \28460 , \7981 , RIbe29290_51);
nand \U$28208 ( \28461 , \28459 , \28460 );
and \U$28209 ( \28462 , \28461 , \14299 );
not \U$28210 ( \28463 , \28461 );
and \U$28211 ( \28464 , \28463 , \7984 );
nor \U$28212 ( \28465 , \28462 , \28464 );
xor \U$28213 ( \28466 , \28456 , \28465 );
not \U$28214 ( \28467 , RIbe28390_19);
not \U$28215 ( \28468 , \6980 );
or \U$28216 ( \28469 , \28467 , \28468 );
nand \U$28217 ( \28470 , \10898 , RIbe28b10_35);
nand \U$28218 ( \28471 , \28469 , \28470 );
and \U$28219 ( \28472 , \28471 , \13167 );
not \U$28220 ( \28473 , \28471 );
and \U$28221 ( \28474 , \28473 , \6992 );
nor \U$28222 ( \28475 , \28472 , \28474 );
xnor \U$28223 ( \28476 , \28466 , \28475 );
not \U$28224 ( \28477 , \28476 );
not \U$28225 ( \28478 , RIbe28480_21);
not \U$28226 ( \28479 , \21608 );
or \U$28227 ( \28480 , \28478 , \28479 );
nand \U$28228 ( \28481 , \7958 , RIbe28408_20);
nand \U$28229 ( \28482 , \28480 , \28481 );
and \U$28230 ( \28483 , \28482 , \6569 );
not \U$28231 ( \28484 , \28482 );
and \U$28232 ( \28485 , \28484 , \7293 );
nor \U$28233 ( \28486 , \28483 , \28485 );
not \U$28234 ( \28487 , RIbe285e8_24);
not \U$28235 ( \28488 , \6868 );
or \U$28236 ( \28489 , \28487 , \28488 );
nand \U$28237 ( \28490 , \7278 , RIbe287c8_28);
nand \U$28238 ( \28491 , \28489 , \28490 );
and \U$28239 ( \28492 , \28491 , \14666 );
not \U$28240 ( \28493 , \28491 );
and \U$28241 ( \28494 , \28493 , \7948 );
nor \U$28242 ( \28495 , \28492 , \28494 );
xor \U$28243 ( \28496 , \28486 , \28495 );
not \U$28244 ( \28497 , RIbe27e68_8);
not \U$28245 ( \28498 , \6880 );
or \U$28246 ( \28499 , \28497 , \28498 );
nand \U$28247 ( \28500 , \6540 , RIbe28660_25);
nand \U$28248 ( \28501 , \28499 , \28500 );
not \U$28249 ( \28502 , \28501 );
not \U$28250 ( \28503 , \9933 );
and \U$28251 ( \28504 , \28502 , \28503 );
and \U$28252 ( \28505 , \28501 , \6891 );
nor \U$28253 ( \28506 , \28504 , \28505 );
not \U$28254 ( \28507 , \28506 );
and \U$28255 ( \28508 , \28496 , \28507 );
not \U$28256 ( \28509 , \28496 );
and \U$28257 ( \28510 , \28509 , \28506 );
nor \U$28258 ( \28511 , \28508 , \28510 );
not \U$28259 ( \28512 , \28511 );
or \U$28260 ( \28513 , \28477 , \28512 );
or \U$28261 ( \28514 , \28511 , \28476 );
nand \U$28262 ( \28515 , \28513 , \28514 );
not \U$28263 ( \28516 , RIbe27fd0_11);
not \U$28264 ( \28517 , \6139 );
or \U$28265 ( \28518 , \28516 , \28517 );
nand \U$28266 ( \28519 , \6617 , RIbe27f58_10);
nand \U$28267 ( \28520 , \28518 , \28519 );
and \U$28268 ( \28521 , \28520 , \5740 );
not \U$28269 ( \28522 , \28520 );
and \U$28270 ( \28523 , \28522 , \7534 );
nor \U$28271 ( \28524 , \28521 , \28523 );
not \U$28272 ( \28525 , RIbe28f48_44);
not \U$28273 ( \28526 , \15313 );
or \U$28274 ( \28527 , \28525 , \28526 );
nand \U$28275 ( \28528 , \7100 , RIbe28ed0_43);
nand \U$28276 ( \28529 , \28527 , \28528 );
and \U$28277 ( \28530 , \28529 , \5457 );
not \U$28278 ( \28531 , \28529 );
and \U$28279 ( \28532 , \28531 , \10272 );
nor \U$28280 ( \28533 , \28530 , \28532 );
xor \U$28281 ( \28534 , \28524 , \28533 );
not \U$28282 ( \28535 , RIbe29c68_72);
not \U$28283 ( \28536 , \4829 );
or \U$28284 ( \28537 , \28535 , \28536 );
nand \U$28285 ( \28538 , \7056 , RIbe29bf0_71);
nand \U$28286 ( \28539 , \28537 , \28538 );
not \U$28287 ( \28540 , \28539 );
not \U$28288 ( \28541 , \4592 );
and \U$28289 ( \28542 , \28540 , \28541 );
and \U$28290 ( \28543 , \28539 , \4592 );
nor \U$28291 ( \28544 , \28542 , \28543 );
xor \U$28292 ( \28545 , \28534 , \28544 );
not \U$28293 ( \28546 , \28545 );
and \U$28294 ( \28547 , \28515 , \28546 );
not \U$28295 ( \28548 , \28515 );
and \U$28296 ( \28549 , \28548 , \28545 );
nor \U$28297 ( \28550 , \28547 , \28549 );
and \U$28298 ( \28551 , \28449 , \28550 );
not \U$28299 ( \28552 , \28449 );
not \U$28300 ( \28553 , \28550 );
and \U$28301 ( \28554 , \28552 , \28553 );
nor \U$28302 ( \28555 , \28551 , \28554 );
and \U$28303 ( \28556 , \28267 , \28555 );
and \U$28304 ( \28557 , \28241 , \28266 );
or \U$28305 ( \28558 , \28556 , \28557 );
not \U$28306 ( \28559 , RIbe29dd0_75);
not \U$28307 ( \28560 , \15313 );
or \U$28308 ( \28561 , \28559 , \28560 );
nand \U$28309 ( \28562 , \8246 , RIbe29c68_72);
nand \U$28310 ( \28563 , \28561 , \28562 );
and \U$28311 ( \28564 , \28563 , \5754 );
not \U$28312 ( \28565 , \28563 );
and \U$28313 ( \28566 , \28565 , \5045 );
nor \U$28314 ( \28567 , \28564 , \28566 );
not \U$28315 ( \28568 , \28567 );
not \U$28316 ( \28569 , RIbe2acd0_107);
not \U$28317 ( \28570 , \4317 );
or \U$28318 ( \28571 , \28569 , \28570 );
not \U$28319 ( \28572 , \14374 );
nand \U$28320 ( \28573 , \28572 , \7858 );
nand \U$28321 ( \28574 , \28571 , \28573 );
and \U$28322 ( \28575 , \28574 , \4007 );
not \U$28323 ( \28576 , \28574 );
and \U$28324 ( \28577 , \28576 , \7865 );
nor \U$28325 ( \28578 , \28575 , \28577 );
or \U$28326 ( \28579 , \28568 , \28578 );
not \U$28327 ( \28580 , RIbe29fb0_79);
not \U$28328 ( \28581 , \20809 );
or \U$28329 ( \28582 , \28580 , \28581 );
nand \U$28330 ( \28583 , RIbe29e48_76, \5052 );
nand \U$28331 ( \28584 , \28582 , \28583 );
and \U$28332 ( \28585 , \28584 , \4586 );
not \U$28333 ( \28586 , \28584 );
and \U$28334 ( \28587 , \28586 , \20465 );
nor \U$28335 ( \28588 , \28585 , \28587 );
nand \U$28336 ( \28589 , \28579 , \28588 );
nand \U$28337 ( \28590 , \28568 , \28578 );
nand \U$28338 ( \28591 , \28589 , \28590 );
not \U$28339 ( \28592 , RIbe27f58_10);
not \U$28340 ( \28593 , \20487 );
or \U$28341 ( \28594 , \28592 , \28593 );
nand \U$28342 ( \28595 , \7278 , RIbe27e68_8);
nand \U$28343 ( \28596 , \28594 , \28595 );
and \U$28344 ( \28597 , \28596 , \6582 );
not \U$28345 ( \28598 , \28596 );
and \U$28346 ( \28599 , \28598 , \8957 );
nor \U$28347 ( \28600 , \28597 , \28599 );
not \U$28348 ( \28601 , RIbe29bf0_71);
not \U$28349 ( \28602 , \12268 );
or \U$28350 ( \28603 , \28601 , \28602 );
nand \U$28351 ( \28604 , RIbe28f48_44, \7087 );
nand \U$28352 ( \28605 , \28603 , \28604 );
and \U$28353 ( \28606 , \28605 , \6620 );
not \U$28354 ( \28607 , \28605 );
and \U$28355 ( \28608 , \28607 , \7535 );
nor \U$28356 ( \28609 , \28606 , \28608 );
nor \U$28357 ( \28610 , \28600 , \28609 );
not \U$28358 ( \28611 , RIbe28ed0_43);
not \U$28359 ( \28612 , \6535 );
or \U$28360 ( \28613 , \28611 , \28612 );
nand \U$28361 ( \28614 , \6540 , RIbe27fd0_11);
nand \U$28362 ( \28615 , \28613 , \28614 );
not \U$28363 ( \28616 , \28615 );
not \U$28364 ( \28617 , \6888 );
and \U$28365 ( \28618 , \28616 , \28617 );
and \U$28366 ( \28619 , \28615 , \6891 );
nor \U$28367 ( \28620 , \28618 , \28619 );
or \U$28368 ( \28621 , \28610 , \28620 );
nand \U$28369 ( \28622 , \28600 , \28609 );
nand \U$28370 ( \28623 , \28621 , \28622 );
xor \U$28371 ( \28624 , \28591 , \28623 );
not \U$28372 ( \28625 , \6572 );
not \U$28373 ( \28626 , RIbe28660_25);
not \U$28374 ( \28627 , \7954 );
or \U$28375 ( \28628 , \28626 , \28627 );
nand \U$28376 ( \28629 , \8202 , RIbe285e8_24);
nand \U$28377 ( \28630 , \28628 , \28629 );
not \U$28378 ( \28631 , \28630 );
or \U$28379 ( \28632 , \28625 , \28631 );
or \U$28380 ( \28633 , \28630 , \6572 );
nand \U$28381 ( \28634 , \28632 , \28633 );
not \U$28382 ( \28635 , RIbe28408_20);
not \U$28383 ( \28636 , \6942 );
or \U$28384 ( \28637 , \28635 , \28636 );
nand \U$28385 ( \28638 , \9891 , RIbe28390_19);
nand \U$28386 ( \28639 , \28637 , \28638 );
and \U$28387 ( \28640 , \28639 , \6950 );
not \U$28388 ( \28641 , \28639 );
and \U$28389 ( \28642 , \28641 , \6948 );
nor \U$28390 ( \28643 , \28640 , \28642 );
or \U$28391 ( \28644 , \28634 , \28643 );
not \U$28392 ( \28645 , RIbe287c8_28);
not \U$28393 ( \28646 , \6980 );
or \U$28394 ( \28647 , \28645 , \28646 );
nand \U$28395 ( \28648 , \10898 , RIbe28480_21);
nand \U$28396 ( \28649 , \28647 , \28648 );
not \U$28397 ( \28650 , \28649 );
not \U$28398 ( \28651 , \6992 );
and \U$28399 ( \28652 , \28650 , \28651 );
and \U$28400 ( \28653 , \28649 , \10902 );
nor \U$28401 ( \28654 , \28652 , \28653 );
not \U$28402 ( \28655 , \28654 );
nand \U$28403 ( \28656 , \28644 , \28655 );
nand \U$28404 ( \28657 , \28643 , \28634 );
nand \U$28405 ( \28658 , \28656 , \28657 );
and \U$28406 ( \28659 , \28624 , \28658 );
and \U$28407 ( \28660 , \28591 , \28623 );
or \U$28408 ( \28661 , \28659 , \28660 );
not \U$28409 ( \28662 , \28661 );
not \U$28410 ( \28663 , RIbe29290_51);
not \U$28411 ( \28664 , \20530 );
or \U$28412 ( \28665 , \28663 , \28664 );
nand \U$28413 ( \28666 , \12212 , RIbe28a20_33);
nand \U$28414 ( \28667 , \28665 , \28666 );
not \U$28415 ( \28668 , \28667 );
not \U$28416 ( \28669 , \13033 );
and \U$28417 ( \28670 , \28668 , \28669 );
and \U$28418 ( \28671 , \28667 , \10943 );
nor \U$28419 ( \28672 , \28670 , \28671 );
and \U$28420 ( \28673 , \20405 , RIbe28b10_35);
and \U$28421 ( \28674 , \13038 , RIbe28b88_36);
nor \U$28422 ( \28675 , \28673 , \28674 );
and \U$28423 ( \28676 , \28675 , \10926 );
not \U$28424 ( \28677 , \28675 );
and \U$28425 ( \28678 , \28677 , \13383 );
nor \U$28426 ( \28679 , \28676 , \28678 );
nand \U$28427 ( \28680 , \28672 , \28679 );
not \U$28428 ( \28681 , \15627 );
not \U$28429 ( \28682 , \9078 );
and \U$28430 ( \28683 , \28681 , \28682 );
and \U$28431 ( \28684 , \12942 , RIbe289a8_32);
nor \U$28432 ( \28685 , \28683 , \28684 );
and \U$28433 ( \28686 , \28685 , \12956 );
not \U$28434 ( \28687 , \28685 );
and \U$28435 ( \28688 , \28687 , \12195 );
nor \U$28436 ( \28689 , \28686 , \28688 );
and \U$28437 ( \28690 , \28680 , \28689 );
nor \U$28438 ( \28691 , \28672 , \28679 );
nor \U$28439 ( \28692 , \28690 , \28691 );
not \U$28440 ( \28693 , \28692 );
not \U$28441 ( \28694 , RIbe29a88_68);
not \U$28442 ( \28695 , \13003 );
or \U$28443 ( \28696 , \28694 , \28695 );
nand \U$28444 ( \28697 , RIbe27d78_6, RIbe2ae38_110);
nand \U$28445 ( \28698 , \28696 , \28697 );
xnor \U$28446 ( \28699 , \28698 , RIbe2aeb0_111);
not \U$28447 ( \28700 , RIbe28fc0_45);
not \U$28448 ( \28701 , \15249 );
or \U$28449 ( \28702 , \28700 , \28701 );
nand \U$28450 ( \28703 , \12794 , RIbe290b0_47);
nand \U$28451 ( \28704 , \28702 , \28703 );
not \U$28452 ( \28705 , \28704 );
not \U$28453 ( \28706 , \12801 );
and \U$28454 ( \28707 , \28705 , \28706 );
and \U$28455 ( \28708 , \28704 , \12893 );
nor \U$28456 ( \28709 , \28707 , \28708 );
xor \U$28457 ( \28710 , \28699 , \28709 );
not \U$28458 ( \28711 , RIbe29650_59);
not \U$28459 ( \28712 , \13010 );
or \U$28460 ( \28713 , \28711 , \28712 );
nand \U$28461 ( \28714 , \12835 , RIbe29038_46);
nand \U$28462 ( \28715 , \28713 , \28714 );
not \U$28463 ( \28716 , \28715 );
not \U$28464 ( \28717 , \12823 );
and \U$28465 ( \28718 , \28716 , \28717 );
and \U$28466 ( \28719 , \28715 , \12863 );
nor \U$28467 ( \28720 , \28718 , \28719 );
and \U$28468 ( \28721 , \28710 , \28720 );
and \U$28469 ( \28722 , \28699 , \28709 );
or \U$28470 ( \28723 , \28721 , \28722 );
not \U$28471 ( \28724 , \28723 );
or \U$28472 ( \28725 , \28693 , \28724 );
not \U$28473 ( \28726 , RIbe281b0_15);
not \U$28474 ( \28727 , \16759 );
or \U$28475 ( \28728 , \28726 , \28727 );
nand \U$28476 ( \28729 , RIbe280c0_13, \13727 );
nand \U$28477 ( \28730 , \28728 , \28729 );
xnor \U$28478 ( \28731 , \28730 , \12723 );
not \U$28479 ( \28732 , RIbe29830_63);
not \U$28480 ( \28733 , \14534 );
or \U$28481 ( \28734 , \28732 , \28733 );
nand \U$28482 ( \28735 , RIbe296c8_60, \12735 );
nand \U$28483 ( \28736 , \28734 , \28735 );
and \U$28484 ( \28737 , \28736 , \21013 );
not \U$28485 ( \28738 , \28736 );
and \U$28486 ( \28739 , \28738 , \14542 );
nor \U$28487 ( \28740 , \28737 , \28739 );
or \U$28488 ( \28741 , \28731 , \28740 );
not \U$28489 ( \28742 , \12751 );
not \U$28490 ( \28743 , \3952 );
and \U$28491 ( \28744 , \28742 , \28743 );
and \U$28492 ( \28745 , \12921 , RIbe29560_57);
nor \U$28493 ( \28746 , \28744 , \28745 );
and \U$28494 ( \28747 , \28746 , \26172 );
not \U$28495 ( \28748 , \28746 );
and \U$28496 ( \28749 , \28748 , \12927 );
nor \U$28497 ( \28750 , \28747 , \28749 );
and \U$28498 ( \28751 , \28741 , \28750 );
and \U$28499 ( \28752 , \28740 , \28731 );
nor \U$28500 ( \28753 , \28751 , \28752 );
not \U$28501 ( \28754 , \28753 );
nand \U$28502 ( \28755 , \28725 , \28754 );
or \U$28503 ( \28756 , \28723 , \28692 );
nand \U$28504 ( \28757 , \28755 , \28756 );
not \U$28505 ( \28758 , \28757 );
or \U$28506 ( \28759 , \28662 , \28758 );
or \U$28507 ( \28760 , \28757 , \28661 );
not \U$28508 ( \28761 , RIbe2b090_115);
not \U$28509 ( \28762 , \1094 );
or \U$28510 ( \28763 , \28761 , \28762 );
nand \U$28511 ( \28764 , \1455 , RIbe2a280_85);
nand \U$28512 ( \28765 , \28763 , \28764 );
and \U$28513 ( \28766 , \28765 , \1309 );
not \U$28514 ( \28767 , \28765 );
and \U$28515 ( \28768 , \28767 , \5125 );
nor \U$28516 ( \28769 , \28766 , \28768 );
not \U$28517 ( \28770 , RIbe2a208_84);
not \U$28518 ( \28771 , \23509 );
or \U$28519 ( \28772 , \28770 , \28771 );
not \U$28520 ( \28773 , \14285 );
nand \U$28521 ( \28774 , \28773 , \5467 );
nand \U$28522 ( \28775 , \28772 , \28774 );
and \U$28523 ( \28776 , \28775 , \1131 );
not \U$28524 ( \28777 , \28775 );
and \U$28525 ( \28778 , \28777 , \1125 );
nor \U$28526 ( \28779 , \28776 , \28778 );
or \U$28527 ( \28780 , \28769 , \28779 );
not \U$28528 ( \28781 , RIbe2a5c8_92);
not \U$28529 ( \28782 , \20674 );
or \U$28530 ( \28783 , \28781 , \28782 );
nand \U$28531 ( \28784 , \2384 , RIbe2a550_91);
nand \U$28532 ( \28785 , \28783 , \28784 );
not \U$28533 ( \28786 , \28785 );
not \U$28534 ( \28787 , \3516 );
and \U$28535 ( \28788 , \28786 , \28787 );
and \U$28536 ( \28789 , \28785 , \1076 );
nor \U$28537 ( \28790 , \28788 , \28789 );
not \U$28538 ( \28791 , \28790 );
nand \U$28539 ( \28792 , \28780 , \28791 );
nand \U$28540 ( \28793 , \28769 , \28779 );
nand \U$28541 ( \28794 , \28792 , \28793 );
not \U$28542 ( \28795 , \28794 );
not \U$28543 ( \28796 , RIbe2a988_100);
not \U$28544 ( \28797 , \8342 );
or \U$28545 ( \28798 , \28796 , \28797 );
nand \U$28546 ( \28799 , \3267 , RIbe2a910_99);
nand \U$28547 ( \28800 , \28798 , \28799 );
and \U$28548 ( \28801 , \28800 , \2576 );
not \U$28549 ( \28802 , \28800 );
and \U$28550 ( \28803 , \28802 , \2380 );
nor \U$28551 ( \28804 , \28801 , \28803 );
not \U$28552 ( \28805 , RIbe2a370_87);
not \U$28553 ( \28806 , \4021 );
or \U$28554 ( \28807 , \28805 , \28806 );
nand \U$28555 ( \28808 , \4027 , RIbe2a2f8_86);
nand \U$28556 ( \28809 , \28807 , \28808 );
and \U$28557 ( \28810 , \28809 , \3471 );
not \U$28558 ( \28811 , \28809 );
and \U$28559 ( \28812 , \28811 , \3448 );
nor \U$28560 ( \28813 , \28810 , \28812 );
not \U$28561 ( \28814 , \28813 );
nand \U$28562 ( \28815 , \28804 , \28814 );
not \U$28563 ( \28816 , RIbe2b5b8_126);
not \U$28564 ( \28817 , \3451 );
or \U$28565 ( \28818 , \28816 , \28817 );
nand \U$28566 ( \28819 , \4011 , RIbe2a3e8_88);
nand \U$28567 ( \28820 , \28818 , \28819 );
and \U$28568 ( \28821 , \28820 , \3461 );
not \U$28569 ( \28822 , \28820 );
and \U$28570 ( \28823 , \28822 , \4346 );
nor \U$28571 ( \28824 , \28821 , \28823 );
not \U$28572 ( \28825 , \28824 );
and \U$28573 ( \28826 , \28815 , \28825 );
not \U$28574 ( \28827 , \28813 );
nor \U$28575 ( \28828 , \28827 , \28804 );
nor \U$28576 ( \28829 , \28826 , \28828 );
not \U$28577 ( \28830 , \28829 );
not \U$28578 ( \28831 , \28830 );
or \U$28579 ( \28832 , \28795 , \28831 );
not \U$28580 ( \28833 , \28794 );
not \U$28581 ( \28834 , \28833 );
not \U$28582 ( \28835 , \28829 );
or \U$28583 ( \28836 , \28834 , \28835 );
not \U$28584 ( \28837 , RIbe2b270_119);
not \U$28585 ( \28838 , \2597 );
or \U$28586 ( \28839 , \28837 , \28838 );
nand \U$28587 ( \28840 , \1147 , RIbe2b108_116);
nand \U$28588 ( \28841 , \28839 , \28840 );
and \U$28589 ( \28842 , \28841 , \1652 );
not \U$28590 ( \28843 , \28841 );
and \U$28591 ( \28844 , \28843 , \1152 );
nor \U$28592 ( \28845 , \28842 , \28844 );
not \U$28593 ( \28846 , \28845 );
not \U$28594 ( \28847 , \28846 );
and \U$28595 ( \28848 , \1807 , RIbe2b1f8_118);
and \U$28596 ( \28849 , \2000 , RIbe2b180_117);
nor \U$28597 ( \28850 , \28848 , \28849 );
and \U$28598 ( \28851 , \28850 , \1813 );
not \U$28599 ( \28852 , \28850 );
and \U$28600 ( \28853 , \28852 , \1011 );
nor \U$28601 ( \28854 , \28851 , \28853 );
not \U$28602 ( \28855 , \28854 );
not \U$28603 ( \28856 , \28855 );
or \U$28604 ( \28857 , \28847 , \28856 );
not \U$28605 ( \28858 , RIbe2afa0_113);
not \U$28606 ( \28859 , \6350 );
or \U$28607 ( \28860 , \28858 , \28859 );
nand \U$28608 ( \28861 , \740 , RIbe2af28_112);
nand \U$28609 ( \28862 , \28860 , \28861 );
not \U$28610 ( \28863 , \28862 );
not \U$28611 ( \28864 , \564 );
and \U$28612 ( \28865 , \28863 , \28864 );
and \U$28613 ( \28866 , \28862 , \4217 );
nor \U$28614 ( \28867 , \28865 , \28866 );
not \U$28615 ( \28868 , \28867 );
nand \U$28616 ( \28869 , \28857 , \28868 );
nand \U$28617 ( \28870 , \28854 , \28845 );
nand \U$28618 ( \28871 , \28869 , \28870 );
nand \U$28619 ( \28872 , \28836 , \28871 );
nand \U$28620 ( \28873 , \28832 , \28872 );
nand \U$28621 ( \28874 , \28760 , \28873 );
nand \U$28622 ( \28875 , \28759 , \28874 );
xor \U$28623 ( \28876 , \28247 , \28249 );
xor \U$28624 ( \28877 , \28876 , \28252 );
not \U$28625 ( \28878 , \28877 );
xor \U$28626 ( \28879 , \27470 , \27479 );
xor \U$28627 ( \28880 , \28879 , \27489 );
not \U$28628 ( \28881 , \28880 );
xor \U$28629 ( \28882 , \27528 , \27539 );
xnor \U$28630 ( \28883 , \28882 , \27552 );
nand \U$28631 ( \28884 , \28881 , \28883 );
not \U$28632 ( \28885 , \28884 );
or \U$28633 ( \28886 , \28878 , \28885 );
not \U$28634 ( \28887 , \28883 );
nand \U$28635 ( \28888 , \28887 , \28880 );
nand \U$28636 ( \28889 , \28886 , \28888 );
xor \U$28637 ( \28890 , \28875 , \28889 );
not \U$28638 ( \28891 , \27567 );
not \U$28639 ( \28892 , \27577 );
not \U$28640 ( \28893 , \27587 );
or \U$28641 ( \28894 , \28892 , \28893 );
or \U$28642 ( \28895 , \27587 , \27577 );
nand \U$28643 ( \28896 , \28894 , \28895 );
not \U$28644 ( \28897 , \28896 );
or \U$28645 ( \28898 , \28891 , \28897 );
or \U$28646 ( \28899 , \28896 , \27567 );
nand \U$28647 ( \28900 , \28898 , \28899 );
xor \U$28648 ( \28901 , \28063 , \28073 );
xor \U$28649 ( \28902 , \28901 , \28053 );
xor \U$28650 ( \28903 , \28900 , \28902 );
not \U$28651 ( \28904 , \27621 );
not \U$28652 ( \28905 , \27600 );
or \U$28653 ( \28906 , \28904 , \28905 );
not \U$28654 ( \28907 , \27600 );
nand \U$28655 ( \28908 , \28907 , \27620 );
nand \U$28656 ( \28909 , \28906 , \28908 );
buf \U$28657 ( \28910 , \27608 );
not \U$28658 ( \28911 , \28910 );
and \U$28659 ( \28912 , \28909 , \28911 );
not \U$28660 ( \28913 , \28909 );
and \U$28661 ( \28914 , \28913 , \28910 );
nor \U$28662 ( \28915 , \28912 , \28914 );
and \U$28663 ( \28916 , \28903 , \28915 );
and \U$28664 ( \28917 , \28900 , \28902 );
or \U$28665 ( \28918 , \28916 , \28917 );
not \U$28666 ( \28919 , \28918 );
not \U$28667 ( \28920 , \28095 );
not \U$28668 ( \28921 , \28085 );
not \U$28669 ( \28922 , \28921 );
or \U$28670 ( \28923 , \28920 , \28922 );
nand \U$28671 ( \28924 , \28094 , \28085 );
nand \U$28672 ( \28925 , \28923 , \28924 );
xor \U$28673 ( \28926 , \28925 , \28106 );
not \U$28674 ( \28927 , \28926 );
xnor \U$28675 ( \28928 , \28126 , \28119 );
xnor \U$28676 ( \28929 , \28928 , \28138 );
not \U$28677 ( \28930 , \28929 );
or \U$28678 ( \28931 , \28927 , \28930 );
and \U$28679 ( \28932 , \28226 , \28215 );
not \U$28680 ( \28933 , \28226 );
and \U$28681 ( \28934 , \28933 , \28216 );
or \U$28682 ( \28935 , \28932 , \28934 );
not \U$28683 ( \28936 , \28206 );
and \U$28684 ( \28937 , \28935 , \28936 );
not \U$28685 ( \28938 , \28935 );
and \U$28686 ( \28939 , \28938 , \28206 );
nor \U$28687 ( \28940 , \28937 , \28939 );
nand \U$28688 ( \28941 , \28931 , \28940 );
not \U$28689 ( \28942 , \28926 );
not \U$28690 ( \28943 , \28929 );
nand \U$28691 ( \28944 , \28942 , \28943 );
nand \U$28692 ( \28945 , \28941 , \28944 );
not \U$28693 ( \28946 , \28945 );
or \U$28694 ( \28947 , \28919 , \28946 );
or \U$28695 ( \28948 , \28945 , \28918 );
nand \U$28696 ( \28949 , \287 , RIbe2ab68_104);
and \U$28697 ( \28950 , \28949 , \300 );
not \U$28698 ( \28951 , \28949 );
and \U$28699 ( \28952 , \28951 , \293 );
nor \U$28700 ( \28953 , \28950 , \28952 );
xor \U$28701 ( \28954 , \27647 , \27658 );
xnor \U$28702 ( \28955 , \28954 , \27638 );
xor \U$28703 ( \28956 , \28953 , \28955 );
xor \U$28704 ( \28957 , \27786 , \27804 );
xor \U$28705 ( \28958 , \28957 , \27795 );
and \U$28706 ( \28959 , \28956 , \28958 );
and \U$28707 ( \28960 , \28953 , \28955 );
or \U$28708 ( \28961 , \28959 , \28960 );
nand \U$28709 ( \28962 , \28948 , \28961 );
nand \U$28710 ( \28963 , \28947 , \28962 );
and \U$28711 ( \28964 , \28890 , \28963 );
and \U$28712 ( \28965 , \28875 , \28889 );
or \U$28713 ( \28966 , \28964 , \28965 );
and \U$28714 ( \28967 , \28558 , \28966 );
not \U$28715 ( \28968 , \28558 );
not \U$28716 ( \28969 , \28966 );
and \U$28717 ( \28970 , \28968 , \28969 );
nor \U$28718 ( \28971 , \28967 , \28970 );
not \U$28719 ( \28972 , \28971 );
or \U$28720 ( \28973 , \28035 , \28972 );
or \U$28721 ( \28974 , \28971 , \28034 );
nand \U$28722 ( \28975 , \28973 , \28974 );
and \U$28723 ( \28976 , \28161 , \293 );
not \U$28724 ( \28977 , \28161 );
and \U$28725 ( \28978 , \28977 , \300 );
or \U$28726 ( \28979 , \28976 , \28978 );
xnor \U$28727 ( \28980 , \28979 , \28155 );
not \U$28728 ( \28981 , \28980 );
not \U$28729 ( \28982 , \28174 );
not \U$28730 ( \28983 , \28193 );
or \U$28731 ( \28984 , \28982 , \28983 );
or \U$28732 ( \28985 , \28193 , \28174 );
nand \U$28733 ( \28986 , \28984 , \28985 );
xnor \U$28734 ( \28987 , \28986 , \28183 );
not \U$28735 ( \28988 , \28987 );
or \U$28736 ( \28989 , \28981 , \28988 );
or \U$28737 ( \28990 , \28987 , \28980 );
nand \U$28738 ( \28991 , \28989 , \28990 );
not \U$28739 ( \28992 , \28991 );
xor \U$28740 ( \28993 , \28740 , \28731 );
xnor \U$28741 ( \28994 , \28993 , \28750 );
not \U$28742 ( \28995 , \28994 );
xor \U$28743 ( \28996 , \28699 , \28709 );
xor \U$28744 ( \28997 , \28996 , \28720 );
not \U$28745 ( \28998 , \28997 );
or \U$28746 ( \28999 , \28995 , \28998 );
xor \U$28747 ( \29000 , \28672 , \28689 );
xor \U$28748 ( \29001 , \29000 , \28679 );
nand \U$28749 ( \29002 , \28999 , \29001 );
not \U$28750 ( \29003 , \28994 );
not \U$28751 ( \29004 , \28997 );
nand \U$28752 ( \29005 , \29003 , \29004 );
and \U$28753 ( \29006 , \29002 , \29005 );
not \U$28754 ( \29007 , \29006 );
or \U$28755 ( \29008 , \28992 , \29007 );
not \U$28756 ( \29009 , \29005 );
not \U$28757 ( \29010 , \29002 );
or \U$28758 ( \29011 , \29009 , \29010 );
not \U$28759 ( \29012 , \28991 );
nand \U$28760 ( \29013 , \29011 , \29012 );
nand \U$28761 ( \29014 , \29008 , \29013 );
not \U$28762 ( \29015 , \29014 );
not \U$28763 ( \29016 , \29015 );
not \U$28764 ( \29017 , \12801 );
not \U$28765 ( \29018 , RIbe29038_46);
not \U$28766 ( \29019 , \13518 );
or \U$28767 ( \29020 , \29018 , \29019 );
nand \U$28768 ( \29021 , \12890 , RIbe28fc0_45);
nand \U$28769 ( \29022 , \29020 , \29021 );
not \U$28770 ( \29023 , \29022 );
or \U$28771 ( \29024 , \29017 , \29023 );
or \U$28772 ( \29025 , \29022 , \12893 );
nand \U$28773 ( \29026 , \29024 , \29025 );
not \U$28774 ( \29027 , RIbe290b0_47);
not \U$28775 ( \29028 , \13003 );
or \U$28776 ( \29029 , \29027 , \29028 );
nand \U$28777 ( \29030 , RIbe29a88_68, RIbe2ae38_110);
nand \U$28778 ( \29031 , \29029 , \29030 );
not \U$28779 ( \29032 , RIbe2aeb0_111);
xor \U$28780 ( \29033 , \29031 , \29032 );
nand \U$28781 ( \29034 , \29033 , \313 );
and \U$28782 ( \29035 , \29026 , \29034 );
nor \U$28783 ( \29036 , \29033 , \1547 );
nor \U$28784 ( \29037 , \29035 , \29036 );
not \U$28785 ( \29038 , \29037 );
not \U$28786 ( \29039 , RIbe28b88_36);
not \U$28787 ( \29040 , \13024 );
or \U$28788 ( \29041 , \29039 , \29040 );
nand \U$28789 ( \29042 , \12971 , RIbe29290_51);
nand \U$28790 ( \29043 , \29041 , \29042 );
not \U$28791 ( \29044 , \29043 );
not \U$28792 ( \29045 , \12218 );
and \U$28793 ( \29046 , \29044 , \29045 );
and \U$28794 ( \29047 , \29043 , \10940 );
nor \U$28795 ( \29048 , \29046 , \29047 );
and \U$28796 ( \29049 , \12920 , RIbe28930_31);
and \U$28797 ( \29050 , \14491 , RIbe29560_57);
nor \U$28798 ( \29051 , \29049 , \29050 );
and \U$28799 ( \29052 , \29051 , \12774 );
not \U$28800 ( \29053 , \29051 );
and \U$28801 ( \29054 , \29053 , \12769 );
nor \U$28802 ( \29055 , \29052 , \29054 );
and \U$28803 ( \29056 , \29048 , \29055 );
not \U$28804 ( \29057 , RIbe28a20_33);
not \U$28805 ( \29058 , \12942 );
or \U$28806 ( \29059 , \29057 , \29058 );
not \U$28807 ( \29060 , \3421 );
nand \U$28808 ( \29061 , \29060 , \12947 );
nand \U$28809 ( \29062 , \29059 , \29061 );
and \U$28810 ( \29063 , \29062 , \12960 );
not \U$28811 ( \29064 , \29062 );
and \U$28812 ( \29065 , \29064 , \12195 );
nor \U$28813 ( \29066 , \29063 , \29065 );
nor \U$28814 ( \29067 , \29056 , \29066 );
nor \U$28815 ( \29068 , \29048 , \29055 );
nor \U$28816 ( \29069 , \29067 , \29068 );
not \U$28817 ( \29070 , \29069 );
or \U$28818 ( \29071 , \29038 , \29070 );
and \U$28819 ( \29072 , \12834 , \5494 );
not \U$28820 ( \29073 , \12834 );
nand \U$28821 ( \29074 , \12828 , RIbe296c8_60);
and \U$28822 ( \29075 , \29073 , \29074 );
or \U$28823 ( \29076 , \29072 , \29075 );
and \U$28824 ( \29077 , \29076 , \20602 );
not \U$28825 ( \29078 , \29076 );
and \U$28826 ( \29079 , \29078 , \16366 );
nor \U$28827 ( \29080 , \29077 , \29079 );
not \U$28828 ( \29081 , \29080 );
not \U$28829 ( \29082 , \12723 );
not \U$28830 ( \29083 , RIbe28228_16);
not \U$28831 ( \29084 , \12707 );
or \U$28832 ( \29085 , \29083 , \29084 );
nand \U$28833 ( \29086 , \13728 , RIbe281b0_15);
nand \U$28834 ( \29087 , \29085 , \29086 );
not \U$28835 ( \29088 , \29087 );
or \U$28836 ( \29089 , \29082 , \29088 );
or \U$28837 ( \29090 , \12706 , \3952 );
not \U$28838 ( \29091 , \12710 );
or \U$28839 ( \29092 , \29091 , \3663 );
nand \U$28840 ( \29093 , \29090 , \29092 , \12716 );
nand \U$28841 ( \29094 , \29089 , \29093 );
not \U$28842 ( \29095 , \29094 );
not \U$28843 ( \29096 , RIbe280c0_13);
not \U$28844 ( \29097 , \15161 );
or \U$28845 ( \29098 , \29096 , \29097 );
nand \U$28846 ( \29099 , \14074 , RIbe29830_63);
nand \U$28847 ( \29100 , \29098 , \29099 );
and \U$28848 ( \29101 , \29100 , \12746 );
not \U$28849 ( \29102 , \29100 );
and \U$28850 ( \29103 , \29102 , \12743 );
nor \U$28851 ( \29104 , \29101 , \29103 );
nand \U$28852 ( \29105 , \29095 , \29104 );
nand \U$28853 ( \29106 , \29081 , \29105 );
not \U$28854 ( \29107 , \29104 );
nand \U$28855 ( \29108 , \29107 , \29094 );
nand \U$28856 ( \29109 , \29106 , \29108 );
nand \U$28857 ( \29110 , \29071 , \29109 );
not \U$28858 ( \29111 , \29069 );
not \U$28859 ( \29112 , \29037 );
nand \U$28860 ( \29113 , \29111 , \29112 );
nand \U$28861 ( \29114 , \29110 , \29113 );
not \U$28862 ( \29115 , \29114 );
not \U$28863 ( \29116 , RIbe27fd0_11);
not \U$28864 ( \29117 , \20487 );
or \U$28865 ( \29118 , \29116 , \29117 );
nand \U$28866 ( \29119 , RIbe27f58_10, \6595 );
nand \U$28867 ( \29120 , \29118 , \29119 );
not \U$28868 ( \29121 , \6582 );
and \U$28869 ( \29122 , \29120 , \29121 );
not \U$28870 ( \29123 , \29120 );
and \U$28871 ( \29124 , \29123 , \7948 );
nor \U$28872 ( \29125 , \29122 , \29124 );
not \U$28873 ( \29126 , RIbe27e68_8);
not \U$28874 ( \29127 , \21608 );
or \U$28875 ( \29128 , \29126 , \29127 );
not \U$28876 ( \29129 , \25899 );
nand \U$28877 ( \29130 , \29129 , \6962 );
nand \U$28878 ( \29131 , \29128 , \29130 );
and \U$28879 ( \29132 , \29131 , \6569 );
not \U$28880 ( \29133 , \29131 );
and \U$28881 ( \29134 , \29133 , \7293 );
nor \U$28882 ( \29135 , \29132 , \29134 );
nand \U$28883 ( \29136 , \29125 , \29135 );
not \U$28884 ( \29137 , \6888 );
not \U$28885 ( \29138 , RIbe28f48_44);
not \U$28886 ( \29139 , \6535 );
or \U$28887 ( \29140 , \29138 , \29139 );
nand \U$28888 ( \29141 , \7075 , RIbe28ed0_43);
nand \U$28889 ( \29142 , \29140 , \29141 );
not \U$28890 ( \29143 , \29142 );
or \U$28891 ( \29144 , \29137 , \29143 );
or \U$28892 ( \29145 , \29142 , \9933 );
nand \U$28893 ( \29146 , \29144 , \29145 );
and \U$28894 ( \29147 , \29136 , \29146 );
nor \U$28895 ( \29148 , \29125 , \29135 );
nor \U$28896 ( \29149 , \29147 , \29148 );
not \U$28897 ( \29150 , \29149 );
not \U$28898 ( \29151 , RIbe29c68_72);
not \U$28899 ( \29152 , \21081 );
or \U$28900 ( \29153 , \29151 , \29152 );
nand \U$28901 ( \29154 , RIbe29bf0_71, \8234 );
nand \U$28902 ( \29155 , \29153 , \29154 );
and \U$28903 ( \29156 , \29155 , \21090 );
not \U$28904 ( \29157 , \29155 );
and \U$28905 ( \29158 , \29157 , \21093 );
nor \U$28906 ( \29159 , \29156 , \29158 );
not \U$28907 ( \29160 , RIbe2a028_80);
not \U$28908 ( \29161 , \20809 );
or \U$28909 ( \29162 , \29160 , \29161 );
nand \U$28910 ( \29163 , \7056 , RIbe29fb0_79);
nand \U$28911 ( \29164 , \29162 , \29163 );
and \U$28912 ( \29165 , \29164 , \20465 );
not \U$28913 ( \29166 , \29164 );
and \U$28914 ( \29167 , \29166 , \4586 );
nor \U$28915 ( \29168 , \29165 , \29167 );
nand \U$28916 ( \29169 , \29159 , \29168 );
not \U$28917 ( \29170 , RIbe29e48_76);
not \U$28918 ( \29171 , \20796 );
or \U$28919 ( \29172 , \29170 , \29171 );
nand \U$28920 ( \29173 , \7099 , RIbe29dd0_75);
nand \U$28921 ( \29174 , \29172 , \29173 );
and \U$28922 ( \29175 , \29174 , \6121 );
not \U$28923 ( \29176 , \29174 );
and \U$28924 ( \29177 , \29176 , \5457 );
nor \U$28925 ( \29178 , \29175 , \29177 );
and \U$28926 ( \29179 , \29169 , \29178 );
nor \U$28927 ( \29180 , \29159 , \29168 );
nor \U$28928 ( \29181 , \29179 , \29180 );
not \U$28929 ( \29182 , \29181 );
or \U$28930 ( \29183 , \29150 , \29182 );
and \U$28931 ( \29184 , \10915 , RIbe28390_19);
and \U$28932 ( \29185 , \13038 , RIbe28b10_35);
nor \U$28933 ( \29186 , \29184 , \29185 );
and \U$28934 ( \29187 , \29186 , \15233 );
not \U$28935 ( \29188 , \29186 );
and \U$28936 ( \29189 , \29188 , \13649 );
nor \U$28937 ( \29190 , \29187 , \29189 );
not \U$28938 ( \29191 , \29190 );
not \U$28939 ( \29192 , \29191 );
not \U$28940 ( \29193 , RIbe28480_21);
not \U$28941 ( \29194 , \6942 );
or \U$28942 ( \29195 , \29193 , \29194 );
nand \U$28943 ( \29196 , RIbe28408_20, \13339 );
nand \U$28944 ( \29197 , \29195 , \29196 );
and \U$28945 ( \29198 , \29197 , \7984 );
not \U$28946 ( \29199 , \29197 );
and \U$28947 ( \29200 , \29199 , \6950 );
nor \U$28948 ( \29201 , \29198 , \29200 );
not \U$28949 ( \29202 , \29201 );
or \U$28950 ( \29203 , \29192 , \29202 );
not \U$28951 ( \29204 , \6993 );
and \U$28952 ( \29205 , \7298 , RIbe285e8_24);
and \U$28953 ( \29206 , \13224 , RIbe287c8_28);
nor \U$28954 ( \29207 , \29205 , \29206 );
not \U$28955 ( \29208 , \29207 );
or \U$28956 ( \29209 , \29204 , \29208 );
or \U$28957 ( \29210 , \29207 , \13167 );
nand \U$28958 ( \29211 , \29209 , \29210 );
nand \U$28959 ( \29212 , \29203 , \29211 );
not \U$28960 ( \29213 , \29191 );
not \U$28961 ( \29214 , \29201 );
nand \U$28962 ( \29215 , \29213 , \29214 );
nand \U$28963 ( \29216 , \29212 , \29215 );
nand \U$28964 ( \29217 , \29183 , \29216 );
not \U$28965 ( \29218 , \29181 );
not \U$28966 ( \29219 , \29149 );
nand \U$28967 ( \29220 , \29218 , \29219 );
nand \U$28968 ( \29221 , \29217 , \29220 );
not \U$28969 ( \29222 , \29221 );
not \U$28970 ( \29223 , \29222 );
or \U$28971 ( \29224 , \29115 , \29223 );
not \U$28972 ( \29225 , \29114 );
nand \U$28973 ( \29226 , \29225 , \29221 );
nand \U$28974 ( \29227 , \29224 , \29226 );
not \U$28975 ( \29228 , RIbe2b108_116);
not \U$28976 ( \29229 , \5476 );
or \U$28977 ( \29230 , \29228 , \29229 );
nand \U$28978 ( \29231 , \4730 , RIbe2b090_115);
nand \U$28979 ( \29232 , \29230 , \29231 );
and \U$28980 ( \29233 , \29232 , \2418 );
not \U$28981 ( \29234 , \29232 );
and \U$28982 ( \29235 , \29234 , \1309 );
nor \U$28983 ( \29236 , \29233 , \29235 );
not \U$28984 ( \29237 , RIbe2af28_112);
not \U$28985 ( \29238 , \4858 );
or \U$28986 ( \29239 , \29237 , \29238 );
nand \U$28987 ( \29240 , \7905 , RIbe2b1f8_118);
nand \U$28988 ( \29241 , \29239 , \29240 );
and \U$28989 ( \29242 , \29241 , \1608 );
not \U$28990 ( \29243 , \29241 );
and \U$28991 ( \29244 , \29243 , \1011 );
nor \U$28992 ( \29245 , \29242 , \29244 );
nand \U$28993 ( \29246 , \29236 , \29245 );
not \U$28994 ( \29247 , RIbe2b180_117);
not \U$28995 ( \29248 , \1143 );
or \U$28996 ( \29249 , \29247 , \29248 );
not \U$28997 ( \29250 , \13109 );
nand \U$28998 ( \29251 , \29250 , \1146 );
nand \U$28999 ( \29252 , \29249 , \29251 );
and \U$29000 ( \29253 , \29252 , \1652 );
not \U$29001 ( \29254 , \29252 );
and \U$29002 ( \29255 , \29254 , \1152 );
nor \U$29003 ( \29256 , \29253 , \29255 );
and \U$29004 ( \29257 , \29246 , \29256 );
nor \U$29005 ( \29258 , \29236 , \29245 );
nor \U$29006 ( \29259 , \29257 , \29258 );
not \U$29007 ( \29260 , \29259 );
not \U$29008 ( \29261 , RIbe2a910_99);
not \U$29009 ( \29262 , \6797 );
or \U$29010 ( \29263 , \29261 , \29262 );
nand \U$29011 ( \29264 , \6800 , RIbe2b5b8_126);
nand \U$29012 ( \29265 , \29263 , \29264 );
and \U$29013 ( \29266 , \29265 , \2887 );
not \U$29014 ( \29267 , \29265 );
and \U$29015 ( \29268 , \29267 , \3290 );
nor \U$29016 ( \29269 , \29266 , \29268 );
not \U$29017 ( \29270 , RIbe2a2f8_86);
not \U$29018 ( \29271 , \4595 );
or \U$29019 ( \29272 , \29270 , \29271 );
nand \U$29020 ( \29273 , \21043 , RIbe2acd0_107);
nand \U$29021 ( \29274 , \29272 , \29273 );
not \U$29022 ( \29275 , \29274 );
not \U$29023 ( \29276 , \7865 );
and \U$29024 ( \29277 , \29275 , \29276 );
and \U$29025 ( \29278 , \29274 , \7865 );
nor \U$29026 ( \29279 , \29277 , \29278 );
nand \U$29027 ( \29280 , \29269 , \29279 );
not \U$29028 ( \29281 , RIbe2a3e8_88);
not \U$29029 ( \29282 , \20764 );
or \U$29030 ( \29283 , \29281 , \29282 );
nand \U$29031 ( \29284 , RIbe2a370_87, \6787 );
nand \U$29032 ( \29285 , \29283 , \29284 );
and \U$29033 ( \29286 , \29285 , \3471 );
not \U$29034 ( \29287 , \29285 );
and \U$29035 ( \29288 , \29287 , \3698 );
nor \U$29036 ( \29289 , \29286 , \29288 );
buf \U$29037 ( \29290 , \29289 );
and \U$29038 ( \29291 , \29280 , \29290 );
nor \U$29039 ( \29292 , \29269 , \29279 );
nor \U$29040 ( \29293 , \29291 , \29292 );
not \U$29041 ( \29294 , \29293 );
or \U$29042 ( \29295 , \29260 , \29294 );
not \U$29043 ( \29296 , RIbe2a550_91);
not \U$29044 ( \29297 , \4050 );
or \U$29045 ( \29298 , \29296 , \29297 );
nand \U$29046 ( \29299 , \2900 , RIbe2a988_100);
nand \U$29047 ( \29300 , \29298 , \29299 );
and \U$29048 ( \29301 , \29300 , \2380 );
not \U$29049 ( \29302 , \29300 );
and \U$29050 ( \29303 , \29302 , \2576 );
nor \U$29051 ( \29304 , \29301 , \29303 );
not \U$29052 ( \29305 , \29304 );
not \U$29053 ( \29306 , RIbe2a280_85);
not \U$29054 ( \29307 , \6380 );
or \U$29055 ( \29308 , \29306 , \29307 );
nand \U$29056 ( \29309 , \1117 , RIbe2a208_84);
nand \U$29057 ( \29310 , \29308 , \29309 );
and \U$29058 ( \29311 , \29310 , \1448 );
not \U$29059 ( \29312 , \29310 );
and \U$29060 ( \29313 , \29312 , \1131 );
nor \U$29061 ( \29314 , \29311 , \29313 );
not \U$29062 ( \29315 , \29314 );
not \U$29063 ( \29316 , \29315 );
or \U$29064 ( \29317 , \29305 , \29316 );
not \U$29065 ( \29318 , \29304 );
not \U$29066 ( \29319 , \29318 );
not \U$29067 ( \29320 , \29314 );
or \U$29068 ( \29321 , \29319 , \29320 );
not \U$29069 ( \29322 , RIbe2a190_83);
not \U$29070 ( \29323 , \2390 );
or \U$29071 ( \29324 , \29322 , \29323 );
nand \U$29072 ( \29325 , \2384 , RIbe2a5c8_92);
nand \U$29073 ( \29326 , \29324 , \29325 );
not \U$29074 ( \29327 , \29326 );
not \U$29075 ( \29328 , \1076 );
and \U$29076 ( \29329 , \29327 , \29328 );
and \U$29077 ( \29330 , \29326 , \7038 );
nor \U$29078 ( \29331 , \29329 , \29330 );
not \U$29079 ( \29332 , \29331 );
nand \U$29080 ( \29333 , \29321 , \29332 );
nand \U$29081 ( \29334 , \29317 , \29333 );
nand \U$29082 ( \29335 , \29295 , \29334 );
not \U$29083 ( \29336 , \29259 );
not \U$29084 ( \29337 , \29293 );
nand \U$29085 ( \29338 , \29336 , \29337 );
nand \U$29086 ( \29339 , \29335 , \29338 );
not \U$29087 ( \29340 , \29339 );
and \U$29088 ( \29341 , \29227 , \29340 );
not \U$29089 ( \29342 , \29227 );
and \U$29090 ( \29343 , \29342 , \29339 );
nor \U$29091 ( \29344 , \29341 , \29343 );
not \U$29092 ( \29345 , \29344 );
or \U$29093 ( \29346 , \29016 , \29345 );
not \U$29094 ( \29347 , RIbe2b630_127);
not \U$29095 ( \29348 , \1237 );
or \U$29096 ( \29349 , \29347 , \29348 );
nand \U$29097 ( \29350 , \552 , RIbe2b018_114);
nand \U$29098 ( \29351 , \29349 , \29350 );
and \U$29099 ( \29352 , \29351 , \1761 );
not \U$29100 ( \29353 , \29351 );
and \U$29101 ( \29354 , \29353 , \424 );
nor \U$29102 ( \29355 , \29352 , \29354 );
not \U$29103 ( \29356 , \29355 );
not \U$29104 ( \29357 , RIbe2ab68_104);
not \U$29105 ( \29358 , \1337 );
or \U$29106 ( \29359 , \29357 , \29358 );
nand \U$29107 ( \29360 , \429 , RIbe2aaf0_103);
nand \U$29108 ( \29361 , \29359 , \29360 );
and \U$29109 ( \29362 , \29361 , \313 );
not \U$29110 ( \29363 , \29361 );
and \U$29111 ( \29364 , \29363 , \306 );
nor \U$29112 ( \29365 , \29362 , \29364 );
not \U$29113 ( \29366 , \29365 );
not \U$29114 ( \29367 , \29366 );
or \U$29115 ( \29368 , \29356 , \29367 );
not \U$29116 ( \29369 , RIbe2aaf0_103);
not \U$29117 ( \29370 , \546 );
or \U$29118 ( \29371 , \29369 , \29370 );
nand \U$29119 ( \29372 , \553 , RIbe2b630_127);
nand \U$29120 ( \29373 , \29371 , \29372 );
not \U$29121 ( \29374 , \29373 );
not \U$29122 ( \29375 , \424 );
and \U$29123 ( \29376 , \29374 , \29375 );
and \U$29124 ( \29377 , \29373 , \424 );
nor \U$29125 ( \29378 , \29376 , \29377 );
nand \U$29126 ( \29379 , \429 , RIbe2ab68_104);
and \U$29127 ( \29380 , \29379 , \306 );
not \U$29128 ( \29381 , \29379 );
and \U$29129 ( \29382 , \29381 , \1232 );
nor \U$29130 ( \29383 , \29380 , \29382 );
and \U$29131 ( \29384 , \29378 , \29383 );
not \U$29132 ( \29385 , \4217 );
not \U$29133 ( \29386 , RIbe2b018_114);
or \U$29134 ( \29387 , \562 , RIbe28c00_37);
nand \U$29135 ( \29388 , \29387 , \662 );
not \U$29136 ( \29389 , \29388 );
or \U$29137 ( \29390 , \29386 , \29389 );
nand \U$29138 ( \29391 , \1179 , RIbe2afa0_113);
nand \U$29139 ( \29392 , \29390 , \29391 );
not \U$29140 ( \29393 , \29392 );
or \U$29141 ( \29394 , \29385 , \29393 );
or \U$29142 ( \29395 , \29392 , \1618 );
nand \U$29143 ( \29396 , \29394 , \29395 );
not \U$29144 ( \29397 , \29396 );
nor \U$29145 ( \29398 , \29384 , \29397 );
nor \U$29146 ( \29399 , \29378 , \29383 );
or \U$29147 ( \29400 , \29398 , \29399 );
not \U$29148 ( \29401 , \29355 );
nand \U$29149 ( \29402 , \29365 , \29401 );
nand \U$29150 ( \29403 , \29400 , \29402 );
nand \U$29151 ( \29404 , \29368 , \29403 );
xor \U$29152 ( \29405 , \28790 , \28779 );
xnor \U$29153 ( \29406 , \29405 , \28769 );
not \U$29154 ( \29407 , \29406 );
not \U$29155 ( \29408 , \28814 );
not \U$29156 ( \29409 , \28825 );
or \U$29157 ( \29410 , \29408 , \29409 );
nand \U$29158 ( \29411 , \28824 , \28813 );
nand \U$29159 ( \29412 , \29410 , \29411 );
not \U$29160 ( \29413 , \28804 );
and \U$29161 ( \29414 , \29412 , \29413 );
not \U$29162 ( \29415 , \29412 );
and \U$29163 ( \29416 , \29415 , \28804 );
nor \U$29164 ( \29417 , \29414 , \29416 );
not \U$29165 ( \29418 , \29417 );
or \U$29166 ( \29419 , \29407 , \29418 );
or \U$29167 ( \29420 , \29406 , \29417 );
not \U$29168 ( \29421 , \28846 );
not \U$29169 ( \29422 , \28868 );
or \U$29170 ( \29423 , \29421 , \29422 );
nand \U$29171 ( \29424 , \28867 , \28845 );
nand \U$29172 ( \29425 , \29423 , \29424 );
and \U$29173 ( \29426 , \29425 , \28855 );
not \U$29174 ( \29427 , \29425 );
and \U$29175 ( \29428 , \29427 , \28854 );
nor \U$29176 ( \29429 , \29426 , \29428 );
not \U$29177 ( \29430 , \29429 );
nand \U$29178 ( \29431 , \29420 , \29430 );
nand \U$29179 ( \29432 , \29419 , \29431 );
xor \U$29180 ( \29433 , \29404 , \29432 );
xor \U$29181 ( \29434 , \28654 , \28643 );
xnor \U$29182 ( \29435 , \29434 , \28634 );
not \U$29183 ( \29436 , \28588 );
not \U$29184 ( \29437 , \29436 );
not \U$29185 ( \29438 , \28568 );
or \U$29186 ( \29439 , \29437 , \29438 );
nand \U$29187 ( \29440 , \28567 , \28588 );
nand \U$29188 ( \29441 , \29439 , \29440 );
xor \U$29189 ( \29442 , \29441 , \28578 );
or \U$29190 ( \29443 , \29435 , \29442 );
xor \U$29191 ( \29444 , \28620 , \28600 );
xor \U$29192 ( \29445 , \29444 , \28609 );
not \U$29193 ( \29446 , \29445 );
nand \U$29194 ( \29447 , \29443 , \29446 );
nand \U$29195 ( \29448 , \29435 , \29442 );
nand \U$29196 ( \29449 , \29447 , \29448 );
xor \U$29197 ( \29450 , \29433 , \29449 );
nand \U$29198 ( \29451 , \29346 , \29450 );
not \U$29199 ( \29452 , \29344 );
nand \U$29200 ( \29453 , \29452 , \29014 );
nand \U$29201 ( \29454 , \29451 , \29453 );
not \U$29202 ( \29455 , RIbe2b090_115);
not \U$29203 ( \29456 , \1111 );
or \U$29204 ( \29457 , \29455 , \29456 );
nand \U$29205 ( \29458 , \20849 , RIbe2a280_85);
nand \U$29206 ( \29459 , \29457 , \29458 );
and \U$29207 ( \29460 , \29459 , \1131 );
not \U$29208 ( \29461 , \29459 );
and \U$29209 ( \29462 , \29461 , \6831 );
nor \U$29210 ( \29463 , \29460 , \29462 );
not \U$29211 ( \29464 , \29463 );
not \U$29212 ( \29465 , RIbe2b270_119);
not \U$29213 ( \29466 , \1631 );
or \U$29214 ( \29467 , \29465 , \29466 );
nand \U$29215 ( \29468 , \1098 , RIbe2b108_116);
nand \U$29216 ( \29469 , \29467 , \29468 );
and \U$29217 ( \29470 , \29469 , \1458 );
not \U$29218 ( \29471 , \29469 );
and \U$29219 ( \29472 , \29471 , \1309 );
nor \U$29220 ( \29473 , \29470 , \29472 );
nand \U$29221 ( \29474 , \29464 , \29473 );
not \U$29222 ( \29475 , RIbe2a208_84);
not \U$29223 ( \29476 , \20674 );
or \U$29224 ( \29477 , \29475 , \29476 );
nand \U$29225 ( \29478 , \2384 , RIbe2a190_83);
nand \U$29226 ( \29479 , \29477 , \29478 );
xor \U$29227 ( \29480 , \29479 , \1076 );
not \U$29228 ( \29481 , \29480 );
and \U$29229 ( \29482 , \29474 , \29481 );
nor \U$29230 ( \29483 , \29464 , \29473 );
nor \U$29231 ( \29484 , \29482 , \29483 );
not \U$29232 ( \29485 , \29484 );
not \U$29233 ( \29486 , \29485 );
not \U$29234 ( \29487 , RIbe2a988_100);
not \U$29235 ( \29488 , \21478 );
or \U$29236 ( \29489 , \29487 , \29488 );
nand \U$29237 ( \29490 , RIbe2a910_99, \6800 );
nand \U$29238 ( \29491 , \29489 , \29490 );
and \U$29239 ( \29492 , \29491 , \2887 );
not \U$29240 ( \29493 , \29491 );
and \U$29241 ( \29494 , \29493 , \3290 );
nor \U$29242 ( \29495 , \29492 , \29494 );
not \U$29243 ( \29496 , RIbe2a5c8_92);
not \U$29244 ( \29497 , \2566 );
and \U$29245 ( \29498 , \29497 , \2568 );
not \U$29246 ( \29499 , \29498 );
or \U$29247 ( \29500 , \29496 , \29499 );
nand \U$29248 ( \29501 , \2901 , RIbe2a550_91);
nand \U$29249 ( \29502 , \29500 , \29501 );
not \U$29250 ( \29503 , \29502 );
not \U$29251 ( \29504 , \2379 );
and \U$29252 ( \29505 , \29503 , \29504 );
and \U$29253 ( \29506 , \29502 , \2576 );
nor \U$29254 ( \29507 , \29505 , \29506 );
nand \U$29255 ( \29508 , \29495 , \29507 );
not \U$29256 ( \29509 , RIbe2b5b8_126);
not \U$29257 ( \29510 , \20625 );
or \U$29258 ( \29511 , \29509 , \29510 );
nand \U$29259 ( \29512 , \7438 , RIbe2a3e8_88);
nand \U$29260 ( \29513 , \29511 , \29512 );
not \U$29261 ( \29514 , \29513 );
not \U$29262 ( \29515 , \3448 );
and \U$29263 ( \29516 , \29514 , \29515 );
and \U$29264 ( \29517 , \29513 , \3698 );
nor \U$29265 ( \29518 , \29516 , \29517 );
not \U$29266 ( \29519 , \29518 );
and \U$29267 ( \29520 , \29508 , \29519 );
nor \U$29268 ( \29521 , \29507 , \29495 );
nor \U$29269 ( \29522 , \29520 , \29521 );
not \U$29270 ( \29523 , \29522 );
not \U$29271 ( \29524 , \29523 );
or \U$29272 ( \29525 , \29486 , \29524 );
nand \U$29273 ( \29526 , \29522 , \29484 );
not \U$29274 ( \29527 , RIbe2afa0_113);
not \U$29275 ( \29528 , \2424 );
or \U$29276 ( \29529 , \29527 , \29528 );
nand \U$29277 ( \29530 , \7905 , RIbe2af28_112);
nand \U$29278 ( \29531 , \29529 , \29530 );
and \U$29279 ( \29532 , \29531 , \1813 );
not \U$29280 ( \29533 , \29531 );
and \U$29281 ( \29534 , \29533 , \1010 );
nor \U$29282 ( \29535 , \29532 , \29534 );
not \U$29283 ( \29536 , \29535 );
not \U$29284 ( \29537 , \29536 );
not \U$29285 ( \29538 , RIbe2b1f8_118);
not \U$29286 ( \29539 , \21344 );
or \U$29287 ( \29540 , \29538 , \29539 );
nand \U$29288 ( \29541 , \1146 , RIbe2b180_117);
nand \U$29289 ( \29542 , \29540 , \29541 );
and \U$29290 ( \29543 , \29542 , \7899 );
not \U$29291 ( \29544 , \29542 );
and \U$29292 ( \29545 , \29544 , \4742 );
nor \U$29293 ( \29546 , \29543 , \29545 );
not \U$29294 ( \29547 , \29546 );
or \U$29295 ( \29548 , \29537 , \29547 );
not \U$29296 ( \29549 , \29546 );
not \U$29297 ( \29550 , \29549 );
not \U$29298 ( \29551 , \29535 );
or \U$29299 ( \29552 , \29550 , \29551 );
not \U$29300 ( \29553 , RIbe2b630_127);
not \U$29301 ( \29554 , \29388 );
or \U$29302 ( \29555 , \29553 , \29554 );
nand \U$29303 ( \29556 , RIbe2b018_114, \740 );
nand \U$29304 ( \29557 , \29555 , \29556 );
not \U$29305 ( \29558 , \29557 );
not \U$29306 ( \29559 , \564 );
and \U$29307 ( \29560 , \29558 , \29559 );
and \U$29308 ( \29561 , \29557 , \564 );
nor \U$29309 ( \29562 , \29560 , \29561 );
not \U$29310 ( \29563 , \29562 );
nand \U$29311 ( \29564 , \29552 , \29563 );
nand \U$29312 ( \29565 , \29548 , \29564 );
nand \U$29313 ( \29566 , \29526 , \29565 );
nand \U$29314 ( \29567 , \29525 , \29566 );
not \U$29315 ( \29568 , RIbe29650_59);
not \U$29316 ( \29569 , \13518 );
or \U$29317 ( \29570 , \29568 , \29569 );
nand \U$29318 ( \29571 , \12890 , RIbe29038_46);
nand \U$29319 ( \29572 , \29570 , \29571 );
and \U$29320 ( \29573 , \29572 , \12801 );
not \U$29321 ( \29574 , \29572 );
and \U$29322 ( \29575 , \29574 , \14103 );
nor \U$29323 ( \29576 , \29573 , \29575 );
not \U$29324 ( \29577 , RIbe28fc0_45);
not \U$29325 ( \29578 , \12811 );
or \U$29326 ( \29579 , \29577 , \29578 );
nand \U$29327 ( \29580 , RIbe290b0_47, RIbe2ae38_110);
nand \U$29328 ( \29581 , \29579 , \29580 );
xnor \U$29329 ( \29582 , \29581 , RIbe2aeb0_111);
nand \U$29330 ( \29583 , \29576 , \29582 );
not \U$29331 ( \29584 , \15263 );
not \U$29332 ( \29585 , RIbe29830_63);
not \U$29333 ( \29586 , \12831 );
or \U$29334 ( \29587 , \29585 , \29586 );
nand \U$29335 ( \29588 , \12835 , RIbe296c8_60);
nand \U$29336 ( \29589 , \29587 , \29588 );
not \U$29337 ( \29590 , \29589 );
or \U$29338 ( \29591 , \29584 , \29590 );
or \U$29339 ( \29592 , \29589 , \12823 );
nand \U$29340 ( \29593 , \29591 , \29592 );
and \U$29341 ( \29594 , \29583 , \29593 );
nor \U$29342 ( \29595 , \29576 , \29582 );
nor \U$29343 ( \29596 , \29594 , \29595 );
not \U$29344 ( \29597 , \29596 );
not \U$29345 ( \29598 , RIbe28b10_35);
not \U$29346 ( \29599 , \20530 );
or \U$29347 ( \29600 , \29598 , \29599 );
nand \U$29348 ( \29601 , \12212 , RIbe28b88_36);
nand \U$29349 ( \29602 , \29600 , \29601 );
xor \U$29350 ( \29603 , \29602 , \10943 );
and \U$29351 ( \29604 , \10915 , RIbe28408_20);
and \U$29352 ( \29605 , \13038 , RIbe28390_19);
nor \U$29353 ( \29606 , \29604 , \29605 );
and \U$29354 ( \29607 , \29606 , \10926 );
not \U$29355 ( \29608 , \29606 );
and \U$29356 ( \29609 , \29608 , \10912 );
nor \U$29357 ( \29610 , \29607 , \29609 );
nand \U$29358 ( \29611 , \29603 , \29610 );
not \U$29359 ( \29612 , \12195 );
not \U$29360 ( \29613 , \15627 );
not \U$29361 ( \29614 , \5177 );
and \U$29362 ( \29615 , \29613 , \29614 );
and \U$29363 ( \29616 , \12942 , RIbe29290_51);
nor \U$29364 ( \29617 , \29615 , \29616 );
not \U$29365 ( \29618 , \29617 );
or \U$29366 ( \29619 , \29612 , \29618 );
or \U$29367 ( \29620 , \12195 , \29617 );
nand \U$29368 ( \29621 , \29619 , \29620 );
and \U$29369 ( \29622 , \29611 , \29621 );
nor \U$29370 ( \29623 , \29610 , \29603 );
nor \U$29371 ( \29624 , \29622 , \29623 );
not \U$29372 ( \29625 , \29624 );
or \U$29373 ( \29626 , \29597 , \29625 );
not \U$29374 ( \29627 , RIbe29560_57);
not \U$29375 ( \29628 , \12871 );
or \U$29376 ( \29629 , \29627 , \29628 );
nand \U$29377 ( \29630 , \12710 , RIbe28228_16);
nand \U$29378 ( \29631 , \29629 , \29630 );
not \U$29379 ( \29632 , \29631 );
not \U$29380 ( \29633 , \13583 );
and \U$29381 ( \29634 , \29632 , \29633 );
and \U$29382 ( \29635 , \29631 , \12723 );
nor \U$29383 ( \29636 , \29634 , \29635 );
not \U$29384 ( \29637 , \29636 );
not \U$29385 ( \29638 , \29637 );
not \U$29386 ( \29639 , RIbe281b0_15);
not \U$29387 ( \29640 , \14071 );
or \U$29388 ( \29641 , \29639 , \29640 );
nand \U$29389 ( \29642 , \12735 , RIbe280c0_13);
nand \U$29390 ( \29643 , \29641 , \29642 );
and \U$29391 ( \29644 , \29643 , \12852 );
not \U$29392 ( \29645 , \29643 );
and \U$29393 ( \29646 , \29645 , \12746 );
nor \U$29394 ( \29647 , \29644 , \29646 );
not \U$29395 ( \29648 , \29647 );
or \U$29396 ( \29649 , \29638 , \29648 );
or \U$29397 ( \29650 , \29647 , \29637 );
not \U$29398 ( \29651 , \12753 );
not \U$29399 ( \29652 , \9078 );
and \U$29400 ( \29653 , \29651 , \29652 );
and \U$29401 ( \29654 , \12921 , RIbe289a8_32);
nor \U$29402 ( \29655 , \29653 , \29654 );
and \U$29403 ( \29656 , \29655 , \12770 );
not \U$29404 ( \29657 , \29655 );
and \U$29405 ( \29658 , \29657 , \12927 );
nor \U$29406 ( \29659 , \29656 , \29658 );
nand \U$29407 ( \29660 , \29650 , \29659 );
nand \U$29408 ( \29661 , \29649 , \29660 );
nand \U$29409 ( \29662 , \29626 , \29661 );
or \U$29410 ( \29663 , \29596 , \29624 );
nand \U$29411 ( \29664 , \29662 , \29663 );
xor \U$29412 ( \29665 , \29567 , \29664 );
not \U$29413 ( \29666 , \6546 );
not \U$29414 ( \29667 , \6541 );
not \U$29415 ( \29668 , \7775 );
and \U$29416 ( \29669 , \29667 , \29668 );
and \U$29417 ( \29670 , \6535 , RIbe29bf0_71);
nor \U$29418 ( \29671 , \29669 , \29670 );
not \U$29419 ( \29672 , \29671 );
or \U$29420 ( \29673 , \29666 , \29672 );
or \U$29421 ( \29674 , \29671 , \15730 );
nand \U$29422 ( \29675 , \29673 , \29674 );
not \U$29423 ( \29676 , RIbe29dd0_75);
not \U$29424 ( \29677 , \6138 );
or \U$29425 ( \29678 , \29676 , \29677 );
nand \U$29426 ( \29679 , \6859 , RIbe29c68_72);
nand \U$29427 ( \29680 , \29678 , \29679 );
and \U$29428 ( \29681 , \29680 , \10969 );
not \U$29429 ( \29682 , \29680 );
and \U$29430 ( \29683 , \29682 , \6141 );
nor \U$29431 ( \29684 , \29681 , \29683 );
xor \U$29432 ( \29685 , \29675 , \29684 );
not \U$29433 ( \29686 , RIbe28ed0_43);
not \U$29434 ( \29687 , \7941 );
or \U$29435 ( \29688 , \29686 , \29687 );
nand \U$29436 ( \29689 , \13436 , RIbe27fd0_11);
nand \U$29437 ( \29690 , \29688 , \29689 );
and \U$29438 ( \29691 , \29690 , \6601 );
not \U$29439 ( \29692 , \29690 );
and \U$29440 ( \29693 , \29692 , \29121 );
nor \U$29441 ( \29694 , \29691 , \29693 );
and \U$29442 ( \29695 , \29685 , \29694 );
and \U$29443 ( \29696 , \29675 , \29684 );
or \U$29444 ( \29697 , \29695 , \29696 );
not \U$29445 ( \29698 , RIbe29fb0_79);
not \U$29446 ( \29699 , \20796 );
or \U$29447 ( \29700 , \29698 , \29699 );
nand \U$29448 ( \29701 , \8246 , RIbe29e48_76);
nand \U$29449 ( \29702 , \29700 , \29701 );
and \U$29450 ( \29703 , \29702 , \5754 );
not \U$29451 ( \29704 , \29702 );
and \U$29452 ( \29705 , \29704 , \5045 );
nor \U$29453 ( \29706 , \29703 , \29705 );
not \U$29454 ( \29707 , RIbe2a370_87);
not \U$29455 ( \29708 , \5058 );
or \U$29456 ( \29709 , \29707 , \29708 );
nand \U$29457 ( \29710 , RIbe2a2f8_86, \7858 );
nand \U$29458 ( \29711 , \29709 , \29710 );
and \U$29459 ( \29712 , \29711 , \7865 );
not \U$29460 ( \29713 , \29711 );
and \U$29461 ( \29714 , \29713 , \4603 );
nor \U$29462 ( \29715 , \29712 , \29714 );
nand \U$29463 ( \29716 , \29706 , \29715 );
not \U$29464 ( \29717 , \20465 );
not \U$29465 ( \29718 , RIbe2acd0_107);
not \U$29466 ( \29719 , \20809 );
or \U$29467 ( \29720 , \29718 , \29719 );
not \U$29468 ( \29721 , \14374 );
nand \U$29469 ( \29722 , \29721 , \5730 );
nand \U$29470 ( \29723 , \29720 , \29722 );
not \U$29471 ( \29724 , \29723 );
or \U$29472 ( \29725 , \29717 , \29724 );
or \U$29473 ( \29726 , \29723 , \20465 );
nand \U$29474 ( \29727 , \29725 , \29726 );
and \U$29475 ( \29728 , \29716 , \29727 );
nor \U$29476 ( \29729 , \29706 , \29715 );
nor \U$29477 ( \29730 , \29728 , \29729 );
not \U$29478 ( \29731 , \29730 );
nor \U$29479 ( \29732 , \29697 , \29731 );
not \U$29480 ( \29733 , RIbe287c8_28);
not \U$29481 ( \29734 , \14633 );
or \U$29482 ( \29735 , \29733 , \29734 );
nand \U$29483 ( \29736 , \10952 , RIbe28480_21);
nand \U$29484 ( \29737 , \29735 , \29736 );
and \U$29485 ( \29738 , \29737 , \6949 );
not \U$29486 ( \29739 , \29737 );
and \U$29487 ( \29740 , \29739 , \6950 );
nor \U$29488 ( \29741 , \29738 , \29740 );
not \U$29489 ( \29742 , \29741 );
not \U$29490 ( \29743 , RIbe27f58_10);
not \U$29491 ( \29744 , \6560 );
or \U$29492 ( \29745 , \29743 , \29744 );
nand \U$29493 ( \29746 , \6963 , RIbe27e68_8);
nand \U$29494 ( \29747 , \29745 , \29746 );
xor \U$29495 ( \29748 , \29747 , \6569 );
not \U$29496 ( \29749 , \29748 );
or \U$29497 ( \29750 , \29742 , \29749 );
and \U$29498 ( \29751 , \7298 , RIbe28660_25);
not \U$29499 ( \29752 , RIbe285e8_24);
nor \U$29500 ( \29753 , \29752 , \6984 );
nor \U$29501 ( \29754 , \29751 , \29753 );
and \U$29502 ( \29755 , \29754 , \8004 );
not \U$29503 ( \29756 , \29754 );
not \U$29504 ( \29757 , \8004 );
and \U$29505 ( \29758 , \29756 , \29757 );
nor \U$29506 ( \29759 , \29755 , \29758 );
nand \U$29507 ( \29760 , \29750 , \29759 );
not \U$29508 ( \29761 , \29741 );
not \U$29509 ( \29762 , \29748 );
nand \U$29510 ( \29763 , \29761 , \29762 );
nand \U$29511 ( \29764 , \29760 , \29763 );
not \U$29512 ( \29765 , \29764 );
or \U$29513 ( \29766 , \29732 , \29765 );
nand \U$29514 ( \29767 , \29697 , \29731 );
nand \U$29515 ( \29768 , \29766 , \29767 );
and \U$29516 ( \29769 , \29665 , \29768 );
and \U$29517 ( \29770 , \29567 , \29664 );
or \U$29518 ( \29771 , \29769 , \29770 );
not \U$29519 ( \29772 , \29159 );
not \U$29520 ( \29773 , \29178 );
or \U$29521 ( \29774 , \29772 , \29773 );
or \U$29522 ( \29775 , \29178 , \29159 );
nand \U$29523 ( \29776 , \29774 , \29775 );
xor \U$29524 ( \29777 , \29776 , \29168 );
not \U$29525 ( \29778 , \29289 );
not \U$29526 ( \29779 , \29279 );
or \U$29527 ( \29780 , \29778 , \29779 );
or \U$29528 ( \29781 , \29289 , \29279 );
nand \U$29529 ( \29782 , \29780 , \29781 );
and \U$29530 ( \29783 , \29782 , \29269 );
not \U$29531 ( \29784 , \29782 );
not \U$29532 ( \29785 , \29269 );
and \U$29533 ( \29786 , \29784 , \29785 );
nor \U$29534 ( \29787 , \29783 , \29786 );
nand \U$29535 ( \29788 , \29777 , \29787 );
not \U$29536 ( \29789 , \29135 );
and \U$29537 ( \29790 , \29125 , \29789 );
not \U$29538 ( \29791 , \29125 );
and \U$29539 ( \29792 , \29791 , \29135 );
or \U$29540 ( \29793 , \29790 , \29792 );
not \U$29541 ( \29794 , \29146 );
and \U$29542 ( \29795 , \29793 , \29794 );
not \U$29543 ( \29796 , \29793 );
and \U$29544 ( \29797 , \29796 , \29146 );
nor \U$29545 ( \29798 , \29795 , \29797 );
not \U$29546 ( \29799 , \29798 );
and \U$29547 ( \29800 , \29788 , \29799 );
nor \U$29548 ( \29801 , \29777 , \29787 );
nor \U$29549 ( \29802 , \29800 , \29801 );
not \U$29550 ( \29803 , \29802 );
xor \U$29551 ( \29804 , \29055 , \29066 );
buf \U$29552 ( \29805 , \29048 );
xor \U$29553 ( \29806 , \29804 , \29805 );
not \U$29554 ( \29807 , \29806 );
not \U$29555 ( \29808 , \29191 );
not \U$29556 ( \29809 , \29214 );
or \U$29557 ( \29810 , \29808 , \29809 );
nand \U$29558 ( \29811 , \29201 , \29190 );
nand \U$29559 ( \29812 , \29810 , \29811 );
not \U$29560 ( \29813 , \29211 );
and \U$29561 ( \29814 , \29812 , \29813 );
not \U$29562 ( \29815 , \29812 );
and \U$29563 ( \29816 , \29815 , \29211 );
nor \U$29564 ( \29817 , \29814 , \29816 );
not \U$29565 ( \29818 , \29817 );
or \U$29566 ( \29819 , \29807 , \29818 );
xor \U$29567 ( \29820 , \29080 , \29094 );
xnor \U$29568 ( \29821 , \29820 , \29107 );
nand \U$29569 ( \29822 , \29819 , \29821 );
not \U$29570 ( \29823 , \29806 );
not \U$29571 ( \29824 , \29817 );
nand \U$29572 ( \29825 , \29823 , \29824 );
nand \U$29573 ( \29826 , \29822 , \29825 );
not \U$29574 ( \29827 , \29826 );
not \U$29575 ( \29828 , \29827 );
or \U$29576 ( \29829 , \29803 , \29828 );
not \U$29577 ( \29830 , \29396 );
not \U$29578 ( \29831 , \29378 );
or \U$29579 ( \29832 , \29830 , \29831 );
or \U$29580 ( \29833 , \29378 , \29396 );
nand \U$29581 ( \29834 , \29832 , \29833 );
not \U$29582 ( \29835 , \29383 );
and \U$29583 ( \29836 , \29834 , \29835 );
not \U$29584 ( \29837 , \29834 );
and \U$29585 ( \29838 , \29837 , \29383 );
nor \U$29586 ( \29839 , \29836 , \29838 );
not \U$29587 ( \29840 , \29331 );
not \U$29588 ( \29841 , \29304 );
or \U$29589 ( \29842 , \29840 , \29841 );
or \U$29590 ( \29843 , \29331 , \29304 );
nand \U$29591 ( \29844 , \29842 , \29843 );
and \U$29592 ( \29845 , \29844 , \29315 );
not \U$29593 ( \29846 , \29844 );
and \U$29594 ( \29847 , \29846 , \29314 );
nor \U$29595 ( \29848 , \29845 , \29847 );
xor \U$29596 ( \29849 , \29839 , \29848 );
xor \U$29597 ( \29850 , \29256 , \29236 );
xor \U$29598 ( \29851 , \29850 , \29245 );
and \U$29599 ( \29852 , \29849 , \29851 );
and \U$29600 ( \29853 , \29839 , \29848 );
or \U$29601 ( \29854 , \29852 , \29853 );
nand \U$29602 ( \29855 , \29829 , \29854 );
not \U$29603 ( \29856 , \29827 );
not \U$29604 ( \29857 , \29802 );
nand \U$29605 ( \29858 , \29856 , \29857 );
nand \U$29606 ( \29859 , \29855 , \29858 );
xor \U$29607 ( \29860 , \29771 , \29859 );
xor \U$29608 ( \29861 , \29442 , \29445 );
xor \U$29609 ( \29862 , \29861 , \29435 );
not \U$29610 ( \29863 , \29862 );
not \U$29611 ( \29864 , \28994 );
not \U$29612 ( \29865 , \29001 );
or \U$29613 ( \29866 , \29864 , \29865 );
or \U$29614 ( \29867 , \29001 , \28994 );
nand \U$29615 ( \29868 , \29866 , \29867 );
and \U$29616 ( \29869 , \29868 , \28997 );
not \U$29617 ( \29870 , \29868 );
and \U$29618 ( \29871 , \29870 , \29004 );
nor \U$29619 ( \29872 , \29869 , \29871 );
not \U$29620 ( \29873 , \29872 );
or \U$29621 ( \29874 , \29863 , \29873 );
not \U$29622 ( \29875 , \29406 );
not \U$29623 ( \29876 , \29875 );
not \U$29624 ( \29877 , \29430 );
or \U$29625 ( \29878 , \29876 , \29877 );
nand \U$29626 ( \29879 , \29429 , \29406 );
nand \U$29627 ( \29880 , \29878 , \29879 );
and \U$29628 ( \29881 , \29880 , \29417 );
not \U$29629 ( \29882 , \29880 );
not \U$29630 ( \29883 , \29417 );
and \U$29631 ( \29884 , \29882 , \29883 );
nor \U$29632 ( \29885 , \29881 , \29884 );
nand \U$29633 ( \29886 , \29874 , \29885 );
not \U$29634 ( \29887 , \29862 );
not \U$29635 ( \29888 , \29872 );
nand \U$29636 ( \29889 , \29887 , \29888 );
nand \U$29637 ( \29890 , \29886 , \29889 );
and \U$29638 ( \29891 , \29860 , \29890 );
and \U$29639 ( \29892 , \29771 , \29859 );
or \U$29640 ( \29893 , \29891 , \29892 );
xor \U$29641 ( \29894 , \29454 , \29893 );
not \U$29642 ( \29895 , \29366 );
not \U$29643 ( \29896 , \29401 );
or \U$29644 ( \29897 , \29895 , \29896 );
nand \U$29645 ( \29898 , \29365 , \29355 );
nand \U$29646 ( \29899 , \29897 , \29898 );
nor \U$29647 ( \29900 , \29398 , \29399 );
xor \U$29648 ( \29901 , \29899 , \29900 );
not \U$29649 ( \29902 , \29901 );
not \U$29650 ( \29903 , \29334 );
not \U$29651 ( \29904 , \29903 );
not \U$29652 ( \29905 , \29337 );
or \U$29653 ( \29906 , \29904 , \29905 );
nand \U$29654 ( \29907 , \29293 , \29334 );
nand \U$29655 ( \29908 , \29906 , \29907 );
xor \U$29656 ( \29909 , \29908 , \29259 );
not \U$29657 ( \29910 , \29909 );
or \U$29658 ( \29911 , \29902 , \29910 );
xor \U$29659 ( \29912 , \29181 , \29219 );
xnor \U$29660 ( \29913 , \29912 , \29216 );
nand \U$29661 ( \29914 , \29911 , \29913 );
or \U$29662 ( \29915 , \29909 , \29901 );
nand \U$29663 ( \29916 , \29914 , \29915 );
xor \U$29664 ( \29917 , \28591 , \28623 );
xor \U$29665 ( \29918 , \29917 , \28658 );
not \U$29666 ( \29919 , \29918 );
and \U$29667 ( \29920 , \28692 , \28753 );
not \U$29668 ( \29921 , \28692 );
and \U$29669 ( \29922 , \29921 , \28754 );
nor \U$29670 ( \29923 , \29920 , \29922 );
not \U$29671 ( \29924 , \29923 );
not \U$29672 ( \29925 , \28723 );
and \U$29673 ( \29926 , \29924 , \29925 );
and \U$29674 ( \29927 , \29923 , \28723 );
nor \U$29675 ( \29928 , \29926 , \29927 );
not \U$29676 ( \29929 , \29928 );
or \U$29677 ( \29930 , \29919 , \29929 );
or \U$29678 ( \29931 , \29928 , \29918 );
nand \U$29679 ( \29932 , \29930 , \29931 );
not \U$29680 ( \29933 , \28833 );
not \U$29681 ( \29934 , \28830 );
or \U$29682 ( \29935 , \29933 , \29934 );
nand \U$29683 ( \29936 , \28794 , \28829 );
nand \U$29684 ( \29937 , \29935 , \29936 );
not \U$29685 ( \29938 , \28871 );
and \U$29686 ( \29939 , \29937 , \29938 );
not \U$29687 ( \29940 , \29937 );
and \U$29688 ( \29941 , \29940 , \28871 );
nor \U$29689 ( \29942 , \29939 , \29941 );
not \U$29690 ( \29943 , \29942 );
and \U$29691 ( \29944 , \29932 , \29943 );
not \U$29692 ( \29945 , \29932 );
and \U$29693 ( \29946 , \29945 , \29942 );
nor \U$29694 ( \29947 , \29944 , \29946 );
xor \U$29695 ( \29948 , \29916 , \29947 );
xor \U$29696 ( \29949 , \28900 , \28902 );
xor \U$29697 ( \29950 , \29949 , \28915 );
not \U$29698 ( \29951 , \28926 );
not \U$29699 ( \29952 , \28940 );
or \U$29700 ( \29953 , \29951 , \29952 );
or \U$29701 ( \29954 , \28926 , \28940 );
nand \U$29702 ( \29955 , \29953 , \29954 );
and \U$29703 ( \29956 , \29955 , \28943 );
not \U$29704 ( \29957 , \29955 );
and \U$29705 ( \29958 , \29957 , \28929 );
nor \U$29706 ( \29959 , \29956 , \29958 );
xor \U$29707 ( \29960 , \29950 , \29959 );
xor \U$29708 ( \29961 , \28953 , \28955 );
xor \U$29709 ( \29962 , \29961 , \28958 );
xor \U$29710 ( \29963 , \29960 , \29962 );
and \U$29711 ( \29964 , \29948 , \29963 );
and \U$29712 ( \29965 , \29916 , \29947 );
or \U$29713 ( \29966 , \29964 , \29965 );
and \U$29714 ( \29967 , \29894 , \29966 );
and \U$29715 ( \29968 , \29454 , \29893 );
or \U$29716 ( \29969 , \29967 , \29968 );
not \U$29717 ( \29970 , \29969 );
xor \U$29718 ( \29971 , \28873 , \28661 );
xor \U$29719 ( \29972 , \29971 , \28757 );
not \U$29720 ( \29973 , \28961 );
not \U$29721 ( \29974 , \29973 );
xor \U$29722 ( \29975 , \28945 , \28918 );
not \U$29723 ( \29976 , \29975 );
or \U$29724 ( \29977 , \29974 , \29976 );
or \U$29725 ( \29978 , \29975 , \29973 );
nand \U$29726 ( \29979 , \29977 , \29978 );
xor \U$29727 ( \29980 , \29972 , \29979 );
not \U$29728 ( \29981 , \27773 );
not \U$29729 ( \29982 , \27666 );
or \U$29730 ( \29983 , \29981 , \29982 );
or \U$29731 ( \29984 , \27773 , \27666 );
nand \U$29732 ( \29985 , \29983 , \29984 );
not \U$29733 ( \29986 , \27878 );
and \U$29734 ( \29987 , \29985 , \29986 );
not \U$29735 ( \29988 , \29985 );
and \U$29736 ( \29989 , \29988 , \27878 );
nor \U$29737 ( \29990 , \29987 , \29989 );
not \U$29738 ( \29991 , \29990 );
xnor \U$29739 ( \29992 , \28229 , \28165 );
xnor \U$29740 ( \29993 , \29992 , \28196 );
not \U$29741 ( \29994 , \28883 );
not \U$29742 ( \29995 , \28880 );
or \U$29743 ( \29996 , \29994 , \29995 );
or \U$29744 ( \29997 , \28880 , \28883 );
nand \U$29745 ( \29998 , \29996 , \29997 );
xnor \U$29746 ( \29999 , \28877 , \29998 );
xor \U$29747 ( \30000 , \29993 , \29999 );
not \U$29748 ( \30001 , \30000 );
or \U$29749 ( \30002 , \29991 , \30001 );
or \U$29750 ( \30003 , \30000 , \29990 );
nand \U$29751 ( \30004 , \30002 , \30003 );
and \U$29752 ( \30005 , \29980 , \30004 );
and \U$29753 ( \30006 , \29972 , \29979 );
or \U$29754 ( \30007 , \30005 , \30006 );
not \U$29755 ( \30008 , \30007 );
nand \U$29756 ( \30009 , \29970 , \30008 );
not \U$29757 ( \30010 , \30009 );
xor \U$29758 ( \30011 , \28875 , \28889 );
xor \U$29759 ( \30012 , \30011 , \28963 );
xor \U$29760 ( \30013 , \27558 , \27880 );
xor \U$29761 ( \30014 , \30013 , \28030 );
xor \U$29762 ( \30015 , \30012 , \30014 );
xor \U$29763 ( \30016 , \28241 , \28266 );
xor \U$29764 ( \30017 , \30016 , \28555 );
xor \U$29765 ( \30018 , \30015 , \30017 );
not \U$29766 ( \30019 , \30018 );
or \U$29767 ( \30020 , \30010 , \30019 );
nand \U$29768 ( \30021 , \29969 , \30007 );
nand \U$29769 ( \30022 , \30020 , \30021 );
xor \U$29770 ( \30023 , \28975 , \30022 );
not \U$29771 ( \30024 , \29222 );
not \U$29772 ( \30025 , \29340 );
or \U$29773 ( \30026 , \30024 , \30025 );
nand \U$29774 ( \30027 , \30026 , \29114 );
nand \U$29775 ( \30028 , \29339 , \29221 );
nand \U$29776 ( \30029 , \30027 , \30028 );
not \U$29777 ( \30030 , \30029 );
xor \U$29778 ( \30031 , \29404 , \29432 );
and \U$29779 ( \30032 , \30031 , \29449 );
and \U$29780 ( \30033 , \29404 , \29432 );
or \U$29781 ( \30034 , \30032 , \30033 );
not \U$29782 ( \30035 , \30034 );
or \U$29783 ( \30036 , \30030 , \30035 );
or \U$29784 ( \30037 , \30034 , \30029 );
not \U$29785 ( \30038 , \28980 );
not \U$29786 ( \30039 , \30038 );
not \U$29787 ( \30040 , \28987 );
or \U$29788 ( \30041 , \30039 , \30040 );
not \U$29789 ( \30042 , \29006 );
or \U$29790 ( \30043 , \28987 , \30038 );
nand \U$29791 ( \30044 , \30042 , \30043 );
nand \U$29792 ( \30045 , \30041 , \30044 );
nand \U$29793 ( \30046 , \30037 , \30045 );
nand \U$29794 ( \30047 , \30036 , \30046 );
xnor \U$29795 ( \30048 , \28076 , \28109 );
xor \U$29796 ( \30049 , \30048 , \28141 );
not \U$29797 ( \30050 , \29928 );
not \U$29798 ( \30051 , \29942 );
or \U$29799 ( \30052 , \30050 , \30051 );
nand \U$29800 ( \30053 , \30052 , \29918 );
not \U$29801 ( \30054 , \29928 );
nand \U$29802 ( \30055 , \30054 , \29943 );
nand \U$29803 ( \30056 , \30053 , \30055 );
xor \U$29804 ( \30057 , \30049 , \30056 );
xor \U$29805 ( \30058 , \29950 , \29959 );
and \U$29806 ( \30059 , \30058 , \29962 );
and \U$29807 ( \30060 , \29950 , \29959 );
or \U$29808 ( \30061 , \30059 , \30060 );
and \U$29809 ( \30062 , \30057 , \30061 );
and \U$29810 ( \30063 , \30049 , \30056 );
or \U$29811 ( \30064 , \30062 , \30063 );
xor \U$29812 ( \30065 , \30047 , \30064 );
and \U$29813 ( \30066 , \29993 , \29999 );
or \U$29814 ( \30067 , \29990 , \30066 );
or \U$29815 ( \30068 , \29999 , \29993 );
nand \U$29816 ( \30069 , \30067 , \30068 );
and \U$29817 ( \30070 , \30065 , \30069 );
and \U$29818 ( \30071 , \30047 , \30064 );
or \U$29819 ( \30072 , \30070 , \30071 );
xor \U$29820 ( \30073 , \30012 , \30014 );
and \U$29821 ( \30074 , \30073 , \30017 );
and \U$29822 ( \30075 , \30012 , \30014 );
or \U$29823 ( \30076 , \30074 , \30075 );
xor \U$29824 ( \30077 , \30072 , \30076 );
not \U$29825 ( \30078 , \28232 );
not \U$29826 ( \30079 , \28144 );
or \U$29827 ( \30080 , \30078 , \30079 );
nand \U$29828 ( \30081 , \30080 , \28042 );
nand \U$29829 ( \30082 , \28145 , \28233 );
nand \U$29830 ( \30083 , \30081 , \30082 );
not \U$29831 ( \30084 , \28245 );
not \U$29832 ( \30085 , \28260 );
or \U$29833 ( \30086 , \30084 , \30085 );
nand \U$29834 ( \30087 , \30086 , \28255 );
not \U$29835 ( \30088 , \28245 );
nand \U$29836 ( \30089 , \30088 , \28261 );
nand \U$29837 ( \30090 , \30087 , \30089 );
xor \U$29838 ( \30091 , \30083 , \30090 );
or \U$29839 ( \30092 , \28550 , \28448 );
nand \U$29840 ( \30093 , \30092 , \28360 );
nand \U$29841 ( \30094 , \28448 , \28550 );
nand \U$29842 ( \30095 , \30093 , \30094 );
xnor \U$29843 ( \30096 , \30091 , \30095 );
not \U$29844 ( \30097 , \27896 );
not \U$29845 ( \30098 , \27968 );
or \U$29846 ( \30099 , \30097 , \30098 );
or \U$29847 ( \30100 , \27896 , \27968 );
nand \U$29848 ( \30101 , \30100 , \28025 );
nand \U$29849 ( \30102 , \30099 , \30101 );
nand \U$29850 ( \30103 , \28274 , \1362 );
not \U$29851 ( \30104 , \30103 );
not \U$29852 ( \30105 , \28289 );
or \U$29853 ( \30106 , \30104 , \30105 );
nand \U$29854 ( \30107 , \28275 , \1663 );
nand \U$29855 ( \30108 , \30106 , \30107 );
or \U$29856 ( \30109 , \28358 , \28338 );
nand \U$29857 ( \30110 , \30109 , \28347 );
nand \U$29858 ( \30111 , \28358 , \28338 );
nand \U$29859 ( \30112 , \30110 , \30111 );
xor \U$29860 ( \30113 , \30108 , \30112 );
or \U$29861 ( \30114 , \28312 , \28303 );
nand \U$29862 ( \30115 , \30114 , \28324 );
nand \U$29863 ( \30116 , \28312 , \28303 );
nand \U$29864 ( \30117 , \30115 , \30116 );
xor \U$29865 ( \30118 , \30113 , \30117 );
not \U$29866 ( \30119 , \30118 );
not \U$29867 ( \30120 , \28456 );
not \U$29868 ( \30121 , \28465 );
or \U$29869 ( \30122 , \30120 , \30121 );
or \U$29870 ( \30123 , \28465 , \28456 );
nand \U$29871 ( \30124 , \30123 , \28475 );
nand \U$29872 ( \30125 , \30122 , \30124 );
not \U$29873 ( \30126 , \30125 );
not \U$29874 ( \30127 , \30126 );
and \U$29875 ( \30128 , \28495 , \28486 );
nor \U$29876 ( \30129 , \30128 , \28506 );
nor \U$29877 ( \30130 , \28495 , \28486 );
nor \U$29878 ( \30131 , \30129 , \30130 );
not \U$29879 ( \30132 , \30131 );
not \U$29880 ( \30133 , \30132 );
or \U$29881 ( \30134 , \30127 , \30133 );
nand \U$29882 ( \30135 , \30125 , \30131 );
nand \U$29883 ( \30136 , \30134 , \30135 );
not \U$29884 ( \30137 , \30136 );
and \U$29885 ( \30138 , \28533 , \28544 );
nor \U$29886 ( \30139 , \30138 , \28524 );
nor \U$29887 ( \30140 , \28544 , \28533 );
nor \U$29888 ( \30141 , \30139 , \30140 );
not \U$29889 ( \30142 , \30141 );
and \U$29890 ( \30143 , \30137 , \30142 );
and \U$29891 ( \30144 , \30136 , \30141 );
nor \U$29892 ( \30145 , \30143 , \30144 );
not \U$29893 ( \30146 , \30145 );
or \U$29894 ( \30147 , \30119 , \30146 );
or \U$29895 ( \30148 , \30118 , \30145 );
nand \U$29896 ( \30149 , \30147 , \30148 );
xor \U$29897 ( \30150 , \28369 , \28378 );
and \U$29898 ( \30151 , \30150 , \28388 );
and \U$29899 ( \30152 , \28369 , \28378 );
or \U$29900 ( \30153 , \30151 , \30152 );
not \U$29901 ( \30154 , \30153 );
not \U$29902 ( \30155 , \30154 );
or \U$29903 ( \30156 , \28415 , \28399 );
not \U$29904 ( \30157 , \28405 );
nand \U$29905 ( \30158 , \30156 , \30157 );
nand \U$29906 ( \30159 , \28415 , \28399 );
nand \U$29907 ( \30160 , \30158 , \30159 );
not \U$29908 ( \30161 , \30160 );
or \U$29909 ( \30162 , \30155 , \30161 );
nand \U$29910 ( \30163 , \30153 , \30158 , \30159 );
nand \U$29911 ( \30164 , \30162 , \30163 );
and \U$29912 ( \30165 , \28437 , \28446 );
nor \U$29913 ( \30166 , \30165 , \28425 );
nor \U$29914 ( \30167 , \28437 , \28446 );
nor \U$29915 ( \30168 , \30166 , \30167 );
and \U$29916 ( \30169 , \30164 , \30168 );
not \U$29917 ( \30170 , \30164 );
not \U$29918 ( \30171 , \30168 );
and \U$29919 ( \30172 , \30170 , \30171 );
nor \U$29920 ( \30173 , \30169 , \30172 );
not \U$29921 ( \30174 , \30173 );
and \U$29922 ( \30175 , \30149 , \30174 );
not \U$29923 ( \30176 , \30149 );
and \U$29924 ( \30177 , \30176 , \30173 );
nor \U$29925 ( \30178 , \30175 , \30177 );
xor \U$29926 ( \30179 , \30102 , \30178 );
and \U$29927 ( \30180 , \1357 , RIbe2ab68_104);
and \U$29928 ( \30181 , \1831 , RIbe2aaf0_103);
nor \U$29929 ( \30182 , \30180 , \30181 );
and \U$29930 ( \30183 , \30182 , \269 );
not \U$29931 ( \30184 , \30182 );
and \U$29932 ( \30185 , \30184 , \6058 );
nor \U$29933 ( \30186 , \30183 , \30185 );
not \U$29934 ( \30187 , \27974 );
nand \U$29935 ( \30188 , \30187 , \27982 );
xor \U$29936 ( \30189 , \30186 , \30188 );
and \U$29937 ( \30190 , \28023 , \28013 );
not \U$29938 ( \30191 , \28003 );
nor \U$29939 ( \30192 , \30190 , \30191 );
nor \U$29940 ( \30193 , \28023 , \28013 );
nor \U$29941 ( \30194 , \30192 , \30193 );
xnor \U$29942 ( \30195 , \30189 , \30194 );
not \U$29943 ( \30196 , RIbe2b1f8_118);
not \U$29944 ( \30197 , \546 );
or \U$29945 ( \30198 , \30196 , \30197 );
nand \U$29946 ( \30199 , \552 , RIbe2b180_117);
nand \U$29947 ( \30200 , \30198 , \30199 );
not \U$29948 ( \30201 , \30200 );
not \U$29949 ( \30202 , \424 );
and \U$29950 ( \30203 , \30201 , \30202 );
and \U$29951 ( \30204 , \30200 , \7124 );
nor \U$29952 ( \30205 , \30203 , \30204 );
not \U$29953 ( \30206 , RIbe2afa0_113);
not \U$29954 ( \30207 , \1773 );
or \U$29955 ( \30208 , \30206 , \30207 );
nand \U$29956 ( \30209 , \429 , RIbe2af28_112);
nand \U$29957 ( \30210 , \30208 , \30209 );
and \U$29958 ( \30211 , \30210 , \306 );
not \U$29959 ( \30212 , \30210 );
and \U$29960 ( \30213 , \30212 , \1547 );
nor \U$29961 ( \30214 , \30211 , \30213 );
xor \U$29962 ( \30215 , \30205 , \30214 );
and \U$29963 ( \30216 , \6311 , RIbe2b630_127);
and \U$29964 ( \30217 , \9816 , RIbe2b018_114);
nor \U$29965 ( \30218 , \30216 , \30217 );
and \U$29966 ( \30219 , \30218 , \293 );
not \U$29967 ( \30220 , \30218 );
and \U$29968 ( \30221 , \30220 , \300 );
nor \U$29969 ( \30222 , \30219 , \30221 );
xor \U$29970 ( \30223 , \30215 , \30222 );
and \U$29971 ( \30224 , \10759 , RIbe2a988_100);
and \U$29972 ( \30225 , \1117 , RIbe2a910_99);
nor \U$29973 ( \30226 , \30224 , \30225 );
and \U$29974 ( \30227 , \30226 , \1131 );
not \U$29975 ( \30228 , \30226 );
and \U$29976 ( \30229 , \30228 , \1125 );
nor \U$29977 ( \30230 , \30227 , \30229 );
not \U$29978 ( \30231 , \4064 );
not \U$29979 ( \30232 , \13089 );
and \U$29980 ( \30233 , \30231 , \30232 );
and \U$29981 ( \30234 , \27613 , RIbe2b5b8_126);
nor \U$29982 ( \30235 , \30233 , \30234 );
and \U$29983 ( \30236 , \30235 , \1277 );
not \U$29984 ( \30237 , \30235 );
and \U$29985 ( \30238 , \30237 , \1076 );
nor \U$29986 ( \30239 , \30236 , \30238 );
xor \U$29987 ( \30240 , \30230 , \30239 );
not \U$29988 ( \30241 , RIbe2a5c8_92);
not \U$29989 ( \30242 , \1632 );
or \U$29990 ( \30243 , \30241 , \30242 );
nand \U$29991 ( \30244 , \1454 , RIbe2a550_91);
nand \U$29992 ( \30245 , \30243 , \30244 );
not \U$29993 ( \30246 , \30245 );
not \U$29994 ( \30247 , \2418 );
and \U$29995 ( \30248 , \30246 , \30247 );
and \U$29996 ( \30249 , \30245 , \1458 );
nor \U$29997 ( \30250 , \30248 , \30249 );
xnor \U$29998 ( \30251 , \30240 , \30250 );
xor \U$29999 ( \30252 , \30223 , \30251 );
not \U$30000 ( \30253 , RIbe2b270_119);
not \U$30001 ( \30254 , \6350 );
or \U$30002 ( \30255 , \30253 , \30254 );
nand \U$30003 ( \30256 , \1179 , RIbe2b108_116);
nand \U$30004 ( \30257 , \30255 , \30256 );
not \U$30005 ( \30258 , \30257 );
not \U$30006 ( \30259 , \564 );
and \U$30007 ( \30260 , \30258 , \30259 );
and \U$30008 ( \30261 , \30257 , \1618 );
nor \U$30009 ( \30262 , \30260 , \30261 );
not \U$30010 ( \30263 , RIbe2a208_84);
not \U$30011 ( \30264 , \1143 );
or \U$30012 ( \30265 , \30263 , \30264 );
nand \U$30013 ( \30266 , \1147 , RIbe2a190_83);
nand \U$30014 ( \30267 , \30265 , \30266 );
and \U$30015 ( \30268 , \30267 , \3993 );
not \U$30016 ( \30269 , \30267 );
and \U$30017 ( \30270 , \30269 , \1157 );
nor \U$30018 ( \30271 , \30268 , \30270 );
xor \U$30019 ( \30272 , \30262 , \30271 );
not \U$30020 ( \30273 , \752 );
not \U$30021 ( \30274 , RIbe2b090_115);
not \U$30022 ( \30275 , \6747 );
or \U$30023 ( \30276 , \30274 , \30275 );
nand \U$30024 ( \30277 , \1203 , RIbe2a280_85);
nand \U$30025 ( \30278 , \30276 , \30277 );
not \U$30026 ( \30279 , \30278 );
or \U$30027 ( \30280 , \30273 , \30279 );
or \U$30028 ( \30281 , \752 , \30278 );
nand \U$30029 ( \30282 , \30280 , \30281 );
xnor \U$30030 ( \30283 , \30272 , \30282 );
xor \U$30031 ( \30284 , \30252 , \30283 );
xor \U$30032 ( \30285 , \30195 , \30284 );
not \U$30033 ( \30286 , RIbe2acd0_107);
not \U$30034 ( \30287 , \3451 );
or \U$30035 ( \30288 , \30286 , \30287 );
nand \U$30036 ( \30289 , \3457 , RIbe2a028_80);
nand \U$30037 ( \30290 , \30288 , \30289 );
and \U$30038 ( \30291 , \30290 , \3461 );
not \U$30039 ( \30292 , \30290 );
and \U$30040 ( \30293 , \30292 , \4346 );
nor \U$30041 ( \30294 , \30291 , \30293 );
not \U$30042 ( \30295 , \30294 );
not \U$30043 ( \30296 , RIbe29fb0_79);
not \U$30044 ( \30297 , \20764 );
or \U$30045 ( \30298 , \30296 , \30297 );
nand \U$30046 ( \30299 , \8368 , RIbe29e48_76);
nand \U$30047 ( \30300 , \30298 , \30299 );
and \U$30048 ( \30301 , \30300 , \3471 );
not \U$30049 ( \30302 , \30300 );
and \U$30050 ( \30303 , \30302 , \4821 );
nor \U$30051 ( \30304 , \30301 , \30303 );
not \U$30052 ( \30305 , \30304 );
or \U$30053 ( \30306 , \30295 , \30305 );
or \U$30054 ( \30307 , \30294 , \30304 );
nand \U$30055 ( \30308 , \30306 , \30307 );
not \U$30056 ( \30309 , RIbe2a370_87);
not \U$30057 ( \30310 , \8342 );
or \U$30058 ( \30311 , \30309 , \30310 );
nand \U$30059 ( \30312 , \3267 , RIbe2a2f8_86);
nand \U$30060 ( \30313 , \30311 , \30312 );
and \U$30061 ( \30314 , \30313 , \4059 );
not \U$30062 ( \30315 , \30313 );
and \U$30063 ( \30316 , \30315 , \7457 );
nor \U$30064 ( \30317 , \30314 , \30316 );
and \U$30065 ( \30318 , \30308 , \30317 );
not \U$30066 ( \30319 , \30308 );
not \U$30067 ( \30320 , \30317 );
and \U$30068 ( \30321 , \30319 , \30320 );
nor \U$30069 ( \30322 , \30318 , \30321 );
not \U$30070 ( \30323 , RIbe29bf0_71);
not \U$30071 ( \30324 , \21097 );
or \U$30072 ( \30325 , \30323 , \30324 );
nand \U$30073 ( \30326 , \22378 , RIbe28f48_44);
nand \U$30074 ( \30327 , \30325 , \30326 );
xor \U$30075 ( \30328 , \30327 , \4592 );
not \U$30076 ( \30329 , \30328 );
not \U$30077 ( \30330 , RIbe28ed0_43);
not \U$30078 ( \30331 , \5455 );
or \U$30079 ( \30332 , \30330 , \30331 );
nand \U$30080 ( \30333 , \6634 , RIbe27fd0_11);
nand \U$30081 ( \30334 , \30332 , \30333 );
not \U$30082 ( \30335 , \10984 );
and \U$30083 ( \30336 , \30334 , \30335 );
not \U$30084 ( \30337 , \30334 );
and \U$30085 ( \30338 , \30337 , \5754 );
nor \U$30086 ( \30339 , \30336 , \30338 );
not \U$30087 ( \30340 , \30339 );
or \U$30088 ( \30341 , \30329 , \30340 );
or \U$30089 ( \30342 , \30339 , \30328 );
nand \U$30090 ( \30343 , \30341 , \30342 );
not \U$30091 ( \30344 , RIbe29dd0_75);
not \U$30092 ( \30345 , \5058 );
or \U$30093 ( \30346 , \30344 , \30345 );
nand \U$30094 ( \30347 , \6418 , RIbe29c68_72);
nand \U$30095 ( \30348 , \30346 , \30347 );
not \U$30096 ( \30349 , \30348 );
not \U$30097 ( \30350 , \4323 );
and \U$30098 ( \30351 , \30349 , \30350 );
and \U$30099 ( \30352 , \30348 , \7865 );
nor \U$30100 ( \30353 , \30351 , \30352 );
and \U$30101 ( \30354 , \30343 , \30353 );
not \U$30102 ( \30355 , \30343 );
not \U$30103 ( \30356 , \30353 );
and \U$30104 ( \30357 , \30355 , \30356 );
nor \U$30105 ( \30358 , \30354 , \30357 );
xor \U$30106 ( \30359 , \30322 , \30358 );
not \U$30107 ( \30360 , RIbe28660_25);
not \U$30108 ( \30361 , \6536 );
or \U$30109 ( \30362 , \30360 , \30361 );
nand \U$30110 ( \30363 , \10348 , RIbe285e8_24);
nand \U$30111 ( \30364 , \30362 , \30363 );
not \U$30112 ( \30365 , \30364 );
not \U$30113 ( \30366 , \6891 );
and \U$30114 ( \30367 , \30365 , \30366 );
and \U$30115 ( \30368 , \30364 , \6548 );
nor \U$30116 ( \30369 , \30367 , \30368 );
not \U$30117 ( \30370 , \30369 );
not \U$30118 ( \30371 , RIbe287c8_28);
not \U$30119 ( \30372 , \6868 );
or \U$30120 ( \30373 , \30371 , \30372 );
nand \U$30121 ( \30374 , \13436 , RIbe28480_21);
nand \U$30122 ( \30375 , \30373 , \30374 );
and \U$30123 ( \30376 , \30375 , \6601 );
not \U$30124 ( \30377 , \30375 );
and \U$30125 ( \30378 , \30377 , \7949 );
nor \U$30126 ( \30379 , \30376 , \30378 );
not \U$30127 ( \30380 , \30379 );
or \U$30128 ( \30381 , \30370 , \30380 );
or \U$30129 ( \30382 , \30379 , \30369 );
nand \U$30130 ( \30383 , \30381 , \30382 );
not \U$30131 ( \30384 , RIbe27f58_10);
not \U$30132 ( \30385 , \8231 );
or \U$30133 ( \30386 , \30384 , \30385 );
nand \U$30134 ( \30387 , \9939 , RIbe27e68_8);
nand \U$30135 ( \30388 , \30386 , \30387 );
and \U$30136 ( \30389 , \30388 , \6144 );
not \U$30137 ( \30390 , \30388 );
and \U$30138 ( \30391 , \30390 , \10972 );
nor \U$30139 ( \30392 , \30389 , \30391 );
xor \U$30140 ( \30393 , \30383 , \30392 );
xor \U$30141 ( \30394 , \30359 , \30393 );
xor \U$30142 ( \30395 , \30285 , \30394 );
xor \U$30143 ( \30396 , \30179 , \30395 );
xor \U$30144 ( \30397 , \30096 , \30396 );
or \U$30145 ( \30398 , \27521 , \27557 );
nand \U$30146 ( \30399 , \30398 , \27492 );
nand \U$30147 ( \30400 , \27521 , \27557 );
nand \U$30148 ( \30401 , \30399 , \30400 );
xor \U$30149 ( \30402 , \27886 , \27890 );
and \U$30150 ( \30403 , \30402 , \27895 );
and \U$30151 ( \30404 , \27886 , \27890 );
or \U$30152 ( \30405 , \30403 , \30404 );
xor \U$30153 ( \30406 , \30401 , \30405 );
xor \U$30154 ( \30407 , \27929 , \27935 );
and \U$30155 ( \30408 , \30407 , \27967 );
and \U$30156 ( \30409 , \27929 , \27935 );
or \U$30157 ( \30410 , \30408 , \30409 );
xor \U$30158 ( \30411 , \30406 , \30410 );
not \U$30159 ( \30412 , RIbe29a88_68);
not \U$30160 ( \30413 , \13010 );
or \U$30161 ( \30414 , \30412 , \30413 );
nand \U$30162 ( \30415 , \12835 , RIbe27d78_6);
nand \U$30163 ( \30416 , \30414 , \30415 );
xnor \U$30164 ( \30417 , \12823 , \30416 );
not \U$30165 ( \30418 , \30417 );
not \U$30166 ( \30419 , RIbe27d00_5);
not \U$30167 ( \30420 , \12787 );
or \U$30168 ( \30421 , \30419 , \30420 );
nand \U$30169 ( \30422 , \12890 , RIbe27c10_3);
nand \U$30170 ( \30423 , \30421 , \30422 );
and \U$30171 ( \30424 , \30423 , \14103 );
not \U$30172 ( \30425 , \30423 );
and \U$30173 ( \30426 , \30425 , \12893 );
nor \U$30174 ( \30427 , \30424 , \30426 );
nand \U$30175 ( \30428 , \13004 , RIbe28e58_42);
nand \U$30176 ( \30429 , RIbe28de0_41, RIbe2ae38_110);
and \U$30177 ( \30430 , \30428 , \30429 );
xor \U$30178 ( \30431 , \30430 , RIbe2aeb0_111);
xor \U$30179 ( \30432 , \30427 , \30431 );
not \U$30180 ( \30433 , \30432 );
or \U$30181 ( \30434 , \30418 , \30433 );
or \U$30182 ( \30435 , \30432 , \30417 );
nand \U$30183 ( \30436 , \30434 , \30435 );
xor \U$30184 ( \30437 , \28294 , \28327 );
and \U$30185 ( \30438 , \30437 , \28359 );
and \U$30186 ( \30439 , \28294 , \28327 );
or \U$30187 ( \30440 , \30438 , \30439 );
xor \U$30188 ( \30441 , \30436 , \30440 );
not \U$30189 ( \30442 , RIbe28b10_35);
not \U$30190 ( \30443 , \7298 );
or \U$30191 ( \30444 , \30442 , \30443 );
nand \U$30192 ( \30445 , \10898 , RIbe28b88_36);
nand \U$30193 ( \30446 , \30444 , \30445 );
xor \U$30194 ( \30447 , \30446 , \6992 );
not \U$30195 ( \30448 , \30447 );
not \U$30196 ( \30449 , \30448 );
not \U$30197 ( \30450 , RIbe29290_51);
not \U$30198 ( \30451 , \7975 );
or \U$30199 ( \30452 , \30450 , \30451 );
nand \U$30200 ( \30453 , \10952 , RIbe28a20_33);
nand \U$30201 ( \30454 , \30452 , \30453 );
and \U$30202 ( \30455 , \30454 , \7985 );
not \U$30203 ( \30456 , \30454 );
and \U$30204 ( \30457 , \30456 , \6949 );
nor \U$30205 ( \30458 , \30455 , \30457 );
not \U$30206 ( \30459 , \30458 );
not \U$30207 ( \30460 , \30459 );
or \U$30208 ( \30461 , \30449 , \30460 );
nand \U$30209 ( \30462 , \30458 , \30447 );
nand \U$30210 ( \30463 , \30461 , \30462 );
not \U$30211 ( \30464 , RIbe28408_20);
not \U$30212 ( \30465 , \6958 );
or \U$30213 ( \30466 , \30464 , \30465 );
nand \U$30214 ( \30467 , \6963 , RIbe28390_19);
nand \U$30215 ( \30468 , \30466 , \30467 );
and \U$30216 ( \30469 , \30468 , \6569 );
not \U$30217 ( \30470 , \30468 );
and \U$30218 ( \30471 , \30470 , \7293 );
nor \U$30219 ( \30472 , \30469 , \30471 );
and \U$30220 ( \30473 , \30463 , \30472 );
not \U$30221 ( \30474 , \30463 );
not \U$30222 ( \30475 , \30472 );
and \U$30223 ( \30476 , \30474 , \30475 );
nor \U$30224 ( \30477 , \30473 , \30476 );
and \U$30225 ( \30478 , \16431 , RIbe289a8_32);
and \U$30226 ( \30479 , \13038 , RIbe28930_31);
nor \U$30227 ( \30480 , \30478 , \30479 );
and \U$30228 ( \30481 , \30480 , \16437 );
not \U$30229 ( \30482 , \30480 );
and \U$30230 ( \30483 , \30482 , \12202 );
nor \U$30231 ( \30484 , \30481 , \30483 );
not \U$30232 ( \30485 , RIbe29560_57);
not \U$30233 ( \30486 , \13024 );
or \U$30234 ( \30487 , \30485 , \30486 );
nand \U$30235 ( \30488 , \12971 , RIbe28228_16);
nand \U$30236 ( \30489 , \30487 , \30488 );
not \U$30237 ( \30490 , \30489 );
not \U$30238 ( \30491 , \10943 );
and \U$30239 ( \30492 , \30490 , \30491 );
and \U$30240 ( \30493 , \30489 , \13030 );
nor \U$30241 ( \30494 , \30492 , \30493 );
xor \U$30242 ( \30495 , \30484 , \30494 );
not \U$30243 ( \30496 , RIbe281b0_15);
not \U$30244 ( \30497 , \13049 );
or \U$30245 ( \30498 , \30496 , \30497 );
nand \U$30246 ( \30499 , \15628 , RIbe280c0_13);
nand \U$30247 ( \30500 , \30498 , \30499 );
not \U$30248 ( \30501 , \30500 );
not \U$30249 ( \30502 , \17005 );
and \U$30250 ( \30503 , \30501 , \30502 );
and \U$30251 ( \30504 , \30500 , \12960 );
nor \U$30252 ( \30505 , \30503 , \30504 );
xor \U$30253 ( \30506 , \30495 , \30505 );
xor \U$30254 ( \30507 , \30477 , \30506 );
not \U$30255 ( \30508 , RIbe29650_59);
not \U$30256 ( \30509 , \15573 );
or \U$30257 ( \30510 , \30508 , \30509 );
nand \U$30258 ( \30511 , \12710 , RIbe29038_46);
nand \U$30259 ( \30512 , \30510 , \30511 );
not \U$30260 ( \30513 , \30512 );
not \U$30261 ( \30514 , \12723 );
and \U$30262 ( \30515 , \30513 , \30514 );
and \U$30263 ( \30516 , \30512 , \12723 );
nor \U$30264 ( \30517 , \30515 , \30516 );
not \U$30265 ( \30518 , \30517 );
not \U$30266 ( \30519 , RIbe28fc0_45);
not \U$30267 ( \30520 , \15161 );
or \U$30268 ( \30521 , \30519 , \30520 );
nand \U$30269 ( \30522 , \12735 , RIbe290b0_47);
nand \U$30270 ( \30523 , \30521 , \30522 );
and \U$30271 ( \30524 , \30523 , \12743 );
not \U$30272 ( \30525 , \30523 );
and \U$30273 ( \30526 , \30525 , \12746 );
nor \U$30274 ( \30527 , \30524 , \30526 );
not \U$30275 ( \30528 , \30527 );
or \U$30276 ( \30529 , \30518 , \30528 );
or \U$30277 ( \30530 , \30517 , \30527 );
nand \U$30278 ( \30531 , \30529 , \30530 );
not \U$30279 ( \30532 , \12752 );
not \U$30280 ( \30533 , RIbe296c8_60);
not \U$30281 ( \30534 , \30533 );
and \U$30282 ( \30535 , \30532 , \30534 );
and \U$30283 ( \30536 , \15615 , RIbe29830_63);
nor \U$30284 ( \30537 , \30535 , \30536 );
and \U$30285 ( \30538 , \30537 , \12774 );
not \U$30286 ( \30539 , \30537 );
and \U$30287 ( \30540 , \30539 , \12769 );
nor \U$30288 ( \30541 , \30538 , \30540 );
and \U$30289 ( \30542 , \30531 , \30541 );
not \U$30290 ( \30543 , \30531 );
not \U$30291 ( \30544 , \30541 );
and \U$30292 ( \30545 , \30543 , \30544 );
nor \U$30293 ( \30546 , \30542 , \30545 );
not \U$30294 ( \30547 , \30546 );
and \U$30295 ( \30548 , \30507 , \30547 );
not \U$30296 ( \30549 , \30507 );
and \U$30297 ( \30550 , \30549 , \30546 );
nor \U$30298 ( \30551 , \30548 , \30550 );
xor \U$30299 ( \30552 , \30441 , \30551 );
xor \U$30300 ( \30553 , \30411 , \30552 );
xor \U$30301 ( \30554 , \27986 , \27993 );
and \U$30302 ( \30555 , \30554 , \28024 );
and \U$30303 ( \30556 , \27986 , \27993 );
or \U$30304 ( \30557 , \30555 , \30556 );
nand \U$30305 ( \30558 , \28545 , \28476 );
and \U$30306 ( \30559 , \30558 , \28511 );
nor \U$30307 ( \30560 , \28476 , \28545 );
nor \U$30308 ( \30561 , \30559 , \30560 );
xor \U$30309 ( \30562 , \30557 , \30561 );
xor \U$30310 ( \30563 , \28389 , \28416 );
and \U$30311 ( \30564 , \30563 , \28447 );
and \U$30312 ( \30565 , \28389 , \28416 );
or \U$30313 ( \30566 , \30564 , \30565 );
xnor \U$30314 ( \30567 , \30562 , \30566 );
xor \U$30315 ( \30568 , \30553 , \30567 );
xnor \U$30316 ( \30569 , \30397 , \30568 );
xor \U$30317 ( \30570 , \30077 , \30569 );
and \U$30318 ( \30571 , \30023 , \30570 );
and \U$30319 ( \30572 , \28975 , \30022 );
or \U$30320 ( \30573 , \30571 , \30572 );
not \U$30321 ( \30574 , \30573 );
not \U$30322 ( \30575 , \30568 );
nand \U$30323 ( \30576 , \30575 , \30096 );
and \U$30324 ( \30577 , \30576 , \30396 );
nor \U$30325 ( \30578 , \30575 , \30096 );
nor \U$30326 ( \30579 , \30577 , \30578 );
not \U$30327 ( \30580 , \30579 );
buf \U$30328 ( \30581 , \30145 );
nand \U$30329 ( \30582 , \30173 , \30581 );
and \U$30330 ( \30583 , \30582 , \30118 );
nor \U$30331 ( \30584 , \30581 , \30173 );
nor \U$30332 ( \30585 , \30583 , \30584 );
not \U$30333 ( \30586 , \30328 );
not \U$30334 ( \30587 , \30586 );
not \U$30335 ( \30588 , \30356 );
or \U$30336 ( \30589 , \30587 , \30588 );
not \U$30337 ( \30590 , \30328 );
not \U$30338 ( \30591 , \30353 );
or \U$30339 ( \30592 , \30590 , \30591 );
nand \U$30340 ( \30593 , \30592 , \30339 );
nand \U$30341 ( \30594 , \30589 , \30593 );
not \U$30342 ( \30595 , \30475 );
not \U$30343 ( \30596 , \30458 );
or \U$30344 ( \30597 , \30595 , \30596 );
not \U$30345 ( \30598 , \30459 );
not \U$30346 ( \30599 , \30472 );
or \U$30347 ( \30600 , \30598 , \30599 );
nand \U$30348 ( \30601 , \30600 , \30448 );
nand \U$30349 ( \30602 , \30597 , \30601 );
xor \U$30350 ( \30603 , \30594 , \30602 );
or \U$30351 ( \30604 , \30379 , \30392 );
not \U$30352 ( \30605 , \30369 );
nand \U$30353 ( \30606 , \30604 , \30605 );
nand \U$30354 ( \30607 , \30379 , \30392 );
nand \U$30355 ( \30608 , \30606 , \30607 );
xnor \U$30356 ( \30609 , \30603 , \30608 );
xor \U$30357 ( \30610 , \30585 , \30609 );
xor \U$30358 ( \30611 , \30195 , \30284 );
and \U$30359 ( \30612 , \30611 , \30394 );
and \U$30360 ( \30613 , \30195 , \30284 );
or \U$30361 ( \30614 , \30612 , \30613 );
xor \U$30362 ( \30615 , \30610 , \30614 );
not \U$30363 ( \30616 , \28969 );
not \U$30364 ( \30617 , \28034 );
or \U$30365 ( \30618 , \30616 , \30617 );
nand \U$30366 ( \30619 , \30618 , \28558 );
nand \U$30367 ( \30620 , \28033 , \28966 );
nand \U$30368 ( \30621 , \30619 , \30620 );
xor \U$30369 ( \30622 , \30615 , \30621 );
not \U$30370 ( \30623 , \30622 );
or \U$30371 ( \30624 , \30580 , \30623 );
or \U$30372 ( \30625 , \30579 , \30622 );
nand \U$30373 ( \30626 , \30624 , \30625 );
xor \U$30374 ( \30627 , \30072 , \30076 );
and \U$30375 ( \30628 , \30627 , \30569 );
and \U$30376 ( \30629 , \30072 , \30076 );
or \U$30377 ( \30630 , \30628 , \30629 );
xor \U$30378 ( \30631 , \30626 , \30630 );
not \U$30379 ( \30632 , \30557 );
not \U$30380 ( \30633 , \30632 );
not \U$30381 ( \30634 , \30561 );
or \U$30382 ( \30635 , \30633 , \30634 );
nand \U$30383 ( \30636 , \30635 , \30566 );
not \U$30384 ( \30637 , \30561 );
nand \U$30385 ( \30638 , \30637 , \30557 );
and \U$30386 ( \30639 , \30636 , \30638 );
not \U$30387 ( \30640 , \30639 );
xor \U$30388 ( \30641 , \30401 , \30405 );
and \U$30389 ( \30642 , \30641 , \30410 );
and \U$30390 ( \30643 , \30401 , \30405 );
or \U$30391 ( \30644 , \30642 , \30643 );
not \U$30392 ( \30645 , \30644 );
and \U$30393 ( \30646 , \30640 , \30645 );
and \U$30394 ( \30647 , \30639 , \30644 );
nor \U$30395 ( \30648 , \30646 , \30647 );
not \U$30396 ( \30649 , \30648 );
xor \U$30397 ( \30650 , \30436 , \30440 );
and \U$30398 ( \30651 , \30650 , \30551 );
and \U$30399 ( \30652 , \30436 , \30440 );
or \U$30400 ( \30653 , \30651 , \30652 );
not \U$30401 ( \30654 , \30653 );
and \U$30402 ( \30655 , \30649 , \30654 );
and \U$30403 ( \30656 , \30648 , \30653 );
nor \U$30404 ( \30657 , \30655 , \30656 );
not \U$30405 ( \30658 , \30427 );
nand \U$30406 ( \30659 , \30658 , \30431 );
and \U$30407 ( \30660 , \30659 , \30417 );
nor \U$30408 ( \30661 , \30658 , \30431 );
nor \U$30409 ( \30662 , \30660 , \30661 );
not \U$30410 ( \30663 , \30662 );
xor \U$30411 ( \30664 , \30484 , \30494 );
and \U$30412 ( \30665 , \30664 , \30505 );
and \U$30413 ( \30666 , \30484 , \30494 );
or \U$30414 ( \30667 , \30665 , \30666 );
not \U$30415 ( \30668 , \30667 );
not \U$30416 ( \30669 , \30517 );
or \U$30417 ( \30670 , \30669 , \30527 );
nand \U$30418 ( \30671 , \30670 , \30544 );
nand \U$30419 ( \30672 , \30669 , \30527 );
nand \U$30420 ( \30673 , \30671 , \30672 );
not \U$30421 ( \30674 , \30673 );
or \U$30422 ( \30675 , \30668 , \30674 );
or \U$30423 ( \30676 , \30673 , \30667 );
nand \U$30424 ( \30677 , \30675 , \30676 );
not \U$30425 ( \30678 , \30677 );
or \U$30426 ( \30679 , \30663 , \30678 );
or \U$30427 ( \30680 , \30677 , \30662 );
nand \U$30428 ( \30681 , \30679 , \30680 );
buf \U$30429 ( \30682 , \30205 );
nand \U$30430 ( \30683 , \30682 , \30222 );
and \U$30431 ( \30684 , \30683 , \30214 );
nor \U$30432 ( \30685 , \30682 , \30222 );
nor \U$30433 ( \30686 , \30684 , \30685 );
not \U$30434 ( \30687 , RIbe2b108_116);
not \U$30435 ( \30688 , \29388 );
or \U$30436 ( \30689 , \30687 , \30688 );
nand \U$30437 ( \30690 , \1179 , RIbe2b090_115);
nand \U$30438 ( \30691 , \30689 , \30690 );
not \U$30439 ( \30692 , \30691 );
not \U$30440 ( \30693 , \564 );
and \U$30441 ( \30694 , \30692 , \30693 );
and \U$30442 ( \30695 , \1618 , \30691 );
nor \U$30443 ( \30696 , \30694 , \30695 );
not \U$30444 ( \30697 , \30696 );
and \U$30445 ( \30698 , \546 , RIbe2b180_117);
and \U$30446 ( \30699 , \552 , RIbe2b270_119);
nor \U$30447 ( \30700 , \30698 , \30699 );
and \U$30448 ( \30701 , \30700 , \424 );
not \U$30449 ( \30702 , \30700 );
and \U$30450 ( \30703 , \30702 , \7123 );
nor \U$30451 ( \30704 , \30701 , \30703 );
not \U$30452 ( \30705 , \30704 );
or \U$30453 ( \30706 , \30697 , \30705 );
or \U$30454 ( \30707 , \30704 , \30696 );
nand \U$30455 ( \30708 , \30706 , \30707 );
not \U$30456 ( \30709 , RIbe2af28_112);
not \U$30457 ( \30710 , \1337 );
or \U$30458 ( \30711 , \30709 , \30710 );
nand \U$30459 ( \30712 , \429 , RIbe2b1f8_118);
nand \U$30460 ( \30713 , \30711 , \30712 );
and \U$30461 ( \30714 , \30713 , \306 );
not \U$30462 ( \30715 , \30713 );
and \U$30463 ( \30716 , \30715 , \313 );
nor \U$30464 ( \30717 , \30714 , \30716 );
and \U$30465 ( \30718 , \30708 , \30717 );
not \U$30466 ( \30719 , \30708 );
not \U$30467 ( \30720 , \30717 );
and \U$30468 ( \30721 , \30719 , \30720 );
nor \U$30469 ( \30722 , \30718 , \30721 );
xor \U$30470 ( \30723 , \30686 , \30722 );
not \U$30471 ( \30724 , RIbe2aaf0_103);
nor \U$30472 ( \30725 , \258 , \257 );
not \U$30473 ( \30726 , \30725 );
or \U$30474 ( \30727 , \30724 , \30726 );
nand \U$30475 ( \30728 , \263 , RIbe2b630_127);
nand \U$30476 ( \30729 , \30727 , \30728 );
not \U$30477 ( \30730 , \30729 );
not \U$30478 ( \30731 , \1362 );
and \U$30479 ( \30732 , \30730 , \30731 );
and \U$30480 ( \30733 , \6058 , \30729 );
nor \U$30481 ( \30734 , \30732 , \30733 );
not \U$30482 ( \30735 , RIbe2b018_114);
not \U$30483 ( \30736 , \1252 );
or \U$30484 ( \30737 , \30735 , \30736 );
nand \U$30485 ( \30738 , \9816 , RIbe2afa0_113);
nand \U$30486 ( \30739 , \30737 , \30738 );
and \U$30487 ( \30740 , \30739 , \293 );
not \U$30488 ( \30741 , \30739 );
and \U$30489 ( \30742 , \30741 , \300 );
nor \U$30490 ( \30743 , \30740 , \30742 );
xnor \U$30491 ( \30744 , \30734 , \30743 );
nand \U$30492 ( \30745 , \330 , RIbe2ab68_104);
and \U$30493 ( \30746 , \30745 , \1374 );
not \U$30494 ( \30747 , \30745 );
and \U$30495 ( \30748 , \30747 , \338 );
or \U$30496 ( \30749 , \30746 , \30748 );
xor \U$30497 ( \30750 , \30744 , \30749 );
xnor \U$30498 ( \30751 , \30723 , \30750 );
not \U$30499 ( \30752 , \30751 );
not \U$30500 ( \30753 , \30752 );
nand \U$30501 ( \30754 , \30317 , \30294 );
and \U$30502 ( \30755 , \30754 , \30304 );
nor \U$30503 ( \30756 , \30317 , \30294 );
nor \U$30504 ( \30757 , \30755 , \30756 );
and \U$30505 ( \30758 , \30230 , \30250 );
nor \U$30506 ( \30759 , \30758 , \30239 );
nor \U$30507 ( \30760 , \30230 , \30250 );
nor \U$30508 ( \30761 , \30759 , \30760 );
not \U$30509 ( \30762 , \30761 );
and \U$30510 ( \30763 , \30757 , \30762 );
not \U$30511 ( \30764 , \30757 );
and \U$30512 ( \30765 , \30764 , \30761 );
or \U$30513 ( \30766 , \30763 , \30765 );
not \U$30514 ( \30767 , \30282 );
not \U$30515 ( \30768 , \30271 );
or \U$30516 ( \30769 , \30767 , \30768 );
or \U$30517 ( \30770 , \30271 , \30282 );
not \U$30518 ( \30771 , \30262 );
nand \U$30519 ( \30772 , \30770 , \30771 );
nand \U$30520 ( \30773 , \30769 , \30772 );
xor \U$30521 ( \30774 , \30766 , \30773 );
not \U$30522 ( \30775 , \30774 );
not \U$30523 ( \30776 , \30775 );
or \U$30524 ( \30777 , \30753 , \30776 );
nand \U$30525 ( \30778 , \30751 , \30774 );
nand \U$30526 ( \30779 , \30777 , \30778 );
and \U$30527 ( \30780 , \2568 , RIbe2a2f8_86);
or \U$30528 ( \30781 , \4284 , \30780 );
not \U$30529 ( \30782 , RIbe2acd0_107);
nand \U$30530 ( \30783 , \30782 , \4284 );
nand \U$30531 ( \30784 , \30781 , \30783 );
and \U$30532 ( \30785 , \30784 , \2379 );
not \U$30533 ( \30786 , \30784 );
and \U$30534 ( \30787 , \30786 , \25477 );
nor \U$30535 ( \30788 , \30785 , \30787 );
not \U$30536 ( \30789 , \30788 );
not \U$30537 ( \30790 , RIbe2a3e8_88);
not \U$30538 ( \30791 , \20674 );
or \U$30539 ( \30792 , \30790 , \30791 );
nand \U$30540 ( \30793 , \2384 , RIbe2a370_87);
nand \U$30541 ( \30794 , \30792 , \30793 );
and \U$30542 ( \30795 , \30794 , \7038 );
not \U$30543 ( \30796 , \30794 );
and \U$30544 ( \30797 , \30796 , \1276 );
nor \U$30545 ( \30798 , \30795 , \30797 );
not \U$30546 ( \30799 , \30798 );
or \U$30547 ( \30800 , \30789 , \30799 );
or \U$30548 ( \30801 , \30798 , \30788 );
nand \U$30549 ( \30802 , \30800 , \30801 );
not \U$30550 ( \30803 , RIbe2a910_99);
not \U$30551 ( \30804 , \23509 );
or \U$30552 ( \30805 , \30803 , \30804 );
nand \U$30553 ( \30806 , \5467 , RIbe2b5b8_126);
nand \U$30554 ( \30807 , \30805 , \30806 );
and \U$30555 ( \30808 , \30807 , \1125 );
not \U$30556 ( \30809 , \30807 );
and \U$30557 ( \30810 , \30809 , \1131 );
nor \U$30558 ( \30811 , \30808 , \30810 );
xor \U$30559 ( \30812 , \30802 , \30811 );
not \U$30560 ( \30813 , \1152 );
not \U$30561 ( \30814 , RIbe2a190_83);
not \U$30562 ( \30815 , \2597 );
or \U$30563 ( \30816 , \30814 , \30815 );
nand \U$30564 ( \30817 , \1147 , RIbe2a5c8_92);
nand \U$30565 ( \30818 , \30816 , \30817 );
not \U$30566 ( \30819 , \30818 );
and \U$30567 ( \30820 , \30813 , \30819 );
and \U$30568 ( \30821 , \30818 , \1153 );
nor \U$30569 ( \30822 , \30820 , \30821 );
and \U$30570 ( \30823 , \5973 , RIbe2a280_85);
and \U$30571 ( \30824 , \1203 , RIbe2a208_84);
nor \U$30572 ( \30825 , \30823 , \30824 );
and \U$30573 ( \30826 , \30825 , \1011 );
not \U$30574 ( \30827 , \30825 );
and \U$30575 ( \30828 , \30827 , \1608 );
nor \U$30576 ( \30829 , \30826 , \30828 );
xor \U$30577 ( \30830 , \30822 , \30829 );
not \U$30578 ( \30831 , RIbe2a550_91);
not \U$30579 ( \30832 , \5476 );
or \U$30580 ( \30833 , \30831 , \30832 );
nand \U$30581 ( \30834 , \1099 , RIbe2a988_100);
nand \U$30582 ( \30835 , \30833 , \30834 );
and \U$30583 ( \30836 , \30835 , \1082 );
not \U$30584 ( \30837 , \30835 );
and \U$30585 ( \30838 , \30837 , \1309 );
nor \U$30586 ( \30839 , \30836 , \30838 );
xor \U$30587 ( \30840 , \30830 , \30839 );
xor \U$30588 ( \30841 , \30812 , \30840 );
not \U$30589 ( \30842 , RIbe29e48_76);
not \U$30590 ( \30843 , \20764 );
or \U$30591 ( \30844 , \30842 , \30843 );
nand \U$30592 ( \30845 , \4026 , RIbe29dd0_75);
nand \U$30593 ( \30846 , \30844 , \30845 );
and \U$30594 ( \30847 , \30846 , \3698 );
not \U$30595 ( \30848 , \30846 );
and \U$30596 ( \30849 , \30848 , \3471 );
nor \U$30597 ( \30850 , \30847 , \30849 );
not \U$30598 ( \30851 , RIbe29c68_72);
not \U$30599 ( \30852 , \6414 );
or \U$30600 ( \30853 , \30851 , \30852 );
nand \U$30601 ( \30854 , \6418 , RIbe29bf0_71);
nand \U$30602 ( \30855 , \30853 , \30854 );
and \U$30603 ( \30856 , \30855 , \4007 );
not \U$30604 ( \30857 , \30855 );
and \U$30605 ( \30858 , \30857 , \4323 );
nor \U$30606 ( \30859 , \30856 , \30858 );
xor \U$30607 ( \30860 , \30850 , \30859 );
not \U$30608 ( \30861 , RIbe2a028_80);
not \U$30609 ( \30862 , \3283 );
not \U$30610 ( \30863 , \30862 );
or \U$30611 ( \30864 , \30861 , \30863 );
nand \U$30612 ( \30865 , \6800 , RIbe29fb0_79);
nand \U$30613 ( \30866 , \30864 , \30865 );
not \U$30614 ( \30867 , \30866 );
not \U$30615 ( \30868 , \2887 );
and \U$30616 ( \30869 , \30867 , \30868 );
and \U$30617 ( \30870 , \30866 , \3461 );
nor \U$30618 ( \30871 , \30869 , \30870 );
xnor \U$30619 ( \30872 , \30860 , \30871 );
xor \U$30620 ( \30873 , \30841 , \30872 );
not \U$30621 ( \30874 , \30873 );
and \U$30622 ( \30875 , \30779 , \30874 );
not \U$30623 ( \30876 , \30779 );
and \U$30624 ( \30877 , \30876 , \30873 );
nor \U$30625 ( \30878 , \30875 , \30877 );
xor \U$30626 ( \30879 , \30681 , \30878 );
and \U$30627 ( \30880 , \30506 , \30546 );
nor \U$30628 ( \30881 , \30880 , \30477 );
nor \U$30629 ( \30882 , \30506 , \30546 );
nor \U$30630 ( \30883 , \30881 , \30882 );
not \U$30631 ( \30884 , \1374 );
not \U$30632 ( \30885 , RIbe28de0_41);
not \U$30633 ( \30886 , \12811 );
or \U$30634 ( \30887 , \30885 , \30886 );
nand \U$30635 ( \30888 , RIbe29920_65, RIbe2ae38_110);
nand \U$30636 ( \30889 , \30887 , \30888 );
not \U$30637 ( \30890 , RIbe2aeb0_111);
and \U$30638 ( \30891 , \30889 , \30890 );
not \U$30639 ( \30892 , \30889 );
and \U$30640 ( \30893 , \30892 , RIbe2aeb0_111);
nor \U$30641 ( \30894 , \30891 , \30893 );
not \U$30642 ( \30895 , \30894 );
not \U$30643 ( \30896 , \30895 );
or \U$30644 ( \30897 , \30884 , \30896 );
or \U$30645 ( \30898 , \30895 , \1379 );
nand \U$30646 ( \30899 , \30897 , \30898 );
not \U$30647 ( \30900 , RIbe27c10_3);
not \U$30648 ( \30901 , \12887 );
or \U$30649 ( \30902 , \30900 , \30901 );
nand \U$30650 ( \30903 , \12794 , RIbe28e58_42);
nand \U$30651 ( \30904 , \30902 , \30903 );
and \U$30652 ( \30905 , \30904 , \14103 );
not \U$30653 ( \30906 , \30904 );
and \U$30654 ( \30907 , \30906 , \12893 );
nor \U$30655 ( \30908 , \30905 , \30907 );
xor \U$30656 ( \30909 , \30899 , \30908 );
not \U$30657 ( \30910 , \12823 );
not \U$30658 ( \30911 , RIbe27d78_6);
not \U$30659 ( \30912 , \12831 );
or \U$30660 ( \30913 , \30911 , \30912 );
nand \U$30661 ( \30914 , RIbe27d00_5, \12834 );
nand \U$30662 ( \30915 , \30913 , \30914 );
not \U$30663 ( \30916 , \30915 );
or \U$30664 ( \30917 , \30910 , \30916 );
or \U$30665 ( \30918 , \30915 , \12863 );
nand \U$30666 ( \30919 , \30917 , \30918 );
not \U$30667 ( \30920 , RIbe290b0_47);
not \U$30668 ( \30921 , \13074 );
or \U$30669 ( \30922 , \30920 , \30921 );
nand \U$30670 ( \30923 , \12735 , RIbe29a88_68);
nand \U$30671 ( \30924 , \30922 , \30923 );
not \U$30672 ( \30925 , \30924 );
not \U$30673 ( \30926 , \12746 );
or \U$30674 ( \30927 , \30925 , \30926 );
or \U$30675 ( \30928 , \30924 , \15169 );
nand \U$30676 ( \30929 , \30927 , \30928 );
xor \U$30677 ( \30930 , \30919 , \30929 );
not \U$30678 ( \30931 , \12723 );
not \U$30679 ( \30932 , RIbe29038_46);
not \U$30680 ( \30933 , \14523 );
or \U$30681 ( \30934 , \30932 , \30933 );
nand \U$30682 ( \30935 , \13728 , RIbe28fc0_45);
nand \U$30683 ( \30936 , \30934 , \30935 );
not \U$30684 ( \30937 , \30936 );
or \U$30685 ( \30938 , \30931 , \30937 );
or \U$30686 ( \30939 , \30936 , \12723 );
nand \U$30687 ( \30940 , \30938 , \30939 );
xor \U$30688 ( \30941 , \30930 , \30940 );
xor \U$30689 ( \30942 , \30909 , \30941 );
not \U$30690 ( \30943 , \12218 );
not \U$30691 ( \30944 , RIbe28228_16);
not \U$30692 ( \30945 , \10936 );
or \U$30693 ( \30946 , \30944 , \30945 );
nand \U$30694 ( \30947 , \12213 , RIbe281b0_15);
nand \U$30695 ( \30948 , \30946 , \30947 );
not \U$30696 ( \30949 , \30948 );
or \U$30697 ( \30950 , \30943 , \30949 );
or \U$30698 ( \30951 , \30948 , \10943 );
nand \U$30699 ( \30952 , \30950 , \30951 );
not \U$30700 ( \30953 , \12752 );
not \U$30701 ( \30954 , \5494 );
and \U$30702 ( \30955 , \30953 , \30954 );
and \U$30703 ( \30956 , \14725 , RIbe296c8_60);
nor \U$30704 ( \30957 , \30955 , \30956 );
and \U$30705 ( \30958 , \30957 , \14000 );
not \U$30706 ( \30959 , \30957 );
and \U$30707 ( \30960 , \30959 , \12774 );
nor \U$30708 ( \30961 , \30958 , \30960 );
xor \U$30709 ( \30962 , \30952 , \30961 );
not \U$30710 ( \30963 , RIbe280c0_13);
not \U$30711 ( \30964 , \12942 );
or \U$30712 ( \30965 , \30963 , \30964 );
nand \U$30713 ( \30966 , \12947 , RIbe29830_63);
nand \U$30714 ( \30967 , \30965 , \30966 );
and \U$30715 ( \30968 , \30967 , \12195 );
not \U$30716 ( \30969 , \30967 );
and \U$30717 ( \30970 , \30969 , \12957 );
nor \U$30718 ( \30971 , \30968 , \30970 );
xor \U$30719 ( \30972 , \30962 , \30971 );
xor \U$30720 ( \30973 , \30942 , \30972 );
xor \U$30721 ( \30974 , \30883 , \30973 );
not \U$30722 ( \30975 , RIbe28a20_33);
not \U$30723 ( \30976 , \6942 );
or \U$30724 ( \30977 , \30975 , \30976 );
nand \U$30725 ( \30978 , \13158 , RIbe289a8_32);
nand \U$30726 ( \30979 , \30977 , \30978 );
and \U$30727 ( \30980 , \30979 , \7984 );
not \U$30728 ( \30981 , \30979 );
and \U$30729 ( \30982 , \30981 , \9896 );
nor \U$30730 ( \30983 , \30980 , \30982 );
not \U$30731 ( \30984 , \30983 );
not \U$30732 ( \30985 , \30984 );
and \U$30733 ( \30986 , \10915 , RIbe28930_31);
and \U$30734 ( \30987 , \13038 , RIbe29560_57);
nor \U$30735 ( \30988 , \30986 , \30987 );
and \U$30736 ( \30989 , \30988 , \15233 );
not \U$30737 ( \30990 , \30988 );
and \U$30738 ( \30991 , \30990 , \10926 );
nor \U$30739 ( \30992 , \30989 , \30991 );
not \U$30740 ( \30993 , \30992 );
not \U$30741 ( \30994 , \30993 );
or \U$30742 ( \30995 , \30985 , \30994 );
nand \U$30743 ( \30996 , \30992 , \30983 );
nand \U$30744 ( \30997 , \30995 , \30996 );
not \U$30745 ( \30998 , \7301 );
not \U$30746 ( \30999 , RIbe28b88_36);
not \U$30747 ( \31000 , \7299 );
or \U$30748 ( \31001 , \30999 , \31000 );
nand \U$30749 ( \31002 , \6985 , RIbe29290_51);
nand \U$30750 ( \31003 , \31001 , \31002 );
not \U$30751 ( \31004 , \31003 );
or \U$30752 ( \31005 , \30998 , \31004 );
or \U$30753 ( \31006 , \31003 , \13168 );
nand \U$30754 ( \31007 , \31005 , \31006 );
xnor \U$30755 ( \31008 , \30997 , \31007 );
not \U$30756 ( \31009 , \31008 );
not \U$30757 ( \31010 , \6572 );
not \U$30758 ( \31011 , RIbe28390_19);
not \U$30759 ( \31012 , \21608 );
or \U$30760 ( \31013 , \31011 , \31012 );
nand \U$30761 ( \31014 , \6962 , RIbe28b10_35);
nand \U$30762 ( \31015 , \31013 , \31014 );
not \U$30763 ( \31016 , \31015 );
and \U$30764 ( \31017 , \31010 , \31016 );
and \U$30765 ( \31018 , \31015 , \6569 );
nor \U$30766 ( \31019 , \31017 , \31018 );
not \U$30767 ( \31020 , RIbe28480_21);
not \U$30768 ( \31021 , \13238 );
or \U$30769 ( \31022 , \31020 , \31021 );
nand \U$30770 ( \31023 , \7278 , RIbe28408_20);
nand \U$30771 ( \31024 , \31022 , \31023 );
and \U$30772 ( \31025 , \31024 , \6601 );
not \U$30773 ( \31026 , \31024 );
and \U$30774 ( \31027 , \31026 , \6602 );
nor \U$30775 ( \31028 , \31025 , \31027 );
and \U$30776 ( \31029 , \31019 , \31028 );
not \U$30777 ( \31030 , \31019 );
not \U$30778 ( \31031 , \31028 );
and \U$30779 ( \31032 , \31030 , \31031 );
or \U$30780 ( \31033 , \31029 , \31032 );
not \U$30781 ( \31034 , RIbe285e8_24);
not \U$30782 ( \31035 , \6536 );
or \U$30783 ( \31036 , \31034 , \31035 );
nand \U$30784 ( \31037 , \10348 , RIbe287c8_28);
nand \U$30785 ( \31038 , \31036 , \31037 );
and \U$30786 ( \31039 , \31038 , \15730 );
not \U$30787 ( \31040 , \31038 );
and \U$30788 ( \31041 , \31040 , \6888 );
nor \U$30789 ( \31042 , \31039 , \31041 );
xnor \U$30790 ( \31043 , \31033 , \31042 );
not \U$30791 ( \31044 , \31043 );
not \U$30792 ( \31045 , \31044 );
or \U$30793 ( \31046 , \31009 , \31045 );
not \U$30794 ( \31047 , \31008 );
nand \U$30795 ( \31048 , \31047 , \31043 );
nand \U$30796 ( \31049 , \31046 , \31048 );
not \U$30797 ( \31050 , RIbe27fd0_11);
not \U$30798 ( \31051 , \5455 );
or \U$30799 ( \31052 , \31050 , \31051 );
nand \U$30800 ( \31053 , \15885 , RIbe27f58_10);
nand \U$30801 ( \31054 , \31052 , \31053 );
and \U$30802 ( \31055 , \31054 , \10272 );
not \U$30803 ( \31056 , \31054 );
and \U$30804 ( \31057 , \31056 , \6640 );
nor \U$30805 ( \31058 , \31055 , \31057 );
not \U$30806 ( \31059 , \31058 );
not \U$30807 ( \31060 , RIbe27e68_8);
not \U$30808 ( \31061 , \6138 );
or \U$30809 ( \31062 , \31060 , \31061 );
nand \U$30810 ( \31063 , \6859 , RIbe28660_25);
nand \U$30811 ( \31064 , \31062 , \31063 );
not \U$30812 ( \31065 , \31064 );
not \U$30813 ( \31066 , \21090 );
and \U$30814 ( \31067 , \31065 , \31066 );
and \U$30815 ( \31068 , \31064 , \5740 );
nor \U$30816 ( \31069 , \31067 , \31068 );
not \U$30817 ( \31070 , \31069 );
or \U$30818 ( \31071 , \31059 , \31070 );
or \U$30819 ( \31072 , \31058 , \31069 );
nand \U$30820 ( \31073 , \31071 , \31072 );
not \U$30821 ( \31074 , RIbe28f48_44);
not \U$30822 ( \31075 , \5727 );
or \U$30823 ( \31076 , \31074 , \31075 );
nand \U$30824 ( \31077 , \5052 , RIbe28ed0_43);
nand \U$30825 ( \31078 , \31076 , \31077 );
and \U$30826 ( \31079 , \31078 , \4586 );
not \U$30827 ( \31080 , \31078 );
and \U$30828 ( \31081 , \31080 , \4592 );
nor \U$30829 ( \31082 , \31079 , \31081 );
not \U$30830 ( \31083 , \31082 );
and \U$30831 ( \31084 , \31073 , \31083 );
not \U$30832 ( \31085 , \31073 );
and \U$30833 ( \31086 , \31085 , \31082 );
nor \U$30834 ( \31087 , \31084 , \31086 );
and \U$30835 ( \31088 , \31049 , \31087 );
not \U$30836 ( \31089 , \31049 );
not \U$30837 ( \31090 , \31087 );
and \U$30838 ( \31091 , \31089 , \31090 );
nor \U$30839 ( \31092 , \31088 , \31091 );
xor \U$30840 ( \31093 , \30974 , \31092 );
xor \U$30841 ( \31094 , \30879 , \31093 );
not \U$30842 ( \31095 , \30126 );
not \U$30843 ( \31096 , \30141 );
or \U$30844 ( \31097 , \31095 , \31096 );
nand \U$30845 ( \31098 , \31097 , \30132 );
or \U$30846 ( \31099 , \30126 , \30141 );
nand \U$30847 ( \31100 , \31098 , \31099 );
xor \U$30848 ( \31101 , \30108 , \30112 );
and \U$30849 ( \31102 , \31101 , \30117 );
and \U$30850 ( \31103 , \30108 , \30112 );
or \U$30851 ( \31104 , \31102 , \31103 );
xor \U$30852 ( \31105 , \31100 , \31104 );
not \U$30853 ( \31106 , \30153 );
not \U$30854 ( \31107 , \30171 );
or \U$30855 ( \31108 , \31106 , \31107 );
not \U$30856 ( \31109 , \30154 );
not \U$30857 ( \31110 , \30168 );
or \U$30858 ( \31111 , \31109 , \31110 );
nand \U$30859 ( \31112 , \31111 , \30160 );
nand \U$30860 ( \31113 , \31108 , \31112 );
xor \U$30861 ( \31114 , \31105 , \31113 );
xor \U$30862 ( \31115 , \30223 , \30251 );
and \U$30863 ( \31116 , \31115 , \30283 );
and \U$30864 ( \31117 , \30223 , \30251 );
or \U$30865 ( \31118 , \31116 , \31117 );
nand \U$30866 ( \31119 , \30358 , \30322 );
and \U$30867 ( \31120 , \31119 , \30393 );
nor \U$30868 ( \31121 , \30322 , \30358 );
nor \U$30869 ( \31122 , \31120 , \31121 );
and \U$30870 ( \31123 , \30188 , \30186 );
nor \U$30871 ( \31124 , \31123 , \30194 );
nor \U$30872 ( \31125 , \30188 , \30186 );
nor \U$30873 ( \31126 , \31124 , \31125 );
and \U$30874 ( \31127 , \31122 , \31126 );
not \U$30875 ( \31128 , \31122 );
not \U$30876 ( \31129 , \31126 );
and \U$30877 ( \31130 , \31128 , \31129 );
nor \U$30878 ( \31131 , \31127 , \31130 );
xor \U$30879 ( \31132 , \31118 , \31131 );
xor \U$30880 ( \31133 , \31114 , \31132 );
xor \U$30881 ( \31134 , \31094 , \31133 );
xor \U$30882 ( \31135 , \30657 , \31134 );
or \U$30883 ( \31136 , \30090 , \30083 );
not \U$30884 ( \31137 , \31136 );
not \U$30885 ( \31138 , \30095 );
or \U$30886 ( \31139 , \31137 , \31138 );
nand \U$30887 ( \31140 , \30090 , \30083 );
nand \U$30888 ( \31141 , \31139 , \31140 );
not \U$30889 ( \31142 , \30178 );
not \U$30890 ( \31143 , \30102 );
nand \U$30891 ( \31144 , \31142 , \31143 );
and \U$30892 ( \31145 , \31144 , \30395 );
nor \U$30893 ( \31146 , \31142 , \31143 );
nor \U$30894 ( \31147 , \31145 , \31146 );
xor \U$30895 ( \31148 , \31141 , \31147 );
xor \U$30896 ( \31149 , \30411 , \30552 );
and \U$30897 ( \31150 , \31149 , \30567 );
and \U$30898 ( \31151 , \30411 , \30552 );
or \U$30899 ( \31152 , \31150 , \31151 );
xnor \U$30900 ( \31153 , \31148 , \31152 );
xnor \U$30901 ( \31154 , \31135 , \31153 );
buf \U$30902 ( \31155 , \31154 );
and \U$30903 ( \31156 , \30631 , \31155 );
not \U$30904 ( \31157 , \30631 );
not \U$30905 ( \31158 , \31155 );
and \U$30906 ( \31159 , \31157 , \31158 );
nor \U$30907 ( \31160 , \31156 , \31159 );
not \U$30908 ( \31161 , \31160 );
not \U$30909 ( \31162 , \31161 );
or \U$30910 ( \31163 , \30574 , \31162 );
not \U$30911 ( \31164 , \30573 );
nand \U$30912 ( \31165 , \31164 , \31160 );
nand \U$30913 ( \31166 , \31163 , \31165 );
not \U$30914 ( \31167 , \31166 );
xor \U$30915 ( \31168 , \30047 , \30064 );
xor \U$30916 ( \31169 , \31168 , \30069 );
xor \U$30917 ( \31170 , \30049 , \30056 );
xor \U$30918 ( \31171 , \31170 , \30061 );
and \U$30919 ( \31172 , \29033 , \306 );
not \U$30920 ( \31173 , \29033 );
and \U$30921 ( \31174 , \31173 , \313 );
nor \U$30922 ( \31175 , \31172 , \31174 );
not \U$30923 ( \31176 , \31175 );
not \U$30924 ( \31177 , \29026 );
or \U$30925 ( \31178 , \31176 , \31177 );
or \U$30926 ( \31179 , \29026 , \31175 );
nand \U$30927 ( \31180 , \31178 , \31179 );
not \U$30928 ( \31181 , \31180 );
not \U$30929 ( \31182 , \29799 );
not \U$30930 ( \31183 , \29777 );
or \U$30931 ( \31184 , \31182 , \31183 );
not \U$30932 ( \31185 , \29777 );
nand \U$30933 ( \31186 , \31185 , \29798 );
nand \U$30934 ( \31187 , \31184 , \31186 );
buf \U$30935 ( \31188 , \29787 );
xor \U$30936 ( \31189 , \31187 , \31188 );
not \U$30937 ( \31190 , \31189 );
not \U$30938 ( \31191 , \31190 );
or \U$30939 ( \31192 , \31181 , \31191 );
and \U$30940 ( \31193 , \29821 , \29806 );
not \U$30941 ( \31194 , \29821 );
and \U$30942 ( \31195 , \31194 , \29823 );
or \U$30943 ( \31196 , \31193 , \31195 );
buf \U$30944 ( \31197 , \29824 );
and \U$30945 ( \31198 , \31196 , \31197 );
not \U$30946 ( \31199 , \31196 );
not \U$30947 ( \31200 , \31197 );
and \U$30948 ( \31201 , \31199 , \31200 );
nor \U$30949 ( \31202 , \31198 , \31201 );
not \U$30950 ( \31203 , \31180 );
nand \U$30951 ( \31204 , \31203 , \31189 );
nand \U$30952 ( \31205 , \31202 , \31204 );
nand \U$30953 ( \31206 , \31192 , \31205 );
not \U$30954 ( \31207 , \31206 );
nand \U$30955 ( \31208 , \23603 , \23580 );
and \U$30956 ( \31209 , \31208 , \23590 );
nor \U$30957 ( \31210 , \23603 , \23580 );
nor \U$30958 ( \31211 , \31209 , \31210 );
nand \U$30959 ( \31212 , \23657 , \424 );
and \U$30960 ( \31213 , \23671 , \31212 );
nor \U$30961 ( \31214 , \23657 , \1764 );
nor \U$30962 ( \31215 , \31213 , \31214 );
nand \U$30963 ( \31216 , \31211 , \31215 );
not \U$30964 ( \31217 , \23708 );
not \U$30965 ( \31218 , \23693 );
or \U$30966 ( \31219 , \31217 , \31218 );
not \U$30967 ( \31220 , \23690 );
not \U$30968 ( \31221 , \23705 );
or \U$30969 ( \31222 , \31220 , \31221 );
nand \U$30970 ( \31223 , \31222 , \23681 );
nand \U$30971 ( \31224 , \31219 , \31223 );
and \U$30972 ( \31225 , \31216 , \31224 );
nor \U$30973 ( \31226 , \31211 , \31215 );
nor \U$30974 ( \31227 , \31225 , \31226 );
not \U$30975 ( \31228 , \31227 );
nand \U$30976 ( \31229 , \23356 , \23347 );
and \U$30977 ( \31230 , \31229 , \23367 );
nor \U$30978 ( \31231 , \23356 , \23347 );
nor \U$30979 ( \31232 , \31230 , \31231 );
nand \U$30980 ( \31233 , \23492 , \23518 );
and \U$30981 ( \31234 , \31233 , \23503 );
nor \U$30982 ( \31235 , \23492 , \23518 );
nor \U$30983 ( \31236 , \31234 , \31235 );
xor \U$30984 ( \31237 , \31232 , \31236 );
nand \U$30985 ( \31238 , \23429 , \23442 );
and \U$30986 ( \31239 , \31238 , \23419 );
nor \U$30987 ( \31240 , \23429 , \23442 );
nor \U$30988 ( \31241 , \31239 , \31240 );
and \U$30989 ( \31242 , \31237 , \31241 );
and \U$30990 ( \31243 , \31232 , \31236 );
or \U$30991 ( \31244 , \31242 , \31243 );
not \U$30992 ( \31245 , \31244 );
or \U$30993 ( \31246 , \31228 , \31245 );
not \U$30994 ( \31247 , \23476 );
not \U$30995 ( \31248 , \23466 );
or \U$30996 ( \31249 , \31247 , \31248 );
nand \U$30997 ( \31250 , \31249 , \23457 );
not \U$30998 ( \31251 , \23466 );
nand \U$30999 ( \31252 , \31251 , \23477 );
nand \U$31000 ( \31253 , \31250 , \31252 );
not \U$31001 ( \31254 , \23621 );
not \U$31002 ( \31255 , \31254 );
not \U$31003 ( \31256 , \23631 );
or \U$31004 ( \31257 , \31255 , \31256 );
or \U$31005 ( \31258 , \23631 , \31254 );
nand \U$31006 ( \31259 , \31258 , \23644 );
nand \U$31007 ( \31260 , \31257 , \31259 );
xor \U$31008 ( \31261 , \31253 , \31260 );
buf \U$31009 ( \31262 , \23546 );
buf \U$31010 ( \31263 , \23555 );
or \U$31011 ( \31264 , \31262 , \31263 );
nand \U$31012 ( \31265 , \31264 , \23565 );
nand \U$31013 ( \31266 , \31263 , \31262 );
nand \U$31014 ( \31267 , \31265 , \31266 );
and \U$31015 ( \31268 , \31261 , \31267 );
and \U$31016 ( \31269 , \31253 , \31260 );
or \U$31017 ( \31270 , \31268 , \31269 );
nand \U$31018 ( \31271 , \31246 , \31270 );
not \U$31019 ( \31272 , \31244 );
not \U$31020 ( \31273 , \31227 );
nand \U$31021 ( \31274 , \31272 , \31273 );
and \U$31022 ( \31275 , \31271 , \31274 );
nand \U$31023 ( \31276 , \31207 , \31275 );
xor \U$31024 ( \31277 , \29480 , \29463 );
xnor \U$31025 ( \31278 , \31277 , \29473 );
not \U$31026 ( \31279 , RIbe2ab68_104);
not \U$31027 ( \31280 , \3244 );
or \U$31028 ( \31281 , \31279 , \31280 );
nand \U$31029 ( \31282 , \1327 , RIbe2aaf0_103);
nand \U$31030 ( \31283 , \31281 , \31282 );
not \U$31031 ( \31284 , \31283 );
not \U$31032 ( \31285 , \1333 );
and \U$31033 ( \31286 , \31284 , \31285 );
and \U$31034 ( \31287 , \31283 , \6340 );
nor \U$31035 ( \31288 , \31286 , \31287 );
buf \U$31036 ( \31289 , \31288 );
nand \U$31037 ( \31290 , \31278 , \31289 );
xor \U$31038 ( \31291 , \29562 , \29546 );
and \U$31039 ( \31292 , \31291 , \29536 );
not \U$31040 ( \31293 , \31291 );
and \U$31041 ( \31294 , \31293 , \29535 );
nor \U$31042 ( \31295 , \31292 , \31294 );
not \U$31043 ( \31296 , \31295 );
and \U$31044 ( \31297 , \31290 , \31296 );
nor \U$31045 ( \31298 , \31278 , \31289 );
nor \U$31046 ( \31299 , \31297 , \31298 );
not \U$31047 ( \31300 , \31299 );
not \U$31048 ( \31301 , \29727 );
not \U$31049 ( \31302 , \29706 );
or \U$31050 ( \31303 , \31301 , \31302 );
or \U$31051 ( \31304 , \29706 , \29727 );
nand \U$31052 ( \31305 , \31303 , \31304 );
not \U$31053 ( \31306 , \29715 );
and \U$31054 ( \31307 , \31305 , \31306 );
not \U$31055 ( \31308 , \31305 );
and \U$31056 ( \31309 , \31308 , \29715 );
nor \U$31057 ( \31310 , \31307 , \31309 );
not \U$31058 ( \31311 , \31310 );
and \U$31059 ( \31312 , \29495 , \29519 );
not \U$31060 ( \31313 , \29495 );
and \U$31061 ( \31314 , \31313 , \29518 );
or \U$31062 ( \31315 , \31312 , \31314 );
xor \U$31063 ( \31316 , \31315 , \29507 );
nand \U$31064 ( \31317 , \31311 , \31316 );
xor \U$31065 ( \31318 , \29675 , \29684 );
xor \U$31066 ( \31319 , \31318 , \29694 );
and \U$31067 ( \31320 , \31317 , \31319 );
nor \U$31068 ( \31321 , \31311 , \31316 );
nor \U$31069 ( \31322 , \31320 , \31321 );
not \U$31070 ( \31323 , \31322 );
or \U$31071 ( \31324 , \31300 , \31323 );
xor \U$31072 ( \31325 , \29636 , \29647 );
xor \U$31073 ( \31326 , \31325 , \29659 );
not \U$31074 ( \31327 , \31326 );
not \U$31075 ( \31328 , \29621 );
not \U$31076 ( \31329 , \29603 );
or \U$31077 ( \31330 , \31328 , \31329 );
or \U$31078 ( \31331 , \29603 , \29621 );
nand \U$31079 ( \31332 , \31330 , \31331 );
xor \U$31080 ( \31333 , \31332 , \29610 );
not \U$31081 ( \31334 , \31333 );
or \U$31082 ( \31335 , \31327 , \31334 );
not \U$31083 ( \31336 , \29741 );
not \U$31084 ( \31337 , \29759 );
or \U$31085 ( \31338 , \31336 , \31337 );
not \U$31086 ( \31339 , \29759 );
not \U$31087 ( \31340 , \29741 );
nand \U$31088 ( \31341 , \31339 , \31340 );
nand \U$31089 ( \31342 , \31338 , \31341 );
and \U$31090 ( \31343 , \31342 , \29762 );
not \U$31091 ( \31344 , \31342 );
and \U$31092 ( \31345 , \31344 , \29748 );
nor \U$31093 ( \31346 , \31343 , \31345 );
nand \U$31094 ( \31347 , \31335 , \31346 );
not \U$31095 ( \31348 , \31333 );
not \U$31096 ( \31349 , \31326 );
nand \U$31097 ( \31350 , \31348 , \31349 );
nand \U$31098 ( \31351 , \31347 , \31350 );
nand \U$31099 ( \31352 , \31324 , \31351 );
not \U$31100 ( \31353 , \31299 );
not \U$31101 ( \31354 , \31322 );
nand \U$31102 ( \31355 , \31353 , \31354 );
nand \U$31103 ( \31356 , \31352 , \31355 );
and \U$31104 ( \31357 , \31276 , \31356 );
nor \U$31105 ( \31358 , \31207 , \31275 );
nor \U$31106 ( \31359 , \31357 , \31358 );
not \U$31107 ( \31360 , \31359 );
xor \U$31108 ( \31361 , \29901 , \29913 );
xnor \U$31109 ( \31362 , \31361 , \29909 );
xor \U$31110 ( \31363 , \29109 , \29069 );
and \U$31111 ( \31364 , \31363 , \29112 );
not \U$31112 ( \31365 , \31363 );
and \U$31113 ( \31366 , \31365 , \29037 );
or \U$31114 ( \31367 , \31364 , \31366 );
not \U$31115 ( \31368 , \31367 );
nand \U$31116 ( \31369 , \31362 , \31368 );
not \U$31117 ( \31370 , \29523 );
not \U$31118 ( \31371 , \29484 );
or \U$31119 ( \31372 , \31370 , \31371 );
nand \U$31120 ( \31373 , \29485 , \29522 );
nand \U$31121 ( \31374 , \31372 , \31373 );
and \U$31122 ( \31375 , \31374 , \29565 );
not \U$31123 ( \31376 , \31374 );
not \U$31124 ( \31377 , \29565 );
and \U$31125 ( \31378 , \31376 , \31377 );
nor \U$31126 ( \31379 , \31375 , \31378 );
not \U$31127 ( \31380 , \31379 );
not \U$31128 ( \31381 , \29731 );
not \U$31129 ( \31382 , \29765 );
or \U$31130 ( \31383 , \31381 , \31382 );
nand \U$31131 ( \31384 , \29764 , \29730 );
nand \U$31132 ( \31385 , \31383 , \31384 );
not \U$31133 ( \31386 , \29697 );
and \U$31134 ( \31387 , \31385 , \31386 );
not \U$31135 ( \31388 , \31385 );
and \U$31136 ( \31389 , \31388 , \29697 );
nor \U$31137 ( \31390 , \31387 , \31389 );
not \U$31138 ( \31391 , \31390 );
not \U$31139 ( \31392 , \31391 );
or \U$31140 ( \31393 , \31380 , \31392 );
or \U$31141 ( \31394 , \31391 , \31379 );
xor \U$31142 ( \31395 , \29839 , \29848 );
xor \U$31143 ( \31396 , \31395 , \29851 );
nand \U$31144 ( \31397 , \31394 , \31396 );
nand \U$31145 ( \31398 , \31393 , \31397 );
and \U$31146 ( \31399 , \31369 , \31398 );
nor \U$31147 ( \31400 , \31362 , \31368 );
nor \U$31148 ( \31401 , \31399 , \31400 );
not \U$31149 ( \31402 , \31401 );
or \U$31150 ( \31403 , \31360 , \31402 );
xor \U$31151 ( \31404 , \29567 , \29664 );
xor \U$31152 ( \31405 , \31404 , \29768 );
not \U$31153 ( \31406 , \29857 );
not \U$31154 ( \31407 , \29827 );
or \U$31155 ( \31408 , \31406 , \31407 );
nand \U$31156 ( \31409 , \29826 , \29802 );
nand \U$31157 ( \31410 , \31408 , \31409 );
xor \U$31158 ( \31411 , \31410 , \29854 );
xor \U$31159 ( \31412 , \31405 , \31411 );
not \U$31160 ( \31413 , \29862 );
not \U$31161 ( \31414 , \29888 );
or \U$31162 ( \31415 , \31413 , \31414 );
nand \U$31163 ( \31416 , \29887 , \29872 );
nand \U$31164 ( \31417 , \31415 , \31416 );
xor \U$31165 ( \31418 , \31417 , \29885 );
and \U$31166 ( \31419 , \31412 , \31418 );
and \U$31167 ( \31420 , \31405 , \31411 );
or \U$31168 ( \31421 , \31419 , \31420 );
nand \U$31169 ( \31422 , \31403 , \31421 );
not \U$31170 ( \31423 , \31401 );
not \U$31171 ( \31424 , \31359 );
nand \U$31172 ( \31425 , \31423 , \31424 );
nand \U$31173 ( \31426 , \31422 , \31425 );
xor \U$31174 ( \31427 , \31171 , \31426 );
not \U$31175 ( \31428 , \29014 );
not \U$31176 ( \31429 , \29344 );
or \U$31177 ( \31430 , \31428 , \31429 );
or \U$31178 ( \31431 , \29014 , \29344 );
nand \U$31179 ( \31432 , \31430 , \31431 );
not \U$31180 ( \31433 , \29450 );
and \U$31181 ( \31434 , \31432 , \31433 );
not \U$31182 ( \31435 , \31432 );
and \U$31183 ( \31436 , \31435 , \29450 );
nor \U$31184 ( \31437 , \31434 , \31436 );
not \U$31185 ( \31438 , \31437 );
xor \U$31186 ( \31439 , \29771 , \29859 );
xor \U$31187 ( \31440 , \31439 , \29890 );
not \U$31188 ( \31441 , \31440 );
not \U$31189 ( \31442 , \31441 );
or \U$31190 ( \31443 , \31438 , \31442 );
xor \U$31191 ( \31444 , \29916 , \29947 );
xor \U$31192 ( \31445 , \31444 , \29963 );
nand \U$31193 ( \31446 , \31443 , \31445 );
not \U$31194 ( \31447 , \31437 );
nand \U$31195 ( \31448 , \31440 , \31447 );
nand \U$31196 ( \31449 , \31446 , \31448 );
and \U$31197 ( \31450 , \31427 , \31449 );
and \U$31198 ( \31451 , \31171 , \31426 );
or \U$31199 ( \31452 , \31450 , \31451 );
xor \U$31200 ( \31453 , \31169 , \31452 );
xor \U$31201 ( \31454 , \30045 , \30029 );
xor \U$31202 ( \31455 , \31454 , \30034 );
xor \U$31203 ( \31456 , \29972 , \29979 );
xor \U$31204 ( \31457 , \31456 , \30004 );
xor \U$31205 ( \31458 , \31455 , \31457 );
xor \U$31206 ( \31459 , \29454 , \29893 );
xor \U$31207 ( \31460 , \31459 , \29966 );
and \U$31208 ( \31461 , \31458 , \31460 );
and \U$31209 ( \31462 , \31455 , \31457 );
or \U$31210 ( \31463 , \31461 , \31462 );
and \U$31211 ( \31464 , \31453 , \31463 );
and \U$31212 ( \31465 , \31169 , \31452 );
or \U$31213 ( \31466 , \31464 , \31465 );
not \U$31214 ( \31467 , \31466 );
not \U$31215 ( \31468 , \31467 );
xor \U$31216 ( \31469 , \28975 , \30022 );
xor \U$31217 ( \31470 , \31469 , \30570 );
nand \U$31218 ( \31471 , \31468 , \31470 );
nor \U$31219 ( \31472 , \31167 , \31471 );
nor \U$31220 ( \31473 , \27461 , \31472 );
nand \U$31221 ( \31474 , \27436 , \31473 );
not \U$31222 ( \31475 , \25625 );
and \U$31223 ( \31476 , \27419 , \27428 );
not \U$31224 ( \31477 , \31476 );
nor \U$31225 ( \31478 , \27386 , \27406 );
not \U$31226 ( \31479 , \31478 );
or \U$31227 ( \31480 , \31477 , \31479 );
not \U$31228 ( \31481 , \27404 );
not \U$31229 ( \31482 , \27401 );
or \U$31230 ( \31483 , \31481 , \31482 );
nand \U$31231 ( \31484 , \27400 , \27397 );
nand \U$31232 ( \31485 , \31483 , \31484 );
not \U$31233 ( \31486 , \31485 );
nor \U$31234 ( \31487 , \31486 , \27257 );
and \U$31235 ( \31488 , \27324 , \27353 );
not \U$31236 ( \31489 , \31488 );
not \U$31237 ( \31490 , \27385 );
or \U$31238 ( \31491 , \31489 , \31490 );
nand \U$31239 ( \31492 , \27384 , \27358 );
nand \U$31240 ( \31493 , \31491 , \31492 );
and \U$31241 ( \31494 , \31487 , \31493 );
not \U$31242 ( \31495 , \27254 );
not \U$31243 ( \31496 , \27160 );
not \U$31244 ( \31497 , \31496 );
or \U$31245 ( \31498 , \31495 , \31497 );
or \U$31246 ( \31499 , \27254 , \31496 );
nand \U$31247 ( \31500 , \31498 , \31499 );
not \U$31248 ( \31501 , \31500 );
nor \U$31249 ( \31502 , \27400 , \27404 );
not \U$31250 ( \31503 , \31502 );
or \U$31251 ( \31504 , \31501 , \31503 );
nand \U$31252 ( \31505 , \31504 , \27255 );
nor \U$31253 ( \31506 , \31494 , \31505 );
nand \U$31254 ( \31507 , \31480 , \31506 );
not \U$31255 ( \31508 , \31507 );
or \U$31256 ( \31509 , \31475 , \31508 );
not \U$31257 ( \31510 , \27151 );
nor \U$31258 ( \31511 , \31510 , \27149 );
not \U$31259 ( \31512 , \31511 );
not \U$31260 ( \31513 , \27147 );
or \U$31261 ( \31514 , \31512 , \31513 );
nand \U$31262 ( \31515 , \27142 , \27145 );
nand \U$31263 ( \31516 , \31514 , \31515 );
not \U$31264 ( \31517 , \31516 );
and \U$31265 ( \31518 , \27076 , \26911 , \27116 );
not \U$31266 ( \31519 , \31518 );
or \U$31267 ( \31520 , \31517 , \31519 );
not \U$31268 ( \31521 , \26717 );
not \U$31269 ( \31522 , \26907 );
not \U$31270 ( \31523 , \31522 );
or \U$31271 ( \31524 , \31521 , \31523 );
and \U$31272 ( \31525 , \27114 , \27115 );
nand \U$31273 ( \31526 , \31524 , \31525 );
not \U$31274 ( \31527 , \31526 );
not \U$31275 ( \31528 , \26717 );
nand \U$31276 ( \31529 , \31528 , \26907 );
not \U$31277 ( \31530 , \31529 );
or \U$31278 ( \31531 , \31527 , \31530 );
not \U$31279 ( \31532 , \27434 );
and \U$31280 ( \31533 , \26917 , \27075 );
nor \U$31281 ( \31534 , \31532 , \31533 );
nand \U$31282 ( \31535 , \31531 , \31534 );
nand \U$31283 ( \31536 , \31520 , \31535 );
not \U$31284 ( \31537 , \25139 );
buf \U$31285 ( \31538 , \27354 );
nand \U$31286 ( \31539 , \27385 , \31500 , \31538 );
nor \U$31287 ( \31540 , \31537 , \31539 );
not \U$31288 ( \31541 , \24658 );
nand \U$31289 ( \31542 , \25624 , \31485 , \27429 );
nor \U$31290 ( \31543 , \31541 , \31542 );
nand \U$31291 ( \31544 , \31536 , \31540 , \31543 );
nand \U$31292 ( \31545 , \31509 , \31544 );
nor \U$31293 ( \31546 , \31474 , \31545 );
not \U$31294 ( \31547 , \31546 );
or \U$31295 ( \31548 , \27432 , \31547 );
xor \U$31296 ( \31549 , \31232 , \31236 );
xor \U$31297 ( \31550 , \31549 , \31241 );
xor \U$31298 ( \31551 , \31253 , \31260 );
xor \U$31299 ( \31552 , \31551 , \31267 );
xor \U$31300 ( \31553 , \31550 , \31552 );
not \U$31301 ( \31554 , \31289 );
not \U$31302 ( \31555 , \31296 );
or \U$31303 ( \31556 , \31554 , \31555 );
not \U$31304 ( \31557 , \31288 );
nand \U$31305 ( \31558 , \31557 , \31295 );
nand \U$31306 ( \31559 , \31556 , \31558 );
buf \U$31307 ( \31560 , \31278 );
xnor \U$31308 ( \31561 , \31559 , \31560 );
xnor \U$31309 ( \31562 , \31553 , \31561 );
not \U$31310 ( \31563 , \23373 );
not \U$31311 ( \31564 , \31563 );
not \U$31312 ( \31565 , \23383 );
or \U$31313 ( \31566 , \31564 , \31565 );
not \U$31314 ( \31567 , \23383 );
nand \U$31315 ( \31568 , \31567 , \23373 );
nand \U$31316 ( \31569 , \23368 , \31568 );
nand \U$31317 ( \31570 , \31566 , \31569 );
nand \U$31318 ( \31571 , \23570 , \23649 );
and \U$31319 ( \31572 , \31571 , \23610 );
nor \U$31320 ( \31573 , \23570 , \23649 );
nor \U$31321 ( \31574 , \31572 , \31573 );
not \U$31322 ( \31575 , \31574 );
xor \U$31323 ( \31576 , \31570 , \31575 );
not \U$31324 ( \31577 , \23447 );
not \U$31325 ( \31578 , \31577 );
not \U$31326 ( \31579 , \23478 );
or \U$31327 ( \31580 , \31578 , \31579 );
nand \U$31328 ( \31581 , \31580 , \23520 );
or \U$31329 ( \31582 , \23478 , \31577 );
and \U$31330 ( \31583 , \31581 , \31582 );
xnor \U$31331 ( \31584 , \31576 , \31583 );
xor \U$31332 ( \31585 , \31562 , \31584 );
xor \U$31333 ( \31586 , \29576 , \29582 );
xor \U$31334 ( \31587 , \31586 , \29593 );
and \U$31335 ( \31588 , \31319 , \31310 );
not \U$31336 ( \31589 , \31319 );
and \U$31337 ( \31590 , \31589 , \31311 );
nor \U$31338 ( \31591 , \31588 , \31590 );
xor \U$31339 ( \31592 , \31591 , \31316 );
xor \U$31340 ( \31593 , \31587 , \31592 );
not \U$31341 ( \31594 , \31333 );
not \U$31342 ( \31595 , \31346 );
or \U$31343 ( \31596 , \31594 , \31595 );
or \U$31344 ( \31597 , \31333 , \31346 );
nand \U$31345 ( \31598 , \31596 , \31597 );
and \U$31346 ( \31599 , \31598 , \31349 );
not \U$31347 ( \31600 , \31598 );
and \U$31348 ( \31601 , \31600 , \31326 );
nor \U$31349 ( \31602 , \31599 , \31601 );
xnor \U$31350 ( \31603 , \31593 , \31602 );
xor \U$31351 ( \31604 , \31585 , \31603 );
nand \U$31352 ( \31605 , \23332 , \23311 );
not \U$31353 ( \31606 , \31605 );
xor \U$31354 ( \31607 , \31215 , \31211 );
xor \U$31355 ( \31608 , \31607 , \31224 );
not \U$31356 ( \31609 , \31608 );
and \U$31357 ( \31610 , \31606 , \31609 );
and \U$31358 ( \31611 , \31605 , \31608 );
nor \U$31359 ( \31612 , \31610 , \31611 );
not \U$31360 ( \31613 , \31612 );
not \U$31361 ( \31614 , \23389 );
not \U$31362 ( \31615 , \23525 );
or \U$31363 ( \31616 , \31614 , \31615 );
nand \U$31364 ( \31617 , \31616 , \23406 );
nand \U$31365 ( \31618 , \23526 , \23388 );
nand \U$31366 ( \31619 , \31617 , \31618 );
not \U$31367 ( \31620 , \31619 );
or \U$31368 ( \31621 , \31613 , \31620 );
or \U$31369 ( \31622 , \31619 , \31612 );
nand \U$31370 ( \31623 , \31621 , \31622 );
not \U$31371 ( \31624 , \31623 );
not \U$31372 ( \31625 , \23404 );
not \U$31373 ( \31626 , \23399 );
or \U$31374 ( \31627 , \31625 , \31626 );
nand \U$31375 ( \31628 , \31627 , \23395 );
or \U$31376 ( \31629 , \23399 , \23404 );
nand \U$31377 ( \31630 , \31628 , \31629 );
xor \U$31378 ( \31631 , \23318 , \23326 );
and \U$31379 ( \31632 , \31631 , \23331 );
and \U$31380 ( \31633 , \23318 , \23326 );
or \U$31381 ( \31634 , \31632 , \31633 );
xor \U$31382 ( \31635 , \31630 , \31634 );
not \U$31383 ( \31636 , \23300 );
not \U$31384 ( \31637 , \31636 );
not \U$31385 ( \31638 , \23304 );
or \U$31386 ( \31639 , \31637 , \31638 );
nand \U$31387 ( \31640 , \31639 , \23310 );
nand \U$31388 ( \31641 , \23305 , \23300 );
nand \U$31389 ( \31642 , \31640 , \31641 );
xnor \U$31390 ( \31643 , \31635 , \31642 );
nand \U$31391 ( \31644 , \31624 , \31643 );
and \U$31392 ( \31645 , \31604 , \31644 );
nor \U$31393 ( \31646 , \31624 , \31643 );
nor \U$31394 ( \31647 , \31645 , \31646 );
not \U$31395 ( \31648 , \23273 );
not \U$31396 ( \31649 , \23265 );
or \U$31397 ( \31650 , \31648 , \31649 );
not \U$31398 ( \31651 , \23265 );
nand \U$31399 ( \31652 , \31651 , \23274 );
nand \U$31400 ( \31653 , \31652 , \23285 );
nand \U$31401 ( \31654 , \31650 , \31653 );
not \U$31402 ( \31655 , \31654 );
and \U$31403 ( \31656 , \23784 , \23719 );
nor \U$31404 ( \31657 , \31656 , \23753 );
nor \U$31405 ( \31658 , \23719 , \23784 );
nor \U$31406 ( \31659 , \31657 , \31658 );
and \U$31407 ( \31660 , \31655 , \31659 );
or \U$31408 ( \31661 , \23333 , \23294 );
and \U$31409 ( \31662 , \31661 , \23530 );
and \U$31410 ( \31663 , \23294 , \23333 );
nor \U$31411 ( \31664 , \31662 , \31663 );
nor \U$31412 ( \31665 , \31660 , \31664 );
nor \U$31413 ( \31666 , \31655 , \31659 );
nor \U$31414 ( \31667 , \31665 , \31666 );
xor \U$31415 ( \31668 , \31647 , \31667 );
xnor \U$31416 ( \31669 , \31270 , \31273 );
and \U$31417 ( \31670 , \31669 , \31244 );
not \U$31418 ( \31671 , \31669 );
and \U$31419 ( \31672 , \31671 , \31272 );
nor \U$31420 ( \31673 , \31670 , \31672 );
xor \U$31421 ( \31674 , \31299 , \31354 );
xnor \U$31422 ( \31675 , \31674 , \31351 );
xor \U$31423 ( \31676 , \31673 , \31675 );
xor \U$31424 ( \31677 , \31180 , \31190 );
xor \U$31425 ( \31678 , \31677 , \31202 );
xor \U$31426 ( \31679 , \31676 , \31678 );
not \U$31427 ( \31680 , \31642 );
not \U$31428 ( \31681 , \31634 );
or \U$31429 ( \31682 , \31680 , \31681 );
or \U$31430 ( \31683 , \31634 , \31642 );
nand \U$31431 ( \31684 , \31683 , \31630 );
nand \U$31432 ( \31685 , \31682 , \31684 );
not \U$31433 ( \31686 , \31582 );
not \U$31434 ( \31687 , \31581 );
or \U$31435 ( \31688 , \31686 , \31687 );
not \U$31436 ( \31689 , \31570 );
nand \U$31437 ( \31690 , \31689 , \31574 );
nand \U$31438 ( \31691 , \31688 , \31690 );
nand \U$31439 ( \31692 , \31575 , \31570 );
nand \U$31440 ( \31693 , \31691 , \31692 );
xor \U$31441 ( \31694 , \31685 , \31693 );
not \U$31442 ( \31695 , \31587 );
not \U$31443 ( \31696 , \31602 );
or \U$31444 ( \31697 , \31695 , \31696 );
or \U$31445 ( \31698 , \31602 , \31587 );
not \U$31446 ( \31699 , \31592 );
nand \U$31447 ( \31700 , \31698 , \31699 );
nand \U$31448 ( \31701 , \31697 , \31700 );
xor \U$31449 ( \31702 , \31694 , \31701 );
not \U$31450 ( \31703 , \31702 );
xor \U$31451 ( \31704 , \29624 , \29661 );
xnor \U$31452 ( \31705 , \31704 , \29596 );
not \U$31453 ( \31706 , \31561 );
not \U$31454 ( \31707 , \31550 );
not \U$31455 ( \31708 , \31707 );
or \U$31456 ( \31709 , \31706 , \31708 );
or \U$31457 ( \31710 , \31707 , \31561 );
nand \U$31458 ( \31711 , \31710 , \31552 );
nand \U$31459 ( \31712 , \31709 , \31711 );
xor \U$31460 ( \31713 , \31705 , \31712 );
not \U$31461 ( \31714 , \31379 );
not \U$31462 ( \31715 , \31714 );
not \U$31463 ( \31716 , \31391 );
or \U$31464 ( \31717 , \31715 , \31716 );
nand \U$31465 ( \31718 , \31390 , \31379 );
nand \U$31466 ( \31719 , \31717 , \31718 );
not \U$31467 ( \31720 , \31396 );
and \U$31468 ( \31721 , \31719 , \31720 );
not \U$31469 ( \31722 , \31719 );
and \U$31470 ( \31723 , \31722 , \31396 );
nor \U$31471 ( \31724 , \31721 , \31723 );
xnor \U$31472 ( \31725 , \31713 , \31724 );
not \U$31473 ( \31726 , \31725 );
or \U$31474 ( \31727 , \31703 , \31726 );
or \U$31475 ( \31728 , \31725 , \31702 );
nand \U$31476 ( \31729 , \31727 , \31728 );
xor \U$31477 ( \31730 , \31679 , \31729 );
xor \U$31478 ( \31731 , \31668 , \31730 );
not \U$31479 ( \31732 , \23731 );
and \U$31480 ( \31733 , \31732 , \23749 );
nor \U$31481 ( \31734 , \31733 , \23737 );
nor \U$31482 ( \31735 , \31732 , \23749 );
nor \U$31483 ( \31736 , \31734 , \31735 );
not \U$31484 ( \31737 , \31736 );
not \U$31485 ( \31738 , \23672 );
nand \U$31486 ( \31739 , \31738 , \23710 );
and \U$31487 ( \31740 , \23650 , \31739 );
and \U$31488 ( \31741 , \23713 , \23672 );
nor \U$31489 ( \31742 , \31740 , \31741 );
not \U$31490 ( \31743 , \31742 );
or \U$31491 ( \31744 , \31737 , \31743 );
not \U$31492 ( \31745 , \23773 );
not \U$31493 ( \31746 , \23780 );
or \U$31494 ( \31747 , \31745 , \31746 );
nand \U$31495 ( \31748 , \31747 , \23763 );
or \U$31496 ( \31749 , \23773 , \23780 );
nand \U$31497 ( \31750 , \31748 , \31749 );
nand \U$31498 ( \31751 , \31744 , \31750 );
not \U$31499 ( \31752 , \31742 );
not \U$31500 ( \31753 , \31736 );
nand \U$31501 ( \31754 , \31752 , \31753 );
nand \U$31502 ( \31755 , \31751 , \31754 );
not \U$31503 ( \31756 , \31608 );
nand \U$31504 ( \31757 , \31756 , \31605 );
not \U$31505 ( \31758 , \31757 );
not \U$31506 ( \31759 , \31619 );
or \U$31507 ( \31760 , \31758 , \31759 );
nand \U$31508 ( \31761 , \23332 , \23311 , \31608 );
nand \U$31509 ( \31762 , \31760 , \31761 );
xor \U$31510 ( \31763 , \31755 , \31762 );
xor \U$31511 ( \31764 , \31562 , \31584 );
and \U$31512 ( \31765 , \31764 , \31603 );
and \U$31513 ( \31766 , \31562 , \31584 );
or \U$31514 ( \31767 , \31765 , \31766 );
xor \U$31515 ( \31768 , \31763 , \31767 );
buf \U$31516 ( \31769 , \31659 );
not \U$31517 ( \31770 , \31769 );
not \U$31518 ( \31771 , \31654 );
not \U$31519 ( \31772 , \31664 );
or \U$31520 ( \31773 , \31771 , \31772 );
or \U$31521 ( \31774 , \31664 , \31654 );
nand \U$31522 ( \31775 , \31773 , \31774 );
not \U$31523 ( \31776 , \31775 );
or \U$31524 ( \31777 , \31770 , \31776 );
or \U$31525 ( \31778 , \31775 , \31769 );
nand \U$31526 ( \31779 , \31777 , \31778 );
not \U$31527 ( \31780 , \31604 );
not \U$31528 ( \31781 , \31623 );
not \U$31529 ( \31782 , \31643 );
and \U$31530 ( \31783 , \31781 , \31782 );
and \U$31531 ( \31784 , \31623 , \31643 );
nor \U$31532 ( \31785 , \31783 , \31784 );
not \U$31533 ( \31786 , \31785 );
or \U$31534 ( \31787 , \31780 , \31786 );
or \U$31535 ( \31788 , \31785 , \31604 );
nand \U$31536 ( \31789 , \31787 , \31788 );
nand \U$31537 ( \31790 , \31779 , \31789 );
xor \U$31538 ( \31791 , \31768 , \31790 );
not \U$31539 ( \31792 , \31742 );
and \U$31540 ( \31793 , \31750 , \31736 );
not \U$31541 ( \31794 , \31750 );
and \U$31542 ( \31795 , \31794 , \31753 );
nor \U$31543 ( \31796 , \31793 , \31795 );
not \U$31544 ( \31797 , \31796 );
not \U$31545 ( \31798 , \31797 );
or \U$31546 ( \31799 , \31792 , \31798 );
not \U$31547 ( \31800 , \31742 );
nand \U$31548 ( \31801 , \31800 , \31796 );
nand \U$31549 ( \31802 , \31799 , \31801 );
not \U$31550 ( \31803 , \31802 );
not \U$31551 ( \31804 , \23535 );
not \U$31552 ( \31805 , \23531 );
or \U$31553 ( \31806 , \31804 , \31805 );
not \U$31554 ( \31807 , \23286 );
not \U$31555 ( \31808 , \23534 );
or \U$31556 ( \31809 , \31807 , \31808 );
nand \U$31557 ( \31810 , \31809 , \23789 );
nand \U$31558 ( \31811 , \31806 , \31810 );
not \U$31559 ( \31812 , \31811 );
or \U$31560 ( \31813 , \31803 , \31812 );
or \U$31561 ( \31814 , \31811 , \31802 );
xor \U$31562 ( \31815 , \23234 , \23238 );
and \U$31563 ( \31816 , \31815 , \23243 );
and \U$31564 ( \31817 , \23234 , \23238 );
or \U$31565 ( \31818 , \31816 , \31817 );
not \U$31566 ( \31819 , \31818 );
nand \U$31567 ( \31820 , \31814 , \31819 );
nand \U$31568 ( \31821 , \31813 , \31820 );
xnor \U$31569 ( \31822 , \31791 , \31821 );
and \U$31570 ( \31823 , \31731 , \31822 );
not \U$31571 ( \31824 , \31823 );
not \U$31572 ( \31825 , \31821 );
not \U$31573 ( \31826 , \31768 );
nand \U$31574 ( \31827 , \31825 , \31826 );
not \U$31575 ( \31828 , \31790 );
and \U$31576 ( \31829 , \31827 , \31828 );
nor \U$31577 ( \31830 , \31825 , \31826 );
nor \U$31578 ( \31831 , \31829 , \31830 );
not \U$31579 ( \31832 , \31831 );
nand \U$31580 ( \31833 , \31647 , \31667 );
and \U$31581 ( \31834 , \31833 , \31730 );
nor \U$31582 ( \31835 , \31647 , \31667 );
nor \U$31583 ( \31836 , \31834 , \31835 );
not \U$31584 ( \31837 , \31836 );
xor \U$31585 ( \31838 , \31685 , \31693 );
and \U$31586 ( \31839 , \31838 , \31701 );
and \U$31587 ( \31840 , \31685 , \31693 );
or \U$31588 ( \31841 , \31839 , \31840 );
not \U$31589 ( \31842 , \31705 );
not \U$31590 ( \31843 , \31712 );
not \U$31591 ( \31844 , \31843 );
or \U$31592 ( \31845 , \31842 , \31844 );
not \U$31593 ( \31846 , \31724 );
nand \U$31594 ( \31847 , \31845 , \31846 );
not \U$31595 ( \31848 , \31705 );
nand \U$31596 ( \31849 , \31848 , \31712 );
nand \U$31597 ( \31850 , \31847 , \31849 );
xor \U$31598 ( \31851 , \31841 , \31850 );
xor \U$31599 ( \31852 , \31673 , \31675 );
and \U$31600 ( \31853 , \31852 , \31678 );
and \U$31601 ( \31854 , \31673 , \31675 );
or \U$31602 ( \31855 , \31853 , \31854 );
xor \U$31603 ( \31856 , \31851 , \31855 );
not \U$31604 ( \31857 , \31856 );
and \U$31605 ( \31858 , \31837 , \31857 );
and \U$31606 ( \31859 , \31836 , \31856 );
nor \U$31607 ( \31860 , \31858 , \31859 );
not \U$31608 ( \31861 , \31860 );
not \U$31609 ( \31862 , \31356 );
not \U$31610 ( \31863 , \31275 );
and \U$31611 ( \31864 , \31862 , \31863 );
and \U$31612 ( \31865 , \31356 , \31275 );
nor \U$31613 ( \31866 , \31864 , \31865 );
and \U$31614 ( \31867 , \31866 , \31207 );
not \U$31615 ( \31868 , \31866 );
not \U$31616 ( \31869 , \31207 );
and \U$31617 ( \31870 , \31868 , \31869 );
nor \U$31618 ( \31871 , \31867 , \31870 );
xor \U$31619 ( \31872 , \31367 , \31398 );
xnor \U$31620 ( \31873 , \31872 , \31362 );
xor \U$31621 ( \31874 , \31871 , \31873 );
xor \U$31622 ( \31875 , \31405 , \31411 );
xor \U$31623 ( \31876 , \31875 , \31418 );
xor \U$31624 ( \31877 , \31874 , \31876 );
not \U$31625 ( \31878 , \31877 );
not \U$31626 ( \31879 , \31725 );
nand \U$31627 ( \31880 , \31879 , \31702 );
not \U$31628 ( \31881 , \31702 );
not \U$31629 ( \31882 , \31881 );
not \U$31630 ( \31883 , \31725 );
or \U$31631 ( \31884 , \31882 , \31883 );
nand \U$31632 ( \31885 , \31884 , \31679 );
nand \U$31633 ( \31886 , \31880 , \31885 );
not \U$31634 ( \31887 , \31886 );
not \U$31635 ( \31888 , \31762 );
not \U$31636 ( \31889 , \31755 );
nand \U$31637 ( \31890 , \31888 , \31889 );
and \U$31638 ( \31891 , \31890 , \31767 );
nor \U$31639 ( \31892 , \31888 , \31889 );
nor \U$31640 ( \31893 , \31891 , \31892 );
not \U$31641 ( \31894 , \31893 );
and \U$31642 ( \31895 , \31887 , \31894 );
and \U$31643 ( \31896 , \31886 , \31893 );
nor \U$31644 ( \31897 , \31895 , \31896 );
not \U$31645 ( \31898 , \31897 );
or \U$31646 ( \31899 , \31878 , \31898 );
or \U$31647 ( \31900 , \31897 , \31877 );
nand \U$31648 ( \31901 , \31899 , \31900 );
not \U$31649 ( \31902 , \31901 );
or \U$31650 ( \31903 , \31861 , \31902 );
or \U$31651 ( \31904 , \31860 , \31901 );
nand \U$31652 ( \31905 , \31903 , \31904 );
not \U$31653 ( \31906 , \31905 );
or \U$31654 ( \31907 , \31832 , \31906 );
or \U$31655 ( \31908 , \31831 , \31905 );
nand \U$31656 ( \31909 , \31907 , \31908 );
not \U$31657 ( \31910 , \31909 );
not \U$31658 ( \31911 , \31910 );
or \U$31659 ( \31912 , \31824 , \31911 );
not \U$31660 ( \31913 , \31823 );
nand \U$31661 ( \31914 , \31913 , \31909 );
nand \U$31662 ( \31915 , \31912 , \31914 );
not \U$31663 ( \31916 , \31831 );
nand \U$31664 ( \31917 , \31916 , \31905 );
not \U$31665 ( \31918 , \31917 );
not \U$31666 ( \31919 , \31856 );
nand \U$31667 ( \31920 , \31836 , \31919 );
and \U$31668 ( \31921 , \31901 , \31920 );
nor \U$31669 ( \31922 , \31836 , \31919 );
nor \U$31670 ( \31923 , \31921 , \31922 );
xor \U$31671 ( \31924 , \31421 , \31401 );
xnor \U$31672 ( \31925 , \31924 , \31424 );
not \U$31673 ( \31926 , \31925 );
not \U$31674 ( \31927 , \31926 );
not \U$31675 ( \31928 , \31893 );
or \U$31676 ( \31929 , \31877 , \31928 );
nand \U$31677 ( \31930 , \31929 , \31886 );
nand \U$31678 ( \31931 , \31877 , \31928 );
nand \U$31679 ( \31932 , \31930 , \31931 );
not \U$31680 ( \31933 , \31932 );
or \U$31681 ( \31934 , \31927 , \31933 );
nand \U$31682 ( \31935 , \31930 , \31931 , \31925 );
nand \U$31683 ( \31936 , \31934 , \31935 );
not \U$31684 ( \31937 , \31850 );
not \U$31685 ( \31938 , \31841 );
or \U$31686 ( \31939 , \31937 , \31938 );
or \U$31687 ( \31940 , \31841 , \31850 );
nand \U$31688 ( \31941 , \31940 , \31855 );
nand \U$31689 ( \31942 , \31939 , \31941 );
xor \U$31690 ( \31943 , \31871 , \31873 );
and \U$31691 ( \31944 , \31943 , \31876 );
and \U$31692 ( \31945 , \31871 , \31873 );
or \U$31693 ( \31946 , \31944 , \31945 );
xor \U$31694 ( \31947 , \31942 , \31946 );
not \U$31695 ( \31948 , \31437 );
not \U$31696 ( \31949 , \31948 );
not \U$31697 ( \31950 , \31441 );
or \U$31698 ( \31951 , \31949 , \31950 );
nand \U$31699 ( \31952 , \31440 , \31437 );
nand \U$31700 ( \31953 , \31951 , \31952 );
xnor \U$31701 ( \31954 , \31953 , \31445 );
xor \U$31702 ( \31955 , \31947 , \31954 );
not \U$31703 ( \31956 , \31955 );
and \U$31704 ( \31957 , \31936 , \31956 );
not \U$31705 ( \31958 , \31936 );
and \U$31706 ( \31959 , \31958 , \31955 );
nor \U$31707 ( \31960 , \31957 , \31959 );
and \U$31708 ( \31961 , \31923 , \31960 );
not \U$31709 ( \31962 , \31923 );
not \U$31710 ( \31963 , \31960 );
and \U$31711 ( \31964 , \31962 , \31963 );
nor \U$31712 ( \31965 , \31961 , \31964 );
not \U$31713 ( \31966 , \31965 );
not \U$31714 ( \31967 , \31966 );
or \U$31715 ( \31968 , \31918 , \31967 );
not \U$31716 ( \31969 , \31917 );
nand \U$31717 ( \31970 , \31965 , \31969 );
nand \U$31718 ( \31971 , \31968 , \31970 );
not \U$31719 ( \31972 , \31923 );
nand \U$31720 ( \31973 , \31972 , \31960 );
not \U$31721 ( \31974 , \31973 );
not \U$31722 ( \31975 , \31974 );
nand \U$31723 ( \31976 , \31955 , \31926 );
and \U$31724 ( \31977 , \31976 , \31932 );
nor \U$31725 ( \31978 , \31955 , \31926 );
nor \U$31726 ( \31979 , \31977 , \31978 );
not \U$31727 ( \31980 , \31979 );
not \U$31728 ( \31981 , \31980 );
xor \U$31729 ( \31982 , \31171 , \31426 );
xor \U$31730 ( \31983 , \31982 , \31449 );
not \U$31731 ( \31984 , \31942 );
nand \U$31732 ( \31985 , \31984 , \31954 );
not \U$31733 ( \31986 , \31985 );
not \U$31734 ( \31987 , \31946 );
or \U$31735 ( \31988 , \31986 , \31987 );
not \U$31736 ( \31989 , \31954 );
nand \U$31737 ( \31990 , \31989 , \31942 );
nand \U$31738 ( \31991 , \31988 , \31990 );
xor \U$31739 ( \31992 , \31983 , \31991 );
xor \U$31740 ( \31993 , \31455 , \31457 );
xor \U$31741 ( \31994 , \31993 , \31460 );
xor \U$31742 ( \31995 , \31992 , \31994 );
not \U$31743 ( \31996 , \31995 );
not \U$31744 ( \31997 , \31996 );
or \U$31745 ( \31998 , \31981 , \31997 );
nand \U$31746 ( \31999 , \31995 , \31979 );
nand \U$31747 ( \32000 , \31998 , \31999 );
not \U$31748 ( \32001 , \32000 );
not \U$31749 ( \32002 , \32001 );
or \U$31750 ( \32003 , \31975 , \32002 );
nand \U$31751 ( \32004 , \32000 , \31973 );
nand \U$31752 ( \32005 , \32003 , \32004 );
xor \U$31753 ( \32006 , \31731 , \31822 );
not \U$31754 ( \32007 , \32006 );
not \U$31755 ( \32008 , \32007 );
not \U$31756 ( \32009 , \31779 );
xor \U$31757 ( \32010 , \31789 , \32009 );
and \U$31758 ( \32011 , \31802 , \31819 );
not \U$31759 ( \32012 , \31802 );
and \U$31760 ( \32013 , \32012 , \31818 );
nor \U$31761 ( \32014 , \32011 , \32013 );
xnor \U$31762 ( \32015 , \32014 , \31811 );
xor \U$31763 ( \32016 , \32010 , \32015 );
xor \U$31764 ( \32017 , \23253 , \23257 );
and \U$31765 ( \32018 , \32017 , \23794 );
and \U$31766 ( \32019 , \23253 , \23257 );
or \U$31767 ( \32020 , \32018 , \32019 );
and \U$31768 ( \32021 , \32016 , \32020 );
and \U$31769 ( \32022 , \32010 , \32015 );
or \U$31770 ( \32023 , \32021 , \32022 );
not \U$31771 ( \32024 , \32023 );
not \U$31772 ( \32025 , \32024 );
or \U$31773 ( \32026 , \32008 , \32025 );
nand \U$31774 ( \32027 , \32006 , \32023 );
nand \U$31775 ( \32028 , \32026 , \32027 );
buf \U$31776 ( \32029 , \32028 );
nand \U$31777 ( \32030 , \31915 , \31971 , \32005 , \32029 );
not \U$31778 ( \32031 , \29969 );
not \U$31779 ( \32032 , \30008 );
and \U$31780 ( \32033 , \32031 , \32032 );
and \U$31781 ( \32034 , \29969 , \30008 );
nor \U$31782 ( \32035 , \32033 , \32034 );
not \U$31783 ( \32036 , \32035 );
xor \U$31784 ( \32037 , \30018 , \32036 );
xor \U$31785 ( \32038 , \31169 , \31452 );
xor \U$31786 ( \32039 , \32038 , \31463 );
xor \U$31787 ( \32040 , \32037 , \32039 );
xor \U$31788 ( \32041 , \31983 , \31991 );
and \U$31789 ( \32042 , \32041 , \31994 );
and \U$31790 ( \32043 , \31983 , \31991 );
or \U$31791 ( \32044 , \32042 , \32043 );
and \U$31792 ( \32045 , \32040 , \32044 );
and \U$31793 ( \32046 , \32037 , \32039 );
or \U$31794 ( \32047 , \32045 , \32046 );
not \U$31795 ( \32048 , \32047 );
not \U$31796 ( \32049 , \31467 );
not \U$31797 ( \32050 , \31470 );
or \U$31798 ( \32051 , \32049 , \32050 );
or \U$31799 ( \32052 , \31467 , \31470 );
nand \U$31800 ( \32053 , \32051 , \32052 );
not \U$31801 ( \32054 , \32053 );
not \U$31802 ( \32055 , \32054 );
or \U$31803 ( \32056 , \32048 , \32055 );
not \U$31804 ( \32057 , \32047 );
nand \U$31805 ( \32058 , \32057 , \32053 );
nand \U$31806 ( \32059 , \32056 , \32058 );
nand \U$31807 ( \32060 , \31980 , \31995 );
not \U$31808 ( \32061 , \32060 );
xor \U$31809 ( \32062 , \32037 , \32039 );
xor \U$31810 ( \32063 , \32062 , \32044 );
not \U$31811 ( \32064 , \32063 );
or \U$31812 ( \32065 , \32061 , \32064 );
or \U$31813 ( \32066 , \32063 , \32060 );
nand \U$31814 ( \32067 , \32065 , \32066 );
xor \U$31815 ( \32068 , \32010 , \32015 );
xor \U$31816 ( \32069 , \32068 , \32020 );
buf \U$31817 ( \32070 , \23795 );
and \U$31818 ( \32071 , \32070 , \23244 );
nor \U$31819 ( \32072 , \32071 , \23248 );
nor \U$31820 ( \32073 , \32070 , \23244 );
nor \U$31821 ( \32074 , \32072 , \32073 );
xor \U$31822 ( \32075 , \32069 , \32074 );
nand \U$31823 ( \32076 , \32059 , \32067 , \32075 );
not \U$31824 ( \32077 , \31166 );
not \U$31825 ( \32078 , \31471 );
and \U$31826 ( \32079 , \32077 , \32078 );
and \U$31827 ( \32080 , \31166 , \31471 );
nor \U$31828 ( \32081 , \32079 , \32080 );
or \U$31829 ( \32082 , \32030 , \32076 , \32081 );
not \U$31830 ( \32083 , \31472 );
nand \U$31831 ( \32084 , \32082 , \32083 );
nand \U$31832 ( \32085 , \31548 , \32084 );
nor \U$31833 ( \32086 , \32069 , \32074 );
nand \U$31834 ( \32087 , \32028 , \32086 );
nand \U$31835 ( \32088 , \31909 , \31823 );
nand \U$31836 ( \32089 , \32006 , \32024 );
nand \U$31837 ( \32090 , \32087 , \32088 , \32089 );
and \U$31838 ( \32091 , \31971 , \32090 );
not \U$31839 ( \32092 , \31969 );
not \U$31840 ( \32093 , \31966 );
or \U$31841 ( \32094 , \32092 , \32093 );
nand \U$31842 ( \32095 , \31974 , \32000 );
nand \U$31843 ( \32096 , \32094 , \32095 );
nor \U$31844 ( \32097 , \32091 , \32096 );
not \U$31845 ( \32098 , \32060 );
nand \U$31846 ( \32099 , \32098 , \32063 );
nand \U$31847 ( \32100 , \32053 , \32047 );
and \U$31848 ( \32101 , \32099 , \32100 );
nand \U$31849 ( \32102 , \32097 , \32101 );
not \U$31850 ( \32103 , \32100 );
nor \U$31851 ( \32104 , \32103 , \32059 );
nor \U$31852 ( \32105 , \32104 , \32081 );
and \U$31853 ( \32106 , \32102 , \32105 );
not \U$31854 ( \32107 , \32063 );
nand \U$31855 ( \32108 , \32107 , \32060 );
not \U$31856 ( \32109 , \32108 );
not \U$31857 ( \32110 , \32088 );
nor \U$31858 ( \32111 , \31915 , \32110 );
not \U$31859 ( \32112 , \32096 );
and \U$31860 ( \32113 , \32111 , \32112 );
not \U$31861 ( \32114 , \32095 );
nor \U$31862 ( \32115 , \32114 , \32005 );
nor \U$31863 ( \32116 , \32113 , \32115 );
not \U$31864 ( \32117 , \32116 );
or \U$31865 ( \32118 , \32109 , \32117 );
nand \U$31866 ( \32119 , \32118 , \32101 );
nand \U$31867 ( \32120 , \32106 , \32119 );
nand \U$31868 ( \32121 , \32085 , \32120 );
not \U$31869 ( \32122 , \32121 );
not \U$31870 ( \32123 , RIbe29c68_72);
not \U$31871 ( \32124 , \30862 );
or \U$31872 ( \32125 , \32123 , \32124 );
nand \U$31873 ( \32126 , RIbe29bf0_71, \3689 );
nand \U$31874 ( \32127 , \32125 , \32126 );
xor \U$31875 ( \32128 , \32127 , \2887 );
not \U$31876 ( \32129 , \4059 );
not \U$31877 ( \32130 , RIbe29e48_76);
not \U$31878 ( \32131 , \7827 );
or \U$31879 ( \32132 , \32130 , \32131 );
nand \U$31880 ( \32133 , \4284 , RIbe29dd0_75);
nand \U$31881 ( \32134 , \32132 , \32133 );
not \U$31882 ( \32135 , \32134 );
and \U$31883 ( \32136 , \32129 , \32135 );
and \U$31884 ( \32137 , \32134 , \2576 );
nor \U$31885 ( \32138 , \32136 , \32137 );
and \U$31886 ( \32139 , \32128 , \32138 );
not \U$31887 ( \32140 , \4065 );
not \U$31888 ( \32141 , \14722 );
and \U$31889 ( \32142 , \32140 , \32141 );
and \U$31890 ( \32143 , \3303 , RIbe2a028_80);
nor \U$31891 ( \32144 , \32142 , \32143 );
and \U$31892 ( \32145 , \32144 , \9083 );
not \U$31893 ( \32146 , \32144 );
and \U$31894 ( \32147 , \32146 , \3516 );
nor \U$31895 ( \32148 , \32145 , \32147 );
or \U$31896 ( \32149 , \32139 , \32148 );
or \U$31897 ( \32150 , \32128 , \32138 );
nand \U$31898 ( \32151 , \32149 , \32150 );
not \U$31899 ( \32152 , \32151 );
not \U$31900 ( \32153 , RIbe2a3e8_88);
not \U$31901 ( \32154 , \1094 );
or \U$31902 ( \32155 , \32153 , \32154 );
nand \U$31903 ( \32156 , \4730 , RIbe2a370_87);
nand \U$31904 ( \32157 , \32155 , \32156 );
and \U$31905 ( \32158 , \32157 , \1309 );
not \U$31906 ( \32159 , \32157 );
and \U$31907 ( \32160 , \32159 , \4251 );
nor \U$31908 ( \32161 , \32158 , \32160 );
not \U$31909 ( \32162 , \32161 );
not \U$31910 ( \32163 , RIbe2a910_99);
not \U$31911 ( \32164 , \1143 );
or \U$31912 ( \32165 , \32163 , \32164 );
nand \U$31913 ( \32166 , \1147 , RIbe2b5b8_126);
nand \U$31914 ( \32167 , \32165 , \32166 );
not \U$31915 ( \32168 , \32167 );
not \U$31916 ( \32169 , \1153 );
and \U$31917 ( \32170 , \32168 , \32169 );
and \U$31918 ( \32171 , \32167 , \8327 );
nor \U$31919 ( \32172 , \32170 , \32171 );
not \U$31920 ( \32173 , \32172 );
not \U$31921 ( \32174 , \32173 );
or \U$31922 ( \32175 , \32162 , \32174 );
not \U$31923 ( \32176 , \32172 );
not \U$31924 ( \32177 , \32161 );
not \U$31925 ( \32178 , \32177 );
or \U$31926 ( \32179 , \32176 , \32178 );
and \U$31927 ( \32180 , \1113 , RIbe2a2f8_86);
and \U$31928 ( \32181 , \20664 , RIbe2acd0_107);
nor \U$31929 ( \32182 , \32180 , \32181 );
and \U$31930 ( \32183 , \32182 , \1131 );
not \U$31931 ( \32184 , \32182 );
and \U$31932 ( \32185 , \32184 , \1448 );
nor \U$31933 ( \32186 , \32183 , \32185 );
not \U$31934 ( \32187 , \32186 );
nand \U$31935 ( \32188 , \32179 , \32187 );
nand \U$31936 ( \32189 , \32175 , \32188 );
not \U$31937 ( \32190 , \32189 );
not \U$31938 ( \32191 , \32190 );
or \U$31939 ( \32192 , \32152 , \32191 );
not \U$31940 ( \32193 , \32151 );
nand \U$31941 ( \32194 , \32193 , \32189 );
nand \U$31942 ( \32195 , \32192 , \32194 );
and \U$31943 ( \32196 , \5973 , RIbe2a550_91);
and \U$31944 ( \32197 , \2000 , RIbe2a988_100);
nor \U$31945 ( \32198 , \32196 , \32197 );
and \U$31946 ( \32199 , \32198 , \1011 );
not \U$31947 ( \32200 , \32198 );
and \U$31948 ( \32201 , \32200 , \1813 );
nor \U$31949 ( \32202 , \32199 , \32201 );
not \U$31950 ( \32203 , \32202 );
not \U$31951 ( \32204 , \1761 );
not \U$31952 ( \32205 , \3774 );
not \U$31953 ( \32206 , \13156 );
and \U$31954 ( \32207 , \32205 , \32206 );
and \U$31955 ( \32208 , \546 , RIbe2a280_85);
nor \U$31956 ( \32209 , \32207 , \32208 );
not \U$31957 ( \32210 , \32209 );
or \U$31958 ( \32211 , \32204 , \32210 );
or \U$31959 ( \32212 , \32209 , \7123 );
nand \U$31960 ( \32213 , \32211 , \32212 );
not \U$31961 ( \32214 , \32213 );
not \U$31962 ( \32215 , \32214 );
and \U$31963 ( \32216 , \32203 , \32215 );
and \U$31964 ( \32217 , \32214 , \32202 );
and \U$31965 ( \32218 , \664 , RIbe2a190_83);
and \U$31966 ( \32219 , \740 , RIbe2a5c8_92);
nor \U$31967 ( \32220 , \32218 , \32219 );
not \U$31968 ( \32221 , \32220 );
not \U$31969 ( \32222 , \1621 );
and \U$31970 ( \32223 , \32221 , \32222 );
and \U$31971 ( \32224 , \672 , \32220 );
nor \U$31972 ( \32225 , \32223 , \32224 );
nor \U$31973 ( \32226 , \32217 , \32225 );
nor \U$31974 ( \32227 , \32216 , \32226 );
xor \U$31975 ( \32228 , \32195 , \32227 );
not \U$31976 ( \32229 , \32228 );
not \U$31977 ( \32230 , RIbe28228_16);
not \U$31978 ( \32231 , \10949 );
or \U$31979 ( \32232 , \32230 , \32231 );
nand \U$31980 ( \32233 , \8269 , RIbe281b0_15);
nand \U$31981 ( \32234 , \32232 , \32233 );
and \U$31982 ( \32235 , \32234 , \7984 );
not \U$31983 ( \32236 , \32234 );
and \U$31984 ( \32237 , \32236 , \9896 );
nor \U$31985 ( \32238 , \32235 , \32237 );
not \U$31986 ( \32239 , RIbe296c8_60);
not \U$31987 ( \32240 , \20530 );
or \U$31988 ( \32241 , \32239 , \32240 );
nand \U$31989 ( \32242 , \12212 , RIbe29650_59);
nand \U$31990 ( \32243 , \32241 , \32242 );
xor \U$31991 ( \32244 , \32243 , \13661 );
nand \U$31992 ( \32245 , \32238 , \32244 );
not \U$31993 ( \32246 , \8077 );
not \U$31994 ( \32247 , RIbe280c0_13);
not \U$31995 ( \32248 , \8276 );
or \U$31996 ( \32249 , \32247 , \32248 );
nand \U$31997 ( \32250 , \10919 , RIbe29830_63);
nand \U$31998 ( \32251 , \32249 , \32250 );
not \U$31999 ( \32252 , \32251 );
or \U$32000 ( \32253 , \32246 , \32252 );
or \U$32001 ( \32254 , \32251 , \25808 );
nand \U$32002 ( \32255 , \32253 , \32254 );
and \U$32003 ( \32256 , \32245 , \32255 );
nor \U$32004 ( \32257 , \32238 , \32244 );
nor \U$32005 ( \32258 , \32256 , \32257 );
not \U$32006 ( \32259 , RIbe27c10_3);
not \U$32007 ( \32260 , \12732 );
or \U$32008 ( \32261 , \32259 , \32260 );
nand \U$32009 ( \32262 , \13077 , RIbe28e58_42);
nand \U$32010 ( \32263 , \32261 , \32262 );
and \U$32011 ( \32264 , \32263 , \12746 );
not \U$32012 ( \32265 , \32263 );
and \U$32013 ( \32266 , \32265 , \13570 );
nor \U$32014 ( \32267 , \32264 , \32266 );
nand \U$32015 ( \32268 , \15249 , RIbe27b98_2);
and \U$32016 ( \32269 , \32268 , \12804 );
not \U$32017 ( \32270 , \32268 );
and \U$32018 ( \32271 , \32270 , \12893 );
nor \U$32019 ( \32272 , \32269 , \32271 );
and \U$32020 ( \32273 , \32267 , \32272 );
not \U$32021 ( \32274 , RIbe28de0_41);
not \U$32022 ( \32275 , \18608 );
or \U$32023 ( \32276 , \32274 , \32275 );
nand \U$32024 ( \32277 , \13012 , RIbe29920_65);
nand \U$32025 ( \32278 , \32276 , \32277 );
not \U$32026 ( \32279 , \32278 );
not \U$32027 ( \32280 , \12823 );
and \U$32028 ( \32281 , \32279 , \32280 );
and \U$32029 ( \32282 , \32278 , \12863 );
nor \U$32030 ( \32283 , \32281 , \32282 );
nor \U$32031 ( \32284 , \32273 , \32283 );
nor \U$32032 ( \32285 , \32267 , \32272 );
nor \U$32033 ( \32286 , \32284 , \32285 );
xor \U$32034 ( \32287 , \32258 , \32286 );
not \U$32035 ( \32288 , RIbe27d78_6);
not \U$32036 ( \32289 , \16383 );
or \U$32037 ( \32290 , \32288 , \32289 );
nand \U$32038 ( \32291 , \12711 , RIbe27d00_5);
nand \U$32039 ( \32292 , \32290 , \32291 );
and \U$32040 ( \32293 , \32292 , \12723 );
not \U$32041 ( \32294 , \32292 );
and \U$32042 ( \32295 , \32294 , \12716 );
nor \U$32043 ( \32296 , \32293 , \32295 );
not \U$32044 ( \32297 , \12752 );
not \U$32045 ( \32298 , \346 );
and \U$32046 ( \32299 , \32297 , \32298 );
and \U$32047 ( \32300 , \13738 , RIbe290b0_47);
nor \U$32048 ( \32301 , \32299 , \32300 );
and \U$32049 ( \32302 , \32301 , \12924 );
not \U$32050 ( \32303 , \32301 );
and \U$32051 ( \32304 , \32303 , \12927 );
nor \U$32052 ( \32305 , \32302 , \32304 );
not \U$32053 ( \32306 , \32305 );
nand \U$32054 ( \32307 , \32296 , \32306 );
not \U$32055 ( \32308 , RIbe29038_46);
not \U$32056 ( \32309 , \15205 );
or \U$32057 ( \32310 , \32308 , \32309 );
nand \U$32058 ( \32311 , \13669 , RIbe28fc0_45);
nand \U$32059 ( \32312 , \32310 , \32311 );
not \U$32060 ( \32313 , \32312 );
not \U$32061 ( \32314 , \12960 );
and \U$32062 ( \32315 , \32313 , \32314 );
and \U$32063 ( \32316 , \32312 , \17005 );
nor \U$32064 ( \32317 , \32315 , \32316 );
not \U$32065 ( \32318 , \32317 );
and \U$32066 ( \32319 , \32307 , \32318 );
nor \U$32067 ( \32320 , \32296 , \32306 );
nor \U$32068 ( \32321 , \32319 , \32320 );
xor \U$32069 ( \32322 , \32287 , \32321 );
not \U$32070 ( \32323 , \32322 );
or \U$32071 ( \32324 , \32229 , \32323 );
not \U$32072 ( \32325 , RIbe28f48_44);
not \U$32073 ( \32326 , \7880 );
or \U$32074 ( \32327 , \32325 , \32326 );
nand \U$32075 ( \32328 , \7438 , RIbe28ed0_43);
nand \U$32076 ( \32329 , \32327 , \32328 );
and \U$32077 ( \32330 , \32329 , \3471 );
not \U$32078 ( \32331 , \32329 );
and \U$32079 ( \32332 , \32331 , \3448 );
nor \U$32080 ( \32333 , \32330 , \32332 );
not \U$32081 ( \32334 , RIbe27fd0_11);
not \U$32082 ( \32335 , \5058 );
or \U$32083 ( \32336 , \32334 , \32335 );
nand \U$32084 ( \32337 , RIbe27f58_10, \4808 );
nand \U$32085 ( \32338 , \32336 , \32337 );
and \U$32086 ( \32339 , \32338 , \4603 );
not \U$32087 ( \32340 , \32338 );
and \U$32088 ( \32341 , \32340 , \4323 );
nor \U$32089 ( \32342 , \32339 , \32341 );
or \U$32090 ( \32343 , \32333 , \32342 );
not \U$32091 ( \32344 , RIbe27e68_8);
not \U$32092 ( \32345 , \21097 );
or \U$32093 ( \32346 , \32344 , \32345 );
not \U$32094 ( \32347 , \25899 );
nand \U$32095 ( \32348 , \32347 , \22378 );
nand \U$32096 ( \32349 , \32346 , \32348 );
and \U$32097 ( \32350 , \32349 , \4592 );
not \U$32098 ( \32351 , \32349 );
and \U$32099 ( \32352 , \32351 , \4586 );
nor \U$32100 ( \32353 , \32350 , \32352 );
not \U$32101 ( \32354 , \32353 );
nand \U$32102 ( \32355 , \32343 , \32354 );
nand \U$32103 ( \32356 , \32333 , \32342 );
nand \U$32104 ( \32357 , \32355 , \32356 );
not \U$32105 ( \32358 , RIbe28930_31);
not \U$32106 ( \32359 , \6980 );
or \U$32107 ( \32360 , \32358 , \32359 );
nand \U$32108 ( \32361 , \6985 , RIbe29560_57);
nand \U$32109 ( \32362 , \32360 , \32361 );
not \U$32110 ( \32363 , \32362 );
not \U$32111 ( \32364 , \7301 );
or \U$32112 ( \32365 , \32363 , \32364 );
or \U$32113 ( \32366 , \32362 , \7301 );
nand \U$32114 ( \32367 , \32365 , \32366 );
not \U$32115 ( \32368 , RIbe28a20_33);
not \U$32116 ( \32369 , \7954 );
or \U$32117 ( \32370 , \32368 , \32369 );
nand \U$32118 ( \32371 , \7958 , RIbe289a8_32);
nand \U$32119 ( \32372 , \32370 , \32371 );
and \U$32120 ( \32373 , \32372 , \7293 );
not \U$32121 ( \32374 , \32372 );
and \U$32122 ( \32375 , \32374 , \6572 );
nor \U$32123 ( \32376 , \32373 , \32375 );
xor \U$32124 ( \32377 , \32367 , \32376 );
not \U$32125 ( \32378 , RIbe28b88_36);
not \U$32126 ( \32379 , \7274 );
or \U$32127 ( \32380 , \32378 , \32379 );
nand \U$32128 ( \32381 , \7483 , RIbe29290_51);
nand \U$32129 ( \32382 , \32380 , \32381 );
and \U$32130 ( \32383 , \32382 , \6582 );
not \U$32131 ( \32384 , \32382 );
and \U$32132 ( \32385 , \32384 , \6583 );
nor \U$32133 ( \32386 , \32383 , \32385 );
and \U$32134 ( \32387 , \32377 , \32386 );
and \U$32135 ( \32388 , \32367 , \32376 );
or \U$32136 ( \32389 , \32387 , \32388 );
xor \U$32137 ( \32390 , \32357 , \32389 );
not \U$32138 ( \32391 , \6547 );
and \U$32139 ( \32392 , \6880 , RIbe28390_19);
and \U$32140 ( \32393 , \6539 , RIbe28b10_35);
nor \U$32141 ( \32394 , \32392 , \32393 );
not \U$32142 ( \32395 , \32394 );
or \U$32143 ( \32396 , \32391 , \32395 );
or \U$32144 ( \32397 , \7935 , \32394 );
nand \U$32145 ( \32398 , \32396 , \32397 );
not \U$32146 ( \32399 , RIbe28480_21);
not \U$32147 ( \32400 , \8231 );
or \U$32148 ( \32401 , \32399 , \32400 );
nand \U$32149 ( \32402 , \6859 , RIbe28408_20);
nand \U$32150 ( \32403 , \32401 , \32402 );
and \U$32151 ( \32404 , \32403 , \5741 );
not \U$32152 ( \32405 , \32403 );
and \U$32153 ( \32406 , \32405 , \6624 );
nor \U$32154 ( \32407 , \32404 , \32406 );
xor \U$32155 ( \32408 , \32398 , \32407 );
not \U$32156 ( \32409 , RIbe285e8_24);
not \U$32157 ( \32410 , \6630 );
or \U$32158 ( \32411 , \32409 , \32410 );
nand \U$32159 ( \32412 , \14239 , RIbe287c8_28);
nand \U$32160 ( \32413 , \32411 , \32412 );
and \U$32161 ( \32414 , \32413 , \6907 );
not \U$32162 ( \32415 , \32413 );
and \U$32163 ( \32416 , \32415 , \6641 );
nor \U$32164 ( \32417 , \32414 , \32416 );
and \U$32165 ( \32418 , \32408 , \32417 );
and \U$32166 ( \32419 , \32398 , \32407 );
or \U$32167 ( \32420 , \32418 , \32419 );
and \U$32168 ( \32421 , \32390 , \32420 );
not \U$32169 ( \32422 , \32390 );
not \U$32170 ( \32423 , \32420 );
and \U$32171 ( \32424 , \32422 , \32423 );
nor \U$32172 ( \32425 , \32421 , \32424 );
nand \U$32173 ( \32426 , \32324 , \32425 );
not \U$32174 ( \32427 , \32322 );
not \U$32175 ( \32428 , \32228 );
nand \U$32176 ( \32429 , \32427 , \32428 );
nand \U$32177 ( \32430 , \32426 , \32429 );
not \U$32178 ( \32431 , \32430 );
not \U$32179 ( \32432 , \32431 );
and \U$32180 ( \32433 , \3160 , RIbe2afa0_113);
and \U$32181 ( \32434 , \329 , RIbe2af28_112);
nor \U$32182 ( \32435 , \32433 , \32434 );
and \U$32183 ( \32436 , \32435 , \1379 );
not \U$32184 ( \32437 , \32435 );
and \U$32185 ( \32438 , \32437 , \338 );
nor \U$32186 ( \32439 , \32436 , \32438 );
not \U$32187 ( \32440 , RIbe2b018_114);
not \U$32188 ( \32441 , \325 );
or \U$32189 ( \32442 , \32440 , \32441 );
nand \U$32190 ( \32443 , \330 , RIbe2afa0_113);
nand \U$32191 ( \32444 , \32442 , \32443 );
and \U$32192 ( \32445 , \32444 , \1379 );
not \U$32193 ( \32446 , \32444 );
and \U$32194 ( \32447 , \32446 , \338 );
nor \U$32195 ( \32448 , \32445 , \32447 );
nand \U$32196 ( \32449 , RIbe29380_53, RIbe2b630_127);
nand \U$32197 ( \32450 , \32448 , \32449 );
xor \U$32198 ( \32451 , \32439 , \32450 );
not \U$32199 ( \32452 , RIbe2b180_117);
buf \U$32200 ( \32453 , \278 );
nor \U$32201 ( \32454 , \1681 , \32453 );
not \U$32202 ( \32455 , \32454 );
or \U$32203 ( \32456 , \32452 , \32455 );
not \U$32204 ( \32457 , \13109 );
nand \U$32205 ( \32458 , \32457 , \1681 );
nand \U$32206 ( \32459 , \32456 , \32458 );
and \U$32207 ( \32460 , \32459 , \293 );
not \U$32208 ( \32461 , \32459 );
and \U$32209 ( \32462 , \32461 , \300 );
nor \U$32210 ( \32463 , \32460 , \32462 );
not \U$32211 ( \32464 , RIbe2b108_116);
not \U$32212 ( \32465 , \1773 );
or \U$32213 ( \32466 , \32464 , \32465 );
nand \U$32214 ( \32467 , \429 , RIbe2b090_115);
nand \U$32215 ( \32468 , \32466 , \32467 );
and \U$32216 ( \32469 , \32468 , \306 );
not \U$32217 ( \32470 , \32468 );
and \U$32218 ( \32471 , \32470 , \312 );
nor \U$32219 ( \32472 , \32469 , \32471 );
xor \U$32220 ( \32473 , \32463 , \32472 );
and \U$32221 ( \32474 , \1659 , RIbe2af28_112);
and \U$32222 ( \32475 , \6325 , RIbe2b1f8_118);
nor \U$32223 ( \32476 , \32474 , \32475 );
and \U$32224 ( \32477 , \32476 , \1362 );
not \U$32225 ( \32478 , \32476 );
and \U$32226 ( \32479 , \32478 , \269 );
nor \U$32227 ( \32480 , \32477 , \32479 );
and \U$32228 ( \32481 , \32473 , \32480 );
and \U$32229 ( \32482 , \32463 , \32472 );
or \U$32230 ( \32483 , \32481 , \32482 );
xor \U$32231 ( \32484 , \32451 , \32483 );
not \U$32232 ( \32485 , \32484 );
not \U$32233 ( \32486 , RIbe27f58_10);
not \U$32234 ( \32487 , \4317 );
or \U$32235 ( \32488 , \32486 , \32487 );
nand \U$32236 ( \32489 , RIbe27e68_8, \7858 );
nand \U$32237 ( \32490 , \32488 , \32489 );
and \U$32238 ( \32491 , \32490 , \4326 );
not \U$32239 ( \32492 , \32490 );
and \U$32240 ( \32493 , \32492 , \7865 );
nor \U$32241 ( \32494 , \32491 , \32493 );
not \U$32242 ( \32495 , RIbe28660_25);
not \U$32243 ( \32496 , \15894 );
or \U$32244 ( \32497 , \32495 , \32496 );
nand \U$32245 ( \32498 , \5731 , RIbe285e8_24);
nand \U$32246 ( \32499 , \32497 , \32498 );
and \U$32247 ( \32500 , \32499 , \4586 );
not \U$32248 ( \32501 , \32499 );
and \U$32249 ( \32502 , \32501 , \20465 );
nor \U$32250 ( \32503 , \32500 , \32502 );
xor \U$32251 ( \32504 , \32494 , \32503 );
not \U$32252 ( \32505 , RIbe28ed0_43);
not \U$32253 ( \32506 , \6783 );
or \U$32254 ( \32507 , \32505 , \32506 );
nand \U$32255 ( \32508 , \4027 , RIbe27fd0_11);
nand \U$32256 ( \32509 , \32507 , \32508 );
and \U$32257 ( \32510 , \32509 , \3471 );
not \U$32258 ( \32511 , \32509 );
and \U$32259 ( \32512 , \32511 , \3448 );
nor \U$32260 ( \32513 , \32510 , \32512 );
xor \U$32261 ( \32514 , \32504 , \32513 );
not \U$32262 ( \32515 , \32514 );
not \U$32263 ( \32516 , RIbe2acd0_107);
not \U$32264 ( \32517 , \23509 );
or \U$32265 ( \32518 , \32516 , \32517 );
nand \U$32266 ( \32519 , \1117 , RIbe2a028_80);
nand \U$32267 ( \32520 , \32518 , \32519 );
and \U$32268 ( \32521 , \32520 , \1132 );
not \U$32269 ( \32522 , \32520 );
and \U$32270 ( \32523 , \32522 , \1125 );
nor \U$32271 ( \32524 , \32521 , \32523 );
not \U$32272 ( \32525 , RIbe2a370_87);
not \U$32273 ( \32526 , \8868 );
or \U$32274 ( \32527 , \32525 , \32526 );
nand \U$32275 ( \32528 , RIbe2a2f8_86, \1098 );
nand \U$32276 ( \32529 , \32527 , \32528 );
and \U$32277 ( \32530 , \32529 , \1082 );
not \U$32278 ( \32531 , \32529 );
and \U$32279 ( \32532 , \32531 , \1309 );
nor \U$32280 ( \32533 , \32530 , \32532 );
and \U$32281 ( \32534 , \32524 , \32533 );
not \U$32282 ( \32535 , \32524 );
not \U$32283 ( \32536 , \32533 );
and \U$32284 ( \32537 , \32535 , \32536 );
nor \U$32285 ( \32538 , \32534 , \32537 );
not \U$32286 ( \32539 , RIbe2b5b8_126);
not \U$32287 ( \32540 , \1143 );
or \U$32288 ( \32541 , \32539 , \32540 );
nand \U$32289 ( \32542 , \1147 , RIbe2a3e8_88);
nand \U$32290 ( \32543 , \32541 , \32542 );
and \U$32291 ( \32544 , \32543 , \3993 );
not \U$32292 ( \32545 , \32543 );
and \U$32293 ( \32546 , \32545 , \1153 );
nor \U$32294 ( \32547 , \32544 , \32546 );
xor \U$32295 ( \32548 , \32538 , \32547 );
not \U$32296 ( \32549 , \32548 );
or \U$32297 ( \32550 , \32515 , \32549 );
or \U$32298 ( \32551 , \32514 , \32548 );
nand \U$32299 ( \32552 , \32550 , \32551 );
and \U$32300 ( \32553 , \8833 , RIbe29fb0_79);
and \U$32301 ( \32554 , \2384 , RIbe29e48_76);
nor \U$32302 ( \32555 , \32553 , \32554 );
and \U$32303 ( \32556 , \32555 , \1076 );
not \U$32304 ( \32557 , \32555 );
and \U$32305 ( \32558 , \32557 , \9083 );
nor \U$32306 ( \32559 , \32556 , \32558 );
not \U$32307 ( \32560 , RIbe29dd0_75);
not \U$32308 ( \32561 , \2898 );
or \U$32309 ( \32562 , \32560 , \32561 );
not \U$32310 ( \32563 , \9801 );
nand \U$32311 ( \32564 , \32563 , \3267 );
nand \U$32312 ( \32565 , \32562 , \32564 );
and \U$32313 ( \32566 , \32565 , \25477 );
not \U$32314 ( \32567 , \32565 );
and \U$32315 ( \32568 , \32567 , \2379 );
nor \U$32316 ( \32569 , \32566 , \32568 );
xor \U$32317 ( \32570 , \32559 , \32569 );
not \U$32318 ( \32571 , RIbe29bf0_71);
not \U$32319 ( \32572 , \3452 );
or \U$32320 ( \32573 , \32571 , \32572 );
nand \U$32321 ( \32574 , \3689 , RIbe28f48_44);
nand \U$32322 ( \32575 , \32573 , \32574 );
and \U$32323 ( \32576 , \32575 , \3290 );
not \U$32324 ( \32577 , \32575 );
and \U$32325 ( \32578 , \32577 , \3461 );
nor \U$32326 ( \32579 , \32576 , \32578 );
xor \U$32327 ( \32580 , \32570 , \32579 );
not \U$32328 ( \32581 , \32580 );
and \U$32329 ( \32582 , \32552 , \32581 );
not \U$32330 ( \32583 , \32552 );
and \U$32331 ( \32584 , \32583 , \32580 );
nor \U$32332 ( \32585 , \32582 , \32584 );
and \U$32333 ( \32586 , \32485 , \32585 );
and \U$32334 ( \32587 , RIbe29380_53, RIbe2b018_114);
not \U$32335 ( \32588 , RIbe2a5c8_92);
not \U$32336 ( \32589 , \1743 );
not \U$32337 ( \32590 , \32589 );
or \U$32338 ( \32591 , \32588 , \32590 );
not \U$32339 ( \32592 , \21491 );
nand \U$32340 ( \32593 , \32592 , \1179 );
nand \U$32341 ( \32594 , \32591 , \32593 );
and \U$32342 ( \32595 , \32594 , \672 );
not \U$32343 ( \32596 , \32594 );
and \U$32344 ( \32597 , \32596 , \564 );
nor \U$32345 ( \32598 , \32595 , \32597 );
and \U$32346 ( \32599 , \546 , RIbe2a208_84);
not \U$32347 ( \32600 , \552 );
nor \U$32348 ( \32601 , \32600 , \14285 );
nor \U$32349 ( \32602 , \32599 , \32601 );
and \U$32350 ( \32603 , \32602 , \424 );
not \U$32351 ( \32604 , \32602 );
and \U$32352 ( \32605 , \32604 , \425 );
nor \U$32353 ( \32606 , \32603 , \32605 );
xor \U$32354 ( \32607 , \32598 , \32606 );
and \U$32355 ( \32608 , \4858 , RIbe2a988_100);
and \U$32356 ( \32609 , \1203 , RIbe2a910_99);
nor \U$32357 ( \32610 , \32608 , \32609 );
and \U$32358 ( \32611 , \32610 , \1608 );
not \U$32359 ( \32612 , \32610 );
and \U$32360 ( \32613 , \32612 , \1011 );
nor \U$32361 ( \32614 , \32611 , \32613 );
xor \U$32362 ( \32615 , \32607 , \32614 );
xor \U$32363 ( \32616 , \32587 , \32615 );
not \U$32364 ( \32617 , RIbe2b270_119);
not \U$32365 ( \32618 , \1252 );
or \U$32366 ( \32619 , \32617 , \32618 );
nand \U$32367 ( \32620 , \1682 , RIbe2b108_116);
nand \U$32368 ( \32621 , \32619 , \32620 );
and \U$32369 ( \32622 , \32621 , \293 );
not \U$32370 ( \32623 , \32621 );
and \U$32371 ( \32624 , \32623 , \300 );
nor \U$32372 ( \32625 , \32622 , \32624 );
not \U$32373 ( \32626 , RIbe2b090_115);
not \U$32374 ( \32627 , \1223 );
or \U$32375 ( \32628 , \32626 , \32627 );
nand \U$32376 ( \32629 , \429 , RIbe2a280_85);
nand \U$32377 ( \32630 , \32628 , \32629 );
and \U$32378 ( \32631 , \32630 , \313 );
not \U$32379 ( \32632 , \32630 );
and \U$32380 ( \32633 , \32632 , \306 );
nor \U$32381 ( \32634 , \32631 , \32633 );
xor \U$32382 ( \32635 , \32625 , \32634 );
not \U$32383 ( \32636 , RIbe2b1f8_118);
not \U$32384 ( \32637 , \260 );
or \U$32385 ( \32638 , \32636 , \32637 );
not \U$32386 ( \32639 , \14248 );
nand \U$32387 ( \32640 , \32639 , \263 );
nand \U$32388 ( \32641 , \32638 , \32640 );
and \U$32389 ( \32642 , \32641 , \1663 );
not \U$32390 ( \32643 , \32641 );
and \U$32391 ( \32644 , \32643 , \6058 );
nor \U$32392 ( \32645 , \32642 , \32644 );
xnor \U$32393 ( \32646 , \32635 , \32645 );
xnor \U$32394 ( \32647 , \32616 , \32646 );
nor \U$32395 ( \32648 , \32586 , \32647 );
nor \U$32396 ( \32649 , \32585 , \32485 );
nor \U$32397 ( \32650 , \32648 , \32649 );
not \U$32398 ( \32651 , \32650 );
or \U$32399 ( \32652 , \32432 , \32651 );
not \U$32400 ( \32653 , RIbe29920_65);
not \U$32401 ( \32654 , \13010 );
or \U$32402 ( \32655 , \32653 , \32654 );
nand \U$32403 ( \32656 , \12835 , RIbe27b98_2);
nand \U$32404 ( \32657 , \32655 , \32656 );
and \U$32405 ( \32658 , \32657 , \12866 );
not \U$32406 ( \32659 , \32657 );
and \U$32407 ( \32660 , \32659 , \12863 );
nor \U$32408 ( \32661 , \32658 , \32660 );
xor \U$32409 ( \32662 , \12998 , \32661 );
not \U$32410 ( \32663 , \12746 );
not \U$32411 ( \32664 , RIbe28e58_42);
not \U$32412 ( \32665 , \12732 );
or \U$32413 ( \32666 , \32664 , \32665 );
nand \U$32414 ( \32667 , \14074 , RIbe28de0_41);
nand \U$32415 ( \32668 , \32666 , \32667 );
not \U$32416 ( \32669 , \32668 );
or \U$32417 ( \32670 , \32663 , \32669 );
or \U$32418 ( \32671 , \32668 , \12746 );
nand \U$32419 ( \32672 , \32670 , \32671 );
and \U$32420 ( \32673 , \32662 , \32672 );
and \U$32421 ( \32674 , \12998 , \32661 );
or \U$32422 ( \32675 , \32673 , \32674 );
and \U$32423 ( \32676 , \8278 , RIbe29830_63);
and \U$32424 ( \32677 , \13038 , RIbe296c8_60);
nor \U$32425 ( \32678 , \32676 , \32677 );
and \U$32426 ( \32679 , \32678 , \25808 );
not \U$32427 ( \32680 , \32678 );
and \U$32428 ( \32681 , \32680 , \16994 );
nor \U$32429 ( \32682 , \32679 , \32681 );
not \U$32430 ( \32683 , RIbe281b0_15);
not \U$32431 ( \32684 , \10949 );
or \U$32432 ( \32685 , \32683 , \32684 );
nand \U$32433 ( \32686 , \7981 , RIbe280c0_13);
nand \U$32434 ( \32687 , \32685 , \32686 );
and \U$32435 ( \32688 , \32687 , \7985 );
not \U$32436 ( \32689 , \32687 );
and \U$32437 ( \32690 , \32689 , \7989 );
nor \U$32438 ( \32691 , \32688 , \32690 );
xor \U$32439 ( \32692 , \32682 , \32691 );
not \U$32440 ( \32693 , RIbe29650_59);
not \U$32441 ( \32694 , \10936 );
or \U$32442 ( \32695 , \32693 , \32694 );
nand \U$32443 ( \32696 , \14511 , RIbe29038_46);
nand \U$32444 ( \32697 , \32695 , \32696 );
and \U$32445 ( \32698 , \32697 , \17297 );
not \U$32446 ( \32699 , \32697 );
and \U$32447 ( \32700 , \32699 , \10940 );
nor \U$32448 ( \32701 , \32698 , \32700 );
and \U$32449 ( \32702 , \32692 , \32701 );
and \U$32450 ( \32703 , \32682 , \32691 );
or \U$32451 ( \32704 , \32702 , \32703 );
xor \U$32452 ( \32705 , \32675 , \32704 );
not \U$32453 ( \32706 , \12753 );
not \U$32454 ( \32707 , \255 );
and \U$32455 ( \32708 , \32706 , \32707 );
and \U$32456 ( \32709 , \12765 , RIbe29a88_68);
nor \U$32457 ( \32710 , \32708 , \32709 );
and \U$32458 ( \32711 , \32710 , \12924 );
not \U$32459 ( \32712 , \32710 );
and \U$32460 ( \32713 , \32712 , \12774 );
nor \U$32461 ( \32714 , \32711 , \32713 );
not \U$32462 ( \32715 , \12195 );
and \U$32463 ( \32716 , \12942 , RIbe28fc0_45);
and \U$32464 ( \32717 , \15628 , RIbe290b0_47);
nor \U$32465 ( \32718 , \32716 , \32717 );
not \U$32466 ( \32719 , \32718 );
or \U$32467 ( \32720 , \32715 , \32719 );
or \U$32468 ( \32721 , \32718 , \12195 );
nand \U$32469 ( \32722 , \32720 , \32721 );
xor \U$32470 ( \32723 , \32714 , \32722 );
not \U$32471 ( \32724 , RIbe27d00_5);
not \U$32472 ( \32725 , \14523 );
or \U$32473 ( \32726 , \32724 , \32725 );
nand \U$32474 ( \32727 , \13728 , RIbe27c10_3);
nand \U$32475 ( \32728 , \32726 , \32727 );
and \U$32476 ( \32729 , \32728 , \12716 );
not \U$32477 ( \32730 , \32728 );
and \U$32478 ( \32731 , \32730 , \12723 );
nor \U$32479 ( \32732 , \32729 , \32731 );
and \U$32480 ( \32733 , \32723 , \32732 );
and \U$32481 ( \32734 , \32714 , \32722 );
or \U$32482 ( \32735 , \32733 , \32734 );
xor \U$32483 ( \32736 , \32705 , \32735 );
xor \U$32484 ( \32737 , \32494 , \32503 );
and \U$32485 ( \32738 , \32737 , \32513 );
and \U$32486 ( \32739 , \32494 , \32503 );
or \U$32487 ( \32740 , \32738 , \32739 );
not \U$32488 ( \32741 , RIbe29560_57);
not \U$32489 ( \32742 , \6980 );
or \U$32490 ( \32743 , \32741 , \32742 );
not \U$32491 ( \32744 , \3952 );
nand \U$32492 ( \32745 , \32744 , \10898 );
nand \U$32493 ( \32746 , \32743 , \32745 );
and \U$32494 ( \32747 , \32746 , \7304 );
not \U$32495 ( \32748 , \32746 );
and \U$32496 ( \32749 , \32748 , \6992 );
nor \U$32497 ( \32750 , \32747 , \32749 );
not \U$32498 ( \32751 , RIbe289a8_32);
not \U$32499 ( \32752 , \8199 );
or \U$32500 ( \32753 , \32751 , \32752 );
nand \U$32501 ( \32754 , \8202 , RIbe28930_31);
nand \U$32502 ( \32755 , \32753 , \32754 );
and \U$32503 ( \32756 , \32755 , \7293 );
not \U$32504 ( \32757 , \32755 );
and \U$32505 ( \32758 , \32757 , \6572 );
nor \U$32506 ( \32759 , \32756 , \32758 );
xor \U$32507 ( \32760 , \32750 , \32759 );
not \U$32508 ( \32761 , RIbe29290_51);
not \U$32509 ( \32762 , \7274 );
or \U$32510 ( \32763 , \32761 , \32762 );
nand \U$32511 ( \32764 , \7483 , RIbe28a20_33);
nand \U$32512 ( \32765 , \32763 , \32764 );
and \U$32513 ( \32766 , \32765 , \6582 );
not \U$32514 ( \32767 , \32765 );
and \U$32515 ( \32768 , \32767 , \7646 );
nor \U$32516 ( \32769 , \32766 , \32768 );
and \U$32517 ( \32770 , \32760 , \32769 );
and \U$32518 ( \32771 , \32750 , \32759 );
or \U$32519 ( \32772 , \32770 , \32771 );
xor \U$32520 ( \32773 , \32740 , \32772 );
not \U$32521 ( \32774 , RIbe28b10_35);
not \U$32522 ( \32775 , \6880 );
or \U$32523 ( \32776 , \32774 , \32775 );
nand \U$32524 ( \32777 , \6884 , RIbe28b88_36);
nand \U$32525 ( \32778 , \32776 , \32777 );
and \U$32526 ( \32779 , \32778 , \6552 );
not \U$32527 ( \32780 , \32778 );
and \U$32528 ( \32781 , \32780 , \6891 );
nor \U$32529 ( \32782 , \32779 , \32781 );
not \U$32530 ( \32783 , RIbe28408_20);
not \U$32531 ( \32784 , \6139 );
or \U$32532 ( \32785 , \32783 , \32784 );
nand \U$32533 ( \32786 , \8235 , RIbe28390_19);
nand \U$32534 ( \32787 , \32785 , \32786 );
and \U$32535 ( \32788 , \32787 , \10969 );
not \U$32536 ( \32789 , \32787 );
and \U$32537 ( \32790 , \32789 , \10972 );
nor \U$32538 ( \32791 , \32788 , \32790 );
xor \U$32539 ( \32792 , \32782 , \32791 );
not \U$32540 ( \32793 , RIbe287c8_28);
not \U$32541 ( \32794 , \5455 );
or \U$32542 ( \32795 , \32793 , \32794 );
nand \U$32543 ( \32796 , \10269 , RIbe28480_21);
nand \U$32544 ( \32797 , \32795 , \32796 );
and \U$32545 ( \32798 , \32797 , \6907 );
not \U$32546 ( \32799 , \32797 );
and \U$32547 ( \32800 , \32799 , \5457 );
nor \U$32548 ( \32801 , \32798 , \32800 );
and \U$32549 ( \32802 , \32792 , \32801 );
and \U$32550 ( \32803 , \32782 , \32791 );
or \U$32551 ( \32804 , \32802 , \32803 );
xor \U$32552 ( \32805 , \32773 , \32804 );
xor \U$32553 ( \32806 , \32736 , \32805 );
xor \U$32554 ( \32807 , \32598 , \32606 );
and \U$32555 ( \32808 , \32807 , \32614 );
and \U$32556 ( \32809 , \32598 , \32606 );
or \U$32557 ( \32810 , \32808 , \32809 );
not \U$32558 ( \32811 , \32536 );
not \U$32559 ( \32812 , \32547 );
or \U$32560 ( \32813 , \32811 , \32812 );
or \U$32561 ( \32814 , \32547 , \32536 );
nand \U$32562 ( \32815 , \32814 , \32524 );
nand \U$32563 ( \32816 , \32813 , \32815 );
xor \U$32564 ( \32817 , \32810 , \32816 );
xor \U$32565 ( \32818 , \32559 , \32569 );
and \U$32566 ( \32819 , \32818 , \32579 );
and \U$32567 ( \32820 , \32559 , \32569 );
or \U$32568 ( \32821 , \32819 , \32820 );
xor \U$32569 ( \32822 , \32817 , \32821 );
xor \U$32570 ( \32823 , \32806 , \32822 );
nand \U$32571 ( \32824 , \32652 , \32823 );
not \U$32572 ( \32825 , \32431 );
not \U$32573 ( \32826 , \32650 );
nand \U$32574 ( \32827 , \32825 , \32826 );
nand \U$32575 ( \32828 , \32824 , \32827 );
not \U$32576 ( \32829 , RIbe2a988_100);
not \U$32577 ( \32830 , \4257 );
or \U$32578 ( \32831 , \32829 , \32830 );
nand \U$32579 ( \32832 , \1147 , RIbe2a910_99);
nand \U$32580 ( \32833 , \32831 , \32832 );
and \U$32581 ( \32834 , \32833 , \3993 );
not \U$32582 ( \32835 , \32833 );
and \U$32583 ( \32836 , \32835 , \1157 );
nor \U$32584 ( \32837 , \32834 , \32836 );
not \U$32585 ( \32838 , \8173 );
not \U$32586 ( \32839 , \14285 );
and \U$32587 ( \32840 , \32838 , \32839 );
and \U$32588 ( \32841 , \664 , RIbe2a208_84);
nor \U$32589 ( \32842 , \32840 , \32841 );
and \U$32590 ( \32843 , \32842 , \564 );
not \U$32591 ( \32844 , \32842 );
and \U$32592 ( \32845 , \32844 , \3959 );
nor \U$32593 ( \32846 , \32843 , \32845 );
xor \U$32594 ( \32847 , \32837 , \32846 );
and \U$32595 ( \32848 , \1807 , RIbe2a5c8_92);
and \U$32596 ( \32849 , \1203 , RIbe2a550_91);
nor \U$32597 ( \32850 , \32848 , \32849 );
and \U$32598 ( \32851 , \32850 , \1608 );
not \U$32599 ( \32852 , \32850 );
and \U$32600 ( \32853 , \32852 , \1011 );
nor \U$32601 ( \32854 , \32851 , \32853 );
and \U$32602 ( \32855 , \32847 , \32854 );
and \U$32603 ( \32856 , \32837 , \32846 );
or \U$32604 ( \32857 , \32855 , \32856 );
and \U$32605 ( \32858 , \27601 , RIbe2a370_87);
and \U$32606 ( \32859 , \5467 , RIbe2a2f8_86);
nor \U$32607 ( \32860 , \32858 , \32859 );
and \U$32608 ( \32861 , \32860 , \2563 );
not \U$32609 ( \32862 , \32860 );
and \U$32610 ( \32863 , \32862 , \1131 );
nor \U$32611 ( \32864 , \32861 , \32863 );
not \U$32612 ( \32865 , RIbe2b5b8_126);
not \U$32613 ( \32866 , \1094 );
or \U$32614 ( \32867 , \32865 , \32866 );
nand \U$32615 ( \32868 , \4730 , RIbe2a3e8_88);
nand \U$32616 ( \32869 , \32867 , \32868 );
and \U$32617 ( \32870 , \32869 , \1309 );
not \U$32618 ( \32871 , \32869 );
and \U$32619 ( \32872 , \32871 , \2418 );
nor \U$32620 ( \32873 , \32870 , \32872 );
or \U$32621 ( \32874 , \32864 , \32873 );
not \U$32622 ( \32875 , \2889 );
not \U$32623 ( \32876 , \14374 );
and \U$32624 ( \32877 , \32875 , \32876 );
and \U$32625 ( \32878 , \4295 , RIbe2acd0_107);
nor \U$32626 ( \32879 , \32877 , \32878 );
and \U$32627 ( \32880 , \32879 , \1277 );
not \U$32628 ( \32881 , \32879 );
and \U$32629 ( \32882 , \32881 , \1076 );
nor \U$32630 ( \32883 , \32880 , \32882 );
not \U$32631 ( \32884 , \32883 );
nand \U$32632 ( \32885 , \32874 , \32884 );
nand \U$32633 ( \32886 , \32864 , \32873 );
nand \U$32634 ( \32887 , \32885 , \32886 );
xor \U$32635 ( \32888 , \32857 , \32887 );
not \U$32636 ( \32889 , \2576 );
not \U$32637 ( \32890 , RIbe29fb0_79);
not \U$32638 ( \32891 , \2898 );
or \U$32639 ( \32892 , \32890 , \32891 );
nand \U$32640 ( \32893 , \3267 , RIbe29e48_76);
nand \U$32641 ( \32894 , \32892 , \32893 );
not \U$32642 ( \32895 , \32894 );
or \U$32643 ( \32896 , \32889 , \32895 );
or \U$32644 ( \32897 , \32894 , \2379 );
nand \U$32645 ( \32898 , \32896 , \32897 );
not \U$32646 ( \32899 , RIbe29dd0_75);
not \U$32647 ( \32900 , \3284 );
or \U$32648 ( \32901 , \32899 , \32900 );
nand \U$32649 ( \32902 , \3689 , RIbe29c68_72);
nand \U$32650 ( \32903 , \32901 , \32902 );
and \U$32651 ( \32904 , \32903 , \3290 );
not \U$32652 ( \32905 , \32903 );
and \U$32653 ( \32906 , \32905 , \3461 );
nor \U$32654 ( \32907 , \32904 , \32906 );
xor \U$32655 ( \32908 , \32898 , \32907 );
not \U$32656 ( \32909 , RIbe29bf0_71);
not \U$32657 ( \32910 , \5094 );
or \U$32658 ( \32911 , \32909 , \32910 );
nand \U$32659 ( \32912 , \4333 , RIbe28f48_44);
nand \U$32660 ( \32913 , \32911 , \32912 );
and \U$32661 ( \32914 , \32913 , \3471 );
not \U$32662 ( \32915 , \32913 );
and \U$32663 ( \32916 , \32915 , \3698 );
nor \U$32664 ( \32917 , \32914 , \32916 );
and \U$32665 ( \32918 , \32908 , \32917 );
and \U$32666 ( \32919 , \32898 , \32907 );
or \U$32667 ( \32920 , \32918 , \32919 );
and \U$32668 ( \32921 , \32888 , \32920 );
and \U$32669 ( \32922 , \32857 , \32887 );
or \U$32670 ( \32923 , \32921 , \32922 );
not \U$32671 ( \32924 , \32923 );
not \U$32672 ( \32925 , \32924 );
not \U$32673 ( \32926 , RIbe28b10_35);
not \U$32674 ( \32927 , \7941 );
or \U$32675 ( \32928 , \32926 , \32927 );
nand \U$32676 ( \32929 , \13436 , RIbe28b88_36);
nand \U$32677 ( \32930 , \32928 , \32929 );
and \U$32678 ( \32931 , \32930 , \6582 );
not \U$32679 ( \32932 , \32930 );
and \U$32680 ( \32933 , \32932 , \7271 );
nor \U$32681 ( \32934 , \32931 , \32933 );
not \U$32682 ( \32935 , RIbe287c8_28);
not \U$32683 ( \32936 , \8231 );
or \U$32684 ( \32937 , \32935 , \32936 );
nand \U$32685 ( \32938 , \7528 , RIbe28480_21);
nand \U$32686 ( \32939 , \32937 , \32938 );
and \U$32687 ( \32940 , \32939 , \6144 );
not \U$32688 ( \32941 , \32939 );
and \U$32689 ( \32942 , \32941 , \6141 );
nor \U$32690 ( \32943 , \32940 , \32942 );
or \U$32691 ( \32944 , \32934 , \32943 );
not \U$32692 ( \32945 , RIbe28408_20);
not \U$32693 ( \32946 , \6536 );
or \U$32694 ( \32947 , \32945 , \32946 );
nand \U$32695 ( \32948 , \7076 , RIbe28390_19);
nand \U$32696 ( \32949 , \32947 , \32948 );
not \U$32697 ( \32950 , \32949 );
not \U$32698 ( \32951 , \9933 );
and \U$32699 ( \32952 , \32950 , \32951 );
and \U$32700 ( \32953 , \32949 , \6891 );
nor \U$32701 ( \32954 , \32952 , \32953 );
not \U$32702 ( \32955 , \32954 );
nand \U$32703 ( \32956 , \32944 , \32955 );
nand \U$32704 ( \32957 , \32934 , \32943 );
nand \U$32705 ( \32958 , \32956 , \32957 );
not \U$32706 ( \32959 , \32958 );
not \U$32707 ( \32960 , RIbe28ed0_43);
not \U$32708 ( \32961 , \4804 );
or \U$32709 ( \32962 , \32960 , \32961 );
nand \U$32710 ( \32963 , \7858 , RIbe27fd0_11);
nand \U$32711 ( \32964 , \32962 , \32963 );
and \U$32712 ( \32965 , \32964 , \4326 );
not \U$32713 ( \32966 , \32964 );
and \U$32714 ( \32967 , \32966 , \4323 );
nor \U$32715 ( \32968 , \32965 , \32967 );
not \U$32716 ( \32969 , \32968 );
not \U$32717 ( \32970 , RIbe27f58_10);
not \U$32718 ( \32971 , \15894 );
or \U$32719 ( \32972 , \32970 , \32971 );
nand \U$32720 ( \32973 , \5731 , RIbe27e68_8);
nand \U$32721 ( \32974 , \32972 , \32973 );
and \U$32722 ( \32975 , \32974 , \4586 );
not \U$32723 ( \32976 , \32974 );
and \U$32724 ( \32977 , \32976 , \4946 );
nor \U$32725 ( \32978 , \32975 , \32977 );
not \U$32726 ( \32979 , \32978 );
or \U$32727 ( \32980 , \32969 , \32979 );
or \U$32728 ( \32981 , \32978 , \32968 );
not \U$32729 ( \32982 , RIbe28660_25);
not \U$32730 ( \32983 , \6630 );
or \U$32731 ( \32984 , \32982 , \32983 );
nand \U$32732 ( \32985 , \10269 , RIbe285e8_24);
nand \U$32733 ( \32986 , \32984 , \32985 );
not \U$32734 ( \32987 , \8252 );
and \U$32735 ( \32988 , \32986 , \32987 );
not \U$32736 ( \32989 , \32986 );
and \U$32737 ( \32990 , \32989 , \5754 );
nor \U$32738 ( \32991 , \32988 , \32990 );
nand \U$32739 ( \32992 , \32981 , \32991 );
nand \U$32740 ( \32993 , \32980 , \32992 );
not \U$32741 ( \32994 , \32993 );
and \U$32742 ( \32995 , \32959 , \32994 );
not \U$32743 ( \32996 , RIbe29560_57);
not \U$32744 ( \32997 , \10949 );
or \U$32745 ( \32998 , \32996 , \32997 );
nand \U$32746 ( \32999 , \8269 , RIbe28228_16);
nand \U$32747 ( \33000 , \32998 , \32999 );
not \U$32748 ( \33001 , \33000 );
not \U$32749 ( \33002 , \7984 );
and \U$32750 ( \33003 , \33001 , \33002 );
and \U$32751 ( \33004 , \33000 , \6948 );
nor \U$32752 ( \33005 , \33003 , \33004 );
not \U$32753 ( \33006 , RIbe29290_51);
not \U$32754 ( \33007 , \7954 );
or \U$32755 ( \33008 , \33006 , \33007 );
nand \U$32756 ( \33009 , \7958 , RIbe28a20_33);
nand \U$32757 ( \33010 , \33008 , \33009 );
xor \U$32758 ( \33011 , \33010 , \6572 );
nand \U$32759 ( \33012 , \33005 , \33011 );
not \U$32760 ( \33013 , RIbe289a8_32);
not \U$32761 ( \33014 , \7299 );
or \U$32762 ( \33015 , \33013 , \33014 );
nand \U$32763 ( \33016 , \6985 , RIbe28930_31);
nand \U$32764 ( \33017 , \33015 , \33016 );
xnor \U$32765 ( \33018 , \33017 , \13168 );
and \U$32766 ( \33019 , \33012 , \33018 );
nor \U$32767 ( \33020 , \33005 , \33011 );
nor \U$32768 ( \33021 , \33019 , \33020 );
nor \U$32769 ( \33022 , \32995 , \33021 );
and \U$32770 ( \33023 , \32993 , \32958 );
nor \U$32771 ( \33024 , \33022 , \33023 );
not \U$32772 ( \33025 , \33024 );
or \U$32773 ( \33026 , \32925 , \33025 );
not \U$32774 ( \33027 , RIbe29920_65);
not \U$32775 ( \33028 , \12787 );
or \U$32776 ( \33029 , \33027 , \33028 );
nand \U$32777 ( \33030 , \12794 , RIbe27b98_2);
nand \U$32778 ( \33031 , \33029 , \33030 );
and \U$32779 ( \33032 , \33031 , \12893 );
not \U$32780 ( \33033 , \33031 );
and \U$32781 ( \33034 , \33033 , \14103 );
nor \U$32782 ( \33035 , \33032 , \33034 );
nand \U$32783 ( \33036 , \33035 , RIbe2aeb0_111);
not \U$32784 ( \33037 , \33036 );
not \U$32785 ( \33038 , RIbe28e58_42);
not \U$32786 ( \33039 , \18608 );
or \U$32787 ( \33040 , \33038 , \33039 );
nand \U$32788 ( \33041 , \12835 , RIbe28de0_41);
nand \U$32789 ( \33042 , \33040 , \33041 );
and \U$32790 ( \33043 , \33042 , \14555 );
not \U$32791 ( \33044 , \33042 );
and \U$32792 ( \33045 , \33044 , \12823 );
nor \U$32793 ( \33046 , \33043 , \33045 );
not \U$32794 ( \33047 , \33046 );
or \U$32795 ( \33048 , \33037 , \33047 );
or \U$32796 ( \33049 , RIbe2aeb0_111, \33035 );
nand \U$32797 ( \33050 , \33048 , \33049 );
not \U$32798 ( \33051 , \33050 );
not \U$32799 ( \33052 , \33051 );
not \U$32800 ( \33053 , RIbe27d00_5);
not \U$32801 ( \33054 , \14071 );
or \U$32802 ( \33055 , \33053 , \33054 );
nand \U$32803 ( \33056 , \13077 , RIbe27c10_3);
nand \U$32804 ( \33057 , \33055 , \33056 );
and \U$32805 ( \33058 , \33057 , \13570 );
not \U$32806 ( \33059 , \33057 );
and \U$32807 ( \33060 , \33059 , \12746 );
nor \U$32808 ( \33061 , \33058 , \33060 );
not \U$32809 ( \33062 , \33061 );
not \U$32810 ( \33063 , \33062 );
not \U$32811 ( \33064 , RIbe29a88_68);
not \U$32812 ( \33065 , \15573 );
or \U$32813 ( \33066 , \33064 , \33065 );
nand \U$32814 ( \33067 , \13728 , RIbe27d78_6);
nand \U$32815 ( \33068 , \33066 , \33067 );
xor \U$32816 ( \33069 , \33068 , \12723 );
not \U$32817 ( \33070 , \33069 );
or \U$32818 ( \33071 , \33063 , \33070 );
not \U$32819 ( \33072 , \13087 );
not \U$32820 ( \33073 , \4545 );
and \U$32821 ( \33074 , \33072 , \33073 );
and \U$32822 ( \33075 , \12765 , RIbe28fc0_45);
nor \U$32823 ( \33076 , \33074 , \33075 );
and \U$32824 ( \33077 , \33076 , \12770 );
not \U$32825 ( \33078 , \33076 );
and \U$32826 ( \33079 , \33078 , \12774 );
nor \U$32827 ( \33080 , \33077 , \33079 );
nand \U$32828 ( \33081 , \33071 , \33080 );
not \U$32829 ( \33082 , \33069 );
nand \U$32830 ( \33083 , \33082 , \33061 );
nand \U$32831 ( \33084 , \33081 , \33083 );
not \U$32832 ( \33085 , \33084 );
not \U$32833 ( \33086 , \33085 );
or \U$32834 ( \33087 , \33052 , \33086 );
not \U$32835 ( \33088 , RIbe29830_63);
not \U$32836 ( \33089 , \10936 );
or \U$32837 ( \33090 , \33088 , \33089 );
nand \U$32838 ( \33091 , \12213 , RIbe296c8_60);
nand \U$32839 ( \33092 , \33090 , \33091 );
not \U$32840 ( \33093 , \33092 );
not \U$32841 ( \33094 , \12218 );
and \U$32842 ( \33095 , \33093 , \33094 );
and \U$32843 ( \33096 , \33092 , \10943 );
nor \U$32844 ( \33097 , \33095 , \33096 );
not \U$32845 ( \33098 , \33097 );
and \U$32846 ( \33099 , \13036 , RIbe281b0_15);
and \U$32847 ( \33100 , \9914 , RIbe280c0_13);
nor \U$32848 ( \33101 , \33099 , \33100 );
and \U$32849 ( \33102 , \33101 , \16059 );
not \U$32850 ( \33103 , \33101 );
and \U$32851 ( \33104 , \33103 , \16994 );
nor \U$32852 ( \33105 , \33102 , \33104 );
or \U$32853 ( \33106 , \33098 , \33105 );
not \U$32854 ( \33107 , \12960 );
not \U$32855 ( \33108 , RIbe29650_59);
not \U$32856 ( \33109 , \12943 );
or \U$32857 ( \33110 , \33108 , \33109 );
nand \U$32858 ( \33111 , \13669 , RIbe29038_46);
nand \U$32859 ( \33112 , \33110 , \33111 );
not \U$32860 ( \33113 , \33112 );
or \U$32861 ( \33114 , \33107 , \33113 );
or \U$32862 ( \33115 , \33112 , \17005 );
nand \U$32863 ( \33116 , \33114 , \33115 );
nand \U$32864 ( \33117 , \33106 , \33116 );
nand \U$32865 ( \33118 , \33105 , \33098 );
nand \U$32866 ( \33119 , \33117 , \33118 );
nand \U$32867 ( \33120 , \33087 , \33119 );
nand \U$32868 ( \33121 , \33084 , \33050 );
nand \U$32869 ( \33122 , \33120 , \33121 );
nand \U$32870 ( \33123 , \33026 , \33122 );
not \U$32871 ( \33124 , \33024 );
nand \U$32872 ( \33125 , \33124 , \32923 );
nand \U$32873 ( \33126 , \33123 , \33125 );
not \U$32874 ( \33127 , \33126 );
not \U$32875 ( \33128 , \33127 );
nand \U$32876 ( \33129 , RIbe29380_53, RIbe2aaf0_103);
not \U$32877 ( \33130 , \33129 );
not \U$32878 ( \33131 , RIbe2b630_127);
not \U$32879 ( \33132 , \12312 );
or \U$32880 ( \33133 , \33131 , \33132 );
nand \U$32881 ( \33134 , \329 , RIbe2b018_114);
nand \U$32882 ( \33135 , \33133 , \33134 );
xor \U$32883 ( \33136 , \33135 , \12321 );
not \U$32884 ( \33137 , \33136 );
or \U$32885 ( \33138 , \33130 , \33137 );
not \U$32886 ( \33139 , RIbe2afa0_113);
not \U$32887 ( \33140 , \260 );
or \U$32888 ( \33141 , \33139 , \33140 );
nand \U$32889 ( \33142 , \6325 , RIbe2af28_112);
nand \U$32890 ( \33143 , \33141 , \33142 );
xnor \U$32891 ( \33144 , \33143 , \1362 );
nand \U$32892 ( \33145 , \33138 , \33144 );
or \U$32893 ( \33146 , \33136 , \33129 );
nand \U$32894 ( \33147 , \33145 , \33146 );
xor \U$32895 ( \33148 , \32449 , \1374 );
xnor \U$32896 ( \33149 , \33148 , \32444 );
xor \U$32897 ( \33150 , \33147 , \33149 );
and \U$32898 ( \33151 , \546 , RIbe2b090_115);
and \U$32899 ( \33152 , \552 , RIbe2a280_85);
nor \U$32900 ( \33153 , \33151 , \33152 );
not \U$32901 ( \33154 , \33153 );
not \U$32902 ( \33155 , \425 );
and \U$32903 ( \33156 , \33154 , \33155 );
and \U$32904 ( \33157 , \33153 , \7123 );
nor \U$32905 ( \33158 , \33156 , \33157 );
not \U$32906 ( \33159 , \33158 );
and \U$32907 ( \33160 , \1679 , RIbe2b1f8_118);
and \U$32908 ( \33161 , \7116 , RIbe2b180_117);
nor \U$32909 ( \33162 , \33160 , \33161 );
and \U$32910 ( \33163 , \33162 , \293 );
not \U$32911 ( \33164 , \33162 );
and \U$32912 ( \33165 , \33164 , \300 );
nor \U$32913 ( \33166 , \33163 , \33165 );
not \U$32914 ( \33167 , \33166 );
or \U$32915 ( \33168 , \33159 , \33167 );
not \U$32916 ( \33169 , RIbe2b270_119);
not \U$32917 ( \33170 , \9239 );
or \U$32918 ( \33171 , \33169 , \33170 );
nand \U$32919 ( \33172 , \428 , RIbe2b108_116);
nand \U$32920 ( \33173 , \33171 , \33172 );
and \U$32921 ( \33174 , \33173 , \306 );
not \U$32922 ( \33175 , \33173 );
and \U$32923 ( \33176 , \33175 , \312 );
nor \U$32924 ( \33177 , \33174 , \33176 );
nand \U$32925 ( \33178 , \33168 , \33177 );
not \U$32926 ( \33179 , \33158 );
not \U$32927 ( \33180 , \33166 );
nand \U$32928 ( \33181 , \33179 , \33180 );
nand \U$32929 ( \33182 , \33178 , \33181 );
and \U$32930 ( \33183 , \33150 , \33182 );
and \U$32931 ( \33184 , \33147 , \33149 );
or \U$32932 ( \33185 , \33183 , \33184 );
not \U$32933 ( \33186 , \33185 );
not \U$32934 ( \33187 , \33186 );
xor \U$32935 ( \33188 , \32128 , \32138 );
and \U$32936 ( \33189 , \33188 , \32148 );
not \U$32937 ( \33190 , \33188 );
not \U$32938 ( \33191 , \32148 );
and \U$32939 ( \33192 , \33190 , \33191 );
nor \U$32940 ( \33193 , \33189 , \33192 );
not \U$32941 ( \33194 , \33193 );
xor \U$32942 ( \33195 , \32342 , \32353 );
xor \U$32943 ( \33196 , \33195 , \32333 );
not \U$32944 ( \33197 , \33196 );
or \U$32945 ( \33198 , \33194 , \33197 );
xor \U$32946 ( \33199 , \32398 , \32407 );
xor \U$32947 ( \33200 , \33199 , \32417 );
nand \U$32948 ( \33201 , \33198 , \33200 );
not \U$32949 ( \33202 , \33196 );
not \U$32950 ( \33203 , \33193 );
nand \U$32951 ( \33204 , \33202 , \33203 );
nand \U$32952 ( \33205 , \33201 , \33204 );
not \U$32953 ( \33206 , \33205 );
not \U$32954 ( \33207 , \33206 );
or \U$32955 ( \33208 , \33187 , \33207 );
xor \U$32956 ( \33209 , \32463 , \32472 );
xor \U$32957 ( \33210 , \33209 , \32480 );
xor \U$32958 ( \33211 , \32213 , \32225 );
xor \U$32959 ( \33212 , \33211 , \32202 );
xor \U$32960 ( \33213 , \33210 , \33212 );
not \U$32961 ( \33214 , \32177 );
not \U$32962 ( \33215 , \32187 );
or \U$32963 ( \33216 , \33214 , \33215 );
nand \U$32964 ( \33217 , \32161 , \32186 );
nand \U$32965 ( \33218 , \33216 , \33217 );
and \U$32966 ( \33219 , \33218 , \32173 );
not \U$32967 ( \33220 , \33218 );
and \U$32968 ( \33221 , \33220 , \32172 );
nor \U$32969 ( \33222 , \33219 , \33221 );
and \U$32970 ( \33223 , \33213 , \33222 );
and \U$32971 ( \33224 , \33210 , \33212 );
or \U$32972 ( \33225 , \33223 , \33224 );
nand \U$32973 ( \33226 , \33208 , \33225 );
not \U$32974 ( \33227 , \33206 );
nand \U$32975 ( \33228 , \33227 , \33185 );
nand \U$32976 ( \33229 , \33226 , \33228 );
not \U$32977 ( \33230 , \33229 );
not \U$32978 ( \33231 , \33230 );
or \U$32979 ( \33232 , \33128 , \33231 );
xor \U$32980 ( \33233 , \32714 , \32722 );
xor \U$32981 ( \33234 , \33233 , \32732 );
xor \U$32982 ( \33235 , \12998 , \32661 );
xor \U$32983 ( \33236 , \33235 , \32672 );
xor \U$32984 ( \33237 , \33234 , \33236 );
not \U$32985 ( \33238 , \32255 );
not \U$32986 ( \33239 , \32244 );
or \U$32987 ( \33240 , \33238 , \33239 );
or \U$32988 ( \33241 , \32255 , \32244 );
nand \U$32989 ( \33242 , \33240 , \33241 );
buf \U$32990 ( \33243 , \32238 );
xnor \U$32991 ( \33244 , \33242 , \33243 );
xor \U$32992 ( \33245 , \32367 , \32376 );
xor \U$32993 ( \33246 , \33245 , \32386 );
or \U$32994 ( \33247 , \33244 , \33246 );
not \U$32995 ( \33248 , \32306 );
not \U$32996 ( \33249 , \32318 );
or \U$32997 ( \33250 , \33248 , \33249 );
nand \U$32998 ( \33251 , \32317 , \32305 );
nand \U$32999 ( \33252 , \33250 , \33251 );
not \U$33000 ( \33253 , \32296 );
and \U$33001 ( \33254 , \33252 , \33253 );
not \U$33002 ( \33255 , \33252 );
and \U$33003 ( \33256 , \33255 , \32296 );
nor \U$33004 ( \33257 , \33254 , \33256 );
nand \U$33005 ( \33258 , \33247 , \33257 );
nand \U$33006 ( \33259 , \33244 , \33246 );
nand \U$33007 ( \33260 , \33258 , \33259 );
xor \U$33008 ( \33261 , \33237 , \33260 );
xor \U$33009 ( \33262 , \32750 , \32759 );
xor \U$33010 ( \33263 , \33262 , \32769 );
xor \U$33011 ( \33264 , \32682 , \32691 );
xor \U$33012 ( \33265 , \33264 , \32701 );
xor \U$33013 ( \33266 , \33263 , \33265 );
xor \U$33014 ( \33267 , \32782 , \32791 );
xor \U$33015 ( \33268 , \33267 , \32801 );
xor \U$33016 ( \33269 , \33266 , \33268 );
and \U$33017 ( \33270 , \33261 , \33269 );
and \U$33018 ( \33271 , \33237 , \33260 );
or \U$33019 ( \33272 , \33270 , \33271 );
nand \U$33020 ( \33273 , \33232 , \33272 );
nand \U$33021 ( \33274 , \33229 , \33126 );
nand \U$33022 ( \33275 , \33273 , \33274 );
xor \U$33023 ( \33276 , \32828 , \33275 );
xor \U$33024 ( \33277 , \32439 , \32450 );
and \U$33025 ( \33278 , \33277 , \32483 );
and \U$33026 ( \33279 , \32439 , \32450 );
or \U$33027 ( \33280 , \33278 , \33279 );
not \U$33028 ( \33281 , \32587 );
not \U$33029 ( \33282 , \32615 );
or \U$33030 ( \33283 , \33281 , \33282 );
or \U$33031 ( \33284 , \32615 , \32587 );
nand \U$33032 ( \33285 , \33284 , \32646 );
nand \U$33033 ( \33286 , \33283 , \33285 );
xor \U$33034 ( \33287 , \33280 , \33286 );
nor \U$33035 ( \33288 , \32580 , \32514 );
or \U$33036 ( \33289 , \33288 , \32548 );
nand \U$33037 ( \33290 , \32580 , \32514 );
nand \U$33038 ( \33291 , \33289 , \33290 );
xnor \U$33039 ( \33292 , \33287 , \33291 );
not \U$33040 ( \33293 , \33292 );
and \U$33041 ( \33294 , \33234 , \33236 );
xor \U$33042 ( \33295 , \33263 , \33265 );
and \U$33043 ( \33296 , \33295 , \33268 );
and \U$33044 ( \33297 , \33263 , \33265 );
or \U$33045 ( \33298 , \33296 , \33297 );
xor \U$33046 ( \33299 , \33294 , \33298 );
not \U$33047 ( \33300 , RIbe28228_16);
not \U$33048 ( \33301 , \6980 );
or \U$33049 ( \33302 , \33300 , \33301 );
nand \U$33050 ( \33303 , \10898 , RIbe281b0_15);
nand \U$33051 ( \33304 , \33302 , \33303 );
and \U$33052 ( \33305 , \33304 , \6992 );
not \U$33053 ( \33306 , \33304 );
and \U$33054 ( \33307 , \33306 , \7304 );
or \U$33055 ( \33308 , \33305 , \33307 );
not \U$33056 ( \33309 , \33308 );
not \U$33057 ( \33310 , RIbe280c0_13);
not \U$33058 ( \33311 , \7974 );
or \U$33059 ( \33312 , \33310 , \33311 );
nand \U$33060 ( \33313 , RIbe29830_63, \13158 );
nand \U$33061 ( \33314 , \33312 , \33313 );
and \U$33062 ( \33315 , \33314 , \7984 );
not \U$33063 ( \33316 , \33314 );
and \U$33064 ( \33317 , \33316 , \14299 );
nor \U$33065 ( \33318 , \33315 , \33317 );
not \U$33066 ( \33319 , \33318 );
and \U$33067 ( \33320 , \8276 , RIbe296c8_60);
and \U$33068 ( \33321 , \13038 , RIbe29650_59);
nor \U$33069 ( \33322 , \33320 , \33321 );
and \U$33070 ( \33323 , \33322 , \7970 );
not \U$33071 ( \33324 , \33322 );
and \U$33072 ( \33325 , \33324 , \7971 );
nor \U$33073 ( \33326 , \33323 , \33325 );
not \U$33074 ( \33327 , \33326 );
not \U$33075 ( \33328 , \33327 );
or \U$33076 ( \33329 , \33319 , \33328 );
not \U$33077 ( \33330 , \33318 );
nand \U$33078 ( \33331 , \33330 , \33326 );
nand \U$33079 ( \33332 , \33329 , \33331 );
not \U$33080 ( \33333 , \33332 );
not \U$33081 ( \33334 , \33333 );
or \U$33082 ( \33335 , \33309 , \33334 );
not \U$33083 ( \33336 , \33308 );
nand \U$33084 ( \33337 , \33332 , \33336 );
nand \U$33085 ( \33338 , \33335 , \33337 );
not \U$33086 ( \33339 , RIbe290b0_47);
not \U$33087 ( \33340 , \12941 );
or \U$33088 ( \33341 , \33339 , \33340 );
nand \U$33089 ( \33342 , \12947 , RIbe29a88_68);
nand \U$33090 ( \33343 , \33341 , \33342 );
not \U$33091 ( \33344 , \33343 );
not \U$33092 ( \33345 , \12956 );
and \U$33093 ( \33346 , \33344 , \33345 );
and \U$33094 ( \33347 , \33343 , \12956 );
nor \U$33095 ( \33348 , \33346 , \33347 );
not \U$33096 ( \33349 , \12751 );
not \U$33097 ( \33350 , RIbe27d00_5);
not \U$33098 ( \33351 , \33350 );
and \U$33099 ( \33352 , \33349 , \33351 );
and \U$33100 ( \33353 , \20520 , RIbe27d78_6);
nor \U$33101 ( \33354 , \33352 , \33353 );
and \U$33102 ( \33355 , \33354 , \26172 );
not \U$33103 ( \33356 , \33354 );
and \U$33104 ( \33357 , \33356 , \12773 );
nor \U$33105 ( \33358 , \33355 , \33357 );
and \U$33106 ( \33359 , \33348 , \33358 );
not \U$33107 ( \33360 , \33348 );
not \U$33108 ( \33361 , \33358 );
and \U$33109 ( \33362 , \33360 , \33361 );
or \U$33110 ( \33363 , \33359 , \33362 );
not \U$33111 ( \33364 , RIbe29038_46);
not \U$33112 ( \33365 , \10936 );
or \U$33113 ( \33366 , \33364 , \33365 );
nand \U$33114 ( \33367 , \12212 , RIbe28fc0_45);
nand \U$33115 ( \33368 , \33366 , \33367 );
and \U$33116 ( \33369 , \33368 , \13030 );
not \U$33117 ( \33370 , \33368 );
and \U$33118 ( \33371 , \33370 , \9902 );
nor \U$33119 ( \33372 , \33369 , \33371 );
not \U$33120 ( \33373 , \33372 );
and \U$33121 ( \33374 , \33363 , \33373 );
not \U$33122 ( \33375 , \33363 );
and \U$33123 ( \33376 , \33375 , \33372 );
nor \U$33124 ( \33377 , \33374 , \33376 );
not \U$33125 ( \33378 , \33377 );
and \U$33126 ( \33379 , \33338 , \33378 );
not \U$33127 ( \33380 , \33338 );
and \U$33128 ( \33381 , \33380 , \33377 );
nor \U$33129 ( \33382 , \33379 , \33381 );
not \U$33130 ( \33383 , RIbe28de0_41);
not \U$33131 ( \33384 , \14071 );
or \U$33132 ( \33385 , \33383 , \33384 );
not \U$33133 ( \33386 , \1636 );
nand \U$33134 ( \33387 , \33386 , \12735 );
nand \U$33135 ( \33388 , \33385 , \33387 );
and \U$33136 ( \33389 , \33388 , \12743 );
not \U$33137 ( \33390 , \33388 );
and \U$33138 ( \33391 , \33390 , \12746 );
nor \U$33139 ( \33392 , \33389 , \33391 );
not \U$33140 ( \33393 , \33392 );
not \U$33141 ( \33394 , \33393 );
nor \U$33142 ( \33395 , \18607 , \1640 );
not \U$33143 ( \33396 , \33395 );
not \U$33144 ( \33397 , \16366 );
and \U$33145 ( \33398 , \33396 , \33397 );
and \U$33146 ( \33399 , \33395 , \15263 );
nor \U$33147 ( \33400 , \33398 , \33399 );
not \U$33148 ( \33401 , \33400 );
not \U$33149 ( \33402 , \33401 );
or \U$33150 ( \33403 , \33394 , \33402 );
nand \U$33151 ( \33404 , \33392 , \33400 );
nand \U$33152 ( \33405 , \33403 , \33404 );
not \U$33153 ( \33406 , \33405 );
not \U$33154 ( \33407 , RIbe27c10_3);
not \U$33155 ( \33408 , \16383 );
or \U$33156 ( \33409 , \33407 , \33408 );
nand \U$33157 ( \33410 , \12711 , RIbe28e58_42);
nand \U$33158 ( \33411 , \33409 , \33410 );
and \U$33159 ( \33412 , \33411 , \12723 );
not \U$33160 ( \33413 , \33411 );
and \U$33161 ( \33414 , \33413 , \12716 );
nor \U$33162 ( \33415 , \33412 , \33414 );
buf \U$33163 ( \33416 , \33415 );
and \U$33164 ( \33417 , \33406 , \33416 );
not \U$33165 ( \33418 , \33406 );
not \U$33166 ( \33419 , \33415 );
and \U$33167 ( \33420 , \33418 , \33419 );
nor \U$33168 ( \33421 , \33417 , \33420 );
not \U$33169 ( \33422 , \33421 );
and \U$33170 ( \33423 , \33382 , \33422 );
not \U$33171 ( \33424 , \33382 );
and \U$33172 ( \33425 , \33424 , \33421 );
nor \U$33173 ( \33426 , \33423 , \33425 );
xor \U$33174 ( \33427 , \33299 , \33426 );
not \U$33175 ( \33428 , \33427 );
not \U$33176 ( \33429 , \33428 );
or \U$33177 ( \33430 , \33293 , \33429 );
nand \U$33178 ( \33431 , RIbe29380_53, RIbe2afa0_113);
nor \U$33179 ( \33432 , \32645 , \32625 );
or \U$33180 ( \33433 , \33432 , \32634 );
nand \U$33181 ( \33434 , \32625 , \32645 );
nand \U$33182 ( \33435 , \33433 , \33434 );
xor \U$33183 ( \33436 , \33431 , \33435 );
not \U$33184 ( \33437 , RIbe2af28_112);
not \U$33185 ( \33438 , \325 );
or \U$33186 ( \33439 , \33437 , \33438 );
nand \U$33187 ( \33440 , \330 , RIbe2b1f8_118);
nand \U$33188 ( \33441 , \33439 , \33440 );
and \U$33189 ( \33442 , \33441 , \1379 );
not \U$33190 ( \33443 , \33441 );
and \U$33191 ( \33444 , \33443 , \1375 );
nor \U$33192 ( \33445 , \33442 , \33444 );
not \U$33193 ( \33446 , \33445 );
not \U$33194 ( \33447 , RIbe2b180_117);
not \U$33195 ( \33448 , \260 );
or \U$33196 ( \33449 , \33447 , \33448 );
nand \U$33197 ( \33450 , \263 , RIbe2b270_119);
nand \U$33198 ( \33451 , \33449 , \33450 );
xor \U$33199 ( \33452 , \33451 , \6058 );
not \U$33200 ( \33453 , \33452 );
and \U$33201 ( \33454 , \6311 , RIbe2b108_116);
and \U$33202 ( \33455 , \7116 , RIbe2b090_115);
nor \U$33203 ( \33456 , \33454 , \33455 );
and \U$33204 ( \33457 , \33456 , \300 );
not \U$33205 ( \33458 , \33456 );
and \U$33206 ( \33459 , \33458 , \293 );
nor \U$33207 ( \33460 , \33457 , \33459 );
not \U$33208 ( \33461 , \33460 );
or \U$33209 ( \33462 , \33453 , \33461 );
or \U$33210 ( \33463 , \33460 , \33452 );
nand \U$33211 ( \33464 , \33462 , \33463 );
not \U$33212 ( \33465 , \33464 );
or \U$33213 ( \33466 , \33446 , \33465 );
or \U$33214 ( \33467 , \33464 , \33445 );
nand \U$33215 ( \33468 , \33466 , \33467 );
xor \U$33216 ( \33469 , \33436 , \33468 );
not \U$33217 ( \33470 , RIbe2a190_83);
not \U$33218 ( \33471 , \546 );
or \U$33219 ( \33472 , \33470 , \33471 );
nand \U$33220 ( \33473 , \1327 , RIbe2a5c8_92);
nand \U$33221 ( \33474 , \33472 , \33473 );
not \U$33222 ( \33475 , \33474 );
not \U$33223 ( \33476 , \424 );
and \U$33224 ( \33477 , \33475 , \33476 );
and \U$33225 ( \33478 , \6340 , \33474 );
nor \U$33226 ( \33479 , \33477 , \33478 );
not \U$33227 ( \33480 , RIbe2a550_91);
not \U$33228 ( \33481 , \32589 );
or \U$33229 ( \33482 , \33480 , \33481 );
nand \U$33230 ( \33483 , \1179 , RIbe2a988_100);
nand \U$33231 ( \33484 , \33482 , \33483 );
not \U$33232 ( \33485 , \33484 );
not \U$33233 ( \33486 , \564 );
and \U$33234 ( \33487 , \33485 , \33486 );
and \U$33235 ( \33488 , \33484 , \1618 );
nor \U$33236 ( \33489 , \33487 , \33488 );
xor \U$33237 ( \33490 , \33479 , \33489 );
not \U$33238 ( \33491 , RIbe2a280_85);
not \U$33239 ( \33492 , \1223 );
or \U$33240 ( \33493 , \33491 , \33492 );
nand \U$33241 ( \33494 , \429 , RIbe2a208_84);
nand \U$33242 ( \33495 , \33493 , \33494 );
and \U$33243 ( \33496 , \33495 , \313 );
not \U$33244 ( \33497 , \33495 );
and \U$33245 ( \33498 , \33497 , \306 );
nor \U$33246 ( \33499 , \33496 , \33498 );
xnor \U$33247 ( \33500 , \33490 , \33499 );
not \U$33248 ( \33501 , \4064 );
not \U$33249 ( \33502 , \15612 );
and \U$33250 ( \33503 , \33501 , \33502 );
and \U$33251 ( \33504 , \8833 , RIbe29e48_76);
nor \U$33252 ( \33505 , \33503 , \33504 );
and \U$33253 ( \33506 , \33505 , \9083 );
not \U$33254 ( \33507 , \33505 );
and \U$33255 ( \33508 , \33507 , \1076 );
nor \U$33256 ( \33509 , \33506 , \33508 );
not \U$33257 ( \33510 , RIbe29c68_72);
not \U$33258 ( \33511 , \7007 );
or \U$33259 ( \33512 , \33510 , \33511 );
nand \U$33260 ( \33513 , \2900 , RIbe29bf0_71);
nand \U$33261 ( \33514 , \33512 , \33513 );
and \U$33262 ( \33515 , \33514 , \4058 );
not \U$33263 ( \33516 , \33514 );
and \U$33264 ( \33517 , \33516 , \2379 );
nor \U$33265 ( \33518 , \33515 , \33517 );
xor \U$33266 ( \33519 , \33509 , \33518 );
and \U$33267 ( \33520 , \1286 , RIbe2a028_80);
and \U$33268 ( \33521 , \1117 , RIbe29fb0_79);
nor \U$33269 ( \33522 , \33520 , \33521 );
and \U$33270 ( \33523 , \33522 , \1131 );
not \U$33271 ( \33524 , \33522 );
and \U$33272 ( \33525 , \33524 , \2563 );
nor \U$33273 ( \33526 , \33523 , \33525 );
xor \U$33274 ( \33527 , \33519 , \33526 );
not \U$33275 ( \33528 , RIbe2a2f8_86);
not \U$33276 ( \33529 , \1298 );
or \U$33277 ( \33530 , \33528 , \33529 );
nand \U$33278 ( \33531 , \1099 , RIbe2acd0_107);
nand \U$33279 ( \33532 , \33530 , \33531 );
and \U$33280 ( \33533 , \33532 , \4251 );
not \U$33281 ( \33534 , \33532 );
and \U$33282 ( \33535 , \33534 , \1309 );
nor \U$33283 ( \33536 , \33533 , \33535 );
not \U$33284 ( \33537 , RIbe2a3e8_88);
not \U$33285 ( \33538 , \4257 );
or \U$33286 ( \33539 , \33537 , \33538 );
nand \U$33287 ( \33540 , \1146 , RIbe2a370_87);
nand \U$33288 ( \33541 , \33539 , \33540 );
and \U$33289 ( \33542 , \33541 , \1652 );
not \U$33290 ( \33543 , \33541 );
and \U$33291 ( \33544 , \33543 , \1153 );
nor \U$33292 ( \33545 , \33542 , \33544 );
and \U$33293 ( \33546 , \33536 , \33545 );
not \U$33294 ( \33547 , \33536 );
not \U$33295 ( \33548 , \33545 );
and \U$33296 ( \33549 , \33547 , \33548 );
or \U$33297 ( \33550 , \33546 , \33549 );
not \U$33298 ( \33551 , \1608 );
not \U$33299 ( \33552 , RIbe2a910_99);
not \U$33300 ( \33553 , \2424 );
or \U$33301 ( \33554 , \33552 , \33553 );
nand \U$33302 ( \33555 , \2000 , RIbe2b5b8_126);
nand \U$33303 ( \33556 , \33554 , \33555 );
not \U$33304 ( \33557 , \33556 );
and \U$33305 ( \33558 , \33551 , \33557 );
and \U$33306 ( \33559 , \33556 , \1813 );
nor \U$33307 ( \33560 , \33558 , \33559 );
xor \U$33308 ( \33561 , \33550 , \33560 );
and \U$33309 ( \33562 , \33527 , \33561 );
not \U$33310 ( \33563 , \33527 );
not \U$33311 ( \33564 , \33561 );
and \U$33312 ( \33565 , \33563 , \33564 );
or \U$33313 ( \33566 , \33562 , \33565 );
xor \U$33314 ( \33567 , \33500 , \33566 );
xor \U$33315 ( \33568 , \33469 , \33567 );
nand \U$33316 ( \33569 , \3701 , RIbe27fd0_11);
or \U$33317 ( \33570 , \33569 , \20767 );
nand \U$33318 ( \33571 , \4026 , RIbe27f58_10);
nand \U$33319 ( \33572 , \33570 , \33571 );
and \U$33320 ( \33573 , \33572 , \3471 );
not \U$33321 ( \33574 , \33572 );
and \U$33322 ( \33575 , \33574 , \3698 );
nor \U$33323 ( \33576 , \33573 , \33575 );
not \U$33324 ( \33577 , RIbe27e68_8);
not \U$33325 ( \33578 , \6414 );
or \U$33326 ( \33579 , \33577 , \33578 );
nand \U$33327 ( \33580 , \4600 , RIbe28660_25);
nand \U$33328 ( \33581 , \33579 , \33580 );
and \U$33329 ( \33582 , \33581 , \4007 );
not \U$33330 ( \33583 , \33581 );
and \U$33331 ( \33584 , \33583 , \4323 );
nor \U$33332 ( \33585 , \33582 , \33584 );
xor \U$33333 ( \33586 , \33576 , \33585 );
not \U$33334 ( \33587 , RIbe28f48_44);
not \U$33335 ( \33588 , \4764 );
or \U$33336 ( \33589 , \33587 , \33588 );
nand \U$33337 ( \33590 , \3458 , RIbe28ed0_43);
nand \U$33338 ( \33591 , \33589 , \33590 );
and \U$33339 ( \33592 , \33591 , \3290 );
not \U$33340 ( \33593 , \33591 );
and \U$33341 ( \33594 , \33593 , \3461 );
nor \U$33342 ( \33595 , \33592 , \33594 );
xor \U$33343 ( \33596 , \33586 , \33595 );
and \U$33344 ( \33597 , \5453 , RIbe28480_21);
not \U$33345 ( \33598 , \33597 );
not \U$33346 ( \33599 , \5750 );
or \U$33347 ( \33600 , \33598 , \33599 );
nand \U$33348 ( \33601 , RIbe28408_20, \6634 );
nand \U$33349 ( \33602 , \33600 , \33601 );
not \U$33350 ( \33603 , \33602 );
not \U$33351 ( \33604 , \10984 );
or \U$33352 ( \33605 , \33603 , \33604 );
or \U$33353 ( \33606 , \33602 , \8252 );
nand \U$33354 ( \33607 , \33605 , \33606 );
not \U$33355 ( \33608 , RIbe28390_19);
not \U$33356 ( \33609 , \6138 );
or \U$33357 ( \33610 , \33608 , \33609 );
nand \U$33358 ( \33611 , \7087 , RIbe28b10_35);
nand \U$33359 ( \33612 , \33610 , \33611 );
and \U$33360 ( \33613 , \33612 , \5741 );
not \U$33361 ( \33614 , \33612 );
and \U$33362 ( \33615 , \33614 , \5740 );
nor \U$33363 ( \33616 , \33613 , \33615 );
xor \U$33364 ( \33617 , \33607 , \33616 );
not \U$33365 ( \33618 , RIbe285e8_24);
not \U$33366 ( \33619 , \5727 );
or \U$33367 ( \33620 , \33618 , \33619 );
nand \U$33368 ( \33621 , \5052 , RIbe287c8_28);
nand \U$33369 ( \33622 , \33620 , \33621 );
and \U$33370 ( \33623 , \33622 , \4586 );
not \U$33371 ( \33624 , \33622 );
and \U$33372 ( \33625 , \33624 , \4946 );
nor \U$33373 ( \33626 , \33623 , \33625 );
xor \U$33374 ( \33627 , \33617 , \33626 );
xor \U$33375 ( \33628 , \33596 , \33627 );
not \U$33376 ( \33629 , RIbe28a20_33);
not \U$33377 ( \33630 , \7941 );
or \U$33378 ( \33631 , \33629 , \33630 );
nand \U$33379 ( \33632 , \6596 , RIbe289a8_32);
nand \U$33380 ( \33633 , \33631 , \33632 );
and \U$33381 ( \33634 , \33633 , \6582 );
not \U$33382 ( \33635 , \33633 );
and \U$33383 ( \33636 , \33635 , \7271 );
nor \U$33384 ( \33637 , \33634 , \33636 );
not \U$33385 ( \33638 , RIbe28930_31);
not \U$33386 ( \33639 , \8199 );
or \U$33387 ( \33640 , \33638 , \33639 );
nand \U$33388 ( \33641 , \7958 , RIbe29560_57);
nand \U$33389 ( \33642 , \33640 , \33641 );
and \U$33390 ( \33643 , \33642 , \7293 );
not \U$33391 ( \33644 , \33642 );
and \U$33392 ( \33645 , \33644 , \6572 );
nor \U$33393 ( \33646 , \33643 , \33645 );
xor \U$33394 ( \33647 , \33637 , \33646 );
not \U$33395 ( \33648 , RIbe28b88_36);
not \U$33396 ( \33649 , \6536 );
or \U$33397 ( \33650 , \33648 , \33649 );
nand \U$33398 ( \33651 , \6540 , RIbe29290_51);
nand \U$33399 ( \33652 , \33650 , \33651 );
and \U$33400 ( \33653 , \33652 , \6546 );
not \U$33401 ( \33654 , \33652 );
and \U$33402 ( \33655 , \33654 , \6891 );
nor \U$33403 ( \33656 , \33653 , \33655 );
xor \U$33404 ( \33657 , \33647 , \33656 );
xor \U$33405 ( \33658 , \33628 , \33657 );
xor \U$33406 ( \33659 , \33568 , \33658 );
nand \U$33407 ( \33660 , \33430 , \33659 );
not \U$33408 ( \33661 , \33292 );
nand \U$33409 ( \33662 , \33661 , \33427 );
nand \U$33410 ( \33663 , \33660 , \33662 );
xor \U$33411 ( \33664 , \33276 , \33663 );
xor \U$33412 ( \33665 , \33294 , \33298 );
and \U$33413 ( \33666 , \33665 , \33426 );
and \U$33414 ( \33667 , \33294 , \33298 );
or \U$33415 ( \33668 , \33666 , \33667 );
not \U$33416 ( \33669 , \33280 );
not \U$33417 ( \33670 , \33286 );
or \U$33418 ( \33671 , \33669 , \33670 );
or \U$33419 ( \33672 , \33286 , \33280 );
nand \U$33420 ( \33673 , \33672 , \33291 );
nand \U$33421 ( \33674 , \33671 , \33673 );
or \U$33422 ( \33675 , \32357 , \32389 );
and \U$33423 ( \33676 , \33675 , \32420 );
and \U$33424 ( \33677 , \32357 , \32389 );
nor \U$33425 ( \33678 , \33676 , \33677 );
not \U$33426 ( \33679 , \33678 );
xor \U$33427 ( \33680 , \32258 , \32286 );
and \U$33428 ( \33681 , \33680 , \32321 );
and \U$33429 ( \33682 , \32258 , \32286 );
or \U$33430 ( \33683 , \33681 , \33682 );
not \U$33431 ( \33684 , \33683 );
or \U$33432 ( \33685 , \33679 , \33684 );
or \U$33433 ( \33686 , \32227 , \32190 );
not \U$33434 ( \33687 , \32190 );
not \U$33435 ( \33688 , \32227 );
or \U$33436 ( \33689 , \33687 , \33688 );
nand \U$33437 ( \33690 , \33689 , \32151 );
nand \U$33438 ( \33691 , \33686 , \33690 );
nand \U$33439 ( \33692 , \33685 , \33691 );
not \U$33440 ( \33693 , \33678 );
not \U$33441 ( \33694 , \33683 );
nand \U$33442 ( \33695 , \33693 , \33694 );
nand \U$33443 ( \33696 , \33692 , \33695 );
xor \U$33444 ( \33697 , \33674 , \33696 );
xor \U$33445 ( \33698 , \33668 , \33697 );
and \U$33446 ( \33699 , \6962 , \5423 );
not \U$33447 ( \33700 , \6962 );
nand \U$33448 ( \33701 , \6557 , RIbe28b88_36);
and \U$33449 ( \33702 , \33700 , \33701 );
or \U$33450 ( \33703 , \33699 , \33702 );
xnor \U$33451 ( \33704 , \33703 , \7293 );
not \U$33452 ( \33705 , \33704 );
and \U$33453 ( \33706 , RIbe28390_19, \6588 );
and \U$33454 ( \33707 , \7482 , \33706 );
not \U$33455 ( \33708 , \7482 );
and \U$33456 ( \33709 , \33708 , RIbe28b10_35);
nor \U$33457 ( \33710 , \33707 , \33709 );
and \U$33458 ( \33711 , \33710 , \7948 );
not \U$33459 ( \33712 , \33710 );
and \U$33460 ( \33713 , \33712 , \29121 );
nor \U$33461 ( \33714 , \33711 , \33713 );
nand \U$33462 ( \33715 , \33705 , \33714 );
not \U$33463 ( \33716 , \33715 );
not \U$33464 ( \33717 , RIbe28480_21);
not \U$33465 ( \33718 , \6536 );
or \U$33466 ( \33719 , \33717 , \33718 );
nand \U$33467 ( \33720 , \6540 , RIbe28408_20);
nand \U$33468 ( \33721 , \33719 , \33720 );
and \U$33469 ( \33722 , \33721 , \15730 );
not \U$33470 ( \33723 , \33721 );
and \U$33471 ( \33724 , \33723 , \13412 );
nor \U$33472 ( \33725 , \33722 , \33724 );
not \U$33473 ( \33726 , \33725 );
or \U$33474 ( \33727 , \33716 , \33726 );
not \U$33475 ( \33728 , \33714 );
nand \U$33476 ( \33729 , \33728 , \33704 );
nand \U$33477 ( \33730 , \33727 , \33729 );
and \U$33478 ( \33731 , \5453 , RIbe27e68_8);
or \U$33479 ( \33732 , \5749 , \33731 );
not \U$33480 ( \33733 , RIbe28660_25);
nand \U$33481 ( \33734 , \33733 , \6633 );
nand \U$33482 ( \33735 , \33732 , \33734 );
and \U$33483 ( \33736 , \33735 , \5754 );
not \U$33484 ( \33737 , \33735 );
not \U$33485 ( \33738 , \5046 );
and \U$33486 ( \33739 , \33737 , \33738 );
nor \U$33487 ( \33740 , \33736 , \33739 );
not \U$33488 ( \33741 , \33740 );
or \U$33489 ( \33742 , \6615 , RIbe287c8_28);
not \U$33490 ( \33743 , RIbe285e8_24);
not \U$33491 ( \33744 , \6134 );
or \U$33492 ( \33745 , \33743 , \33744 );
not \U$33493 ( \33746 , \8234 );
nand \U$33494 ( \33747 , \33745 , \33746 );
nand \U$33495 ( \33748 , \33742 , \33747 );
not \U$33496 ( \33749 , \33748 );
not \U$33497 ( \33750 , \21093 );
and \U$33498 ( \33751 , \33749 , \33750 );
and \U$33499 ( \33752 , \21093 , \33748 );
nor \U$33500 ( \33753 , \33751 , \33752 );
nand \U$33501 ( \33754 , \33741 , \33753 );
not \U$33502 ( \33755 , \33754 );
not \U$33503 ( \33756 , RIbe27fd0_11);
not \U$33504 ( \33757 , \6427 );
or \U$33505 ( \33758 , \33756 , \33757 );
nand \U$33506 ( \33759 , \7056 , RIbe27f58_10);
nand \U$33507 ( \33760 , \33758 , \33759 );
and \U$33508 ( \33761 , \33760 , \4586 );
not \U$33509 ( \33762 , \33760 );
and \U$33510 ( \33763 , \33762 , \4592 );
nor \U$33511 ( \33764 , \33761 , \33763 );
not \U$33512 ( \33765 , \33764 );
or \U$33513 ( \33766 , \33755 , \33765 );
not \U$33514 ( \33767 , \33753 );
nand \U$33515 ( \33768 , \33767 , \33740 );
nand \U$33516 ( \33769 , \33766 , \33768 );
or \U$33517 ( \33770 , \33730 , \33769 );
and \U$33518 ( \33771 , \13036 , RIbe28228_16);
and \U$33519 ( \33772 , \10919 , RIbe281b0_15);
nor \U$33520 ( \33773 , \33771 , \33772 );
and \U$33521 ( \33774 , \33773 , \8077 );
not \U$33522 ( \33775 , \33773 );
and \U$33523 ( \33776 , \33775 , \7970 );
nor \U$33524 ( \33777 , \33774 , \33776 );
not \U$33525 ( \33778 , \33777 );
not \U$33526 ( \33779 , RIbe28930_31);
not \U$33527 ( \33780 , \10949 );
or \U$33528 ( \33781 , \33779 , \33780 );
nand \U$33529 ( \33782 , \7981 , RIbe29560_57);
nand \U$33530 ( \33783 , \33781 , \33782 );
and \U$33531 ( \33784 , \33783 , \6948 );
not \U$33532 ( \33785 , \33783 );
and \U$33533 ( \33786 , \33785 , \7988 );
nor \U$33534 ( \33787 , \33784 , \33786 );
not \U$33535 ( \33788 , \33787 );
not \U$33536 ( \33789 , \33788 );
or \U$33537 ( \33790 , \33778 , \33789 );
or \U$33538 ( \33791 , \33788 , \33777 );
not \U$33539 ( \33792 , RIbe28a20_33);
not \U$33540 ( \33793 , \6980 );
or \U$33541 ( \33794 , \33792 , \33793 );
nand \U$33542 ( \33795 , \13224 , RIbe289a8_32);
nand \U$33543 ( \33796 , \33794 , \33795 );
and \U$33544 ( \33797 , \33796 , \6993 );
not \U$33545 ( \33798 , \33796 );
and \U$33546 ( \33799 , \33798 , \7661 );
nor \U$33547 ( \33800 , \33797 , \33799 );
nand \U$33548 ( \33801 , \33791 , \33800 );
nand \U$33549 ( \33802 , \33790 , \33801 );
and \U$33550 ( \33803 , \33770 , \33802 );
and \U$33551 ( \33804 , \33769 , \33730 );
nor \U$33552 ( \33805 , \33803 , \33804 );
not \U$33553 ( \33806 , \33805 );
not \U$33554 ( \33807 , RIbe29c68_72);
not \U$33555 ( \33808 , \20764 );
or \U$33556 ( \33809 , \33807 , \33808 );
nand \U$33557 ( \33810 , \8368 , RIbe29bf0_71);
nand \U$33558 ( \33811 , \33809 , \33810 );
not \U$33559 ( \33812 , \33811 );
not \U$33560 ( \33813 , \3698 );
and \U$33561 ( \33814 , \33812 , \33813 );
and \U$33562 ( \33815 , \33811 , \3698 );
nor \U$33563 ( \33816 , \33814 , \33815 );
not \U$33564 ( \33817 , \33816 );
not \U$33565 ( \33818 , RIbe29e48_76);
not \U$33566 ( \33819 , \3284 );
or \U$33567 ( \33820 , \33818 , \33819 );
nand \U$33568 ( \33821 , \3689 , RIbe29dd0_75);
nand \U$33569 ( \33822 , \33820 , \33821 );
xor \U$33570 ( \33823 , \33822 , \2887 );
not \U$33571 ( \33824 , \33823 );
or \U$33572 ( \33825 , \33817 , \33824 );
not \U$33573 ( \33826 , RIbe28f48_44);
not \U$33574 ( \33827 , \6414 );
or \U$33575 ( \33828 , \33826 , \33827 );
nand \U$33576 ( \33829 , \4600 , RIbe28ed0_43);
nand \U$33577 ( \33830 , \33828 , \33829 );
and \U$33578 ( \33831 , \33830 , \4326 );
not \U$33579 ( \33832 , \33830 );
and \U$33580 ( \33833 , \33832 , \4323 );
nor \U$33581 ( \33834 , \33831 , \33833 );
nand \U$33582 ( \33835 , \33825 , \33834 );
not \U$33583 ( \33836 , \33823 );
not \U$33584 ( \33837 , \33816 );
nand \U$33585 ( \33838 , \33836 , \33837 );
and \U$33586 ( \33839 , \1098 , RIbe2b5b8_126);
not \U$33587 ( \33840 , \1098 );
and \U$33588 ( \33841 , \1629 , RIbe2a910_99);
and \U$33589 ( \33842 , \33840 , \33841 );
nor \U$33590 ( \33843 , \33839 , \33842 );
not \U$33591 ( \33844 , \33843 );
not \U$33592 ( \33845 , \1309 );
and \U$33593 ( \33846 , \33844 , \33845 );
and \U$33594 ( \33847 , \33843 , \1309 );
nor \U$33595 ( \33848 , \33846 , \33847 );
not \U$33596 ( \33849 , RIbe2a190_83);
not \U$33597 ( \33850 , \23339 );
or \U$33598 ( \33851 , \33849 , \33850 );
nand \U$33599 ( \33852 , \1202 , RIbe2a5c8_92);
nand \U$33600 ( \33853 , \33851 , \33852 );
not \U$33601 ( \33854 , \33853 );
not \U$33602 ( \33855 , \1813 );
and \U$33603 ( \33856 , \33854 , \33855 );
and \U$33604 ( \33857 , \33853 , \1813 );
nor \U$33605 ( \33858 , \33856 , \33857 );
and \U$33606 ( \33859 , \33848 , \33858 );
not \U$33607 ( \33860 , \1652 );
and \U$33608 ( \33861 , \1146 , RIbe2a988_100);
not \U$33609 ( \33862 , \1146 );
and \U$33610 ( \33863 , \1140 , RIbe2a550_91);
and \U$33611 ( \33864 , \33862 , \33863 );
nor \U$33612 ( \33865 , \33861 , \33864 );
not \U$33613 ( \33866 , \33865 );
or \U$33614 ( \33867 , \33860 , \33866 );
or \U$33615 ( \33868 , \33865 , \7899 );
nand \U$33616 ( \33869 , \33867 , \33868 );
not \U$33617 ( \33870 , \33869 );
nor \U$33618 ( \33871 , \33859 , \33870 );
nor \U$33619 ( \33872 , \33858 , \33848 );
nor \U$33620 ( \33873 , \33871 , \33872 );
and \U$33621 ( \33874 , \33835 , \33838 , \33873 );
not \U$33622 ( \33875 , \24063 );
not \U$33623 ( \33876 , RIbe2a2f8_86);
not \U$33624 ( \33877 , RIbe295d8_58);
not \U$33625 ( \33878 , RIbe29740_61);
or \U$33626 ( \33879 , \33877 , \33878 );
or \U$33627 ( \33880 , RIbe29740_61, RIbe295d8_58);
nand \U$33628 ( \33881 , \33879 , \33880 );
nor \U$33629 ( \33882 , \33876 , \33881 );
or \U$33630 ( \33883 , \33882 , \2384 );
not \U$33631 ( \33884 , RIbe2acd0_107);
nand \U$33632 ( \33885 , \33884 , \2383 );
nand \U$33633 ( \33886 , \33883 , \33885 );
not \U$33634 ( \33887 , \33886 );
or \U$33635 ( \33888 , \33875 , \33887 );
or \U$33636 ( \33889 , \33886 , \1276 );
nand \U$33637 ( \33890 , \33888 , \33889 );
not \U$33638 ( \33891 , \33890 );
not \U$33639 ( \33892 , RIbe2a3e8_88);
not \U$33640 ( \33893 , \1112 );
or \U$33641 ( \33894 , \33892 , \33893 );
nand \U$33642 ( \33895 , \20664 , RIbe2a370_87);
nand \U$33643 ( \33896 , \33894 , \33895 );
and \U$33644 ( \33897 , \33896 , \6831 );
not \U$33645 ( \33898 , \33896 );
and \U$33646 ( \33899 , \33898 , \1131 );
nor \U$33647 ( \33900 , \33897 , \33899 );
not \U$33648 ( \33901 , \33900 );
not \U$33649 ( \33902 , \33901 );
or \U$33650 ( \33903 , \33891 , \33902 );
or \U$33651 ( \33904 , \33901 , \33890 );
and \U$33652 ( \33905 , \2900 , RIbe29fb0_79);
not \U$33653 ( \33906 , \2900 );
and \U$33654 ( \33907 , \2568 , RIbe2a028_80);
and \U$33655 ( \33908 , \33906 , \33907 );
nor \U$33656 ( \33909 , \33905 , \33908 );
not \U$33657 ( \33910 , \33909 );
not \U$33658 ( \33911 , \2573 );
and \U$33659 ( \33912 , \33910 , \33911 );
and \U$33660 ( \33913 , \33909 , \2380 );
nor \U$33661 ( \33914 , \33912 , \33913 );
not \U$33662 ( \33915 , \33914 );
nand \U$33663 ( \33916 , \33904 , \33915 );
nand \U$33664 ( \33917 , \33903 , \33916 );
not \U$33665 ( \33918 , \33917 );
nor \U$33666 ( \33919 , \33874 , \33918 );
and \U$33667 ( \33920 , \33835 , \33838 );
nor \U$33668 ( \33921 , \33920 , \33873 );
nor \U$33669 ( \33922 , \33919 , \33921 );
not \U$33670 ( \33923 , \33922 );
or \U$33671 ( \33924 , \33806 , \33923 );
not \U$33672 ( \33925 , \12893 );
not \U$33673 ( \33926 , RIbe28de0_41);
not \U$33674 ( \33927 , \13518 );
or \U$33675 ( \33928 , \33926 , \33927 );
nand \U$33676 ( \33929 , \12890 , RIbe29920_65);
nand \U$33677 ( \33930 , \33928 , \33929 );
not \U$33678 ( \33931 , \33930 );
or \U$33679 ( \33932 , \33925 , \33931 );
or \U$33680 ( \33933 , \33930 , \12893 );
nand \U$33681 ( \33934 , \33932 , \33933 );
and \U$33682 ( \33935 , \12811 , RIbe27b98_2);
nor \U$33683 ( \33936 , \33935 , \30890 );
nand \U$33684 ( \33937 , \33934 , \33936 );
not \U$33685 ( \33938 , \33937 );
not \U$33686 ( \33939 , \33938 );
not \U$33687 ( \33940 , RIbe29038_46);
not \U$33688 ( \33941 , RIbe2b4c8_124);
not \U$33689 ( \33942 , RIbe2b540_125);
or \U$33690 ( \33943 , \33941 , \33942 );
or \U$33691 ( \33944 , RIbe2b540_125, RIbe2b4c8_124);
nand \U$33692 ( \33945 , \33943 , \33944 );
nor \U$33693 ( \33946 , \33940 , \33945 );
or \U$33694 ( \33947 , \14491 , \33946 );
nand \U$33695 ( \33948 , \19749 , \1931 );
nand \U$33696 ( \33949 , \33947 , \33948 );
and \U$33697 ( \33950 , \33949 , \14000 );
not \U$33698 ( \33951 , \33949 );
and \U$33699 ( \33952 , \33951 , \12774 );
nor \U$33700 ( \33953 , \33950 , \33952 );
not \U$33701 ( \33954 , \33953 );
not \U$33702 ( \33955 , RIbe296c8_60);
not \U$33703 ( \33956 , RIbe2ad48_108);
not \U$33704 ( \33957 , RIbe2adc0_109);
or \U$33705 ( \33958 , \33956 , \33957 );
or \U$33706 ( \33959 , RIbe2adc0_109, RIbe2ad48_108);
nand \U$33707 ( \33960 , \33958 , \33959 );
nor \U$33708 ( \33961 , \33955 , \33960 );
or \U$33709 ( \33962 , \13669 , \33961 );
nand \U$33710 ( \33963 , \15628 , \5494 );
nand \U$33711 ( \33964 , \33962 , \33963 );
and \U$33712 ( \33965 , \33964 , \12195 );
not \U$33713 ( \33966 , \33964 );
and \U$33714 ( \33967 , \33966 , \12956 );
nor \U$33715 ( \33968 , \33965 , \33967 );
nand \U$33716 ( \33969 , \33954 , \33968 );
not \U$33717 ( \33970 , \33969 );
not \U$33718 ( \33971 , RIbe280c0_13);
not \U$33719 ( \33972 , \10936 );
or \U$33720 ( \33973 , \33971 , \33972 );
nand \U$33721 ( \33974 , \14511 , RIbe29830_63);
nand \U$33722 ( \33975 , \33973 , \33974 );
and \U$33723 ( \33976 , \33975 , \17297 );
not \U$33724 ( \33977 , \33975 );
and \U$33725 ( \33978 , \33977 , \13030 );
nor \U$33726 ( \33979 , \33976 , \33978 );
not \U$33727 ( \33980 , \33979 );
or \U$33728 ( \33981 , \33970 , \33980 );
not \U$33729 ( \33982 , \33968 );
nand \U$33730 ( \33983 , \33982 , \33953 );
nand \U$33731 ( \33984 , \33981 , \33983 );
not \U$33732 ( \33985 , \33984 );
or \U$33733 ( \33986 , \33939 , \33985 );
not \U$33734 ( \33987 , \33937 );
not \U$33735 ( \33988 , \33984 );
not \U$33736 ( \33989 , \33988 );
or \U$33737 ( \33990 , \33987 , \33989 );
not \U$33738 ( \33991 , \21013 );
and \U$33739 ( \33992 , \12735 , RIbe27d00_5);
not \U$33740 ( \33993 , \12735 );
and \U$33741 ( \33994 , \12729 , RIbe27d78_6);
and \U$33742 ( \33995 , \33993 , \33994 );
nor \U$33743 ( \33996 , \33992 , \33995 );
not \U$33744 ( \33997 , \33996 );
or \U$33745 ( \33998 , \33991 , \33997 );
or \U$33746 ( \33999 , \33996 , \15166 );
nand \U$33747 ( \34000 , \33998 , \33999 );
and \U$33748 ( \34001 , \12828 , RIbe27c10_3);
or \U$33749 ( \34002 , \12835 , \34001 );
nand \U$33750 ( \34003 , \12835 , \3299 );
nand \U$33751 ( \34004 , \34002 , \34003 );
and \U$33752 ( \34005 , \34004 , \12823 );
not \U$33753 ( \34006 , \34004 );
and \U$33754 ( \34007 , \34006 , \13705 );
nor \U$33755 ( \34008 , \34005 , \34007 );
xor \U$33756 ( \34009 , \34000 , \34008 );
not \U$33757 ( \34010 , RIbe290b0_47);
not \U$33758 ( \34011 , \12707 );
or \U$33759 ( \34012 , \34010 , \34011 );
nand \U$33760 ( \34013 , \12711 , RIbe29a88_68);
nand \U$33761 ( \34014 , \34012 , \34013 );
and \U$33762 ( \34015 , \34014 , \12879 );
not \U$33763 ( \34016 , \34014 );
and \U$33764 ( \34017 , \34016 , \12723 );
nor \U$33765 ( \34018 , \34015 , \34017 );
and \U$33766 ( \34019 , \34009 , \34018 );
and \U$33767 ( \34020 , \34000 , \34008 );
or \U$33768 ( \34021 , \34019 , \34020 );
nand \U$33769 ( \34022 , \33990 , \34021 );
nand \U$33770 ( \34023 , \33986 , \34022 );
nand \U$33771 ( \34024 , \33924 , \34023 );
not \U$33772 ( \34025 , \33805 );
not \U$33773 ( \34026 , \33922 );
nand \U$33774 ( \34027 , \34025 , \34026 );
nand \U$33775 ( \34028 , \34024 , \34027 );
xor \U$33776 ( \34029 , \32283 , \32272 );
xor \U$33777 ( \34030 , \34029 , \32267 );
not \U$33778 ( \34031 , \34030 );
not \U$33779 ( \34032 , \34031 );
xor \U$33780 ( \34033 , \33069 , \33061 );
xnor \U$33781 ( \34034 , \34033 , \33080 );
xor \U$33782 ( \34035 , RIbe2aeb0_111, \12801 );
xor \U$33783 ( \34036 , \34035 , \33031 );
xnor \U$33784 ( \34037 , \34036 , \33046 );
not \U$33785 ( \34038 , \34037 );
and \U$33786 ( \34039 , \34034 , \34038 );
not \U$33787 ( \34040 , \34039 );
or \U$33788 ( \34041 , \34032 , \34040 );
xor \U$33789 ( \34042 , \33011 , \33018 );
xor \U$33790 ( \34043 , \34042 , \33005 );
not \U$33791 ( \34044 , \34043 );
not \U$33792 ( \34045 , \33116 );
not \U$33793 ( \34046 , \33097 );
or \U$33794 ( \34047 , \34045 , \34046 );
or \U$33795 ( \34048 , \33097 , \33116 );
nand \U$33796 ( \34049 , \34047 , \34048 );
not \U$33797 ( \34050 , \33105 );
and \U$33798 ( \34051 , \34049 , \34050 );
not \U$33799 ( \34052 , \34049 );
and \U$33800 ( \34053 , \34052 , \33105 );
nor \U$33801 ( \34054 , \34051 , \34053 );
not \U$33802 ( \34055 , \34054 );
not \U$33803 ( \34056 , \34055 );
or \U$33804 ( \34057 , \34044 , \34056 );
or \U$33805 ( \34058 , \34043 , \34055 );
not \U$33806 ( \34059 , \32955 );
not \U$33807 ( \34060 , \32934 );
not \U$33808 ( \34061 , \34060 );
or \U$33809 ( \34062 , \34059 , \34061 );
nand \U$33810 ( \34063 , \32934 , \32954 );
nand \U$33811 ( \34064 , \34062 , \34063 );
and \U$33812 ( \34065 , \34064 , \32943 );
not \U$33813 ( \34066 , \34064 );
not \U$33814 ( \34067 , \32943 );
and \U$33815 ( \34068 , \34066 , \34067 );
nor \U$33816 ( \34069 , \34065 , \34068 );
nand \U$33817 ( \34070 , \34058 , \34069 );
nand \U$33818 ( \34071 , \34057 , \34070 );
not \U$33819 ( \34072 , \34038 );
not \U$33820 ( \34073 , \34034 );
or \U$33821 ( \34074 , \34072 , \34073 );
nand \U$33822 ( \34075 , \34074 , \34030 );
nand \U$33823 ( \34076 , \34071 , \34075 );
nand \U$33824 ( \34077 , \34041 , \34076 );
xor \U$33825 ( \34078 , \34028 , \34077 );
not \U$33826 ( \34079 , RIbe2aaf0_103);
not \U$33827 ( \34080 , \325 );
or \U$33828 ( \34081 , \34079 , \34080 );
nand \U$33829 ( \34082 , \330 , RIbe2b630_127);
nand \U$33830 ( \34083 , \34081 , \34082 );
not \U$33831 ( \34084 , \34083 );
not \U$33832 ( \34085 , \1374 );
and \U$33833 ( \34086 , \34084 , \34085 );
and \U$33834 ( \34087 , \34083 , \1374 );
nor \U$33835 ( \34088 , \34086 , \34087 );
not \U$33836 ( \34089 , RIbe2b018_114);
not \U$33837 ( \34090 , \30725 );
or \U$33838 ( \34091 , \34089 , \34090 );
nand \U$33839 ( \34092 , \263 , RIbe2afa0_113);
nand \U$33840 ( \34093 , \34091 , \34092 );
not \U$33841 ( \34094 , \34093 );
not \U$33842 ( \34095 , \1362 );
and \U$33843 ( \34096 , \34094 , \34095 );
and \U$33844 ( \34097 , \34093 , \6058 );
nor \U$33845 ( \34098 , \34096 , \34097 );
nand \U$33846 ( \34099 , \34088 , \34098 );
not \U$33847 ( \34100 , \300 );
not \U$33848 ( \34101 , RIbe2af28_112);
not \U$33849 ( \34102 , \6311 );
or \U$33850 ( \34103 , \34101 , \34102 );
nand \U$33851 ( \34104 , \3897 , RIbe2b1f8_118);
nand \U$33852 ( \34105 , \34103 , \34104 );
not \U$33853 ( \34106 , \34105 );
or \U$33854 ( \34107 , \34100 , \34106 );
nand \U$33855 ( \34108 , \3895 , RIbe2af28_112);
nand \U$33856 ( \34109 , \34108 , \34104 , \293 );
nand \U$33857 ( \34110 , \34107 , \34109 );
and \U$33858 ( \34111 , \34099 , \34110 );
nor \U$33859 ( \34112 , \34088 , \34098 );
nor \U$33860 ( \34113 , \34111 , \34112 );
and \U$33861 ( \34114 , \740 , \13156 );
not \U$33862 ( \34115 , \740 );
not \U$33863 ( \34116 , RIbe29308_52);
not \U$33864 ( \34117 , RIbe28c00_37);
or \U$33865 ( \34118 , \34116 , \34117 );
or \U$33866 ( \34119 , RIbe28c00_37, RIbe29308_52);
nand \U$33867 ( \34120 , \34118 , \34119 );
not \U$33868 ( \34121 , \34120 );
nand \U$33869 ( \34122 , \34121 , RIbe2a280_85);
and \U$33870 ( \34123 , \34115 , \34122 );
or \U$33871 ( \34124 , \34114 , \34123 );
not \U$33872 ( \34125 , \34124 );
not \U$33873 ( \34126 , \670 );
and \U$33874 ( \34127 , \34125 , \34126 );
and \U$33875 ( \34128 , \34124 , \670 );
nor \U$33876 ( \34129 , \34127 , \34128 );
not \U$33877 ( \34130 , RIbe2b108_116);
not \U$33878 ( \34131 , \546 );
or \U$33879 ( \34132 , \34130 , \34131 );
nand \U$33880 ( \34133 , \552 , RIbe2b090_115);
nand \U$33881 ( \34134 , \34132 , \34133 );
not \U$33882 ( \34135 , \34134 );
not \U$33883 ( \34136 , \424 );
and \U$33884 ( \34137 , \34135 , \34136 );
and \U$33885 ( \34138 , \34134 , \7124 );
nor \U$33886 ( \34139 , \34137 , \34138 );
and \U$33887 ( \34140 , \34129 , \34139 );
not \U$33888 ( \34141 , \34140 );
not \U$33889 ( \34142 , RIbe2b180_117);
not \U$33890 ( \34143 , \383 );
or \U$33891 ( \34144 , \34142 , \34143 );
nand \U$33892 ( \34145 , \429 , RIbe2b270_119);
nand \U$33893 ( \34146 , \34144 , \34145 );
and \U$33894 ( \34147 , \34146 , \313 );
not \U$33895 ( \34148 , \34146 );
and \U$33896 ( \34149 , \34148 , \306 );
nor \U$33897 ( \34150 , \34147 , \34149 );
not \U$33898 ( \34151 , \34150 );
and \U$33899 ( \34152 , \34141 , \34151 );
nor \U$33900 ( \34153 , \34139 , \34129 );
nor \U$33901 ( \34154 , \34152 , \34153 );
nand \U$33902 ( \34155 , \34113 , \34154 );
not \U$33903 ( \34156 , \34155 );
xor \U$33904 ( \34157 , \32898 , \32907 );
xor \U$33905 ( \34158 , \34157 , \32917 );
not \U$33906 ( \34159 , \34158 );
xor \U$33907 ( \34160 , \32991 , \32978 );
xnor \U$33908 ( \34161 , \34160 , \32968 );
and \U$33909 ( \34162 , \34159 , \34161 );
not \U$33910 ( \34163 , \32864 );
not \U$33911 ( \34164 , \32883 );
or \U$33912 ( \34165 , \34163 , \34164 );
or \U$33913 ( \34166 , \32883 , \32864 );
nand \U$33914 ( \34167 , \34165 , \34166 );
not \U$33915 ( \34168 , \32873 );
and \U$33916 ( \34169 , \34167 , \34168 );
not \U$33917 ( \34170 , \34167 );
and \U$33918 ( \34171 , \34170 , \32873 );
nor \U$33919 ( \34172 , \34169 , \34171 );
nor \U$33920 ( \34173 , \34162 , \34172 );
nor \U$33921 ( \34174 , \34159 , \34161 );
nor \U$33922 ( \34175 , \34173 , \34174 );
not \U$33923 ( \34176 , \34175 );
not \U$33924 ( \34177 , \34176 );
or \U$33925 ( \34178 , \34156 , \34177 );
not \U$33926 ( \34179 , \34155 );
not \U$33927 ( \34180 , \34179 );
not \U$33928 ( \34181 , \34175 );
or \U$33929 ( \34182 , \34180 , \34181 );
xor \U$33930 ( \34183 , \33158 , \33177 );
xor \U$33931 ( \34184 , \34183 , \33180 );
not \U$33932 ( \34185 , \34184 );
xor \U$33933 ( \34186 , \33129 , \33136 );
xor \U$33934 ( \34187 , \34186 , \33144 );
nand \U$33935 ( \34188 , \34185 , \34187 );
not \U$33936 ( \34189 , \34187 );
not \U$33937 ( \34190 , \34189 );
not \U$33938 ( \34191 , \34184 );
or \U$33939 ( \34192 , \34190 , \34191 );
xor \U$33940 ( \34193 , \32837 , \32846 );
xor \U$33941 ( \34194 , \34193 , \32854 );
nand \U$33942 ( \34195 , \34192 , \34194 );
nand \U$33943 ( \34196 , \34188 , \34195 );
nand \U$33944 ( \34197 , \34182 , \34196 );
nand \U$33945 ( \34198 , \34178 , \34197 );
and \U$33946 ( \34199 , \34078 , \34198 );
and \U$33947 ( \34200 , \34028 , \34077 );
or \U$33948 ( \34201 , \34199 , \34200 );
xor \U$33949 ( \34202 , \33237 , \33260 );
xor \U$33950 ( \34203 , \34202 , \33269 );
not \U$33951 ( \34204 , \34203 );
not \U$33952 ( \34205 , \33185 );
not \U$33953 ( \34206 , \33206 );
or \U$33954 ( \34207 , \34205 , \34206 );
nand \U$33955 ( \34208 , \33205 , \33186 );
nand \U$33956 ( \34209 , \34207 , \34208 );
not \U$33957 ( \34210 , \33225 );
and \U$33958 ( \34211 , \34209 , \34210 );
not \U$33959 ( \34212 , \34209 );
and \U$33960 ( \34213 , \34212 , \33225 );
nor \U$33961 ( \34214 , \34211 , \34213 );
not \U$33962 ( \34215 , \34214 );
not \U$33963 ( \34216 , \34215 );
or \U$33964 ( \34217 , \34204 , \34216 );
not \U$33965 ( \34218 , \34214 );
not \U$33966 ( \34219 , \34203 );
not \U$33967 ( \34220 , \34219 );
or \U$33968 ( \34221 , \34218 , \34220 );
xnor \U$33969 ( \34222 , \32484 , \32647 );
xnor \U$33970 ( \34223 , \34222 , \32585 );
nand \U$33971 ( \34224 , \34221 , \34223 );
nand \U$33972 ( \34225 , \34217 , \34224 );
xor \U$33973 ( \34226 , \34201 , \34225 );
xor \U$33974 ( \34227 , \33147 , \33149 );
xor \U$33975 ( \34228 , \34227 , \33182 );
not \U$33976 ( \34229 , \33021 );
xor \U$33977 ( \34230 , \32993 , \32958 );
not \U$33978 ( \34231 , \34230 );
or \U$33979 ( \34232 , \34229 , \34231 );
or \U$33980 ( \34233 , \33021 , \34230 );
nand \U$33981 ( \34234 , \34232 , \34233 );
xor \U$33982 ( \34235 , \34228 , \34234 );
xor \U$33983 ( \34236 , \32857 , \32887 );
xor \U$33984 ( \34237 , \34236 , \32920 );
and \U$33985 ( \34238 , \34235 , \34237 );
and \U$33986 ( \34239 , \34228 , \34234 );
or \U$33987 ( \34240 , \34238 , \34239 );
xor \U$33988 ( \34241 , \33210 , \33212 );
xor \U$33989 ( \34242 , \34241 , \33222 );
not \U$33990 ( \34243 , \33196 );
not \U$33991 ( \34244 , \33200 );
or \U$33992 ( \34245 , \34243 , \34244 );
or \U$33993 ( \34246 , \33200 , \33196 );
nand \U$33994 ( \34247 , \34245 , \34246 );
and \U$33995 ( \34248 , \34247 , \33203 );
not \U$33996 ( \34249 , \34247 );
and \U$33997 ( \34250 , \34249 , \33193 );
nor \U$33998 ( \34251 , \34248 , \34250 );
xor \U$33999 ( \34252 , \34242 , \34251 );
not \U$34000 ( \34253 , \33244 );
xor \U$34001 ( \34254 , \33257 , \34253 );
xnor \U$34002 ( \34255 , \34254 , \33246 );
and \U$34003 ( \34256 , \34252 , \34255 );
and \U$34004 ( \34257 , \34242 , \34251 );
or \U$34005 ( \34258 , \34256 , \34257 );
xor \U$34006 ( \34259 , \34240 , \34258 );
xnor \U$34007 ( \34260 , \32322 , \32425 );
and \U$34008 ( \34261 , \34260 , \32428 );
not \U$34009 ( \34262 , \34260 );
and \U$34010 ( \34263 , \34262 , \32228 );
nor \U$34011 ( \34264 , \34261 , \34263 );
and \U$34012 ( \34265 , \34259 , \34264 );
and \U$34013 ( \34266 , \34240 , \34258 );
or \U$34014 ( \34267 , \34265 , \34266 );
and \U$34015 ( \34268 , \34226 , \34267 );
and \U$34016 ( \34269 , \34201 , \34225 );
or \U$34017 ( \34270 , \34268 , \34269 );
xor \U$34018 ( \34271 , \33698 , \34270 );
and \U$34019 ( \34272 , \33678 , \33683 );
not \U$34020 ( \34273 , \33678 );
and \U$34021 ( \34274 , \34273 , \33694 );
nor \U$34022 ( \34275 , \34272 , \34274 );
xnor \U$34023 ( \34276 , \34275 , \33691 );
not \U$34024 ( \34277 , \32431 );
not \U$34025 ( \34278 , \32826 );
or \U$34026 ( \34279 , \34277 , \34278 );
nand \U$34027 ( \34280 , \32430 , \32650 );
nand \U$34028 ( \34281 , \34279 , \34280 );
xnor \U$34029 ( \34282 , \34281 , \32823 );
xor \U$34030 ( \34283 , \34276 , \34282 );
not \U$34031 ( \34284 , \33292 );
not \U$34032 ( \34285 , \33427 );
or \U$34033 ( \34286 , \34284 , \34285 );
or \U$34034 ( \34287 , \33427 , \33292 );
nand \U$34035 ( \34288 , \34286 , \34287 );
xnor \U$34036 ( \34289 , \33659 , \34288 );
and \U$34037 ( \34290 , \34283 , \34289 );
and \U$34038 ( \34291 , \34276 , \34282 );
or \U$34039 ( \34292 , \34290 , \34291 );
xnor \U$34040 ( \34293 , \34271 , \34292 );
and \U$34041 ( \34294 , \33664 , \34293 );
xor \U$34042 ( \34295 , \32810 , \32816 );
and \U$34043 ( \34296 , \34295 , \32821 );
and \U$34044 ( \34297 , \32810 , \32816 );
or \U$34045 ( \34298 , \34296 , \34297 );
not \U$34046 ( \34299 , \34298 );
not \U$34047 ( \34300 , \34299 );
xor \U$34048 ( \34301 , \32740 , \32772 );
and \U$34049 ( \34302 , \34301 , \32804 );
and \U$34050 ( \34303 , \32740 , \32772 );
or \U$34051 ( \34304 , \34302 , \34303 );
xor \U$34052 ( \34305 , \32675 , \32704 );
and \U$34053 ( \34306 , \34305 , \32735 );
and \U$34054 ( \34307 , \32675 , \32704 );
or \U$34055 ( \34308 , \34306 , \34307 );
and \U$34056 ( \34309 , \34304 , \34308 );
not \U$34057 ( \34310 , \34304 );
not \U$34058 ( \34311 , \34308 );
and \U$34059 ( \34312 , \34310 , \34311 );
nor \U$34060 ( \34313 , \34309 , \34312 );
not \U$34061 ( \34314 , \34313 );
or \U$34062 ( \34315 , \34300 , \34314 );
or \U$34063 ( \34316 , \34313 , \34299 );
nand \U$34064 ( \34317 , \34315 , \34316 );
or \U$34065 ( \34318 , \32736 , \32822 );
nand \U$34066 ( \34319 , \34318 , \32805 );
nand \U$34067 ( \34320 , \32736 , \32822 );
nand \U$34068 ( \34321 , \34319 , \34320 );
or \U$34069 ( \34322 , \33658 , \33469 );
nand \U$34070 ( \34323 , \34322 , \33567 );
nand \U$34071 ( \34324 , \33658 , \33469 );
nand \U$34072 ( \34325 , \34323 , \34324 );
xor \U$34073 ( \34326 , \34321 , \34325 );
or \U$34074 ( \34327 , \33637 , \33646 );
nand \U$34075 ( \34328 , \34327 , \33656 );
nand \U$34076 ( \34329 , \33646 , \33637 );
nand \U$34077 ( \34330 , \34328 , \34329 );
xor \U$34078 ( \34331 , \33576 , \33585 );
and \U$34079 ( \34332 , \34331 , \33595 );
and \U$34080 ( \34333 , \33576 , \33585 );
or \U$34081 ( \34334 , \34332 , \34333 );
xor \U$34082 ( \34335 , \34330 , \34334 );
xor \U$34083 ( \34336 , \33607 , \33616 );
and \U$34084 ( \34337 , \34336 , \33626 );
and \U$34085 ( \34338 , \33607 , \33616 );
or \U$34086 ( \34339 , \34337 , \34338 );
xor \U$34087 ( \34340 , \34335 , \34339 );
not \U$34088 ( \34341 , \33326 );
not \U$34089 ( \34342 , \33318 );
or \U$34090 ( \34343 , \34341 , \34342 );
nand \U$34091 ( \34344 , \34343 , \33308 );
nand \U$34092 ( \34345 , \33330 , \33327 );
nand \U$34093 ( \34346 , \34344 , \34345 );
not \U$34094 ( \34347 , \34346 );
not \U$34095 ( \34348 , \34347 );
and \U$34096 ( \34349 , \33372 , \33361 );
nor \U$34097 ( \34350 , \34349 , \33348 );
nor \U$34098 ( \34351 , \33372 , \33361 );
nor \U$34099 ( \34352 , \34350 , \34351 );
not \U$34100 ( \34353 , \34352 );
not \U$34101 ( \34354 , \34353 );
or \U$34102 ( \34355 , \34348 , \34354 );
nand \U$34103 ( \34356 , \34346 , \34352 );
nand \U$34104 ( \34357 , \34355 , \34356 );
not \U$34105 ( \34358 , \33392 );
not \U$34106 ( \34359 , \33419 );
or \U$34107 ( \34360 , \34358 , \34359 );
not \U$34108 ( \34361 , \33393 );
not \U$34109 ( \34362 , \33415 );
or \U$34110 ( \34363 , \34361 , \34362 );
nand \U$34111 ( \34364 , \34363 , \33401 );
nand \U$34112 ( \34365 , \34360 , \34364 );
not \U$34113 ( \34366 , \34365 );
and \U$34114 ( \34367 , \34357 , \34366 );
not \U$34115 ( \34368 , \34357 );
and \U$34116 ( \34369 , \34368 , \34365 );
nor \U$34117 ( \34370 , \34367 , \34369 );
xor \U$34118 ( \34371 , \34340 , \34370 );
and \U$34119 ( \34372 , \33548 , \33560 );
nor \U$34120 ( \34373 , \34372 , \33536 );
nor \U$34121 ( \34374 , \33548 , \33560 );
nor \U$34122 ( \34375 , \34373 , \34374 );
buf \U$34123 ( \34376 , \33479 );
and \U$34124 ( \34377 , \33499 , \34376 );
nor \U$34125 ( \34378 , \34377 , \33489 );
nor \U$34126 ( \34379 , \33499 , \34376 );
nor \U$34127 ( \34380 , \34378 , \34379 );
xor \U$34128 ( \34381 , \34375 , \34380 );
not \U$34129 ( \34382 , \33518 );
and \U$34130 ( \34383 , \33526 , \34382 );
nor \U$34131 ( \34384 , \34383 , \33509 );
nor \U$34132 ( \34385 , \33526 , \34382 );
nor \U$34133 ( \34386 , \34384 , \34385 );
xor \U$34134 ( \34387 , \34381 , \34386 );
and \U$34135 ( \34388 , \34371 , \34387 );
not \U$34136 ( \34389 , \34371 );
not \U$34137 ( \34390 , \34387 );
and \U$34138 ( \34391 , \34389 , \34390 );
nor \U$34139 ( \34392 , \34388 , \34391 );
xor \U$34140 ( \34393 , \34326 , \34392 );
xor \U$34141 ( \34394 , \34317 , \34393 );
not \U$34142 ( \34395 , RIbe27f58_10);
not \U$34143 ( \34396 , \7880 );
or \U$34144 ( \34397 , \34395 , \34396 );
nand \U$34145 ( \34398 , \6787 , RIbe27e68_8);
nand \U$34146 ( \34399 , \34397 , \34398 );
and \U$34147 ( \34400 , \34399 , \3471 );
not \U$34148 ( \34401 , \34399 );
and \U$34149 ( \34402 , \34401 , \3448 );
nor \U$34150 ( \34403 , \34400 , \34402 );
not \U$34151 ( \34404 , \34403 );
not \U$34152 ( \34405 , RIbe28660_25);
not \U$34153 ( \34406 , \6413 );
or \U$34154 ( \34407 , \34405 , \34406 );
nand \U$34155 ( \34408 , \21043 , RIbe285e8_24);
nand \U$34156 ( \34409 , \34407 , \34408 );
not \U$34157 ( \34410 , \34409 );
not \U$34158 ( \34411 , \4323 );
and \U$34159 ( \34412 , \34410 , \34411 );
and \U$34160 ( \34413 , \34409 , \7865 );
nor \U$34161 ( \34414 , \34412 , \34413 );
not \U$34162 ( \34415 , \34414 );
or \U$34163 ( \34416 , \34404 , \34415 );
or \U$34164 ( \34417 , \34414 , \34403 );
nand \U$34165 ( \34418 , \34416 , \34417 );
not \U$34166 ( \34419 , RIbe28ed0_43);
not \U$34167 ( \34420 , \3451 );
or \U$34168 ( \34421 , \34419 , \34420 );
nand \U$34169 ( \34422 , \4011 , RIbe27fd0_11);
nand \U$34170 ( \34423 , \34421 , \34422 );
not \U$34171 ( \34424 , \34423 );
not \U$34172 ( \34425 , \2887 );
and \U$34173 ( \34426 , \34424 , \34425 );
and \U$34174 ( \34427 , \34423 , \2887 );
nor \U$34175 ( \34428 , \34426 , \34427 );
and \U$34176 ( \34429 , \34418 , \34428 );
not \U$34177 ( \34430 , \34418 );
not \U$34178 ( \34431 , \34428 );
and \U$34179 ( \34432 , \34430 , \34431 );
nor \U$34180 ( \34433 , \34429 , \34432 );
not \U$34181 ( \34434 , RIbe28b10_35);
not \U$34182 ( \34435 , \6138 );
or \U$34183 ( \34436 , \34434 , \34435 );
nand \U$34184 ( \34437 , \6616 , RIbe28b88_36);
nand \U$34185 ( \34438 , \34436 , \34437 );
and \U$34186 ( \34439 , \34438 , \7535 );
not \U$34187 ( \34440 , \34438 );
and \U$34188 ( \34441 , \34440 , \6623 );
nor \U$34189 ( \34442 , \34439 , \34441 );
not \U$34190 ( \34443 , \34442 );
not \U$34191 ( \34444 , RIbe28408_20);
not \U$34192 ( \34445 , \5455 );
or \U$34193 ( \34446 , \34444 , \34445 );
nand \U$34194 ( \34447 , \6634 , RIbe28390_19);
nand \U$34195 ( \34448 , \34446 , \34447 );
not \U$34196 ( \34449 , \34448 );
not \U$34197 ( \34450 , \6641 );
and \U$34198 ( \34451 , \34449 , \34450 );
and \U$34199 ( \34452 , \34448 , \6118 );
nor \U$34200 ( \34453 , \34451 , \34452 );
not \U$34201 ( \34454 , \34453 );
not \U$34202 ( \34455 , \34454 );
or \U$34203 ( \34456 , \34443 , \34455 );
not \U$34204 ( \34457 , \34442 );
nand \U$34205 ( \34458 , \34457 , \34453 );
nand \U$34206 ( \34459 , \34456 , \34458 );
not \U$34207 ( \34460 , RIbe287c8_28);
not \U$34208 ( \34461 , \4829 );
or \U$34209 ( \34462 , \34460 , \34461 );
nand \U$34210 ( \34463 , \5052 , RIbe28480_21);
nand \U$34211 ( \34464 , \34462 , \34463 );
and \U$34212 ( \34465 , \34464 , \4946 );
not \U$34213 ( \34466 , \34464 );
and \U$34214 ( \34467 , \34466 , \4586 );
nor \U$34215 ( \34468 , \34465 , \34467 );
xor \U$34216 ( \34469 , \34459 , \34468 );
xor \U$34217 ( \34470 , \34433 , \34469 );
not \U$34218 ( \34471 , \2889 );
not \U$34219 ( \34472 , \9801 );
and \U$34220 ( \34473 , \34471 , \34472 );
and \U$34221 ( \34474 , \8833 , RIbe29dd0_75);
nor \U$34222 ( \34475 , \34473 , \34474 );
and \U$34223 ( \34476 , \34475 , \3516 );
not \U$34224 ( \34477 , \34475 );
and \U$34225 ( \34478 , \34477 , \1277 );
nor \U$34226 ( \34479 , \34476 , \34478 );
not \U$34227 ( \34480 , RIbe29bf0_71);
not \U$34228 ( \34481 , \2898 );
or \U$34229 ( \34482 , \34480 , \34481 );
nand \U$34230 ( \34483 , \4284 , RIbe28f48_44);
nand \U$34231 ( \34484 , \34482 , \34483 );
and \U$34232 ( \34485 , \34484 , \2379 );
not \U$34233 ( \34486 , \34484 );
and \U$34234 ( \34487 , \34486 , \7457 );
nor \U$34235 ( \34488 , \34485 , \34487 );
and \U$34236 ( \34489 , \34479 , \34488 );
not \U$34237 ( \34490 , \34479 );
not \U$34238 ( \34491 , \34488 );
and \U$34239 ( \34492 , \34490 , \34491 );
or \U$34240 ( \34493 , \34489 , \34492 );
and \U$34241 ( \34494 , \1112 , RIbe29fb0_79);
and \U$34242 ( \34495 , \1117 , RIbe29e48_76);
nor \U$34243 ( \34496 , \34494 , \34495 );
and \U$34244 ( \34497 , \34496 , \1132 );
not \U$34245 ( \34498 , \34496 );
and \U$34246 ( \34499 , \34498 , \1125 );
nor \U$34247 ( \34500 , \34497 , \34499 );
and \U$34248 ( \34501 , \34493 , \34500 );
not \U$34249 ( \34502 , \34493 );
not \U$34250 ( \34503 , \34500 );
and \U$34251 ( \34504 , \34502 , \34503 );
nor \U$34252 ( \34505 , \34501 , \34504 );
xor \U$34253 ( \34506 , \34470 , \34505 );
nand \U$34254 ( \34507 , RIbe29380_53, RIbe2af28_112);
xor \U$34255 ( \34508 , \34507 , \33431 );
nand \U$34256 ( \34509 , \33452 , \33445 );
and \U$34257 ( \34510 , \34509 , \33460 );
nor \U$34258 ( \34511 , \33445 , \33452 );
nor \U$34259 ( \34512 , \34510 , \34511 );
xor \U$34260 ( \34513 , \34508 , \34512 );
xor \U$34261 ( \34514 , \34506 , \34513 );
not \U$34262 ( \34515 , RIbe2b270_119);
not \U$34263 ( \34516 , \260 );
or \U$34264 ( \34517 , \34515 , \34516 );
nand \U$34265 ( \34518 , \263 , RIbe2b108_116);
nand \U$34266 ( \34519 , \34517 , \34518 );
not \U$34267 ( \34520 , \34519 );
not \U$34268 ( \34521 , \1361 );
and \U$34269 ( \34522 , \34520 , \34521 );
and \U$34270 ( \34523 , \34519 , \6058 );
nor \U$34271 ( \34524 , \34522 , \34523 );
not \U$34272 ( \34525 , RIbe2b090_115);
not \U$34273 ( \34526 , \1252 );
or \U$34274 ( \34527 , \34525 , \34526 );
nand \U$34275 ( \34528 , \9816 , RIbe2a280_85);
nand \U$34276 ( \34529 , \34527 , \34528 );
and \U$34277 ( \34530 , \34529 , \293 );
not \U$34278 ( \34531 , \34529 );
and \U$34279 ( \34532 , \34531 , \300 );
nor \U$34280 ( \34533 , \34530 , \34532 );
xor \U$34281 ( \34534 , \34524 , \34533 );
not \U$34282 ( \34535 , RIbe2b1f8_118);
not \U$34283 ( \34536 , \325 );
or \U$34284 ( \34537 , \34535 , \34536 );
not \U$34285 ( \34538 , \14248 );
nand \U$34286 ( \34539 , \34538 , \329 );
nand \U$34287 ( \34540 , \34537 , \34539 );
and \U$34288 ( \34541 , \34540 , \4172 );
not \U$34289 ( \34542 , \34540 );
and \U$34290 ( \34543 , \34542 , \1375 );
nor \U$34291 ( \34544 , \34541 , \34543 );
xor \U$34292 ( \34545 , \34534 , \34544 );
not \U$34293 ( \34546 , RIbe2a370_87);
not \U$34294 ( \34547 , \2597 );
or \U$34295 ( \34548 , \34546 , \34547 );
nand \U$34296 ( \34549 , \1146 , RIbe2a2f8_86);
nand \U$34297 ( \34550 , \34548 , \34549 );
not \U$34298 ( \34551 , \34550 );
not \U$34299 ( \34552 , \1153 );
and \U$34300 ( \34553 , \34551 , \34552 );
and \U$34301 ( \34554 , \34550 , \3994 );
nor \U$34302 ( \34555 , \34553 , \34554 );
not \U$34303 ( \34556 , RIbe2acd0_107);
not \U$34304 ( \34557 , \1632 );
or \U$34305 ( \34558 , \34556 , \34557 );
nand \U$34306 ( \34559 , \1099 , RIbe2a028_80);
nand \U$34307 ( \34560 , \34558 , \34559 );
and \U$34308 ( \34561 , \34560 , \1309 );
not \U$34309 ( \34562 , \34560 );
and \U$34310 ( \34563 , \34562 , \5125 );
nor \U$34311 ( \34564 , \34561 , \34563 );
xnor \U$34312 ( \34565 , \34555 , \34564 );
not \U$34313 ( \34566 , RIbe2b5b8_126);
not \U$34314 ( \34567 , \1003 );
or \U$34315 ( \34568 , \34566 , \34567 );
nand \U$34316 ( \34569 , \7905 , RIbe2a3e8_88);
nand \U$34317 ( \34570 , \34568 , \34569 );
and \U$34318 ( \34571 , \34570 , \1608 );
not \U$34319 ( \34572 , \34570 );
and \U$34320 ( \34573 , \34572 , \1011 );
nor \U$34321 ( \34574 , \34571 , \34573 );
xnor \U$34322 ( \34575 , \34565 , \34574 );
xor \U$34323 ( \34576 , \34545 , \34575 );
not \U$34324 ( \34577 , RIbe2a208_84);
not \U$34325 ( \34578 , \1337 );
or \U$34326 ( \34579 , \34577 , \34578 );
not \U$34327 ( \34580 , \14285 );
nand \U$34328 ( \34581 , \34580 , \429 );
nand \U$34329 ( \34582 , \34579 , \34581 );
and \U$34330 ( \34583 , \34582 , \313 );
not \U$34331 ( \34584 , \34582 );
and \U$34332 ( \34585 , \34584 , \306 );
nor \U$34333 ( \34586 , \34583 , \34585 );
not \U$34334 ( \34587 , RIbe2a988_100);
not \U$34335 ( \34588 , \664 );
or \U$34336 ( \34589 , \34587 , \34588 );
nand \U$34337 ( \34590 , RIbe2a910_99, \1180 );
nand \U$34338 ( \34591 , \34589 , \34590 );
xor \U$34339 ( \34592 , \34591 , \564 );
xor \U$34340 ( \34593 , \34586 , \34592 );
and \U$34341 ( \34594 , \1756 , RIbe2a5c8_92);
and \U$34342 ( \34595 , \552 , RIbe2a550_91);
nor \U$34343 ( \34596 , \34594 , \34595 );
and \U$34344 ( \34597 , \34596 , \1764 );
not \U$34345 ( \34598 , \34596 );
and \U$34346 ( \34599 , \34598 , \1245 );
nor \U$34347 ( \34600 , \34597 , \34599 );
xor \U$34348 ( \34601 , \34593 , \34600 );
xor \U$34349 ( \34602 , \34576 , \34601 );
xor \U$34350 ( \34603 , \34514 , \34602 );
not \U$34351 ( \34604 , \34603 );
not \U$34352 ( \34605 , RIbe28e58_42);
not \U$34353 ( \34606 , \15573 );
or \U$34354 ( \34607 , \34605 , \34606 );
not \U$34355 ( \34608 , \2890 );
nand \U$34356 ( \34609 , \34608 , \12711 );
nand \U$34357 ( \34610 , \34607 , \34609 );
and \U$34358 ( \34611 , \34610 , \12723 );
not \U$34359 ( \34612 , \34610 );
and \U$34360 ( \34613 , \34612 , \12716 );
nor \U$34361 ( \34614 , \34611 , \34613 );
not \U$34362 ( \34615 , \34614 );
and \U$34363 ( \34616 , \12729 , RIbe29920_65);
or \U$34364 ( \34617 , \14074 , \34616 );
nand \U$34365 ( \34618 , \13077 , \1640 );
nand \U$34366 ( \34619 , \34617 , \34618 );
and \U$34367 ( \34620 , \34619 , \12746 );
not \U$34368 ( \34621 , \34619 );
and \U$34369 ( \34622 , \34621 , \12743 );
nor \U$34370 ( \34623 , \34620 , \34622 );
and \U$34371 ( \34624 , \34623 , \19783 );
not \U$34372 ( \34625 , \34623 );
and \U$34373 ( \34626 , \34625 , \13595 );
nor \U$34374 ( \34627 , \34624 , \34626 );
xor \U$34375 ( \34628 , \34615 , \34627 );
not \U$34376 ( \34629 , \33338 );
not \U$34377 ( \34630 , \33421 );
or \U$34378 ( \34631 , \34629 , \34630 );
nand \U$34379 ( \34632 , \33377 , \33406 , \33419 );
nand \U$34380 ( \34633 , \33377 , \33332 , \33336 );
nand \U$34381 ( \34634 , \34632 , \34633 );
nand \U$34382 ( \34635 , \33377 , \33405 , \33416 );
nand \U$34383 ( \34636 , \33377 , \33333 , \33308 );
nand \U$34384 ( \34637 , \34635 , \34636 );
nor \U$34385 ( \34638 , \34634 , \34637 );
nand \U$34386 ( \34639 , \34631 , \34638 );
xor \U$34387 ( \34640 , \34628 , \34639 );
and \U$34388 ( \34641 , \13092 , RIbe27d00_5);
and \U$34389 ( \34642 , \13086 , RIbe27c10_3);
nor \U$34390 ( \34643 , \34641 , \34642 );
and \U$34391 ( \34644 , \34643 , \12927 );
not \U$34392 ( \34645 , \34643 );
and \U$34393 ( \34646 , \34645 , \12770 );
nor \U$34394 ( \34647 , \34644 , \34646 );
not \U$34395 ( \34648 , \34647 );
and \U$34396 ( \34649 , \15205 , RIbe29a88_68);
not \U$34397 ( \34650 , \12947 );
nor \U$34398 ( \34651 , \34650 , \255 );
nor \U$34399 ( \34652 , \34649 , \34651 );
and \U$34400 ( \34653 , \34652 , \17005 );
not \U$34401 ( \34654 , \34652 );
and \U$34402 ( \34655 , \34654 , \12195 );
nor \U$34403 ( \34656 , \34653 , \34655 );
not \U$34404 ( \34657 , \34656 );
or \U$34405 ( \34658 , \34648 , \34657 );
or \U$34406 ( \34659 , \34647 , \34656 );
nand \U$34407 ( \34660 , \34658 , \34659 );
not \U$34408 ( \34661 , RIbe28fc0_45);
not \U$34409 ( \34662 , \10936 );
or \U$34410 ( \34663 , \34661 , \34662 );
nand \U$34411 ( \34664 , \12213 , RIbe290b0_47);
nand \U$34412 ( \34665 , \34663 , \34664 );
not \U$34413 ( \34666 , \34665 );
not \U$34414 ( \34667 , \13030 );
and \U$34415 ( \34668 , \34666 , \34667 );
and \U$34416 ( \34669 , \34665 , \13661 );
nor \U$34417 ( \34670 , \34668 , \34669 );
not \U$34418 ( \34671 , \34670 );
and \U$34419 ( \34672 , \34660 , \34671 );
not \U$34420 ( \34673 , \34660 );
and \U$34421 ( \34674 , \34673 , \34670 );
nor \U$34422 ( \34675 , \34672 , \34674 );
not \U$34423 ( \34676 , \34675 );
not \U$34424 ( \34677 , RIbe29830_63);
not \U$34425 ( \34678 , \6942 );
or \U$34426 ( \34679 , \34677 , \34678 );
nand \U$34427 ( \34680 , \13158 , RIbe296c8_60);
nand \U$34428 ( \34681 , \34679 , \34680 );
and \U$34429 ( \34682 , \34681 , \6948 );
not \U$34430 ( \34683 , \34681 );
and \U$34431 ( \34684 , \34683 , \6950 );
nor \U$34432 ( \34685 , \34682 , \34684 );
not \U$34433 ( \34686 , \34685 );
not \U$34434 ( \34687 , \34686 );
and \U$34435 ( \34688 , \10915 , RIbe29650_59);
and \U$34436 ( \34689 , \13038 , RIbe29038_46);
nor \U$34437 ( \34690 , \34688 , \34689 );
and \U$34438 ( \34691 , \34690 , \13383 );
not \U$34439 ( \34692 , \34690 );
and \U$34440 ( \34693 , \34692 , \16994 );
nor \U$34441 ( \34694 , \34691 , \34693 );
not \U$34442 ( \34695 , \34694 );
not \U$34443 ( \34696 , \34695 );
or \U$34444 ( \34697 , \34687 , \34696 );
nand \U$34445 ( \34698 , \34694 , \34685 );
nand \U$34446 ( \34699 , \34697 , \34698 );
not \U$34447 ( \34700 , RIbe281b0_15);
not \U$34448 ( \34701 , \7298 );
or \U$34449 ( \34702 , \34700 , \34701 );
nand \U$34450 ( \34703 , \13792 , RIbe280c0_13);
nand \U$34451 ( \34704 , \34702 , \34703 );
and \U$34452 ( \34705 , \34704 , \7304 );
not \U$34453 ( \34706 , \34704 );
and \U$34454 ( \34707 , \34706 , \6992 );
nor \U$34455 ( \34708 , \34705 , \34707 );
xnor \U$34456 ( \34709 , \34699 , \34708 );
not \U$34457 ( \34710 , \34709 );
or \U$34458 ( \34711 , \34676 , \34710 );
or \U$34459 ( \34712 , \34675 , \34709 );
nand \U$34460 ( \34713 , \34711 , \34712 );
not \U$34461 ( \34714 , RIbe29560_57);
not \U$34462 ( \34715 , \13327 );
or \U$34463 ( \34716 , \34714 , \34715 );
not \U$34464 ( \34717 , \3952 );
nand \U$34465 ( \34718 , \34717 , \7958 );
nand \U$34466 ( \34719 , \34716 , \34718 );
and \U$34467 ( \34720 , \34719 , \6572 );
not \U$34468 ( \34721 , \34719 );
and \U$34469 ( \34722 , \34721 , \7293 );
nor \U$34470 ( \34723 , \34720 , \34722 );
not \U$34471 ( \34724 , RIbe289a8_32);
not \U$34472 ( \34725 , \7941 );
or \U$34473 ( \34726 , \34724 , \34725 );
nand \U$34474 ( \34727 , RIbe28930_31, \6596 );
nand \U$34475 ( \34728 , \34726 , \34727 );
and \U$34476 ( \34729 , \34728 , \13956 );
not \U$34477 ( \34730 , \34728 );
and \U$34478 ( \34731 , \34730 , \7948 );
nor \U$34479 ( \34732 , \34729 , \34731 );
not \U$34480 ( \34733 , \34732 );
xor \U$34481 ( \34734 , \34723 , \34733 );
not \U$34482 ( \34735 , RIbe29290_51);
not \U$34483 ( \34736 , \6536 );
or \U$34484 ( \34737 , \34735 , \34736 );
nand \U$34485 ( \34738 , \7076 , RIbe28a20_33);
nand \U$34486 ( \34739 , \34737 , \34738 );
xnor \U$34487 ( \34740 , \34739 , \6891 );
xor \U$34488 ( \34741 , \34734 , \34740 );
not \U$34489 ( \34742 , \34741 );
and \U$34490 ( \34743 , \34713 , \34742 );
not \U$34491 ( \34744 , \34713 );
and \U$34492 ( \34745 , \34744 , \34741 );
nor \U$34493 ( \34746 , \34743 , \34745 );
xnor \U$34494 ( \34747 , \34640 , \34746 );
not \U$34495 ( \34748 , \34747 );
xor \U$34496 ( \34749 , \33431 , \33435 );
and \U$34497 ( \34750 , \34749 , \33468 );
and \U$34498 ( \34751 , \33431 , \33435 );
or \U$34499 ( \34752 , \34750 , \34751 );
not \U$34500 ( \34753 , \33500 );
not \U$34501 ( \34754 , \33564 );
or \U$34502 ( \34755 , \34753 , \34754 );
or \U$34503 ( \34756 , \33564 , \33500 );
nand \U$34504 ( \34757 , \34756 , \33527 );
nand \U$34505 ( \34758 , \34755 , \34757 );
xor \U$34506 ( \34759 , \34752 , \34758 );
xor \U$34507 ( \34760 , \33596 , \33627 );
and \U$34508 ( \34761 , \34760 , \33657 );
and \U$34509 ( \34762 , \33596 , \33627 );
or \U$34510 ( \34763 , \34761 , \34762 );
xor \U$34511 ( \34764 , \34759 , \34763 );
not \U$34512 ( \34765 , \34764 );
and \U$34513 ( \34766 , \34748 , \34765 );
and \U$34514 ( \34767 , \34747 , \34764 );
nor \U$34515 ( \34768 , \34766 , \34767 );
not \U$34516 ( \34769 , \34768 );
or \U$34517 ( \34770 , \34604 , \34769 );
or \U$34518 ( \34771 , \34603 , \34768 );
nand \U$34519 ( \34772 , \34770 , \34771 );
xor \U$34520 ( \34773 , \34394 , \34772 );
and \U$34521 ( \34774 , \34021 , \33984 );
not \U$34522 ( \34775 , \34021 );
and \U$34523 ( \34776 , \34775 , \33988 );
nor \U$34524 ( \34777 , \34774 , \34776 );
and \U$34525 ( \34778 , \34777 , \33937 );
not \U$34526 ( \34779 , \34777 );
and \U$34527 ( \34780 , \34779 , \33938 );
nor \U$34528 ( \34781 , \34778 , \34780 );
xor \U$34529 ( \34782 , \33873 , \33917 );
nand \U$34530 ( \34783 , \33837 , \33836 );
nand \U$34531 ( \34784 , \33835 , \34783 );
xnor \U$34532 ( \34785 , \34782 , \34784 );
not \U$34533 ( \34786 , \34785 );
nand \U$34534 ( \34787 , \34781 , \34786 );
xor \U$34535 ( \34788 , \33769 , \33730 );
xor \U$34536 ( \34789 , \34788 , \33802 );
and \U$34537 ( \34790 , \34787 , \34789 );
nor \U$34538 ( \34791 , \34781 , \34786 );
nor \U$34539 ( \34792 , \34790 , \34791 );
and \U$34540 ( \34793 , \33119 , \33085 );
not \U$34541 ( \34794 , \33119 );
and \U$34542 ( \34795 , \34794 , \33084 );
or \U$34543 ( \34796 , \34793 , \34795 );
xor \U$34544 ( \34797 , \34796 , \33051 );
or \U$34545 ( \34798 , \34792 , \34797 );
not \U$34546 ( \34799 , \34797 );
not \U$34547 ( \34800 , \34792 );
or \U$34548 ( \34801 , \34799 , \34800 );
xor \U$34549 ( \34802 , \34172 , \34158 );
and \U$34550 ( \34803 , \34802 , \34161 );
not \U$34551 ( \34804 , \34802 );
not \U$34552 ( \34805 , \34161 );
and \U$34553 ( \34806 , \34804 , \34805 );
nor \U$34554 ( \34807 , \34803 , \34806 );
not \U$34555 ( \34808 , \34807 );
or \U$34556 ( \34809 , \34113 , \34154 );
nand \U$34557 ( \34810 , \34809 , \34155 );
not \U$34558 ( \34811 , \34810 );
not \U$34559 ( \34812 , \34184 );
not \U$34560 ( \34813 , \34194 );
or \U$34561 ( \34814 , \34812 , \34813 );
or \U$34562 ( \34815 , \34184 , \34194 );
nand \U$34563 ( \34816 , \34814 , \34815 );
and \U$34564 ( \34817 , \34816 , \34189 );
not \U$34565 ( \34818 , \34816 );
and \U$34566 ( \34819 , \34818 , \34187 );
nor \U$34567 ( \34820 , \34817 , \34819 );
nand \U$34568 ( \34821 , \34811 , \34820 );
not \U$34569 ( \34822 , \34821 );
or \U$34570 ( \34823 , \34808 , \34822 );
not \U$34571 ( \34824 , \34820 );
nand \U$34572 ( \34825 , \34824 , \34810 );
nand \U$34573 ( \34826 , \34823 , \34825 );
nand \U$34574 ( \34827 , \34801 , \34826 );
nand \U$34575 ( \34828 , \34798 , \34827 );
not \U$34576 ( \34829 , \34828 );
and \U$34577 ( \34830 , \1161 , RIbe2a208_84);
and \U$34578 ( \34831 , \7905 , RIbe2a190_83);
nor \U$34579 ( \34832 , \34830 , \34831 );
and \U$34580 ( \34833 , \34832 , \1011 );
not \U$34581 ( \34834 , \34832 );
and \U$34582 ( \34835 , \34834 , \1813 );
nor \U$34583 ( \34836 , \34833 , \34835 );
not \U$34584 ( \34837 , RIbe2a5c8_92);
not \U$34585 ( \34838 , \1143 );
or \U$34586 ( \34839 , \34837 , \34838 );
not \U$34587 ( \34840 , \21491 );
nand \U$34588 ( \34841 , \34840 , \1147 );
nand \U$34589 ( \34842 , \34839 , \34841 );
and \U$34590 ( \34843 , \34842 , \1153 );
not \U$34591 ( \34844 , \34842 );
and \U$34592 ( \34845 , \34844 , \1154 );
nor \U$34593 ( \34846 , \34843 , \34845 );
and \U$34594 ( \34847 , \34836 , \34846 );
not \U$34595 ( \34848 , RIbe2b090_115);
not \U$34596 ( \34849 , \6350 );
or \U$34597 ( \34850 , \34848 , \34849 );
nand \U$34598 ( \34851 , \1180 , RIbe2a280_85);
nand \U$34599 ( \34852 , \34850 , \34851 );
not \U$34600 ( \34853 , \34852 );
not \U$34601 ( \34854 , \4217 );
and \U$34602 ( \34855 , \34853 , \34854 );
and \U$34603 ( \34856 , \34852 , \1618 );
nor \U$34604 ( \34857 , \34855 , \34856 );
nor \U$34605 ( \34858 , \34847 , \34857 );
nor \U$34606 ( \34859 , \34836 , \34846 );
nor \U$34607 ( \34860 , \34858 , \34859 );
not \U$34608 ( \34861 , RIbe2b5b8_126);
not \U$34609 ( \34862 , \1112 );
or \U$34610 ( \34863 , \34861 , \34862 );
nand \U$34611 ( \34864 , \5467 , RIbe2a3e8_88);
nand \U$34612 ( \34865 , \34863 , \34864 );
and \U$34613 ( \34866 , \34865 , \1131 );
not \U$34614 ( \34867 , \34865 );
and \U$34615 ( \34868 , \34867 , \3491 );
nor \U$34616 ( \34869 , \34866 , \34868 );
not \U$34617 ( \34870 , RIbe2a988_100);
not \U$34618 ( \34871 , \5476 );
or \U$34619 ( \34872 , \34870 , \34871 );
nand \U$34620 ( \34873 , \4730 , RIbe2a910_99);
nand \U$34621 ( \34874 , \34872 , \34873 );
and \U$34622 ( \34875 , \34874 , \1309 );
not \U$34623 ( \34876 , \34874 );
and \U$34624 ( \34877 , \34876 , \4251 );
nor \U$34625 ( \34878 , \34875 , \34877 );
or \U$34626 ( \34879 , \34869 , \34878 );
not \U$34627 ( \34880 , \4064 );
not \U$34628 ( \34881 , \12755 );
and \U$34629 ( \34882 , \34880 , \34881 );
and \U$34630 ( \34883 , \8833 , RIbe2a370_87);
nor \U$34631 ( \34884 , \34882 , \34883 );
and \U$34632 ( \34885 , \34884 , \3516 );
not \U$34633 ( \34886 , \34884 );
and \U$34634 ( \34887 , \34886 , \1277 );
nor \U$34635 ( \34888 , \34885 , \34887 );
nand \U$34636 ( \34889 , \34879 , \34888 );
nand \U$34637 ( \34890 , \34869 , \34878 );
nand \U$34638 ( \34891 , \34889 , \34890 );
not \U$34639 ( \34892 , \34891 );
nand \U$34640 ( \34893 , \34860 , \34892 );
not \U$34641 ( \34894 , RIbe2acd0_107);
not \U$34642 ( \34895 , \8342 );
or \U$34643 ( \34896 , \34894 , \34895 );
nand \U$34644 ( \34897 , \4284 , RIbe2a028_80);
nand \U$34645 ( \34898 , \34896 , \34897 );
and \U$34646 ( \34899 , \34898 , \4058 );
not \U$34647 ( \34900 , \34898 );
and \U$34648 ( \34901 , \34900 , \2576 );
nor \U$34649 ( \34902 , \34899 , \34901 );
not \U$34650 ( \34903 , \34902 );
not \U$34651 ( \34904 , RIbe29fb0_79);
not \U$34652 ( \34905 , \3451 );
or \U$34653 ( \34906 , \34904 , \34905 );
nand \U$34654 ( \34907 , \4011 , RIbe29e48_76);
nand \U$34655 ( \34908 , \34906 , \34907 );
and \U$34656 ( \34909 , \34908 , \4346 );
not \U$34657 ( \34910 , \34908 );
and \U$34658 ( \34911 , \34910 , \2887 );
nor \U$34659 ( \34912 , \34909 , \34911 );
not \U$34660 ( \34913 , \34912 );
or \U$34661 ( \34914 , \34903 , \34913 );
or \U$34662 ( \34915 , \34912 , \34902 );
not \U$34663 ( \34916 , RIbe29dd0_75);
not \U$34664 ( \34917 , \6783 );
or \U$34665 ( \34918 , \34916 , \34917 );
nand \U$34666 ( \34919 , \4332 , RIbe29c68_72);
nand \U$34667 ( \34920 , \34918 , \34919 );
and \U$34668 ( \34921 , \34920 , \3471 );
not \U$34669 ( \34922 , \34920 );
and \U$34670 ( \34923 , \34922 , \3448 );
nor \U$34671 ( \34924 , \34921 , \34923 );
nand \U$34672 ( \34925 , \34915 , \34924 );
nand \U$34673 ( \34926 , \34914 , \34925 );
and \U$34674 ( \34927 , \34893 , \34926 );
nor \U$34675 ( \34928 , \34860 , \34892 );
nor \U$34676 ( \34929 , \34927 , \34928 );
not \U$34677 ( \34930 , \34929 );
not \U$34678 ( \34931 , RIbe289a8_32);
not \U$34679 ( \34932 , \6942 );
or \U$34680 ( \34933 , \34931 , \34932 );
nand \U$34681 ( \34934 , \7981 , RIbe28930_31);
nand \U$34682 ( \34935 , \34933 , \34934 );
and \U$34683 ( \34936 , \34935 , \6948 );
not \U$34684 ( \34937 , \34935 );
and \U$34685 ( \34938 , \34937 , \12234 );
nor \U$34686 ( \34939 , \34936 , \34938 );
not \U$34687 ( \34940 , \34939 );
not \U$34688 ( \34941 , RIbe28b10_35);
not \U$34689 ( \34942 , \8199 );
or \U$34690 ( \34943 , \34941 , \34942 );
nand \U$34691 ( \34944 , \8202 , RIbe28b88_36);
nand \U$34692 ( \34945 , \34943 , \34944 );
xor \U$34693 ( \34946 , \34945 , \6572 );
not \U$34694 ( \34947 , \34946 );
nand \U$34695 ( \34948 , \34940 , \34947 );
not \U$34696 ( \34949 , \34946 );
not \U$34697 ( \34950 , \34939 );
or \U$34698 ( \34951 , \34949 , \34950 );
not \U$34699 ( \34952 , \7301 );
not \U$34700 ( \34953 , RIbe29290_51);
not \U$34701 ( \34954 , \7298 );
or \U$34702 ( \34955 , \34953 , \34954 );
nand \U$34703 ( \34956 , \13224 , RIbe28a20_33);
nand \U$34704 ( \34957 , \34955 , \34956 );
not \U$34705 ( \34958 , \34957 );
or \U$34706 ( \34959 , \34952 , \34958 );
or \U$34707 ( \34960 , \34957 , \6992 );
nand \U$34708 ( \34961 , \34959 , \34960 );
nand \U$34709 ( \34962 , \34951 , \34961 );
nand \U$34710 ( \34963 , \34948 , \34962 );
not \U$34711 ( \34964 , RIbe28408_20);
not \U$34712 ( \34965 , \6868 );
or \U$34713 ( \34966 , \34964 , \34965 );
nand \U$34714 ( \34967 , \13436 , RIbe28390_19);
nand \U$34715 ( \34968 , \34966 , \34967 );
and \U$34716 ( \34969 , \34968 , \6873 );
not \U$34717 ( \34970 , \34968 );
and \U$34718 ( \34971 , \34970 , \7948 );
nor \U$34719 ( \34972 , \34969 , \34971 );
not \U$34720 ( \34973 , \34972 );
not \U$34721 ( \34974 , \34973 );
not \U$34722 ( \34975 , RIbe28660_25);
not \U$34723 ( \34976 , \8231 );
or \U$34724 ( \34977 , \34975 , \34976 );
nand \U$34725 ( \34978 , \8235 , RIbe285e8_24);
nand \U$34726 ( \34979 , \34977 , \34978 );
and \U$34727 ( \34980 , \34979 , \6141 );
not \U$34728 ( \34981 , \34979 );
and \U$34729 ( \34982 , \34981 , \7534 );
nor \U$34730 ( \34983 , \34980 , \34982 );
not \U$34731 ( \34984 , \34983 );
not \U$34732 ( \34985 , \34984 );
or \U$34733 ( \34986 , \34974 , \34985 );
not \U$34734 ( \34987 , \34972 );
not \U$34735 ( \34988 , \34983 );
or \U$34736 ( \34989 , \34987 , \34988 );
not \U$34737 ( \34990 , \13412 );
not \U$34738 ( \34991 , RIbe287c8_28);
not \U$34739 ( \34992 , \6536 );
or \U$34740 ( \34993 , \34991 , \34992 );
nand \U$34741 ( \34994 , \6540 , RIbe28480_21);
nand \U$34742 ( \34995 , \34993 , \34994 );
not \U$34743 ( \34996 , \34995 );
or \U$34744 ( \34997 , \34990 , \34996 );
or \U$34745 ( \34998 , \6891 , \34995 );
nand \U$34746 ( \34999 , \34997 , \34998 );
nand \U$34747 ( \35000 , \34989 , \34999 );
nand \U$34748 ( \35001 , \34986 , \35000 );
or \U$34749 ( \35002 , \34963 , \35001 );
not \U$34750 ( \35003 , RIbe29bf0_71);
not \U$34751 ( \35004 , \4595 );
or \U$34752 ( \35005 , \35003 , \35004 );
nand \U$34753 ( \35006 , \4600 , RIbe28f48_44);
nand \U$34754 ( \35007 , \35005 , \35006 );
not \U$34755 ( \35008 , \35007 );
not \U$34756 ( \35009 , \4323 );
and \U$34757 ( \35010 , \35008 , \35009 );
and \U$34758 ( \35011 , \35007 , \4323 );
nor \U$34759 ( \35012 , \35010 , \35011 );
not \U$34760 ( \35013 , \35012 );
not \U$34761 ( \35014 , \35013 );
not \U$34762 ( \35015 , RIbe27f58_10);
not \U$34763 ( \35016 , \6630 );
or \U$34764 ( \35017 , \35015 , \35016 );
nand \U$34765 ( \35018 , \14239 , RIbe27e68_8);
nand \U$34766 ( \35019 , \35017 , \35018 );
xor \U$34767 ( \35020 , \35019 , \5754 );
not \U$34768 ( \35021 , \35020 );
not \U$34769 ( \35022 , \35021 );
or \U$34770 ( \35023 , \35014 , \35022 );
not \U$34771 ( \35024 , \35012 );
not \U$34772 ( \35025 , \35020 );
or \U$34773 ( \35026 , \35024 , \35025 );
not \U$34774 ( \35027 , RIbe28ed0_43);
not \U$34775 ( \35028 , \4830 );
or \U$34776 ( \35029 , \35027 , \35028 );
nand \U$34777 ( \35030 , \5052 , RIbe27fd0_11);
nand \U$34778 ( \35031 , \35029 , \35030 );
and \U$34779 ( \35032 , \35031 , \4586 );
not \U$34780 ( \35033 , \35031 );
and \U$34781 ( \35034 , \35033 , \4946 );
nor \U$34782 ( \35035 , \35032 , \35034 );
nand \U$34783 ( \35036 , \35026 , \35035 );
nand \U$34784 ( \35037 , \35023 , \35036 );
and \U$34785 ( \35038 , \35002 , \35037 );
and \U$34786 ( \35039 , \34963 , \35001 );
nor \U$34787 ( \35040 , \35038 , \35039 );
not \U$34788 ( \35041 , \35040 );
or \U$34789 ( \35042 , \34930 , \35041 );
not \U$34790 ( \35043 , RIbe29920_65);
not \U$34791 ( \35044 , \13690 );
or \U$34792 ( \35045 , \35043 , \35044 );
nand \U$34793 ( \35046 , RIbe27b98_2, RIbe2ae38_110);
nand \U$34794 ( \35047 , \35045 , \35046 );
xnor \U$34795 ( \35048 , \35047 , RIbe2aeb0_111);
not \U$34796 ( \35049 , RIbe28e58_42);
not \U$34797 ( \35050 , \12887 );
or \U$34798 ( \35051 , \35049 , \35050 );
nand \U$34799 ( \35052 , \12794 , RIbe28de0_41);
nand \U$34800 ( \35053 , \35051 , \35052 );
not \U$34801 ( \35054 , \35053 );
not \U$34802 ( \35055 , \12998 );
and \U$34803 ( \35056 , \35054 , \35055 );
and \U$34804 ( \35057 , \35053 , \12801 );
nor \U$34805 ( \35058 , \35056 , \35057 );
xor \U$34806 ( \35059 , \35048 , \35058 );
not \U$34807 ( \35060 , RIbe27d00_5);
not \U$34808 ( \35061 , \13590 );
or \U$34809 ( \35062 , \35060 , \35061 );
nand \U$34810 ( \35063 , \12835 , RIbe27c10_3);
nand \U$34811 ( \35064 , \35062 , \35063 );
not \U$34812 ( \35065 , \35064 );
not \U$34813 ( \35066 , \12823 );
and \U$34814 ( \35067 , \35065 , \35066 );
and \U$34815 ( \35068 , \35064 , \12823 );
nor \U$34816 ( \35069 , \35067 , \35068 );
and \U$34817 ( \35070 , \35059 , \35069 );
and \U$34818 ( \35071 , \35048 , \35058 );
or \U$34819 ( \35072 , \35070 , \35071 );
not \U$34820 ( \35073 , \35072 );
and \U$34821 ( \35074 , \13478 , RIbe29560_57);
and \U$34822 ( \35075 , \13380 , RIbe28228_16);
nor \U$34823 ( \35076 , \35074 , \35075 );
and \U$34824 ( \35077 , \35076 , \7970 );
not \U$34825 ( \35078 , \35076 );
and \U$34826 ( \35079 , \35078 , \10912 );
nor \U$34827 ( \35080 , \35077 , \35079 );
not \U$34828 ( \35081 , RIbe29830_63);
not \U$34829 ( \35082 , \13049 );
or \U$34830 ( \35083 , \35081 , \35082 );
nand \U$34831 ( \35084 , \12948 , RIbe296c8_60);
nand \U$34832 ( \35085 , \35083 , \35084 );
not \U$34833 ( \35086 , \35085 );
not \U$34834 ( \35087 , \12957 );
and \U$34835 ( \35088 , \35086 , \35087 );
and \U$34836 ( \35089 , \35085 , \12957 );
nor \U$34837 ( \35090 , \35088 , \35089 );
xor \U$34838 ( \35091 , \35080 , \35090 );
not \U$34839 ( \35092 , RIbe281b0_15);
not \U$34840 ( \35093 , \13024 );
or \U$34841 ( \35094 , \35092 , \35093 );
nand \U$34842 ( \35095 , \14511 , RIbe280c0_13);
nand \U$34843 ( \35096 , \35094 , \35095 );
not \U$34844 ( \35097 , \35096 );
not \U$34845 ( \35098 , \13030 );
and \U$34846 ( \35099 , \35097 , \35098 );
and \U$34847 ( \35100 , \35096 , \13033 );
nor \U$34848 ( \35101 , \35099 , \35100 );
and \U$34849 ( \35102 , \35091 , \35101 );
and \U$34850 ( \35103 , \35080 , \35090 );
or \U$34851 ( \35104 , \35102 , \35103 );
not \U$34852 ( \35105 , \35104 );
or \U$34853 ( \35106 , \35073 , \35105 );
not \U$34854 ( \35107 , RIbe28fc0_45);
not \U$34855 ( \35108 , \14523 );
or \U$34856 ( \35109 , \35107 , \35108 );
nand \U$34857 ( \35110 , \12711 , RIbe290b0_47);
nand \U$34858 ( \35111 , \35109 , \35110 );
and \U$34859 ( \35112 , \35111 , \13068 );
not \U$34860 ( \35113 , \35111 );
and \U$34861 ( \35114 , \35113 , \13583 );
nor \U$34862 ( \35115 , \35112 , \35114 );
not \U$34863 ( \35116 , \12752 );
not \U$34864 ( \35117 , \2355 );
and \U$34865 ( \35118 , \35116 , \35117 );
and \U$34866 ( \35119 , \13092 , RIbe29650_59);
nor \U$34867 ( \35120 , \35118 , \35119 );
and \U$34868 ( \35121 , \35120 , \12770 );
not \U$34869 ( \35122 , \35120 );
and \U$34870 ( \35123 , \35122 , \12927 );
nor \U$34871 ( \35124 , \35121 , \35123 );
xor \U$34872 ( \35125 , \35115 , \35124 );
not \U$34873 ( \35126 , RIbe29a88_68);
not \U$34874 ( \35127 , \12732 );
or \U$34875 ( \35128 , \35126 , \35127 );
nand \U$34876 ( \35129 , \13077 , RIbe27d78_6);
nand \U$34877 ( \35130 , \35128 , \35129 );
and \U$34878 ( \35131 , \35130 , \12743 );
not \U$34879 ( \35132 , \35130 );
and \U$34880 ( \35133 , \35132 , \12742 );
nor \U$34881 ( \35134 , \35131 , \35133 );
and \U$34882 ( \35135 , \35125 , \35134 );
and \U$34883 ( \35136 , \35115 , \35124 );
or \U$34884 ( \35137 , \35135 , \35136 );
nand \U$34885 ( \35138 , \35106 , \35137 );
not \U$34886 ( \35139 , \35072 );
not \U$34887 ( \35140 , \35104 );
nand \U$34888 ( \35141 , \35139 , \35140 );
nand \U$34889 ( \35142 , \35138 , \35141 );
nand \U$34890 ( \35143 , \35042 , \35142 );
or \U$34891 ( \35144 , \35040 , \34929 );
and \U$34892 ( \35145 , \35143 , \35144 );
xor \U$34893 ( \35146 , \34098 , \34110 );
xor \U$34894 ( \35147 , \35146 , \34088 );
not \U$34895 ( \35148 , \35147 );
nand \U$34896 ( \35149 , RIbe29380_53, RIbe2ab68_104);
nand \U$34897 ( \35150 , \35148 , \35149 );
and \U$34898 ( \35151 , \3895 , RIbe2afa0_113);
and \U$34899 ( \35152 , \7116 , RIbe2af28_112);
nor \U$34900 ( \35153 , \35151 , \35152 );
and \U$34901 ( \35154 , \35153 , \300 );
not \U$34902 ( \35155 , \35153 );
and \U$34903 ( \35156 , \35155 , \293 );
nor \U$34904 ( \35157 , \35154 , \35156 );
not \U$34905 ( \35158 , \35157 );
and \U$34906 ( \35159 , \546 , RIbe2b270_119);
and \U$34907 ( \35160 , \552 , RIbe2b108_116);
nor \U$34908 ( \35161 , \35159 , \35160 );
and \U$34909 ( \35162 , \35161 , \424 );
not \U$34910 ( \35163 , \35161 );
and \U$34911 ( \35164 , \35163 , \425 );
nor \U$34912 ( \35165 , \35162 , \35164 );
not \U$34913 ( \35166 , \35165 );
or \U$34914 ( \35167 , \35158 , \35166 );
or \U$34915 ( \35168 , \35165 , \35157 );
not \U$34916 ( \35169 , RIbe2b1f8_118);
not \U$34917 ( \35170 , \1773 );
or \U$34918 ( \35171 , \35169 , \35170 );
nand \U$34919 ( \35172 , \429 , RIbe2b180_117);
nand \U$34920 ( \35173 , \35171 , \35172 );
and \U$34921 ( \35174 , \35173 , \1547 );
not \U$34922 ( \35175 , \35173 );
and \U$34923 ( \35176 , \35175 , \306 );
nor \U$34924 ( \35177 , \35174 , \35176 );
not \U$34925 ( \35178 , \35177 );
nand \U$34926 ( \35179 , \35168 , \35178 );
nand \U$34927 ( \35180 , \35167 , \35179 );
and \U$34928 ( \35181 , \35150 , \35180 );
nor \U$34929 ( \35182 , \35148 , \35149 );
nor \U$34930 ( \35183 , \35181 , \35182 );
not \U$34931 ( \35184 , \33764 );
and \U$34932 ( \35185 , \33753 , \33740 );
not \U$34933 ( \35186 , \33753 );
and \U$34934 ( \35187 , \35186 , \33741 );
nor \U$34935 ( \35188 , \35185 , \35187 );
not \U$34936 ( \35189 , \35188 );
or \U$34937 ( \35190 , \35184 , \35189 );
or \U$34938 ( \35191 , \33764 , \35188 );
nand \U$34939 ( \35192 , \35190 , \35191 );
not \U$34940 ( \35193 , \35192 );
not \U$34941 ( \35194 , \33725 );
not \U$34942 ( \35195 , \33714 );
not \U$34943 ( \35196 , \33704 );
and \U$34944 ( \35197 , \35195 , \35196 );
and \U$34945 ( \35198 , \33714 , \33704 );
nor \U$34946 ( \35199 , \35197 , \35198 );
not \U$34947 ( \35200 , \35199 );
and \U$34948 ( \35201 , \35194 , \35200 );
and \U$34949 ( \35202 , \33725 , \35199 );
nor \U$34950 ( \35203 , \35201 , \35202 );
nand \U$34951 ( \35204 , \35193 , \35203 );
not \U$34952 ( \35205 , \35204 );
not \U$34953 ( \35206 , \33816 );
not \U$34954 ( \35207 , \33834 );
or \U$34955 ( \35208 , \35206 , \35207 );
or \U$34956 ( \35209 , \33816 , \33834 );
nand \U$34957 ( \35210 , \35208 , \35209 );
and \U$34958 ( \35211 , \35210 , \33836 );
not \U$34959 ( \35212 , \35210 );
and \U$34960 ( \35213 , \35212 , \33823 );
nor \U$34961 ( \35214 , \35211 , \35213 );
not \U$34962 ( \35215 , \35214 );
or \U$34963 ( \35216 , \35205 , \35215 );
not \U$34964 ( \35217 , \35203 );
nand \U$34965 ( \35218 , \35192 , \35217 );
nand \U$34966 ( \35219 , \35216 , \35218 );
not \U$34967 ( \35220 , \35219 );
nand \U$34968 ( \35221 , \35183 , \35220 );
xor \U$34969 ( \35222 , \34129 , \34139 );
xnor \U$34970 ( \35223 , \35222 , \34150 );
not \U$34971 ( \35224 , \35223 );
and \U$34972 ( \35225 , \33848 , \33869 );
not \U$34973 ( \35226 , \33848 );
and \U$34974 ( \35227 , \35226 , \33870 );
or \U$34975 ( \35228 , \35225 , \35227 );
xor \U$34976 ( \35229 , \35228 , \33858 );
not \U$34977 ( \35230 , \35229 );
not \U$34978 ( \35231 , \35230 );
or \U$34979 ( \35232 , \35224 , \35231 );
not \U$34980 ( \35233 , \35229 );
not \U$34981 ( \35234 , \35223 );
not \U$34982 ( \35235 , \35234 );
or \U$34983 ( \35236 , \35233 , \35235 );
not \U$34984 ( \35237 , \33900 );
not \U$34985 ( \35238 , \33890 );
not \U$34986 ( \35239 , \33914 );
or \U$34987 ( \35240 , \35238 , \35239 );
or \U$34988 ( \35241 , \33914 , \33890 );
nand \U$34989 ( \35242 , \35240 , \35241 );
not \U$34990 ( \35243 , \35242 );
or \U$34991 ( \35244 , \35237 , \35243 );
or \U$34992 ( \35245 , \35242 , \33900 );
nand \U$34993 ( \35246 , \35244 , \35245 );
buf \U$34994 ( \35247 , \35246 );
nand \U$34995 ( \35248 , \35236 , \35247 );
nand \U$34996 ( \35249 , \35232 , \35248 );
and \U$34997 ( \35250 , \35221 , \35249 );
nor \U$34998 ( \35251 , \35220 , \35183 );
nor \U$34999 ( \35252 , \35250 , \35251 );
nand \U$35000 ( \35253 , \35145 , \35252 );
or \U$35001 ( \35254 , \33777 , \33787 );
nand \U$35002 ( \35255 , \33787 , \33777 );
nand \U$35003 ( \35256 , \35254 , \35255 );
not \U$35004 ( \35257 , \33800 );
and \U$35005 ( \35258 , \35256 , \35257 );
not \U$35006 ( \35259 , \35256 );
and \U$35007 ( \35260 , \35259 , \33800 );
nor \U$35008 ( \35261 , \35258 , \35260 );
not \U$35009 ( \35262 , \33953 );
not \U$35010 ( \35263 , \33968 );
or \U$35011 ( \35264 , \35262 , \35263 );
or \U$35012 ( \35265 , \33953 , \33968 );
nand \U$35013 ( \35266 , \35264 , \35265 );
not \U$35014 ( \35267 , \33979 );
and \U$35015 ( \35268 , \35266 , \35267 );
not \U$35016 ( \35269 , \35266 );
and \U$35017 ( \35270 , \35269 , \33979 );
nor \U$35018 ( \35271 , \35268 , \35270 );
and \U$35019 ( \35272 , \35261 , \35271 );
xor \U$35020 ( \35273 , \34000 , \34008 );
xor \U$35021 ( \35274 , \35273 , \34018 );
not \U$35022 ( \35275 , \35274 );
nor \U$35023 ( \35276 , \35272 , \35275 );
nor \U$35024 ( \35277 , \35261 , \35271 );
nor \U$35025 ( \35278 , \35276 , \35277 );
not \U$35026 ( \35279 , \34034 );
not \U$35027 ( \35280 , \34037 );
and \U$35028 ( \35281 , \35279 , \35280 );
and \U$35029 ( \35282 , \34034 , \34037 );
nor \U$35030 ( \35283 , \35281 , \35282 );
and \U$35031 ( \35284 , \35278 , \35283 );
not \U$35032 ( \35285 , \34069 );
not \U$35033 ( \35286 , \35285 );
not \U$35034 ( \35287 , \34055 );
or \U$35035 ( \35288 , \35286 , \35287 );
nand \U$35036 ( \35289 , \34054 , \34069 );
nand \U$35037 ( \35290 , \35288 , \35289 );
not \U$35038 ( \35291 , \34043 );
and \U$35039 ( \35292 , \35290 , \35291 );
not \U$35040 ( \35293 , \35290 );
and \U$35041 ( \35294 , \35293 , \34043 );
nor \U$35042 ( \35295 , \35292 , \35294 );
or \U$35043 ( \35296 , \35284 , \35295 );
or \U$35044 ( \35297 , \35283 , \35278 );
nand \U$35045 ( \35298 , \35296 , \35297 );
and \U$35046 ( \35299 , \35253 , \35298 );
nor \U$35047 ( \35300 , \35252 , \35145 );
nor \U$35048 ( \35301 , \35299 , \35300 );
not \U$35049 ( \35302 , \35301 );
not \U$35050 ( \35303 , \35302 );
or \U$35051 ( \35304 , \34829 , \35303 );
not \U$35052 ( \35305 , \35301 );
not \U$35053 ( \35306 , \34828 );
not \U$35054 ( \35307 , \35306 );
or \U$35055 ( \35308 , \35305 , \35307 );
xor \U$35056 ( \35309 , \34228 , \34234 );
xor \U$35057 ( \35310 , \35309 , \34237 );
not \U$35058 ( \35311 , \35310 );
and \U$35059 ( \35312 , \34039 , \34031 );
not \U$35060 ( \35313 , \34039 );
and \U$35061 ( \35314 , \35313 , \34030 );
nor \U$35062 ( \35315 , \35312 , \35314 );
not \U$35063 ( \35316 , \34071 );
and \U$35064 ( \35317 , \35315 , \35316 );
not \U$35065 ( \35318 , \35315 );
and \U$35066 ( \35319 , \35318 , \34071 );
nor \U$35067 ( \35320 , \35317 , \35319 );
not \U$35068 ( \35321 , \35320 );
not \U$35069 ( \35322 , \35321 );
or \U$35070 ( \35323 , \35311 , \35322 );
not \U$35071 ( \35324 , \35320 );
not \U$35072 ( \35325 , \35310 );
not \U$35073 ( \35326 , \35325 );
or \U$35074 ( \35327 , \35324 , \35326 );
xor \U$35075 ( \35328 , \34242 , \34251 );
xor \U$35076 ( \35329 , \35328 , \34255 );
nand \U$35077 ( \35330 , \35327 , \35329 );
nand \U$35078 ( \35331 , \35323 , \35330 );
nand \U$35079 ( \35332 , \35308 , \35331 );
nand \U$35080 ( \35333 , \35304 , \35332 );
not \U$35081 ( \35334 , \35333 );
not \U$35082 ( \35335 , \33126 );
not \U$35083 ( \35336 , \33230 );
or \U$35084 ( \35337 , \35335 , \35336 );
nand \U$35085 ( \35338 , \33229 , \33127 );
nand \U$35086 ( \35339 , \35337 , \35338 );
xnor \U$35087 ( \35340 , \35339 , \33272 );
nand \U$35088 ( \35341 , \35334 , \35340 );
not \U$35089 ( \35342 , \35341 );
xor \U$35090 ( \35343 , \32924 , \33024 );
xor \U$35091 ( \35344 , \35343 , \33122 );
not \U$35092 ( \35345 , \35344 );
not \U$35093 ( \35346 , \34219 );
not \U$35094 ( \35347 , \34215 );
or \U$35095 ( \35348 , \35346 , \35347 );
nand \U$35096 ( \35349 , \34203 , \34214 );
nand \U$35097 ( \35350 , \35348 , \35349 );
not \U$35098 ( \35351 , \34223 );
and \U$35099 ( \35352 , \35350 , \35351 );
not \U$35100 ( \35353 , \35350 );
and \U$35101 ( \35354 , \35353 , \34223 );
nor \U$35102 ( \35355 , \35352 , \35354 );
nand \U$35103 ( \35356 , \35345 , \35355 );
not \U$35104 ( \35357 , \35356 );
xor \U$35105 ( \35358 , \34240 , \34258 );
xor \U$35106 ( \35359 , \35358 , \34264 );
not \U$35107 ( \35360 , \35359 );
or \U$35108 ( \35361 , \35357 , \35360 );
not \U$35109 ( \35362 , \35355 );
nand \U$35110 ( \35363 , \35362 , \35344 );
nand \U$35111 ( \35364 , \35361 , \35363 );
not \U$35112 ( \35365 , \35364 );
or \U$35113 ( \35366 , \35342 , \35365 );
not \U$35114 ( \35367 , \35340 );
nand \U$35115 ( \35368 , \35367 , \35333 );
nand \U$35116 ( \35369 , \35366 , \35368 );
xor \U$35117 ( \35370 , \34773 , \35369 );
xor \U$35118 ( \35371 , \34201 , \34225 );
xor \U$35119 ( \35372 , \35371 , \34267 );
not \U$35120 ( \35373 , \35372 );
xor \U$35121 ( \35374 , \34276 , \34282 );
xor \U$35122 ( \35375 , \35374 , \34289 );
nor \U$35123 ( \35376 , \35373 , \35375 );
and \U$35124 ( \35377 , \35370 , \35376 );
and \U$35125 ( \35378 , \34773 , \35369 );
or \U$35126 ( \35379 , \35377 , \35378 );
or \U$35127 ( \35380 , \34294 , \35379 );
nor \U$35128 ( \35381 , \34270 , \33698 );
not \U$35129 ( \35382 , \35381 );
not \U$35130 ( \35383 , \34292 );
and \U$35131 ( \35384 , \35382 , \35383 );
and \U$35132 ( \35385 , \34270 , \33698 );
nor \U$35133 ( \35386 , \35384 , \35385 );
xor \U$35134 ( \35387 , \34752 , \34758 );
and \U$35135 ( \35388 , \35387 , \34763 );
and \U$35136 ( \35389 , \34752 , \34758 );
or \U$35137 ( \35390 , \35388 , \35389 );
not \U$35138 ( \35391 , \34299 );
not \U$35139 ( \35392 , \34311 );
or \U$35140 ( \35393 , \35391 , \35392 );
nand \U$35141 ( \35394 , \35393 , \34304 );
nand \U$35142 ( \35395 , \34308 , \34298 );
nand \U$35143 ( \35396 , \35394 , \35395 );
xor \U$35144 ( \35397 , \35390 , \35396 );
not \U$35145 ( \35398 , \34628 );
not \U$35146 ( \35399 , \34639 );
or \U$35147 ( \35400 , \35398 , \35399 );
or \U$35148 ( \35401 , \34639 , \34628 );
nand \U$35149 ( \35402 , \35401 , \34746 );
nand \U$35150 ( \35403 , \35400 , \35402 );
xnor \U$35151 ( \35404 , \35397 , \35403 );
not \U$35152 ( \35405 , \34533 );
and \U$35153 ( \35406 , \34544 , \35405 );
nor \U$35154 ( \35407 , \35406 , \34524 );
nor \U$35155 ( \35408 , \34544 , \35405 );
nor \U$35156 ( \35409 , \35407 , \35408 );
nand \U$35157 ( \35410 , RIbe29380_53, RIbe2b1f8_118);
and \U$35158 ( \35411 , \12312 , RIbe2b180_117);
and \U$35159 ( \35412 , \329 , RIbe2b270_119);
nor \U$35160 ( \35413 , \35411 , \35412 );
and \U$35161 ( \35414 , \35413 , \338 );
not \U$35162 ( \35415 , \35413 );
and \U$35163 ( \35416 , \35415 , \337 );
nor \U$35164 ( \35417 , \35414 , \35416 );
xor \U$35165 ( \35418 , \35410 , \35417 );
and \U$35166 ( \35419 , \1659 , RIbe2b108_116);
and \U$35167 ( \35420 , \263 , RIbe2b090_115);
nor \U$35168 ( \35421 , \35419 , \35420 );
and \U$35169 ( \35422 , \35421 , \1362 );
not \U$35170 ( \35423 , \35421 );
and \U$35171 ( \35424 , \35423 , \1663 );
or \U$35172 ( \35425 , \35422 , \35424 );
xor \U$35173 ( \35426 , \35418 , \35425 );
or \U$35174 ( \35427 , \35409 , \35426 );
nand \U$35175 ( \35428 , \35426 , \35409 );
nand \U$35176 ( \35429 , \35427 , \35428 );
not \U$35177 ( \35430 , \35429 );
not \U$35178 ( \35431 , \35430 );
not \U$35179 ( \35432 , \34488 );
not \U$35180 ( \35433 , \34500 );
or \U$35181 ( \35434 , \35432 , \35433 );
nand \U$35182 ( \35435 , \35434 , \34479 );
nand \U$35183 ( \35436 , \34503 , \34491 );
nand \U$35184 ( \35437 , \35435 , \35436 );
not \U$35185 ( \35438 , \35437 );
not \U$35186 ( \35439 , \35438 );
not \U$35187 ( \35440 , \34600 );
and \U$35188 ( \35441 , \35440 , \34586 );
nor \U$35189 ( \35442 , \35441 , \34592 );
nor \U$35190 ( \35443 , \35440 , \34586 );
nor \U$35191 ( \35444 , \35442 , \35443 );
not \U$35192 ( \35445 , \35444 );
not \U$35193 ( \35446 , \35445 );
or \U$35194 ( \35447 , \35439 , \35446 );
nand \U$35195 ( \35448 , \35444 , \35437 );
nand \U$35196 ( \35449 , \35447 , \35448 );
not \U$35197 ( \35450 , \34564 );
and \U$35198 ( \35451 , \35450 , \34574 );
nor \U$35199 ( \35452 , \35451 , \34555 );
nor \U$35200 ( \35453 , \35450 , \34574 );
nor \U$35201 ( \35454 , \35452 , \35453 );
and \U$35202 ( \35455 , \35449 , \35454 );
not \U$35203 ( \35456 , \35449 );
not \U$35204 ( \35457 , \35454 );
and \U$35205 ( \35458 , \35456 , \35457 );
nor \U$35206 ( \35459 , \35455 , \35458 );
or \U$35207 ( \35460 , \35431 , \35459 );
nand \U$35208 ( \35461 , \35459 , \35429 );
nand \U$35209 ( \35462 , \35460 , \35461 );
not \U$35210 ( \35463 , RIbe29e48_76);
not \U$35211 ( \35464 , \8823 );
or \U$35212 ( \35465 , \35463 , \35464 );
nand \U$35213 ( \35466 , \20849 , RIbe29dd0_75);
nand \U$35214 ( \35467 , \35465 , \35466 );
not \U$35215 ( \35468 , \35467 );
not \U$35216 ( \35469 , \1448 );
and \U$35217 ( \35470 , \35468 , \35469 );
and \U$35218 ( \35471 , \35467 , \6831 );
nor \U$35219 ( \35472 , \35470 , \35471 );
not \U$35220 ( \35473 , RIbe29c68_72);
not \U$35221 ( \35474 , \2583 );
or \U$35222 ( \35475 , \35473 , \35474 );
nand \U$35223 ( \35476 , \2384 , RIbe29bf0_71);
nand \U$35224 ( \35477 , \35475 , \35476 );
and \U$35225 ( \35478 , \35477 , \1277 );
not \U$35226 ( \35479 , \35477 );
and \U$35227 ( \35480 , \35479 , \1076 );
nor \U$35228 ( \35481 , \35478 , \35480 );
xnor \U$35229 ( \35482 , \35472 , \35481 );
not \U$35230 ( \35483 , RIbe2a028_80);
not \U$35231 ( \35484 , \1632 );
or \U$35232 ( \35485 , \35483 , \35484 );
nand \U$35233 ( \35486 , \2817 , RIbe29fb0_79);
nand \U$35234 ( \35487 , \35485 , \35486 );
not \U$35235 ( \35488 , \35487 );
not \U$35236 ( \35489 , \1458 );
and \U$35237 ( \35490 , \35488 , \35489 );
and \U$35238 ( \35491 , \35487 , \1082 );
nor \U$35239 ( \35492 , \35490 , \35491 );
xor \U$35240 ( \35493 , \35482 , \35492 );
not \U$35241 ( \35494 , \35493 );
not \U$35242 ( \35495 , \35494 );
and \U$35243 ( \35496 , \5365 , RIbe2a280_85);
and \U$35244 ( \35497 , \1682 , RIbe2a208_84);
nor \U$35245 ( \35498 , \35496 , \35497 );
and \U$35246 ( \35499 , \35498 , \300 );
not \U$35247 ( \35500 , \35498 );
and \U$35248 ( \35501 , \35500 , \293 );
nor \U$35249 ( \35502 , \35499 , \35501 );
not \U$35250 ( \35503 , \428 );
or \U$35251 ( \35504 , \35503 , RIbe2a5c8_92);
not \U$35252 ( \35505 , RIbe2a190_83);
not \U$35253 ( \35506 , \380 );
or \U$35254 ( \35507 , \35505 , \35506 );
nand \U$35255 ( \35508 , \35507 , \35503 );
nand \U$35256 ( \35509 , \35504 , \35508 );
and \U$35257 ( \35510 , \35509 , \306 );
not \U$35258 ( \35511 , \35509 );
and \U$35259 ( \35512 , \35511 , \313 );
nor \U$35260 ( \35513 , \35510 , \35512 );
not \U$35261 ( \35514 , \35513 );
not \U$35262 ( \35515 , \35514 );
not \U$35263 ( \35516 , RIbe2a550_91);
not \U$35264 ( \35517 , \546 );
or \U$35265 ( \35518 , \35516 , \35517 );
nand \U$35266 ( \35519 , \552 , RIbe2a988_100);
nand \U$35267 ( \35520 , \35518 , \35519 );
not \U$35268 ( \35521 , \35520 );
not \U$35269 ( \35522 , \424 );
and \U$35270 ( \35523 , \35521 , \35522 );
and \U$35271 ( \35524 , \35520 , \7124 );
nor \U$35272 ( \35525 , \35523 , \35524 );
not \U$35273 ( \35526 , \35525 );
or \U$35274 ( \35527 , \35515 , \35526 );
or \U$35275 ( \35528 , \35525 , \35514 );
nand \U$35276 ( \35529 , \35527 , \35528 );
xnor \U$35277 ( \35530 , \35502 , \35529 );
not \U$35278 ( \35531 , \35530 );
and \U$35279 ( \35532 , \1146 , RIbe2acd0_107);
not \U$35280 ( \35533 , \1146 );
and \U$35281 ( \35534 , \1140 , RIbe2a2f8_86);
and \U$35282 ( \35535 , \35533 , \35534 );
nor \U$35283 ( \35536 , \35532 , \35535 );
and \U$35284 ( \35537 , \35536 , \1153 );
not \U$35285 ( \35538 , \35536 );
and \U$35286 ( \35539 , \35538 , \1794 );
nor \U$35287 ( \35540 , \35537 , \35539 );
not \U$35288 ( \35541 , \3959 );
not \U$35289 ( \35542 , \6345 );
not \U$35290 ( \35543 , \13531 );
and \U$35291 ( \35544 , \35542 , \35543 );
and \U$35292 ( \35545 , \7363 , RIbe2a910_99);
nor \U$35293 ( \35546 , \35544 , \35545 );
not \U$35294 ( \35547 , \35546 );
or \U$35295 ( \35548 , \35541 , \35547 );
or \U$35296 ( \35549 , \35546 , \3959 );
nand \U$35297 ( \35550 , \35548 , \35549 );
xor \U$35298 ( \35551 , \35540 , \35550 );
not \U$35299 ( \35552 , \1813 );
not \U$35300 ( \35553 , RIbe2a3e8_88);
not \U$35301 ( \35554 , \6747 );
or \U$35302 ( \35555 , \35553 , \35554 );
nand \U$35303 ( \35556 , \1203 , RIbe2a370_87);
nand \U$35304 ( \35557 , \35555 , \35556 );
not \U$35305 ( \35558 , \35557 );
or \U$35306 ( \35559 , \35552 , \35558 );
or \U$35307 ( \35560 , \35557 , \752 );
nand \U$35308 ( \35561 , \35559 , \35560 );
xor \U$35309 ( \35562 , \35551 , \35561 );
not \U$35310 ( \35563 , \35562 );
or \U$35311 ( \35564 , \35531 , \35563 );
or \U$35312 ( \35565 , \35562 , \35530 );
nand \U$35313 ( \35566 , \35564 , \35565 );
not \U$35314 ( \35567 , \35566 );
not \U$35315 ( \35568 , \35567 );
or \U$35316 ( \35569 , \35495 , \35568 );
nand \U$35317 ( \35570 , \35566 , \35493 );
nand \U$35318 ( \35571 , \35569 , \35570 );
not \U$35319 ( \35572 , \35571 );
and \U$35320 ( \35573 , \35462 , \35572 );
not \U$35321 ( \35574 , \35462 );
and \U$35322 ( \35575 , \35574 , \35571 );
nor \U$35323 ( \35576 , \35573 , \35575 );
not \U$35324 ( \35577 , \35576 );
not \U$35325 ( \35578 , \34353 );
not \U$35326 ( \35579 , \34346 );
or \U$35327 ( \35580 , \35578 , \35579 );
not \U$35328 ( \35581 , \34352 );
not \U$35329 ( \35582 , \34347 );
or \U$35330 ( \35583 , \35581 , \35582 );
nand \U$35331 ( \35584 , \35583 , \34365 );
nand \U$35332 ( \35585 , \35580 , \35584 );
not \U$35333 ( \35586 , \35585 );
not \U$35334 ( \35587 , \35586 );
xor \U$35335 ( \35588 , \34330 , \34334 );
and \U$35336 ( \35589 , \35588 , \34339 );
and \U$35337 ( \35590 , \34330 , \34334 );
or \U$35338 ( \35591 , \35589 , \35590 );
not \U$35339 ( \35592 , \35591 );
or \U$35340 ( \35593 , \35587 , \35592 );
or \U$35341 ( \35594 , \35591 , \35586 );
nand \U$35342 ( \35595 , \35593 , \35594 );
not \U$35343 ( \35596 , \35595 );
xor \U$35344 ( \35597 , \34375 , \34380 );
and \U$35345 ( \35598 , \35597 , \34386 );
and \U$35346 ( \35599 , \34375 , \34380 );
or \U$35347 ( \35600 , \35598 , \35599 );
not \U$35348 ( \35601 , \35600 );
and \U$35349 ( \35602 , \35596 , \35601 );
and \U$35350 ( \35603 , \35595 , \35600 );
nor \U$35351 ( \35604 , \35602 , \35603 );
xor \U$35352 ( \35605 , \34507 , \33431 );
and \U$35353 ( \35606 , \35605 , \34512 );
and \U$35354 ( \35607 , \34507 , \33431 );
or \U$35355 ( \35608 , \35606 , \35607 );
xor \U$35356 ( \35609 , \34433 , \34469 );
and \U$35357 ( \35610 , \35609 , \34505 );
and \U$35358 ( \35611 , \34433 , \34469 );
or \U$35359 ( \35612 , \35610 , \35611 );
not \U$35360 ( \35613 , \35612 );
xor \U$35361 ( \35614 , \35608 , \35613 );
xor \U$35362 ( \35615 , \34545 , \34575 );
and \U$35363 ( \35616 , \35615 , \34601 );
and \U$35364 ( \35617 , \34545 , \34575 );
or \U$35365 ( \35618 , \35616 , \35617 );
xor \U$35366 ( \35619 , \35614 , \35618 );
xor \U$35367 ( \35620 , \35604 , \35619 );
xor \U$35368 ( \35621 , \35577 , \35620 );
nand \U$35369 ( \35622 , \34670 , \34647 );
and \U$35370 ( \35623 , \35622 , \34656 );
nor \U$35371 ( \35624 , \34670 , \34647 );
nor \U$35372 ( \35625 , \35623 , \35624 );
not \U$35373 ( \35626 , \34685 );
not \U$35374 ( \35627 , \34695 );
or \U$35375 ( \35628 , \35626 , \35627 );
nand \U$35376 ( \35629 , \35628 , \34708 );
nand \U$35377 ( \35630 , \34686 , \34694 );
nand \U$35378 ( \35631 , \35629 , \35630 );
xor \U$35379 ( \35632 , \35625 , \35631 );
nand \U$35380 ( \35633 , \34614 , \14555 );
and \U$35381 ( \35634 , \35633 , \34623 );
nor \U$35382 ( \35635 , \34614 , \18364 );
nor \U$35383 ( \35636 , \35634 , \35635 );
xnor \U$35384 ( \35637 , \35632 , \35636 );
not \U$35385 ( \35638 , \3456 );
and \U$35386 ( \35639 , RIbe27fd0_11, \3281 );
and \U$35387 ( \35640 , \35638 , \35639 );
not \U$35388 ( \35641 , \35638 );
and \U$35389 ( \35642 , \35641 , RIbe27f58_10);
nor \U$35390 ( \35643 , \35640 , \35642 );
and \U$35391 ( \35644 , \35643 , \2887 );
not \U$35392 ( \35645 , \35643 );
and \U$35393 ( \35646 , \35645 , \4346 );
nor \U$35394 ( \35647 , \35644 , \35646 );
nand \U$35395 ( \35648 , \3701 , RIbe27e68_8);
not \U$35396 ( \35649 , \35648 );
not \U$35397 ( \35650 , \4025 );
or \U$35398 ( \35651 , \35649 , \35650 );
nand \U$35399 ( \35652 , \6787 , \25899 );
nand \U$35400 ( \35653 , \35651 , \35652 );
not \U$35401 ( \35654 , \35653 );
not \U$35402 ( \35655 , \3471 );
and \U$35403 ( \35656 , \35654 , \35655 );
and \U$35404 ( \35657 , \35653 , \3471 );
nor \U$35405 ( \35658 , \35656 , \35657 );
xor \U$35406 ( \35659 , \35647 , \35658 );
not \U$35407 ( \35660 , RIbe28f48_44);
not \U$35408 ( \35661 , \2898 );
or \U$35409 ( \35662 , \35660 , \35661 );
nand \U$35410 ( \35663 , \2901 , RIbe28ed0_43);
nand \U$35411 ( \35664 , \35662 , \35663 );
and \U$35412 ( \35665 , \35664 , \2380 );
not \U$35413 ( \35666 , \35664 );
and \U$35414 ( \35667 , \35666 , \6468 );
nor \U$35415 ( \35668 , \35665 , \35667 );
xnor \U$35416 ( \35669 , \35659 , \35668 );
not \U$35417 ( \35670 , \35669 );
not \U$35418 ( \35671 , \35670 );
not \U$35419 ( \35672 , RIbe28930_31);
not \U$35420 ( \35673 , \7941 );
or \U$35421 ( \35674 , \35672 , \35673 );
not \U$35422 ( \35675 , \28220 );
nand \U$35423 ( \35676 , \35675 , \6596 );
nand \U$35424 ( \35677 , \35674 , \35676 );
and \U$35425 ( \35678 , \35677 , \7948 );
not \U$35426 ( \35679 , \35677 );
and \U$35427 ( \35680 , \35679 , \7488 );
nor \U$35428 ( \35681 , \35678 , \35680 );
not \U$35429 ( \35682 , \35681 );
not \U$35430 ( \35683 , RIbe28a20_33);
not \U$35431 ( \35684 , \6535 );
or \U$35432 ( \35685 , \35683 , \35684 );
nand \U$35433 ( \35686 , \7075 , RIbe289a8_32);
nand \U$35434 ( \35687 , \35685 , \35686 );
not \U$35435 ( \35688 , \35687 );
not \U$35436 ( \35689 , \6891 );
and \U$35437 ( \35690 , \35688 , \35689 );
and \U$35438 ( \35691 , \35687 , \13412 );
nor \U$35439 ( \35692 , \35690 , \35691 );
not \U$35440 ( \35693 , \35692 );
or \U$35441 ( \35694 , \35682 , \35693 );
or \U$35442 ( \35695 , \35681 , \35692 );
nand \U$35443 ( \35696 , \35694 , \35695 );
not \U$35444 ( \35697 , RIbe28b88_36);
not \U$35445 ( \35698 , \12268 );
or \U$35446 ( \35699 , \35697 , \35698 );
nand \U$35447 ( \35700 , \9939 , RIbe29290_51);
nand \U$35448 ( \35701 , \35699 , \35700 );
and \U$35449 ( \35702 , \35701 , \6620 );
not \U$35450 ( \35703 , \35701 );
and \U$35451 ( \35704 , \35703 , \5740 );
nor \U$35452 ( \35705 , \35702 , \35704 );
not \U$35453 ( \35706 , \35705 );
and \U$35454 ( \35707 , \35696 , \35706 );
not \U$35455 ( \35708 , \35696 );
and \U$35456 ( \35709 , \35708 , \35705 );
nor \U$35457 ( \35710 , \35707 , \35709 );
not \U$35458 ( \35711 , \35710 );
not \U$35459 ( \35712 , \35711 );
or \U$35460 ( \35713 , \35671 , \35712 );
nand \U$35461 ( \35714 , \35669 , \35710 );
nand \U$35462 ( \35715 , \35713 , \35714 );
not \U$35463 ( \35716 , RIbe28480_21);
not \U$35464 ( \35717 , \15894 );
or \U$35465 ( \35718 , \35716 , \35717 );
nand \U$35466 ( \35719 , \22378 , RIbe28408_20);
nand \U$35467 ( \35720 , \35718 , \35719 );
and \U$35468 ( \35721 , \35720 , \20465 );
not \U$35469 ( \35722 , \35720 );
and \U$35470 ( \35723 , \35722 , \4586 );
nor \U$35471 ( \35724 , \35721 , \35723 );
not \U$35472 ( \35725 , \35724 );
not \U$35473 ( \35726 , RIbe28390_19);
not \U$35474 ( \35727 , \15313 );
or \U$35475 ( \35728 , \35726 , \35727 );
nand \U$35476 ( \35729 , \6634 , RIbe28b10_35);
nand \U$35477 ( \35730 , \35728 , \35729 );
not \U$35478 ( \35731 , \35730 );
not \U$35479 ( \35732 , \10984 );
and \U$35480 ( \35733 , \35731 , \35732 );
and \U$35481 ( \35734 , \35730 , \8252 );
nor \U$35482 ( \35735 , \35733 , \35734 );
not \U$35483 ( \35736 , \35735 );
not \U$35484 ( \35737 , \35736 );
or \U$35485 ( \35738 , \35725 , \35737 );
not \U$35486 ( \35739 , \35724 );
nand \U$35487 ( \35740 , \35735 , \35739 );
nand \U$35488 ( \35741 , \35738 , \35740 );
not \U$35489 ( \35742 , RIbe285e8_24);
not \U$35490 ( \35743 , \4804 );
or \U$35491 ( \35744 , \35742 , \35743 );
nand \U$35492 ( \35745 , \6418 , RIbe287c8_28);
nand \U$35493 ( \35746 , \35744 , \35745 );
xor \U$35494 ( \35747 , \35746 , \4323 );
and \U$35495 ( \35748 , \35741 , \35747 );
not \U$35496 ( \35749 , \35741 );
xnor \U$35497 ( \35750 , \35746 , \4323 );
and \U$35498 ( \35751 , \35749 , \35750 );
nor \U$35499 ( \35752 , \35748 , \35751 );
buf \U$35500 ( \35753 , \35752 );
and \U$35501 ( \35754 , \35715 , \35753 );
not \U$35502 ( \35755 , \35715 );
not \U$35503 ( \35756 , \35753 );
and \U$35504 ( \35757 , \35755 , \35756 );
nor \U$35505 ( \35758 , \35754 , \35757 );
not \U$35506 ( \35759 , \35758 );
xor \U$35507 ( \35760 , \35637 , \35759 );
and \U$35508 ( \35761 , \12704 , RIbe28de0_41);
or \U$35509 ( \35762 , \13728 , \35761 );
nand \U$35510 ( \35763 , \13728 , \1636 );
nand \U$35511 ( \35764 , \35762 , \35763 );
and \U$35512 ( \35765 , \35764 , \12723 );
not \U$35513 ( \35766 , \35764 );
and \U$35514 ( \35767 , \35766 , \12879 );
nor \U$35515 ( \35768 , \35765 , \35767 );
not \U$35516 ( \35769 , \13087 );
not \U$35517 ( \35770 , \3299 );
and \U$35518 ( \35771 , \35769 , \35770 );
and \U$35519 ( \35772 , \14726 , RIbe27c10_3);
nor \U$35520 ( \35773 , \35771 , \35772 );
and \U$35521 ( \35774 , \35773 , \12770 );
not \U$35522 ( \35775 , \35773 );
and \U$35523 ( \35776 , \35775 , \12927 );
nor \U$35524 ( \35777 , \35774 , \35776 );
xor \U$35525 ( \35778 , \35768 , \35777 );
nand \U$35526 ( \35779 , \13074 , RIbe27b98_2);
and \U$35527 ( \35780 , \35779 , \12743 );
not \U$35528 ( \35781 , \35779 );
and \U$35529 ( \35782 , \35781 , \12746 );
nor \U$35530 ( \35783 , \35780 , \35782 );
and \U$35531 ( \35784 , \35778 , \35783 );
not \U$35532 ( \35785 , \35778 );
not \U$35533 ( \35786 , \35783 );
and \U$35534 ( \35787 , \35785 , \35786 );
nor \U$35535 ( \35788 , \35784 , \35787 );
not \U$35536 ( \35789 , \35788 );
not \U$35537 ( \35790 , \35789 );
not \U$35538 ( \35791 , RIbe290b0_47);
not \U$35539 ( \35792 , \10936 );
or \U$35540 ( \35793 , \35791 , \35792 );
nand \U$35541 ( \35794 , \12971 , RIbe29a88_68);
nand \U$35542 ( \35795 , \35793 , \35794 );
not \U$35543 ( \35796 , \35795 );
not \U$35544 ( \35797 , \9903 );
and \U$35545 ( \35798 , \35796 , \35797 );
and \U$35546 ( \35799 , \35795 , \10940 );
nor \U$35547 ( \35800 , \35798 , \35799 );
and \U$35548 ( \35801 , \13049 , RIbe27d78_6);
and \U$35549 ( \35802 , \12947 , RIbe27d00_5);
nor \U$35550 ( \35803 , \35801 , \35802 );
and \U$35551 ( \35804 , \35803 , \12956 );
not \U$35552 ( \35805 , \35803 );
and \U$35553 ( \35806 , \35805 , \12195 );
nor \U$35554 ( \35807 , \35804 , \35806 );
xor \U$35555 ( \35808 , \35800 , \35807 );
and \U$35556 ( \35809 , \10915 , RIbe29038_46);
and \U$35557 ( \35810 , \14771 , RIbe28fc0_45);
nor \U$35558 ( \35811 , \35809 , \35810 );
and \U$35559 ( \35812 , \35811 , \13384 );
not \U$35560 ( \35813 , \35811 );
and \U$35561 ( \35814 , \35813 , \13650 );
nor \U$35562 ( \35815 , \35812 , \35814 );
xor \U$35563 ( \35816 , \35808 , \35815 );
not \U$35564 ( \35817 , \35816 );
not \U$35565 ( \35818 , \35817 );
or \U$35566 ( \35819 , \35790 , \35818 );
nand \U$35567 ( \35820 , \35816 , \35788 );
nand \U$35568 ( \35821 , \35819 , \35820 );
not \U$35569 ( \35822 , \6985 );
not \U$35570 ( \35823 , \35822 );
not \U$35571 ( \35824 , \28330 );
and \U$35572 ( \35825 , \35823 , \35824 );
and \U$35573 ( \35826 , \7299 , RIbe280c0_13);
nor \U$35574 ( \35827 , \35825 , \35826 );
and \U$35575 ( \35828 , \35827 , \13227 );
not \U$35576 ( \35829 , \35827 );
and \U$35577 ( \35830 , \35829 , \13168 );
nor \U$35578 ( \35831 , \35828 , \35830 );
not \U$35579 ( \35832 , \35831 );
not \U$35580 ( \35833 , \35832 );
not \U$35581 ( \35834 , RIbe296c8_60);
not \U$35582 ( \35835 , \7975 );
or \U$35583 ( \35836 , \35834 , \35835 );
nand \U$35584 ( \35837 , \7981 , RIbe29650_59);
nand \U$35585 ( \35838 , \35836 , \35837 );
and \U$35586 ( \35839 , \35838 , \6950 );
not \U$35587 ( \35840 , \35838 );
and \U$35588 ( \35841 , \35840 , \7984 );
nor \U$35589 ( \35842 , \35839 , \35841 );
not \U$35590 ( \35843 , \35842 );
not \U$35591 ( \35844 , \35843 );
or \U$35592 ( \35845 , \35833 , \35844 );
nand \U$35593 ( \35846 , \35842 , \35831 );
nand \U$35594 ( \35847 , \35845 , \35846 );
not \U$35595 ( \35848 , RIbe28228_16);
not \U$35596 ( \35849 , \13327 );
or \U$35597 ( \35850 , \35848 , \35849 );
nand \U$35598 ( \35851 , \6963 , RIbe281b0_15);
nand \U$35599 ( \35852 , \35850 , \35851 );
and \U$35600 ( \35853 , \35852 , \6572 );
not \U$35601 ( \35854 , \35852 );
and \U$35602 ( \35855 , \35854 , \7293 );
nor \U$35603 ( \35856 , \35853 , \35855 );
xor \U$35604 ( \35857 , \35847 , \35856 );
not \U$35605 ( \35858 , \35857 );
and \U$35606 ( \35859 , \35821 , \35858 );
not \U$35607 ( \35860 , \35821 );
and \U$35608 ( \35861 , \35860 , \35857 );
nor \U$35609 ( \35862 , \35859 , \35861 );
not \U$35610 ( \35863 , \35862 );
nand \U$35611 ( \35864 , \34741 , \34709 );
and \U$35612 ( \35865 , \35864 , \34675 );
nor \U$35613 ( \35866 , \34709 , \34741 );
nor \U$35614 ( \35867 , \35865 , \35866 );
not \U$35615 ( \35868 , \35867 );
or \U$35616 ( \35869 , \35863 , \35868 );
not \U$35617 ( \35870 , \35862 );
not \U$35618 ( \35871 , \35867 );
nand \U$35619 ( \35872 , \35870 , \35871 );
nand \U$35620 ( \35873 , \35869 , \35872 );
xnor \U$35621 ( \35874 , \35760 , \35873 );
xnor \U$35622 ( \35875 , \35621 , \35874 );
xor \U$35623 ( \35876 , \35404 , \35875 );
not \U$35624 ( \35877 , \33696 );
not \U$35625 ( \35878 , \33674 );
or \U$35626 ( \35879 , \35877 , \35878 );
or \U$35627 ( \35880 , \33674 , \33696 );
nand \U$35628 ( \35881 , \35880 , \33668 );
nand \U$35629 ( \35882 , \35879 , \35881 );
xor \U$35630 ( \35883 , \34321 , \34325 );
and \U$35631 ( \35884 , \35883 , \34392 );
and \U$35632 ( \35885 , \34321 , \34325 );
or \U$35633 ( \35886 , \35884 , \35885 );
xor \U$35634 ( \35887 , \35882 , \35886 );
not \U$35635 ( \35888 , \34764 );
nand \U$35636 ( \35889 , \34747 , \35888 );
and \U$35637 ( \35890 , \35889 , \34603 );
nor \U$35638 ( \35891 , \34747 , \35888 );
nor \U$35639 ( \35892 , \35890 , \35891 );
not \U$35640 ( \35893 , \35892 );
xnor \U$35641 ( \35894 , \35887 , \35893 );
xor \U$35642 ( \35895 , \35876 , \35894 );
xor \U$35643 ( \35896 , \35386 , \35895 );
nand \U$35644 ( \35897 , \34732 , \34723 );
and \U$35645 ( \35898 , \35897 , \34740 );
nor \U$35646 ( \35899 , \34723 , \34732 );
nor \U$35647 ( \35900 , \35898 , \35899 );
not \U$35648 ( \35901 , \35900 );
not \U$35649 ( \35902 , \34414 );
not \U$35650 ( \35903 , \34428 );
or \U$35651 ( \35904 , \35902 , \35903 );
nand \U$35652 ( \35905 , \35904 , \34403 );
not \U$35653 ( \35906 , \34414 );
nand \U$35654 ( \35907 , \35906 , \34431 );
nand \U$35655 ( \35908 , \35905 , \35907 );
nand \U$35656 ( \35909 , \34442 , \34468 );
and \U$35657 ( \35910 , \35909 , \34454 );
nor \U$35658 ( \35911 , \34442 , \34468 );
nor \U$35659 ( \35912 , \35910 , \35911 );
and \U$35660 ( \35913 , \35908 , \35912 );
not \U$35661 ( \35914 , \35908 );
not \U$35662 ( \35915 , \35912 );
and \U$35663 ( \35916 , \35914 , \35915 );
nor \U$35664 ( \35917 , \35913 , \35916 );
xor \U$35665 ( \35918 , \35901 , \35917 );
nand \U$35666 ( \35919 , \34370 , \34387 );
and \U$35667 ( \35920 , \35919 , \34340 );
nor \U$35668 ( \35921 , \34370 , \34387 );
nor \U$35669 ( \35922 , \35920 , \35921 );
xor \U$35670 ( \35923 , \35918 , \35922 );
nand \U$35671 ( \35924 , \34506 , \34513 );
and \U$35672 ( \35925 , \35924 , \34602 );
nor \U$35673 ( \35926 , \34506 , \34513 );
nor \U$35674 ( \35927 , \35925 , \35926 );
xor \U$35675 ( \35928 , \35923 , \35927 );
not \U$35676 ( \35929 , \33275 );
not \U$35677 ( \35930 , \33663 );
or \U$35678 ( \35931 , \35929 , \35930 );
not \U$35679 ( \35932 , \33660 );
nand \U$35680 ( \35933 , \33662 , \33273 , \33274 );
or \U$35681 ( \35934 , \35932 , \35933 );
nand \U$35682 ( \35935 , \35934 , \32828 );
nand \U$35683 ( \35936 , \35931 , \35935 );
xor \U$35684 ( \35937 , \35928 , \35936 );
xor \U$35685 ( \35938 , \34317 , \34393 );
and \U$35686 ( \35939 , \35938 , \34772 );
and \U$35687 ( \35940 , \34317 , \34393 );
or \U$35688 ( \35941 , \35939 , \35940 );
not \U$35689 ( \35942 , \35941 );
xnor \U$35690 ( \35943 , \35937 , \35942 );
xor \U$35691 ( \35944 , \35896 , \35943 );
not \U$35692 ( \35945 , \35944 );
and \U$35693 ( \35946 , \35380 , \35945 );
and \U$35694 ( \35947 , \35379 , \34294 );
nor \U$35695 ( \35948 , \35946 , \35947 );
not \U$35696 ( \35949 , \35948 );
not \U$35697 ( \35950 , \35882 );
not \U$35698 ( \35951 , \35893 );
or \U$35699 ( \35952 , \35950 , \35951 );
not \U$35700 ( \35953 , \35882 );
not \U$35701 ( \35954 , \35953 );
not \U$35702 ( \35955 , \35892 );
or \U$35703 ( \35956 , \35954 , \35955 );
nand \U$35704 ( \35957 , \35956 , \35886 );
nand \U$35705 ( \35958 , \35952 , \35957 );
nand \U$35706 ( \35959 , \35758 , \35867 );
and \U$35707 ( \35960 , \35959 , \35862 );
nor \U$35708 ( \35961 , \35758 , \35867 );
nor \U$35709 ( \35962 , \35960 , \35961 );
not \U$35710 ( \35963 , \35962 );
nand \U$35711 ( \35964 , \35600 , \35586 );
not \U$35712 ( \35965 , \35964 );
not \U$35713 ( \35966 , \35591 );
or \U$35714 ( \35967 , \35965 , \35966 );
not \U$35715 ( \35968 , \35600 );
nand \U$35716 ( \35969 , \35968 , \35585 );
nand \U$35717 ( \35970 , \35967 , \35969 );
not \U$35718 ( \35971 , \35608 );
not \U$35719 ( \35972 , \35612 );
or \U$35720 ( \35973 , \35971 , \35972 );
nand \U$35721 ( \35974 , \35973 , \35618 );
not \U$35722 ( \35975 , \35608 );
nand \U$35723 ( \35976 , \35975 , \35613 );
nand \U$35724 ( \35977 , \35974 , \35976 );
xor \U$35725 ( \35978 , \35970 , \35977 );
not \U$35726 ( \35979 , \35978 );
or \U$35727 ( \35980 , \35963 , \35979 );
not \U$35728 ( \35981 , \35978 );
not \U$35729 ( \35982 , \35962 );
nand \U$35730 ( \35983 , \35981 , \35982 );
nand \U$35731 ( \35984 , \35980 , \35983 );
not \U$35732 ( \35985 , \35454 );
not \U$35733 ( \35986 , \35438 );
or \U$35734 ( \35987 , \35985 , \35986 );
nand \U$35735 ( \35988 , \35987 , \35445 );
nand \U$35736 ( \35989 , \35437 , \35457 );
and \U$35737 ( \35990 , \35988 , \35989 );
not \U$35738 ( \35991 , \35990 );
not \U$35739 ( \35992 , \35912 );
not \U$35740 ( \35993 , \35900 );
or \U$35741 ( \35994 , \35992 , \35993 );
nand \U$35742 ( \35995 , \35994 , \35908 );
nand \U$35743 ( \35996 , \35915 , \35901 );
nand \U$35744 ( \35997 , \35995 , \35996 );
not \U$35745 ( \35998 , \35997 );
not \U$35746 ( \35999 , \35636 );
not \U$35747 ( \36000 , \35625 );
or \U$35748 ( \36001 , \35999 , \36000 );
nand \U$35749 ( \36002 , \36001 , \35631 );
or \U$35750 ( \36003 , \35625 , \35636 );
nand \U$35751 ( \36004 , \36002 , \36003 );
not \U$35752 ( \36005 , \36004 );
not \U$35753 ( \36006 , \36005 );
or \U$35754 ( \36007 , \35998 , \36006 );
or \U$35755 ( \36008 , \36005 , \35997 );
nand \U$35756 ( \36009 , \36007 , \36008 );
not \U$35757 ( \36010 , \36009 );
or \U$35758 ( \36011 , \35991 , \36010 );
or \U$35759 ( \36012 , \36009 , \35990 );
nand \U$35760 ( \36013 , \36011 , \36012 );
not \U$35761 ( \36014 , RIbe29a88_68);
not \U$35762 ( \36015 , \13024 );
or \U$35763 ( \36016 , \36014 , \36015 );
nand \U$35764 ( \36017 , \14511 , RIbe27d78_6);
nand \U$35765 ( \36018 , \36016 , \36017 );
not \U$35766 ( \36019 , \36018 );
not \U$35767 ( \36020 , \12218 );
and \U$35768 ( \36021 , \36019 , \36020 );
and \U$35769 ( \36022 , \36018 , \13033 );
nor \U$35770 ( \36023 , \36021 , \36022 );
not \U$35771 ( \36024 , RIbe27d00_5);
not \U$35772 ( \36025 , \12942 );
or \U$35773 ( \36026 , \36024 , \36025 );
nand \U$35774 ( \36027 , \13669 , RIbe27c10_3);
nand \U$35775 ( \36028 , \36026 , \36027 );
and \U$35776 ( \36029 , \36028 , \12195 );
not \U$35777 ( \36030 , \36028 );
and \U$35778 ( \36031 , \36030 , \12957 );
nor \U$35779 ( \36032 , \36029 , \36031 );
xnor \U$35780 ( \36033 , \36023 , \36032 );
and \U$35781 ( \36034 , \8278 , RIbe28fc0_45);
and \U$35782 ( \36035 , \13643 , RIbe290b0_47);
nor \U$35783 ( \36036 , \36034 , \36035 );
and \U$35784 ( \36037 , \36036 , \13646 );
not \U$35785 ( \36038 , \36036 );
and \U$35786 ( \36039 , \36038 , \8077 );
nor \U$35787 ( \36040 , \36037 , \36039 );
buf \U$35788 ( \36041 , \36040 );
not \U$35789 ( \36042 , \36041 );
and \U$35790 ( \36043 , \36033 , \36042 );
not \U$35791 ( \36044 , \36033 );
and \U$35792 ( \36045 , \36044 , \36041 );
nor \U$35793 ( \36046 , \36043 , \36045 );
not \U$35794 ( \36047 , \36046 );
not \U$35795 ( \36048 , RIbe28e58_42);
not \U$35796 ( \36049 , \15615 );
or \U$35797 ( \36050 , \36048 , \36049 );
nand \U$35798 ( \36051 , \14491 , RIbe28de0_41);
nand \U$35799 ( \36052 , \36050 , \36051 );
not \U$35800 ( \36053 , \36052 );
not \U$35801 ( \36054 , \14000 );
and \U$35802 ( \36055 , \36053 , \36054 );
and \U$35803 ( \36056 , \36052 , \26172 );
nor \U$35804 ( \36057 , \36055 , \36056 );
xor \U$35805 ( \36058 , \15166 , \36057 );
not \U$35806 ( \36059 , RIbe29920_65);
not \U$35807 ( \36060 , \12707 );
or \U$35808 ( \36061 , \36059 , \36060 );
nand \U$35809 ( \36062 , \12711 , RIbe27b98_2);
nand \U$35810 ( \36063 , \36061 , \36062 );
xnor \U$35811 ( \36064 , \36063 , \13068 );
xor \U$35812 ( \36065 , \36058 , \36064 );
not \U$35813 ( \36066 , \36065 );
or \U$35814 ( \36067 , \36047 , \36066 );
or \U$35815 ( \36068 , \36046 , \36065 );
nand \U$35816 ( \36069 , \36067 , \36068 );
not \U$35817 ( \36070 , \36069 );
not \U$35818 ( \36071 , \36070 );
not \U$35819 ( \36072 , \35817 );
not \U$35820 ( \36073 , \35857 );
or \U$35821 ( \36074 , \36072 , \36073 );
not \U$35822 ( \36075 , \35788 );
nand \U$35823 ( \36076 , \36074 , \36075 );
not \U$35824 ( \36077 , \35817 );
nand \U$35825 ( \36078 , \36077 , \35858 );
nand \U$35826 ( \36079 , \36076 , \36078 );
not \U$35827 ( \36080 , \36079 );
or \U$35828 ( \36081 , \36071 , \36080 );
nand \U$35829 ( \36082 , \36069 , \36076 , \36078 );
nand \U$35830 ( \36083 , \36081 , \36082 );
xor \U$35831 ( \36084 , \36013 , \36083 );
not \U$35832 ( \36085 , \35670 );
not \U$35833 ( \36086 , \35752 );
or \U$35834 ( \36087 , \36085 , \36086 );
nand \U$35835 ( \36088 , \36087 , \35711 );
not \U$35836 ( \36089 , \35752 );
nand \U$35837 ( \36090 , \36089 , \35669 );
nand \U$35838 ( \36091 , \36088 , \36090 );
xor \U$35839 ( \36092 , \35428 , \36091 );
not \U$35840 ( \36093 , \35530 );
nand \U$35841 ( \36094 , \36093 , \35494 );
not \U$35842 ( \36095 , \35493 );
not \U$35843 ( \36096 , \35530 );
or \U$35844 ( \36097 , \36095 , \36096 );
nand \U$35845 ( \36098 , \36097 , \35562 );
nand \U$35846 ( \36099 , \36094 , \36098 );
xor \U$35847 ( \36100 , \36092 , \36099 );
xor \U$35848 ( \36101 , \36084 , \36100 );
xor \U$35849 ( \36102 , \35984 , \36101 );
not \U$35850 ( \36103 , \35459 );
not \U$35851 ( \36104 , \36103 );
not \U$35852 ( \36105 , \35431 );
or \U$35853 ( \36106 , \36104 , \36105 );
or \U$35854 ( \36107 , \36103 , \35431 );
nand \U$35855 ( \36108 , \36107 , \35571 );
nand \U$35856 ( \36109 , \36106 , \36108 );
not \U$35857 ( \36110 , \36109 );
not \U$35858 ( \36111 , \36110 );
not \U$35859 ( \36112 , \35525 );
not \U$35860 ( \36113 , \35513 );
or \U$35861 ( \36114 , \36112 , \36113 );
nand \U$35862 ( \36115 , \36114 , \35502 );
not \U$35863 ( \36116 , \35525 );
nand \U$35864 ( \36117 , \36116 , \35514 );
nand \U$35865 ( \36118 , \36115 , \36117 );
xor \U$35866 ( \36119 , \35540 , \35550 );
and \U$35867 ( \36120 , \36119 , \35561 );
and \U$35868 ( \36121 , \35540 , \35550 );
or \U$35869 ( \36122 , \36120 , \36121 );
xor \U$35870 ( \36123 , \36118 , \36122 );
nand \U$35871 ( \36124 , \35492 , \35472 );
and \U$35872 ( \36125 , \36124 , \35481 );
nor \U$35873 ( \36126 , \35492 , \35472 );
nor \U$35874 ( \36127 , \36125 , \36126 );
xor \U$35875 ( \36128 , \36123 , \36127 );
not \U$35876 ( \36129 , \35647 );
nand \U$35877 ( \36130 , \36129 , \35658 );
not \U$35878 ( \36131 , \36130 );
not \U$35879 ( \36132 , \35668 );
or \U$35880 ( \36133 , \36131 , \36132 );
not \U$35881 ( \36134 , \35658 );
nand \U$35882 ( \36135 , \36134 , \35647 );
nand \U$35883 ( \36136 , \36133 , \36135 );
or \U$35884 ( \36137 , \35705 , \35681 );
not \U$35885 ( \36138 , \35692 );
nand \U$35886 ( \36139 , \36137 , \36138 );
nand \U$35887 ( \36140 , \35705 , \35681 );
nand \U$35888 ( \36141 , \36139 , \36140 );
xor \U$35889 ( \36142 , \36136 , \36141 );
not \U$35890 ( \36143 , \35750 );
not \U$35891 ( \36144 , \35739 );
or \U$35892 ( \36145 , \36143 , \36144 );
not \U$35893 ( \36146 , \35724 );
not \U$35894 ( \36147 , \35747 );
or \U$35895 ( \36148 , \36146 , \36147 );
nand \U$35896 ( \36149 , \36148 , \35736 );
nand \U$35897 ( \36150 , \36145 , \36149 );
xnor \U$35898 ( \36151 , \36142 , \36150 );
xor \U$35899 ( \36152 , \36128 , \36151 );
nand \U$35900 ( \36153 , \35815 , \35800 );
buf \U$35901 ( \36154 , \35807 );
and \U$35902 ( \36155 , \36153 , \36154 );
nor \U$35903 ( \36156 , \35815 , \35800 );
nor \U$35904 ( \36157 , \36155 , \36156 );
not \U$35905 ( \36158 , \36157 );
not \U$35906 ( \36159 , \35768 );
not \U$35907 ( \36160 , \36159 );
not \U$35908 ( \36161 , \35783 );
or \U$35909 ( \36162 , \36160 , \36161 );
nand \U$35910 ( \36163 , \36162 , \35777 );
nand \U$35911 ( \36164 , \35786 , \35768 );
nand \U$35912 ( \36165 , \36163 , \36164 );
not \U$35913 ( \36166 , \36165 );
or \U$35914 ( \36167 , \36158 , \36166 );
or \U$35915 ( \36168 , \36157 , \36165 );
nand \U$35916 ( \36169 , \36167 , \36168 );
not \U$35917 ( \36170 , \36169 );
and \U$35918 ( \36171 , \35856 , \35843 );
nor \U$35919 ( \36172 , \36171 , \35831 );
nor \U$35920 ( \36173 , \35856 , \35843 );
nor \U$35921 ( \36174 , \36172 , \36173 );
not \U$35922 ( \36175 , \36174 );
and \U$35923 ( \36176 , \36170 , \36175 );
and \U$35924 ( \36177 , \36169 , \36174 );
nor \U$35925 ( \36178 , \36176 , \36177 );
xor \U$35926 ( \36179 , \36152 , \36178 );
not \U$35927 ( \36180 , \36179 );
not \U$35928 ( \36181 , \36180 );
or \U$35929 ( \36182 , \36111 , \36181 );
nand \U$35930 ( \36183 , \36179 , \36109 );
nand \U$35931 ( \36184 , \36182 , \36183 );
xor \U$35932 ( \36185 , \35410 , \35417 );
and \U$35933 ( \36186 , \36185 , \35425 );
and \U$35934 ( \36187 , \35410 , \35417 );
or \U$35935 ( \36188 , \36186 , \36187 );
not \U$35936 ( \36189 , RIbe2a5c8_92);
not \U$35937 ( \36190 , \9239 );
or \U$35938 ( \36191 , \36189 , \36190 );
not \U$35939 ( \36192 , \21491 );
nand \U$35940 ( \36193 , \36192 , \428 );
nand \U$35941 ( \36194 , \36191 , \36193 );
and \U$35942 ( \36195 , \36194 , \306 );
not \U$35943 ( \36196 , \36194 );
and \U$35944 ( \36197 , \36196 , \312 );
nor \U$35945 ( \36198 , \36195 , \36197 );
not \U$35946 ( \36199 , \36198 );
and \U$35947 ( \36200 , \546 , RIbe2a988_100);
and \U$35948 ( \36201 , \552 , RIbe2a910_99);
nor \U$35949 ( \36202 , \36200 , \36201 );
not \U$35950 ( \36203 , \36202 );
not \U$35951 ( \36204 , \1761 );
and \U$35952 ( \36205 , \36203 , \36204 );
and \U$35953 ( \36206 , \1245 , \36202 );
nor \U$35954 ( \36207 , \36205 , \36206 );
not \U$35955 ( \36208 , \36207 );
or \U$35956 ( \36209 , \36199 , \36208 );
or \U$35957 ( \36210 , \36207 , \36198 );
nand \U$35958 ( \36211 , \36209 , \36210 );
and \U$35959 ( \36212 , \5365 , RIbe2a208_84);
and \U$35960 ( \36213 , \1256 , RIbe2a190_83);
nor \U$35961 ( \36214 , \36212 , \36213 );
and \U$35962 ( \36215 , \36214 , \300 );
not \U$35963 ( \36216 , \36214 );
and \U$35964 ( \36217 , \36216 , \293 );
nor \U$35965 ( \36218 , \36215 , \36217 );
and \U$35966 ( \36219 , \36211 , \36218 );
not \U$35967 ( \36220 , \36211 );
not \U$35968 ( \36221 , \36218 );
and \U$35969 ( \36222 , \36220 , \36221 );
nor \U$35970 ( \36223 , \36219 , \36222 );
xor \U$35971 ( \36224 , \36188 , \36223 );
nand \U$35972 ( \36225 , RIbe29380_53, RIbe2b180_117);
not \U$35973 ( \36226 , RIbe2b270_119);
not \U$35974 ( \36227 , \12312 );
or \U$35975 ( \36228 , \36226 , \36227 );
nand \U$35976 ( \36229 , \329 , RIbe2b108_116);
nand \U$35977 ( \36230 , \36228 , \36229 );
not \U$35978 ( \36231 , \36230 );
not \U$35979 ( \36232 , \12321 );
and \U$35980 ( \36233 , \36231 , \36232 );
and \U$35981 ( \36234 , \36230 , \12321 );
nor \U$35982 ( \36235 , \36233 , \36234 );
xor \U$35983 ( \36236 , \36225 , \36235 );
not \U$35984 ( \36237 , RIbe2b090_115);
not \U$35985 ( \36238 , \260 );
or \U$35986 ( \36239 , \36237 , \36238 );
nand \U$35987 ( \36240 , \263 , RIbe2a280_85);
nand \U$35988 ( \36241 , \36239 , \36240 );
xnor \U$35989 ( \36242 , \36241 , \1362 );
xnor \U$35990 ( \36243 , \36236 , \36242 );
xnor \U$35991 ( \36244 , \36224 , \36243 );
not \U$35992 ( \36245 , RIbe28660_25);
not \U$35993 ( \36246 , \7880 );
or \U$35994 ( \36247 , \36245 , \36246 );
nand \U$35995 ( \36248 , \8368 , RIbe285e8_24);
nand \U$35996 ( \36249 , \36247 , \36248 );
and \U$35997 ( \36250 , \36249 , \4821 );
not \U$35998 ( \36251 , \36249 );
and \U$35999 ( \36252 , \36251 , \3471 );
nor \U$36000 ( \36253 , \36250 , \36252 );
not \U$36001 ( \36254 , \36253 );
not \U$36002 ( \36255 , \36254 );
not \U$36003 ( \36256 , RIbe27f58_10);
not \U$36004 ( \36257 , \30862 );
or \U$36005 ( \36258 , \36256 , \36257 );
nand \U$36006 ( \36259 , RIbe27e68_8, \3689 );
nand \U$36007 ( \36260 , \36258 , \36259 );
and \U$36008 ( \36261 , \36260 , \3290 );
not \U$36009 ( \36262 , \36260 );
and \U$36010 ( \36263 , \36262 , \2887 );
nor \U$36011 ( \36264 , \36261 , \36263 );
not \U$36012 ( \36265 , \36264 );
not \U$36013 ( \36266 , \36265 );
or \U$36014 ( \36267 , \36255 , \36266 );
nand \U$36015 ( \36268 , \36253 , \36264 );
nand \U$36016 ( \36269 , \36267 , \36268 );
not \U$36017 ( \36270 , RIbe28ed0_43);
not \U$36018 ( \36271 , \7827 );
or \U$36019 ( \36272 , \36270 , \36271 );
nand \U$36020 ( \36273 , \2900 , RIbe27fd0_11);
nand \U$36021 ( \36274 , \36272 , \36273 );
not \U$36022 ( \36275 , \36274 );
not \U$36023 ( \36276 , \2379 );
and \U$36024 ( \36277 , \36275 , \36276 );
and \U$36025 ( \36278 , \36274 , \2379 );
nor \U$36026 ( \36279 , \36277 , \36278 );
not \U$36027 ( \36280 , \36279 );
and \U$36028 ( \36281 , \36269 , \36280 );
not \U$36029 ( \36282 , \36269 );
and \U$36030 ( \36283 , \36282 , \36279 );
nor \U$36031 ( \36284 , \36281 , \36283 );
not \U$36032 ( \36285 , RIbe29bf0_71);
not \U$36033 ( \36286 , \27613 );
or \U$36034 ( \36287 , \36285 , \36286 );
nand \U$36035 ( \36288 , \2384 , RIbe28f48_44);
nand \U$36036 ( \36289 , \36287 , \36288 );
not \U$36037 ( \36290 , \36289 );
not \U$36038 ( \36291 , \3516 );
and \U$36039 ( \36292 , \36290 , \36291 );
and \U$36040 ( \36293 , \36289 , \1076 );
nor \U$36041 ( \36294 , \36292 , \36293 );
not \U$36042 ( \36295 , \36294 );
not \U$36043 ( \36296 , RIbe29dd0_75);
not \U$36044 ( \36297 , \2554 );
or \U$36045 ( \36298 , \36296 , \36297 );
nand \U$36046 ( \36299 , \5467 , RIbe29c68_72);
nand \U$36047 ( \36300 , \36298 , \36299 );
and \U$36048 ( \36301 , \36300 , \1131 );
not \U$36049 ( \36302 , \36300 );
and \U$36050 ( \36303 , \36302 , \3491 );
nor \U$36051 ( \36304 , \36301 , \36303 );
not \U$36052 ( \36305 , \36304 );
or \U$36053 ( \36306 , \36295 , \36305 );
or \U$36054 ( \36307 , \36294 , \36304 );
nand \U$36055 ( \36308 , \36306 , \36307 );
not \U$36056 ( \36309 , RIbe29fb0_79);
not \U$36057 ( \36310 , \1094 );
or \U$36058 ( \36311 , \36309 , \36310 );
nand \U$36059 ( \36312 , \4730 , RIbe29e48_76);
nand \U$36060 ( \36313 , \36311 , \36312 );
and \U$36061 ( \36314 , \36313 , \5125 );
not \U$36062 ( \36315 , \36313 );
and \U$36063 ( \36316 , \36315 , \1309 );
nor \U$36064 ( \36317 , \36314 , \36316 );
not \U$36065 ( \36318 , \36317 );
and \U$36066 ( \36319 , \36308 , \36318 );
not \U$36067 ( \36320 , \36308 );
and \U$36068 ( \36321 , \36320 , \36317 );
nor \U$36069 ( \36322 , \36319 , \36321 );
xor \U$36070 ( \36323 , \36284 , \36322 );
not \U$36071 ( \36324 , \36323 );
not \U$36072 ( \36325 , RIbe2acd0_107);
not \U$36073 ( \36326 , \1142 );
or \U$36074 ( \36327 , \36325 , \36326 );
not \U$36075 ( \36328 , \14374 );
nand \U$36076 ( \36329 , \36328 , \1146 );
nand \U$36077 ( \36330 , \36327 , \36329 );
and \U$36078 ( \36331 , \36330 , \1157 );
not \U$36079 ( \36332 , \36330 );
and \U$36080 ( \36333 , \36332 , \7899 );
nor \U$36081 ( \36334 , \36331 , \36333 );
not \U$36082 ( \36335 , \36334 );
not \U$36083 ( \36336 , \36335 );
not \U$36084 ( \36337 , \6345 );
not \U$36085 ( \36338 , \13089 );
and \U$36086 ( \36339 , \36337 , \36338 );
and \U$36087 ( \36340 , \6350 , RIbe2b5b8_126);
nor \U$36088 ( \36341 , \36339 , \36340 );
and \U$36089 ( \36342 , \36341 , \4217 );
not \U$36090 ( \36343 , \36341 );
and \U$36091 ( \36344 , \36343 , \3959 );
nor \U$36092 ( \36345 , \36342 , \36344 );
not \U$36093 ( \36346 , \36345 );
not \U$36094 ( \36347 , \36346 );
or \U$36095 ( \36348 , \36336 , \36347 );
or \U$36096 ( \36349 , \36335 , \36346 );
nand \U$36097 ( \36350 , \36348 , \36349 );
and \U$36098 ( \36351 , \1002 , RIbe2a370_87);
and \U$36099 ( \36352 , \7905 , RIbe2a2f8_86);
nor \U$36100 ( \36353 , \36351 , \36352 );
and \U$36101 ( \36354 , \36353 , \1010 );
not \U$36102 ( \36355 , \36353 );
and \U$36103 ( \36356 , \36355 , \1813 );
nor \U$36104 ( \36357 , \36354 , \36356 );
buf \U$36105 ( \36358 , \36357 );
xor \U$36106 ( \36359 , \36350 , \36358 );
not \U$36107 ( \36360 , \36359 );
and \U$36108 ( \36361 , \36324 , \36360 );
and \U$36109 ( \36362 , \36359 , \36323 );
nor \U$36110 ( \36363 , \36361 , \36362 );
xor \U$36111 ( \36364 , \36244 , \36363 );
not \U$36112 ( \36365 , RIbe28408_20);
not \U$36113 ( \36366 , \5727 );
or \U$36114 ( \36367 , \36365 , \36366 );
nand \U$36115 ( \36368 , \22378 , RIbe28390_19);
nand \U$36116 ( \36369 , \36367 , \36368 );
and \U$36117 ( \36370 , \36369 , \4586 );
not \U$36118 ( \36371 , \36369 );
and \U$36119 ( \36372 , \36371 , \4592 );
nor \U$36120 ( \36373 , \36370 , \36372 );
not \U$36121 ( \36374 , RIbe28b10_35);
not \U$36122 ( \36375 , \15313 );
or \U$36123 ( \36376 , \36374 , \36375 );
nand \U$36124 ( \36377 , \10269 , RIbe28b88_36);
nand \U$36125 ( \36378 , \36376 , \36377 );
and \U$36126 ( \36379 , \36378 , \32987 );
not \U$36127 ( \36380 , \36378 );
and \U$36128 ( \36381 , \36380 , \5457 );
nor \U$36129 ( \36382 , \36379 , \36381 );
xor \U$36130 ( \36383 , \36373 , \36382 );
not \U$36131 ( \36384 , RIbe287c8_28);
not \U$36132 ( \36385 , \4804 );
or \U$36133 ( \36386 , \36384 , \36385 );
nand \U$36134 ( \36387 , \4600 , RIbe28480_21);
nand \U$36135 ( \36388 , \36386 , \36387 );
and \U$36136 ( \36389 , \36388 , \4007 );
not \U$36137 ( \36390 , \36388 );
and \U$36138 ( \36391 , \36390 , \4323 );
nor \U$36139 ( \36392 , \36389 , \36391 );
xor \U$36140 ( \36393 , \36383 , \36392 );
not \U$36141 ( \36394 , RIbe29830_63);
not \U$36142 ( \36395 , \7298 );
or \U$36143 ( \36396 , \36394 , \36395 );
nand \U$36144 ( \36397 , \6985 , RIbe296c8_60);
nand \U$36145 ( \36398 , \36396 , \36397 );
or \U$36146 ( \36399 , \36398 , \8004 );
nand \U$36147 ( \36400 , \36398 , \6992 );
nand \U$36148 ( \36401 , \36399 , \36400 );
not \U$36149 ( \36402 , RIbe29650_59);
not \U$36150 ( \36403 , \7974 );
or \U$36151 ( \36404 , \36402 , \36403 );
nand \U$36152 ( \36405 , RIbe29038_46, \7981 );
nand \U$36153 ( \36406 , \36404 , \36405 );
and \U$36154 ( \36407 , \36406 , \6948 );
not \U$36155 ( \36408 , \36406 );
and \U$36156 ( \36409 , \36408 , \7985 );
nor \U$36157 ( \36410 , \36407 , \36409 );
and \U$36158 ( \36411 , \36401 , \36410 );
not \U$36159 ( \36412 , \36401 );
not \U$36160 ( \36413 , \36410 );
and \U$36161 ( \36414 , \36412 , \36413 );
nor \U$36162 ( \36415 , \36411 , \36414 );
not \U$36163 ( \36416 , \36415 );
not \U$36164 ( \36417 , RIbe281b0_15);
not \U$36165 ( \36418 , \6958 );
or \U$36166 ( \36419 , \36417 , \36418 );
nand \U$36167 ( \36420 , \6963 , RIbe280c0_13);
nand \U$36168 ( \36421 , \36419 , \36420 );
and \U$36169 ( \36422 , \36421 , \6572 );
not \U$36170 ( \36423 , \36421 );
and \U$36171 ( \36424 , \36423 , \7293 );
nor \U$36172 ( \36425 , \36422 , \36424 );
not \U$36173 ( \36426 , \36425 );
not \U$36174 ( \36427 , \36426 );
and \U$36175 ( \36428 , \36416 , \36427 );
and \U$36176 ( \36429 , \36415 , \36426 );
nor \U$36177 ( \36430 , \36428 , \36429 );
xor \U$36178 ( \36431 , \36393 , \36430 );
and \U$36179 ( \36432 , \6536 , RIbe289a8_32);
and \U$36180 ( \36433 , \6540 , RIbe28930_31);
nor \U$36181 ( \36434 , \36432 , \36433 );
and \U$36182 ( \36435 , \36434 , \13412 );
not \U$36183 ( \36436 , \36434 );
and \U$36184 ( \36437 , \36436 , \6552 );
nor \U$36185 ( \36438 , \36435 , \36437 );
not \U$36186 ( \36439 , RIbe29560_57);
not \U$36187 ( \36440 , \13238 );
or \U$36188 ( \36441 , \36439 , \36440 );
nand \U$36189 ( \36442 , \6596 , RIbe28228_16);
nand \U$36190 ( \36443 , \36441 , \36442 );
and \U$36191 ( \36444 , \36443 , \6601 );
not \U$36192 ( \36445 , \36443 );
and \U$36193 ( \36446 , \36445 , \21238 );
nor \U$36194 ( \36447 , \36444 , \36446 );
xor \U$36195 ( \36448 , \36438 , \36447 );
not \U$36196 ( \36449 , \6141 );
not \U$36197 ( \36450 , RIbe29290_51);
not \U$36198 ( \36451 , \8231 );
or \U$36199 ( \36452 , \36450 , \36451 );
nand \U$36200 ( \36453 , \7528 , RIbe28a20_33);
nand \U$36201 ( \36454 , \36452 , \36453 );
not \U$36202 ( \36455 , \36454 );
or \U$36203 ( \36456 , \36449 , \36455 );
or \U$36204 ( \36457 , \36454 , \6141 );
nand \U$36205 ( \36458 , \36456 , \36457 );
xor \U$36206 ( \36459 , \36448 , \36458 );
and \U$36207 ( \36460 , \36431 , \36459 );
not \U$36208 ( \36461 , \36431 );
not \U$36209 ( \36462 , \36459 );
and \U$36210 ( \36463 , \36461 , \36462 );
nor \U$36211 ( \36464 , \36460 , \36463 );
xor \U$36212 ( \36465 , \36364 , \36464 );
not \U$36213 ( \36466 , \36465 );
and \U$36214 ( \36467 , \36184 , \36466 );
not \U$36215 ( \36468 , \36184 );
and \U$36216 ( \36469 , \36468 , \36465 );
nor \U$36217 ( \36470 , \36467 , \36469 );
xor \U$36218 ( \36471 , \36102 , \36470 );
xor \U$36219 ( \36472 , \35958 , \36471 );
and \U$36220 ( \36473 , \35874 , \35576 );
not \U$36221 ( \36474 , \35874 );
and \U$36222 ( \36475 , \36474 , \35577 );
nor \U$36223 ( \36476 , \36473 , \36475 );
and \U$36224 ( \36477 , \35604 , \35619 );
or \U$36225 ( \36478 , \36476 , \36477 );
or \U$36226 ( \36479 , \35619 , \35604 );
nand \U$36227 ( \36480 , \36478 , \36479 );
xor \U$36228 ( \36481 , \36472 , \36480 );
not \U$36229 ( \36482 , \36481 );
not \U$36230 ( \36483 , \36482 );
xor \U$36231 ( \36484 , \35918 , \35922 );
and \U$36232 ( \36485 , \36484 , \35927 );
and \U$36233 ( \36486 , \35918 , \35922 );
or \U$36234 ( \36487 , \36485 , \36486 );
not \U$36235 ( \36488 , \35396 );
not \U$36236 ( \36489 , \35403 );
or \U$36237 ( \36490 , \36488 , \36489 );
or \U$36238 ( \36491 , \35403 , \35396 );
nand \U$36239 ( \36492 , \36491 , \35390 );
nand \U$36240 ( \36493 , \36490 , \36492 );
not \U$36241 ( \36494 , \36493 );
xor \U$36242 ( \36495 , \36487 , \36494 );
and \U$36243 ( \36496 , \35873 , \35759 );
not \U$36244 ( \36497 , \35873 );
and \U$36245 ( \36498 , \36497 , \35758 );
nor \U$36246 ( \36499 , \36496 , \36498 );
nand \U$36247 ( \36500 , \35637 , \35576 );
and \U$36248 ( \36501 , \36499 , \36500 );
nor \U$36249 ( \36502 , \35576 , \35637 );
nor \U$36250 ( \36503 , \36501 , \36502 );
xor \U$36251 ( \36504 , \36495 , \36503 );
not \U$36252 ( \36505 , \36504 );
nand \U$36253 ( \36506 , \33663 , \33275 );
nand \U$36254 ( \36507 , \35935 , \36506 , \35928 );
not \U$36255 ( \36508 , \36507 );
not \U$36256 ( \36509 , \35941 );
or \U$36257 ( \36510 , \36508 , \36509 );
not \U$36258 ( \36511 , \35928 );
nand \U$36259 ( \36512 , \36511 , \35936 );
nand \U$36260 ( \36513 , \36510 , \36512 );
not \U$36261 ( \36514 , \36513 );
or \U$36262 ( \36515 , \36505 , \36514 );
or \U$36263 ( \36516 , \36513 , \36504 );
nand \U$36264 ( \36517 , \36515 , \36516 );
xor \U$36265 ( \36518 , \35404 , \35875 );
and \U$36266 ( \36519 , \36518 , \35894 );
and \U$36267 ( \36520 , \35404 , \35875 );
or \U$36268 ( \36521 , \36519 , \36520 );
and \U$36269 ( \36522 , \36517 , \36521 );
not \U$36270 ( \36523 , \36517 );
not \U$36271 ( \36524 , \36521 );
and \U$36272 ( \36525 , \36523 , \36524 );
nor \U$36273 ( \36526 , \36522 , \36525 );
not \U$36274 ( \36527 , \36526 );
not \U$36275 ( \36528 , \36527 );
or \U$36276 ( \36529 , \36483 , \36528 );
nand \U$36277 ( \36530 , \36526 , \36481 );
nand \U$36278 ( \36531 , \36529 , \36530 );
xor \U$36279 ( \36532 , \35386 , \35895 );
and \U$36280 ( \36533 , \36532 , \35943 );
and \U$36281 ( \36534 , \35386 , \35895 );
or \U$36282 ( \36535 , \36533 , \36534 );
not \U$36283 ( \36536 , \36535 );
not \U$36284 ( \36537 , \36536 );
and \U$36285 ( \36538 , \36531 , \36537 );
not \U$36286 ( \36539 , \36531 );
and \U$36287 ( \36540 , \36539 , \36536 );
nor \U$36288 ( \36541 , \36538 , \36540 );
not \U$36289 ( \36542 , \36541 );
not \U$36290 ( \36543 , \36542 );
or \U$36291 ( \36544 , \35949 , \36543 );
not \U$36292 ( \36545 , \35948 );
nand \U$36293 ( \36546 , \36541 , \36545 );
nand \U$36294 ( \36547 , \36544 , \36546 );
not \U$36295 ( \36548 , \36504 );
not \U$36296 ( \36549 , \36521 );
or \U$36297 ( \36550 , \36548 , \36549 );
not \U$36298 ( \36551 , \36507 );
not \U$36299 ( \36552 , \35941 );
or \U$36300 ( \36553 , \36551 , \36552 );
nand \U$36301 ( \36554 , \36553 , \36512 );
nand \U$36302 ( \36555 , \36550 , \36554 );
not \U$36303 ( \36556 , \36504 );
nand \U$36304 ( \36557 , \36556 , \36524 );
nand \U$36305 ( \36558 , \36555 , \36557 );
not \U$36306 ( \36559 , \36280 );
not \U$36307 ( \36560 , \36264 );
or \U$36308 ( \36561 , \36559 , \36560 );
not \U$36309 ( \36562 , \36265 );
not \U$36310 ( \36563 , \36279 );
or \U$36311 ( \36564 , \36562 , \36563 );
nand \U$36312 ( \36565 , \36564 , \36254 );
nand \U$36313 ( \36566 , \36561 , \36565 );
xor \U$36314 ( \36567 , \36373 , \36382 );
and \U$36315 ( \36568 , \36567 , \36392 );
and \U$36316 ( \36569 , \36373 , \36382 );
or \U$36317 ( \36570 , \36568 , \36569 );
xor \U$36318 ( \36571 , \36566 , \36570 );
xor \U$36319 ( \36572 , \36438 , \36447 );
and \U$36320 ( \36573 , \36572 , \36458 );
and \U$36321 ( \36574 , \36438 , \36447 );
or \U$36322 ( \36575 , \36573 , \36574 );
not \U$36323 ( \36576 , \36575 );
and \U$36324 ( \36577 , \36571 , \36576 );
nor \U$36325 ( \36578 , \36571 , \36576 );
nor \U$36326 ( \36579 , \36577 , \36578 );
xor \U$36327 ( \36580 , \36128 , \36151 );
and \U$36328 ( \36581 , \36580 , \36178 );
and \U$36329 ( \36582 , \36128 , \36151 );
or \U$36330 ( \36583 , \36581 , \36582 );
xor \U$36331 ( \36584 , \36579 , \36583 );
xor \U$36332 ( \36585 , \36244 , \36363 );
and \U$36333 ( \36586 , \36585 , \36464 );
and \U$36334 ( \36587 , \36244 , \36363 );
or \U$36335 ( \36588 , \36586 , \36587 );
xor \U$36336 ( \36589 , \36584 , \36588 );
xor \U$36337 ( \36590 , \36487 , \36494 );
and \U$36338 ( \36591 , \36590 , \36503 );
and \U$36339 ( \36592 , \36487 , \36494 );
or \U$36340 ( \36593 , \36591 , \36592 );
xor \U$36341 ( \36594 , \36589 , \36593 );
or \U$36342 ( \36595 , \36101 , \35984 );
and \U$36343 ( \36596 , \36595 , \36470 );
and \U$36344 ( \36597 , \35984 , \36101 );
nor \U$36345 ( \36598 , \36596 , \36597 );
xor \U$36346 ( \36599 , \36594 , \36598 );
not \U$36347 ( \36600 , \36599 );
not \U$36348 ( \36601 , \36600 );
xor \U$36349 ( \36602 , \35958 , \36471 );
and \U$36350 ( \36603 , \36602 , \36480 );
and \U$36351 ( \36604 , \35958 , \36471 );
or \U$36352 ( \36605 , \36603 , \36604 );
not \U$36353 ( \36606 , \36605 );
not \U$36354 ( \36607 , \36606 );
or \U$36355 ( \36608 , \36601 , \36607 );
nand \U$36356 ( \36609 , \36605 , \36599 );
nand \U$36357 ( \36610 , \36608 , \36609 );
not \U$36358 ( \36611 , \36046 );
nand \U$36359 ( \36612 , \36611 , \36065 );
not \U$36360 ( \36613 , \36612 );
not \U$36361 ( \36614 , \36079 );
or \U$36362 ( \36615 , \36613 , \36614 );
not \U$36363 ( \36616 , \36065 );
nand \U$36364 ( \36617 , \36616 , \36046 );
nand \U$36365 ( \36618 , \36615 , \36617 );
not \U$36366 ( \36619 , \35997 );
and \U$36367 ( \36620 , \35990 , \36619 );
nor \U$36368 ( \36621 , \36620 , \36005 );
nor \U$36369 ( \36622 , \35990 , \36619 );
nor \U$36370 ( \36623 , \36621 , \36622 );
xor \U$36371 ( \36624 , \36618 , \36623 );
xor \U$36372 ( \36625 , \35428 , \36091 );
and \U$36373 ( \36626 , \36625 , \36099 );
and \U$36374 ( \36627 , \35428 , \36091 );
or \U$36375 ( \36628 , \36626 , \36627 );
not \U$36376 ( \36629 , \36628 );
xnor \U$36377 ( \36630 , \36624 , \36629 );
not \U$36378 ( \36631 , \36118 );
nand \U$36379 ( \36632 , \36127 , \36631 );
and \U$36380 ( \36633 , \36632 , \36122 );
nor \U$36381 ( \36634 , \36127 , \36631 );
nor \U$36382 ( \36635 , \36633 , \36634 );
or \U$36383 ( \36636 , \36150 , \36141 );
and \U$36384 ( \36637 , \36636 , \36136 );
and \U$36385 ( \36638 , \36150 , \36141 );
nor \U$36386 ( \36639 , \36637 , \36638 );
xor \U$36387 ( \36640 , \36635 , \36639 );
nand \U$36388 ( \36641 , \36174 , \36157 );
and \U$36389 ( \36642 , \36641 , \36165 );
nor \U$36390 ( \36643 , \36174 , \36157 );
nor \U$36391 ( \36644 , \36642 , \36643 );
xor \U$36392 ( \36645 , \36640 , \36644 );
not \U$36393 ( \36646 , \36223 );
and \U$36394 ( \36647 , \36646 , \36188 );
nor \U$36395 ( \36648 , \36647 , \36243 );
nor \U$36396 ( \36649 , \36646 , \36188 );
nor \U$36397 ( \36650 , \36648 , \36649 );
not \U$36398 ( \36651 , \36284 );
not \U$36399 ( \36652 , \36322 );
and \U$36400 ( \36653 , \36651 , \36652 );
nor \U$36401 ( \36654 , \36653 , \36359 );
and \U$36402 ( \36655 , \36284 , \36322 );
nor \U$36403 ( \36656 , \36654 , \36655 );
not \U$36404 ( \36657 , \36656 );
not \U$36405 ( \36658 , \36657 );
xor \U$36406 ( \36659 , \36650 , \36658 );
or \U$36407 ( \36660 , \36459 , \36393 );
not \U$36408 ( \36661 , \36430 );
nand \U$36409 ( \36662 , \36660 , \36661 );
nand \U$36410 ( \36663 , \36459 , \36393 );
nand \U$36411 ( \36664 , \36662 , \36663 );
xnor \U$36412 ( \36665 , \36659 , \36664 );
xor \U$36413 ( \36666 , \36645 , \36665 );
and \U$36414 ( \36667 , \5730 , RIbe28b10_35);
not \U$36415 ( \36668 , \5730 );
and \U$36416 ( \36669 , \4826 , RIbe28390_19);
and \U$36417 ( \36670 , \36668 , \36669 );
nor \U$36418 ( \36671 , \36667 , \36670 );
and \U$36419 ( \36672 , \36671 , \20465 );
not \U$36420 ( \36673 , \36671 );
and \U$36421 ( \36674 , \36673 , \4586 );
nor \U$36422 ( \36675 , \36672 , \36674 );
not \U$36423 ( \36676 , RIbe28480_21);
not \U$36424 ( \36677 , \21040 );
or \U$36425 ( \36678 , \36676 , \36677 );
not \U$36426 ( \36679 , \4598 );
nand \U$36427 ( \36680 , \36679 , RIbe28408_20);
nand \U$36428 ( \36681 , \36678 , \36680 );
and \U$36429 ( \36682 , \36681 , \7865 );
not \U$36430 ( \36683 , \36681 );
and \U$36431 ( \36684 , \36683 , \4005 );
nor \U$36432 ( \36685 , \36682 , \36684 );
xor \U$36433 ( \36686 , \36675 , \36685 );
not \U$36434 ( \36687 , RIbe285e8_24);
not \U$36435 ( \36688 , \6783 );
or \U$36436 ( \36689 , \36687 , \36688 );
nand \U$36437 ( \36690 , \20767 , RIbe287c8_28);
nand \U$36438 ( \36691 , \36689 , \36690 );
and \U$36439 ( \36692 , \36691 , \3471 );
not \U$36440 ( \36693 , \36691 );
and \U$36441 ( \36694 , \36693 , \4821 );
nor \U$36442 ( \36695 , \36692 , \36694 );
xnor \U$36443 ( \36696 , \36686 , \36695 );
not \U$36444 ( \36697 , \6572 );
not \U$36445 ( \36698 , RIbe280c0_13);
not \U$36446 ( \36699 , \21608 );
or \U$36447 ( \36700 , \36698 , \36699 );
nand \U$36448 ( \36701 , RIbe29830_63, \6962 );
nand \U$36449 ( \36702 , \36700 , \36701 );
not \U$36450 ( \36703 , \36702 );
or \U$36451 ( \36704 , \36697 , \36703 );
or \U$36452 ( \36705 , \36702 , \6569 );
nand \U$36453 ( \36706 , \36704 , \36705 );
not \U$36454 ( \36707 , \8004 );
not \U$36455 ( \36708 , RIbe296c8_60);
not \U$36456 ( \36709 , \7298 );
or \U$36457 ( \36710 , \36708 , \36709 );
nand \U$36458 ( \36711 , \13792 , RIbe29650_59);
nand \U$36459 ( \36712 , \36710 , \36711 );
not \U$36460 ( \36713 , \36712 );
or \U$36461 ( \36714 , \36707 , \36713 );
or \U$36462 ( \36715 , \6992 , \36712 );
nand \U$36463 ( \36716 , \36714 , \36715 );
xor \U$36464 ( \36717 , \36706 , \36716 );
not \U$36465 ( \36718 , RIbe28228_16);
not \U$36466 ( \36719 , \7941 );
or \U$36467 ( \36720 , \36718 , \36719 );
nand \U$36468 ( \36721 , \6596 , RIbe281b0_15);
nand \U$36469 ( \36722 , \36720 , \36721 );
and \U$36470 ( \36723 , \36722 , \6582 );
not \U$36471 ( \36724 , \36722 );
and \U$36472 ( \36725 , \36724 , \7646 );
nor \U$36473 ( \36726 , \36723 , \36725 );
xor \U$36474 ( \36727 , \36717 , \36726 );
xor \U$36475 ( \36728 , \36696 , \36727 );
not \U$36476 ( \36729 , \6551 );
not \U$36477 ( \36730 , RIbe28930_31);
not \U$36478 ( \36731 , \6535 );
or \U$36479 ( \36732 , \36730 , \36731 );
nand \U$36480 ( \36733 , \6540 , RIbe29560_57);
nand \U$36481 ( \36734 , \36732 , \36733 );
not \U$36482 ( \36735 , \36734 );
or \U$36483 ( \36736 , \36729 , \36735 );
or \U$36484 ( \36737 , \36734 , \13412 );
nand \U$36485 ( \36738 , \36736 , \36737 );
not \U$36486 ( \36739 , \36738 );
not \U$36487 ( \36740 , RIbe28a20_33);
not \U$36488 ( \36741 , \6856 );
or \U$36489 ( \36742 , \36740 , \36741 );
nand \U$36490 ( \36743 , \6616 , RIbe289a8_32);
nand \U$36491 ( \36744 , \36742 , \36743 );
and \U$36492 ( \36745 , \36744 , \5740 );
not \U$36493 ( \36746 , \36744 );
and \U$36494 ( \36747 , \36746 , \7534 );
nor \U$36495 ( \36748 , \36745 , \36747 );
not \U$36496 ( \36749 , \36748 );
or \U$36497 ( \36750 , \36739 , \36749 );
or \U$36498 ( \36751 , \36738 , \36748 );
nand \U$36499 ( \36752 , \36750 , \36751 );
not \U$36500 ( \36753 , RIbe28b88_36);
not \U$36501 ( \36754 , \6630 );
or \U$36502 ( \36755 , \36753 , \36754 );
nand \U$36503 ( \36756 , \15885 , RIbe29290_51);
nand \U$36504 ( \36757 , \36755 , \36756 );
not \U$36505 ( \36758 , \36757 );
not \U$36506 ( \36759 , \10984 );
and \U$36507 ( \36760 , \36758 , \36759 );
and \U$36508 ( \36761 , \36757 , \6641 );
nor \U$36509 ( \36762 , \36760 , \36761 );
not \U$36510 ( \36763 , \36762 );
and \U$36511 ( \36764 , \36752 , \36763 );
not \U$36512 ( \36765 , \36752 );
and \U$36513 ( \36766 , \36765 , \36762 );
nor \U$36514 ( \36767 , \36764 , \36766 );
xor \U$36515 ( \36768 , \36728 , \36767 );
not \U$36516 ( \36769 , \36768 );
xor \U$36517 ( \36770 , \15166 , \36057 );
and \U$36518 ( \36771 , \36770 , \36064 );
and \U$36519 ( \36772 , \15166 , \36057 );
or \U$36520 ( \36773 , \36771 , \36772 );
not \U$36521 ( \36774 , \36773 );
nand \U$36522 ( \36775 , \36023 , \36040 );
and \U$36523 ( \36776 , \36775 , \36032 );
nor \U$36524 ( \36777 , \36023 , \36040 );
nor \U$36525 ( \36778 , \36776 , \36777 );
not \U$36526 ( \36779 , \36778 );
not \U$36527 ( \36780 , \36779 );
or \U$36528 ( \36781 , \36774 , \36780 );
not \U$36529 ( \36782 , \36773 );
nand \U$36530 ( \36783 , \36782 , \36778 );
nand \U$36531 ( \36784 , \36781 , \36783 );
not \U$36532 ( \36785 , \36784 );
nand \U$36533 ( \36786 , \36425 , \36410 );
not \U$36534 ( \36787 , \36786 );
not \U$36535 ( \36788 , \36401 );
or \U$36536 ( \36789 , \36787 , \36788 );
nand \U$36537 ( \36790 , \36426 , \36413 );
nand \U$36538 ( \36791 , \36789 , \36790 );
not \U$36539 ( \36792 , \36791 );
not \U$36540 ( \36793 , \36792 );
and \U$36541 ( \36794 , \36785 , \36793 );
and \U$36542 ( \36795 , \36784 , \36792 );
nor \U$36543 ( \36796 , \36794 , \36795 );
not \U$36544 ( \36797 , \36796 );
or \U$36545 ( \36798 , \36769 , \36797 );
or \U$36546 ( \36799 , \36796 , \36768 );
nand \U$36547 ( \36800 , \36798 , \36799 );
not \U$36548 ( \36801 , RIbe27c10_3);
not \U$36549 ( \36802 , \13049 );
or \U$36550 ( \36803 , \36801 , \36802 );
nand \U$36551 ( \36804 , \12948 , RIbe28e58_42);
nand \U$36552 ( \36805 , \36803 , \36804 );
and \U$36553 ( \36806 , \36805 , \12195 );
not \U$36554 ( \36807 , \36805 );
and \U$36555 ( \36808 , \36807 , \17005 );
nor \U$36556 ( \36809 , \36806 , \36808 );
not \U$36557 ( \36810 , \12752 );
not \U$36558 ( \36811 , \1636 );
and \U$36559 ( \36812 , \36810 , \36811 );
and \U$36560 ( \36813 , \14725 , RIbe28de0_41);
nor \U$36561 ( \36814 , \36812 , \36813 );
and \U$36562 ( \36815 , \36814 , \12924 );
not \U$36563 ( \36816 , \36814 );
and \U$36564 ( \36817 , \36816 , \12774 );
nor \U$36565 ( \36818 , \36815 , \36817 );
xor \U$36566 ( \36819 , \36809 , \36818 );
nand \U$36567 ( \36820 , \19262 , RIbe27b98_2);
and \U$36568 ( \36821 , \36820 , \12723 );
not \U$36569 ( \36822 , \36820 );
and \U$36570 ( \36823 , \36822 , \12879 );
nor \U$36571 ( \36824 , \36821 , \36823 );
xnor \U$36572 ( \36825 , \36819 , \36824 );
not \U$36573 ( \36826 , \36825 );
and \U$36574 ( \36827 , \10915 , RIbe290b0_47);
and \U$36575 ( \36828 , \14771 , RIbe29a88_68);
nor \U$36576 ( \36829 , \36827 , \36828 );
and \U$36577 ( \36830 , \36829 , \13650 );
not \U$36578 ( \36831 , \36829 );
and \U$36579 ( \36832 , \36831 , \7970 );
nor \U$36580 ( \36833 , \36830 , \36832 );
not \U$36581 ( \36834 , \10940 );
not \U$36582 ( \36835 , RIbe27d78_6);
not \U$36583 ( \36836 , \13024 );
or \U$36584 ( \36837 , \36835 , \36836 );
nand \U$36585 ( \36838 , \12212 , RIbe27d00_5);
nand \U$36586 ( \36839 , \36837 , \36838 );
not \U$36587 ( \36840 , \36839 );
or \U$36588 ( \36841 , \36834 , \36840 );
or \U$36589 ( \36842 , \36839 , \9903 );
nand \U$36590 ( \36843 , \36841 , \36842 );
xnor \U$36591 ( \36844 , \36833 , \36843 );
not \U$36592 ( \36845 , \6948 );
not \U$36593 ( \36846 , RIbe29038_46);
not \U$36594 ( \36847 , \10949 );
or \U$36595 ( \36848 , \36846 , \36847 );
nand \U$36596 ( \36849 , \13339 , RIbe28fc0_45);
nand \U$36597 ( \36850 , \36848 , \36849 );
not \U$36598 ( \36851 , \36850 );
or \U$36599 ( \36852 , \36845 , \36851 );
or \U$36600 ( \36853 , \36850 , \6949 );
nand \U$36601 ( \36854 , \36852 , \36853 );
buf \U$36602 ( \36855 , \36854 );
not \U$36603 ( \36856 , \36855 );
and \U$36604 ( \36857 , \36844 , \36856 );
not \U$36605 ( \36858 , \36844 );
and \U$36606 ( \36859 , \36858 , \36855 );
nor \U$36607 ( \36860 , \36857 , \36859 );
not \U$36608 ( \36861 , \36860 );
and \U$36609 ( \36862 , \36826 , \36861 );
and \U$36610 ( \36863 , \36825 , \36860 );
nor \U$36611 ( \36864 , \36862 , \36863 );
xor \U$36612 ( \36865 , \36800 , \36864 );
nand \U$36613 ( \36866 , \36235 , \36225 );
and \U$36614 ( \36867 , \36242 , \36866 );
nor \U$36615 ( \36868 , \36235 , \36225 );
nor \U$36616 ( \36869 , \36867 , \36868 );
nand \U$36617 ( \36870 , RIbe29380_53, RIbe2b270_119);
and \U$36618 ( \36871 , \324 , RIbe2b108_116);
and \U$36619 ( \36872 , \329 , RIbe2b090_115);
nor \U$36620 ( \36873 , \36871 , \36872 );
and \U$36621 ( \36874 , \36873 , \1378 );
not \U$36622 ( \36875 , \36873 );
and \U$36623 ( \36876 , \36875 , \1374 );
nor \U$36624 ( \36877 , \36874 , \36876 );
or \U$36625 ( \36878 , \36870 , \36877 );
nand \U$36626 ( \36879 , \36877 , \36870 );
nand \U$36627 ( \36880 , \36878 , \36879 );
not \U$36628 ( \36881 , \36880 );
xor \U$36629 ( \36882 , \36869 , \36881 );
and \U$36630 ( \36883 , \260 , RIbe2a280_85);
and \U$36631 ( \36884 , \264 , RIbe2a208_84);
nor \U$36632 ( \36885 , \36883 , \36884 );
and \U$36633 ( \36886 , \36885 , \270 );
not \U$36634 ( \36887 , \36885 );
and \U$36635 ( \36888 , \36887 , \1663 );
nor \U$36636 ( \36889 , \36886 , \36888 );
not \U$36637 ( \36890 , RIbe2a550_91);
not \U$36638 ( \36891 , \9239 );
or \U$36639 ( \36892 , \36890 , \36891 );
not \U$36640 ( \36893 , \13552 );
nand \U$36641 ( \36894 , \36893 , \429 );
nand \U$36642 ( \36895 , \36892 , \36894 );
and \U$36643 ( \36896 , \36895 , \3175 );
not \U$36644 ( \36897 , \36895 );
and \U$36645 ( \36898 , \36897 , \306 );
nor \U$36646 ( \36899 , \36896 , \36898 );
not \U$36647 ( \36900 , \36899 );
not \U$36648 ( \36901 , \36900 );
and \U$36649 ( \36902 , \3895 , RIbe2a190_83);
and \U$36650 ( \36903 , \9816 , RIbe2a5c8_92);
nor \U$36651 ( \36904 , \36902 , \36903 );
and \U$36652 ( \36905 , \36904 , \300 );
not \U$36653 ( \36906 , \36904 );
and \U$36654 ( \36907 , \36906 , \293 );
nor \U$36655 ( \36908 , \36905 , \36907 );
not \U$36656 ( \36909 , \36908 );
not \U$36657 ( \36910 , \36909 );
or \U$36658 ( \36911 , \36901 , \36910 );
nand \U$36659 ( \36912 , \36908 , \36899 );
nand \U$36660 ( \36913 , \36911 , \36912 );
xnor \U$36661 ( \36914 , \36889 , \36913 );
xor \U$36662 ( \36915 , \36882 , \36914 );
not \U$36663 ( \36916 , \36915 );
nand \U$36664 ( \36917 , \36334 , \36357 );
and \U$36665 ( \36918 , \36917 , \36345 );
nor \U$36666 ( \36919 , \36334 , \36357 );
nor \U$36667 ( \36920 , \36918 , \36919 );
not \U$36668 ( \36921 , \36304 );
and \U$36669 ( \36922 , \36317 , \36921 );
nor \U$36670 ( \36923 , \36922 , \36294 );
nor \U$36671 ( \36924 , \36317 , \36921 );
nor \U$36672 ( \36925 , \36923 , \36924 );
xor \U$36673 ( \36926 , \36920 , \36925 );
not \U$36674 ( \36927 , \36221 );
not \U$36675 ( \36928 , \36207 );
and \U$36676 ( \36929 , \36927 , \36928 );
and \U$36677 ( \36930 , \36221 , \36207 );
not \U$36678 ( \36931 , \36198 );
nor \U$36679 ( \36932 , \36930 , \36931 );
nor \U$36680 ( \36933 , \36929 , \36932 );
xor \U$36681 ( \36934 , \36926 , \36933 );
not \U$36682 ( \36935 , \36934 );
not \U$36683 ( \36936 , \36935 );
or \U$36684 ( \36937 , \36916 , \36936 );
not \U$36685 ( \36938 , \36915 );
nand \U$36686 ( \36939 , \36938 , \36934 );
nand \U$36687 ( \36940 , \36937 , \36939 );
not \U$36688 ( \36941 , RIbe29e48_76);
not \U$36689 ( \36942 , \1631 );
or \U$36690 ( \36943 , \36941 , \36942 );
nand \U$36691 ( \36944 , RIbe29dd0_75, \1098 );
nand \U$36692 ( \36945 , \36943 , \36944 );
and \U$36693 ( \36946 , \36945 , \1309 );
not \U$36694 ( \36947 , \36945 );
and \U$36695 ( \36948 , \36947 , \1458 );
nor \U$36696 ( \36949 , \36946 , \36948 );
not \U$36697 ( \36950 , \36949 );
not \U$36698 ( \36951 , RIbe29c68_72);
not \U$36699 ( \36952 , \1111 );
or \U$36700 ( \36953 , \36951 , \36952 );
nand \U$36701 ( \36954 , \1116 , RIbe29bf0_71);
nand \U$36702 ( \36955 , \36953 , \36954 );
not \U$36703 ( \36956 , \36955 );
not \U$36704 ( \36957 , \1123 );
and \U$36705 ( \36958 , \36956 , \36957 );
and \U$36706 ( \36959 , \1125 , \36955 );
nor \U$36707 ( \36960 , \36958 , \36959 );
not \U$36708 ( \36961 , \36960 );
or \U$36709 ( \36962 , \36950 , \36961 );
not \U$36710 ( \36963 , \36960 );
not \U$36711 ( \36964 , \36949 );
nand \U$36712 ( \36965 , \36963 , \36964 );
nand \U$36713 ( \36966 , \36962 , \36965 );
not \U$36714 ( \36967 , RIbe2a028_80);
not \U$36715 ( \36968 , \21344 );
or \U$36716 ( \36969 , \36967 , \36968 );
nand \U$36717 ( \36970 , \1146 , RIbe29fb0_79);
nand \U$36718 ( \36971 , \36969 , \36970 );
and \U$36719 ( \36972 , \36971 , \4742 );
not \U$36720 ( \36973 , \36971 );
and \U$36721 ( \36974 , \36973 , \7899 );
nor \U$36722 ( \36975 , \36972 , \36974 );
not \U$36723 ( \36976 , \36975 );
and \U$36724 ( \36977 , \36966 , \36976 );
not \U$36725 ( \36978 , \36966 );
and \U$36726 ( \36979 , \36978 , \36975 );
nor \U$36727 ( \36980 , \36977 , \36979 );
not \U$36728 ( \36981 , \36980 );
not \U$36729 ( \36982 , RIbe27e68_8);
not \U$36730 ( \36983 , \21478 );
or \U$36731 ( \36984 , \36982 , \36983 );
nand \U$36732 ( \36985 , \3456 , RIbe28660_25);
nand \U$36733 ( \36986 , \36984 , \36985 );
and \U$36734 ( \36987 , \36986 , \3290 );
not \U$36735 ( \36988 , \36986 );
and \U$36736 ( \36989 , \36988 , \2887 );
nor \U$36737 ( \36990 , \36987 , \36989 );
not \U$36738 ( \36991 , \36990 );
not \U$36739 ( \36992 , RIbe27fd0_11);
not \U$36740 ( \36993 , \29498 );
or \U$36741 ( \36994 , \36992 , \36993 );
nand \U$36742 ( \36995 , RIbe27f58_10, \2900 );
nand \U$36743 ( \36996 , \36994 , \36995 );
and \U$36744 ( \36997 , \36996 , \2379 );
not \U$36745 ( \36998 , \36996 );
and \U$36746 ( \36999 , \36998 , \2573 );
nor \U$36747 ( \37000 , \36997 , \36999 );
not \U$36748 ( \37001 , \37000 );
or \U$36749 ( \37002 , \36991 , \37001 );
or \U$36750 ( \37003 , \36990 , \37000 );
nand \U$36751 ( \37004 , \37002 , \37003 );
not \U$36752 ( \37005 , \2385 );
not \U$36753 ( \37006 , \6757 );
and \U$36754 ( \37007 , \37005 , \37006 );
and \U$36755 ( \37008 , \8833 , RIbe28f48_44);
nor \U$36756 ( \37009 , \37007 , \37008 );
and \U$36757 ( \37010 , \37009 , \1274 );
not \U$36758 ( \37011 , \37009 );
and \U$36759 ( \37012 , \37011 , \3516 );
nor \U$36760 ( \37013 , \37010 , \37012 );
and \U$36761 ( \37014 , \37004 , \37013 );
not \U$36762 ( \37015 , \37004 );
not \U$36763 ( \37016 , \37013 );
and \U$36764 ( \37017 , \37015 , \37016 );
nor \U$36765 ( \37018 , \37014 , \37017 );
not \U$36766 ( \37019 , \37018 );
or \U$36767 ( \37020 , \36981 , \37019 );
or \U$36768 ( \37021 , \37018 , \36980 );
nand \U$36769 ( \37022 , \37020 , \37021 );
not \U$36770 ( \37023 , \6345 );
not \U$36771 ( \37024 , \12917 );
and \U$36772 ( \37025 , \37023 , \37024 );
and \U$36773 ( \37026 , \664 , RIbe2a3e8_88);
nor \U$36774 ( \37027 , \37025 , \37026 );
and \U$36775 ( \37028 , \37027 , \3959 );
not \U$36776 ( \37029 , \37027 );
and \U$36777 ( \37030 , \37029 , \564 );
nor \U$36778 ( \37031 , \37028 , \37030 );
not \U$36779 ( \37032 , RIbe2a910_99);
not \U$36780 ( \37033 , \545 );
or \U$36781 ( \37034 , \37032 , \37033 );
nand \U$36782 ( \37035 , \552 , RIbe2b5b8_126);
nand \U$36783 ( \37036 , \37034 , \37035 );
not \U$36784 ( \37037 , \37036 );
not \U$36785 ( \37038 , \424 );
and \U$36786 ( \37039 , \37037 , \37038 );
and \U$36787 ( \37040 , \37036 , \424 );
nor \U$36788 ( \37041 , \37039 , \37040 );
xor \U$36789 ( \37042 , \37031 , \37041 );
not \U$36790 ( \37043 , RIbe2a2f8_86);
not \U$36791 ( \37044 , \1002 );
or \U$36792 ( \37045 , \37043 , \37044 );
nand \U$36793 ( \37046 , \1165 , RIbe2acd0_107);
nand \U$36794 ( \37047 , \37045 , \37046 );
not \U$36795 ( \37048 , \37047 );
not \U$36796 ( \37049 , \1813 );
and \U$36797 ( \37050 , \37048 , \37049 );
and \U$36798 ( \37051 , \37047 , \1608 );
nor \U$36799 ( \37052 , \37050 , \37051 );
xnor \U$36800 ( \37053 , \37042 , \37052 );
not \U$36801 ( \37054 , \37053 );
and \U$36802 ( \37055 , \37022 , \37054 );
not \U$36803 ( \37056 , \37022 );
and \U$36804 ( \37057 , \37056 , \37053 );
nor \U$36805 ( \37058 , \37055 , \37057 );
buf \U$36806 ( \37059 , \37058 );
not \U$36807 ( \37060 , \37059 );
and \U$36808 ( \37061 , \36940 , \37060 );
not \U$36809 ( \37062 , \36940 );
and \U$36810 ( \37063 , \37062 , \37059 );
nor \U$36811 ( \37064 , \37061 , \37063 );
and \U$36812 ( \37065 , \36865 , \37064 );
not \U$36813 ( \37066 , \36865 );
not \U$36814 ( \37067 , \37064 );
and \U$36815 ( \37068 , \37066 , \37067 );
nor \U$36816 ( \37069 , \37065 , \37068 );
xor \U$36817 ( \37070 , \36666 , \37069 );
xor \U$36818 ( \37071 , \36630 , \37070 );
not \U$36819 ( \37072 , \36083 );
not \U$36820 ( \37073 , \36013 );
nand \U$36821 ( \37074 , \37072 , \37073 );
and \U$36822 ( \37075 , \37074 , \36100 );
and \U$36823 ( \37076 , \36013 , \36083 );
nor \U$36824 ( \37077 , \37075 , \37076 );
or \U$36825 ( \37078 , \35977 , \35970 );
and \U$36826 ( \37079 , \37078 , \35982 );
and \U$36827 ( \37080 , \35970 , \35977 );
nor \U$36828 ( \37081 , \37079 , \37080 );
xor \U$36829 ( \37082 , \37077 , \37081 );
and \U$36830 ( \37083 , \36465 , \36110 );
buf \U$36831 ( \37084 , \36179 );
nor \U$36832 ( \37085 , \37083 , \37084 );
nor \U$36833 ( \37086 , \36465 , \36110 );
nor \U$36834 ( \37087 , \37085 , \37086 );
xor \U$36835 ( \37088 , \37082 , \37087 );
xor \U$36836 ( \37089 , \37071 , \37088 );
not \U$36837 ( \37090 , \37089 );
and \U$36838 ( \37091 , \36610 , \37090 );
not \U$36839 ( \37092 , \36610 );
and \U$36840 ( \37093 , \37092 , \37089 );
nor \U$36841 ( \37094 , \37091 , \37093 );
xor \U$36842 ( \37095 , \36558 , \37094 );
not \U$36843 ( \37096 , \36482 );
not \U$36844 ( \37097 , \36535 );
or \U$36845 ( \37098 , \37096 , \37097 );
not \U$36846 ( \37099 , \36526 );
nand \U$36847 ( \37100 , \37098 , \37099 );
not \U$36848 ( \37101 , \36482 );
nand \U$36849 ( \37102 , \37101 , \36536 );
nand \U$36850 ( \37103 , \37100 , \37102 );
xor \U$36851 ( \37104 , \37095 , \37103 );
nand \U$36852 ( \37105 , \36547 , \37104 );
xor \U$36853 ( \37106 , \36706 , \36716 );
and \U$36854 ( \37107 , \37106 , \36726 );
and \U$36855 ( \37108 , \36706 , \36716 );
or \U$36856 ( \37109 , \37107 , \37108 );
or \U$36857 ( \37110 , \36824 , \36818 );
nand \U$36858 ( \37111 , \37110 , \36809 );
nand \U$36859 ( \37112 , \36824 , \36818 );
nand \U$36860 ( \37113 , \37111 , \37112 );
not \U$36861 ( \37114 , \37113 );
xor \U$36862 ( \37115 , \37109 , \37114 );
not \U$36863 ( \37116 , \36854 );
not \U$36864 ( \37117 , \36843 );
or \U$36865 ( \37118 , \37116 , \37117 );
or \U$36866 ( \37119 , \36843 , \36854 );
nand \U$36867 ( \37120 , \37119 , \36833 );
nand \U$36868 ( \37121 , \37118 , \37120 );
xnor \U$36869 ( \37122 , \37115 , \37121 );
nand \U$36870 ( \37123 , \37058 , \36915 );
and \U$36871 ( \37124 , \37123 , \36935 );
nor \U$36872 ( \37125 , \37058 , \36915 );
nor \U$36873 ( \37126 , \37124 , \37125 );
not \U$36874 ( \37127 , \37126 );
xor \U$36875 ( \37128 , \37122 , \37127 );
and \U$36876 ( \37129 , RIbe29380_53, RIbe2b108_116);
and \U$36877 ( \37130 , \3160 , RIbe2b090_115);
and \U$36878 ( \37131 , \330 , RIbe2a280_85);
nor \U$36879 ( \37132 , \37130 , \37131 );
and \U$36880 ( \37133 , \37132 , \1374 );
not \U$36881 ( \37134 , \37132 );
and \U$36882 ( \37135 , \37134 , \1375 );
nor \U$36883 ( \37136 , \37133 , \37135 );
xor \U$36884 ( \37137 , \37129 , \37136 );
xor \U$36885 ( \37138 , \37137 , \36879 );
not \U$36886 ( \37139 , \36889 );
not \U$36887 ( \37140 , \36908 );
or \U$36888 ( \37141 , \37139 , \37140 );
or \U$36889 ( \37142 , \36889 , \36908 );
nand \U$36890 ( \37143 , \37142 , \36900 );
nand \U$36891 ( \37144 , \37141 , \37143 );
not \U$36892 ( \37145 , \37144 );
not \U$36893 ( \37146 , \37145 );
and \U$36894 ( \37147 , \36964 , \36975 );
nor \U$36895 ( \37148 , \37147 , \36960 );
nor \U$36896 ( \37149 , \36975 , \36964 );
nor \U$36897 ( \37150 , \37148 , \37149 );
nand \U$36898 ( \37151 , \37041 , \37052 );
not \U$36899 ( \37152 , \37031 );
and \U$36900 ( \37153 , \37151 , \37152 );
nor \U$36901 ( \37154 , \37041 , \37052 );
nor \U$36902 ( \37155 , \37153 , \37154 );
and \U$36903 ( \37156 , \37150 , \37155 );
not \U$36904 ( \37157 , \37150 );
not \U$36905 ( \37158 , \37155 );
and \U$36906 ( \37159 , \37157 , \37158 );
nor \U$36907 ( \37160 , \37156 , \37159 );
not \U$36908 ( \37161 , \37160 );
or \U$36909 ( \37162 , \37146 , \37161 );
or \U$36910 ( \37163 , \37160 , \37145 );
nand \U$36911 ( \37164 , \37162 , \37163 );
xor \U$36912 ( \37165 , \37138 , \37164 );
not \U$36913 ( \37166 , \36695 );
nand \U$36914 ( \37167 , \37166 , \36685 );
buf \U$36915 ( \37168 , \36675 );
and \U$36916 ( \37169 , \37167 , \37168 );
nor \U$36917 ( \37170 , \37166 , \36685 );
nor \U$36918 ( \37171 , \37169 , \37170 );
not \U$36919 ( \37172 , \37171 );
not \U$36920 ( \37173 , \37000 );
not \U$36921 ( \37174 , \37173 );
not \U$36922 ( \37175 , \36990 );
or \U$36923 ( \37176 , \37174 , \37175 );
or \U$36924 ( \37177 , \37173 , \36990 );
nand \U$36925 ( \37178 , \37177 , \37016 );
nand \U$36926 ( \37179 , \37176 , \37178 );
xor \U$36927 ( \37180 , \37172 , \37179 );
nand \U$36928 ( \37181 , \36748 , \36762 );
and \U$36929 ( \37182 , \37181 , \36738 );
nor \U$36930 ( \37183 , \36748 , \36762 );
nor \U$36931 ( \37184 , \37182 , \37183 );
and \U$36932 ( \37185 , \37180 , \37184 );
not \U$36933 ( \37186 , \37180 );
not \U$36934 ( \37187 , \37184 );
and \U$36935 ( \37188 , \37186 , \37187 );
or \U$36936 ( \37189 , \37185 , \37188 );
xor \U$36937 ( \37190 , \37165 , \37189 );
xor \U$36938 ( \37191 , \37128 , \37190 );
not \U$36939 ( \37192 , \37191 );
xor \U$36940 ( \37193 , \36635 , \36639 );
and \U$36941 ( \37194 , \37193 , \36644 );
and \U$36942 ( \37195 , \36635 , \36639 );
or \U$36943 ( \37196 , \37194 , \37195 );
not \U$36944 ( \37197 , \37196 );
not \U$36945 ( \37198 , \36650 );
not \U$36946 ( \37199 , \36656 );
or \U$36947 ( \37200 , \37198 , \37199 );
nand \U$36948 ( \37201 , \37200 , \36664 );
not \U$36949 ( \37202 , \36650 );
nand \U$36950 ( \37203 , \37202 , \36657 );
nand \U$36951 ( \37204 , \37201 , \37203 );
not \U$36952 ( \37205 , \37204 );
or \U$36953 ( \37206 , \37197 , \37205 );
or \U$36954 ( \37207 , \37204 , \37196 );
nand \U$36955 ( \37208 , \37206 , \37207 );
not \U$36956 ( \37209 , \36860 );
nand \U$36957 ( \37210 , \37209 , \36825 );
and \U$36958 ( \37211 , \37210 , \36768 );
nor \U$36959 ( \37212 , \36825 , \37209 );
nor \U$36960 ( \37213 , \37211 , \37212 );
buf \U$36961 ( \37214 , \37213 );
xnor \U$36962 ( \37215 , \37208 , \37214 );
not \U$36963 ( \37216 , \37215 );
and \U$36964 ( \37217 , \37192 , \37216 );
xor \U$36965 ( \37218 , \36920 , \36925 );
and \U$36966 ( \37219 , \37218 , \36933 );
and \U$36967 ( \37220 , \36920 , \36925 );
or \U$36968 ( \37221 , \37219 , \37220 );
buf \U$36969 ( \37222 , \37221 );
not \U$36970 ( \37223 , \37222 );
or \U$36971 ( \37224 , \36575 , \36566 );
nand \U$36972 ( \37225 , \37224 , \36570 );
nand \U$36973 ( \37226 , \36575 , \36566 );
nand \U$36974 ( \37227 , \37225 , \37226 );
not \U$36975 ( \37228 , \36773 );
not \U$36976 ( \37229 , \36778 );
or \U$36977 ( \37230 , \37228 , \37229 );
nand \U$36978 ( \37231 , \37230 , \36791 );
nand \U$36979 ( \37232 , \36779 , \36782 );
nand \U$36980 ( \37233 , \37231 , \37232 );
xor \U$36981 ( \37234 , \37227 , \37233 );
not \U$36982 ( \37235 , \37234 );
or \U$36983 ( \37236 , \37223 , \37235 );
or \U$36984 ( \37237 , \37234 , \37222 );
nand \U$36985 ( \37238 , \37236 , \37237 );
xor \U$36986 ( \37239 , \36869 , \36881 );
and \U$36987 ( \37240 , \37239 , \36914 );
and \U$36988 ( \37241 , \36869 , \36881 );
or \U$36989 ( \37242 , \37240 , \37241 );
not \U$36990 ( \37243 , \37242 );
xor \U$36991 ( \37244 , \36696 , \36727 );
and \U$36992 ( \37245 , \37244 , \36767 );
and \U$36993 ( \37246 , \36696 , \36727 );
or \U$36994 ( \37247 , \37245 , \37246 );
not \U$36995 ( \37248 , \36980 );
nand \U$36996 ( \37249 , \37248 , \37018 );
and \U$36997 ( \37250 , \37249 , \37053 );
nor \U$36998 ( \37251 , \37018 , \37248 );
nor \U$36999 ( \37252 , \37250 , \37251 );
not \U$37000 ( \37253 , \37252 );
and \U$37001 ( \37254 , \37247 , \37253 );
not \U$37002 ( \37255 , \37247 );
and \U$37003 ( \37256 , \37255 , \37252 );
nor \U$37004 ( \37257 , \37254 , \37256 );
not \U$37005 ( \37258 , \37257 );
or \U$37006 ( \37259 , \37243 , \37258 );
or \U$37007 ( \37260 , \37257 , \37242 );
nand \U$37008 ( \37261 , \37259 , \37260 );
xor \U$37009 ( \37262 , \37238 , \37261 );
not \U$37010 ( \37263 , RIbe27f58_10);
not \U$37011 ( \37264 , \29498 );
or \U$37012 ( \37265 , \37263 , \37264 );
nand \U$37013 ( \37266 , \2900 , RIbe27e68_8);
nand \U$37014 ( \37267 , \37265 , \37266 );
and \U$37015 ( \37268 , \37267 , \3272 );
not \U$37016 ( \37269 , \37267 );
and \U$37017 ( \37270 , \37269 , \2379 );
nor \U$37018 ( \37271 , \37268 , \37270 );
not \U$37019 ( \37272 , \37271 );
not \U$37020 ( \37273 , RIbe28660_25);
not \U$37021 ( \37274 , \3451 );
or \U$37022 ( \37275 , \37273 , \37274 );
nand \U$37023 ( \37276 , RIbe285e8_24, \6800 );
nand \U$37024 ( \37277 , \37275 , \37276 );
and \U$37025 ( \37278 , \37277 , \2887 );
not \U$37026 ( \37279 , \37277 );
and \U$37027 ( \37280 , \37279 , \4346 );
nor \U$37028 ( \37281 , \37278 , \37280 );
not \U$37029 ( \37282 , \37281 );
nand \U$37030 ( \37283 , \37272 , \37282 );
nand \U$37031 ( \37284 , \37281 , \37271 );
nand \U$37032 ( \37285 , \37283 , \37284 );
not \U$37033 ( \37286 , \4064 );
not \U$37034 ( \37287 , \7360 );
and \U$37035 ( \37288 , \37286 , \37287 );
and \U$37036 ( \37289 , \2390 , RIbe28ed0_43);
nor \U$37037 ( \37290 , \37288 , \37289 );
and \U$37038 ( \37291 , \37290 , \3516 );
not \U$37039 ( \37292 , \37290 );
and \U$37040 ( \37293 , \37292 , \1277 );
nor \U$37041 ( \37294 , \37291 , \37293 );
and \U$37042 ( \37295 , \37285 , \37294 );
not \U$37043 ( \37296 , \37285 );
not \U$37044 ( \37297 , \37294 );
and \U$37045 ( \37298 , \37296 , \37297 );
nor \U$37046 ( \37299 , \37295 , \37298 );
not \U$37047 ( \37300 , RIbe29290_51);
not \U$37048 ( \37301 , \5455 );
or \U$37049 ( \37302 , \37300 , \37301 );
nand \U$37050 ( \37303 , \7100 , RIbe28a20_33);
nand \U$37051 ( \37304 , \37302 , \37303 );
and \U$37052 ( \37305 , \37304 , \5754 );
not \U$37053 ( \37306 , \37304 );
and \U$37054 ( \37307 , \37306 , \6907 );
nor \U$37055 ( \37308 , \37305 , \37307 );
buf \U$37056 ( \37309 , \37308 );
not \U$37057 ( \37310 , \37309 );
not \U$37058 ( \37311 , \37310 );
not \U$37059 ( \37312 , \6541 );
not \U$37060 ( \37313 , \3952 );
and \U$37061 ( \37314 , \37312 , \37313 );
and \U$37062 ( \37315 , \6535 , RIbe29560_57);
nor \U$37063 ( \37316 , \37314 , \37315 );
and \U$37064 ( \37317 , \37316 , \6891 );
not \U$37065 ( \37318 , \37316 );
and \U$37066 ( \37319 , \37318 , \6546 );
nor \U$37067 ( \37320 , \37317 , \37319 );
not \U$37068 ( \37321 , RIbe289a8_32);
not \U$37069 ( \37322 , \13894 );
or \U$37070 ( \37323 , \37321 , \37322 );
nand \U$37071 ( \37324 , RIbe28930_31, \21084 );
nand \U$37072 ( \37325 , \37323 , \37324 );
and \U$37073 ( \37326 , \37325 , \6141 );
not \U$37074 ( \37327 , \37325 );
and \U$37075 ( \37328 , \37327 , \5741 );
nor \U$37076 ( \37329 , \37326 , \37328 );
and \U$37077 ( \37330 , \37320 , \37329 );
not \U$37078 ( \37331 , \37320 );
not \U$37079 ( \37332 , \37329 );
and \U$37080 ( \37333 , \37331 , \37332 );
nor \U$37081 ( \37334 , \37330 , \37333 );
not \U$37082 ( \37335 , \37334 );
or \U$37083 ( \37336 , \37311 , \37335 );
not \U$37084 ( \37337 , \37334 );
nand \U$37085 ( \37338 , \37337 , \37309 );
nand \U$37086 ( \37339 , \37336 , \37338 );
xor \U$37087 ( \37340 , \37299 , \37339 );
not \U$37088 ( \37341 , RIbe28408_20);
not \U$37089 ( \37342 , \4804 );
or \U$37090 ( \37343 , \37341 , \37342 );
nand \U$37091 ( \37344 , \6418 , RIbe28390_19);
nand \U$37092 ( \37345 , \37343 , \37344 );
not \U$37093 ( \37346 , \37345 );
not \U$37094 ( \37347 , \4323 );
and \U$37095 ( \37348 , \37346 , \37347 );
and \U$37096 ( \37349 , \37345 , \4323 );
nor \U$37097 ( \37350 , \37348 , \37349 );
not \U$37098 ( \37351 , RIbe28b10_35);
not \U$37099 ( \37352 , \15894 );
or \U$37100 ( \37353 , \37351 , \37352 );
nand \U$37101 ( \37354 , \22378 , RIbe28b88_36);
nand \U$37102 ( \37355 , \37353 , \37354 );
and \U$37103 ( \37356 , \37355 , \4586 );
not \U$37104 ( \37357 , \37355 );
and \U$37105 ( \37358 , \37357 , \4592 );
nor \U$37106 ( \37359 , \37356 , \37358 );
xor \U$37107 ( \37360 , \37350 , \37359 );
not \U$37108 ( \37361 , RIbe287c8_28);
not \U$37109 ( \37362 , \6783 );
or \U$37110 ( \37363 , \37361 , \37362 );
nand \U$37111 ( \37364 , \4333 , RIbe28480_21);
nand \U$37112 ( \37365 , \37363 , \37364 );
and \U$37113 ( \37366 , \37365 , \4821 );
not \U$37114 ( \37367 , \37365 );
and \U$37115 ( \37368 , \37367 , \3471 );
nor \U$37116 ( \37369 , \37366 , \37368 );
xor \U$37117 ( \37370 , \37360 , \37369 );
xor \U$37118 ( \37371 , \37340 , \37370 );
not \U$37119 ( \37372 , \37371 );
not \U$37120 ( \37373 , RIbe28e58_42);
not \U$37121 ( \37374 , \12943 );
or \U$37122 ( \37375 , \37373 , \37374 );
nand \U$37123 ( \37376 , \12947 , RIbe28de0_41);
nand \U$37124 ( \37377 , \37375 , \37376 );
not \U$37125 ( \37378 , \37377 );
not \U$37126 ( \37379 , \17005 );
and \U$37127 ( \37380 , \37378 , \37379 );
and \U$37128 ( \37381 , \37377 , \12956 );
nor \U$37129 ( \37382 , \37380 , \37381 );
not \U$37130 ( \37383 , \37382 );
xor \U$37131 ( \37384 , \12769 , \12723 );
not \U$37132 ( \37385 , \12752 );
not \U$37133 ( \37386 , \1640 );
and \U$37134 ( \37387 , \37385 , \37386 );
and \U$37135 ( \37388 , \15615 , RIbe29920_65);
nor \U$37136 ( \37389 , \37387 , \37388 );
xor \U$37137 ( \37390 , \37384 , \37389 );
not \U$37138 ( \37391 , \37390 );
and \U$37139 ( \37392 , \37383 , \37391 );
and \U$37140 ( \37393 , \37382 , \37390 );
nor \U$37141 ( \37394 , \37392 , \37393 );
not \U$37142 ( \37395 , \37394 );
not \U$37143 ( \37396 , \29757 );
not \U$37144 ( \37397 , \6984 );
not \U$37145 ( \37398 , \2355 );
and \U$37146 ( \37399 , \37397 , \37398 );
and \U$37147 ( \37400 , \7298 , RIbe29650_59);
nor \U$37148 ( \37401 , \37399 , \37400 );
not \U$37149 ( \37402 , \37401 );
or \U$37150 ( \37403 , \37396 , \37402 );
or \U$37151 ( \37404 , \37401 , \7304 );
nand \U$37152 ( \37405 , \37403 , \37404 );
not \U$37153 ( \37406 , RIbe29830_63);
not \U$37154 ( \37407 , \6958 );
or \U$37155 ( \37408 , \37406 , \37407 );
nand \U$37156 ( \37409 , \6963 , RIbe296c8_60);
nand \U$37157 ( \37410 , \37408 , \37409 );
and \U$37158 ( \37411 , \37410 , \7293 );
not \U$37159 ( \37412 , \37410 );
and \U$37160 ( \37413 , \37412 , \6572 );
nor \U$37161 ( \37414 , \37411 , \37413 );
xor \U$37162 ( \37415 , \37405 , \37414 );
not \U$37163 ( \37416 , RIbe281b0_15);
not \U$37164 ( \37417 , \7941 );
or \U$37165 ( \37418 , \37416 , \37417 );
nand \U$37166 ( \37419 , \6596 , RIbe280c0_13);
nand \U$37167 ( \37420 , \37418 , \37419 );
and \U$37168 ( \37421 , \37420 , \7948 );
not \U$37169 ( \37422 , \37420 );
and \U$37170 ( \37423 , \37422 , \7646 );
nor \U$37171 ( \37424 , \37421 , \37423 );
xor \U$37172 ( \37425 , \37415 , \37424 );
not \U$37173 ( \37426 , \37425 );
or \U$37174 ( \37427 , \37395 , \37426 );
or \U$37175 ( \37428 , \37425 , \37394 );
nand \U$37176 ( \37429 , \37427 , \37428 );
and \U$37177 ( \37430 , \10915 , RIbe29a88_68);
and \U$37178 ( \37431 , \10919 , RIbe27d78_6);
nor \U$37179 ( \37432 , \37430 , \37431 );
and \U$37180 ( \37433 , \37432 , \8077 );
not \U$37181 ( \37434 , \37432 );
and \U$37182 ( \37435 , \37434 , \16994 );
nor \U$37183 ( \37436 , \37433 , \37435 );
not \U$37184 ( \37437 , \37436 );
not \U$37185 ( \37438 , RIbe27d00_5);
not \U$37186 ( \37439 , \10936 );
or \U$37187 ( \37440 , \37438 , \37439 );
nand \U$37188 ( \37441 , \12971 , RIbe27c10_3);
nand \U$37189 ( \37442 , \37440 , \37441 );
not \U$37190 ( \37443 , \37442 );
not \U$37191 ( \37444 , \13030 );
and \U$37192 ( \37445 , \37443 , \37444 );
and \U$37193 ( \37446 , \37442 , \10940 );
nor \U$37194 ( \37447 , \37445 , \37446 );
not \U$37195 ( \37448 , \37447 );
or \U$37196 ( \37449 , \37437 , \37448 );
or \U$37197 ( \37450 , \37447 , \37436 );
nand \U$37198 ( \37451 , \37449 , \37450 );
not \U$37199 ( \37452 , RIbe28fc0_45);
not \U$37200 ( \37453 , \6942 );
or \U$37201 ( \37454 , \37452 , \37453 );
nand \U$37202 ( \37455 , \8269 , RIbe290b0_47);
nand \U$37203 ( \37456 , \37454 , \37455 );
and \U$37204 ( \37457 , \37456 , \14299 );
not \U$37205 ( \37458 , \37456 );
and \U$37206 ( \37459 , \37458 , \6948 );
nor \U$37207 ( \37460 , \37457 , \37459 );
xnor \U$37208 ( \37461 , \37451 , \37460 );
and \U$37209 ( \37462 , \37429 , \37461 );
not \U$37210 ( \37463 , \37429 );
not \U$37211 ( \37464 , \37461 );
and \U$37212 ( \37465 , \37463 , \37464 );
nor \U$37213 ( \37466 , \37462 , \37465 );
not \U$37214 ( \37467 , \37466 );
or \U$37215 ( \37468 , \37372 , \37467 );
not \U$37216 ( \37469 , \37466 );
not \U$37217 ( \37470 , \37371 );
nand \U$37218 ( \37471 , \37469 , \37470 );
nand \U$37219 ( \37472 , \37468 , \37471 );
not \U$37220 ( \37473 , RIbe2a5c8_92);
not \U$37221 ( \37474 , \32454 );
or \U$37222 ( \37475 , \37473 , \37474 );
nand \U$37223 ( \37476 , \1681 , RIbe2a550_91);
nand \U$37224 ( \37477 , \37475 , \37476 );
not \U$37225 ( \37478 , \37477 );
not \U$37226 ( \37479 , \300 );
and \U$37227 ( \37480 , \37478 , \37479 );
and \U$37228 ( \37481 , \37477 , \300 );
nor \U$37229 ( \37482 , \37480 , \37481 );
not \U$37230 ( \37483 , \37482 );
not \U$37231 ( \37484 , RIbe2a988_100);
not \U$37232 ( \37485 , \9239 );
or \U$37233 ( \37486 , \37484 , \37485 );
nand \U$37234 ( \37487 , RIbe2a910_99, \428 );
nand \U$37235 ( \37488 , \37486 , \37487 );
and \U$37236 ( \37489 , \37488 , \306 );
not \U$37237 ( \37490 , \37488 );
and \U$37238 ( \37491 , \37490 , \312 );
nor \U$37239 ( \37492 , \37489 , \37491 );
not \U$37240 ( \37493 , \37492 );
or \U$37241 ( \37494 , \37483 , \37493 );
or \U$37242 ( \37495 , \37492 , \37482 );
nand \U$37243 ( \37496 , \37494 , \37495 );
not \U$37244 ( \37497 , RIbe2a208_84);
not \U$37245 ( \37498 , \30725 );
or \U$37246 ( \37499 , \37497 , \37498 );
nand \U$37247 ( \37500 , \263 , RIbe2a190_83);
nand \U$37248 ( \37501 , \37499 , \37500 );
xor \U$37249 ( \37502 , \37501 , \1362 );
not \U$37250 ( \37503 , \37502 );
and \U$37251 ( \37504 , \37496 , \37503 );
not \U$37252 ( \37505 , \37496 );
and \U$37253 ( \37506 , \37505 , \37502 );
nor \U$37254 ( \37507 , \37504 , \37506 );
not \U$37255 ( \37508 , \37507 );
not \U$37256 ( \37509 , RIbe2acd0_107);
not \U$37257 ( \37510 , \23339 );
or \U$37258 ( \37511 , \37509 , \37510 );
nand \U$37259 ( \37512 , \1202 , RIbe2a028_80);
nand \U$37260 ( \37513 , \37511 , \37512 );
nor \U$37261 ( \37514 , \37513 , \750 );
not \U$37262 ( \37515 , \37514 );
nand \U$37263 ( \37516 , \37513 , \1813 );
nand \U$37264 ( \37517 , \37515 , \37516 );
not \U$37265 ( \37518 , RIbe2b5b8_126);
not \U$37266 ( \37519 , \546 );
or \U$37267 ( \37520 , \37518 , \37519 );
nand \U$37268 ( \37521 , \552 , RIbe2a3e8_88);
nand \U$37269 ( \37522 , \37520 , \37521 );
xor \U$37270 ( \37523 , \37522 , \424 );
xor \U$37271 ( \37524 , \37517 , \37523 );
not \U$37272 ( \37525 , \1621 );
not \U$37273 ( \37526 , \6345 );
not \U$37274 ( \37527 , \12755 );
and \U$37275 ( \37528 , \37526 , \37527 );
and \U$37276 ( \37529 , \664 , RIbe2a370_87);
nor \U$37277 ( \37530 , \37528 , \37529 );
not \U$37278 ( \37531 , \37530 );
or \U$37279 ( \37532 , \37525 , \37531 );
or \U$37280 ( \37533 , \672 , \37530 );
nand \U$37281 ( \37534 , \37532 , \37533 );
xor \U$37282 ( \37535 , \37524 , \37534 );
not \U$37283 ( \37536 , \37535 );
or \U$37284 ( \37537 , \37508 , \37536 );
or \U$37285 ( \37538 , \37535 , \37507 );
nand \U$37286 ( \37539 , \37537 , \37538 );
not \U$37287 ( \37540 , RIbe29bf0_71);
not \U$37288 ( \37541 , \6380 );
or \U$37289 ( \37542 , \37540 , \37541 );
nand \U$37290 ( \37543 , \1117 , RIbe28f48_44);
nand \U$37291 ( \37544 , \37542 , \37543 );
and \U$37292 ( \37545 , \37544 , \1132 );
not \U$37293 ( \37546 , \37544 );
and \U$37294 ( \37547 , \37546 , \1448 );
nor \U$37295 ( \37548 , \37545 , \37547 );
not \U$37296 ( \37549 , \37548 );
not \U$37297 ( \37550 , \37549 );
not \U$37298 ( \37551 , RIbe29dd0_75);
not \U$37299 ( \37552 , \1094 );
or \U$37300 ( \37553 , \37551 , \37552 );
nand \U$37301 ( \37554 , \1099 , RIbe29c68_72);
nand \U$37302 ( \37555 , \37553 , \37554 );
and \U$37303 ( \37556 , \37555 , \5125 );
not \U$37304 ( \37557 , \37555 );
and \U$37305 ( \37558 , \37557 , \1309 );
nor \U$37306 ( \37559 , \37556 , \37558 );
not \U$37307 ( \37560 , \37559 );
not \U$37308 ( \37561 , \37560 );
or \U$37309 ( \37562 , \37550 , \37561 );
nand \U$37310 ( \37563 , \37548 , \37559 );
nand \U$37311 ( \37564 , \37562 , \37563 );
not \U$37312 ( \37565 , RIbe29fb0_79);
not \U$37313 ( \37566 , \1143 );
or \U$37314 ( \37567 , \37565 , \37566 );
nand \U$37315 ( \37568 , \1147 , RIbe29e48_76);
nand \U$37316 ( \37569 , \37567 , \37568 );
not \U$37317 ( \37570 , \37569 );
not \U$37318 ( \37571 , \1153 );
and \U$37319 ( \37572 , \37570 , \37571 );
and \U$37320 ( \37573 , \37569 , \3994 );
nor \U$37321 ( \37574 , \37572 , \37573 );
xnor \U$37322 ( \37575 , \37564 , \37574 );
not \U$37323 ( \37576 , \37575 );
and \U$37324 ( \37577 , \37539 , \37576 );
not \U$37325 ( \37578 , \37539 );
and \U$37326 ( \37579 , \37578 , \37575 );
nor \U$37327 ( \37580 , \37577 , \37579 );
not \U$37328 ( \37581 , \37580 );
and \U$37329 ( \37582 , \37472 , \37581 );
not \U$37330 ( \37583 , \37472 );
and \U$37331 ( \37584 , \37583 , \37580 );
nor \U$37332 ( \37585 , \37582 , \37584 );
xnor \U$37333 ( \37586 , \37262 , \37585 );
nor \U$37334 ( \37587 , \37217 , \37586 );
and \U$37335 ( \37588 , \37215 , \37191 );
nor \U$37336 ( \37589 , \37587 , \37588 );
not \U$37337 ( \37590 , \36618 );
nand \U$37338 ( \37591 , \37590 , \36629 );
not \U$37339 ( \37592 , \36623 );
and \U$37340 ( \37593 , \37591 , \37592 );
and \U$37341 ( \37594 , \36618 , \36628 );
nor \U$37342 ( \37595 , \37593 , \37594 );
not \U$37343 ( \37596 , \36864 );
not \U$37344 ( \37597 , \36768 );
and \U$37345 ( \37598 , \37596 , \37597 );
and \U$37346 ( \37599 , \36768 , \36864 );
nor \U$37347 ( \37600 , \37598 , \37599 );
buf \U$37348 ( \37601 , \36796 );
nand \U$37349 ( \37602 , \37600 , \37601 );
and \U$37350 ( \37603 , \37602 , \37064 );
nor \U$37351 ( \37604 , \37600 , \37601 );
nor \U$37352 ( \37605 , \37603 , \37604 );
xor \U$37353 ( \37606 , \37595 , \37605 );
xor \U$37354 ( \37607 , \36579 , \36583 );
and \U$37355 ( \37608 , \37607 , \36588 );
and \U$37356 ( \37609 , \36579 , \36583 );
or \U$37357 ( \37610 , \37608 , \37609 );
and \U$37358 ( \37611 , \37606 , \37610 );
and \U$37359 ( \37612 , \37595 , \37605 );
or \U$37360 ( \37613 , \37611 , \37612 );
and \U$37361 ( \37614 , \37589 , \37613 );
not \U$37362 ( \37615 , \37589 );
not \U$37363 ( \37616 , \37613 );
and \U$37364 ( \37617 , \37615 , \37616 );
nor \U$37365 ( \37618 , \37614 , \37617 );
xor \U$37366 ( \37619 , \37138 , \37164 );
and \U$37367 ( \37620 , \37619 , \37189 );
and \U$37368 ( \37621 , \37138 , \37164 );
or \U$37369 ( \37622 , \37620 , \37621 );
nand \U$37370 ( \37623 , \37482 , \37502 );
and \U$37371 ( \37624 , \37623 , \37492 );
nor \U$37372 ( \37625 , \37482 , \37502 );
nor \U$37373 ( \37626 , \37624 , \37625 );
not \U$37374 ( \37627 , \37626 );
not \U$37375 ( \37628 , \37627 );
not \U$37376 ( \37629 , \37517 );
nand \U$37377 ( \37630 , \37629 , \37523 );
not \U$37378 ( \37631 , \37630 );
not \U$37379 ( \37632 , \37534 );
or \U$37380 ( \37633 , \37631 , \37632 );
not \U$37381 ( \37634 , \37523 );
nand \U$37382 ( \37635 , \37634 , \37517 );
nand \U$37383 ( \37636 , \37633 , \37635 );
not \U$37384 ( \37637 , \37636 );
not \U$37385 ( \37638 , \37637 );
or \U$37386 ( \37639 , \37628 , \37638 );
nand \U$37387 ( \37640 , \37636 , \37626 );
nand \U$37388 ( \37641 , \37639 , \37640 );
not \U$37389 ( \37642 , \37641 );
and \U$37390 ( \37643 , \37574 , \37559 );
nor \U$37391 ( \37644 , \37643 , \37549 );
not \U$37392 ( \37645 , \37560 );
nor \U$37393 ( \37646 , \37645 , \37574 );
nor \U$37394 ( \37647 , \37644 , \37646 );
not \U$37395 ( \37648 , \37647 );
and \U$37396 ( \37649 , \37642 , \37648 );
and \U$37397 ( \37650 , \37641 , \37647 );
nor \U$37398 ( \37651 , \37649 , \37650 );
nand \U$37399 ( \37652 , \37308 , \37329 );
and \U$37400 ( \37653 , \37652 , \37320 );
nor \U$37401 ( \37654 , \37308 , \37329 );
nor \U$37402 ( \37655 , \37653 , \37654 );
not \U$37403 ( \37656 , \37655 );
not \U$37404 ( \37657 , \37656 );
or \U$37405 ( \37658 , \37271 , \37282 );
nand \U$37406 ( \37659 , \37658 , \37294 );
nand \U$37407 ( \37660 , \37282 , \37271 );
nand \U$37408 ( \37661 , \37659 , \37660 );
not \U$37409 ( \37662 , \37661 );
not \U$37410 ( \37663 , \37662 );
or \U$37411 ( \37664 , \37657 , \37663 );
nand \U$37412 ( \37665 , \37655 , \37661 );
nand \U$37413 ( \37666 , \37664 , \37665 );
nand \U$37414 ( \37667 , \37350 , \37369 );
and \U$37415 ( \37668 , \37667 , \37359 );
nor \U$37416 ( \37669 , \37350 , \37369 );
nor \U$37417 ( \37670 , \37668 , \37669 );
and \U$37418 ( \37671 , \37666 , \37670 );
not \U$37419 ( \37672 , \37666 );
not \U$37420 ( \37673 , \37670 );
and \U$37421 ( \37674 , \37672 , \37673 );
nor \U$37422 ( \37675 , \37671 , \37674 );
xor \U$37423 ( \37676 , \37651 , \37675 );
not \U$37424 ( \37677 , \13068 );
and \U$37425 ( \37678 , \37389 , \12774 );
not \U$37426 ( \37679 , \37389 );
and \U$37427 ( \37680 , \37679 , \12924 );
nor \U$37428 ( \37681 , \37678 , \37680 );
not \U$37429 ( \37682 , \37681 );
or \U$37430 ( \37683 , \37677 , \37682 );
not \U$37431 ( \37684 , \37382 );
nand \U$37432 ( \37685 , \37683 , \37684 );
not \U$37433 ( \37686 , \37681 );
nand \U$37434 ( \37687 , \37686 , \12723 );
nand \U$37435 ( \37688 , \37685 , \37687 );
not \U$37436 ( \37689 , \37436 );
not \U$37437 ( \37690 , \37460 );
or \U$37438 ( \37691 , \37689 , \37690 );
or \U$37439 ( \37692 , \37460 , \37436 );
not \U$37440 ( \37693 , \37447 );
nand \U$37441 ( \37694 , \37692 , \37693 );
nand \U$37442 ( \37695 , \37691 , \37694 );
xor \U$37443 ( \37696 , \37688 , \37695 );
xor \U$37444 ( \37697 , \37405 , \37414 );
and \U$37445 ( \37698 , \37697 , \37424 );
and \U$37446 ( \37699 , \37405 , \37414 );
or \U$37447 ( \37700 , \37698 , \37699 );
xor \U$37448 ( \37701 , \37696 , \37700 );
xor \U$37449 ( \37702 , \37676 , \37701 );
xor \U$37450 ( \37703 , \37622 , \37702 );
nand \U$37451 ( \37704 , RIbe29380_53, RIbe2b090_115);
not \U$37452 ( \37705 , RIbe2a280_85);
not \U$37453 ( \37706 , \324 );
or \U$37454 ( \37707 , \37705 , \37706 );
nand \U$37455 ( \37708 , \329 , RIbe2a208_84);
nand \U$37456 ( \37709 , \37707 , \37708 );
not \U$37457 ( \37710 , \37709 );
not \U$37458 ( \37711 , \12321 );
and \U$37459 ( \37712 , \37710 , \37711 );
and \U$37460 ( \37713 , \37709 , \1374 );
nor \U$37461 ( \37714 , \37712 , \37713 );
xor \U$37462 ( \37715 , \37704 , \37714 );
not \U$37463 ( \37716 , \300 );
not \U$37464 ( \37717 , RIbe2a550_91);
not \U$37465 ( \37718 , \1679 );
or \U$37466 ( \37719 , \37717 , \37718 );
nand \U$37467 ( \37720 , \1531 , RIbe2a988_100);
nand \U$37468 ( \37721 , \37719 , \37720 );
not \U$37469 ( \37722 , \37721 );
or \U$37470 ( \37723 , \37716 , \37722 );
or \U$37471 ( \37724 , \37721 , \300 );
nand \U$37472 ( \37725 , \37723 , \37724 );
not \U$37473 ( \37726 , RIbe2a190_83);
not \U$37474 ( \37727 , \260 );
or \U$37475 ( \37728 , \37726 , \37727 );
nand \U$37476 ( \37729 , \263 , RIbe2a5c8_92);
nand \U$37477 ( \37730 , \37728 , \37729 );
not \U$37478 ( \37731 , \37730 );
not \U$37479 ( \37732 , \6058 );
and \U$37480 ( \37733 , \37731 , \37732 );
and \U$37481 ( \37734 , \6058 , \37730 );
nor \U$37482 ( \37735 , \37733 , \37734 );
and \U$37483 ( \37736 , \37725 , \37735 );
not \U$37484 ( \37737 , \37725 );
not \U$37485 ( \37738 , \37735 );
and \U$37486 ( \37739 , \37737 , \37738 );
or \U$37487 ( \37740 , \37736 , \37739 );
xnor \U$37488 ( \37741 , \37715 , \37740 );
not \U$37489 ( \37742 , \6583 );
not \U$37490 ( \37743 , RIbe280c0_13);
not \U$37491 ( \37744 , \20487 );
or \U$37492 ( \37745 , \37743 , \37744 );
nand \U$37493 ( \37746 , \7278 , RIbe29830_63);
nand \U$37494 ( \37747 , \37745 , \37746 );
not \U$37495 ( \37748 , \37747 );
and \U$37496 ( \37749 , \37742 , \37748 );
and \U$37497 ( \37750 , \37747 , \9868 );
nor \U$37498 ( \37751 , \37749 , \37750 );
not \U$37499 ( \37752 , RIbe296c8_60);
not \U$37500 ( \37753 , \21608 );
or \U$37501 ( \37754 , \37752 , \37753 );
nand \U$37502 ( \37755 , \7958 , RIbe29650_59);
nand \U$37503 ( \37756 , \37754 , \37755 );
and \U$37504 ( \37757 , \37756 , \7293 );
not \U$37505 ( \37758 , \37756 );
and \U$37506 ( \37759 , \37758 , \6572 );
nor \U$37507 ( \37760 , \37757 , \37759 );
xor \U$37508 ( \37761 , \37751 , \37760 );
not \U$37509 ( \37762 , RIbe28228_16);
not \U$37510 ( \37763 , \6536 );
or \U$37511 ( \37764 , \37762 , \37763 );
nand \U$37512 ( \37765 , \10348 , RIbe281b0_15);
nand \U$37513 ( \37766 , \37764 , \37765 );
and \U$37514 ( \37767 , \37766 , \15730 );
not \U$37515 ( \37768 , \37766 );
and \U$37516 ( \37769 , \37768 , \6891 );
nor \U$37517 ( \37770 , \37767 , \37769 );
xor \U$37518 ( \37771 , \37761 , \37770 );
not \U$37519 ( \37772 , \37771 );
not \U$37520 ( \37773 , RIbe28930_31);
not \U$37521 ( \37774 , \6138 );
or \U$37522 ( \37775 , \37773 , \37774 );
nand \U$37523 ( \37776 , \8235 , RIbe29560_57);
nand \U$37524 ( \37777 , \37775 , \37776 );
and \U$37525 ( \37778 , \37777 , \6623 );
not \U$37526 ( \37779 , \37777 );
and \U$37527 ( \37780 , \37779 , \10972 );
nor \U$37528 ( \37781 , \37778 , \37780 );
not \U$37529 ( \37782 , RIbe28b88_36);
not \U$37530 ( \37783 , \4829 );
or \U$37531 ( \37784 , \37782 , \37783 );
nand \U$37532 ( \37785 , \7056 , RIbe29290_51);
nand \U$37533 ( \37786 , \37784 , \37785 );
and \U$37534 ( \37787 , \37786 , \4586 );
not \U$37535 ( \37788 , \37786 );
and \U$37536 ( \37789 , \37788 , \4946 );
nor \U$37537 ( \37790 , \37787 , \37789 );
xor \U$37538 ( \37791 , \37781 , \37790 );
not \U$37539 ( \37792 , RIbe28a20_33);
not \U$37540 ( \37793 , \15313 );
or \U$37541 ( \37794 , \37792 , \37793 );
nand \U$37542 ( \37795 , \7100 , RIbe289a8_32);
nand \U$37543 ( \37796 , \37794 , \37795 );
and \U$37544 ( \37797 , \37796 , \6121 );
not \U$37545 ( \37798 , \37796 );
and \U$37546 ( \37799 , \37798 , \8252 );
nor \U$37547 ( \37800 , \37797 , \37799 );
xor \U$37548 ( \37801 , \37791 , \37800 );
not \U$37549 ( \37802 , \37801 );
or \U$37550 ( \37803 , \37772 , \37802 );
or \U$37551 ( \37804 , \37801 , \37771 );
nand \U$37552 ( \37805 , \37803 , \37804 );
not \U$37553 ( \37806 , RIbe28480_21);
not \U$37554 ( \37807 , \5094 );
or \U$37555 ( \37808 , \37806 , \37807 );
nand \U$37556 ( \37809 , \7438 , RIbe28408_20);
nand \U$37557 ( \37810 , \37808 , \37809 );
and \U$37558 ( \37811 , \37810 , \3471 );
not \U$37559 ( \37812 , \37810 );
and \U$37560 ( \37813 , \37812 , \3448 );
nor \U$37561 ( \37814 , \37811 , \37813 );
not \U$37562 ( \37815 , \37814 );
not \U$37563 ( \37816 , \37815 );
not \U$37564 ( \37817 , RIbe28390_19);
not \U$37565 ( \37818 , \5058 );
or \U$37566 ( \37819 , \37817 , \37818 );
nand \U$37567 ( \37820 , \4600 , RIbe28b10_35);
nand \U$37568 ( \37821 , \37819 , \37820 );
and \U$37569 ( \37822 , \37821 , \7865 );
not \U$37570 ( \37823 , \37821 );
and \U$37571 ( \37824 , \37823 , \4603 );
nor \U$37572 ( \37825 , \37822 , \37824 );
not \U$37573 ( \37826 , \37825 );
not \U$37574 ( \37827 , \37826 );
or \U$37575 ( \37828 , \37816 , \37827 );
nand \U$37576 ( \37829 , \37825 , \37814 );
nand \U$37577 ( \37830 , \37828 , \37829 );
not \U$37578 ( \37831 , RIbe285e8_24);
not \U$37579 ( \37832 , \3285 );
or \U$37580 ( \37833 , \37831 , \37832 );
nand \U$37581 ( \37834 , \3689 , RIbe287c8_28);
nand \U$37582 ( \37835 , \37833 , \37834 );
and \U$37583 ( \37836 , \37835 , \3461 );
not \U$37584 ( \37837 , \37835 );
and \U$37585 ( \37838 , \37837 , \3290 );
nor \U$37586 ( \37839 , \37836 , \37838 );
and \U$37587 ( \37840 , \37830 , \37839 );
not \U$37588 ( \37841 , \37830 );
not \U$37589 ( \37842 , \37839 );
and \U$37590 ( \37843 , \37841 , \37842 );
nor \U$37591 ( \37844 , \37840 , \37843 );
and \U$37592 ( \37845 , \37805 , \37844 );
not \U$37593 ( \37846 , \37805 );
not \U$37594 ( \37847 , \37844 );
and \U$37595 ( \37848 , \37846 , \37847 );
nor \U$37596 ( \37849 , \37845 , \37848 );
xor \U$37597 ( \37850 , \37741 , \37849 );
not \U$37598 ( \37851 , RIbe2a028_80);
not \U$37599 ( \37852 , \23339 );
or \U$37600 ( \37853 , \37851 , \37852 );
nand \U$37601 ( \37854 , \1202 , RIbe29fb0_79);
nand \U$37602 ( \37855 , \37853 , \37854 );
and \U$37603 ( \37856 , \37855 , \1011 );
not \U$37604 ( \37857 , \37855 );
and \U$37605 ( \37858 , \37857 , \1608 );
nor \U$37606 ( \37859 , \37856 , \37858 );
not \U$37607 ( \37860 , RIbe29e48_76);
not \U$37608 ( \37861 , \4257 );
or \U$37609 ( \37862 , \37860 , \37861 );
nand \U$37610 ( \37863 , RIbe29dd0_75, \1146 );
nand \U$37611 ( \37864 , \37862 , \37863 );
and \U$37612 ( \37865 , \37864 , \1154 );
not \U$37613 ( \37866 , \37864 );
and \U$37614 ( \37867 , \37866 , \1153 );
nor \U$37615 ( \37868 , \37865 , \37867 );
xor \U$37616 ( \37869 , \37859 , \37868 );
not \U$37617 ( \37870 , RIbe29c68_72);
not \U$37618 ( \37871 , \1094 );
or \U$37619 ( \37872 , \37870 , \37871 );
nand \U$37620 ( \37873 , RIbe29bf0_71, \1099 );
nand \U$37621 ( \37874 , \37872 , \37873 );
and \U$37622 ( \37875 , \37874 , \1309 );
not \U$37623 ( \37876 , \37874 );
and \U$37624 ( \37877 , \37876 , \4251 );
nor \U$37625 ( \37878 , \37875 , \37877 );
xor \U$37626 ( \37879 , \37869 , \37878 );
not \U$37627 ( \37880 , \37879 );
not \U$37628 ( \37881 , \37880 );
not \U$37629 ( \37882 , \2889 );
not \U$37630 ( \37883 , \7180 );
and \U$37631 ( \37884 , \37882 , \37883 );
and \U$37632 ( \37885 , \2390 , RIbe27fd0_11);
nor \U$37633 ( \37886 , \37884 , \37885 );
and \U$37634 ( \37887 , \37886 , \7038 );
not \U$37635 ( \37888 , \37886 );
and \U$37636 ( \37889 , \37888 , \9083 );
nor \U$37637 ( \37890 , \37887 , \37889 );
not \U$37638 ( \37891 , RIbe27e68_8);
not \U$37639 ( \37892 , \3476 );
or \U$37640 ( \37893 , \37891 , \37892 );
not \U$37641 ( \37894 , \25899 );
nand \U$37642 ( \37895 , \37894 , \2900 );
nand \U$37643 ( \37896 , \37893 , \37895 );
and \U$37644 ( \37897 , \37896 , \4059 );
not \U$37645 ( \37898 , \37896 );
and \U$37646 ( \37899 , \37898 , \2380 );
nor \U$37647 ( \37900 , \37897 , \37899 );
and \U$37648 ( \37901 , \37890 , \37900 );
not \U$37649 ( \37902 , \37890 );
not \U$37650 ( \37903 , \37900 );
and \U$37651 ( \37904 , \37902 , \37903 );
or \U$37652 ( \37905 , \37901 , \37904 );
not \U$37653 ( \37906 , RIbe28f48_44);
not \U$37654 ( \37907 , \1112 );
or \U$37655 ( \37908 , \37906 , \37907 );
nand \U$37656 ( \37909 , RIbe28ed0_43, \5467 );
nand \U$37657 ( \37910 , \37908 , \37909 );
not \U$37658 ( \37911 , \37910 );
not \U$37659 ( \37912 , \1125 );
and \U$37660 ( \37913 , \37911 , \37912 );
and \U$37661 ( \37914 , \37910 , \3491 );
nor \U$37662 ( \37915 , \37913 , \37914 );
and \U$37663 ( \37916 , \37905 , \37915 );
not \U$37664 ( \37917 , \37905 );
not \U$37665 ( \37918 , \37915 );
and \U$37666 ( \37919 , \37917 , \37918 );
nor \U$37667 ( \37920 , \37916 , \37919 );
not \U$37668 ( \37921 , \37920 );
not \U$37669 ( \37922 , \37921 );
or \U$37670 ( \37923 , \37881 , \37922 );
nand \U$37671 ( \37924 , \37920 , \37879 );
nand \U$37672 ( \37925 , \37923 , \37924 );
not \U$37673 ( \37926 , RIbe2a2f8_86);
not \U$37674 ( \37927 , \6350 );
or \U$37675 ( \37928 , \37926 , \37927 );
nand \U$37676 ( \37929 , \740 , RIbe2acd0_107);
nand \U$37677 ( \37930 , \37928 , \37929 );
not \U$37678 ( \37931 , \37930 );
not \U$37679 ( \37932 , \564 );
and \U$37680 ( \37933 , \37931 , \37932 );
and \U$37681 ( \37934 , \37930 , \564 );
nor \U$37682 ( \37935 , \37933 , \37934 );
not \U$37683 ( \37936 , \37935 );
not \U$37684 ( \37937 , \37936 );
not \U$37685 ( \37938 , RIbe2a3e8_88);
not \U$37686 ( \37939 , \546 );
or \U$37687 ( \37940 , \37938 , \37939 );
nand \U$37688 ( \37941 , \552 , RIbe2a370_87);
nand \U$37689 ( \37942 , \37940 , \37941 );
and \U$37690 ( \37943 , \37942 , \1761 );
not \U$37691 ( \37944 , \37942 );
and \U$37692 ( \37945 , \37944 , \6340 );
nor \U$37693 ( \37946 , \37943 , \37945 );
not \U$37694 ( \37947 , \37946 );
not \U$37695 ( \37948 , \37947 );
or \U$37696 ( \37949 , \37937 , \37948 );
nand \U$37697 ( \37950 , \37946 , \37935 );
nand \U$37698 ( \37951 , \37949 , \37950 );
not \U$37699 ( \37952 , RIbe2a910_99);
not \U$37700 ( \37953 , \1337 );
or \U$37701 ( \37954 , \37952 , \37953 );
nand \U$37702 ( \37955 , \429 , RIbe2b5b8_126);
nand \U$37703 ( \37956 , \37954 , \37955 );
not \U$37704 ( \37957 , \37956 );
not \U$37705 ( \37958 , \1232 );
and \U$37706 ( \37959 , \37957 , \37958 );
and \U$37707 ( \37960 , \37956 , \3175 );
nor \U$37708 ( \37961 , \37959 , \37960 );
and \U$37709 ( \37962 , \37951 , \37961 );
not \U$37710 ( \37963 , \37951 );
not \U$37711 ( \37964 , \37961 );
and \U$37712 ( \37965 , \37963 , \37964 );
nor \U$37713 ( \37966 , \37962 , \37965 );
and \U$37714 ( \37967 , \37925 , \37966 );
not \U$37715 ( \37968 , \37925 );
not \U$37716 ( \37969 , \37966 );
and \U$37717 ( \37970 , \37968 , \37969 );
nor \U$37718 ( \37971 , \37967 , \37970 );
xor \U$37719 ( \37972 , \37850 , \37971 );
xor \U$37720 ( \37973 , \37703 , \37972 );
not \U$37721 ( \37974 , \37973 );
not \U$37722 ( \37975 , \37974 );
not \U$37723 ( \37976 , \37221 );
nand \U$37724 ( \37977 , \37976 , \37227 );
not \U$37725 ( \37978 , \37221 );
not \U$37726 ( \37979 , \37227 );
not \U$37727 ( \37980 , \37979 );
or \U$37728 ( \37981 , \37978 , \37980 );
nand \U$37729 ( \37982 , \37981 , \37233 );
nand \U$37730 ( \37983 , \37977 , \37982 );
not \U$37731 ( \37984 , \37242 );
not \U$37732 ( \37985 , \37252 );
or \U$37733 ( \37986 , \37984 , \37985 );
nand \U$37734 ( \37987 , \37986 , \37247 );
not \U$37735 ( \37988 , \37242 );
nand \U$37736 ( \37989 , \37988 , \37253 );
nand \U$37737 ( \37990 , \37987 , \37989 );
xor \U$37738 ( \37991 , \37983 , \37990 );
nand \U$37739 ( \37992 , \37466 , \37580 );
and \U$37740 ( \37993 , \37992 , \37371 );
nor \U$37741 ( \37994 , \37580 , \37466 );
nor \U$37742 ( \37995 , \37993 , \37994 );
and \U$37743 ( \37996 , \37991 , \37995 );
not \U$37744 ( \37997 , \37991 );
not \U$37745 ( \37998 , \37995 );
and \U$37746 ( \37999 , \37997 , \37998 );
nor \U$37747 ( \38000 , \37996 , \37999 );
not \U$37748 ( \38001 , \37187 );
not \U$37749 ( \38002 , \37172 );
or \U$37750 ( \38003 , \38001 , \38002 );
not \U$37751 ( \38004 , \37184 );
not \U$37752 ( \38005 , \37171 );
or \U$37753 ( \38006 , \38004 , \38005 );
nand \U$37754 ( \38007 , \38006 , \37179 );
nand \U$37755 ( \38008 , \38003 , \38007 );
not \U$37756 ( \38009 , \37121 );
not \U$37757 ( \38010 , \37109 );
or \U$37758 ( \38011 , \38009 , \38010 );
or \U$37759 ( \38012 , \37109 , \37121 );
nand \U$37760 ( \38013 , \38012 , \37113 );
nand \U$37761 ( \38014 , \38011 , \38013 );
and \U$37762 ( \38015 , \38008 , \38014 );
not \U$37763 ( \38016 , \38008 );
not \U$37764 ( \38017 , \38014 );
and \U$37765 ( \38018 , \38016 , \38017 );
nor \U$37766 ( \38019 , \38015 , \38018 );
not \U$37767 ( \38020 , \37155 );
not \U$37768 ( \38021 , \37150 );
or \U$37769 ( \38022 , \38020 , \38021 );
nand \U$37770 ( \38023 , \38022 , \37144 );
not \U$37771 ( \38024 , \37150 );
nand \U$37772 ( \38025 , \38024 , \37158 );
nand \U$37773 ( \38026 , \38023 , \38025 );
not \U$37774 ( \38027 , \38026 );
and \U$37775 ( \38028 , \38019 , \38027 );
not \U$37776 ( \38029 , \38019 );
and \U$37777 ( \38030 , \38029 , \38026 );
nor \U$37778 ( \38031 , \38028 , \38030 );
not \U$37779 ( \38032 , \38031 );
nand \U$37780 ( \38033 , \13738 , RIbe27b98_2);
xnor \U$37781 ( \38034 , \38033 , \12924 );
not \U$37782 ( \38035 , \12960 );
not \U$37783 ( \38036 , RIbe28de0_41);
not \U$37784 ( \38037 , \15205 );
or \U$37785 ( \38038 , \38036 , \38037 );
nand \U$37786 ( \38039 , \13669 , RIbe29920_65);
nand \U$37787 ( \38040 , \38038 , \38039 );
not \U$37788 ( \38041 , \38040 );
or \U$37789 ( \38042 , \38035 , \38041 );
or \U$37790 ( \38043 , \38040 , \12960 );
nand \U$37791 ( \38044 , \38042 , \38043 );
xor \U$37792 ( \38045 , \38034 , \38044 );
not \U$37793 ( \38046 , RIbe27c10_3);
not \U$37794 ( \38047 , \13024 );
or \U$37795 ( \38048 , \38046 , \38047 );
nand \U$37796 ( \38049 , \14511 , RIbe28e58_42);
nand \U$37797 ( \38050 , \38048 , \38049 );
and \U$37798 ( \38051 , \38050 , \14756 );
not \U$37799 ( \38052 , \38050 );
and \U$37800 ( \38053 , \38052 , \9904 );
nor \U$37801 ( \38054 , \38051 , \38053 );
xnor \U$37802 ( \38055 , \38045 , \38054 );
not \U$37803 ( \38056 , \38055 );
not \U$37804 ( \38057 , RIbe29038_46);
not \U$37805 ( \38058 , \7298 );
or \U$37806 ( \38059 , \38057 , \38058 );
nand \U$37807 ( \38060 , \13224 , RIbe28fc0_45);
nand \U$37808 ( \38061 , \38059 , \38060 );
and \U$37809 ( \38062 , \38061 , \7660 );
not \U$37810 ( \38063 , \38061 );
and \U$37811 ( \38064 , \38063 , \13168 );
nor \U$37812 ( \38065 , \38062 , \38064 );
not \U$37813 ( \38066 , RIbe290b0_47);
not \U$37814 ( \38067 , \10949 );
or \U$37815 ( \38068 , \38066 , \38067 );
nand \U$37816 ( \38069 , \7981 , RIbe29a88_68);
nand \U$37817 ( \38070 , \38068 , \38069 );
and \U$37818 ( \38071 , \38070 , \14299 );
not \U$37819 ( \38072 , \38070 );
and \U$37820 ( \38073 , \38072 , \7984 );
nor \U$37821 ( \38074 , \38071 , \38073 );
xor \U$37822 ( \38075 , \38065 , \38074 );
and \U$37823 ( \38076 , \10916 , RIbe27d78_6);
and \U$37824 ( \38077 , \14771 , RIbe27d00_5);
nor \U$37825 ( \38078 , \38076 , \38077 );
and \U$37826 ( \38079 , \38078 , \15233 );
not \U$37827 ( \38080 , \38078 );
and \U$37828 ( \38081 , \38080 , \18797 );
nor \U$37829 ( \38082 , \38079 , \38081 );
xor \U$37830 ( \38083 , \38075 , \38082 );
not \U$37831 ( \38084 , \38083 );
or \U$37832 ( \38085 , \38056 , \38084 );
or \U$37833 ( \38086 , \38055 , \38083 );
nand \U$37834 ( \38087 , \38085 , \38086 );
not \U$37835 ( \38088 , \38087 );
not \U$37836 ( \38089 , \38088 );
not \U$37837 ( \38090 , \37461 );
not \U$37838 ( \38091 , \37394 );
or \U$37839 ( \38092 , \38090 , \38091 );
nand \U$37840 ( \38093 , \38092 , \37425 );
not \U$37841 ( \38094 , \37394 );
nand \U$37842 ( \38095 , \38094 , \37464 );
nand \U$37843 ( \38096 , \38093 , \38095 );
not \U$37844 ( \38097 , \38096 );
or \U$37845 ( \38098 , \38089 , \38097 );
nand \U$37846 ( \38099 , \38087 , \38093 , \38095 );
nand \U$37847 ( \38100 , \38098 , \38099 );
not \U$37848 ( \38101 , \38100 );
or \U$37849 ( \38102 , \38032 , \38101 );
or \U$37850 ( \38103 , \38031 , \38100 );
nand \U$37851 ( \38104 , \38102 , \38103 );
xor \U$37852 ( \38105 , \37129 , \37136 );
and \U$37853 ( \38106 , \38105 , \36879 );
and \U$37854 ( \38107 , \37129 , \37136 );
or \U$37855 ( \38108 , \38106 , \38107 );
or \U$37856 ( \38109 , \37575 , \37507 );
not \U$37857 ( \38110 , \37535 );
nand \U$37858 ( \38111 , \38109 , \38110 );
nand \U$37859 ( \38112 , \37575 , \37507 );
nand \U$37860 ( \38113 , \38111 , \38112 );
xor \U$37861 ( \38114 , \38108 , \38113 );
xor \U$37862 ( \38115 , \37299 , \37339 );
and \U$37863 ( \38116 , \38115 , \37370 );
and \U$37864 ( \38117 , \37299 , \37339 );
or \U$37865 ( \38118 , \38116 , \38117 );
xor \U$37866 ( \38119 , \38114 , \38118 );
not \U$37867 ( \38120 , \38119 );
and \U$37868 ( \38121 , \38104 , \38120 );
not \U$37869 ( \38122 , \38104 );
and \U$37870 ( \38123 , \38122 , \38119 );
nor \U$37871 ( \38124 , \38121 , \38123 );
xor \U$37872 ( \38125 , \38000 , \38124 );
not \U$37873 ( \38126 , \38125 );
or \U$37874 ( \38127 , \37975 , \38126 );
or \U$37875 ( \38128 , \37974 , \38125 );
nand \U$37876 ( \38129 , \38127 , \38128 );
and \U$37877 ( \38130 , \37618 , \38129 );
not \U$37878 ( \38131 , \37618 );
not \U$37879 ( \38132 , \38129 );
and \U$37880 ( \38133 , \38131 , \38132 );
nor \U$37881 ( \38134 , \38130 , \38133 );
xor \U$37882 ( \38135 , \37215 , \37191 );
not \U$37883 ( \38136 , \37586 );
and \U$37884 ( \38137 , \38135 , \38136 );
not \U$37885 ( \38138 , \38135 );
and \U$37886 ( \38139 , \38138 , \37586 );
nor \U$37887 ( \38140 , \38137 , \38139 );
not \U$37888 ( \38141 , \38140 );
xor \U$37889 ( \38142 , \37077 , \37081 );
and \U$37890 ( \38143 , \38142 , \37087 );
and \U$37891 ( \38144 , \37077 , \37081 );
or \U$37892 ( \38145 , \38143 , \38144 );
xor \U$37893 ( \38146 , \36645 , \36665 );
and \U$37894 ( \38147 , \38146 , \37069 );
and \U$37895 ( \38148 , \36645 , \36665 );
or \U$37896 ( \38149 , \38147 , \38148 );
nand \U$37897 ( \38150 , \38145 , \38149 );
not \U$37898 ( \38151 , \38150 );
or \U$37899 ( \38152 , \38141 , \38151 );
not \U$37900 ( \38153 , \38149 );
not \U$37901 ( \38154 , \38145 );
nand \U$37902 ( \38155 , \38153 , \38154 );
nand \U$37903 ( \38156 , \38152 , \38155 );
not \U$37904 ( \38157 , \37213 );
not \U$37905 ( \38158 , \37196 );
or \U$37906 ( \38159 , \38157 , \38158 );
nand \U$37907 ( \38160 , \38159 , \37204 );
or \U$37908 ( \38161 , \37196 , \37213 );
nand \U$37909 ( \38162 , \38160 , \38161 );
not \U$37910 ( \38163 , \37122 );
not \U$37911 ( \38164 , \37127 );
or \U$37912 ( \38165 , \38163 , \38164 );
not \U$37913 ( \38166 , \37122 );
not \U$37914 ( \38167 , \38166 );
not \U$37915 ( \38168 , \37126 );
or \U$37916 ( \38169 , \38167 , \38168 );
nand \U$37917 ( \38170 , \38169 , \37190 );
nand \U$37918 ( \38171 , \38165 , \38170 );
xor \U$37919 ( \38172 , \38162 , \38171 );
or \U$37920 ( \38173 , \37261 , \37238 );
and \U$37921 ( \38174 , \37585 , \38173 );
and \U$37922 ( \38175 , \37238 , \37261 );
nor \U$37923 ( \38176 , \38174 , \38175 );
xnor \U$37924 ( \38177 , \38172 , \38176 );
and \U$37925 ( \38178 , \38156 , \38177 );
not \U$37926 ( \38179 , \38156 );
not \U$37927 ( \38180 , \38177 );
and \U$37928 ( \38181 , \38179 , \38180 );
nor \U$37929 ( \38182 , \38178 , \38181 );
xor \U$37930 ( \38183 , \38134 , \38182 );
not \U$37931 ( \38184 , \38183 );
xor \U$37932 ( \38185 , \37595 , \37605 );
xor \U$37933 ( \38186 , \38185 , \37610 );
xor \U$37934 ( \38187 , \36630 , \37070 );
and \U$37935 ( \38188 , \38187 , \37088 );
and \U$37936 ( \38189 , \36630 , \37070 );
or \U$37937 ( \38190 , \38188 , \38189 );
xor \U$37938 ( \38191 , \38186 , \38190 );
xor \U$37939 ( \38192 , \36589 , \36593 );
and \U$37940 ( \38193 , \38192 , \36598 );
and \U$37941 ( \38194 , \36589 , \36593 );
or \U$37942 ( \38195 , \38193 , \38194 );
and \U$37943 ( \38196 , \38191 , \38195 );
and \U$37944 ( \38197 , \38186 , \38190 );
or \U$37945 ( \38198 , \38196 , \38197 );
not \U$37946 ( \38199 , \38198 );
and \U$37947 ( \38200 , \38184 , \38199 );
and \U$37948 ( \38201 , \38183 , \38198 );
nor \U$37949 ( \38202 , \38200 , \38201 );
not \U$37950 ( \38203 , \38202 );
not \U$37951 ( \38204 , \38203 );
xor \U$37952 ( \38205 , \38149 , \38154 );
xor \U$37953 ( \38206 , \38205 , \38140 );
xor \U$37954 ( \38207 , \38186 , \38190 );
xor \U$37955 ( \38208 , \38207 , \38195 );
xor \U$37956 ( \38209 , \38206 , \38208 );
nand \U$37957 ( \38210 , \36599 , \37089 );
and \U$37958 ( \38211 , \38210 , \36605 );
nor \U$37959 ( \38212 , \36599 , \37089 );
nor \U$37960 ( \38213 , \38211 , \38212 );
and \U$37961 ( \38214 , \38209 , \38213 );
and \U$37962 ( \38215 , \38206 , \38208 );
or \U$37963 ( \38216 , \38214 , \38215 );
buf \U$37964 ( \38217 , \38216 );
not \U$37965 ( \38218 , \38217 );
or \U$37966 ( \38219 , \38204 , \38218 );
not \U$37967 ( \38220 , \38216 );
nand \U$37968 ( \38221 , \38220 , \38202 );
nand \U$37969 ( \38222 , \38219 , \38221 );
xor \U$37970 ( \38223 , \34773 , \35369 );
xor \U$37971 ( \38224 , \38223 , \35376 );
xor \U$37972 ( \38225 , \33664 , \34293 );
or \U$37973 ( \38226 , \38224 , \38225 );
not \U$37974 ( \38227 , \35364 );
not \U$37975 ( \38228 , \35333 );
not \U$37976 ( \38229 , \35340 );
and \U$37977 ( \38230 , \38228 , \38229 );
and \U$37978 ( \38231 , \35333 , \35340 );
nor \U$37979 ( \38232 , \38230 , \38231 );
not \U$37980 ( \38233 , \38232 );
or \U$37981 ( \38234 , \38227 , \38233 );
or \U$37982 ( \38235 , \35364 , \38232 );
nand \U$37983 ( \38236 , \38234 , \38235 );
not \U$37984 ( \38237 , \35321 );
not \U$37985 ( \38238 , \35325 );
or \U$37986 ( \38239 , \38237 , \38238 );
nand \U$37987 ( \38240 , \35310 , \35320 );
nand \U$37988 ( \38241 , \38239 , \38240 );
and \U$37989 ( \38242 , \38241 , \35329 );
not \U$37990 ( \38243 , \38241 );
not \U$37991 ( \38244 , \35329 );
and \U$37992 ( \38245 , \38243 , \38244 );
nor \U$37993 ( \38246 , \38242 , \38245 );
xor \U$37994 ( \38247 , \34026 , \34023 );
xnor \U$37995 ( \38248 , \38247 , \33805 );
not \U$37996 ( \38249 , \38248 );
xor \U$37997 ( \38250 , \34155 , \34196 );
xnor \U$37998 ( \38251 , \38250 , \34176 );
nand \U$37999 ( \38252 , \38249 , \38251 );
and \U$38000 ( \38253 , \38246 , \38252 );
not \U$38001 ( \38254 , \38251 );
and \U$38002 ( \38255 , \38254 , \38248 );
nor \U$38003 ( \38256 , \38253 , \38255 );
not \U$38004 ( \38257 , \38256 );
not \U$38005 ( \38258 , \38257 );
xor \U$38006 ( \38259 , \34028 , \34077 );
xor \U$38007 ( \38260 , \38259 , \34198 );
not \U$38008 ( \38261 , \38260 );
or \U$38009 ( \38262 , \38258 , \38261 );
not \U$38010 ( \38263 , \38260 );
not \U$38011 ( \38264 , \38263 );
not \U$38012 ( \38265 , \38256 );
or \U$38013 ( \38266 , \38264 , \38265 );
not \U$38014 ( \38267 , \30908 );
nand \U$38015 ( \38268 , \5151 , \30894 );
not \U$38016 ( \38269 , \38268 );
or \U$38017 ( \38270 , \38267 , \38269 );
nand \U$38018 ( \38271 , \30895 , \338 );
nand \U$38019 ( \38272 , \38270 , \38271 );
not \U$38020 ( \38273 , \38272 );
or \U$38021 ( \38274 , \30952 , \30961 );
nand \U$38022 ( \38275 , \38274 , \30971 );
nand \U$38023 ( \38276 , \30952 , \30961 );
nand \U$38024 ( \38277 , \38275 , \38276 );
not \U$38025 ( \38278 , \38277 );
or \U$38026 ( \38279 , \38273 , \38278 );
or \U$38027 ( \38280 , \38277 , \38272 );
xor \U$38028 ( \38281 , \30919 , \30929 );
and \U$38029 ( \38282 , \38281 , \30940 );
and \U$38030 ( \38283 , \30919 , \30929 );
or \U$38031 ( \38284 , \38282 , \38283 );
nand \U$38032 ( \38285 , \38280 , \38284 );
nand \U$38033 ( \38286 , \38279 , \38285 );
not \U$38034 ( \38287 , \38286 );
not \U$38035 ( \38288 , \31031 );
not \U$38036 ( \38289 , \31019 );
or \U$38037 ( \38290 , \38288 , \38289 );
nand \U$38038 ( \38291 , \38290 , \31042 );
not \U$38039 ( \38292 , \31019 );
nand \U$38040 ( \38293 , \38292 , \31028 );
nand \U$38041 ( \38294 , \38291 , \38293 );
not \U$38042 ( \38295 , \38294 );
not \U$38043 ( \38296 , \30984 );
not \U$38044 ( \38297 , \30992 );
or \U$38045 ( \38298 , \38296 , \38297 );
not \U$38046 ( \38299 , \30983 );
not \U$38047 ( \38300 , \30993 );
or \U$38048 ( \38301 , \38299 , \38300 );
nand \U$38049 ( \38302 , \38301 , \31007 );
nand \U$38050 ( \38303 , \38298 , \38302 );
not \U$38051 ( \38304 , \38303 );
or \U$38052 ( \38305 , \38295 , \38304 );
not \U$38053 ( \38306 , \38294 );
not \U$38054 ( \38307 , \38306 );
not \U$38055 ( \38308 , \38303 );
not \U$38056 ( \38309 , \38308 );
or \U$38057 ( \38310 , \38307 , \38309 );
not \U$38058 ( \38311 , \31058 );
and \U$38059 ( \38312 , \31083 , \38311 );
nor \U$38060 ( \38313 , \38312 , \31069 );
nor \U$38061 ( \38314 , \31083 , \38311 );
nor \U$38062 ( \38315 , \38313 , \38314 );
not \U$38063 ( \38316 , \38315 );
nand \U$38064 ( \38317 , \38310 , \38316 );
nand \U$38065 ( \38318 , \38305 , \38317 );
not \U$38066 ( \38319 , \38318 );
or \U$38067 ( \38320 , \38287 , \38319 );
or \U$38068 ( \38321 , \38286 , \38318 );
and \U$38069 ( \38322 , \30811 , \30798 );
not \U$38070 ( \38323 , \30788 );
nor \U$38071 ( \38324 , \38322 , \38323 );
nor \U$38072 ( \38325 , \30811 , \30798 );
nor \U$38073 ( \38326 , \38324 , \38325 );
not \U$38074 ( \38327 , \38326 );
xor \U$38075 ( \38328 , \30822 , \30829 );
and \U$38076 ( \38329 , \38328 , \30839 );
and \U$38077 ( \38330 , \30822 , \30829 );
or \U$38078 ( \38331 , \38329 , \38330 );
not \U$38079 ( \38332 , \38331 );
or \U$38080 ( \38333 , \38327 , \38332 );
nand \U$38081 ( \38334 , \30850 , \30871 );
and \U$38082 ( \38335 , \38334 , \30859 );
nor \U$38083 ( \38336 , \30850 , \30871 );
nor \U$38084 ( \38337 , \38335 , \38336 );
not \U$38085 ( \38338 , \38337 );
nand \U$38086 ( \38339 , \38333 , \38338 );
or \U$38087 ( \38340 , \38331 , \38326 );
nand \U$38088 ( \38341 , \38339 , \38340 );
nand \U$38089 ( \38342 , \38321 , \38341 );
nand \U$38090 ( \38343 , \38320 , \38342 );
not \U$38091 ( \38344 , \38343 );
not \U$38092 ( \38345 , \34961 );
not \U$38093 ( \38346 , \34939 );
or \U$38094 ( \38347 , \38345 , \38346 );
or \U$38095 ( \38348 , \34961 , \34939 );
nand \U$38096 ( \38349 , \38347 , \38348 );
and \U$38097 ( \38350 , \38349 , \34947 );
not \U$38098 ( \38351 , \38349 );
and \U$38099 ( \38352 , \38351 , \34946 );
nor \U$38100 ( \38353 , \38350 , \38352 );
not \U$38101 ( \38354 , \38353 );
xor \U$38102 ( \38355 , \35080 , \35090 );
xor \U$38103 ( \38356 , \38355 , \35101 );
nand \U$38104 ( \38357 , \38354 , \38356 );
not \U$38105 ( \38358 , \38357 );
not \U$38106 ( \38359 , \34972 );
not \U$38107 ( \38360 , \34999 );
or \U$38108 ( \38361 , \38359 , \38360 );
not \U$38109 ( \38362 , \34999 );
nand \U$38110 ( \38363 , \38362 , \34973 );
nand \U$38111 ( \38364 , \38361 , \38363 );
and \U$38112 ( \38365 , \38364 , \34983 );
not \U$38113 ( \38366 , \38364 );
and \U$38114 ( \38367 , \38366 , \34984 );
or \U$38115 ( \38368 , \38365 , \38367 );
not \U$38116 ( \38369 , \38368 );
or \U$38117 ( \38370 , \38358 , \38369 );
not \U$38118 ( \38371 , \38356 );
nand \U$38119 ( \38372 , \38371 , \38353 );
nand \U$38120 ( \38373 , \38370 , \38372 );
not \U$38121 ( \38374 , \38373 );
xor \U$38122 ( \38375 , \33936 , \33934 );
not \U$38123 ( \38376 , \38375 );
xor \U$38124 ( \38377 , \35048 , \35058 );
xor \U$38125 ( \38378 , \38377 , \35069 );
not \U$38126 ( \38379 , \38378 );
xor \U$38127 ( \38380 , \35115 , \35124 );
xor \U$38128 ( \38381 , \38380 , \35134 );
nand \U$38129 ( \38382 , \38379 , \38381 );
nand \U$38130 ( \38383 , \38376 , \38382 );
not \U$38131 ( \38384 , \38383 );
or \U$38132 ( \38385 , \38374 , \38384 );
not \U$38133 ( \38386 , \38382 );
nand \U$38134 ( \38387 , \38386 , \38375 );
nand \U$38135 ( \38388 , \38385 , \38387 );
not \U$38136 ( \38389 , \38388 );
or \U$38137 ( \38390 , \38344 , \38389 );
or \U$38138 ( \38391 , \38388 , \38343 );
not \U$38139 ( \38392 , \30704 );
and \U$38140 ( \38393 , \38392 , \30720 );
nor \U$38141 ( \38394 , \38393 , \30696 );
nor \U$38142 ( \38395 , \38392 , \30720 );
nor \U$38143 ( \38396 , \38394 , \38395 );
not \U$38144 ( \38397 , \38396 );
not \U$38145 ( \38398 , \38397 );
and \U$38146 ( \38399 , \1357 , RIbe2b630_127);
and \U$38147 ( \38400 , \1831 , RIbe2b018_114);
nor \U$38148 ( \38401 , \38399 , \38400 );
and \U$38149 ( \38402 , \38401 , \269 );
not \U$38150 ( \38403 , \38401 );
and \U$38151 ( \38404 , \38403 , \1362 );
or \U$38152 ( \38405 , \38402 , \38404 );
not \U$38153 ( \38406 , \38405 );
or \U$38154 ( \38407 , \38398 , \38406 );
not \U$38155 ( \38408 , \38405 );
not \U$38156 ( \38409 , \38408 );
not \U$38157 ( \38410 , \38396 );
or \U$38158 ( \38411 , \38409 , \38410 );
and \U$38159 ( \38412 , \30734 , \30749 );
not \U$38160 ( \38413 , \30743 );
nor \U$38161 ( \38414 , \38412 , \38413 );
nor \U$38162 ( \38415 , \30734 , \30749 );
or \U$38163 ( \38416 , \38414 , \38415 );
nand \U$38164 ( \38417 , \38411 , \38416 );
nand \U$38165 ( \38418 , \38407 , \38417 );
and \U$38166 ( \38419 , \326 , RIbe2ab68_104);
and \U$38167 ( \38420 , \330 , RIbe2aaf0_103);
nor \U$38168 ( \38421 , \38419 , \38420 );
and \U$38169 ( \38422 , \38421 , \339 );
not \U$38170 ( \38423 , \38421 );
and \U$38171 ( \38424 , \38423 , \1378 );
nor \U$38172 ( \38425 , \38422 , \38424 );
xor \U$38173 ( \38426 , \35177 , \35165 );
xnor \U$38174 ( \38427 , \38426 , \35157 );
xor \U$38175 ( \38428 , \38425 , \38427 );
xor \U$38176 ( \38429 , \34846 , \34857 );
xnor \U$38177 ( \38430 , \38429 , \34836 );
and \U$38178 ( \38431 , \38428 , \38430 );
and \U$38179 ( \38432 , \38425 , \38427 );
or \U$38180 ( \38433 , \38431 , \38432 );
xor \U$38181 ( \38434 , \38418 , \38433 );
xor \U$38182 ( \38435 , \34869 , \34888 );
xor \U$38183 ( \38436 , \38435 , \34878 );
xor \U$38184 ( \38437 , \34912 , \34924 );
xor \U$38185 ( \38438 , \38437 , \34902 );
xor \U$38186 ( \38439 , \38436 , \38438 );
and \U$38187 ( \38440 , \35035 , \35020 );
not \U$38188 ( \38441 , \35035 );
and \U$38189 ( \38442 , \38441 , \35021 );
or \U$38190 ( \38443 , \38440 , \38442 );
and \U$38191 ( \38444 , \38443 , \35013 );
not \U$38192 ( \38445 , \38443 );
and \U$38193 ( \38446 , \38445 , \35012 );
nor \U$38194 ( \38447 , \38444 , \38446 );
and \U$38195 ( \38448 , \38439 , \38447 );
and \U$38196 ( \38449 , \38436 , \38438 );
or \U$38197 ( \38450 , \38448 , \38449 );
and \U$38198 ( \38451 , \38434 , \38450 );
and \U$38199 ( \38452 , \38418 , \38433 );
or \U$38200 ( \38453 , \38451 , \38452 );
nand \U$38201 ( \38454 , \38391 , \38453 );
nand \U$38202 ( \38455 , \38390 , \38454 );
not \U$38203 ( \38456 , \35217 );
not \U$38204 ( \38457 , \35193 );
or \U$38205 ( \38458 , \38456 , \38457 );
nand \U$38206 ( \38459 , \35192 , \35203 );
nand \U$38207 ( \38460 , \38458 , \38459 );
and \U$38208 ( \38461 , \38460 , \35214 );
not \U$38209 ( \38462 , \38460 );
not \U$38210 ( \38463 , \35214 );
and \U$38211 ( \38464 , \38462 , \38463 );
nor \U$38212 ( \38465 , \38461 , \38464 );
not \U$38213 ( \38466 , \35246 );
not \U$38214 ( \38467 , \35234 );
or \U$38215 ( \38468 , \38466 , \38467 );
not \U$38216 ( \38469 , \35246 );
nand \U$38217 ( \38470 , \38469 , \35223 );
nand \U$38218 ( \38471 , \38468 , \38470 );
and \U$38219 ( \38472 , \38471 , \35230 );
not \U$38220 ( \38473 , \38471 );
and \U$38221 ( \38474 , \38473 , \35229 );
nor \U$38222 ( \38475 , \38472 , \38474 );
or \U$38223 ( \38476 , \38465 , \38475 );
and \U$38224 ( \38477 , \35271 , \35274 );
not \U$38225 ( \38478 , \35271 );
and \U$38226 ( \38479 , \38478 , \35275 );
or \U$38227 ( \38480 , \38477 , \38479 );
not \U$38228 ( \38481 , \35261 );
and \U$38229 ( \38482 , \38480 , \38481 );
not \U$38230 ( \38483 , \38480 );
and \U$38231 ( \38484 , \38483 , \35261 );
nor \U$38232 ( \38485 , \38482 , \38484 );
nand \U$38233 ( \38486 , \38476 , \38485 );
nand \U$38234 ( \38487 , \38475 , \38465 );
nand \U$38235 ( \38488 , \38486 , \38487 );
xor \U$38236 ( \38489 , \35149 , \35180 );
xnor \U$38237 ( \38490 , \38489 , \35147 );
not \U$38238 ( \38491 , \34860 );
and \U$38239 ( \38492 , \34926 , \34891 );
not \U$38240 ( \38493 , \34926 );
and \U$38241 ( \38494 , \38493 , \34892 );
nor \U$38242 ( \38495 , \38492 , \38494 );
not \U$38243 ( \38496 , \38495 );
or \U$38244 ( \38497 , \38491 , \38496 );
or \U$38245 ( \38498 , \38495 , \34860 );
nand \U$38246 ( \38499 , \38497 , \38498 );
xor \U$38247 ( \38500 , \38490 , \38499 );
xor \U$38248 ( \38501 , \34963 , \35001 );
xor \U$38249 ( \38502 , \38501 , \35037 );
and \U$38250 ( \38503 , \38500 , \38502 );
and \U$38251 ( \38504 , \38490 , \38499 );
or \U$38252 ( \38505 , \38503 , \38504 );
xor \U$38253 ( \38506 , \38488 , \38505 );
not \U$38254 ( \38507 , \34789 );
not \U$38255 ( \38508 , \34786 );
or \U$38256 ( \38509 , \38507 , \38508 );
not \U$38257 ( \38510 , \34789 );
nand \U$38258 ( \38511 , \38510 , \34785 );
nand \U$38259 ( \38512 , \38509 , \38511 );
buf \U$38260 ( \38513 , \34781 );
not \U$38261 ( \38514 , \38513 );
and \U$38262 ( \38515 , \38512 , \38514 );
not \U$38263 ( \38516 , \38512 );
and \U$38264 ( \38517 , \38516 , \38513 );
nor \U$38265 ( \38518 , \38515 , \38517 );
and \U$38266 ( \38519 , \38506 , \38518 );
and \U$38267 ( \38520 , \38488 , \38505 );
or \U$38268 ( \38521 , \38519 , \38520 );
xor \U$38269 ( \38522 , \38455 , \38521 );
not \U$38270 ( \38523 , \35249 );
not \U$38271 ( \38524 , \35220 );
or \U$38272 ( \38525 , \38523 , \38524 );
not \U$38273 ( \38526 , \35249 );
nand \U$38274 ( \38527 , \38526 , \35219 );
nand \U$38275 ( \38528 , \38525 , \38527 );
not \U$38276 ( \38529 , \38528 );
not \U$38277 ( \38530 , \35183 );
or \U$38278 ( \38531 , \38529 , \38530 );
or \U$38279 ( \38532 , \38528 , \35183 );
nand \U$38280 ( \38533 , \38531 , \38532 );
xor \U$38281 ( \38534 , \35278 , \35283 );
not \U$38282 ( \38535 , \38534 );
not \U$38283 ( \38536 , \35295 );
or \U$38284 ( \38537 , \38535 , \38536 );
or \U$38285 ( \38538 , \38534 , \35295 );
nand \U$38286 ( \38539 , \38537 , \38538 );
xor \U$38287 ( \38540 , \38533 , \38539 );
xor \U$38288 ( \38541 , \34810 , \34820 );
xnor \U$38289 ( \38542 , \38541 , \34807 );
and \U$38290 ( \38543 , \38540 , \38542 );
and \U$38291 ( \38544 , \38533 , \38539 );
or \U$38292 ( \38545 , \38543 , \38544 );
and \U$38293 ( \38546 , \38522 , \38545 );
and \U$38294 ( \38547 , \38455 , \38521 );
or \U$38295 ( \38548 , \38546 , \38547 );
nand \U$38296 ( \38549 , \38266 , \38548 );
nand \U$38297 ( \38550 , \38262 , \38549 );
xor \U$38298 ( \38551 , \38236 , \38550 );
not \U$38299 ( \38552 , \35372 );
not \U$38300 ( \38553 , \35375 );
or \U$38301 ( \38554 , \38552 , \38553 );
or \U$38302 ( \38555 , \35375 , \35372 );
nand \U$38303 ( \38556 , \38554 , \38555 );
and \U$38304 ( \38557 , \38551 , \38556 );
and \U$38305 ( \38558 , \38236 , \38550 );
or \U$38306 ( \38559 , \38557 , \38558 );
nand \U$38307 ( \38560 , \38226 , \38559 );
nand \U$38308 ( \38561 , \38224 , \38225 );
nand \U$38309 ( \38562 , \38560 , \38561 );
not \U$38310 ( \38563 , \35945 );
xor \U$38311 ( \38564 , \35379 , \34294 );
not \U$38312 ( \38565 , \38564 );
not \U$38313 ( \38566 , \38565 );
or \U$38314 ( \38567 , \38563 , \38566 );
nand \U$38315 ( \38568 , \38564 , \35944 );
nand \U$38316 ( \38569 , \38567 , \38568 );
xor \U$38317 ( \38570 , \38562 , \38569 );
xor \U$38318 ( \38571 , \38206 , \38208 );
xor \U$38319 ( \38572 , \38571 , \38213 );
nand \U$38320 ( \38573 , \37094 , \36558 );
and \U$38321 ( \38574 , \38572 , \38573 );
not \U$38322 ( \38575 , \38572 );
not \U$38323 ( \38576 , \38573 );
and \U$38324 ( \38577 , \38575 , \38576 );
nor \U$38325 ( \38578 , \38574 , \38577 );
nand \U$38326 ( \38579 , \38222 , \38570 , \38578 );
nor \U$38327 ( \38580 , \37105 , \38579 );
xor \U$38328 ( \38581 , \34797 , \34792 );
xor \U$38329 ( \38582 , \38581 , \34826 );
nand \U$38330 ( \38583 , \30750 , \30686 );
and \U$38331 ( \38584 , \38583 , \30722 );
nor \U$38332 ( \38585 , \30750 , \30686 );
nor \U$38333 ( \38586 , \38584 , \38585 );
and \U$38334 ( \38587 , \31087 , \31043 );
nor \U$38335 ( \38588 , \38587 , \31008 );
nor \U$38336 ( \38589 , \31043 , \31087 );
nor \U$38337 ( \38590 , \38588 , \38589 );
xor \U$38338 ( \38591 , \38586 , \38590 );
xor \U$38339 ( \38592 , \30812 , \30840 );
and \U$38340 ( \38593 , \38592 , \30872 );
and \U$38341 ( \38594 , \30812 , \30840 );
or \U$38342 ( \38595 , \38593 , \38594 );
and \U$38343 ( \38596 , \38591 , \38595 );
and \U$38344 ( \38597 , \38586 , \38590 );
or \U$38345 ( \38598 , \38596 , \38597 );
not \U$38346 ( \38599 , \30602 );
not \U$38347 ( \38600 , \30594 );
or \U$38348 ( \38601 , \38599 , \38600 );
or \U$38349 ( \38602 , \30594 , \30602 );
nand \U$38350 ( \38603 , \38602 , \30608 );
nand \U$38351 ( \38604 , \38601 , \38603 );
not \U$38352 ( \38605 , \38604 );
not \U$38353 ( \38606 , \30662 );
not \U$38354 ( \38607 , \30667 );
or \U$38355 ( \38608 , \38606 , \38607 );
nand \U$38356 ( \38609 , \38608 , \30673 );
or \U$38357 ( \38610 , \30662 , \30667 );
nand \U$38358 ( \38611 , \38609 , \38610 );
not \U$38359 ( \38612 , \38611 );
and \U$38360 ( \38613 , \38605 , \38612 );
not \U$38361 ( \38614 , \30761 );
not \U$38362 ( \38615 , \30757 );
or \U$38363 ( \38616 , \38614 , \38615 );
nand \U$38364 ( \38617 , \38616 , \30773 );
not \U$38365 ( \38618 , \30757 );
nand \U$38366 ( \38619 , \38618 , \30762 );
and \U$38367 ( \38620 , \38617 , \38619 );
nor \U$38368 ( \38621 , \38613 , \38620 );
nor \U$38369 ( \38622 , \38605 , \38612 );
nor \U$38370 ( \38623 , \38621 , \38622 );
nand \U$38371 ( \38624 , \38598 , \38623 );
not \U$38372 ( \38625 , \38378 );
not \U$38373 ( \38626 , \38381 );
or \U$38374 ( \38627 , \38625 , \38626 );
or \U$38375 ( \38628 , \38381 , \38378 );
nand \U$38376 ( \38629 , \38627 , \38628 );
xor \U$38377 ( \38630 , \30909 , \30941 );
and \U$38378 ( \38631 , \38630 , \30972 );
and \U$38379 ( \38632 , \30909 , \30941 );
or \U$38380 ( \38633 , \38631 , \38632 );
xor \U$38381 ( \38634 , \38629 , \38633 );
xor \U$38382 ( \38635 , \38353 , \38356 );
xnor \U$38383 ( \38636 , \38635 , \38368 );
and \U$38384 ( \38637 , \38634 , \38636 );
and \U$38385 ( \38638 , \38629 , \38633 );
or \U$38386 ( \38639 , \38637 , \38638 );
and \U$38387 ( \38640 , \38624 , \38639 );
nor \U$38388 ( \38641 , \38623 , \38598 );
nor \U$38389 ( \38642 , \38640 , \38641 );
not \U$38390 ( \38643 , \38642 );
not \U$38391 ( \38644 , \38643 );
not \U$38392 ( \38645 , \38326 );
not \U$38393 ( \38646 , \38338 );
or \U$38394 ( \38647 , \38645 , \38646 );
not \U$38395 ( \38648 , \38326 );
nand \U$38396 ( \38649 , \38648 , \38337 );
nand \U$38397 ( \38650 , \38647 , \38649 );
not \U$38398 ( \38651 , \38650 );
not \U$38399 ( \38652 , \38331 );
and \U$38400 ( \38653 , \38651 , \38652 );
and \U$38401 ( \38654 , \38650 , \38331 );
nor \U$38402 ( \38655 , \38653 , \38654 );
not \U$38403 ( \38656 , \38655 );
xor \U$38404 ( \38657 , \38272 , \38277 );
xnor \U$38405 ( \38658 , \38657 , \38284 );
not \U$38406 ( \38659 , \38658 );
or \U$38407 ( \38660 , \38656 , \38659 );
not \U$38408 ( \38661 , \38294 );
not \U$38409 ( \38662 , \38308 );
or \U$38410 ( \38663 , \38661 , \38662 );
nand \U$38411 ( \38664 , \38303 , \38306 );
nand \U$38412 ( \38665 , \38663 , \38664 );
not \U$38413 ( \38666 , \38665 );
not \U$38414 ( \38667 , \38315 );
and \U$38415 ( \38668 , \38666 , \38667 );
and \U$38416 ( \38669 , \38665 , \38315 );
nor \U$38417 ( \38670 , \38668 , \38669 );
not \U$38418 ( \38671 , \38670 );
nand \U$38419 ( \38672 , \38660 , \38671 );
not \U$38420 ( \38673 , \38658 );
not \U$38421 ( \38674 , \38655 );
nand \U$38422 ( \38675 , \38673 , \38674 );
and \U$38423 ( \38676 , \38672 , \38675 );
and \U$38424 ( \38677 , \35137 , \35104 );
not \U$38425 ( \38678 , \35137 );
and \U$38426 ( \38679 , \38678 , \35140 );
or \U$38427 ( \38680 , \38677 , \38679 );
xor \U$38428 ( \38681 , \38680 , \35072 );
nand \U$38429 ( \38682 , \38676 , \38681 );
xor \U$38430 ( \38683 , \38405 , \38416 );
xnor \U$38431 ( \38684 , \38683 , \38397 );
not \U$38432 ( \38685 , \38684 );
xor \U$38433 ( \38686 , \38425 , \38427 );
xor \U$38434 ( \38687 , \38686 , \38430 );
not \U$38435 ( \38688 , \38687 );
not \U$38436 ( \38689 , \38688 );
or \U$38437 ( \38690 , \38685 , \38689 );
xor \U$38438 ( \38691 , \38436 , \38438 );
xor \U$38439 ( \38692 , \38691 , \38447 );
nand \U$38440 ( \38693 , \38690 , \38692 );
not \U$38441 ( \38694 , \38684 );
nand \U$38442 ( \38695 , \38687 , \38694 );
nand \U$38443 ( \38696 , \38693 , \38695 );
and \U$38444 ( \38697 , \38682 , \38696 );
nor \U$38445 ( \38698 , \38676 , \38681 );
nor \U$38446 ( \38699 , \38697 , \38698 );
not \U$38447 ( \38700 , \38699 );
not \U$38448 ( \38701 , \38700 );
or \U$38449 ( \38702 , \38644 , \38701 );
not \U$38450 ( \38703 , \38382 );
not \U$38451 ( \38704 , \38375 );
and \U$38452 ( \38705 , \38703 , \38704 );
and \U$38453 ( \38706 , \38382 , \38375 );
nor \U$38454 ( \38707 , \38705 , \38706 );
and \U$38455 ( \38708 , \38707 , \38373 );
not \U$38456 ( \38709 , \38707 );
not \U$38457 ( \38710 , \38373 );
and \U$38458 ( \38711 , \38709 , \38710 );
nor \U$38459 ( \38712 , \38708 , \38711 );
not \U$38460 ( \38713 , \38712 );
xor \U$38461 ( \38714 , \38490 , \38499 );
xor \U$38462 ( \38715 , \38714 , \38502 );
not \U$38463 ( \38716 , \38715 );
not \U$38464 ( \38717 , \38716 );
or \U$38465 ( \38718 , \38713 , \38717 );
not \U$38466 ( \38719 , \38485 );
not \U$38467 ( \38720 , \38719 );
not \U$38468 ( \38721 , \38475 );
or \U$38469 ( \38722 , \38720 , \38721 );
not \U$38470 ( \38723 , \38475 );
nand \U$38471 ( \38724 , \38723 , \38485 );
nand \U$38472 ( \38725 , \38722 , \38724 );
buf \U$38473 ( \38726 , \38465 );
and \U$38474 ( \38727 , \38725 , \38726 );
not \U$38475 ( \38728 , \38725 );
not \U$38476 ( \38729 , \38726 );
and \U$38477 ( \38730 , \38728 , \38729 );
nor \U$38478 ( \38731 , \38727 , \38730 );
nand \U$38479 ( \38732 , \38718 , \38731 );
not \U$38480 ( \38733 , \38712 );
nand \U$38481 ( \38734 , \38733 , \38715 );
nand \U$38482 ( \38735 , \38732 , \38734 );
nand \U$38483 ( \38736 , \38642 , \38699 );
nand \U$38484 ( \38737 , \38735 , \38736 );
nand \U$38485 ( \38738 , \38702 , \38737 );
xor \U$38486 ( \38739 , \38582 , \38738 );
not \U$38487 ( \38740 , \34929 );
not \U$38488 ( \38741 , \35040 );
not \U$38489 ( \38742 , \35142 );
or \U$38490 ( \38743 , \38741 , \38742 );
or \U$38491 ( \38744 , \35142 , \35040 );
nand \U$38492 ( \38745 , \38743 , \38744 );
not \U$38493 ( \38746 , \38745 );
or \U$38494 ( \38747 , \38740 , \38746 );
or \U$38495 ( \38748 , \38745 , \34929 );
nand \U$38496 ( \38749 , \38747 , \38748 );
xor \U$38497 ( \38750 , \38488 , \38505 );
xor \U$38498 ( \38751 , \38750 , \38518 );
xor \U$38499 ( \38752 , \38749 , \38751 );
xor \U$38500 ( \38753 , \38533 , \38539 );
xor \U$38501 ( \38754 , \38753 , \38542 );
and \U$38502 ( \38755 , \38752 , \38754 );
and \U$38503 ( \38756 , \38749 , \38751 );
or \U$38504 ( \38757 , \38755 , \38756 );
and \U$38505 ( \38758 , \38739 , \38757 );
and \U$38506 ( \38759 , \38582 , \38738 );
or \U$38507 ( \38760 , \38758 , \38759 );
xor \U$38508 ( \38761 , \35344 , \35359 );
xor \U$38509 ( \38762 , \38761 , \35362 );
xor \U$38510 ( \38763 , \38760 , \38762 );
buf \U$38511 ( \38764 , \35252 );
xor \U$38512 ( \38765 , \35298 , \38764 );
xor \U$38513 ( \38766 , \38765 , \35145 );
and \U$38514 ( \38767 , \38248 , \38251 );
not \U$38515 ( \38768 , \38248 );
and \U$38516 ( \38769 , \38768 , \38254 );
nor \U$38517 ( \38770 , \38767 , \38769 );
not \U$38518 ( \38771 , \38770 );
not \U$38519 ( \38772 , \38246 );
or \U$38520 ( \38773 , \38771 , \38772 );
or \U$38521 ( \38774 , \38246 , \38770 );
nand \U$38522 ( \38775 , \38773 , \38774 );
xor \U$38523 ( \38776 , \38766 , \38775 );
xor \U$38524 ( \38777 , \38455 , \38521 );
xor \U$38525 ( \38778 , \38777 , \38545 );
and \U$38526 ( \38779 , \38776 , \38778 );
and \U$38527 ( \38780 , \38766 , \38775 );
or \U$38528 ( \38781 , \38779 , \38780 );
and \U$38529 ( \38782 , \38763 , \38781 );
and \U$38530 ( \38783 , \38760 , \38762 );
or \U$38531 ( \38784 , \38782 , \38783 );
not \U$38532 ( \38785 , \38784 );
xor \U$38533 ( \38786 , \34828 , \35302 );
xnor \U$38534 ( \38787 , \38786 , \35331 );
not \U$38535 ( \38788 , \38787 );
and \U$38536 ( \38789 , \38548 , \38263 );
not \U$38537 ( \38790 , \38548 );
and \U$38538 ( \38791 , \38790 , \38260 );
or \U$38539 ( \38792 , \38789 , \38791 );
xnor \U$38540 ( \38793 , \38256 , \38792 );
nand \U$38541 ( \38794 , \38788 , \38793 );
nand \U$38542 ( \38795 , \38785 , \38794 );
xor \U$38543 ( \38796 , \38236 , \38550 );
xor \U$38544 ( \38797 , \38796 , \38556 );
and \U$38545 ( \38798 , \38795 , \38797 );
not \U$38546 ( \38799 , \38794 );
and \U$38547 ( \38800 , \38799 , \38784 );
nor \U$38548 ( \38801 , \38798 , \38800 );
xor \U$38549 ( \38802 , \38559 , \38225 );
not \U$38550 ( \38803 , \38224 );
and \U$38551 ( \38804 , \38802 , \38803 );
not \U$38552 ( \38805 , \38802 );
and \U$38553 ( \38806 , \38805 , \38224 );
nor \U$38554 ( \38807 , \38804 , \38806 );
xnor \U$38555 ( \38808 , \38801 , \38807 );
not \U$38556 ( \38809 , \38134 );
nand \U$38557 ( \38810 , \38809 , \38180 );
and \U$38558 ( \38811 , \38810 , \38156 );
nor \U$38559 ( \38812 , \38809 , \38180 );
nor \U$38560 ( \38813 , \38811 , \38812 );
not \U$38561 ( \38814 , \38813 );
not \U$38562 ( \38815 , \37589 );
not \U$38563 ( \38816 , \37613 );
or \U$38564 ( \38817 , \38815 , \38816 );
nand \U$38565 ( \38818 , \38817 , \38129 );
not \U$38566 ( \38819 , \37589 );
nand \U$38567 ( \38820 , \38819 , \37616 );
and \U$38568 ( \38821 , \38818 , \38820 );
not \U$38569 ( \38822 , \37637 );
not \U$38570 ( \38823 , \37647 );
or \U$38571 ( \38824 , \38822 , \38823 );
nand \U$38572 ( \38825 , \38824 , \37627 );
not \U$38573 ( \38826 , \37647 );
nand \U$38574 ( \38827 , \38826 , \37636 );
nand \U$38575 ( \38828 , \38825 , \38827 );
xor \U$38576 ( \38829 , \37688 , \37695 );
and \U$38577 ( \38830 , \38829 , \37700 );
and \U$38578 ( \38831 , \37688 , \37695 );
or \U$38579 ( \38832 , \38830 , \38831 );
xor \U$38580 ( \38833 , \38828 , \38832 );
not \U$38581 ( \38834 , \37661 );
not \U$38582 ( \38835 , \37656 );
or \U$38583 ( \38836 , \38834 , \38835 );
not \U$38584 ( \38837 , \37670 );
not \U$38585 ( \38838 , \37656 );
nand \U$38586 ( \38839 , \38838 , \37662 );
nand \U$38587 ( \38840 , \38837 , \38839 );
nand \U$38588 ( \38841 , \38836 , \38840 );
xor \U$38589 ( \38842 , \38833 , \38841 );
not \U$38590 ( \38843 , \37741 );
and \U$38591 ( \38844 , \37849 , \38843 );
nor \U$38592 ( \38845 , \38844 , \37971 );
nor \U$38593 ( \38846 , \37849 , \38843 );
nor \U$38594 ( \38847 , \38845 , \38846 );
not \U$38595 ( \38848 , \38847 );
xor \U$38596 ( \38849 , \38065 , \38074 );
and \U$38597 ( \38850 , \38849 , \38082 );
and \U$38598 ( \38851 , \38065 , \38074 );
or \U$38599 ( \38852 , \38850 , \38851 );
not \U$38600 ( \38853 , \37760 );
not \U$38601 ( \38854 , \37751 );
not \U$38602 ( \38855 , \38854 );
or \U$38603 ( \38856 , \38853 , \38855 );
or \U$38604 ( \38857 , \38854 , \37760 );
nand \U$38605 ( \38858 , \38857 , \37770 );
nand \U$38606 ( \38859 , \38856 , \38858 );
xor \U$38607 ( \38860 , \38852 , \38859 );
nand \U$38608 ( \38861 , \38054 , \38034 );
not \U$38609 ( \38862 , \38861 );
not \U$38610 ( \38863 , \38044 );
or \U$38611 ( \38864 , \38862 , \38863 );
or \U$38612 ( \38865 , \38034 , \38054 );
nand \U$38613 ( \38866 , \38864 , \38865 );
not \U$38614 ( \38867 , \38866 );
and \U$38615 ( \38868 , \38860 , \38867 );
not \U$38616 ( \38869 , \38860 );
and \U$38617 ( \38870 , \38869 , \38866 );
nor \U$38618 ( \38871 , \38868 , \38870 );
not \U$38619 ( \38872 , \38871 );
not \U$38620 ( \38873 , \38872 );
nand \U$38621 ( \38874 , \37675 , \37651 );
nand \U$38622 ( \38875 , \37701 , \38874 );
or \U$38623 ( \38876 , \37675 , \37651 );
and \U$38624 ( \38877 , \38875 , \38876 );
not \U$38625 ( \38878 , \38877 );
or \U$38626 ( \38879 , \38873 , \38878 );
not \U$38627 ( \38880 , \38876 );
not \U$38628 ( \38881 , \38875 );
or \U$38629 ( \38882 , \38880 , \38881 );
nand \U$38630 ( \38883 , \38882 , \38871 );
nand \U$38631 ( \38884 , \38879 , \38883 );
not \U$38632 ( \38885 , \38884 );
or \U$38633 ( \38886 , \38848 , \38885 );
or \U$38634 ( \38887 , \38884 , \38847 );
nand \U$38635 ( \38888 , \38886 , \38887 );
xor \U$38636 ( \38889 , \38842 , \38888 );
and \U$38637 ( \38890 , \37740 , \37714 );
not \U$38638 ( \38891 , \37740 );
not \U$38639 ( \38892 , \37714 );
and \U$38640 ( \38893 , \38891 , \38892 );
nor \U$38641 ( \38894 , \38890 , \38893 );
nand \U$38642 ( \38895 , \38894 , \37704 );
not \U$38643 ( \38896 , \37879 );
not \U$38644 ( \38897 , \37969 );
or \U$38645 ( \38898 , \38896 , \38897 );
not \U$38646 ( \38899 , \37966 );
not \U$38647 ( \38900 , \37880 );
or \U$38648 ( \38901 , \38899 , \38900 );
not \U$38649 ( \38902 , \37920 );
nand \U$38650 ( \38903 , \38901 , \38902 );
nand \U$38651 ( \38904 , \38898 , \38903 );
xor \U$38652 ( \38905 , \38895 , \38904 );
not \U$38653 ( \38906 , \37844 );
not \U$38654 ( \38907 , \37771 );
or \U$38655 ( \38908 , \38906 , \38907 );
nand \U$38656 ( \38909 , \38908 , \37801 );
not \U$38657 ( \38910 , \37771 );
nand \U$38658 ( \38911 , \38910 , \37847 );
nand \U$38659 ( \38912 , \38909 , \38911 );
xor \U$38660 ( \38913 , \38905 , \38912 );
not \U$38661 ( \38914 , \37714 );
not \U$38662 ( \38915 , \37735 );
or \U$38663 ( \38916 , \38914 , \38915 );
nand \U$38664 ( \38917 , \38916 , \37725 );
nand \U$38665 ( \38918 , \37738 , \38892 );
nand \U$38666 ( \38919 , \38917 , \38918 );
xor \U$38667 ( \38920 , \37859 , \37868 );
and \U$38668 ( \38921 , \38920 , \37878 );
and \U$38669 ( \38922 , \37859 , \37868 );
or \U$38670 ( \38923 , \38921 , \38922 );
xor \U$38671 ( \38924 , \38919 , \38923 );
not \U$38672 ( \38925 , \37947 );
not \U$38673 ( \38926 , \37961 );
or \U$38674 ( \38927 , \38925 , \38926 );
nand \U$38675 ( \38928 , \38927 , \37936 );
nand \U$38676 ( \38929 , \37964 , \37946 );
nand \U$38677 ( \38930 , \38928 , \38929 );
xor \U$38678 ( \38931 , \38924 , \38930 );
not \U$38679 ( \38932 , \37915 );
not \U$38680 ( \38933 , \37900 );
or \U$38681 ( \38934 , \38932 , \38933 );
nand \U$38682 ( \38935 , \38934 , \37890 );
nand \U$38683 ( \38936 , \37903 , \37918 );
nand \U$38684 ( \38937 , \38935 , \38936 );
xor \U$38685 ( \38938 , \37781 , \37790 );
and \U$38686 ( \38939 , \38938 , \37800 );
and \U$38687 ( \38940 , \37781 , \37790 );
or \U$38688 ( \38941 , \38939 , \38940 );
xor \U$38689 ( \38942 , \38937 , \38941 );
not \U$38690 ( \38943 , \37815 );
not \U$38691 ( \38944 , \37839 );
or \U$38692 ( \38945 , \38943 , \38944 );
nand \U$38693 ( \38946 , \38945 , \37826 );
not \U$38694 ( \38947 , \37815 );
nand \U$38695 ( \38948 , \38947 , \37842 );
nand \U$38696 ( \38949 , \38946 , \38948 );
xor \U$38697 ( \38950 , \38942 , \38949 );
xor \U$38698 ( \38951 , \38931 , \38950 );
and \U$38699 ( \38952 , RIbe29380_53, RIbe2a280_85);
not \U$38700 ( \38953 , RIbe2a370_87);
not \U$38701 ( \38954 , \546 );
or \U$38702 ( \38955 , \38953 , \38954 );
nand \U$38703 ( \38956 , \3775 , RIbe2a2f8_86);
nand \U$38704 ( \38957 , \38955 , \38956 );
and \U$38705 ( \38958 , \38957 , \1761 );
not \U$38706 ( \38959 , \38957 );
and \U$38707 ( \38960 , \38959 , \424 );
nor \U$38708 ( \38961 , \38958 , \38960 );
not \U$38709 ( \38962 , \38961 );
not \U$38710 ( \38963 , \38962 );
not \U$38711 ( \38964 , RIbe2acd0_107);
not \U$38712 ( \38965 , \32589 );
or \U$38713 ( \38966 , \38964 , \38965 );
nand \U$38714 ( \38967 , \1179 , RIbe2a028_80);
nand \U$38715 ( \38968 , \38966 , \38967 );
xor \U$38716 ( \38969 , \38968 , \564 );
not \U$38717 ( \38970 , \38969 );
not \U$38718 ( \38971 , \38970 );
or \U$38719 ( \38972 , \38963 , \38971 );
nand \U$38720 ( \38973 , \38961 , \38969 );
nand \U$38721 ( \38974 , \38972 , \38973 );
not \U$38722 ( \38975 , RIbe2b5b8_126);
not \U$38723 ( \38976 , \1223 );
or \U$38724 ( \38977 , \38975 , \38976 );
nand \U$38725 ( \38978 , \429 , RIbe2a3e8_88);
nand \U$38726 ( \38979 , \38977 , \38978 );
and \U$38727 ( \38980 , \38979 , \1232 );
not \U$38728 ( \38981 , \38979 );
and \U$38729 ( \38982 , \38981 , \306 );
nor \U$38730 ( \38983 , \38980 , \38982 );
xnor \U$38731 ( \38984 , \38974 , \38983 );
xor \U$38732 ( \38985 , \38952 , \38984 );
and \U$38733 ( \38986 , \261 , RIbe2a5c8_92);
and \U$38734 ( \38987 , \264 , RIbe2a550_91);
nor \U$38735 ( \38988 , \38986 , \38987 );
and \U$38736 ( \38989 , \38988 , \270 );
not \U$38737 ( \38990 , \38988 );
and \U$38738 ( \38991 , \38990 , \1663 );
nor \U$38739 ( \38992 , \38989 , \38991 );
and \U$38740 ( \38993 , \5365 , RIbe2a988_100);
and \U$38741 ( \38994 , \3897 , RIbe2a910_99);
nor \U$38742 ( \38995 , \38993 , \38994 );
and \U$38743 ( \38996 , \38995 , \293 );
not \U$38744 ( \38997 , \38995 );
and \U$38745 ( \38998 , \38997 , \300 );
nor \U$38746 ( \38999 , \38996 , \38998 );
and \U$38747 ( \39000 , \38992 , \38999 );
not \U$38748 ( \39001 , \38992 );
not \U$38749 ( \39002 , \38999 );
and \U$38750 ( \39003 , \39001 , \39002 );
or \U$38751 ( \39004 , \39000 , \39003 );
and \U$38752 ( \39005 , \3160 , RIbe2a208_84);
and \U$38753 ( \39006 , \330 , RIbe2a190_83);
nor \U$38754 ( \39007 , \39005 , \39006 );
and \U$38755 ( \39008 , \39007 , \1375 );
not \U$38756 ( \39009 , \39007 );
and \U$38757 ( \39010 , \39009 , \1379 );
nor \U$38758 ( \39011 , \39008 , \39010 );
not \U$38759 ( \39012 , \39011 );
xor \U$38760 ( \39013 , \39004 , \39012 );
xor \U$38761 ( \39014 , \38985 , \39013 );
xor \U$38762 ( \39015 , \38951 , \39014 );
xor \U$38763 ( \39016 , \38913 , \39015 );
xor \U$38764 ( \39017 , \12957 , \12769 );
and \U$38765 ( \39018 , \13049 , RIbe29920_65);
and \U$38766 ( \39019 , \12947 , RIbe27b98_2);
nor \U$38767 ( \39020 , \39018 , \39019 );
xnor \U$38768 ( \39021 , \39017 , \39020 );
not \U$38769 ( \39022 , RIbe28e58_42);
not \U$38770 ( \39023 , \13024 );
or \U$38771 ( \39024 , \39022 , \39023 );
nand \U$38772 ( \39025 , \12971 , RIbe28de0_41);
nand \U$38773 ( \39026 , \39024 , \39025 );
and \U$38774 ( \39027 , \39026 , \12219 );
not \U$38775 ( \39028 , \39026 );
and \U$38776 ( \39029 , \39028 , \9904 );
nor \U$38777 ( \39030 , \39027 , \39029 );
buf \U$38778 ( \39031 , \39030 );
xor \U$38779 ( \39032 , \39021 , \39031 );
not \U$38780 ( \39033 , \1157 );
not \U$38781 ( \39034 , RIbe29dd0_75);
not \U$38782 ( \39035 , \1142 );
or \U$38783 ( \39036 , \39034 , \39035 );
not \U$38784 ( \39037 , \9801 );
nand \U$38785 ( \39038 , \39037 , \1146 );
nand \U$38786 ( \39039 , \39036 , \39038 );
not \U$38787 ( \39040 , \39039 );
or \U$38788 ( \39041 , \39033 , \39040 );
or \U$38789 ( \39042 , \39039 , \1153 );
nand \U$38790 ( \39043 , \39041 , \39042 );
and \U$38791 ( \39044 , \1807 , RIbe29fb0_79);
and \U$38792 ( \39045 , \1165 , RIbe29e48_76);
nor \U$38793 ( \39046 , \39044 , \39045 );
and \U$38794 ( \39047 , \39046 , \1813 );
not \U$38795 ( \39048 , \39046 );
and \U$38796 ( \39049 , \39048 , \1010 );
nor \U$38797 ( \39050 , \39047 , \39049 );
xor \U$38798 ( \39051 , \39043 , \39050 );
not \U$38799 ( \39052 , RIbe29bf0_71);
not \U$38800 ( \39053 , \8868 );
or \U$38801 ( \39054 , \39052 , \39053 );
nand \U$38802 ( \39055 , \4730 , RIbe28f48_44);
nand \U$38803 ( \39056 , \39054 , \39055 );
and \U$38804 ( \39057 , \39056 , \1309 );
not \U$38805 ( \39058 , \39056 );
and \U$38806 ( \39059 , \39058 , \1082 );
nor \U$38807 ( \39060 , \39057 , \39059 );
xor \U$38808 ( \39061 , \39051 , \39060 );
not \U$38809 ( \39062 , RIbe28660_25);
not \U$38810 ( \39063 , \7827 );
or \U$38811 ( \39064 , \39062 , \39063 );
nand \U$38812 ( \39065 , \4284 , RIbe285e8_24);
nand \U$38813 ( \39066 , \39064 , \39065 );
and \U$38814 ( \39067 , \39066 , \4287 );
not \U$38815 ( \39068 , \39066 );
and \U$38816 ( \39069 , \39068 , \4783 );
nor \U$38817 ( \39070 , \39067 , \39069 );
not \U$38818 ( \39071 , \2889 );
not \U$38819 ( \39072 , \6347 );
and \U$38820 ( \39073 , \39071 , \39072 );
and \U$38821 ( \39074 , \27614 , RIbe27f58_10);
nor \U$38822 ( \39075 , \39073 , \39074 );
and \U$38823 ( \39076 , \39075 , \3516 );
not \U$38824 ( \39077 , \39075 );
and \U$38825 ( \39078 , \39077 , \1277 );
nor \U$38826 ( \39079 , \39076 , \39078 );
xor \U$38827 ( \39080 , \39070 , \39079 );
and \U$38828 ( \39081 , \1286 , RIbe28ed0_43);
and \U$38829 ( \39082 , \1117 , RIbe27fd0_11);
nor \U$38830 ( \39083 , \39081 , \39082 );
and \U$38831 ( \39084 , \39083 , \6831 );
not \U$38832 ( \39085 , \39083 );
and \U$38833 ( \39086 , \39085 , \1131 );
nor \U$38834 ( \39087 , \39084 , \39086 );
xor \U$38835 ( \39088 , \39080 , \39087 );
xor \U$38836 ( \39089 , \39061 , \39088 );
not \U$38837 ( \39090 , RIbe28408_20);
not \U$38838 ( \39091 , \7880 );
or \U$38839 ( \39092 , \39090 , \39091 );
nand \U$38840 ( \39093 , \4027 , RIbe28390_19);
nand \U$38841 ( \39094 , \39092 , \39093 );
and \U$38842 ( \39095 , \39094 , \3471 );
not \U$38843 ( \39096 , \39094 );
and \U$38844 ( \39097 , \39096 , \3448 );
nor \U$38845 ( \39098 , \39095 , \39097 );
not \U$38846 ( \39099 , \39098 );
not \U$38847 ( \39100 , \39099 );
not \U$38848 ( \39101 , RIbe28b10_35);
not \U$38849 ( \39102 , \5058 );
or \U$38850 ( \39103 , \39101 , \39102 );
nand \U$38851 ( \39104 , \4600 , RIbe28b88_36);
nand \U$38852 ( \39105 , \39103 , \39104 );
and \U$38853 ( \39106 , \39105 , \4323 );
not \U$38854 ( \39107 , \39105 );
and \U$38855 ( \39108 , \39107 , \4326 );
nor \U$38856 ( \39109 , \39106 , \39108 );
not \U$38857 ( \39110 , \39109 );
not \U$38858 ( \39111 , \39110 );
or \U$38859 ( \39112 , \39100 , \39111 );
nand \U$38860 ( \39113 , \39109 , \39098 );
nand \U$38861 ( \39114 , \39112 , \39113 );
not \U$38862 ( \39115 , RIbe287c8_28);
not \U$38863 ( \39116 , \3452 );
or \U$38864 ( \39117 , \39115 , \39116 );
nand \U$38865 ( \39118 , \3458 , RIbe28480_21);
nand \U$38866 ( \39119 , \39117 , \39118 );
and \U$38867 ( \39120 , \39119 , \3461 );
not \U$38868 ( \39121 , \39119 );
and \U$38869 ( \39122 , \39121 , \4346 );
nor \U$38870 ( \39123 , \39120 , \39122 );
not \U$38871 ( \39124 , \39123 );
and \U$38872 ( \39125 , \39114 , \39124 );
not \U$38873 ( \39126 , \39114 );
and \U$38874 ( \39127 , \39126 , \39123 );
nor \U$38875 ( \39128 , \39125 , \39127 );
xor \U$38876 ( \39129 , \39089 , \39128 );
xor \U$38877 ( \39130 , \39032 , \39129 );
not \U$38878 ( \39131 , RIbe29830_63);
not \U$38879 ( \39132 , \7274 );
or \U$38880 ( \39133 , \39131 , \39132 );
nand \U$38881 ( \39134 , \6596 , RIbe296c8_60);
nand \U$38882 ( \39135 , \39133 , \39134 );
and \U$38883 ( \39136 , \39135 , \7948 );
not \U$38884 ( \39137 , \39135 );
and \U$38885 ( \39138 , \39137 , \6602 );
nor \U$38886 ( \39139 , \39136 , \39138 );
not \U$38887 ( \39140 , RIbe29650_59);
not \U$38888 ( \39141 , \6958 );
or \U$38889 ( \39142 , \39140 , \39141 );
nand \U$38890 ( \39143 , \6963 , RIbe29038_46);
nand \U$38891 ( \39144 , \39142 , \39143 );
and \U$38892 ( \39145 , \39144 , \7293 );
not \U$38893 ( \39146 , \39144 );
and \U$38894 ( \39147 , \39146 , \6569 );
nor \U$38895 ( \39148 , \39145 , \39147 );
xor \U$38896 ( \39149 , \39139 , \39148 );
not \U$38897 ( \39150 , RIbe281b0_15);
not \U$38898 ( \39151 , \6536 );
or \U$38899 ( \39152 , \39150 , \39151 );
nand \U$38900 ( \39153 , \10348 , RIbe280c0_13);
nand \U$38901 ( \39154 , \39152 , \39153 );
and \U$38902 ( \39155 , \39154 , \15730 );
not \U$38903 ( \39156 , \39154 );
and \U$38904 ( \39157 , \39156 , \6891 );
nor \U$38905 ( \39158 , \39155 , \39157 );
xor \U$38906 ( \39159 , \39149 , \39158 );
and \U$38907 ( \39160 , \10916 , RIbe27d00_5);
and \U$38908 ( \39161 , \15228 , RIbe27c10_3);
nor \U$38909 ( \39162 , \39160 , \39161 );
and \U$38910 ( \39163 , \39162 , \16059 );
not \U$38911 ( \39164 , \39162 );
and \U$38912 ( \39165 , \39164 , \18797 );
nor \U$38913 ( \39166 , \39163 , \39165 );
not \U$38914 ( \39167 , RIbe29a88_68);
not \U$38915 ( \39168 , \10949 );
or \U$38916 ( \39169 , \39167 , \39168 );
nand \U$38917 ( \39170 , \10952 , RIbe27d78_6);
nand \U$38918 ( \39171 , \39169 , \39170 );
and \U$38919 ( \39172 , \39171 , \14299 );
not \U$38920 ( \39173 , \39171 );
and \U$38921 ( \39174 , \39173 , \7989 );
nor \U$38922 ( \39175 , \39172 , \39174 );
xor \U$38923 ( \39176 , \39166 , \39175 );
not \U$38924 ( \39177 , RIbe28fc0_45);
not \U$38925 ( \39178 , \7299 );
or \U$38926 ( \39179 , \39177 , \39178 );
nand \U$38927 ( \39180 , \9875 , RIbe290b0_47);
nand \U$38928 ( \39181 , \39179 , \39180 );
not \U$38929 ( \39182 , \39181 );
not \U$38930 ( \39183 , \6992 );
and \U$38931 ( \39184 , \39182 , \39183 );
and \U$38932 ( \39185 , \39181 , \6992 );
nor \U$38933 ( \39186 , \39184 , \39185 );
xnor \U$38934 ( \39187 , \39176 , \39186 );
xor \U$38935 ( \39188 , \39159 , \39187 );
not \U$38936 ( \39189 , \6624 );
not \U$38937 ( \39190 , RIbe29560_57);
not \U$38938 ( \39191 , \6856 );
or \U$38939 ( \39192 , \39190 , \39191 );
nand \U$38940 ( \39193 , \8235 , RIbe28228_16);
nand \U$38941 ( \39194 , \39192 , \39193 );
not \U$38942 ( \39195 , \39194 );
or \U$38943 ( \39196 , \39189 , \39195 );
or \U$38944 ( \39197 , \39194 , \9944 );
nand \U$38945 ( \39198 , \39196 , \39197 );
not \U$38946 ( \39199 , \39198 );
not \U$38947 ( \39200 , RIbe289a8_32);
not \U$38948 ( \39201 , \5455 );
or \U$38949 ( \39202 , \39200 , \39201 );
nand \U$38950 ( \39203 , \8247 , RIbe28930_31);
nand \U$38951 ( \39204 , \39202 , \39203 );
not \U$38952 ( \39205 , \39204 );
not \U$38953 ( \39206 , \6637 );
and \U$38954 ( \39207 , \39205 , \39206 );
and \U$38955 ( \39208 , \39204 , \5754 );
nor \U$38956 ( \39209 , \39207 , \39208 );
not \U$38957 ( \39210 , \39209 );
or \U$38958 ( \39211 , \39199 , \39210 );
or \U$38959 ( \39212 , \39209 , \39198 );
nand \U$38960 ( \39213 , \39211 , \39212 );
not \U$38961 ( \39214 , RIbe29290_51);
not \U$38962 ( \39215 , \4830 );
or \U$38963 ( \39216 , \39214 , \39215 );
nand \U$38964 ( \39217 , \5052 , RIbe28a20_33);
nand \U$38965 ( \39218 , \39216 , \39217 );
not \U$38966 ( \39219 , \39218 );
not \U$38967 ( \39220 , \4592 );
and \U$38968 ( \39221 , \39219 , \39220 );
and \U$38969 ( \39222 , \39218 , \4592 );
nor \U$38970 ( \39223 , \39221 , \39222 );
not \U$38971 ( \39224 , \39223 );
and \U$38972 ( \39225 , \39213 , \39224 );
not \U$38973 ( \39226 , \39213 );
and \U$38974 ( \39227 , \39226 , \39223 );
nor \U$38975 ( \39228 , \39225 , \39227 );
xor \U$38976 ( \39229 , \39188 , \39228 );
xor \U$38977 ( \39230 , \39130 , \39229 );
xor \U$38978 ( \39231 , \39016 , \39230 );
xor \U$38979 ( \39232 , \38889 , \39231 );
nor \U$38980 ( \39233 , \37990 , \37983 );
or \U$38981 ( \39234 , \37995 , \39233 );
nand \U$38982 ( \39235 , \37990 , \37983 );
nand \U$38983 ( \39236 , \39234 , \39235 );
not \U$38984 ( \39237 , \38031 );
not \U$38985 ( \39238 , \38100 );
not \U$38986 ( \39239 , \39238 );
or \U$38987 ( \39240 , \39237 , \39239 );
nand \U$38988 ( \39241 , \39240 , \38119 );
not \U$38989 ( \39242 , \38031 );
nand \U$38990 ( \39243 , \39242 , \38100 );
nand \U$38991 ( \39244 , \39241 , \39243 );
xor \U$38992 ( \39245 , \39236 , \39244 );
xor \U$38993 ( \39246 , \37622 , \37702 );
and \U$38994 ( \39247 , \39246 , \37972 );
and \U$38995 ( \39248 , \37622 , \37702 );
or \U$38996 ( \39249 , \39247 , \39248 );
xor \U$38997 ( \39250 , \39245 , \39249 );
not \U$38998 ( \39251 , \39250 );
and \U$38999 ( \39252 , \39232 , \39251 );
not \U$39000 ( \39253 , \39232 );
and \U$39001 ( \39254 , \39253 , \39250 );
nor \U$39002 ( \39255 , \39252 , \39254 );
not \U$39003 ( \39256 , \39255 );
and \U$39004 ( \39257 , \38821 , \39256 );
not \U$39005 ( \39258 , \38821 );
not \U$39006 ( \39259 , \39256 );
and \U$39007 ( \39260 , \39258 , \39259 );
or \U$39008 ( \39261 , \39257 , \39260 );
nor \U$39009 ( \39262 , \38026 , \38008 );
or \U$39010 ( \39263 , \39262 , \38017 );
nand \U$39011 ( \39264 , \38026 , \38008 );
nand \U$39012 ( \39265 , \39263 , \39264 );
not \U$39013 ( \39266 , \38083 );
nand \U$39014 ( \39267 , \39266 , \38055 );
not \U$39015 ( \39268 , \39267 );
not \U$39016 ( \39269 , \38096 );
or \U$39017 ( \39270 , \39268 , \39269 );
not \U$39018 ( \39271 , \38055 );
nand \U$39019 ( \39272 , \39271 , \38083 );
nand \U$39020 ( \39273 , \39270 , \39272 );
xor \U$39021 ( \39274 , \39265 , \39273 );
xor \U$39022 ( \39275 , \38108 , \38113 );
and \U$39023 ( \39276 , \39275 , \38118 );
and \U$39024 ( \39277 , \38108 , \38113 );
or \U$39025 ( \39278 , \39276 , \39277 );
xor \U$39026 ( \39279 , \39274 , \39278 );
nor \U$39027 ( \39280 , \38171 , \38162 );
or \U$39028 ( \39281 , \38176 , \39280 );
nand \U$39029 ( \39282 , \38171 , \38162 );
nand \U$39030 ( \39283 , \39281 , \39282 );
and \U$39031 ( \39284 , \39279 , \39283 );
not \U$39032 ( \39285 , \39279 );
not \U$39033 ( \39286 , \39283 );
and \U$39034 ( \39287 , \39285 , \39286 );
nor \U$39035 ( \39288 , \39284 , \39287 );
nand \U$39036 ( \39289 , \38124 , \38000 );
and \U$39037 ( \39290 , \37973 , \39289 );
nor \U$39038 ( \39291 , \38124 , \38000 );
nor \U$39039 ( \39292 , \39290 , \39291 );
xor \U$39040 ( \39293 , \39288 , \39292 );
and \U$39041 ( \39294 , \39261 , \39293 );
not \U$39042 ( \39295 , \39261 );
not \U$39043 ( \39296 , \39293 );
and \U$39044 ( \39297 , \39295 , \39296 );
nor \U$39045 ( \39298 , \39294 , \39297 );
not \U$39046 ( \39299 , \39298 );
not \U$39047 ( \39300 , \39299 );
or \U$39048 ( \39301 , \38814 , \39300 );
or \U$39049 ( \39302 , \39299 , \38813 );
nand \U$39050 ( \39303 , \39301 , \39302 );
not \U$39051 ( \39304 , \39303 );
not \U$39052 ( \39305 , \38198 );
nand \U$39053 ( \39306 , \39305 , \38183 );
not \U$39054 ( \39307 , \39306 );
and \U$39055 ( \39308 , \39304 , \39307 );
and \U$39056 ( \39309 , \39303 , \39306 );
nor \U$39057 ( \39310 , \39308 , \39309 );
nor \U$39058 ( \39311 , \38808 , \39310 );
and \U$39059 ( \39312 , \38580 , \39311 );
not \U$39060 ( \39313 , \39312 );
xor \U$39061 ( \39314 , \38318 , \38286 );
xor \U$39062 ( \39315 , \38341 , \39314 );
xor \U$39063 ( \39316 , \38418 , \38433 );
xor \U$39064 ( \39317 , \39316 , \38450 );
xor \U$39065 ( \39318 , \39315 , \39317 );
not \U$39066 ( \39319 , \38712 );
not \U$39067 ( \39320 , \38715 );
or \U$39068 ( \39321 , \39319 , \39320 );
or \U$39069 ( \39322 , \38715 , \38712 );
nand \U$39070 ( \39323 , \39321 , \39322 );
and \U$39071 ( \39324 , \39323 , \38731 );
not \U$39072 ( \39325 , \39323 );
not \U$39073 ( \39326 , \38731 );
and \U$39074 ( \39327 , \39325 , \39326 );
nor \U$39075 ( \39328 , \39324 , \39327 );
and \U$39076 ( \39329 , \39318 , \39328 );
and \U$39077 ( \39330 , \39315 , \39317 );
or \U$39078 ( \39331 , \39329 , \39330 );
not \U$39079 ( \39332 , \39331 );
not \U$39080 ( \39333 , \39332 );
xor \U$39081 ( \39334 , \38388 , \38343 );
xnor \U$39082 ( \39335 , \39334 , \38453 );
not \U$39083 ( \39336 , \39335 );
not \U$39084 ( \39337 , \39336 );
not \U$39085 ( \39338 , \31126 );
not \U$39086 ( \39339 , \31122 );
or \U$39087 ( \39340 , \39338 , \39339 );
nand \U$39088 ( \39341 , \39340 , \31118 );
not \U$39089 ( \39342 , \31122 );
nand \U$39090 ( \39343 , \39342 , \31129 );
nand \U$39091 ( \39344 , \39341 , \39343 );
not \U$39092 ( \39345 , \39344 );
not \U$39093 ( \39346 , \31104 );
not \U$39094 ( \39347 , \31100 );
or \U$39095 ( \39348 , \39346 , \39347 );
or \U$39096 ( \39349 , \31100 , \31104 );
nand \U$39097 ( \39350 , \39349 , \31113 );
nand \U$39098 ( \39351 , \39348 , \39350 );
not \U$39099 ( \39352 , \39351 );
and \U$39100 ( \39353 , \39345 , \39352 );
nand \U$39101 ( \39354 , \31092 , \30883 );
and \U$39102 ( \39355 , \39354 , \30973 );
nor \U$39103 ( \39356 , \31092 , \30883 );
nor \U$39104 ( \39357 , \39355 , \39356 );
nor \U$39105 ( \39358 , \39353 , \39357 );
nor \U$39106 ( \39359 , \39352 , \39345 );
nor \U$39107 ( \39360 , \39358 , \39359 );
xor \U$39108 ( \39361 , \38586 , \38590 );
xor \U$39109 ( \39362 , \39361 , \38595 );
not \U$39110 ( \39363 , \38604 );
not \U$39111 ( \39364 , \38620 );
or \U$39112 ( \39365 , \39363 , \39364 );
or \U$39113 ( \39366 , \38620 , \38604 );
nand \U$39114 ( \39367 , \39365 , \39366 );
and \U$39115 ( \39368 , \39367 , \38611 );
not \U$39116 ( \39369 , \39367 );
and \U$39117 ( \39370 , \39369 , \38612 );
nor \U$39118 ( \39371 , \39368 , \39370 );
not \U$39119 ( \39372 , \39371 );
nand \U$39120 ( \39373 , \39362 , \39372 );
xor \U$39121 ( \39374 , \38629 , \38633 );
xor \U$39122 ( \39375 , \39374 , \38636 );
and \U$39123 ( \39376 , \39373 , \39375 );
nor \U$39124 ( \39377 , \39372 , \39362 );
nor \U$39125 ( \39378 , \39376 , \39377 );
xor \U$39126 ( \39379 , \39360 , \39378 );
not \U$39127 ( \39380 , \38658 );
not \U$39128 ( \39381 , \38671 );
or \U$39129 ( \39382 , \39380 , \39381 );
nand \U$39130 ( \39383 , \38670 , \38673 );
nand \U$39131 ( \39384 , \39382 , \39383 );
and \U$39132 ( \39385 , \39384 , \38674 );
not \U$39133 ( \39386 , \39384 );
and \U$39134 ( \39387 , \39386 , \38655 );
nor \U$39135 ( \39388 , \39385 , \39387 );
not \U$39136 ( \39389 , \39388 );
and \U$39137 ( \39390 , \30873 , \30775 );
nor \U$39138 ( \39391 , \39390 , \30751 );
nor \U$39139 ( \39392 , \30775 , \30873 );
nor \U$39140 ( \39393 , \39391 , \39392 );
nand \U$39141 ( \39394 , \39389 , \39393 );
not \U$39142 ( \39395 , \38694 );
not \U$39143 ( \39396 , \38688 );
or \U$39144 ( \39397 , \39395 , \39396 );
nand \U$39145 ( \39398 , \38687 , \38684 );
nand \U$39146 ( \39399 , \39397 , \39398 );
xor \U$39147 ( \39400 , \39399 , \38692 );
and \U$39148 ( \39401 , \39394 , \39400 );
nor \U$39149 ( \39402 , \39389 , \39393 );
nor \U$39150 ( \39403 , \39401 , \39402 );
and \U$39151 ( \39404 , \39379 , \39403 );
and \U$39152 ( \39405 , \39360 , \39378 );
or \U$39153 ( \39406 , \39404 , \39405 );
not \U$39154 ( \39407 , \39406 );
or \U$39155 ( \39408 , \39337 , \39407 );
not \U$39156 ( \39409 , \39406 );
nand \U$39157 ( \39410 , \39409 , \39335 );
nand \U$39158 ( \39411 , \39408 , \39410 );
not \U$39159 ( \39412 , \39411 );
or \U$39160 ( \39413 , \39333 , \39412 );
or \U$39161 ( \39414 , \39411 , \39332 );
nand \U$39162 ( \39415 , \39413 , \39414 );
xor \U$39163 ( \39416 , \38700 , \38643 );
and \U$39164 ( \39417 , \39416 , \38735 );
not \U$39165 ( \39418 , \39416 );
not \U$39166 ( \39419 , \38735 );
and \U$39167 ( \39420 , \39418 , \39419 );
nor \U$39168 ( \39421 , \39417 , \39420 );
nand \U$39169 ( \39422 , \39415 , \39421 );
xor \U$39170 ( \39423 , \38676 , \38681 );
xor \U$39171 ( \39424 , \39423 , \38696 );
not \U$39172 ( \39425 , \30644 );
nand \U$39173 ( \39426 , \30639 , \39425 );
and \U$39174 ( \39427 , \39426 , \30653 );
nor \U$39175 ( \39428 , \30639 , \39425 );
nor \U$39176 ( \39429 , \39427 , \39428 );
not \U$39177 ( \39430 , \39429 );
nand \U$39178 ( \39431 , \30585 , \30609 );
and \U$39179 ( \39432 , \39431 , \30614 );
nor \U$39180 ( \39433 , \30585 , \30609 );
nor \U$39181 ( \39434 , \39432 , \39433 );
not \U$39182 ( \39435 , \39434 );
or \U$39183 ( \39436 , \39430 , \39435 );
xor \U$39184 ( \39437 , \30681 , \30878 );
and \U$39185 ( \39438 , \39437 , \31093 );
and \U$39186 ( \39439 , \30681 , \30878 );
or \U$39187 ( \39440 , \39438 , \39439 );
nand \U$39188 ( \39441 , \39436 , \39440 );
or \U$39189 ( \39442 , \39434 , \39429 );
nand \U$39190 ( \39443 , \39441 , \39442 );
xor \U$39191 ( \39444 , \39424 , \39443 );
not \U$39192 ( \39445 , \39344 );
not \U$39193 ( \39446 , \39352 );
and \U$39194 ( \39447 , \39445 , \39446 );
and \U$39195 ( \39448 , \39344 , \39352 );
nor \U$39196 ( \39449 , \39447 , \39448 );
xor \U$39197 ( \39450 , \39357 , \39449 );
not \U$39198 ( \39451 , \39375 );
xor \U$39199 ( \39452 , \39362 , \39371 );
not \U$39200 ( \39453 , \39452 );
or \U$39201 ( \39454 , \39451 , \39453 );
or \U$39202 ( \39455 , \39452 , \39375 );
nand \U$39203 ( \39456 , \39454 , \39455 );
xor \U$39204 ( \39457 , \39450 , \39456 );
not \U$39205 ( \39458 , \39400 );
not \U$39206 ( \39459 , \39388 );
not \U$39207 ( \39460 , \39393 );
and \U$39208 ( \39461 , \39459 , \39460 );
and \U$39209 ( \39462 , \39388 , \39393 );
nor \U$39210 ( \39463 , \39461 , \39462 );
not \U$39211 ( \39464 , \39463 );
or \U$39212 ( \39465 , \39458 , \39464 );
or \U$39213 ( \39466 , \39463 , \39400 );
nand \U$39214 ( \39467 , \39465 , \39466 );
and \U$39215 ( \39468 , \39457 , \39467 );
and \U$39216 ( \39469 , \39450 , \39456 );
or \U$39217 ( \39470 , \39468 , \39469 );
and \U$39218 ( \39471 , \39444 , \39470 );
and \U$39219 ( \39472 , \39424 , \39443 );
or \U$39220 ( \39473 , \39471 , \39472 );
not \U$39221 ( \39474 , \39473 );
xor \U$39222 ( \39475 , \38749 , \38751 );
xor \U$39223 ( \39476 , \39475 , \38754 );
not \U$39224 ( \39477 , \39476 );
and \U$39225 ( \39478 , \39474 , \39477 );
xor \U$39226 ( \39479 , \39315 , \39317 );
xor \U$39227 ( \39480 , \39479 , \39328 );
not \U$39228 ( \39481 , \39480 );
xor \U$39229 ( \39482 , \38598 , \38623 );
xnor \U$39230 ( \39483 , \39482 , \38639 );
nand \U$39231 ( \39484 , \39481 , \39483 );
xor \U$39232 ( \39485 , \39360 , \39378 );
xor \U$39233 ( \39486 , \39485 , \39403 );
not \U$39234 ( \39487 , \39486 );
and \U$39235 ( \39488 , \39484 , \39487 );
nor \U$39236 ( \39489 , \39481 , \39483 );
nor \U$39237 ( \39490 , \39488 , \39489 );
nor \U$39238 ( \39491 , \39478 , \39490 );
and \U$39239 ( \39492 , \39476 , \39473 );
nor \U$39240 ( \39493 , \39491 , \39492 );
xor \U$39241 ( \39494 , \39422 , \39493 );
xor \U$39242 ( \39495 , \38582 , \38738 );
xor \U$39243 ( \39496 , \39495 , \38757 );
not \U$39244 ( \39497 , \39409 );
not \U$39245 ( \39498 , \39336 );
or \U$39246 ( \39499 , \39497 , \39498 );
not \U$39247 ( \39500 , \39335 );
not \U$39248 ( \39501 , \39406 );
or \U$39249 ( \39502 , \39500 , \39501 );
nand \U$39250 ( \39503 , \39502 , \39331 );
nand \U$39251 ( \39504 , \39499 , \39503 );
and \U$39252 ( \39505 , \39496 , \39504 );
not \U$39253 ( \39506 , \39496 );
not \U$39254 ( \39507 , \39504 );
and \U$39255 ( \39508 , \39506 , \39507 );
nor \U$39256 ( \39509 , \39505 , \39508 );
xor \U$39257 ( \39510 , \38766 , \38775 );
xor \U$39258 ( \39511 , \39510 , \38778 );
xnor \U$39259 ( \39512 , \39509 , \39511 );
and \U$39260 ( \39513 , \39494 , \39512 );
and \U$39261 ( \39514 , \39422 , \39493 );
or \U$39262 ( \39515 , \39513 , \39514 );
not \U$39263 ( \39516 , \39515 );
not \U$39264 ( \39517 , \39516 );
xor \U$39265 ( \39518 , \38787 , \38257 );
xnor \U$39266 ( \39519 , \39518 , \38792 );
xor \U$39267 ( \39520 , \38760 , \38762 );
xor \U$39268 ( \39521 , \39520 , \38781 );
xor \U$39269 ( \39522 , \39519 , \39521 );
not \U$39270 ( \39523 , \39504 );
not \U$39271 ( \39524 , \39496 );
or \U$39272 ( \39525 , \39523 , \39524 );
not \U$39273 ( \39526 , \39496 );
nand \U$39274 ( \39527 , \39526 , \39507 );
nand \U$39275 ( \39528 , \39511 , \39527 );
nand \U$39276 ( \39529 , \39525 , \39528 );
xnor \U$39277 ( \39530 , \39522 , \39529 );
not \U$39278 ( \39531 , \39530 );
or \U$39279 ( \39532 , \39517 , \39531 );
xor \U$39280 ( \39533 , \39519 , \39521 );
xor \U$39281 ( \39534 , \39533 , \39529 );
nand \U$39282 ( \39535 , \39534 , \39515 );
nand \U$39283 ( \39536 , \39532 , \39535 );
xor \U$39284 ( \39537 , \39421 , \39332 );
xnor \U$39285 ( \39538 , \39537 , \39411 );
not \U$39286 ( \39539 , \39490 );
xor \U$39287 ( \39540 , \39476 , \39473 );
not \U$39288 ( \39541 , \39540 );
or \U$39289 ( \39542 , \39539 , \39541 );
or \U$39290 ( \39543 , \39490 , \39540 );
nand \U$39291 ( \39544 , \39542 , \39543 );
xor \U$39292 ( \39545 , \39538 , \39544 );
not \U$39293 ( \39546 , \31152 );
not \U$39294 ( \39547 , \31141 );
and \U$39295 ( \39548 , \39546 , \39547 );
nor \U$39296 ( \39549 , \39548 , \31147 );
nor \U$39297 ( \39550 , \39546 , \39547 );
nor \U$39298 ( \39551 , \39549 , \39550 );
not \U$39299 ( \39552 , \39551 );
not \U$39300 ( \39553 , \39552 );
or \U$39301 ( \39554 , \31132 , \31114 );
and \U$39302 ( \39555 , \31094 , \39554 );
and \U$39303 ( \39556 , \31114 , \31132 );
nor \U$39304 ( \39557 , \39555 , \39556 );
not \U$39305 ( \39558 , \39557 );
not \U$39306 ( \39559 , \39558 );
or \U$39307 ( \39560 , \39553 , \39559 );
xor \U$39308 ( \39561 , \39450 , \39456 );
xor \U$39309 ( \39562 , \39561 , \39467 );
nand \U$39310 ( \39563 , \39557 , \39551 );
nand \U$39311 ( \39564 , \39562 , \39563 );
nand \U$39312 ( \39565 , \39560 , \39564 );
xor \U$39313 ( \39566 , \39424 , \39443 );
xor \U$39314 ( \39567 , \39566 , \39470 );
xor \U$39315 ( \39568 , \39565 , \39567 );
xor \U$39316 ( \39569 , \39483 , \39480 );
xor \U$39317 ( \39570 , \39569 , \39486 );
and \U$39318 ( \39571 , \39568 , \39570 );
and \U$39319 ( \39572 , \39565 , \39567 );
or \U$39320 ( \39573 , \39571 , \39572 );
and \U$39321 ( \39574 , \39545 , \39573 );
and \U$39322 ( \39575 , \39538 , \39544 );
or \U$39323 ( \39576 , \39574 , \39575 );
not \U$39324 ( \39577 , \39576 );
xor \U$39325 ( \39578 , \39422 , \39493 );
xor \U$39326 ( \39579 , \39578 , \39512 );
not \U$39327 ( \39580 , \39579 );
or \U$39328 ( \39581 , \39577 , \39580 );
or \U$39329 ( \39582 , \39576 , \39579 );
nand \U$39330 ( \39583 , \39581 , \39582 );
nand \U$39331 ( \39584 , \39536 , \39583 );
not \U$39332 ( \39585 , \39584 );
xnor \U$39333 ( \39586 , \39434 , \39429 );
not \U$39334 ( \39587 , \39586 );
not \U$39335 ( \39588 , \39440 );
and \U$39336 ( \39589 , \39587 , \39588 );
and \U$39337 ( \39590 , \39586 , \39440 );
nor \U$39338 ( \39591 , \39589 , \39590 );
not \U$39339 ( \39592 , \30621 );
not \U$39340 ( \39593 , \30615 );
and \U$39341 ( \39594 , \39592 , \39593 );
nor \U$39342 ( \39595 , \39594 , \30579 );
and \U$39343 ( \39596 , \30615 , \30621 );
nor \U$39344 ( \39597 , \39595 , \39596 );
xor \U$39345 ( \39598 , \39591 , \39597 );
not \U$39346 ( \39599 , \31134 );
nand \U$39347 ( \39600 , \30657 , \39599 );
and \U$39348 ( \39601 , \39600 , \31153 );
nor \U$39349 ( \39602 , \39599 , \30657 );
nor \U$39350 ( \39603 , \39601 , \39602 );
and \U$39351 ( \39604 , \39598 , \39603 );
and \U$39352 ( \39605 , \39591 , \39597 );
or \U$39353 ( \39606 , \39604 , \39605 );
not \U$39354 ( \39607 , \39606 );
xor \U$39355 ( \39608 , \39565 , \39567 );
xor \U$39356 ( \39609 , \39608 , \39570 );
nand \U$39357 ( \39610 , \39607 , \39609 );
xor \U$39358 ( \39611 , \39538 , \39544 );
xor \U$39359 ( \39612 , \39611 , \39573 );
xor \U$39360 ( \39613 , \39610 , \39612 );
not \U$39361 ( \39614 , \39613 );
not \U$39362 ( \39615 , \39606 );
not \U$39363 ( \39616 , \39609 );
or \U$39364 ( \39617 , \39615 , \39616 );
or \U$39365 ( \39618 , \39609 , \39606 );
nand \U$39366 ( \39619 , \39617 , \39618 );
not \U$39367 ( \39620 , \39619 );
xor \U$39368 ( \39621 , \39557 , \39551 );
xnor \U$39369 ( \39622 , \39621 , \39562 );
or \U$39370 ( \39623 , \30630 , \30626 );
and \U$39371 ( \39624 , \39623 , \31155 );
and \U$39372 ( \39625 , \30626 , \30630 );
nor \U$39373 ( \39626 , \39624 , \39625 );
xor \U$39374 ( \39627 , \39622 , \39626 );
xor \U$39375 ( \39628 , \39591 , \39597 );
xor \U$39376 ( \39629 , \39628 , \39603 );
and \U$39377 ( \39630 , \39627 , \39629 );
and \U$39378 ( \39631 , \39622 , \39626 );
or \U$39379 ( \39632 , \39630 , \39631 );
not \U$39380 ( \39633 , \39632 );
or \U$39381 ( \39634 , \39620 , \39633 );
or \U$39382 ( \39635 , \39632 , \39619 );
nand \U$39383 ( \39636 , \39634 , \39635 );
buf \U$39384 ( \39637 , \39636 );
nand \U$39385 ( \39638 , \39585 , \39614 , \39637 );
not \U$39386 ( \39639 , \11048 );
not \U$39387 ( \39640 , \11054 );
and \U$39388 ( \39641 , \39639 , \39640 );
and \U$39389 ( \39642 , \11048 , \11054 );
nor \U$39390 ( \39643 , \39641 , \39642 );
xnor \U$39391 ( \39644 , \39643 , \10625 );
not \U$39392 ( \39645 , \39644 );
xor \U$39393 ( \39646 , \12337 , \12368 );
xor \U$39394 ( \39647 , \39646 , \12399 );
and \U$39395 ( \39648 , \12186 , \12151 );
not \U$39396 ( \39649 , \12186 );
and \U$39397 ( \39650 , \39649 , \12150 );
nor \U$39398 ( \39651 , \39648 , \39650 );
xor \U$39399 ( \39652 , \12120 , \39651 );
xor \U$39400 ( \39653 , \39647 , \39652 );
and \U$39401 ( \39654 , \12303 , \12261 );
not \U$39402 ( \39655 , \12303 );
and \U$39403 ( \39656 , \39655 , \12260 );
nor \U$39404 ( \39657 , \39654 , \39656 );
and \U$39405 ( \39658 , \39657 , \12225 );
not \U$39406 ( \39659 , \39657 );
and \U$39407 ( \39660 , \39659 , \12224 );
nor \U$39408 ( \39661 , \39658 , \39660 );
and \U$39409 ( \39662 , \39653 , \39661 );
and \U$39410 ( \39663 , \39647 , \39652 );
or \U$39411 ( \39664 , \39662 , \39663 );
xor \U$39412 ( \39665 , \12041 , \12052 );
xor \U$39413 ( \39666 , \39665 , \12063 );
xor \U$39414 ( \39667 , \39664 , \39666 );
not \U$39415 ( \39668 , \12487 );
not \U$39416 ( \39669 , \12478 );
not \U$39417 ( \39670 , \12492 );
or \U$39418 ( \39671 , \39669 , \39670 );
nand \U$39419 ( \39672 , \12495 , \12491 );
nand \U$39420 ( \39673 , \39671 , \39672 );
not \U$39421 ( \39674 , \39673 );
or \U$39422 ( \39675 , \39668 , \39674 );
or \U$39423 ( \39676 , \39673 , \12487 );
nand \U$39424 ( \39677 , \39675 , \39676 );
and \U$39425 ( \39678 , \39667 , \39677 );
and \U$39426 ( \39679 , \39664 , \39666 );
or \U$39427 ( \39680 , \39678 , \39679 );
and \U$39428 ( \39681 , \10916 , RIbe27c10_3);
and \U$39429 ( \39682 , \15228 , RIbe28e58_42);
nor \U$39430 ( \39683 , \39681 , \39682 );
and \U$39431 ( \39684 , \39683 , \16437 );
not \U$39432 ( \39685 , \39683 );
and \U$39433 ( \39686 , \39685 , \8077 );
nor \U$39434 ( \39687 , \39684 , \39686 );
nand \U$39435 ( \39688 , \13049 , RIbe27b98_2);
and \U$39436 ( \39689 , \39688 , \12195 );
not \U$39437 ( \39690 , \39688 );
and \U$39438 ( \39691 , \39690 , \17005 );
nor \U$39439 ( \39692 , \39689 , \39691 );
nand \U$39440 ( \39693 , \39687 , \39692 );
not \U$39441 ( \39694 , \12971 );
not \U$39442 ( \39695 , RIbe29920_65);
or \U$39443 ( \39696 , \39694 , \39695 );
not \U$39444 ( \39697 , \13024 );
or \U$39445 ( \39698 , \39697 , \2890 );
nand \U$39446 ( \39699 , \39696 , \39698 );
not \U$39447 ( \39700 , \39699 );
not \U$39448 ( \39701 , \9903 );
or \U$39449 ( \39702 , \39700 , \39701 );
or \U$39450 ( \39703 , \39699 , \10940 );
nand \U$39451 ( \39704 , \39702 , \39703 );
and \U$39452 ( \39705 , \39693 , \39704 );
nor \U$39453 ( \39706 , \39692 , \39687 );
nor \U$39454 ( \39707 , \39705 , \39706 );
not \U$39455 ( \39708 , \39707 );
not \U$39456 ( \39709 , \39708 );
not \U$39457 ( \39710 , RIbe28228_16);
not \U$39458 ( \39711 , \8231 );
or \U$39459 ( \39712 , \39710 , \39711 );
nand \U$39460 ( \39713 , \9939 , RIbe281b0_15);
nand \U$39461 ( \39714 , \39712 , \39713 );
and \U$39462 ( \39715 , \39714 , \5740 );
not \U$39463 ( \39716 , \39714 );
and \U$39464 ( \39717 , \39716 , \7501 );
nor \U$39465 ( \39718 , \39715 , \39717 );
not \U$39466 ( \39719 , RIbe296c8_60);
not \U$39467 ( \39720 , \7941 );
or \U$39468 ( \39721 , \39719 , \39720 );
nand \U$39469 ( \39722 , \7483 , RIbe29650_59);
nand \U$39470 ( \39723 , \39721 , \39722 );
and \U$39471 ( \39724 , \39723 , \8957 );
not \U$39472 ( \39725 , \39723 );
and \U$39473 ( \39726 , \39725 , \6582 );
nor \U$39474 ( \39727 , \39724 , \39726 );
and \U$39475 ( \39728 , \39718 , \39727 );
not \U$39476 ( \39729 , \13412 );
not \U$39477 ( \39730 , RIbe280c0_13);
not \U$39478 ( \39731 , \6536 );
or \U$39479 ( \39732 , \39730 , \39731 );
nand \U$39480 ( \39733 , \7076 , RIbe29830_63);
nand \U$39481 ( \39734 , \39732 , \39733 );
not \U$39482 ( \39735 , \39734 );
or \U$39483 ( \39736 , \39729 , \39735 );
or \U$39484 ( \39737 , \39734 , \9933 );
nand \U$39485 ( \39738 , \39736 , \39737 );
not \U$39486 ( \39739 , \39738 );
nor \U$39487 ( \39740 , \39728 , \39739 );
nor \U$39488 ( \39741 , \39718 , \39727 );
nor \U$39489 ( \39742 , \39740 , \39741 );
not \U$39490 ( \39743 , \39742 );
not \U$39491 ( \39744 , \39743 );
or \U$39492 ( \39745 , \39709 , \39744 );
not \U$39493 ( \39746 , \39742 );
not \U$39494 ( \39747 , \39707 );
or \U$39495 ( \39748 , \39746 , \39747 );
not \U$39496 ( \39749 , RIbe27d78_6);
not \U$39497 ( \39750 , \10949 );
or \U$39498 ( \39751 , \39749 , \39750 );
nand \U$39499 ( \39752 , \10952 , RIbe27d00_5);
nand \U$39500 ( \39753 , \39751 , \39752 );
not \U$39501 ( \39754 , \39753 );
not \U$39502 ( \39755 , \7989 );
and \U$39503 ( \39756 , \39754 , \39755 );
and \U$39504 ( \39757 , \39753 , \6949 );
nor \U$39505 ( \39758 , \39756 , \39757 );
not \U$39506 ( \39759 , \39758 );
not \U$39507 ( \39760 , RIbe29038_46);
not \U$39508 ( \39761 , \6561 );
or \U$39509 ( \39762 , \39760 , \39761 );
nand \U$39510 ( \39763 , \7958 , RIbe28fc0_45);
nand \U$39511 ( \39764 , \39762 , \39763 );
not \U$39512 ( \39765 , \39764 );
not \U$39513 ( \39766 , \6572 );
and \U$39514 ( \39767 , \39765 , \39766 );
and \U$39515 ( \39768 , \39764 , \6569 );
nor \U$39516 ( \39769 , \39767 , \39768 );
not \U$39517 ( \39770 , \39769 );
or \U$39518 ( \39771 , \39759 , \39770 );
not \U$39519 ( \39772 , \13168 );
not \U$39520 ( \39773 , RIbe290b0_47);
not \U$39521 ( \39774 , \7298 );
or \U$39522 ( \39775 , \39773 , \39774 );
nand \U$39523 ( \39776 , \10898 , RIbe29a88_68);
nand \U$39524 ( \39777 , \39775 , \39776 );
not \U$39525 ( \39778 , \39777 );
or \U$39526 ( \39779 , \39772 , \39778 );
or \U$39527 ( \39780 , \39777 , \6992 );
nand \U$39528 ( \39781 , \39779 , \39780 );
nand \U$39529 ( \39782 , \39771 , \39781 );
or \U$39530 ( \39783 , \39758 , \39769 );
nand \U$39531 ( \39784 , \39782 , \39783 );
nand \U$39532 ( \39785 , \39748 , \39784 );
nand \U$39533 ( \39786 , \39745 , \39785 );
not \U$39534 ( \39787 , \39786 );
not \U$39535 ( \39788 , \39787 );
nand \U$39536 ( \39789 , RIbe29380_53, RIbe2a208_84);
not \U$39537 ( \39790 , \39789 );
not \U$39538 ( \39791 , RIbe2a190_83);
not \U$39539 ( \39792 , \325 );
or \U$39540 ( \39793 , \39791 , \39792 );
nand \U$39541 ( \39794 , \330 , RIbe2a5c8_92);
nand \U$39542 ( \39795 , \39793 , \39794 );
not \U$39543 ( \39796 , \39795 );
not \U$39544 ( \39797 , \1379 );
and \U$39545 ( \39798 , \39796 , \39797 );
and \U$39546 ( \39799 , \39795 , \4172 );
nor \U$39547 ( \39800 , \39798 , \39799 );
not \U$39548 ( \39801 , \39800 );
or \U$39549 ( \39802 , \39790 , \39801 );
and \U$39550 ( \39803 , \1357 , RIbe2a550_91);
and \U$39551 ( \39804 , \263 , RIbe2a988_100);
nor \U$39552 ( \39805 , \39803 , \39804 );
and \U$39553 ( \39806 , \39805 , \6058 );
not \U$39554 ( \39807 , \39805 );
and \U$39555 ( \39808 , \39807 , \1363 );
nor \U$39556 ( \39809 , \39806 , \39808 );
nand \U$39557 ( \39810 , \39802 , \39809 );
or \U$39558 ( \39811 , \39800 , \39789 );
nand \U$39559 ( \39812 , \39810 , \39811 );
not \U$39560 ( \39813 , RIbe29c68_72);
not \U$39561 ( \39814 , \1143 );
or \U$39562 ( \39815 , \39813 , \39814 );
nand \U$39563 ( \39816 , \1147 , RIbe29bf0_71);
nand \U$39564 ( \39817 , \39815 , \39816 );
and \U$39565 ( \39818 , \39817 , \3993 );
not \U$39566 ( \39819 , \39817 );
and \U$39567 ( \39820 , \39819 , \1157 );
nor \U$39568 ( \39821 , \39818 , \39820 );
and \U$39569 ( \39822 , \1807 , RIbe29e48_76);
and \U$39570 ( \39823 , \1203 , RIbe29dd0_75);
nor \U$39571 ( \39824 , \39822 , \39823 );
and \U$39572 ( \39825 , \39824 , \1813 );
not \U$39573 ( \39826 , \39824 );
and \U$39574 ( \39827 , \39826 , \1011 );
nor \U$39575 ( \39828 , \39825 , \39827 );
or \U$39576 ( \39829 , \39821 , \39828 );
not \U$39577 ( \39830 , RIbe2a028_80);
not \U$39578 ( \39831 , \32589 );
or \U$39579 ( \39832 , \39830 , \39831 );
nand \U$39580 ( \39833 , \1179 , RIbe29fb0_79);
nand \U$39581 ( \39834 , \39832 , \39833 );
not \U$39582 ( \39835 , \39834 );
not \U$39583 ( \39836 , \564 );
and \U$39584 ( \39837 , \39835 , \39836 );
and \U$39585 ( \39838 , \39834 , \564 );
nor \U$39586 ( \39839 , \39837 , \39838 );
not \U$39587 ( \39840 , \39839 );
nand \U$39588 ( \39841 , \39829 , \39840 );
nand \U$39589 ( \39842 , \39821 , \39828 );
nand \U$39590 ( \39843 , \39841 , \39842 );
xor \U$39591 ( \39844 , \39812 , \39843 );
and \U$39592 ( \39845 , \283 , RIbe2a910_99);
and \U$39593 ( \39846 , \3897 , RIbe2b5b8_126);
nor \U$39594 ( \39847 , \39845 , \39846 );
and \U$39595 ( \39848 , \39847 , \300 );
not \U$39596 ( \39849 , \39847 );
and \U$39597 ( \39850 , \39849 , \293 );
nor \U$39598 ( \39851 , \39848 , \39850 );
not \U$39599 ( \39852 , \39851 );
not \U$39600 ( \39853 , RIbe2a2f8_86);
not \U$39601 ( \39854 , \1756 );
or \U$39602 ( \39855 , \39853 , \39854 );
nand \U$39603 ( \39856 , \552 , RIbe2acd0_107);
nand \U$39604 ( \39857 , \39855 , \39856 );
not \U$39605 ( \39858 , \39857 );
not \U$39606 ( \39859 , \424 );
and \U$39607 ( \39860 , \39858 , \39859 );
and \U$39608 ( \39861 , \39857 , \424 );
nor \U$39609 ( \39862 , \39860 , \39861 );
not \U$39610 ( \39863 , \39862 );
not \U$39611 ( \39864 , \39863 );
or \U$39612 ( \39865 , \39852 , \39864 );
or \U$39613 ( \39866 , \39863 , \39851 );
not \U$39614 ( \39867 , \1547 );
not \U$39615 ( \39868 , RIbe2a3e8_88);
not \U$39616 ( \39869 , \1223 );
or \U$39617 ( \39870 , \39868 , \39869 );
nand \U$39618 ( \39871 , \429 , RIbe2a370_87);
nand \U$39619 ( \39872 , \39870 , \39871 );
not \U$39620 ( \39873 , \39872 );
or \U$39621 ( \39874 , \39867 , \39873 );
or \U$39622 ( \39875 , \39872 , \312 );
nand \U$39623 ( \39876 , \39874 , \39875 );
nand \U$39624 ( \39877 , \39866 , \39876 );
nand \U$39625 ( \39878 , \39865 , \39877 );
and \U$39626 ( \39879 , \39844 , \39878 );
and \U$39627 ( \39880 , \39812 , \39843 );
or \U$39628 ( \39881 , \39879 , \39880 );
not \U$39629 ( \39882 , \39881 );
not \U$39630 ( \39883 , \39882 );
and \U$39631 ( \39884 , \39788 , \39883 );
and \U$39632 ( \39885 , \39787 , \39882 );
not \U$39633 ( \39886 , RIbe28b88_36);
not \U$39634 ( \39887 , \4804 );
or \U$39635 ( \39888 , \39886 , \39887 );
nand \U$39636 ( \39889 , \4600 , RIbe29290_51);
nand \U$39637 ( \39890 , \39888 , \39889 );
xor \U$39638 ( \39891 , \39890 , \4323 );
not \U$39639 ( \39892 , RIbe28a20_33);
not \U$39640 ( \39893 , \5727 );
or \U$39641 ( \39894 , \39892 , \39893 );
nand \U$39642 ( \39895 , \7056 , RIbe289a8_32);
nand \U$39643 ( \39896 , \39894 , \39895 );
not \U$39644 ( \39897 , \39896 );
not \U$39645 ( \39898 , \4946 );
and \U$39646 ( \39899 , \39897 , \39898 );
and \U$39647 ( \39900 , \39896 , \4592 );
nor \U$39648 ( \39901 , \39899 , \39900 );
and \U$39649 ( \39902 , \39891 , \39901 );
not \U$39650 ( \39903 , RIbe28930_31);
not \U$39651 ( \39904 , \5455 );
or \U$39652 ( \39905 , \39903 , \39904 );
nand \U$39653 ( \39906 , \8247 , RIbe29560_57);
nand \U$39654 ( \39907 , \39905 , \39906 );
and \U$39655 ( \39908 , \39907 , \5754 );
not \U$39656 ( \39909 , \39907 );
and \U$39657 ( \39910 , \39909 , \6117 );
nor \U$39658 ( \39911 , \39908 , \39910 );
nor \U$39659 ( \39912 , \39902 , \39911 );
nor \U$39660 ( \39913 , \39891 , \39901 );
nor \U$39661 ( \39914 , \39912 , \39913 );
not \U$39662 ( \39915 , RIbe28f48_44);
not \U$39663 ( \39916 , \1094 );
or \U$39664 ( \39917 , \39915 , \39916 );
nand \U$39665 ( \39918 , \4730 , RIbe28ed0_43);
nand \U$39666 ( \39919 , \39917 , \39918 );
and \U$39667 ( \39920 , \39919 , \1309 );
not \U$39668 ( \39921 , \39919 );
and \U$39669 ( \39922 , \39921 , \4251 );
nor \U$39670 ( \39923 , \39920 , \39922 );
not \U$39671 ( \39924 , \39923 );
and \U$39672 ( \39925 , \6380 , RIbe27fd0_11);
and \U$39673 ( \39926 , \20663 , RIbe27f58_10);
nor \U$39674 ( \39927 , \39925 , \39926 );
and \U$39675 ( \39928 , \39927 , \1448 );
not \U$39676 ( \39929 , \39927 );
and \U$39677 ( \39930 , \39929 , \1132 );
nor \U$39678 ( \39931 , \39928 , \39930 );
not \U$39679 ( \39932 , \39931 );
and \U$39680 ( \39933 , \39924 , \39932 );
and \U$39681 ( \39934 , \4295 , RIbe27e68_8);
and \U$39682 ( \39935 , \2384 , RIbe28660_25);
nor \U$39683 ( \39936 , \39934 , \39935 );
and \U$39684 ( \39937 , \39936 , \1274 );
not \U$39685 ( \39938 , \39936 );
and \U$39686 ( \39939 , \39938 , \1076 );
nor \U$39687 ( \39940 , \39937 , \39939 );
nor \U$39688 ( \39941 , \39933 , \39940 );
nor \U$39689 ( \39942 , \39924 , \39932 );
nor \U$39690 ( \39943 , \39941 , \39942 );
nand \U$39691 ( \39944 , \39914 , \39943 );
not \U$39692 ( \39945 , RIbe285e8_24);
not \U$39693 ( \39946 , \2898 );
or \U$39694 ( \39947 , \39945 , \39946 );
nand \U$39695 ( \39948 , \3267 , RIbe287c8_28);
nand \U$39696 ( \39949 , \39947 , \39948 );
and \U$39697 ( \39950 , \39949 , \2380 );
not \U$39698 ( \39951 , \39949 );
and \U$39699 ( \39952 , \39951 , \2379 );
nor \U$39700 ( \39953 , \39950 , \39952 );
not \U$39701 ( \39954 , RIbe28480_21);
not \U$39702 ( \39955 , \3284 );
or \U$39703 ( \39956 , \39954 , \39955 );
nand \U$39704 ( \39957 , \4011 , RIbe28408_20);
nand \U$39705 ( \39958 , \39956 , \39957 );
and \U$39706 ( \39959 , \39958 , \2887 );
not \U$39707 ( \39960 , \39958 );
and \U$39708 ( \39961 , \39960 , \3290 );
nor \U$39709 ( \39962 , \39959 , \39961 );
not \U$39710 ( \39963 , \39962 );
or \U$39711 ( \39964 , \39953 , \39963 );
not \U$39712 ( \39965 , RIbe28390_19);
not \U$39713 ( \39966 , \7880 );
or \U$39714 ( \39967 , \39965 , \39966 );
nand \U$39715 ( \39968 , \4332 , RIbe28b10_35);
nand \U$39716 ( \39969 , \39967 , \39968 );
and \U$39717 ( \39970 , \39969 , \3471 );
not \U$39718 ( \39971 , \39969 );
and \U$39719 ( \39972 , \39971 , \3448 );
nor \U$39720 ( \39973 , \39970 , \39972 );
nand \U$39721 ( \39974 , \39964 , \39973 );
nand \U$39722 ( \39975 , \39963 , \39953 );
nand \U$39723 ( \39976 , \39974 , \39975 );
and \U$39724 ( \39977 , \39944 , \39976 );
nor \U$39725 ( \39978 , \39914 , \39943 );
nor \U$39726 ( \39979 , \39977 , \39978 );
nor \U$39727 ( \39980 , \39885 , \39979 );
nor \U$39728 ( \39981 , \39884 , \39980 );
not \U$39729 ( \39982 , \39981 );
xor \U$39730 ( \39983 , \12131 , \12140 );
xor \U$39731 ( \39984 , \39983 , \12147 );
xor \U$39732 ( \39985 , \12172 , \12162 );
xor \U$39733 ( \39986 , \39985 , \12183 );
or \U$39734 ( \39987 , \39984 , \39986 );
not \U$39735 ( \39988 , \12117 );
not \U$39736 ( \39989 , \12098 );
or \U$39737 ( \39990 , \39988 , \39989 );
nand \U$39738 ( \39991 , \12116 , \12097 );
nand \U$39739 ( \39992 , \39990 , \39991 );
xnor \U$39740 ( \39993 , \39992 , \12107 );
and \U$39741 ( \39994 , \39987 , \39993 );
and \U$39742 ( \39995 , \39984 , \39986 );
nor \U$39743 ( \39996 , \39994 , \39995 );
not \U$39744 ( \39997 , \12366 );
not \U$39745 ( \39998 , \12345 );
or \U$39746 ( \39999 , \39997 , \39998 );
or \U$39747 ( \40000 , \12345 , \12366 );
nand \U$39748 ( \40001 , \39999 , \40000 );
xnor \U$39749 ( \40002 , \40001 , \12354 );
xor \U$39750 ( \40003 , \12309 , \12325 );
xnor \U$39751 ( \40004 , \40003 , \12334 );
nand \U$39752 ( \40005 , \40002 , \40004 );
xor \U$39753 ( \40006 , \12378 , \12388 );
xor \U$39754 ( \40007 , \40006 , \12396 );
and \U$39755 ( \40008 , \40005 , \40007 );
nor \U$39756 ( \40009 , \40004 , \40002 );
nor \U$39757 ( \40010 , \40008 , \40009 );
or \U$39758 ( \40011 , \39996 , \40010 );
not \U$39759 ( \40012 , \40010 );
not \U$39760 ( \40013 , \39996 );
or \U$39761 ( \40014 , \40012 , \40013 );
xor \U$39762 ( \40015 , \12195 , \12206 );
xor \U$39763 ( \40016 , \40015 , \12221 );
not \U$39764 ( \40017 , \40016 );
not \U$39765 ( \40018 , \40017 );
xor \U$39766 ( \40019 , \12257 , \12236 );
not \U$39767 ( \40020 , \12245 );
xor \U$39768 ( \40021 , \40019 , \40020 );
not \U$39769 ( \40022 , \40021 );
not \U$39770 ( \40023 , \40022 );
or \U$39771 ( \40024 , \40018 , \40023 );
not \U$39772 ( \40025 , \40021 );
not \U$39773 ( \40026 , \40016 );
or \U$39774 ( \40027 , \40025 , \40026 );
xor \U$39775 ( \40028 , \12277 , \12300 );
xor \U$39776 ( \40029 , \40028 , \12288 );
nand \U$39777 ( \40030 , \40027 , \40029 );
nand \U$39778 ( \40031 , \40024 , \40030 );
nand \U$39779 ( \40032 , \40014 , \40031 );
nand \U$39780 ( \40033 , \40011 , \40032 );
not \U$39781 ( \40034 , \40033 );
not \U$39782 ( \40035 , \40034 );
or \U$39783 ( \40036 , \39982 , \40035 );
xor \U$39784 ( \40037 , \12406 , \12408 );
xor \U$39785 ( \40038 , \40037 , \12420 );
not \U$39786 ( \40039 , \40038 );
not \U$39787 ( \40040 , \40039 );
not \U$39788 ( \40041 , \12429 );
not \U$39789 ( \40042 , \12448 );
or \U$39790 ( \40043 , \40041 , \40042 );
or \U$39791 ( \40044 , \12429 , \12448 );
nand \U$39792 ( \40045 , \40043 , \40044 );
and \U$39793 ( \40046 , \40045 , \12440 );
not \U$39794 ( \40047 , \40045 );
and \U$39795 ( \40048 , \40047 , \12451 );
nor \U$39796 ( \40049 , \40046 , \40048 );
not \U$39797 ( \40050 , \40049 );
or \U$39798 ( \40051 , \40040 , \40050 );
xor \U$39799 ( \40052 , \12461 , \12463 );
xor \U$39800 ( \40053 , \40052 , \12466 );
nand \U$39801 ( \40054 , \40051 , \40053 );
not \U$39802 ( \40055 , \40049 );
nand \U$39803 ( \40056 , \40055 , \40038 );
nand \U$39804 ( \40057 , \40054 , \40056 );
nand \U$39805 ( \40058 , \40036 , \40057 );
not \U$39806 ( \40059 , \39981 );
nand \U$39807 ( \40060 , \40059 , \40033 );
and \U$39808 ( \40061 , \40058 , \40060 );
xor \U$39809 ( \40062 , \12190 , \12305 );
xnor \U$39810 ( \40063 , \40062 , \12402 );
not \U$39811 ( \40064 , \40063 );
xor \U$39812 ( \40065 , \12423 , \12453 );
xor \U$39813 ( \40066 , \40065 , \12469 );
nand \U$39814 ( \40067 , \40064 , \40066 );
nand \U$39815 ( \40068 , \40061 , \40067 );
and \U$39816 ( \40069 , \39680 , \40068 );
nor \U$39817 ( \40070 , \40061 , \40067 );
nor \U$39818 ( \40071 , \40069 , \40070 );
not \U$39819 ( \40072 , \40071 );
not \U$39820 ( \40073 , \40072 );
not \U$39821 ( \40074 , \40073 );
xor \U$39822 ( \40075 , \12527 , \12522 );
xnor \U$39823 ( \40076 , \40075 , \12512 );
not \U$39824 ( \40077 , \40076 );
or \U$39825 ( \40078 , \40074 , \40077 );
not \U$39826 ( \40079 , \12088 );
not \U$39827 ( \40080 , \12080 );
or \U$39828 ( \40081 , \40079 , \40080 );
or \U$39829 ( \40082 , \12080 , \12088 );
nand \U$39830 ( \40083 , \40081 , \40082 );
xor \U$39831 ( \40084 , \12404 , \12472 );
xor \U$39832 ( \40085 , \40084 , \12497 );
xor \U$39833 ( \40086 , \40083 , \40085 );
not \U$39834 ( \40087 , \12038 );
xnor \U$39835 ( \40088 , \12066 , \12070 );
not \U$39836 ( \40089 , \40088 );
or \U$39837 ( \40090 , \40087 , \40089 );
or \U$39838 ( \40091 , \12038 , \40088 );
nand \U$39839 ( \40092 , \40090 , \40091 );
and \U$39840 ( \40093 , \40086 , \40092 );
and \U$39841 ( \40094 , \40083 , \40085 );
or \U$39842 ( \40095 , \40093 , \40094 );
nand \U$39843 ( \40096 , \40078 , \40095 );
not \U$39844 ( \40097 , \40073 );
not \U$39845 ( \40098 , \40076 );
nand \U$39846 ( \40099 , \40097 , \40098 );
nand \U$39847 ( \40100 , \40096 , \40099 );
not \U$39848 ( \40101 , \40100 );
or \U$39849 ( \40102 , \39645 , \40101 );
not \U$39850 ( \40103 , \39644 );
nand \U$39851 ( \40104 , \40103 , \40099 , \40096 );
nand \U$39852 ( \40105 , \40102 , \40104 );
nor \U$39853 ( \40106 , \12531 , \12505 );
not \U$39854 ( \40107 , \40106 );
nand \U$39855 ( \40108 , \12531 , \12505 );
nand \U$39856 ( \40109 , \40107 , \40108 );
not \U$39857 ( \40110 , \12536 );
and \U$39858 ( \40111 , \40109 , \40110 );
not \U$39859 ( \40112 , \40109 );
and \U$39860 ( \40113 , \40112 , \12536 );
nor \U$39861 ( \40114 , \40111 , \40113 );
not \U$39862 ( \40115 , \40114 );
and \U$39863 ( \40116 , \40105 , \40115 );
not \U$39864 ( \40117 , \40105 );
and \U$39865 ( \40118 , \40117 , \40114 );
nor \U$39866 ( \40119 , \40116 , \40118 );
not \U$39867 ( \40120 , \12073 );
not \U$39868 ( \40121 , \12089 );
not \U$39869 ( \40122 , \12500 );
or \U$39870 ( \40123 , \40121 , \40122 );
or \U$39871 ( \40124 , \12500 , \12089 );
nand \U$39872 ( \40125 , \40123 , \40124 );
not \U$39873 ( \40126 , \40125 );
or \U$39874 ( \40127 , \40120 , \40126 );
or \U$39875 ( \40128 , \40125 , \12073 );
nand \U$39876 ( \40129 , \40127 , \40128 );
not \U$39877 ( \40130 , \39996 );
not \U$39878 ( \40131 , \40031 );
or \U$39879 ( \40132 , \40130 , \40131 );
buf \U$39880 ( \40133 , \39996 );
or \U$39881 ( \40134 , \40133 , \40031 );
nand \U$39882 ( \40135 , \40132 , \40134 );
not \U$39883 ( \40136 , \40135 );
not \U$39884 ( \40137 , \40010 );
and \U$39885 ( \40138 , \40136 , \40137 );
and \U$39886 ( \40139 , \40010 , \40135 );
nor \U$39887 ( \40140 , \40138 , \40139 );
not \U$39888 ( \40141 , \40140 );
not \U$39889 ( \40142 , \39786 );
not \U$39890 ( \40143 , \39979 );
or \U$39891 ( \40144 , \40142 , \40143 );
or \U$39892 ( \40145 , \39786 , \39979 );
nand \U$39893 ( \40146 , \40144 , \40145 );
xor \U$39894 ( \40147 , \39881 , \40146 );
nand \U$39895 ( \40148 , \40141 , \40147 );
not \U$39896 ( \40149 , \40148 );
xor \U$39897 ( \40150 , \39984 , \39986 );
xor \U$39898 ( \40151 , \40150 , \39993 );
not \U$39899 ( \40152 , \40151 );
xor \U$39900 ( \40153 , \40004 , \40007 );
xor \U$39901 ( \40154 , \40153 , \40002 );
not \U$39902 ( \40155 , \40154 );
and \U$39903 ( \40156 , \40152 , \40155 );
not \U$39904 ( \40157 , \40021 );
not \U$39905 ( \40158 , \40017 );
or \U$39906 ( \40159 , \40157 , \40158 );
nand \U$39907 ( \40160 , \40022 , \40016 );
nand \U$39908 ( \40161 , \40159 , \40160 );
not \U$39909 ( \40162 , \40029 );
and \U$39910 ( \40163 , \40161 , \40162 );
not \U$39911 ( \40164 , \40161 );
and \U$39912 ( \40165 , \40164 , \40029 );
nor \U$39913 ( \40166 , \40163 , \40165 );
nor \U$39914 ( \40167 , \40156 , \40166 );
and \U$39915 ( \40168 , \40154 , \40151 );
nor \U$39916 ( \40169 , \40167 , \40168 );
not \U$39917 ( \40170 , \39123 );
not \U$39918 ( \40171 , \39099 );
or \U$39919 ( \40172 , \40170 , \40171 );
nand \U$39920 ( \40173 , \40172 , \39110 );
nand \U$39921 ( \40174 , \39098 , \39124 );
nand \U$39922 ( \40175 , \40173 , \40174 );
xor \U$39923 ( \40176 , \39070 , \39079 );
and \U$39924 ( \40177 , \40176 , \39087 );
and \U$39925 ( \40178 , \39070 , \39079 );
or \U$39926 ( \40179 , \40177 , \40178 );
xor \U$39927 ( \40180 , \40175 , \40179 );
not \U$39928 ( \40181 , \39223 );
not \U$39929 ( \40182 , \39209 );
or \U$39930 ( \40183 , \40181 , \40182 );
nand \U$39931 ( \40184 , \40183 , \39198 );
not \U$39932 ( \40185 , \39209 );
nand \U$39933 ( \40186 , \40185 , \39224 );
nand \U$39934 ( \40187 , \40184 , \40186 );
and \U$39935 ( \40188 , \40180 , \40187 );
and \U$39936 ( \40189 , \40175 , \40179 );
or \U$39937 ( \40190 , \40188 , \40189 );
not \U$39938 ( \40191 , \40190 );
nand \U$39939 ( \40192 , \39031 , \12927 );
and \U$39940 ( \40193 , \39020 , \12956 );
not \U$39941 ( \40194 , \39020 );
and \U$39942 ( \40195 , \40194 , \12195 );
nor \U$39943 ( \40196 , \40193 , \40195 );
and \U$39944 ( \40197 , \40192 , \40196 );
nor \U$39945 ( \40198 , \39030 , \12927 );
nor \U$39946 ( \40199 , \40197 , \40198 );
not \U$39947 ( \40200 , \40199 );
not \U$39948 ( \40201 , \40200 );
not \U$39949 ( \40202 , \39166 );
not \U$39950 ( \40203 , \39175 );
and \U$39951 ( \40204 , \40202 , \40203 );
nor \U$39952 ( \40205 , \40204 , \39186 );
and \U$39953 ( \40206 , \39166 , \39175 );
nor \U$39954 ( \40207 , \40205 , \40206 );
not \U$39955 ( \40208 , \40207 );
not \U$39956 ( \40209 , \40208 );
or \U$39957 ( \40210 , \40201 , \40209 );
not \U$39958 ( \40211 , \40199 );
not \U$39959 ( \40212 , \40207 );
or \U$39960 ( \40213 , \40211 , \40212 );
xor \U$39961 ( \40214 , \39139 , \39148 );
and \U$39962 ( \40215 , \40214 , \39158 );
and \U$39963 ( \40216 , \39139 , \39148 );
or \U$39964 ( \40217 , \40215 , \40216 );
nand \U$39965 ( \40218 , \40213 , \40217 );
nand \U$39966 ( \40219 , \40210 , \40218 );
not \U$39967 ( \40220 , \40219 );
and \U$39968 ( \40221 , \40191 , \40220 );
not \U$39969 ( \40222 , \39002 );
not \U$39970 ( \40223 , \39012 );
or \U$39971 ( \40224 , \40222 , \40223 );
nand \U$39972 ( \40225 , \39011 , \38999 );
nand \U$39973 ( \40226 , \40225 , \38992 );
nand \U$39974 ( \40227 , \40224 , \40226 );
and \U$39975 ( \40228 , \38983 , \38962 );
nor \U$39976 ( \40229 , \40228 , \38969 );
nor \U$39977 ( \40230 , \38983 , \38962 );
nor \U$39978 ( \40231 , \40229 , \40230 );
not \U$39979 ( \40232 , \40231 );
or \U$39980 ( \40233 , \40227 , \40232 );
xor \U$39981 ( \40234 , \39043 , \39050 );
and \U$39982 ( \40235 , \40234 , \39060 );
and \U$39983 ( \40236 , \39043 , \39050 );
or \U$39984 ( \40237 , \40235 , \40236 );
nand \U$39985 ( \40238 , \40233 , \40237 );
nand \U$39986 ( \40239 , \40227 , \40232 );
and \U$39987 ( \40240 , \40238 , \40239 );
nor \U$39988 ( \40241 , \40221 , \40240 );
and \U$39989 ( \40242 , \40219 , \40190 );
nor \U$39990 ( \40243 , \40241 , \40242 );
and \U$39991 ( \40244 , \40169 , \40243 );
xor \U$39992 ( \40245 , \39862 , \39876 );
xor \U$39993 ( \40246 , \40245 , \39851 );
xor \U$39994 ( \40247 , \39789 , \39800 );
xnor \U$39995 ( \40248 , \40247 , \39809 );
nand \U$39996 ( \40249 , \40246 , \40248 );
and \U$39997 ( \40250 , \39940 , \39931 );
not \U$39998 ( \40251 , \39940 );
and \U$39999 ( \40252 , \40251 , \39932 );
or \U$40000 ( \40253 , \40250 , \40252 );
and \U$40001 ( \40254 , \40253 , \39924 );
not \U$40002 ( \40255 , \40253 );
and \U$40003 ( \40256 , \40255 , \39923 );
nor \U$40004 ( \40257 , \40254 , \40256 );
not \U$40005 ( \40258 , \40257 );
not \U$40006 ( \40259 , \40258 );
xor \U$40007 ( \40260 , \39962 , \39973 );
xnor \U$40008 ( \40261 , \40260 , \39953 );
not \U$40009 ( \40262 , \40261 );
or \U$40010 ( \40263 , \40259 , \40262 );
not \U$40011 ( \40264 , \40261 );
not \U$40012 ( \40265 , \40264 );
not \U$40013 ( \40266 , \40257 );
or \U$40014 ( \40267 , \40265 , \40266 );
and \U$40015 ( \40268 , \39821 , \39839 );
not \U$40016 ( \40269 , \39821 );
and \U$40017 ( \40270 , \40269 , \39840 );
or \U$40018 ( \40271 , \40268 , \40270 );
xor \U$40019 ( \40272 , \40271 , \39828 );
nand \U$40020 ( \40273 , \40267 , \40272 );
nand \U$40021 ( \40274 , \40263 , \40273 );
xor \U$40022 ( \40275 , \40249 , \40274 );
not \U$40023 ( \40276 , \39718 );
not \U$40024 ( \40277 , \39738 );
not \U$40025 ( \40278 , \39727 );
or \U$40026 ( \40279 , \40277 , \40278 );
or \U$40027 ( \40280 , \39727 , \39738 );
nand \U$40028 ( \40281 , \40279 , \40280 );
not \U$40029 ( \40282 , \40281 );
or \U$40030 ( \40283 , \40276 , \40282 );
or \U$40031 ( \40284 , \40281 , \39718 );
nand \U$40032 ( \40285 , \40283 , \40284 );
xor \U$40033 ( \40286 , \39769 , \39781 );
xor \U$40034 ( \40287 , \40286 , \39758 );
xor \U$40035 ( \40288 , \40285 , \40287 );
xor \U$40036 ( \40289 , \39901 , \39911 );
not \U$40037 ( \40290 , \39891 );
xor \U$40038 ( \40291 , \40289 , \40290 );
and \U$40039 ( \40292 , \40288 , \40291 );
and \U$40040 ( \40293 , \40285 , \40287 );
or \U$40041 ( \40294 , \40292 , \40293 );
and \U$40042 ( \40295 , \40275 , \40294 );
and \U$40043 ( \40296 , \40249 , \40274 );
or \U$40044 ( \40297 , \40295 , \40296 );
not \U$40045 ( \40298 , \40297 );
nor \U$40046 ( \40299 , \40244 , \40298 );
nor \U$40047 ( \40300 , \40169 , \40243 );
nor \U$40048 ( \40301 , \40299 , \40300 );
not \U$40049 ( \40302 , \40301 );
or \U$40050 ( \40303 , \40149 , \40302 );
xor \U$40051 ( \40304 , \39812 , \39843 );
xor \U$40052 ( \40305 , \40304 , \39878 );
xor \U$40053 ( \40306 , \39707 , \39743 );
xnor \U$40054 ( \40307 , \40306 , \39784 );
xor \U$40055 ( \40308 , \40305 , \40307 );
xor \U$40056 ( \40309 , \39976 , \39914 );
xor \U$40057 ( \40310 , \40309 , \39943 );
and \U$40058 ( \40311 , \40308 , \40310 );
and \U$40059 ( \40312 , \40305 , \40307 );
or \U$40060 ( \40313 , \40311 , \40312 );
xor \U$40061 ( \40314 , \39647 , \39652 );
xor \U$40062 ( \40315 , \40314 , \39661 );
xor \U$40063 ( \40316 , \40313 , \40315 );
not \U$40064 ( \40317 , \40049 );
not \U$40065 ( \40318 , \40053 );
or \U$40066 ( \40319 , \40317 , \40318 );
not \U$40067 ( \40320 , \40053 );
nand \U$40068 ( \40321 , \40320 , \40055 );
nand \U$40069 ( \40322 , \40319 , \40321 );
and \U$40070 ( \40323 , \40322 , \40038 );
not \U$40071 ( \40324 , \40322 );
and \U$40072 ( \40325 , \40324 , \40039 );
nor \U$40073 ( \40326 , \40323 , \40325 );
and \U$40074 ( \40327 , \40316 , \40326 );
and \U$40075 ( \40328 , \40313 , \40315 );
or \U$40076 ( \40329 , \40327 , \40328 );
nand \U$40077 ( \40330 , \40303 , \40329 );
not \U$40078 ( \40331 , \40301 );
not \U$40079 ( \40332 , \40148 );
nand \U$40080 ( \40333 , \40331 , \40332 );
nand \U$40081 ( \40334 , \40330 , \40333 );
not \U$40082 ( \40335 , \40063 );
not \U$40083 ( \40336 , \40066 );
or \U$40084 ( \40337 , \40335 , \40336 );
or \U$40085 ( \40338 , \40066 , \40063 );
nand \U$40086 ( \40339 , \40337 , \40338 );
not \U$40087 ( \40340 , \40057 );
not \U$40088 ( \40341 , \40340 );
not \U$40089 ( \40342 , \39981 );
not \U$40090 ( \40343 , \40033 );
or \U$40091 ( \40344 , \40342 , \40343 );
or \U$40092 ( \40345 , \40033 , \39981 );
nand \U$40093 ( \40346 , \40344 , \40345 );
not \U$40094 ( \40347 , \40346 );
or \U$40095 ( \40348 , \40341 , \40347 );
or \U$40096 ( \40349 , \40346 , \40340 );
nand \U$40097 ( \40350 , \40348 , \40349 );
xor \U$40098 ( \40351 , \40339 , \40350 );
xor \U$40099 ( \40352 , \39664 , \39666 );
xor \U$40100 ( \40353 , \40352 , \39677 );
and \U$40101 ( \40354 , \40351 , \40353 );
and \U$40102 ( \40355 , \40339 , \40350 );
or \U$40103 ( \40356 , \40354 , \40355 );
xor \U$40104 ( \40357 , \40334 , \40356 );
xor \U$40105 ( \40358 , \40083 , \40085 );
xor \U$40106 ( \40359 , \40358 , \40092 );
and \U$40107 ( \40360 , \40357 , \40359 );
and \U$40108 ( \40361 , \40334 , \40356 );
or \U$40109 ( \40362 , \40360 , \40361 );
xor \U$40110 ( \40363 , \40129 , \40362 );
and \U$40111 ( \40364 , \40095 , \40072 );
not \U$40112 ( \40365 , \40095 );
and \U$40113 ( \40366 , \40365 , \40071 );
nor \U$40114 ( \40367 , \40364 , \40366 );
and \U$40115 ( \40368 , \40367 , \40098 );
not \U$40116 ( \40369 , \40367 );
and \U$40117 ( \40370 , \40369 , \40076 );
nor \U$40118 ( \40371 , \40368 , \40370 );
and \U$40119 ( \40372 , \40363 , \40371 );
and \U$40120 ( \40373 , \40129 , \40362 );
or \U$40121 ( \40374 , \40372 , \40373 );
buf \U$40122 ( \40375 , \40374 );
nand \U$40123 ( \40376 , \40119 , \40375 );
not \U$40124 ( \40377 , \40376 );
not \U$40125 ( \40378 , \40377 );
nand \U$40126 ( \40379 , \40114 , \39644 );
buf \U$40127 ( \40380 , \40100 );
and \U$40128 ( \40381 , \40379 , \40380 );
nor \U$40129 ( \40382 , \40114 , \39644 );
nor \U$40130 ( \40383 , \40381 , \40382 );
not \U$40131 ( \40384 , \40383 );
xor \U$40132 ( \40385 , \12036 , \12539 );
xor \U$40133 ( \40386 , \40385 , \12545 );
not \U$40134 ( \40387 , \40386 );
or \U$40135 ( \40388 , \40384 , \40387 );
or \U$40136 ( \40389 , \40383 , \40386 );
nand \U$40137 ( \40390 , \40388 , \40389 );
not \U$40138 ( \40391 , \40390 );
not \U$40139 ( \40392 , \40391 );
or \U$40140 ( \40393 , \40378 , \40392 );
nand \U$40141 ( \40394 , \40390 , \40376 );
nand \U$40142 ( \40395 , \40393 , \40394 );
xor \U$40143 ( \40396 , \39680 , \40061 );
xor \U$40144 ( \40397 , \40396 , \40067 );
not \U$40145 ( \40398 , \40240 );
xor \U$40146 ( \40399 , \40219 , \40190 );
not \U$40147 ( \40400 , \40399 );
or \U$40148 ( \40401 , \40398 , \40400 );
or \U$40149 ( \40402 , \40399 , \40240 );
nand \U$40150 ( \40403 , \40401 , \40402 );
xor \U$40151 ( \40404 , \40249 , \40274 );
xor \U$40152 ( \40405 , \40404 , \40294 );
and \U$40153 ( \40406 , \40403 , \40405 );
xor \U$40154 ( \40407 , \38919 , \38923 );
and \U$40155 ( \40408 , \40407 , \38930 );
and \U$40156 ( \40409 , \38919 , \38923 );
or \U$40157 ( \40410 , \40408 , \40409 );
xor \U$40158 ( \40411 , \38937 , \38941 );
and \U$40159 ( \40412 , \40411 , \38949 );
and \U$40160 ( \40413 , \38937 , \38941 );
or \U$40161 ( \40414 , \40412 , \40413 );
xor \U$40162 ( \40415 , \40410 , \40414 );
not \U$40163 ( \40416 , \38859 );
not \U$40164 ( \40417 , \38852 );
or \U$40165 ( \40418 , \40416 , \40417 );
or \U$40166 ( \40419 , \38852 , \38859 );
nand \U$40167 ( \40420 , \40419 , \38866 );
nand \U$40168 ( \40421 , \40418 , \40420 );
and \U$40169 ( \40422 , \40415 , \40421 );
and \U$40170 ( \40423 , \40410 , \40414 );
or \U$40171 ( \40424 , \40422 , \40423 );
xor \U$40172 ( \40425 , \38952 , \38984 );
and \U$40173 ( \40426 , \40425 , \39013 );
and \U$40174 ( \40427 , \38952 , \38984 );
or \U$40175 ( \40428 , \40426 , \40427 );
xor \U$40176 ( \40429 , \39061 , \39088 );
and \U$40177 ( \40430 , \40429 , \39128 );
and \U$40178 ( \40431 , \39061 , \39088 );
or \U$40179 ( \40432 , \40430 , \40431 );
xor \U$40180 ( \40433 , \40428 , \40432 );
xor \U$40181 ( \40434 , \39159 , \39187 );
and \U$40182 ( \40435 , \40434 , \39228 );
and \U$40183 ( \40436 , \39159 , \39187 );
or \U$40184 ( \40437 , \40435 , \40436 );
and \U$40185 ( \40438 , \40433 , \40437 );
and \U$40186 ( \40439 , \40428 , \40432 );
or \U$40187 ( \40440 , \40438 , \40439 );
xor \U$40188 ( \40441 , \40424 , \40440 );
buf \U$40189 ( \40442 , \39687 );
not \U$40190 ( \40443 , \40442 );
not \U$40191 ( \40444 , \39692 );
not \U$40192 ( \40445 , \39704 );
or \U$40193 ( \40446 , \40444 , \40445 );
or \U$40194 ( \40447 , \39704 , \39692 );
nand \U$40195 ( \40448 , \40446 , \40447 );
not \U$40196 ( \40449 , \40448 );
or \U$40197 ( \40450 , \40443 , \40449 );
or \U$40198 ( \40451 , \40448 , \40442 );
nand \U$40199 ( \40452 , \40450 , \40451 );
not \U$40200 ( \40453 , \40258 );
not \U$40201 ( \40454 , \40264 );
or \U$40202 ( \40455 , \40453 , \40454 );
nand \U$40203 ( \40456 , \40261 , \40257 );
nand \U$40204 ( \40457 , \40455 , \40456 );
and \U$40205 ( \40458 , \40457 , \40272 );
not \U$40206 ( \40459 , \40457 );
not \U$40207 ( \40460 , \40272 );
and \U$40208 ( \40461 , \40459 , \40460 );
nor \U$40209 ( \40462 , \40458 , \40461 );
xor \U$40210 ( \40463 , \40452 , \40462 );
xor \U$40211 ( \40464 , \40285 , \40287 );
xor \U$40212 ( \40465 , \40464 , \40291 );
and \U$40213 ( \40466 , \40463 , \40465 );
and \U$40214 ( \40467 , \40452 , \40462 );
or \U$40215 ( \40468 , \40466 , \40467 );
and \U$40216 ( \40469 , \40441 , \40468 );
and \U$40217 ( \40470 , \40424 , \40440 );
or \U$40218 ( \40471 , \40469 , \40470 );
xor \U$40219 ( \40472 , \40406 , \40471 );
or \U$40220 ( \40473 , \40248 , \40246 );
nand \U$40221 ( \40474 , \40473 , \40249 );
xor \U$40222 ( \40475 , \40175 , \40179 );
xor \U$40223 ( \40476 , \40475 , \40187 );
xor \U$40224 ( \40477 , \40474 , \40476 );
xor \U$40225 ( \40478 , \40227 , \40237 );
xnor \U$40226 ( \40479 , \40478 , \40231 );
and \U$40227 ( \40480 , \40477 , \40479 );
and \U$40228 ( \40481 , \40474 , \40476 );
or \U$40229 ( \40482 , \40480 , \40481 );
xor \U$40230 ( \40483 , \40305 , \40307 );
xor \U$40231 ( \40484 , \40483 , \40310 );
xor \U$40232 ( \40485 , \40482 , \40484 );
not \U$40233 ( \40486 , \40166 );
xor \U$40234 ( \40487 , \40154 , \40151 );
not \U$40235 ( \40488 , \40487 );
or \U$40236 ( \40489 , \40486 , \40488 );
or \U$40237 ( \40490 , \40487 , \40166 );
nand \U$40238 ( \40491 , \40489 , \40490 );
and \U$40239 ( \40492 , \40485 , \40491 );
and \U$40240 ( \40493 , \40482 , \40484 );
or \U$40241 ( \40494 , \40492 , \40493 );
and \U$40242 ( \40495 , \40472 , \40494 );
and \U$40243 ( \40496 , \40406 , \40471 );
or \U$40244 ( \40497 , \40495 , \40496 );
not \U$40245 ( \40498 , \40147 );
not \U$40246 ( \40499 , \40140 );
or \U$40247 ( \40500 , \40498 , \40499 );
or \U$40248 ( \40501 , \40140 , \40147 );
nand \U$40249 ( \40502 , \40500 , \40501 );
buf \U$40250 ( \40503 , \40169 );
not \U$40251 ( \40504 , \40503 );
not \U$40252 ( \40505 , \40243 );
not \U$40253 ( \40506 , \40297 );
or \U$40254 ( \40507 , \40505 , \40506 );
or \U$40255 ( \40508 , \40243 , \40297 );
nand \U$40256 ( \40509 , \40507 , \40508 );
not \U$40257 ( \40510 , \40509 );
or \U$40258 ( \40511 , \40504 , \40510 );
or \U$40259 ( \40512 , \40503 , \40509 );
nand \U$40260 ( \40513 , \40511 , \40512 );
xor \U$40261 ( \40514 , \40502 , \40513 );
xor \U$40262 ( \40515 , \40313 , \40315 );
xor \U$40263 ( \40516 , \40515 , \40326 );
and \U$40264 ( \40517 , \40514 , \40516 );
and \U$40265 ( \40518 , \40502 , \40513 );
or \U$40266 ( \40519 , \40517 , \40518 );
xor \U$40267 ( \40520 , \40497 , \40519 );
xor \U$40268 ( \40521 , \40339 , \40350 );
xor \U$40269 ( \40522 , \40521 , \40353 );
and \U$40270 ( \40523 , \40520 , \40522 );
and \U$40271 ( \40524 , \40497 , \40519 );
or \U$40272 ( \40525 , \40523 , \40524 );
xor \U$40273 ( \40526 , \40397 , \40525 );
xor \U$40274 ( \40527 , \40334 , \40356 );
xor \U$40275 ( \40528 , \40527 , \40359 );
and \U$40276 ( \40529 , \40526 , \40528 );
and \U$40277 ( \40530 , \40397 , \40525 );
or \U$40278 ( \40531 , \40529 , \40530 );
xor \U$40279 ( \40532 , \40129 , \40362 );
xor \U$40280 ( \40533 , \40532 , \40371 );
nand \U$40281 ( \40534 , \40531 , \40533 );
not \U$40282 ( \40535 , \40534 );
not \U$40283 ( \40536 , \40375 );
not \U$40284 ( \40537 , \40119 );
not \U$40285 ( \40538 , \40537 );
or \U$40286 ( \40539 , \40536 , \40538 );
not \U$40287 ( \40540 , \40374 );
nand \U$40288 ( \40541 , \40540 , \40119 );
nand \U$40289 ( \40542 , \40539 , \40541 );
not \U$40290 ( \40543 , \40542 );
or \U$40291 ( \40544 , \40535 , \40543 );
or \U$40292 ( \40545 , \40534 , \40542 );
nand \U$40293 ( \40546 , \40544 , \40545 );
nand \U$40294 ( \40547 , \40395 , \40546 );
and \U$40295 ( \40548 , \40301 , \40148 );
not \U$40296 ( \40549 , \40301 );
and \U$40297 ( \40550 , \40549 , \40332 );
nor \U$40298 ( \40551 , \40548 , \40550 );
xor \U$40299 ( \40552 , \40329 , \40551 );
not \U$40300 ( \40553 , \38841 );
not \U$40301 ( \40554 , \38832 );
or \U$40302 ( \40555 , \40553 , \40554 );
or \U$40303 ( \40556 , \38841 , \38832 );
nand \U$40304 ( \40557 , \40556 , \38828 );
nand \U$40305 ( \40558 , \40555 , \40557 );
xor \U$40306 ( \40559 , \38895 , \38904 );
and \U$40307 ( \40560 , \40559 , \38912 );
and \U$40308 ( \40561 , \38895 , \38904 );
or \U$40309 ( \40562 , \40560 , \40561 );
xor \U$40310 ( \40563 , \40558 , \40562 );
xor \U$40311 ( \40564 , \39032 , \39129 );
and \U$40312 ( \40565 , \40564 , \39229 );
and \U$40313 ( \40566 , \39032 , \39129 );
or \U$40314 ( \40567 , \40565 , \40566 );
and \U$40315 ( \40568 , \40563 , \40567 );
and \U$40316 ( \40569 , \40558 , \40562 );
or \U$40317 ( \40570 , \40568 , \40569 );
and \U$40318 ( \40571 , \40199 , \40207 );
not \U$40319 ( \40572 , \40199 );
and \U$40320 ( \40573 , \40572 , \40208 );
nor \U$40321 ( \40574 , \40571 , \40573 );
xor \U$40322 ( \40575 , \40574 , \40217 );
xor \U$40323 ( \40576 , \38931 , \38950 );
and \U$40324 ( \40577 , \40576 , \39014 );
and \U$40325 ( \40578 , \38931 , \38950 );
or \U$40326 ( \40579 , \40577 , \40578 );
xor \U$40327 ( \40580 , \40575 , \40579 );
xor \U$40328 ( \40581 , \40474 , \40476 );
xor \U$40329 ( \40582 , \40581 , \40479 );
and \U$40330 ( \40583 , \40580 , \40582 );
and \U$40331 ( \40584 , \40575 , \40579 );
or \U$40332 ( \40585 , \40583 , \40584 );
xor \U$40333 ( \40586 , \40570 , \40585 );
xor \U$40334 ( \40587 , \40410 , \40414 );
xor \U$40335 ( \40588 , \40587 , \40421 );
xor \U$40336 ( \40589 , \40428 , \40432 );
xor \U$40337 ( \40590 , \40589 , \40437 );
xor \U$40338 ( \40591 , \40588 , \40590 );
xor \U$40339 ( \40592 , \40452 , \40462 );
xor \U$40340 ( \40593 , \40592 , \40465 );
and \U$40341 ( \40594 , \40591 , \40593 );
and \U$40342 ( \40595 , \40588 , \40590 );
or \U$40343 ( \40596 , \40594 , \40595 );
and \U$40344 ( \40597 , \40586 , \40596 );
and \U$40345 ( \40598 , \40570 , \40585 );
or \U$40346 ( \40599 , \40597 , \40598 );
xor \U$40347 ( \40600 , \40403 , \40405 );
xor \U$40348 ( \40601 , \40424 , \40440 );
xor \U$40349 ( \40602 , \40601 , \40468 );
xor \U$40350 ( \40603 , \40600 , \40602 );
xor \U$40351 ( \40604 , \40482 , \40484 );
xor \U$40352 ( \40605 , \40604 , \40491 );
and \U$40353 ( \40606 , \40603 , \40605 );
and \U$40354 ( \40607 , \40600 , \40602 );
or \U$40355 ( \40608 , \40606 , \40607 );
xor \U$40356 ( \40609 , \40599 , \40608 );
xor \U$40357 ( \40610 , \40502 , \40513 );
xor \U$40358 ( \40611 , \40610 , \40516 );
and \U$40359 ( \40612 , \40609 , \40611 );
and \U$40360 ( \40613 , \40599 , \40608 );
or \U$40361 ( \40614 , \40612 , \40613 );
xor \U$40362 ( \40615 , \40552 , \40614 );
xor \U$40363 ( \40616 , \40497 , \40519 );
xor \U$40364 ( \40617 , \40616 , \40522 );
and \U$40365 ( \40618 , \40615 , \40617 );
and \U$40366 ( \40619 , \40552 , \40614 );
or \U$40367 ( \40620 , \40618 , \40619 );
xor \U$40368 ( \40621 , \40397 , \40525 );
xor \U$40369 ( \40622 , \40621 , \40528 );
and \U$40370 ( \40623 , \40620 , \40622 );
xor \U$40371 ( \40624 , \40531 , \40533 );
xor \U$40372 ( \40625 , \40623 , \40624 );
xor \U$40373 ( \40626 , \40620 , \40622 );
xor \U$40374 ( \40627 , \40406 , \40471 );
xor \U$40375 ( \40628 , \40627 , \40494 );
xor \U$40376 ( \40629 , \39265 , \39273 );
and \U$40377 ( \40630 , \40629 , \39278 );
and \U$40378 ( \40631 , \39265 , \39273 );
or \U$40379 ( \40632 , \40630 , \40631 );
not \U$40380 ( \40633 , \40632 );
not \U$40381 ( \40634 , \40633 );
and \U$40382 ( \40635 , \38847 , \38871 );
nor \U$40383 ( \40636 , \40635 , \38877 );
nor \U$40384 ( \40637 , \38847 , \38871 );
nor \U$40385 ( \40638 , \40636 , \40637 );
not \U$40386 ( \40639 , \40638 );
or \U$40387 ( \40640 , \40634 , \40639 );
xor \U$40388 ( \40641 , \38913 , \39015 );
and \U$40389 ( \40642 , \40641 , \39230 );
and \U$40390 ( \40643 , \38913 , \39015 );
or \U$40391 ( \40644 , \40642 , \40643 );
nand \U$40392 ( \40645 , \40640 , \40644 );
not \U$40393 ( \40646 , \40638 );
nand \U$40394 ( \40647 , \40646 , \40632 );
nand \U$40395 ( \40648 , \40645 , \40647 );
xor \U$40396 ( \40649 , \40558 , \40562 );
xor \U$40397 ( \40650 , \40649 , \40567 );
xor \U$40398 ( \40651 , \40575 , \40579 );
xor \U$40399 ( \40652 , \40651 , \40582 );
xor \U$40400 ( \40653 , \40650 , \40652 );
xor \U$40401 ( \40654 , \40588 , \40590 );
xor \U$40402 ( \40655 , \40654 , \40593 );
and \U$40403 ( \40656 , \40653 , \40655 );
and \U$40404 ( \40657 , \40650 , \40652 );
or \U$40405 ( \40658 , \40656 , \40657 );
xor \U$40406 ( \40659 , \40648 , \40658 );
xor \U$40407 ( \40660 , \40600 , \40602 );
xor \U$40408 ( \40661 , \40660 , \40605 );
and \U$40409 ( \40662 , \40659 , \40661 );
and \U$40410 ( \40663 , \40648 , \40658 );
or \U$40411 ( \40664 , \40662 , \40663 );
xor \U$40412 ( \40665 , \40628 , \40664 );
xor \U$40413 ( \40666 , \40599 , \40608 );
xor \U$40414 ( \40667 , \40666 , \40611 );
and \U$40415 ( \40668 , \40665 , \40667 );
and \U$40416 ( \40669 , \40628 , \40664 );
or \U$40417 ( \40670 , \40668 , \40669 );
xor \U$40418 ( \40671 , \40552 , \40614 );
xor \U$40419 ( \40672 , \40671 , \40617 );
and \U$40420 ( \40673 , \40670 , \40672 );
xor \U$40421 ( \40674 , \40626 , \40673 );
nand \U$40422 ( \40675 , \40625 , \40674 );
nor \U$40423 ( \40676 , \40547 , \40675 );
xor \U$40424 ( \40677 , \40670 , \40672 );
xor \U$40425 ( \40678 , \40570 , \40585 );
xor \U$40426 ( \40679 , \40678 , \40596 );
xor \U$40427 ( \40680 , \39236 , \39244 );
and \U$40428 ( \40681 , \40680 , \39249 );
and \U$40429 ( \40682 , \39236 , \39244 );
or \U$40430 ( \40683 , \40681 , \40682 );
xor \U$40431 ( \40684 , \38842 , \38888 );
and \U$40432 ( \40685 , \40684 , \39231 );
and \U$40433 ( \40686 , \38842 , \38888 );
or \U$40434 ( \40687 , \40685 , \40686 );
xor \U$40435 ( \40688 , \40683 , \40687 );
xor \U$40436 ( \40689 , \40650 , \40652 );
xor \U$40437 ( \40690 , \40689 , \40655 );
and \U$40438 ( \40691 , \40688 , \40690 );
and \U$40439 ( \40692 , \40683 , \40687 );
or \U$40440 ( \40693 , \40691 , \40692 );
xor \U$40441 ( \40694 , \40679 , \40693 );
xor \U$40442 ( \40695 , \40648 , \40658 );
xor \U$40443 ( \40696 , \40695 , \40661 );
and \U$40444 ( \40697 , \40694 , \40696 );
and \U$40445 ( \40698 , \40679 , \40693 );
or \U$40446 ( \40699 , \40697 , \40698 );
xor \U$40447 ( \40700 , \40628 , \40664 );
xor \U$40448 ( \40701 , \40700 , \40667 );
and \U$40449 ( \40702 , \40699 , \40701 );
xor \U$40450 ( \40703 , \40677 , \40702 );
not \U$40451 ( \40704 , \40703 );
nor \U$40452 ( \40705 , \12548 , \12029 );
not \U$40453 ( \40706 , \40705 );
nand \U$40454 ( \40707 , \12548 , \12029 );
nand \U$40455 ( \40708 , \40706 , \40707 );
not \U$40456 ( \40709 , \40708 );
not \U$40457 ( \40710 , \40383 );
nand \U$40458 ( \40711 , \40710 , \40386 );
not \U$40459 ( \40712 , \40711 );
and \U$40460 ( \40713 , \40709 , \40712 );
and \U$40461 ( \40714 , \40708 , \40711 );
nor \U$40462 ( \40715 , \40713 , \40714 );
nor \U$40463 ( \40716 , \40704 , \40715 );
nand \U$40464 ( \40717 , \40676 , \40716 );
xor \U$40465 ( \40718 , \39519 , \39521 );
and \U$40466 ( \40719 , \40718 , \39529 );
and \U$40467 ( \40720 , \39519 , \39521 );
or \U$40468 ( \40721 , \40719 , \40720 );
xor \U$40469 ( \40722 , \38799 , \38784 );
xor \U$40470 ( \40723 , \38797 , \40722 );
xor \U$40471 ( \40724 , \40721 , \40723 );
not \U$40472 ( \40725 , \39279 );
not \U$40473 ( \40726 , \40725 );
not \U$40474 ( \40727 , \39292 );
or \U$40475 ( \40728 , \40726 , \40727 );
not \U$40476 ( \40729 , \39286 );
nand \U$40477 ( \40730 , \40728 , \40729 );
not \U$40478 ( \40731 , \39292 );
nand \U$40479 ( \40732 , \40731 , \39279 );
nand \U$40480 ( \40733 , \40730 , \40732 );
nand \U$40481 ( \40734 , \39232 , \39250 );
xor \U$40482 ( \40735 , \40632 , \40646 );
xnor \U$40483 ( \40736 , \40735 , \40644 );
nand \U$40484 ( \40737 , \40734 , \40736 );
and \U$40485 ( \40738 , \40733 , \40737 );
nor \U$40486 ( \40739 , \40734 , \40736 );
nor \U$40487 ( \40740 , \40738 , \40739 );
not \U$40488 ( \40741 , \40740 );
xor \U$40489 ( \40742 , \40679 , \40693 );
xor \U$40490 ( \40743 , \40742 , \40696 );
nand \U$40491 ( \40744 , \40741 , \40743 );
not \U$40492 ( \40745 , \40744 );
not \U$40493 ( \40746 , \40745 );
xor \U$40494 ( \40747 , \40699 , \40701 );
not \U$40495 ( \40748 , \40747 );
not \U$40496 ( \40749 , \40748 );
or \U$40497 ( \40750 , \40746 , \40749 );
nand \U$40498 ( \40751 , \40747 , \40744 );
nand \U$40499 ( \40752 , \40750 , \40751 );
and \U$40500 ( \40753 , \40724 , \40752 );
nor \U$40501 ( \40754 , \38813 , \39298 );
xor \U$40502 ( \40755 , \40683 , \40687 );
xor \U$40503 ( \40756 , \40755 , \40690 );
and \U$40504 ( \40757 , \39293 , \39255 );
or \U$40505 ( \40758 , \40757 , \38821 );
nand \U$40506 ( \40759 , \39296 , \39256 );
nand \U$40507 ( \40760 , \40758 , \40759 );
xor \U$40508 ( \40761 , \40756 , \40760 );
xor \U$40509 ( \40762 , \40736 , \40734 );
xor \U$40510 ( \40763 , \40762 , \40733 );
xor \U$40511 ( \40764 , \40761 , \40763 );
xor \U$40512 ( \40765 , \40754 , \40764 );
xor \U$40513 ( \40766 , \40756 , \40760 );
and \U$40514 ( \40767 , \40766 , \40763 );
and \U$40515 ( \40768 , \40756 , \40760 );
or \U$40516 ( \40769 , \40767 , \40768 );
not \U$40517 ( \40770 , \40769 );
not \U$40518 ( \40771 , \40740 );
not \U$40519 ( \40772 , \40743 );
or \U$40520 ( \40773 , \40771 , \40772 );
or \U$40521 ( \40774 , \40740 , \40743 );
nand \U$40522 ( \40775 , \40773 , \40774 );
not \U$40523 ( \40776 , \40775 );
not \U$40524 ( \40777 , \40776 );
or \U$40525 ( \40778 , \40770 , \40777 );
not \U$40526 ( \40779 , \40769 );
nand \U$40527 ( \40780 , \40779 , \40775 );
nand \U$40528 ( \40781 , \40778 , \40780 );
nand \U$40529 ( \40782 , \40765 , \40781 );
not \U$40530 ( \40783 , \40782 );
nand \U$40531 ( \40784 , \30573 , \31160 );
xor \U$40532 ( \40785 , \39622 , \39626 );
xor \U$40533 ( \40786 , \40785 , \39629 );
xor \U$40534 ( \40787 , \40784 , \40786 );
nand \U$40535 ( \40788 , \40753 , \40783 , \40787 );
nor \U$40536 ( \40789 , \39313 , \39638 , \40717 , \40788 );
not \U$40537 ( \40790 , \40789 );
or \U$40538 ( \40791 , \32122 , \40790 );
not \U$40539 ( \40792 , \40717 );
nor \U$40540 ( \40793 , \39584 , \39613 );
not \U$40541 ( \40794 , \40793 );
not \U$40542 ( \40795 , \39636 );
nor \U$40543 ( \40796 , \40786 , \40784 );
not \U$40544 ( \40797 , \40796 );
or \U$40545 ( \40798 , \40795 , \40797 );
not \U$40546 ( \40799 , \39632 );
nand \U$40547 ( \40800 , \40799 , \39619 );
nand \U$40548 ( \40801 , \40798 , \40800 );
not \U$40549 ( \40802 , \40801 );
or \U$40550 ( \40803 , \40794 , \40802 );
not \U$40551 ( \40804 , \39612 );
nor \U$40552 ( \40805 , \40804 , \39610 );
and \U$40553 ( \40806 , \39585 , \40805 );
not \U$40554 ( \40807 , \39536 );
not \U$40555 ( \40808 , \39579 );
buf \U$40556 ( \40809 , \39576 );
nand \U$40557 ( \40810 , \40808 , \40809 );
or \U$40558 ( \40811 , \40807 , \40810 );
nand \U$40559 ( \40812 , \39516 , \39534 );
nand \U$40560 ( \40813 , \40811 , \40812 );
nor \U$40561 ( \40814 , \40806 , \40813 );
nand \U$40562 ( \40815 , \40803 , \40814 );
nand \U$40563 ( \40816 , \40792 , \40815 , \40753 );
not \U$40564 ( \40817 , \40547 );
not \U$40565 ( \40818 , \40675 );
and \U$40566 ( \40819 , \40721 , \40723 );
not \U$40567 ( \40820 , \40819 );
not \U$40568 ( \40821 , \40752 );
or \U$40569 ( \40822 , \40820 , \40821 );
nand \U$40570 ( \40823 , \40747 , \40745 );
nand \U$40571 ( \40824 , \40822 , \40823 );
nand \U$40572 ( \40825 , \40817 , \40818 , \40716 , \40824 );
nand \U$40573 ( \40826 , \40816 , \40825 );
buf \U$40574 ( \40827 , \40783 );
not \U$40575 ( \40828 , \40827 );
not \U$40576 ( \40829 , \39312 );
or \U$40577 ( \40830 , \40828 , \40829 );
nand \U$40578 ( \40831 , \40830 , \40823 );
and \U$40579 ( \40832 , \40826 , \40831 );
not \U$40580 ( \40833 , \39310 );
and \U$40581 ( \40834 , \40764 , \40754 );
not \U$40582 ( \40835 , \40834 );
not \U$40583 ( \40836 , \40781 );
or \U$40584 ( \40837 , \40835 , \40836 );
buf \U$40585 ( \40838 , \40775 );
buf \U$40586 ( \40839 , \40769 );
nand \U$40587 ( \40840 , \40838 , \40839 );
nand \U$40588 ( \40841 , \40837 , \40840 );
not \U$40589 ( \40842 , \39303 );
nor \U$40590 ( \40843 , \40842 , \39306 );
nor \U$40591 ( \40844 , \40841 , \40843 );
not \U$40592 ( \40845 , \40844 );
or \U$40593 ( \40846 , \40833 , \40845 );
not \U$40594 ( \40847 , \40841 );
and \U$40595 ( \40848 , \40847 , \40782 );
not \U$40596 ( \40849 , \40752 );
nor \U$40597 ( \40850 , \40848 , \40849 );
nand \U$40598 ( \40851 , \40846 , \40850 );
nor \U$40599 ( \40852 , \40851 , \40717 );
not \U$40600 ( \40853 , \40852 );
not \U$40601 ( \40854 , \38222 );
not \U$40602 ( \40855 , \40854 );
not \U$40603 ( \40856 , \38578 );
and \U$40604 ( \40857 , \37095 , \37103 );
not \U$40605 ( \40858 , \40857 );
or \U$40606 ( \40859 , \40856 , \40858 );
not \U$40607 ( \40860 , \38572 );
nand \U$40608 ( \40861 , \40860 , \38576 );
nand \U$40609 ( \40862 , \40859 , \40861 );
nand \U$40610 ( \40863 , \40855 , \40862 );
or \U$40611 ( \40864 , \38217 , \38202 );
and \U$40612 ( \40865 , \40844 , \40863 , \40864 );
nor \U$40613 ( \40866 , \38807 , \38801 );
nand \U$40614 ( \40867 , \38580 , \40866 );
and \U$40615 ( \40868 , \38562 , \38569 );
not \U$40616 ( \40869 , \40868 );
not \U$40617 ( \40870 , \36547 );
or \U$40618 ( \40871 , \40869 , \40870 );
not \U$40619 ( \40872 , \36541 );
nand \U$40620 ( \40873 , \40872 , \36545 );
nand \U$40621 ( \40874 , \40871 , \40873 );
and \U$40622 ( \40875 , \38572 , \38573 );
not \U$40623 ( \40876 , \38572 );
and \U$40624 ( \40877 , \40876 , \38576 );
nor \U$40625 ( \40878 , \40875 , \40877 );
and \U$40626 ( \40879 , \37104 , \38222 , \40878 );
nand \U$40627 ( \40880 , \40874 , \40879 );
nand \U$40628 ( \40881 , \40865 , \40867 , \40880 );
not \U$40629 ( \40882 , \40881 );
or \U$40630 ( \40883 , \40853 , \40882 );
not \U$40631 ( \40884 , \40711 );
nand \U$40632 ( \40885 , \40884 , \40708 );
not \U$40633 ( \40886 , \40885 );
nand \U$40634 ( \40887 , \40390 , \40377 );
not \U$40635 ( \40888 , \40887 );
not \U$40636 ( \40889 , \40395 );
not \U$40637 ( \40890 , \40889 );
or \U$40638 ( \40891 , \40888 , \40890 );
buf \U$40639 ( \40892 , \40715 );
not \U$40640 ( \40893 , \40892 );
nand \U$40641 ( \40894 , \40891 , \40893 );
not \U$40642 ( \40895 , \40894 );
or \U$40643 ( \40896 , \40886 , \40895 );
and \U$40644 ( \40897 , \40626 , \40673 );
and \U$40645 ( \40898 , \40625 , \40897 );
and \U$40646 ( \40899 , \40623 , \40624 );
nor \U$40647 ( \40900 , \40898 , \40899 );
not \U$40648 ( \40901 , \40900 );
and \U$40649 ( \40902 , \40677 , \40702 );
nand \U$40650 ( \40903 , \40674 , \40625 , \40902 );
not \U$40651 ( \40904 , \40903 );
or \U$40652 ( \40905 , \40901 , \40904 );
buf \U$40653 ( \40906 , \40546 );
nand \U$40654 ( \40907 , \40905 , \40906 );
not \U$40655 ( \40908 , \40534 );
nand \U$40656 ( \40909 , \40908 , \40542 );
and \U$40657 ( \40910 , \40887 , \40885 , \40909 );
nand \U$40658 ( \40911 , \40907 , \40910 );
nand \U$40659 ( \40912 , \40896 , \40911 );
nand \U$40660 ( \40913 , \40883 , \40912 );
nor \U$40661 ( \40914 , \40832 , \40913 );
nand \U$40662 ( \40915 , \40791 , \40914 );
not \U$40663 ( \40916 , \40915 );
or \U$40664 ( \40917 , \12700 , \40916 );
not \U$40665 ( \40918 , \12611 );
not \U$40666 ( \40919 , \12027 );
buf \U$40667 ( \40920 , \10585 );
not \U$40668 ( \40921 , \40920 );
not \U$40669 ( \40922 , \9736 );
not \U$40670 ( \40923 , \10210 );
not \U$40671 ( \40924 , \10202 );
and \U$40672 ( \40925 , \40923 , \40924 );
and \U$40673 ( \40926 , \10590 , \11089 );
and \U$40674 ( \40927 , \10214 , \40926 );
nor \U$40675 ( \40928 , \40925 , \40927 );
or \U$40676 ( \40929 , \40922 , \40928 );
not \U$40677 ( \40930 , \9732 );
nand \U$40678 ( \40931 , \40930 , \9334 );
nand \U$40679 ( \40932 , \40929 , \40931 );
not \U$40680 ( \40933 , \40932 );
or \U$40681 ( \40934 , \40921 , \40933 );
not \U$40682 ( \40935 , \12551 );
nor \U$40683 ( \40936 , \40935 , \12549 );
and \U$40684 ( \40937 , \11091 , \40936 );
not \U$40685 ( \40938 , \10584 );
nor \U$40686 ( \40939 , \40938 , \10216 );
nor \U$40687 ( \40940 , \40937 , \40939 );
nand \U$40688 ( \40941 , \40934 , \40940 );
not \U$40689 ( \40942 , \40941 );
or \U$40690 ( \40943 , \40919 , \40942 );
and \U$40691 ( \40944 , \11740 , \11745 );
not \U$40692 ( \40945 , \40944 );
not \U$40693 ( \40946 , \11738 );
or \U$40694 ( \40947 , \40945 , \40946 );
not \U$40695 ( \40948 , \11734 );
nand \U$40696 ( \40949 , \40948 , \11434 );
nand \U$40697 ( \40950 , \40947 , \40949 );
not \U$40698 ( \40951 , \40950 );
not \U$40699 ( \40952 , \11906 );
or \U$40700 ( \40953 , \40951 , \40952 );
not \U$40701 ( \40954 , \11901 );
nand \U$40702 ( \40955 , \40954 , \11896 );
nand \U$40703 ( \40956 , \40953 , \40955 );
and \U$40704 ( \40957 , \40956 , \12026 );
and \U$40705 ( \40958 , \12020 , \11912 );
nor \U$40706 ( \40959 , \40957 , \40958 );
nand \U$40707 ( \40960 , \40943 , \40959 );
not \U$40708 ( \40961 , \40960 );
or \U$40709 ( \40962 , \40918 , \40961 );
nand \U$40710 ( \40963 , \12606 , \12610 );
nand \U$40711 ( \40964 , \40962 , \40963 );
and \U$40712 ( \40965 , \12698 , \40964 );
not \U$40713 ( \40966 , \12669 );
nand \U$40714 ( \40967 , \12649 , \12650 );
not \U$40715 ( \40968 , \40967 );
and \U$40716 ( \40969 , \40966 , \40968 );
and \U$40717 ( \40970 , \12653 , \12668 );
nor \U$40718 ( \40971 , \40969 , \40970 );
not \U$40719 ( \40972 , \40971 );
not \U$40720 ( \40973 , \12697 );
and \U$40721 ( \40974 , \40972 , \40973 );
and \U$40722 ( \40975 , \12672 , \12687 );
and \U$40723 ( \40976 , \40975 , \12696 );
nor \U$40724 ( \40977 , \40974 , \40976 );
not \U$40725 ( \40978 , \40977 );
nor \U$40726 ( \40979 , \40965 , \40978 );
nand \U$40727 ( \40980 , \40917 , \40979 );
not \U$40728 ( \40981 , \40980 );
or \U$40729 ( \40982 , \6298 , \40981 );
not \U$40730 ( \40983 , \5315 );
not \U$40731 ( \40984 , \5338 );
or \U$40732 ( \40985 , \40983 , \40984 );
not \U$40733 ( \40986 , \5339 );
not \U$40734 ( \40987 , \40986 );
nand \U$40735 ( \40988 , \5310 , \5027 );
not \U$40736 ( \40989 , \40988 );
and \U$40737 ( \40990 , \40987 , \40989 );
not \U$40738 ( \40991 , \6275 );
nor \U$40739 ( \40992 , \40991 , \6273 );
and \U$40740 ( \40993 , \40992 , \5939 );
nand \U$40741 ( \40994 , \5938 , \5937 );
not \U$40742 ( \40995 , \40994 );
nor \U$40743 ( \40996 , \40993 , \40995 );
or \U$40744 ( \40997 , \40996 , \5635 );
not \U$40745 ( \40998 , \5341 );
nand \U$40746 ( \40999 , \40998 , \5634 );
nand \U$40747 ( \41000 , \40997 , \40999 );
and \U$40748 ( \41001 , \41000 , \5340 );
nor \U$40749 ( \41002 , \40990 , \41001 );
nand \U$40750 ( \41003 , \40985 , \41002 );
not \U$40751 ( \41004 , \41003 );
not \U$40752 ( \41005 , \6295 );
or \U$40753 ( \41006 , \41004 , \41005 );
nand \U$40754 ( \41007 , \6294 , \6293 );
nand \U$40755 ( \41008 , \41006 , \41007 );
and \U$40756 ( \41009 , \41008 , \6292 );
nor \U$40757 ( \41010 , \6282 , \6291 );
nor \U$40758 ( \41011 , \41009 , \41010 );
not \U$40759 ( \41012 , \41011 );
not \U$40760 ( \41013 , \4143 );
and \U$40761 ( \41014 , \41012 , \41013 );
not \U$40762 ( \41015 , \6296 );
not \U$40763 ( \41016 , \41015 );
not \U$40764 ( \41017 , \12690 );
nand \U$40765 ( \41018 , \41017 , \12691 );
nor \U$40766 ( \41019 , \4143 , \41018 );
not \U$40767 ( \41020 , \41019 );
or \U$40768 ( \41021 , \41016 , \41020 );
and \U$40769 ( \41022 , \4127 , \4135 );
not \U$40770 ( \41023 , \4142 );
not \U$40771 ( \41024 , \3619 );
nand \U$40772 ( \41025 , \41024 , \4118 );
or \U$40773 ( \41026 , \41023 , \41025 );
not \U$40774 ( \41027 , \4141 );
nand \U$40775 ( \41028 , \41027 , \4137 );
nand \U$40776 ( \41029 , \41026 , \41028 );
and \U$40777 ( \41030 , \41029 , \4136 );
nor \U$40778 ( \41031 , \41022 , \41030 );
nand \U$40779 ( \41032 , \41021 , \41031 );
nor \U$40780 ( \41033 , \41014 , \41032 );
nand \U$40781 ( \41034 , \40982 , \41033 );
not \U$40782 ( \41035 , \41034 );
or \U$40783 ( \41036 , \3150 , \41035 );
not \U$40784 ( \41037 , \2937 );
nand \U$40785 ( \41038 , \41037 , \2943 );
or \U$40786 ( \41039 , \2728 , \41038 );
not \U$40787 ( \41040 , \2718 );
nand \U$40788 ( \41041 , \41040 , \2724 );
nand \U$40789 ( \41042 , \41039 , \41041 );
not \U$40790 ( \41043 , \41042 );
or \U$40791 ( \41044 , \41043 , \2516 );
not \U$40792 ( \41045 , \2515 );
nand \U$40793 ( \41046 , \41045 , \2302 );
nand \U$40794 ( \41047 , \41044 , \41046 );
and \U$40795 ( \41048 , \2297 , \41047 );
not \U$40796 ( \41049 , \2024 );
nand \U$40797 ( \41050 , \41049 , \2166 );
or \U$40798 ( \41051 , \2296 , \41050 );
or \U$40799 ( \41052 , \2293 , \2295 );
nand \U$40800 ( \41053 , \41051 , \41052 );
nor \U$40801 ( \41054 , \41048 , \41053 );
not \U$40802 ( \41055 , \41054 );
not \U$40803 ( \41056 , \3148 );
and \U$40804 ( \41057 , \41055 , \41056 );
not \U$40805 ( \41058 , \3137 );
nand \U$40806 ( \41059 , \41058 , \3135 );
not \U$40807 ( \41060 , \41059 );
not \U$40808 ( \41061 , \3146 );
and \U$40809 ( \41062 , \41060 , \41061 );
not \U$40810 ( \41063 , \3144 );
nand \U$40811 ( \41064 , \41063 , \3145 );
not \U$40812 ( \41065 , \41064 );
nor \U$40813 ( \41066 , \41062 , \41065 );
or \U$40814 ( \41067 , \41066 , \3113 );
or \U$40815 ( \41068 , \3027 , \2955 );
and \U$40816 ( \41069 , \3076 , \3111 );
and \U$40817 ( \41070 , \3071 , \41069 );
not \U$40818 ( \41071 , \3061 );
nand \U$40819 ( \41072 , \41071 , \3067 );
not \U$40820 ( \41073 , \41072 );
nor \U$40821 ( \41074 , \41070 , \41073 );
or \U$40822 ( \41075 , \3028 , \41074 );
nand \U$40823 ( \41076 , \41067 , \41068 , \41075 );
nor \U$40824 ( \41077 , \41057 , \41076 );
nand \U$40825 ( \41078 , \41036 , \41077 );
not \U$40826 ( \41079 , \41078 );
or \U$40827 ( \41080 , \1071 , \41079 );
not \U$40828 ( \41081 , \1064 );
nand \U$40829 ( \41082 , \41081 , \1066 );
nand \U$40830 ( \41083 , \41080 , \41082 );
not \U$40831 ( \41084 , \41083 );
or \U$40832 ( \41085 , \941 , \41084 );
not \U$40833 ( \41086 , \904 );
nand \U$40834 ( \41087 , \41086 , \858 );
not \U$40835 ( \41088 , \41087 );
and \U$40836 ( \41089 , \939 , \41088 );
not \U$40837 ( \41090 , \934 );
nor \U$40838 ( \41091 , \41090 , \932 );
and \U$40839 ( \41092 , \41091 , \927 );
and \U$40840 ( \41093 , \913 , \926 );
nor \U$40841 ( \41094 , \41089 , \41092 , \41093 );
nand \U$40842 ( \41095 , \41085 , \41094 );
nor \U$40843 ( \41096 , \537 , \41095 );
not \U$40844 ( \41097 , \41096 );
not \U$40845 ( \41098 , \536 );
nand \U$40846 ( \41099 , \41098 , \41095 );
nand \U$40847 ( \41100 , \41097 , \41099 );
xor \U$40848 ( \41101 , \41083 , \908 );
buf \U$40849 ( \41102 , \41078 );
xor \U$40850 ( \41103 , \41102 , \1070 );
nand \U$40851 ( \41104 , \41101 , \41103 );
not \U$40852 ( \41105 , \2517 );
not \U$40853 ( \41106 , \2729 );
not \U$40854 ( \41107 , \41033 );
not \U$40855 ( \41108 , \2948 );
not \U$40856 ( \41109 , \41108 );
and \U$40857 ( \41110 , \41107 , \41109 );
and \U$40858 ( \41111 , \6297 , \2948 );
and \U$40859 ( \41112 , \40980 , \41111 );
nor \U$40860 ( \41113 , \41110 , \41112 );
nand \U$40861 ( \41114 , \41113 , \41038 );
not \U$40862 ( \41115 , \41114 );
or \U$40863 ( \41116 , \41106 , \41115 );
nand \U$40864 ( \41117 , \41116 , \41041 );
not \U$40865 ( \41118 , \41117 );
or \U$40866 ( \41119 , \41105 , \41118 );
nand \U$40867 ( \41120 , \41119 , \41046 );
not \U$40868 ( \41121 , \2167 );
and \U$40869 ( \41122 , \41120 , \41121 );
not \U$40870 ( \41123 , \41120 );
and \U$40871 ( \41124 , \41123 , \2167 );
or \U$40872 ( \41125 , \41122 , \41124 );
nor \U$40873 ( \41126 , \41104 , \41125 );
and \U$40874 ( \41127 , \41100 , \41126 );
not \U$40875 ( \41128 , \41127 );
not \U$40876 ( \41129 , \536 );
not \U$40877 ( \41130 , \41095 );
or \U$40878 ( \41131 , \41129 , \41130 );
not \U$40879 ( \41132 , \492 );
nand \U$40880 ( \41133 , \41132 , \532 );
nand \U$40881 ( \41134 , \41131 , \41133 );
nand \U$40882 ( \41135 , RIbe29380_53, RIbe28e58_42);
not \U$40883 ( \41136 , \41135 );
nand \U$40884 ( \41137 , \261 , RIbe27b98_2);
and \U$40885 ( \41138 , \41137 , \271 );
not \U$40886 ( \41139 , \41137 );
and \U$40887 ( \41140 , \41139 , \272 );
nor \U$40888 ( \41141 , \41138 , \41140 );
not \U$40889 ( \41142 , \41141 );
or \U$40890 ( \41143 , \41136 , \41142 );
or \U$40891 ( \41144 , \41141 , \41135 );
nand \U$40892 ( \41145 , \41143 , \41144 );
not \U$40893 ( \41146 , \41145 );
and \U$40894 ( \41147 , \327 , RIbe28de0_41);
and \U$40895 ( \41148 , \331 , RIbe29920_65);
nor \U$40896 ( \41149 , \41147 , \41148 );
and \U$40897 ( \41150 , \41149 , \342 );
not \U$40898 ( \41151 , \41149 );
and \U$40899 ( \41152 , \41151 , \339 );
nor \U$40900 ( \41153 , \41150 , \41152 );
not \U$40901 ( \41154 , \41153 );
and \U$40902 ( \41155 , \41146 , \41154 );
and \U$40903 ( \41156 , \41145 , \41153 );
nor \U$40904 ( \41157 , \41155 , \41156 );
xor \U$40905 ( \41158 , \513 , \293 );
and \U$40906 ( \41159 , \41158 , \521 );
and \U$40907 ( \41160 , \513 , \293 );
or \U$40908 ( \41161 , \41159 , \41160 );
or \U$40909 ( \41162 , \41157 , \41161 );
nand \U$40910 ( \41163 , \41157 , \41161 );
nand \U$40911 ( \41164 , \41162 , \41163 );
not \U$40912 ( \41165 , \41164 );
xor \U$40913 ( \41166 , \499 , \500 );
and \U$40914 ( \41167 , \41166 , \505 );
and \U$40915 ( \41168 , \499 , \500 );
or \U$40916 ( \41169 , \41167 , \41168 );
xor \U$40917 ( \41170 , \41165 , \41169 );
xor \U$40918 ( \41171 , \499 , \500 );
xor \U$40919 ( \41172 , \41171 , \505 );
and \U$40920 ( \41173 , \522 , \41172 );
xor \U$40921 ( \41174 , \499 , \500 );
xor \U$40922 ( \41175 , \41174 , \505 );
and \U$40923 ( \41176 , \526 , \41175 );
and \U$40924 ( \41177 , \522 , \526 );
or \U$40925 ( \41178 , \41173 , \41176 , \41177 );
xor \U$40926 ( \41179 , \41170 , \41178 );
not \U$40927 ( \41180 , \528 );
nand \U$40928 ( \41181 , \41180 , \497 );
xor \U$40929 ( \41182 , \41179 , \41181 );
and \U$40930 ( \41183 , \41134 , \41182 );
not \U$40931 ( \41184 , \41134 );
not \U$40932 ( \41185 , \41182 );
and \U$40933 ( \41186 , \41184 , \41185 );
nor \U$40934 ( \41187 , \41183 , \41186 );
buf \U$40935 ( \41188 , \11739 );
not \U$40936 ( \41189 , \41188 );
not \U$40937 ( \41190 , \41189 );
not \U$40938 ( \41191 , \11746 );
not \U$40939 ( \41192 , \11092 );
not \U$40940 ( \41193 , \40915 );
not \U$40941 ( \41194 , \12555 );
nor \U$40942 ( \41195 , \41193 , \41194 );
not \U$40943 ( \41196 , \41195 );
or \U$40944 ( \41197 , \41192 , \41196 );
not \U$40945 ( \41198 , \40941 );
nand \U$40946 ( \41199 , \41197 , \41198 );
not \U$40947 ( \41200 , \41199 );
or \U$40948 ( \41201 , \41191 , \41200 );
not \U$40949 ( \41202 , \40944 );
nand \U$40950 ( \41203 , \41201 , \41202 );
buf \U$40951 ( \41204 , \41203 );
not \U$40952 ( \41205 , \41204 );
or \U$40953 ( \41206 , \41190 , \41205 );
or \U$40954 ( \41207 , \41189 , \41204 );
nand \U$40955 ( \41208 , \41206 , \41207 );
buf \U$40956 ( \41209 , \41199 );
xor \U$40957 ( \41210 , \11746 , \41209 );
and \U$40958 ( \41211 , \11092 , \12612 );
not \U$40959 ( \41212 , \41211 );
not \U$40960 ( \41213 , \40915 );
or \U$40961 ( \41214 , \41212 , \41213 );
not \U$40962 ( \41215 , \40964 );
nand \U$40963 ( \41216 , \41214 , \41215 );
not \U$40964 ( \41217 , \12651 );
and \U$40965 ( \41218 , \41216 , \41217 );
not \U$40966 ( \41219 , \41216 );
and \U$40967 ( \41220 , \41219 , \12651 );
nor \U$40968 ( \41221 , \41218 , \41220 );
nand \U$40969 ( \41222 , \41210 , \41221 );
buf \U$40970 ( \41223 , \40915 );
and \U$40971 ( \41224 , \41223 , \11092 , \12555 );
buf \U$40972 ( \41225 , \12027 );
and \U$40973 ( \41226 , \41224 , \41225 );
buf \U$40974 ( \41227 , \40960 );
nor \U$40975 ( \41228 , \41226 , \41227 );
xor \U$40976 ( \41229 , \41228 , \12611 );
nor \U$40977 ( \41230 , \41222 , \41229 );
not \U$40978 ( \41231 , \5939 );
not \U$40979 ( \41232 , \6279 );
not \U$40980 ( \41233 , \12699 );
not \U$40981 ( \41234 , \40915 );
or \U$40982 ( \41235 , \41233 , \41234 );
and \U$40983 ( \41236 , \12698 , \40964 );
nand \U$40984 ( \41237 , \40977 , \41018 );
nor \U$40985 ( \41238 , \41236 , \41237 );
nand \U$40986 ( \41239 , \41235 , \41238 );
not \U$40987 ( \41240 , \41239 );
or \U$40988 ( \41241 , \41232 , \41240 );
not \U$40989 ( \41242 , \6273 );
nand \U$40990 ( \41243 , \41242 , \6275 );
nand \U$40991 ( \41244 , \41241 , \41243 );
not \U$40992 ( \41245 , \41244 );
or \U$40993 ( \41246 , \41231 , \41245 );
nand \U$40994 ( \41247 , \41246 , \40994 );
and \U$40995 ( \41248 , \41247 , \5636 );
not \U$40996 ( \41249 , \41247 );
and \U$40997 ( \41250 , \41249 , \5635 );
nor \U$40998 ( \41251 , \41248 , \41250 );
not \U$40999 ( \41252 , \10214 );
buf \U$41000 ( \41253 , \11090 );
not \U$41001 ( \41254 , \41253 );
nor \U$41002 ( \41255 , \41252 , \41254 );
not \U$41003 ( \41256 , \41255 );
not \U$41004 ( \41257 , \12555 );
not \U$41005 ( \41258 , \40915 );
or \U$41006 ( \41259 , \41257 , \41258 );
not \U$41007 ( \41260 , \40936 );
nand \U$41008 ( \41261 , \41259 , \41260 );
not \U$41009 ( \41262 , \41261 );
or \U$41010 ( \41263 , \41256 , \41262 );
buf \U$41011 ( \41264 , \40928 );
nand \U$41012 ( \41265 , \41263 , \41264 );
not \U$41013 ( \41266 , \41265 );
not \U$41014 ( \41267 , \41266 );
not \U$41015 ( \41268 , \9736 );
or \U$41016 ( \41269 , \41267 , \41268 );
nand \U$41017 ( \41270 , \41265 , \40922 );
nand \U$41018 ( \41271 , \41269 , \41270 );
and \U$41019 ( \41272 , \41208 , \41230 , \41251 , \41271 );
not \U$41020 ( \41273 , \41188 );
not \U$41021 ( \41274 , \41203 );
or \U$41022 ( \41275 , \41273 , \41274 );
nand \U$41023 ( \41276 , \41275 , \40949 );
nand \U$41024 ( \41277 , \11906 , \41276 );
nand \U$41025 ( \41278 , \41277 , \40955 );
nand \U$41026 ( \41279 , \41278 , \12026 );
nand \U$41027 ( \41280 , \41272 , \41279 );
not \U$41028 ( \41281 , \12026 );
not \U$41029 ( \41282 , \41281 );
not \U$41030 ( \41283 , \41278 );
not \U$41031 ( \41284 , \41283 );
or \U$41032 ( \41285 , \41282 , \41284 );
and \U$41033 ( \41286 , \41276 , \11906 );
not \U$41034 ( \41287 , \41276 );
not \U$41035 ( \41288 , \11906 );
and \U$41036 ( \41289 , \41287 , \41288 );
nor \U$41037 ( \41290 , \41286 , \41289 );
nand \U$41038 ( \41291 , \41285 , \41290 );
nor \U$41039 ( \41292 , \41280 , \41291 );
not \U$41040 ( \41293 , \938 );
not \U$41041 ( \41294 , \908 );
not \U$41042 ( \41295 , \41083 );
or \U$41043 ( \41296 , \41294 , \41295 );
nand \U$41044 ( \41297 , \41296 , \41087 );
not \U$41045 ( \41298 , \41297 );
or \U$41046 ( \41299 , \41293 , \41298 );
or \U$41047 ( \41300 , \938 , \41297 );
nand \U$41048 ( \41301 , \41299 , \41300 );
nand \U$41049 ( \41302 , \41187 , \41292 , \41301 );
nor \U$41050 ( \41303 , \41128 , \41302 );
not \U$41051 ( \41304 , \41303 );
not \U$41052 ( \41305 , \40818 );
not \U$41053 ( \41306 , \40752 );
not \U$41054 ( \41307 , \40867 );
nand \U$41055 ( \41308 , \40880 , \40863 , \40864 );
nor \U$41056 ( \41309 , \41307 , \41308 );
buf \U$41057 ( \41310 , \39310 );
or \U$41058 ( \41311 , \41309 , \41310 );
not \U$41059 ( \41312 , \40843 );
nand \U$41060 ( \41313 , \41311 , \41312 );
not \U$41061 ( \41314 , \41313 );
not \U$41062 ( \41315 , \40827 );
or \U$41063 ( \41316 , \41314 , \41315 );
nand \U$41064 ( \41317 , \41316 , \40847 );
not \U$41065 ( \41318 , \41317 );
or \U$41066 ( \41319 , \41306 , \41318 );
not \U$41067 ( \41320 , \32121 );
not \U$41068 ( \41321 , \41320 );
buf \U$41069 ( \41322 , \39313 );
nor \U$41070 ( \41323 , \41322 , \39638 , \40788 );
and \U$41071 ( \41324 , \41321 , \41323 );
not \U$41072 ( \41325 , \40815 );
not \U$41073 ( \41326 , \40753 );
or \U$41074 ( \41327 , \41325 , \41326 );
not \U$41075 ( \41328 , \40824 );
nand \U$41076 ( \41329 , \41327 , \41328 );
nand \U$41077 ( \41330 , \40831 , \41329 );
not \U$41078 ( \41331 , \41330 );
nor \U$41079 ( \41332 , \41324 , \41331 );
nand \U$41080 ( \41333 , \41319 , \41332 );
buf \U$41081 ( \41334 , \40703 );
nand \U$41082 ( \41335 , \41333 , \41334 );
not \U$41083 ( \41336 , \40902 );
nand \U$41084 ( \41337 , \41335 , \41336 );
not \U$41085 ( \41338 , \41337 );
or \U$41086 ( \41339 , \41305 , \41338 );
nand \U$41087 ( \41340 , \41339 , \40900 );
xor \U$41088 ( \41341 , \41340 , \40906 );
not \U$41089 ( \41342 , \40674 );
or \U$41090 ( \41343 , \41342 , \41335 );
nor \U$41091 ( \41344 , \41342 , \41336 );
nor \U$41092 ( \41345 , \41344 , \40897 );
nand \U$41093 ( \41346 , \41343 , \41345 );
not \U$41094 ( \41347 , \41346 );
not \U$41095 ( \41348 , \40625 );
not \U$41096 ( \41349 , \41348 );
and \U$41097 ( \41350 , \41347 , \41349 );
and \U$41098 ( \41351 , \41346 , \41348 );
nor \U$41099 ( \41352 , \41350 , \41351 );
nand \U$41100 ( \41353 , \41335 , \41336 );
and \U$41101 ( \41354 , \41353 , \41342 );
not \U$41102 ( \41355 , \41353 );
and \U$41103 ( \41356 , \41355 , \40674 );
nor \U$41104 ( \41357 , \41354 , \41356 );
nor \U$41105 ( \41358 , \41352 , \41357 );
nand \U$41106 ( \41359 , \41341 , \41358 );
buf \U$41107 ( \41360 , \37105 );
buf \U$41108 ( \41361 , \38578 );
not \U$41109 ( \41362 , \41361 );
nor \U$41110 ( \41363 , \41360 , \41362 );
not \U$41111 ( \41364 , \41363 );
not \U$41112 ( \41365 , \38570 );
not \U$41113 ( \41366 , \38808 );
not \U$41114 ( \41367 , \41366 );
not \U$41115 ( \41368 , \40724 );
not \U$41116 ( \41369 , \32120 );
not \U$41117 ( \41370 , \32085 );
or \U$41118 ( \41371 , \41369 , \41370 );
and \U$41119 ( \41372 , \39585 , \39614 , \40787 , \39637 );
nand \U$41120 ( \41373 , \41371 , \41372 );
nand \U$41121 ( \41374 , \41373 , \41325 );
not \U$41122 ( \41375 , \41374 );
or \U$41123 ( \41376 , \41368 , \41375 );
not \U$41124 ( \41377 , \40819 );
nand \U$41125 ( \41378 , \41376 , \41377 );
not \U$41126 ( \41379 , \41378 );
or \U$41127 ( \41380 , \41367 , \41379 );
not \U$41128 ( \41381 , \40866 );
nand \U$41129 ( \41382 , \41380 , \41381 );
not \U$41130 ( \41383 , \41382 );
or \U$41131 ( \41384 , \41365 , \41383 );
not \U$41132 ( \41385 , \40868 );
nand \U$41133 ( \41386 , \41384 , \41385 );
not \U$41134 ( \41387 , \41386 );
or \U$41135 ( \41388 , \41364 , \41387 );
buf \U$41136 ( \41389 , \37104 );
not \U$41137 ( \41390 , \40873 );
and \U$41138 ( \41391 , \41389 , \41390 , \41361 );
nor \U$41139 ( \41392 , \41391 , \40862 );
nand \U$41140 ( \41393 , \41388 , \41392 );
buf \U$41141 ( \41394 , \40854 );
xor \U$41142 ( \41395 , \41393 , \41394 );
nor \U$41143 ( \41396 , \41359 , \41395 );
not \U$41144 ( \41397 , \41378 );
buf \U$41145 ( \41398 , \41322 );
nor \U$41146 ( \41399 , \41397 , \41398 );
and \U$41147 ( \41400 , \41399 , \40827 );
nor \U$41148 ( \41401 , \41400 , \41317 );
not \U$41149 ( \41402 , \41401 );
not \U$41150 ( \41403 , \40849 );
and \U$41151 ( \41404 , \41402 , \41403 );
and \U$41152 ( \41405 , \41401 , \40849 );
nor \U$41153 ( \41406 , \41404 , \41405 );
not \U$41154 ( \41407 , \41334 );
not \U$41155 ( \41408 , \41333 );
not \U$41156 ( \41409 , \41408 );
or \U$41157 ( \41410 , \41407 , \41409 );
or \U$41158 ( \41411 , \41408 , \41334 );
nand \U$41159 ( \41412 , \41410 , \41411 );
nand \U$41160 ( \41413 , \41406 , \41412 );
not \U$41161 ( \41414 , \41413 );
buf \U$41162 ( \41415 , \40781 );
not \U$41163 ( \41416 , \41415 );
not \U$41164 ( \41417 , \41416 );
buf \U$41165 ( \41418 , \40834 );
not \U$41166 ( \41419 , \41418 );
not \U$41167 ( \41420 , \41398 );
not \U$41168 ( \41421 , \41420 );
not \U$41169 ( \41422 , \41378 );
or \U$41170 ( \41423 , \41421 , \41422 );
not \U$41171 ( \41424 , \41313 );
nand \U$41172 ( \41425 , \41423 , \41424 );
buf \U$41173 ( \41426 , \40765 );
nand \U$41174 ( \41427 , \41425 , \41426 );
nand \U$41175 ( \41428 , \41419 , \41427 );
not \U$41176 ( \41429 , \41428 );
or \U$41177 ( \41430 , \41417 , \41429 );
nor \U$41178 ( \41431 , \41416 , \41418 );
nand \U$41179 ( \41432 , \41427 , \41431 );
nand \U$41180 ( \41433 , \41430 , \41432 );
nand \U$41181 ( \41434 , \41414 , \41433 );
buf \U$41182 ( \41435 , \36547 );
and \U$41183 ( \41436 , \41435 , \38570 );
not \U$41184 ( \41437 , \41436 );
not \U$41185 ( \41438 , \41382 );
or \U$41186 ( \41439 , \41437 , \41438 );
not \U$41187 ( \41440 , \40874 );
nand \U$41188 ( \41441 , \41439 , \41440 );
or \U$41189 ( \41442 , \41389 , \41441 );
xor \U$41190 ( \41443 , \41425 , \41426 );
nand \U$41191 ( \41444 , \41442 , \41443 );
not \U$41192 ( \41445 , \41444 );
nand \U$41193 ( \41446 , \41441 , \41389 );
xor \U$41194 ( \41447 , \5939 , \41244 );
nand \U$41195 ( \41448 , \41445 , \41446 , \41447 );
nor \U$41196 ( \41449 , \41434 , \41448 );
not \U$41197 ( \41450 , \12696 );
not \U$41198 ( \41451 , \41450 );
not \U$41199 ( \41452 , \41216 );
not \U$41200 ( \41453 , \12670 );
or \U$41201 ( \41454 , \41452 , \41453 );
nand \U$41202 ( \41455 , \41454 , \40971 );
and \U$41203 ( \41456 , \41455 , \12688 );
nor \U$41204 ( \41457 , \41456 , \40975 );
not \U$41205 ( \41458 , \41457 );
or \U$41206 ( \41459 , \41451 , \41458 );
or \U$41207 ( \41460 , \41457 , \41450 );
nand \U$41208 ( \41461 , \41459 , \41460 );
nor \U$41209 ( \41462 , \41360 , \38579 );
not \U$41210 ( \41463 , \41462 );
not \U$41211 ( \41464 , \41382 );
or \U$41212 ( \41465 , \41463 , \41464 );
not \U$41213 ( \41466 , \41308 );
nand \U$41214 ( \41467 , \41465 , \41466 );
not \U$41215 ( \41468 , \41467 );
not \U$41216 ( \41469 , \41310 );
and \U$41217 ( \41470 , \41468 , \41469 );
and \U$41218 ( \41471 , \41467 , \41310 );
nor \U$41219 ( \41472 , \41470 , \41471 );
nor \U$41220 ( \41473 , \41461 , \41472 );
and \U$41221 ( \41474 , \41396 , \41449 , \41473 );
buf \U$41222 ( \41475 , \41474 );
not \U$41223 ( \41476 , \3147 );
not \U$41224 ( \41477 , \2949 );
not \U$41225 ( \41478 , \41034 );
or \U$41226 ( \41479 , \41477 , \41478 );
buf \U$41227 ( \41480 , \41054 );
nand \U$41228 ( \41481 , \41479 , \41480 );
not \U$41229 ( \41482 , \41481 );
or \U$41230 ( \41483 , \41476 , \41482 );
nand \U$41231 ( \41484 , \41483 , \41066 );
and \U$41232 ( \41485 , \41484 , \3112 );
nor \U$41233 ( \41486 , \41485 , \41069 );
not \U$41234 ( \41487 , \3071 );
and \U$41235 ( \41488 , \41486 , \41487 );
not \U$41236 ( \41489 , \41486 );
and \U$41237 ( \41490 , \41489 , \3071 );
nor \U$41238 ( \41491 , \41488 , \41490 );
not \U$41239 ( \41492 , \3146 );
not \U$41240 ( \41493 , \41492 );
not \U$41241 ( \41494 , \3138 );
not \U$41242 ( \41495 , \41494 );
not \U$41243 ( \41496 , \41481 );
or \U$41244 ( \41497 , \41495 , \41496 );
nand \U$41245 ( \41498 , \41497 , \41059 );
not \U$41246 ( \41499 , \41498 );
or \U$41247 ( \41500 , \41493 , \41499 );
nand \U$41248 ( \41501 , \41500 , \41064 );
xor \U$41249 ( \41502 , \41501 , \3112 );
and \U$41250 ( \41503 , \41475 , \41491 , \41502 );
not \U$41251 ( \41504 , \40986 );
not \U$41252 ( \41505 , \5314 );
nand \U$41253 ( \41506 , \41247 , \5636 );
nand \U$41254 ( \41507 , \41506 , \40999 );
not \U$41255 ( \41508 , \41507 );
or \U$41256 ( \41509 , \41505 , \41508 );
nand \U$41257 ( \41510 , \41509 , \40988 );
not \U$41258 ( \41511 , \41510 );
or \U$41259 ( \41512 , \41504 , \41511 );
not \U$41260 ( \41513 , \41510 );
nand \U$41261 ( \41514 , \41513 , \5339 );
nand \U$41262 ( \41515 , \41512 , \41514 );
not \U$41263 ( \41516 , \6280 );
not \U$41264 ( \41517 , \41239 );
or \U$41265 ( \41518 , \41516 , \41517 );
not \U$41266 ( \41519 , \41003 );
nand \U$41267 ( \41520 , \41518 , \41519 );
xor \U$41268 ( \41521 , \41520 , \6295 );
xor \U$41269 ( \41522 , \41034 , \2948 );
not \U$41270 ( \41523 , \41015 );
not \U$41271 ( \41524 , \41239 );
or \U$41272 ( \41525 , \41523 , \41524 );
nand \U$41273 ( \41526 , \41525 , \41011 );
xor \U$41274 ( \41527 , \41526 , \4122 );
nand \U$41275 ( \41528 , \41521 , \41522 , \41527 );
not \U$41276 ( \41529 , \6295 );
not \U$41277 ( \41530 , \41520 );
or \U$41278 ( \41531 , \41529 , \41530 );
nand \U$41279 ( \41532 , \41531 , \41007 );
xnor \U$41280 ( \41533 , \41532 , \6292 );
nor \U$41281 ( \41534 , \41528 , \41533 );
not \U$41282 ( \41535 , \4122 );
not \U$41283 ( \41536 , \41526 );
or \U$41284 ( \41537 , \41535 , \41536 );
nand \U$41285 ( \41538 , \41537 , \41025 );
and \U$41286 ( \41539 , \41538 , \4142 );
not \U$41287 ( \41540 , \41538 );
and \U$41288 ( \41541 , \41540 , \41023 );
nor \U$41289 ( \41542 , \41539 , \41541 );
and \U$41290 ( \41543 , \41534 , \41542 );
not \U$41291 ( \41544 , \4142 );
not \U$41292 ( \41545 , \41538 );
or \U$41293 ( \41546 , \41544 , \41545 );
nand \U$41294 ( \41547 , \41546 , \41028 );
xor \U$41295 ( \41548 , \41547 , \4136 );
nand \U$41296 ( \41549 , \41506 , \40999 , \5314 );
not \U$41297 ( \41550 , \40999 );
not \U$41298 ( \41551 , \41506 );
or \U$41299 ( \41552 , \41550 , \41551 );
not \U$41300 ( \41553 , \5314 );
nand \U$41301 ( \41554 , \41552 , \41553 );
nand \U$41302 ( \41555 , \41549 , \41554 );
and \U$41303 ( \41556 , \41543 , \41548 , \41555 );
and \U$41304 ( \41557 , \41515 , \41556 );
or \U$41305 ( \41558 , \41486 , \41487 );
nand \U$41306 ( \41559 , \41558 , \41072 );
not \U$41307 ( \41560 , \41559 );
not \U$41308 ( \41561 , \3028 );
and \U$41309 ( \41562 , \41560 , \41561 );
and \U$41310 ( \41563 , \41559 , \3028 );
nor \U$41311 ( \41564 , \41562 , \41563 );
not \U$41312 ( \41565 , \41564 );
nand \U$41313 ( \41566 , \41503 , \41557 , \41565 );
nor \U$41314 ( \41567 , \41304 , \41566 );
nand \U$41315 ( \41568 , \327 , RIbe27b98_2);
and \U$41316 ( \41569 , \41568 , \342 );
not \U$41317 ( \41570 , \41568 );
and \U$41318 ( \41571 , \41570 , \339 );
nor \U$41319 ( \41572 , \41569 , \41571 );
nand \U$41320 ( \41573 , RIbe29380_53, RIbe29920_65);
or \U$41321 ( \41574 , \41572 , \41573 );
nand \U$41322 ( \41575 , \41572 , \41573 );
nand \U$41323 ( \41576 , \41574 , \41575 );
not \U$41324 ( \41577 , RIbe29380_53);
nor \U$41325 ( \41578 , \41577 , \2890 );
xor \U$41326 ( \41579 , \271 , \41578 );
and \U$41327 ( \41580 , \327 , RIbe29920_65);
and \U$41328 ( \41581 , \331 , RIbe27b98_2);
nor \U$41329 ( \41582 , \41580 , \41581 );
and \U$41330 ( \41583 , \41582 , \339 );
not \U$41331 ( \41584 , \41582 );
and \U$41332 ( \41585 , \41584 , \342 );
nor \U$41333 ( \41586 , \41583 , \41585 );
and \U$41334 ( \41587 , \41579 , \41586 );
and \U$41335 ( \41588 , \271 , \41578 );
or \U$41336 ( \41589 , \41587 , \41588 );
xor \U$41337 ( \41590 , \41576 , \41589 );
or \U$41338 ( \41591 , \41153 , \41135 );
not \U$41339 ( \41592 , \41135 );
not \U$41340 ( \41593 , \41153 );
or \U$41341 ( \41594 , \41592 , \41593 );
nand \U$41342 ( \41595 , \41594 , \41141 );
nand \U$41343 ( \41596 , \41591 , \41595 );
xor \U$41344 ( \41597 , \271 , \41578 );
xor \U$41345 ( \41598 , \41597 , \41586 );
xor \U$41346 ( \41599 , \41596 , \41598 );
and \U$41347 ( \41600 , \41599 , \41163 );
and \U$41348 ( \41601 , \41596 , \41598 );
or \U$41349 ( \41602 , \41600 , \41601 );
xor \U$41350 ( \41603 , \41590 , \41602 );
xor \U$41351 ( \41604 , \41165 , \41169 );
and \U$41352 ( \41605 , \41604 , \41178 );
and \U$41353 ( \41606 , \41165 , \41169 );
or \U$41354 ( \41607 , \41605 , \41606 );
not \U$41355 ( \41608 , \41607 );
xor \U$41356 ( \41609 , \41596 , \41598 );
xor \U$41357 ( \41610 , \41609 , \41163 );
not \U$41358 ( \41611 , \41610 );
and \U$41359 ( \41612 , \41608 , \41611 );
and \U$41360 ( \41613 , \41607 , \41610 );
nor \U$41361 ( \41614 , \41612 , \41613 );
not \U$41362 ( \41615 , \41614 );
not \U$41363 ( \41616 , \41615 );
not \U$41364 ( \41617 , \940 );
nand \U$41365 ( \41618 , \41182 , \536 );
nor \U$41366 ( \41619 , \41617 , \41618 );
not \U$41367 ( \41620 , \41619 );
not \U$41368 ( \41621 , \41083 );
or \U$41369 ( \41622 , \41620 , \41621 );
or \U$41370 ( \41623 , \41094 , \41618 );
or \U$41371 ( \41624 , \41133 , \41185 );
or \U$41372 ( \41625 , \41181 , \41179 );
nand \U$41373 ( \41626 , \41623 , \41624 , \41625 );
not \U$41374 ( \41627 , \41626 );
nand \U$41375 ( \41628 , \41622 , \41627 );
not \U$41376 ( \41629 , \41628 );
or \U$41377 ( \41630 , \41616 , \41629 );
not \U$41378 ( \41631 , \41607 );
nand \U$41379 ( \41632 , \41631 , \41610 );
nand \U$41380 ( \41633 , \41630 , \41632 );
xor \U$41381 ( \41634 , \41603 , \41633 );
xnor \U$41382 ( \41635 , \41614 , \41628 );
not \U$41383 ( \41636 , \27447 );
buf \U$41384 ( \41637 , \27440 );
not \U$41385 ( \41638 , \41637 );
not \U$41386 ( \41639 , \25624 );
not \U$41387 ( \41640 , \27430 );
not \U$41388 ( \41641 , \27157 );
not \U$41389 ( \41642 , \41641 );
not \U$41390 ( \41643 , \20403 );
or \U$41391 ( \41644 , \41642 , \41643 );
nor \U$41392 ( \41645 , \31536 , \27435 );
nand \U$41393 ( \41646 , \41644 , \41645 );
not \U$41394 ( \41647 , \41646 );
or \U$41395 ( \41648 , \41640 , \41647 );
not \U$41396 ( \41649 , \31507 );
nand \U$41397 ( \41650 , \41648 , \41649 );
not \U$41398 ( \41651 , \41650 );
or \U$41399 ( \41652 , \41639 , \41651 );
not \U$41400 ( \41653 , \27438 );
nand \U$41401 ( \41654 , \41652 , \41653 );
not \U$41402 ( \41655 , \41654 );
or \U$41403 ( \41656 , \41638 , \41655 );
nand \U$41404 ( \41657 , \41656 , \27443 );
not \U$41405 ( \41658 , \41657 );
or \U$41406 ( \41659 , \41636 , \41658 );
not \U$41407 ( \41660 , \27450 );
nand \U$41408 ( \41661 , \41659 , \41660 );
buf \U$41409 ( \41662 , \27448 );
xor \U$41410 ( \41663 , \41661 , \41662 );
not \U$41411 ( \41664 , \32075 );
not \U$41412 ( \41665 , \31545 );
not \U$41413 ( \41666 , \27461 );
buf \U$41414 ( \41667 , \27436 );
nand \U$41415 ( \41668 , \41665 , \41666 , \27431 , \41667 );
not \U$41416 ( \41669 , \41668 );
or \U$41417 ( \41670 , \41664 , \41669 );
not \U$41418 ( \41671 , \32086 );
nand \U$41419 ( \41672 , \41670 , \41671 );
buf \U$41420 ( \41673 , \32029 );
xor \U$41421 ( \41674 , \41672 , \41673 );
xor \U$41422 ( \41675 , \41657 , \27447 );
xor \U$41423 ( \41676 , \41668 , \32075 );
and \U$41424 ( \41677 , \41674 , \41675 , \41676 );
nand \U$41425 ( \41678 , \41663 , \41677 );
not \U$41426 ( \41679 , \41678 );
not \U$41427 ( \41680 , \39637 );
not \U$41428 ( \41681 , \40787 );
not \U$41429 ( \41682 , \32121 );
or \U$41430 ( \41683 , \41681 , \41682 );
not \U$41431 ( \41684 , \40796 );
nand \U$41432 ( \41685 , \41683 , \41684 );
not \U$41433 ( \41686 , \41685 );
or \U$41434 ( \41687 , \41680 , \41686 );
nand \U$41435 ( \41688 , \41687 , \40800 );
and \U$41436 ( \41689 , \41688 , \39614 );
nor \U$41437 ( \41690 , \41689 , \40805 );
buf \U$41438 ( \41691 , \39583 );
xnor \U$41439 ( \41692 , \41690 , \41691 );
nand \U$41440 ( \41693 , \41679 , \41692 );
and \U$41441 ( \41694 , \41688 , \39613 );
not \U$41442 ( \41695 , \41688 );
and \U$41443 ( \41696 , \41695 , \39614 );
nor \U$41444 ( \41697 , \41694 , \41696 );
not \U$41445 ( \41698 , \41697 );
xor \U$41446 ( \41699 , \41685 , \39637 );
buf \U$41447 ( \41700 , \41374 );
xor \U$41448 ( \41701 , \41700 , \40724 );
and \U$41449 ( \41702 , \41699 , \41701 );
buf \U$41450 ( \41703 , \41378 );
and \U$41451 ( \41704 , \41703 , \41366 );
not \U$41452 ( \41705 , \41703 );
and \U$41453 ( \41706 , \41705 , \38808 );
nor \U$41454 ( \41707 , \41704 , \41706 );
not \U$41455 ( \41708 , \15749 );
not \U$41456 ( \41709 , \15380 );
buf \U$41457 ( \41710 , \15762 );
not \U$41458 ( \41711 , \41710 );
not \U$41459 ( \41712 , \14450 );
not \U$41460 ( \41713 , \19509 );
not \U$41461 ( \41714 , \41713 );
not \U$41462 ( \41715 , \19517 );
not \U$41463 ( \41716 , \20400 );
or \U$41464 ( \41717 , \41715 , \41716 );
not \U$41465 ( \41718 , \19498 );
nand \U$41466 ( \41719 , \41717 , \41718 );
and \U$41467 ( \41720 , \19500 , \19502 );
nand \U$41468 ( \41721 , \41719 , \41720 );
buf \U$41469 ( \41722 , \18128 );
nand \U$41470 ( \41723 , \41721 , \41722 , \19504 );
not \U$41471 ( \41724 , \41723 );
or \U$41472 ( \41725 , \41714 , \41724 );
not \U$41473 ( \41726 , \14717 );
nand \U$41474 ( \41727 , \41725 , \41726 );
not \U$41475 ( \41728 , \41727 );
or \U$41476 ( \41729 , \41712 , \41728 );
not \U$41477 ( \41730 , \14719 );
nand \U$41478 ( \41731 , \41729 , \41730 );
not \U$41479 ( \41732 , \41731 );
or \U$41480 ( \41733 , \41711 , \41732 );
nand \U$41481 ( \41734 , \41733 , \15765 );
not \U$41482 ( \41735 , \41734 );
or \U$41483 ( \41736 , \41709 , \41735 );
not \U$41484 ( \41737 , \15768 );
nand \U$41485 ( \41738 , \41736 , \41737 );
not \U$41486 ( \41739 , \41738 );
or \U$41487 ( \41740 , \41708 , \41739 );
not \U$41488 ( \41741 , \16924 );
nand \U$41489 ( \41742 , \41740 , \41741 );
buf \U$41490 ( \41743 , \16919 );
and \U$41491 ( \41744 , \41742 , \41743 );
not \U$41492 ( \41745 , \16930 );
nor \U$41493 ( \41746 , \41744 , \41745 );
buf \U$41494 ( \41747 , \16903 );
not \U$41495 ( \41748 , \41747 );
and \U$41496 ( \41749 , \41746 , \41748 );
not \U$41497 ( \41750 , \41746 );
and \U$41498 ( \41751 , \41750 , \41747 );
nor \U$41499 ( \41752 , \41749 , \41751 );
not \U$41500 ( \41753 , \41752 );
not \U$41501 ( \41754 , \18104 );
not \U$41502 ( \41755 , \18099 );
not \U$41503 ( \41756 , \19501 );
not \U$41504 ( \41757 , \41719 );
or \U$41505 ( \41758 , \41756 , \41757 );
not \U$41506 ( \41759 , \18088 );
nand \U$41507 ( \41760 , \41758 , \41759 );
not \U$41508 ( \41761 , \41760 );
or \U$41509 ( \41762 , \41755 , \41761 );
nand \U$41510 ( \41763 , \41762 , \18102 );
not \U$41511 ( \41764 , \41763 );
or \U$41512 ( \41765 , \41754 , \41764 );
not \U$41513 ( \41766 , \17869 );
nand \U$41514 ( \41767 , \41765 , \41766 );
buf \U$41515 ( \41768 , \17656 );
xnor \U$41516 ( \41769 , \41767 , \41768 );
not \U$41517 ( \41770 , \41769 );
xnor \U$41518 ( \41771 , \41763 , \18104 );
not \U$41519 ( \41772 , \41771 );
buf \U$41520 ( \41773 , \17441 );
and \U$41521 ( \41774 , \41767 , \41768 );
nor \U$41522 ( \41775 , \41774 , \17871 );
xnor \U$41523 ( \41776 , \41773 , \41775 );
not \U$41524 ( \41777 , \18106 );
and \U$41525 ( \41778 , \19500 , \19501 );
nand \U$41526 ( \41779 , \41719 , \41778 );
nand \U$41527 ( \41780 , \41777 , \41779 );
xor \U$41528 ( \41781 , \41780 , \18127 );
nand \U$41529 ( \41782 , \41770 , \41772 , \41776 , \41781 );
nor \U$41530 ( \41783 , \41753 , \41782 );
nand \U$41531 ( \41784 , \41698 , \41702 , \41707 , \41783 );
nor \U$41532 ( \41785 , \41693 , \41784 );
and \U$41533 ( \41786 , \41661 , \41662 );
not \U$41534 ( \41787 , \27455 );
nor \U$41535 ( \41788 , \41786 , \41787 );
not \U$41536 ( \41789 , \41788 );
not \U$41537 ( \41790 , \27446 );
and \U$41538 ( \41791 , \41789 , \41790 );
and \U$41539 ( \41792 , \41788 , \27446 );
nor \U$41540 ( \41793 , \41791 , \41792 );
not \U$41541 ( \41794 , \41793 );
not \U$41542 ( \41795 , \41742 );
not \U$41543 ( \41796 , \41795 );
not \U$41544 ( \41797 , \41743 );
and \U$41545 ( \41798 , \41796 , \41797 );
and \U$41546 ( \41799 , \41795 , \41743 );
nor \U$41547 ( \41800 , \41798 , \41799 );
not \U$41548 ( \41801 , \41800 );
and \U$41549 ( \41802 , \19506 , \19507 );
not \U$41550 ( \41803 , \41802 );
buf \U$41551 ( \41804 , \41731 );
not \U$41552 ( \41805 , \41804 );
or \U$41553 ( \41806 , \41803 , \41805 );
not \U$41554 ( \41807 , \15769 );
and \U$41555 ( \41808 , \19506 , \41807 );
not \U$41556 ( \41809 , \15767 );
and \U$41557 ( \41810 , \19506 , \41809 );
nor \U$41558 ( \41811 , \41808 , \41810 , \16935 );
nand \U$41559 ( \41812 , \41806 , \41811 );
xor \U$41560 ( \41813 , \41812 , \16936 );
buf \U$41561 ( \41814 , \20403 );
buf \U$41562 ( \41815 , \27155 );
xor \U$41563 ( \41816 , \41814 , \41815 );
buf \U$41564 ( \41817 , \41727 );
and \U$41565 ( \41818 , \41817 , \14450 );
not \U$41566 ( \41819 , \41817 );
and \U$41567 ( \41820 , \41819 , \19510 );
nor \U$41568 ( \41821 , \41818 , \41820 );
not \U$41569 ( \41822 , \41713 );
and \U$41570 ( \41823 , \41780 , \18127 );
not \U$41571 ( \41824 , \19504 );
nor \U$41572 ( \41825 , \41823 , \41824 );
not \U$41573 ( \41826 , \41825 );
or \U$41574 ( \41827 , \41822 , \41826 );
or \U$41575 ( \41828 , \41713 , \41825 );
nand \U$41576 ( \41829 , \41827 , \41828 );
nand \U$41577 ( \41830 , \41816 , \41821 , \41829 );
xnor \U$41578 ( \41831 , \41804 , \41710 );
nor \U$41579 ( \41832 , \41830 , \41831 );
nand \U$41580 ( \41833 , \41813 , \41832 );
buf \U$41581 ( \41834 , \41734 );
not \U$41582 ( \41835 , \41834 );
not \U$41583 ( \41836 , \15380 );
not \U$41584 ( \41837 , \41836 );
and \U$41585 ( \41838 , \41835 , \41837 );
and \U$41586 ( \41839 , \41834 , \41836 );
nor \U$41587 ( \41840 , \41838 , \41839 );
nor \U$41588 ( \41841 , \41833 , \41840 );
not \U$41589 ( \41842 , \15749 );
not \U$41590 ( \41843 , \41738 );
not \U$41591 ( \41844 , \41843 );
or \U$41592 ( \41845 , \41842 , \41844 );
or \U$41593 ( \41846 , \41843 , \15749 );
nand \U$41594 ( \41847 , \41845 , \41846 );
nand \U$41595 ( \41848 , \41841 , \41847 );
not \U$41596 ( \41849 , \41848 );
buf \U$41597 ( \41850 , \19467 );
buf \U$41598 ( \41851 , \19451 );
not \U$41599 ( \41852 , \41851 );
not \U$41600 ( \41853 , \19375 );
not \U$41601 ( \41854 , \19516 );
not \U$41602 ( \41855 , \20400 );
or \U$41603 ( \41856 , \41854 , \41855 );
nand \U$41604 ( \41857 , \41856 , \19303 );
not \U$41605 ( \41858 , \41857 );
or \U$41606 ( \41859 , \41853 , \41858 );
nand \U$41607 ( \41860 , \41859 , \19377 );
not \U$41608 ( \41861 , \41860 );
or \U$41609 ( \41862 , \41852 , \41861 );
nand \U$41610 ( \41863 , \41862 , \19472 );
xor \U$41611 ( \41864 , \41850 , \41863 );
not \U$41612 ( \41865 , \18849 );
not \U$41613 ( \41866 , \19481 );
nand \U$41614 ( \41867 , \20400 , \19515 , \19516 );
nand \U$41615 ( \41868 , \41866 , \41867 );
not \U$41616 ( \41869 , \41868 );
or \U$41617 ( \41870 , \41865 , \41869 );
not \U$41618 ( \41871 , \19487 );
nand \U$41619 ( \41872 , \41870 , \41871 );
buf \U$41620 ( \41873 , \18690 );
and \U$41621 ( \41874 , \41872 , \41873 );
not \U$41622 ( \41875 , \41872 );
not \U$41623 ( \41876 , \41873 );
and \U$41624 ( \41877 , \41875 , \41876 );
nor \U$41625 ( \41878 , \41874 , \41877 );
xnor \U$41626 ( \41879 , \41868 , \18849 );
xnor \U$41627 ( \41880 , \41719 , \19501 );
nor \U$41628 ( \41881 , \41879 , \41880 );
and \U$41629 ( \41882 , \41878 , \41881 );
and \U$41630 ( \41883 , \41864 , \41882 );
not \U$41631 ( \41884 , \41850 );
not \U$41632 ( \41885 , \41863 );
or \U$41633 ( \41886 , \41884 , \41885 );
nand \U$41634 ( \41887 , \41886 , \19475 );
buf \U$41635 ( \41888 , \19514 );
and \U$41636 ( \41889 , \41887 , \41888 );
not \U$41637 ( \41890 , \41887 );
not \U$41638 ( \41891 , \41888 );
and \U$41639 ( \41892 , \41890 , \41891 );
nor \U$41640 ( \41893 , \41889 , \41892 );
not \U$41641 ( \41894 , \41873 );
not \U$41642 ( \41895 , \41872 );
or \U$41643 ( \41896 , \41894 , \41895 );
not \U$41644 ( \41897 , \19489 );
nand \U$41645 ( \41898 , \41896 , \41897 );
xor \U$41646 ( \41899 , \18513 , \41898 );
and \U$41647 ( \41900 , \41883 , \41893 , \41899 );
not \U$41648 ( \41901 , \18513 );
not \U$41649 ( \41902 , \41898 );
or \U$41650 ( \41903 , \41901 , \41902 );
nand \U$41651 ( \41904 , \41903 , \19494 );
buf \U$41652 ( \41905 , \18520 );
xor \U$41653 ( \41906 , \41904 , \41905 );
and \U$41654 ( \41907 , \20371 , \20018 );
not \U$41655 ( \41908 , \41907 );
not \U$41656 ( \41909 , \20371 );
not \U$41657 ( \41910 , \20018 );
and \U$41658 ( \41911 , \41909 , \41910 );
or \U$41659 ( \41912 , \20368 , \20369 );
not \U$41660 ( \41913 , \20360 );
not \U$41661 ( \41914 , \20354 );
nand \U$41662 ( \41915 , \41914 , \20325 );
nand \U$41663 ( \41916 , \41913 , \41915 );
not \U$41664 ( \41917 , \41916 );
not \U$41665 ( \41918 , \20358 );
and \U$41666 ( \41919 , \41917 , \41918 );
and \U$41667 ( \41920 , \41916 , \20358 );
nor \U$41668 ( \41921 , \41919 , \41920 );
not \U$41669 ( \41922 , \20325 );
and \U$41670 ( \41923 , \41922 , \20354 );
not \U$41671 ( \41924 , \20324 );
or \U$41672 ( \41925 , \20322 , \20323 );
not \U$41673 ( \41926 , \20319 );
not \U$41674 ( \41927 , \20320 );
and \U$41675 ( \41928 , \41926 , \41927 );
not \U$41676 ( \41929 , \20321 );
and \U$41677 ( \41930 , \30890 , \20278 );
not \U$41678 ( \41931 , \20279 );
nand \U$41679 ( \41932 , \41931 , \20271 );
_DC gfa ( \41933_nGfa , 1'b0 , 1'b1 );
_DC gf9 ( \41934_nGf9 , 1'b0 , 1'b1 );
nand \U$41684 ( \41935 , \41933_nGfa , \41934_nGf9 );
nor \U$41685 ( \41936 , \41930 , \41932 , \41935 );
nand \U$41686 ( \41937 , \20315 , \41936 , \20267 , \20302 );
nor \U$41687 ( \41938 , \41928 , \41929 , \41937 );
nand \U$41688 ( \41939 , \41925 , \41938 );
nor \U$41689 ( \41940 , \41923 , \41924 , \41939 );
nand \U$41690 ( \41941 , \41921 , \41915 , \20006 , \41940 );
or \U$41691 ( \41942 , \20365 , \20366 );
nand \U$41692 ( \41943 , \41942 , \20367 );
nor \U$41693 ( \41944 , \41941 , \41943 );
nand \U$41694 ( \41945 , \41912 , \41944 , \20370 );
nor \U$41695 ( \41946 , \41911 , \41945 );
nand \U$41696 ( \41947 , \41908 , \41946 );
not \U$41697 ( \41948 , \41947 );
not \U$41698 ( \41949 , \20006 );
not \U$41699 ( \41950 , \41907 );
or \U$41700 ( \41951 , \41949 , \41950 );
nand \U$41701 ( \41952 , \41951 , \20384 );
and \U$41702 ( \41953 , \41952 , \19911 );
not \U$41703 ( \41954 , \41952 );
and \U$41704 ( \41955 , \41954 , \19910 );
nor \U$41705 ( \41956 , \41953 , \41955 );
nand \U$41706 ( \41957 , \41948 , \41956 );
not \U$41707 ( \41958 , \19911 );
not \U$41708 ( \41959 , \41952 );
or \U$41709 ( \41960 , \41958 , \41959 );
nand \U$41710 ( \41961 , \41960 , \20387 );
xnor \U$41711 ( \41962 , \41961 , \20050 );
nor \U$41712 ( \41963 , \41957 , \41962 );
not \U$41713 ( \41964 , \20050 );
not \U$41714 ( \41965 , \41961 );
or \U$41715 ( \41966 , \41964 , \41965 );
nand \U$41716 ( \41967 , \41966 , \20391 );
xor \U$41717 ( \41968 , \41967 , \20034 );
and \U$41718 ( \41969 , \41963 , \41968 );
xor \U$41719 ( \41970 , \20395 , \19623 );
nand \U$41720 ( \41971 , \41969 , \41970 );
xnor \U$41721 ( \41972 , \20400 , \19516 );
nor \U$41722 ( \41973 , \41971 , \41972 );
xor \U$41723 ( \41974 , \41857 , \19375 );
nand \U$41724 ( \41975 , \41973 , \41974 );
xnor \U$41725 ( \41976 , \41860 , \41851 );
nor \U$41726 ( \41977 , \41975 , \41976 );
nand \U$41727 ( \41978 , \41900 , \41906 , \41977 );
xnor \U$41728 ( \41979 , \41760 , \18099 );
nor \U$41729 ( \41980 , \41978 , \41979 );
and \U$41730 ( \41981 , \41801 , \41849 , \41980 );
nand \U$41731 ( \41982 , \41794 , \41981 );
not \U$41732 ( \41983 , \32067 );
buf \U$41733 ( \41984 , \32030 );
not \U$41734 ( \41985 , \41984 );
not \U$41735 ( \41986 , \41985 );
and \U$41736 ( \41987 , \41668 , \32075 );
not \U$41737 ( \41988 , \41987 );
or \U$41738 ( \41989 , \41986 , \41988 );
not \U$41739 ( \41990 , \32097 );
nand \U$41740 ( \41991 , \41990 , \32116 );
nand \U$41741 ( \41992 , \41989 , \41991 );
not \U$41742 ( \41993 , \41992 );
or \U$41743 ( \41994 , \41983 , \41993 );
nand \U$41744 ( \41995 , \41994 , \32099 );
xnor \U$41745 ( \41996 , \41995 , \32059 );
xor \U$41746 ( \41997 , \41992 , \32067 );
xor \U$41747 ( \41998 , \32121 , \40787 );
not \U$41748 ( \41999 , \32081 );
nor \U$41749 ( \42000 , \41984 , \32076 );
not \U$41750 ( \42001 , \42000 );
not \U$41751 ( \42002 , \41668 );
or \U$41752 ( \42003 , \42001 , \42002 );
not \U$41753 ( \42004 , \32104 );
nand \U$41754 ( \42005 , \42004 , \32119 , \32102 );
nand \U$41755 ( \42006 , \42003 , \42005 );
not \U$41756 ( \42007 , \42006 );
or \U$41757 ( \42008 , \41999 , \42007 );
or \U$41758 ( \42009 , \42006 , \32081 );
nand \U$41759 ( \42010 , \42008 , \42009 );
not \U$41760 ( \42011 , \27147 );
not \U$41761 ( \42012 , \41815 );
not \U$41762 ( \42013 , \20403 );
or \U$41763 ( \42014 , \42012 , \42013 );
not \U$41764 ( \42015 , \31511 );
nand \U$41765 ( \42016 , \42014 , \42015 );
not \U$41766 ( \42017 , \42016 );
or \U$41767 ( \42018 , \42011 , \42017 );
nand \U$41768 ( \42019 , \42018 , \31515 );
not \U$41769 ( \42020 , \42019 );
not \U$41770 ( \42021 , \42020 );
not \U$41771 ( \42022 , \27117 );
and \U$41772 ( \42023 , \42021 , \42022 );
and \U$41773 ( \42024 , \42020 , \27117 );
nor \U$41774 ( \42025 , \42023 , \42024 );
buf \U$41775 ( \42026 , \42016 );
xnor \U$41776 ( \42027 , \27147 , \42026 );
nor \U$41777 ( \42028 , \42025 , \42027 );
and \U$41778 ( \42029 , \41998 , \42010 , \42028 );
not \U$41779 ( \42030 , \31915 );
not \U$41780 ( \42031 , \42030 );
and \U$41781 ( \42032 , \41673 , \32075 );
not \U$41782 ( \42033 , \42032 );
not \U$41783 ( \42034 , \41668 );
or \U$41784 ( \42035 , \42033 , \42034 );
and \U$41785 ( \42036 , \32087 , \32089 );
nand \U$41786 ( \42037 , \42035 , \42036 );
not \U$41787 ( \42038 , \42037 );
or \U$41788 ( \42039 , \42031 , \42038 );
or \U$41789 ( \42040 , \42037 , \42030 );
nand \U$41790 ( \42041 , \42039 , \42040 );
nand \U$41791 ( \42042 , \41997 , \42029 , \42041 );
nor \U$41792 ( \42043 , \41996 , \42042 );
buf \U$41793 ( \42044 , \27385 );
not \U$41794 ( \42045 , \42044 );
not \U$41795 ( \42046 , \31538 );
buf \U$41796 ( \42047 , \27429 );
not \U$41797 ( \42048 , \42047 );
not \U$41798 ( \42049 , \41646 );
or \U$41799 ( \42050 , \42048 , \42049 );
not \U$41800 ( \42051 , \31476 );
nand \U$41801 ( \42052 , \42050 , \42051 );
not \U$41802 ( \42053 , \42052 );
or \U$41803 ( \42054 , \42046 , \42053 );
not \U$41804 ( \42055 , \31488 );
nand \U$41805 ( \42056 , \42054 , \42055 );
not \U$41806 ( \42057 , \42056 );
or \U$41807 ( \42058 , \42045 , \42057 );
nand \U$41808 ( \42059 , \42058 , \31492 );
not \U$41809 ( \42060 , \42059 );
not \U$41810 ( \42061 , \31485 );
or \U$41811 ( \42062 , \42060 , \42061 );
not \U$41812 ( \42063 , \31502 );
nand \U$41813 ( \42064 , \42062 , \42063 );
not \U$41814 ( \42065 , \31500 );
xor \U$41815 ( \42066 , \42064 , \42065 );
not \U$41816 ( \42067 , \41654 );
not \U$41817 ( \42068 , \42067 );
not \U$41818 ( \42069 , \41637 );
and \U$41819 ( \42070 , \42068 , \42069 );
and \U$41820 ( \42071 , \42067 , \41637 );
nor \U$41821 ( \42072 , \42070 , \42071 );
buf \U$41822 ( \42073 , \42052 );
xor \U$41823 ( \42074 , \42073 , \31538 );
xor \U$41824 ( \42075 , \41650 , \25624 );
buf \U$41825 ( \42076 , \41646 );
xor \U$41826 ( \42077 , \42076 , \42047 );
nand \U$41827 ( \42078 , \42074 , \42075 , \42077 );
nor \U$41828 ( \42079 , \42072 , \42078 );
buf \U$41829 ( \42080 , \26912 );
not \U$41830 ( \42081 , \42080 );
not \U$41831 ( \42082 , \27117 );
not \U$41832 ( \42083 , \42019 );
or \U$41833 ( \42084 , \42082 , \42083 );
not \U$41834 ( \42085 , \31525 );
nand \U$41835 ( \42086 , \42084 , \42085 );
not \U$41836 ( \42087 , \42086 );
or \U$41837 ( \42088 , \42081 , \42087 );
nand \U$41838 ( \42089 , \42088 , \31529 );
buf \U$41839 ( \42090 , \27077 );
xor \U$41840 ( \42091 , \42089 , \42090 );
and \U$41841 ( \42092 , \42059 , \31485 );
not \U$41842 ( \42093 , \42059 );
and \U$41843 ( \42094 , \42093 , \31486 );
nor \U$41844 ( \42095 , \42092 , \42094 );
xor \U$41845 ( \42096 , \42080 , \42086 );
xor \U$41846 ( \42097 , \42056 , \42044 );
and \U$41847 ( \42098 , \42096 , \42097 );
nand \U$41848 ( \42099 , \42079 , \42091 , \42095 , \42098 );
nor \U$41849 ( \42100 , \42066 , \42099 );
buf \U$41850 ( \42101 , \31971 );
not \U$41851 ( \42102 , \42101 );
not \U$41852 ( \42103 , \31915 );
not \U$41853 ( \42104 , \42037 );
or \U$41854 ( \42105 , \42103 , \42104 );
not \U$41855 ( \42106 , \32110 );
nand \U$41856 ( \42107 , \42105 , \42106 );
not \U$41857 ( \42108 , \42107 );
or \U$41858 ( \42109 , \42102 , \42108 );
nand \U$41859 ( \42110 , \31966 , \31969 );
nand \U$41860 ( \42111 , \42109 , \42110 );
not \U$41861 ( \42112 , \32005 );
xnor \U$41862 ( \42113 , \42111 , \42112 );
xor \U$41863 ( \42114 , \42101 , \42107 );
nand \U$41864 ( \42115 , \42043 , \42100 , \42113 , \42114 );
nor \U$41865 ( \42116 , \41982 , \42115 );
not \U$41866 ( \42117 , \40807 );
not \U$41867 ( \42118 , \42117 );
not \U$41868 ( \42119 , \42118 );
not \U$41869 ( \42120 , \41691 );
not \U$41870 ( \42121 , \41690 );
not \U$41871 ( \42122 , \42121 );
or \U$41872 ( \42123 , \42120 , \42122 );
nand \U$41873 ( \42124 , \42123 , \40810 );
not \U$41874 ( \42125 , \42124 );
or \U$41875 ( \42126 , \42119 , \42125 );
and \U$41876 ( \42127 , \42121 , \41691 );
nand \U$41877 ( \42128 , \42117 , \40810 );
nor \U$41878 ( \42129 , \42127 , \42128 );
not \U$41879 ( \42130 , \42129 );
nand \U$41880 ( \42131 , \42126 , \42130 );
nand \U$41881 ( \42132 , \41785 , \42116 , \42131 );
not \U$41882 ( \42133 , \42132 );
xor \U$41883 ( \42134 , \38570 , \41382 );
buf \U$41884 ( \42135 , \42134 );
nand \U$41885 ( \42136 , \42133 , \42135 );
buf \U$41886 ( \42137 , \42136 );
not \U$41887 ( \42138 , \42137 );
and \U$41888 ( \42139 , \41114 , \2729 );
not \U$41889 ( \42140 , \41114 );
and \U$41890 ( \42141 , \42140 , \2728 );
nor \U$41891 ( \42142 , \42139 , \42141 );
not \U$41892 ( \42143 , \40906 );
not \U$41893 ( \42144 , \41340 );
or \U$41894 ( \42145 , \42143 , \42144 );
nand \U$41895 ( \42146 , \42145 , \40909 );
not \U$41896 ( \42147 , \40889 );
xor \U$41897 ( \42148 , \42146 , \42147 );
not \U$41898 ( \42149 , \41265 );
not \U$41899 ( \42150 , \9736 );
or \U$41900 ( \42151 , \42149 , \42150 );
nand \U$41901 ( \42152 , \42151 , \40931 );
nand \U$41902 ( \42153 , \42152 , \40920 );
not \U$41903 ( \42154 , \41253 );
not \U$41904 ( \42155 , \41261 );
or \U$41905 ( \42156 , \42154 , \42155 );
not \U$41906 ( \42157 , \40926 );
nand \U$41907 ( \42158 , \42156 , \42157 );
xor \U$41908 ( \42159 , \42158 , \41252 );
and \U$41909 ( \42160 , \41261 , \41254 );
not \U$41910 ( \42161 , \41261 );
and \U$41911 ( \42162 , \42161 , \41253 );
nor \U$41912 ( \42163 , \42160 , \42162 );
nor \U$41913 ( \42164 , \42159 , \42163 );
not \U$41914 ( \42165 , \41217 );
not \U$41915 ( \42166 , \41216 );
or \U$41916 ( \42167 , \42165 , \42166 );
nand \U$41917 ( \42168 , \42167 , \40967 );
not \U$41918 ( \42169 , \42168 );
buf \U$41919 ( \42170 , \12669 );
not \U$41920 ( \42171 , \42170 );
and \U$41921 ( \42172 , \42169 , \42171 );
and \U$41922 ( \42173 , \42168 , \42170 );
nor \U$41923 ( \42174 , \42172 , \42173 );
not \U$41924 ( \42175 , \12688 );
xor \U$41925 ( \42176 , \41455 , \42175 );
nor \U$41926 ( \42177 , \42174 , \42176 );
and \U$41927 ( \42178 , \42153 , \42164 , \42177 );
not \U$41928 ( \42179 , \42152 );
not \U$41929 ( \42180 , \40920 );
and \U$41930 ( \42181 , \42179 , \42180 );
and \U$41931 ( \42182 , \41333 , \41334 );
not \U$41932 ( \42183 , \42182 );
not \U$41933 ( \42184 , \40676 );
or \U$41934 ( \42185 , \42183 , \42184 );
not \U$41935 ( \42186 , \40909 );
not \U$41936 ( \42187 , \40907 );
or \U$41937 ( \42188 , \42186 , \42187 );
nand \U$41938 ( \42189 , \42188 , \42147 );
and \U$41939 ( \42190 , \42189 , \40887 );
nand \U$41940 ( \42191 , \42185 , \42190 );
buf \U$41941 ( \42192 , \40892 );
not \U$41942 ( \42193 , \42192 );
and \U$41943 ( \42194 , \42191 , \42193 );
not \U$41944 ( \42195 , \42191 );
and \U$41945 ( \42196 , \42195 , \42192 );
nor \U$41946 ( \42197 , \42194 , \42196 );
not \U$41947 ( \42198 , \12555 );
not \U$41948 ( \42199 , \41223 );
not \U$41949 ( \42200 , \42199 );
or \U$41950 ( \42201 , \42198 , \42200 );
not \U$41951 ( \42202 , \42199 );
nand \U$41952 ( \42203 , \42202 , \41194 );
nand \U$41953 ( \42204 , \42201 , \42203 );
nand \U$41954 ( \42205 , \42197 , \42204 );
nor \U$41955 ( \42206 , \42181 , \42205 );
and \U$41956 ( \42207 , \42148 , \42178 , \42206 );
buf \U$41957 ( \42208 , \42207 );
not \U$41958 ( \42209 , \40857 );
nand \U$41959 ( \42210 , \42209 , \41446 );
not \U$41960 ( \42211 , \42210 );
not \U$41961 ( \42212 , \41362 );
and \U$41962 ( \42213 , \42211 , \42212 );
and \U$41963 ( \42214 , \42210 , \41362 );
nor \U$41964 ( \42215 , \42213 , \42214 );
xor \U$41965 ( \42216 , \41386 , \41435 );
not \U$41966 ( \42217 , \6279 );
not \U$41967 ( \42218 , \42217 );
buf \U$41968 ( \42219 , \41239 );
not \U$41969 ( \42220 , \42219 );
or \U$41970 ( \42221 , \42218 , \42220 );
or \U$41971 ( \42222 , \42219 , \42217 );
nand \U$41972 ( \42223 , \42221 , \42222 );
nand \U$41973 ( \42224 , \42216 , \42223 );
nor \U$41974 ( \42225 , \42215 , \42224 );
buf \U$41975 ( \42226 , \42225 );
and \U$41976 ( \42227 , \42142 , \42208 , \42226 );
not \U$41977 ( \42228 , \938 );
and \U$41978 ( \42229 , \41297 , \42228 );
nor \U$41979 ( \42230 , \42229 , \41091 );
xnor \U$41980 ( \42231 , \42230 , \927 );
and \U$41981 ( \42232 , \41498 , \41492 );
not \U$41982 ( \42233 , \41498 );
and \U$41983 ( \42234 , \42233 , \3146 );
nor \U$41984 ( \42235 , \42232 , \42234 );
xnor \U$41985 ( \42236 , \2516 , \41117 );
buf \U$41986 ( \42237 , \42236 );
and \U$41987 ( \42238 , \41481 , \41494 );
not \U$41988 ( \42239 , \41481 );
and \U$41989 ( \42240 , \42239 , \3138 );
nor \U$41990 ( \42241 , \42238 , \42240 );
nand \U$41991 ( \42242 , \42235 , \42237 , \42241 );
not \U$41992 ( \42243 , \41121 );
not \U$41993 ( \42244 , \41120 );
or \U$41994 ( \42245 , \42243 , \42244 );
nand \U$41995 ( \42246 , \42245 , \41050 );
not \U$41996 ( \42247 , \2296 );
and \U$41997 ( \42248 , \42246 , \42247 );
not \U$41998 ( \42249 , \42246 );
and \U$41999 ( \42250 , \42249 , \2296 );
or \U$42000 ( \42251 , \42248 , \42250 );
nor \U$42001 ( \42252 , \42242 , \42251 );
nand \U$42002 ( \42253 , \42138 , \42227 , \42231 , \42252 );
not \U$42003 ( \42254 , \42253 );
nand \U$42004 ( \42255 , \41567 , \41634 , \41635 , \42254 );
not \U$42005 ( \42256 , \41575 );
not \U$42006 ( \42257 , \342 );
and \U$42007 ( \42258 , \42256 , \42257 );
and \U$42008 ( \42259 , \41575 , \342 );
nor \U$42009 ( \42260 , \42258 , \42259 );
not \U$42010 ( \42261 , \42260 );
nand \U$42011 ( \42262 , RIbe27b98_2, RIbe29380_53);
not \U$42012 ( \42263 , \42262 );
and \U$42013 ( \42264 , \41576 , \41589 );
not \U$42014 ( \42265 , \42264 );
or \U$42015 ( \42266 , \42263 , \42265 );
or \U$42016 ( \42267 , \42264 , \42262 );
nand \U$42017 ( \42268 , \42266 , \42267 );
not \U$42018 ( \42269 , \42268 );
or \U$42019 ( \42270 , \42261 , \42269 );
or \U$42020 ( \42271 , \42268 , \42260 );
nand \U$42021 ( \42272 , \42270 , \42271 );
not \U$42022 ( \42273 , \42272 );
xor \U$42023 ( \42274 , \41590 , \41602 );
and \U$42024 ( \42275 , \42274 , \41633 );
and \U$42025 ( \42276 , \41590 , \41602 );
nor \U$42026 ( \42277 , \42275 , \42276 );
not \U$42027 ( \42278 , \42277 );
or \U$42028 ( \42279 , \42273 , \42278 );
or \U$42029 ( \42280 , \42277 , \42272 );
nand \U$42030 ( \42281 , \42279 , \42280 );
not \U$42031 ( \42282 , \42281 );
and \U$42032 ( \42283 , \42255 , \42282 );
not \U$42033 ( \42284 , \42255 );
and \U$42034 ( \42285 , \42284 , \42281 );
nor \U$42035 ( \42286 , \42283 , \42285 );
buf \U$42036 ( \42287 , \42286 );
nand \U$42037 ( \42288 , \41567 , \41635 , \42254 );
not \U$42038 ( \42289 , \41634 );
and \U$42039 ( \42290 , \42288 , \42289 );
not \U$42040 ( \42291 , \42288 );
and \U$42041 ( \42292 , \42291 , \41634 );
nor \U$42042 ( \42293 , \42290 , \42292 );
buf \U$42043 ( \42294 , \42293 );
not \U$42044 ( \42295 , \41125 );
and \U$42045 ( \42296 , \41556 , \41515 , \42295 );
nor \U$42046 ( \42297 , \41564 , \41104 );
and \U$42047 ( \42298 , \41292 , \41301 );
nand \U$42048 ( \42299 , \42296 , \42297 , \42298 , \41503 );
not \U$42049 ( \42300 , \42299 );
buf \U$42050 ( \42301 , \41187 );
not \U$42051 ( \42302 , \42253 );
and \U$42052 ( \42303 , \42300 , \42301 , \41100 , \42302 );
and \U$42053 ( \42304 , \42303 , \41635 );
not \U$42054 ( \42305 , \42303 );
not \U$42055 ( \42306 , \41635 );
and \U$42056 ( \42307 , \42305 , \42306 );
nor \U$42057 ( \42308 , \42304 , \42307 );
buf \U$42058 ( \42309 , \42308 );
not \U$42059 ( \42310 , \42253 );
nand \U$42060 ( \42311 , \42310 , \42300 , \41100 );
not \U$42061 ( \42312 , \42301 );
and \U$42062 ( \42313 , \42311 , \42312 );
not \U$42063 ( \42314 , \42311 );
and \U$42064 ( \42315 , \42314 , \42301 );
nor \U$42065 ( \42316 , \42313 , \42315 );
buf \U$42066 ( \42317 , \42316 );
nor \U$42067 ( \42318 , \42299 , \42253 );
not \U$42068 ( \42319 , \42318 );
not \U$42069 ( \42320 , \41100 );
not \U$42070 ( \42321 , \42320 );
or \U$42071 ( \42322 , \42319 , \42321 );
or \U$42072 ( \42323 , \42320 , \42318 );
nand \U$42073 ( \42324 , \42322 , \42323 );
buf \U$42074 ( \42325 , \42324 );
not \U$42075 ( \42326 , \42132 );
nand \U$42076 ( \42327 , \41283 , \41281 );
nand \U$42077 ( \42328 , \42326 , \42327 );
not \U$42078 ( \42329 , \42328 );
and \U$42079 ( \42330 , \41272 , \41279 , \41290 );
and \U$42080 ( \42331 , \42241 , \42236 , \42135 );
and \U$42081 ( \42332 , \42331 , \42235 );
and \U$42082 ( \42333 , \42246 , \42247 );
not \U$42083 ( \42334 , \42246 );
and \U$42084 ( \42335 , \42334 , \2296 );
nor \U$42085 ( \42336 , \42333 , \42335 );
nand \U$42086 ( \42337 , \42329 , \42330 , \42332 , \42336 );
not \U$42087 ( \42338 , \42337 );
and \U$42088 ( \42339 , \42142 , \40986 );
nand \U$42089 ( \42340 , \41543 , \41555 , \42339 );
not \U$42090 ( \42341 , \42340 );
and \U$42091 ( \42342 , \42142 , \5339 );
nand \U$42092 ( \42343 , \41543 , \41555 , \42342 );
not \U$42093 ( \42344 , \42343 );
or \U$42094 ( \42345 , \42341 , \42344 );
nand \U$42095 ( \42346 , \41513 , \41548 );
nand \U$42096 ( \42347 , \42340 , \42346 );
nand \U$42097 ( \42348 , \42345 , \42347 );
nand \U$42098 ( \42349 , \41510 , \41548 );
not \U$42099 ( \42350 , \42349 );
not \U$42100 ( \42351 , \42343 );
or \U$42101 ( \42352 , \42350 , \42351 );
nand \U$42102 ( \42353 , \42352 , \41491 );
nor \U$42103 ( \42354 , \42348 , \42353 );
nand \U$42104 ( \42355 , \41475 , \41502 , \42295 );
nand \U$42105 ( \42356 , \42208 , \42226 );
nor \U$42106 ( \42357 , \42355 , \42356 );
nand \U$42107 ( \42358 , \42349 , \42346 );
nand \U$42108 ( \42359 , \42338 , \42354 , \42357 , \42358 );
not \U$42109 ( \42360 , \42359 );
not \U$42110 ( \42361 , \41565 );
not \U$42111 ( \42362 , \42361 );
not \U$42112 ( \42363 , \41301 );
nor \U$42113 ( \42364 , \41104 , \42363 );
nand \U$42114 ( \42365 , \42360 , \42362 , \42364 );
buf \U$42115 ( \42366 , \42231 );
not \U$42116 ( \42367 , \42366 );
and \U$42117 ( \42368 , \42365 , \42367 );
not \U$42118 ( \42369 , \42365 );
and \U$42119 ( \42370 , \42369 , \42366 );
nor \U$42120 ( \42371 , \42368 , \42370 );
buf \U$42121 ( \42372 , \42371 );
not \U$42122 ( \42373 , \42359 );
buf \U$42123 ( \42374 , \42297 );
nand \U$42124 ( \42375 , \42373 , \42374 );
and \U$42125 ( \42376 , \42375 , \42363 );
not \U$42126 ( \42377 , \42375 );
and \U$42127 ( \42378 , \42377 , \41301 );
nor \U$42128 ( \42379 , \42376 , \42378 );
buf \U$42129 ( \42380 , \42379 );
not \U$42130 ( \42381 , \42337 );
nand \U$42131 ( \42382 , \42381 , \42357 , \42358 );
not \U$42132 ( \42383 , \42382 );
buf \U$42133 ( \42384 , \42354 );
nand \U$42134 ( \42385 , \42383 , \42384 , \42362 , \41103 );
not \U$42135 ( \42386 , \41101 );
and \U$42136 ( \42387 , \42385 , \42386 );
not \U$42137 ( \42388 , \42385 );
and \U$42138 ( \42389 , \42388 , \41101 );
nor \U$42139 ( \42390 , \42387 , \42389 );
buf \U$42140 ( \42391 , \42390 );
not \U$42141 ( \42392 , \42359 );
nand \U$42142 ( \42393 , \42392 , \42362 );
not \U$42143 ( \42394 , \41103 );
and \U$42144 ( \42395 , \42393 , \42394 );
not \U$42145 ( \42396 , \42393 );
and \U$42146 ( \42397 , \42396 , \41103 );
nor \U$42147 ( \42398 , \42395 , \42397 );
buf \U$42148 ( \42399 , \42398 );
buf \U$42149 ( \42400 , \42359 );
and \U$42150 ( \42401 , \42400 , \42361 );
not \U$42151 ( \42402 , \42400 );
and \U$42152 ( \42403 , \42402 , \42362 );
nor \U$42153 ( \42404 , \42401 , \42403 );
buf \U$42154 ( \42405 , \42404 );
not \U$42155 ( \42406 , \42348 );
not \U$42156 ( \42407 , \42357 );
not \U$42157 ( \42408 , \42343 );
not \U$42158 ( \42409 , \42349 );
nor \U$42159 ( \42410 , \42408 , \42409 );
nor \U$42160 ( \42411 , \42407 , \42410 );
not \U$42161 ( \42412 , \42358 );
nor \U$42162 ( \42413 , \42412 , \42337 );
nand \U$42163 ( \42414 , \42406 , \42411 , \42413 );
not \U$42164 ( \42415 , \41491 );
and \U$42165 ( \42416 , \42414 , \42415 );
not \U$42166 ( \42417 , \42414 );
not \U$42167 ( \42418 , \42415 );
and \U$42168 ( \42419 , \42417 , \42418 );
nor \U$42169 ( \42420 , \42416 , \42419 );
buf \U$42170 ( \42421 , \42420 );
not \U$42171 ( \42422 , \42337 );
and \U$42172 ( \42423 , \41475 , \42208 , \42226 );
buf \U$42173 ( \42424 , \42423 );
not \U$42174 ( \42425 , \42340 );
nand \U$42175 ( \42426 , \42425 , \42409 , \42295 );
not \U$42176 ( \42427 , \42346 );
nand \U$42177 ( \42428 , \42427 , \42408 , \42295 );
nand \U$42178 ( \42429 , \42426 , \42428 );
nand \U$42179 ( \42430 , \42422 , \42424 , \42429 );
not \U$42180 ( \42431 , \41502 );
and \U$42181 ( \42432 , \42430 , \42431 );
not \U$42182 ( \42433 , \42430 );
not \U$42183 ( \42434 , \42431 );
and \U$42184 ( \42435 , \42433 , \42434 );
nor \U$42185 ( \42436 , \42432 , \42435 );
buf \U$42186 ( \42437 , \42436 );
buf \U$42187 ( \42438 , \41251 );
not \U$42188 ( \42439 , \41281 );
not \U$42189 ( \42440 , \41278 );
or \U$42190 ( \42441 , \42439 , \42440 );
nand \U$42191 ( \42442 , \41277 , \40955 , \12026 );
nand \U$42192 ( \42443 , \42441 , \42442 );
not \U$42193 ( \42444 , \41290 );
nand \U$42194 ( \42445 , \41208 , \41230 , \41271 );
nor \U$42195 ( \42446 , \42444 , \42445 );
nand \U$42196 ( \42447 , \42443 , \42446 );
nor \U$42197 ( \42448 , \42136 , \42447 );
nand \U$42198 ( \42449 , \42423 , \42438 , \42448 );
not \U$42199 ( \42450 , \42449 );
and \U$42200 ( \42451 , \42429 , \42237 );
not \U$42201 ( \42452 , \42241 );
buf \U$42202 ( \42453 , \42251 );
nor \U$42203 ( \42454 , \42452 , \42453 );
nand \U$42204 ( \42455 , \42450 , \42451 , \42454 );
xnor \U$42205 ( \42456 , \42455 , \42235 );
buf \U$42206 ( \42457 , \42456 );
nand \U$42207 ( \42458 , \42423 , \42448 );
not \U$42208 ( \42459 , \42458 );
not \U$42209 ( \42460 , \42453 );
and \U$42210 ( \42461 , \42451 , \42459 , \42460 , \42438 );
and \U$42211 ( \42462 , \42461 , \42241 );
not \U$42212 ( \42463 , \42461 );
not \U$42213 ( \42464 , \42241 );
and \U$42214 ( \42465 , \42463 , \42464 );
nor \U$42215 ( \42466 , \42462 , \42465 );
buf \U$42216 ( \42467 , \42466 );
nand \U$42217 ( \42468 , \42451 , \42448 , \42438 , \42424 );
and \U$42218 ( \42469 , \42468 , \42453 );
not \U$42219 ( \42470 , \42468 );
and \U$42220 ( \42471 , \42470 , \42460 );
nor \U$42221 ( \42472 , \42469 , \42471 );
buf \U$42222 ( \42473 , \42472 );
not \U$42223 ( \42474 , \42136 );
and \U$42224 ( \42475 , \41474 , \42225 , \42207 , \41555 );
nand \U$42225 ( \42476 , \42474 , \42475 , \41292 );
not \U$42226 ( \42477 , \42476 );
and \U$42227 ( \42478 , \41548 , \41543 , \42142 );
buf \U$42228 ( \42479 , \41515 );
nand \U$42229 ( \42480 , \42477 , \42478 , \42479 , \42237 );
and \U$42230 ( \42481 , \42480 , \41125 );
not \U$42231 ( \42482 , \42480 );
and \U$42232 ( \42483 , \42482 , \42295 );
nor \U$42233 ( \42484 , \42481 , \42483 );
buf \U$42234 ( \42485 , \42484 );
nor \U$42235 ( \42486 , \42136 , \41280 , \41291 );
nand \U$42236 ( \42487 , \41515 , \42475 , \42486 );
buf \U$42237 ( \42488 , \42487 );
not \U$42238 ( \42489 , \42488 );
nand \U$42239 ( \42490 , \42489 , \42478 );
not \U$42240 ( \42491 , \42237 );
and \U$42241 ( \42492 , \42490 , \42491 );
not \U$42242 ( \42493 , \42490 );
and \U$42243 ( \42494 , \42493 , \42237 );
nor \U$42244 ( \42495 , \42492 , \42494 );
buf \U$42245 ( \42496 , \42495 );
not \U$42246 ( \42497 , \41533 );
buf \U$42247 ( \42498 , \42497 );
buf \U$42248 ( \42499 , \41521 );
not \U$42249 ( \42500 , \42499 );
nor \U$42250 ( \42501 , \42487 , \42500 );
nand \U$42251 ( \42502 , \42498 , \42501 );
not \U$42252 ( \42503 , \42502 );
buf \U$42253 ( \42504 , \41527 );
buf \U$42254 ( \42505 , \41522 );
not \U$42255 ( \42506 , \41548 );
buf \U$42256 ( \42507 , \41542 );
not \U$42257 ( \42508 , \42507 );
nor \U$42258 ( \42509 , \42506 , \42508 );
nand \U$42259 ( \42510 , \42503 , \42504 , \42505 , \42509 );
not \U$42260 ( \42511 , \42142 );
and \U$42261 ( \42512 , \42510 , \42511 );
not \U$42262 ( \42513 , \42510 );
and \U$42263 ( \42514 , \42513 , \42142 );
nor \U$42264 ( \42515 , \42512 , \42514 );
buf \U$42265 ( \42516 , \42515 );
nand \U$42266 ( \42517 , \42497 , \42504 );
nor \U$42267 ( \42518 , \42506 , \42508 , \42517 );
and \U$42268 ( \42519 , \42501 , \42518 );
xor \U$42269 ( \42520 , \42505 , \42519 );
buf \U$42270 ( \42521 , \42520 );
nand \U$42271 ( \42522 , \42507 , \42498 , \42504 , \42501 );
and \U$42272 ( \42523 , \42522 , \42506 );
not \U$42273 ( \42524 , \42522 );
and \U$42274 ( \42525 , \42524 , \41548 );
nor \U$42275 ( \42526 , \42523 , \42525 );
buf \U$42276 ( \42527 , \42526 );
nand \U$42277 ( \42528 , \42503 , \42504 );
and \U$42278 ( \42529 , \42528 , \42508 );
not \U$42279 ( \42530 , \42528 );
and \U$42280 ( \42531 , \42530 , \42507 );
nor \U$42281 ( \42532 , \42529 , \42531 );
buf \U$42282 ( \42533 , \42532 );
xnor \U$42283 ( \42534 , \42502 , \42504 );
buf \U$42284 ( \42535 , \42534 );
buf \U$42285 ( \42536 , \42501 );
and \U$42286 ( \42537 , \42536 , \42498 );
not \U$42287 ( \42538 , \42536 );
not \U$42288 ( \42539 , \42498 );
and \U$42289 ( \42540 , \42538 , \42539 );
nor \U$42290 ( \42541 , \42537 , \42540 );
buf \U$42291 ( \42542 , \42541 );
not \U$42292 ( \42543 , \42488 );
not \U$42293 ( \42544 , \42543 );
not \U$42294 ( \42545 , \42500 );
or \U$42295 ( \42546 , \42544 , \42545 );
or \U$42296 ( \42547 , \42500 , \42543 );
nand \U$42297 ( \42548 , \42546 , \42547 );
buf \U$42298 ( \42549 , \42548 );
xnor \U$42299 ( \42550 , \42476 , \42479 );
buf \U$42300 ( \42551 , \42550 );
xnor \U$42301 ( \42552 , \41555 , \42449 );
buf \U$42302 ( \42553 , \42552 );
not \U$42303 ( \42554 , \42438 );
and \U$42304 ( \42555 , \42458 , \42554 );
not \U$42305 ( \42556 , \42458 );
and \U$42306 ( \42557 , \42556 , \42438 );
nor \U$42307 ( \42558 , \42555 , \42557 );
buf \U$42308 ( \42559 , \42558 );
buf \U$42309 ( \42560 , \42215 );
not \U$42310 ( \42561 , \42124 );
not \U$42311 ( \42562 , \42118 );
or \U$42312 ( \42563 , \42561 , \42562 );
nand \U$42313 ( \42564 , \42563 , \42130 );
nand \U$42314 ( \42565 , \41707 , \41702 );
nor \U$42315 ( \42566 , \42565 , \41697 );
and \U$42316 ( \42567 , \42564 , \42566 );
nor \U$42317 ( \42568 , \41413 , \41444 );
not \U$42318 ( \42569 , \41782 );
nand \U$42319 ( \42570 , \42569 , \41692 );
not \U$42320 ( \42571 , \41753 );
nand \U$42321 ( \42572 , \42134 , \42571 , \41981 );
nor \U$42322 ( \42573 , \42570 , \42572 );
nand \U$42323 ( \42574 , \42567 , \42568 , \42573 );
nor \U$42324 ( \42575 , \42560 , \42574 );
buf \U$42325 ( \42576 , \41396 );
buf \U$42326 ( \42577 , \42216 );
and \U$42327 ( \42578 , \42043 , \42100 , \42113 , \42114 );
nor \U$42328 ( \42579 , \41678 , \41793 );
and \U$42329 ( \42580 , \42578 , \42579 );
nand \U$42330 ( \42581 , \42577 , \42580 );
not \U$42331 ( \42582 , \41472 );
nand \U$42332 ( \42583 , \41433 , \42582 , \41446 );
nor \U$42333 ( \42584 , \42581 , \42583 );
nand \U$42334 ( \42585 , \42575 , \42576 , \42584 );
buf \U$42335 ( \42586 , \42585 );
not \U$42336 ( \42587 , \42586 );
and \U$42337 ( \42588 , \41457 , \41450 );
not \U$42338 ( \42589 , \41457 );
and \U$42339 ( \42590 , \42589 , \12696 );
nor \U$42340 ( \42591 , \42588 , \42590 );
and \U$42341 ( \42592 , \42208 , \42446 , \42443 );
nand \U$42342 ( \42593 , \42587 , \42591 , \42223 , \42592 );
not \U$42343 ( \42594 , \41447 );
and \U$42344 ( \42595 , \42593 , \42594 );
not \U$42345 ( \42596 , \42593 );
and \U$42346 ( \42597 , \42596 , \41447 );
nor \U$42347 ( \42598 , \42595 , \42597 );
buf \U$42348 ( \42599 , \42598 );
not \U$42349 ( \42600 , \42447 );
nand \U$42350 ( \42601 , \42600 , \42587 , \42591 , \42208 );
not \U$42351 ( \42602 , \42223 );
and \U$42352 ( \42603 , \42601 , \42602 );
not \U$42353 ( \42604 , \42601 );
and \U$42354 ( \42605 , \42604 , \42223 );
nor \U$42355 ( \42606 , \42603 , \42605 );
buf \U$42356 ( \42607 , \42606 );
nand \U$42357 ( \42608 , \42587 , \42592 );
not \U$42358 ( \42609 , \42591 );
and \U$42359 ( \42610 , \42608 , \42609 );
not \U$42360 ( \42611 , \42608 );
and \U$42361 ( \42612 , \42611 , \42591 );
nor \U$42362 ( \42613 , \42610 , \42612 );
buf \U$42363 ( \42614 , \42613 );
not \U$42364 ( \42615 , \42585 );
buf \U$42365 ( \42616 , \42146 );
xnor \U$42366 ( \42617 , \40889 , \42616 );
not \U$42367 ( \42618 , \42205 );
and \U$42368 ( \42619 , \42617 , \42618 );
nand \U$42369 ( \42620 , \42615 , \42619 );
nor \U$42370 ( \42621 , \42620 , \42163 );
nor \U$42371 ( \42622 , \42159 , \42174 );
buf \U$42372 ( \42623 , \42152 );
xor \U$42373 ( \42624 , \42623 , \40920 );
and \U$42374 ( \42625 , \42443 , \42446 , \42624 );
nand \U$42375 ( \42626 , \42621 , \42622 , \42625 );
buf \U$42376 ( \42627 , \42176 );
and \U$42377 ( \42628 , \42626 , \42627 );
not \U$42378 ( \42629 , \42626 );
not \U$42379 ( \42630 , \42627 );
and \U$42380 ( \42631 , \42629 , \42630 );
nor \U$42381 ( \42632 , \42628 , \42631 );
buf \U$42382 ( \42633 , \42632 );
not \U$42383 ( \42634 , \42620 );
not \U$42384 ( \42635 , \42159 );
not \U$42385 ( \42636 , \42163 );
nand \U$42386 ( \42637 , \42634 , \42625 , \42635 , \42636 );
and \U$42387 ( \42638 , \42637 , \42174 );
not \U$42388 ( \42639 , \42637 );
not \U$42389 ( \42640 , \42174 );
and \U$42390 ( \42641 , \42639 , \42640 );
nor \U$42391 ( \42642 , \42638 , \42641 );
buf \U$42392 ( \42643 , \42642 );
not \U$42393 ( \42644 , \42164 );
not \U$42394 ( \42645 , \41271 );
nor \U$42395 ( \42646 , \42644 , \42645 );
nand \U$42396 ( \42647 , \42617 , \42624 , \42646 , \42618 );
nor \U$42397 ( \42648 , \42585 , \42647 );
buf \U$42398 ( \42649 , \41210 );
and \U$42399 ( \42650 , \42648 , \42649 );
buf \U$42400 ( \42651 , \41208 );
not \U$42401 ( \42652 , \42443 );
buf \U$42402 ( \42653 , \41290 );
not \U$42403 ( \42654 , \41229 );
nand \U$42404 ( \42655 , \42653 , \42654 );
nor \U$42405 ( \42656 , \42652 , \42655 );
and \U$42406 ( \42657 , \42650 , \42651 , \42656 );
and \U$42407 ( \42658 , \42657 , \41221 );
not \U$42408 ( \42659 , \42657 );
not \U$42409 ( \42660 , \41221 );
and \U$42410 ( \42661 , \42659 , \42660 );
nor \U$42411 ( \42662 , \42658 , \42661 );
buf \U$42412 ( \42663 , \42662 );
nand \U$42413 ( \42664 , \42650 , \42653 , \42651 , \42443 );
not \U$42414 ( \42665 , \42654 );
and \U$42415 ( \42666 , \42664 , \42665 );
not \U$42416 ( \42667 , \42664 );
and \U$42417 ( \42668 , \42667 , \42654 );
nor \U$42418 ( \42669 , \42666 , \42668 );
buf \U$42419 ( \42670 , \42669 );
and \U$42420 ( \42671 , \42648 , \42651 , \42649 , \42653 );
not \U$42421 ( \42672 , \42671 );
not \U$42422 ( \42673 , \42652 );
or \U$42423 ( \42674 , \42672 , \42673 );
or \U$42424 ( \42675 , \42652 , \42671 );
nand \U$42425 ( \42676 , \42674 , \42675 );
buf \U$42426 ( \42677 , \42676 );
not \U$42427 ( \42678 , \42647 );
nand \U$42428 ( \42679 , \42678 , \42587 , \42649 , \42651 );
not \U$42429 ( \42680 , \42653 );
and \U$42430 ( \42681 , \42679 , \42680 );
not \U$42431 ( \42682 , \42679 );
and \U$42432 ( \42683 , \42682 , \42653 );
nor \U$42433 ( \42684 , \42681 , \42683 );
buf \U$42434 ( \42685 , \42684 );
xor \U$42435 ( \42686 , \42650 , \42651 );
buf \U$42436 ( \42687 , \42686 );
xor \U$42437 ( \42688 , \42648 , \42649 );
buf \U$42438 ( \42689 , \42688 );
not \U$42439 ( \42690 , \42620 );
nand \U$42440 ( \42691 , \42690 , \41271 , \42635 , \42636 );
not \U$42441 ( \42692 , \42624 );
and \U$42442 ( \42693 , \42691 , \42692 );
not \U$42443 ( \42694 , \42691 );
and \U$42444 ( \42695 , \42694 , \42624 );
nor \U$42445 ( \42696 , \42693 , \42695 );
buf \U$42446 ( \42697 , \42696 );
nand \U$42447 ( \42698 , \42621 , \42635 );
and \U$42448 ( \42699 , \42698 , \42645 );
not \U$42449 ( \42700 , \42698 );
and \U$42450 ( \42701 , \42700 , \41271 );
nor \U$42451 ( \42702 , \42699 , \42701 );
buf \U$42452 ( \42703 , \42702 );
and \U$42453 ( \42704 , \42621 , \42635 );
not \U$42454 ( \42705 , \42621 );
and \U$42455 ( \42706 , \42705 , \42159 );
nor \U$42456 ( \42707 , \42704 , \42706 );
buf \U$42457 ( \42708 , \42707 );
and \U$42458 ( \42709 , \42620 , \42163 );
not \U$42459 ( \42710 , \42620 );
and \U$42460 ( \42711 , \42710 , \42636 );
nor \U$42461 ( \42712 , \42709 , \42711 );
buf \U$42462 ( \42713 , \42712 );
buf \U$42463 ( \42714 , \42197 );
buf \U$42464 ( \42715 , \42617 );
and \U$42465 ( \42716 , \42587 , \42714 , \42715 );
and \U$42466 ( \42717 , \42716 , \42204 );
not \U$42467 ( \42718 , \42716 );
not \U$42468 ( \42719 , \42204 );
and \U$42469 ( \42720 , \42718 , \42719 );
nor \U$42470 ( \42721 , \42717 , \42720 );
buf \U$42471 ( \42722 , \42721 );
nand \U$42472 ( \42723 , \42587 , \42715 );
not \U$42473 ( \42724 , \42714 );
and \U$42474 ( \42725 , \42723 , \42724 );
not \U$42475 ( \42726 , \42723 );
and \U$42476 ( \42727 , \42726 , \42714 );
nor \U$42477 ( \42728 , \42725 , \42727 );
buf \U$42478 ( \42729 , \42728 );
not \U$42479 ( \42730 , \42715 );
and \U$42480 ( \42731 , \42586 , \42730 );
not \U$42481 ( \42732 , \42586 );
and \U$42482 ( \42733 , \42732 , \42715 );
nor \U$42483 ( \42734 , \42731 , \42733 );
buf \U$42484 ( \42735 , \42734 );
not \U$42485 ( \42736 , \42560 );
not \U$42486 ( \42737 , \41693 );
not \U$42487 ( \42738 , \42115 );
and \U$42488 ( \42739 , \42737 , \42738 , \42216 );
not \U$42489 ( \42740 , \42135 );
nor \U$42490 ( \42741 , \42740 , \41784 , \41982 );
nand \U$42491 ( \42742 , \42739 , \42131 , \42741 );
xnor \U$42492 ( \42743 , \41441 , \41389 );
nor \U$42493 ( \42744 , \42742 , \42743 );
nand \U$42494 ( \42745 , \42736 , \42744 );
buf \U$42495 ( \42746 , \41395 );
nor \U$42496 ( \42747 , \42745 , \42746 );
buf \U$42497 ( \42748 , \42747 );
not \U$42498 ( \42749 , \41352 );
not \U$42499 ( \42750 , \41416 );
not \U$42500 ( \42751 , \41428 );
or \U$42501 ( \42752 , \42750 , \42751 );
or \U$42502 ( \42753 , \41428 , \41416 );
nand \U$42503 ( \42754 , \42752 , \42753 );
not \U$42504 ( \42755 , \41443 );
nor \U$42505 ( \42756 , \41413 , \42755 );
not \U$42506 ( \42757 , \41357 );
and \U$42507 ( \42758 , \42754 , \42756 , \42582 , \42757 );
nand \U$42508 ( \42759 , \42748 , \42749 , \42758 );
xnor \U$42509 ( \42760 , \42759 , \41341 );
buf \U$42510 ( \42761 , \42760 );
nand \U$42511 ( \42762 , \42748 , \42758 );
not \U$42512 ( \42763 , \42749 );
and \U$42513 ( \42764 , \42762 , \42763 );
not \U$42514 ( \42765 , \42762 );
and \U$42515 ( \42766 , \42765 , \42749 );
nor \U$42516 ( \42767 , \42764 , \42766 );
buf \U$42517 ( \42768 , \42767 );
not \U$42518 ( \42769 , \41412 );
nor \U$42519 ( \42770 , \42757 , \42769 );
not \U$42520 ( \42771 , \42770 );
nand \U$42521 ( \42772 , \42582 , \42747 );
nor \U$42522 ( \42773 , \42772 , \42755 );
nand \U$42523 ( \42774 , \42754 , \42773 );
buf \U$42524 ( \42775 , \41406 );
not \U$42525 ( \42776 , \42775 );
nor \U$42526 ( \42777 , \42774 , \42776 );
not \U$42527 ( \42778 , \42777 );
or \U$42528 ( \42779 , \42771 , \42778 );
not \U$42529 ( \42780 , \41357 );
not \U$42530 ( \42781 , \41413 );
nand \U$42531 ( \42782 , \42781 , \42754 , \42773 );
nand \U$42532 ( \42783 , \42780 , \42782 );
nand \U$42533 ( \42784 , \42779 , \42783 );
buf \U$42534 ( \42785 , \42784 );
and \U$42535 ( \42786 , \42777 , \41412 );
not \U$42536 ( \42787 , \42777 );
and \U$42537 ( \42788 , \42787 , \42769 );
nor \U$42538 ( \42789 , \42786 , \42788 );
buf \U$42539 ( \42790 , \42789 );
and \U$42540 ( \42791 , \42774 , \42776 );
not \U$42541 ( \42792 , \42774 );
and \U$42542 ( \42793 , \42792 , \42775 );
nor \U$42543 ( \42794 , \42791 , \42793 );
buf \U$42544 ( \42795 , \42794 );
buf \U$42545 ( \42796 , \42773 );
and \U$42546 ( \42797 , \42796 , \42754 );
not \U$42547 ( \42798 , \42796 );
not \U$42548 ( \42799 , \42754 );
and \U$42549 ( \42800 , \42798 , \42799 );
nor \U$42550 ( \42801 , \42797 , \42800 );
buf \U$42551 ( \42802 , \42801 );
and \U$42552 ( \42803 , \42772 , \42755 );
not \U$42553 ( \42804 , \42772 );
and \U$42554 ( \42805 , \42804 , \41443 );
nor \U$42555 ( \42806 , \42803 , \42805 );
buf \U$42556 ( \42807 , \42806 );
and \U$42557 ( \42808 , \42748 , \42582 );
not \U$42558 ( \42809 , \42748 );
and \U$42559 ( \42810 , \42809 , \41472 );
nor \U$42560 ( \42811 , \42808 , \42810 );
buf \U$42561 ( \42812 , \42811 );
and \U$42562 ( \42813 , \42745 , \42746 );
not \U$42563 ( \42814 , \42745 );
not \U$42564 ( \42815 , \42746 );
and \U$42565 ( \42816 , \42814 , \42815 );
nor \U$42566 ( \42817 , \42813 , \42816 );
buf \U$42567 ( \42818 , \42817 );
not \U$42568 ( \42819 , \42560 );
and \U$42569 ( \42820 , \42744 , \42819 );
not \U$42570 ( \42821 , \42744 );
and \U$42571 ( \42822 , \42821 , \42560 );
nor \U$42572 ( \42823 , \42820 , \42822 );
buf \U$42573 ( \42824 , \42823 );
xor \U$42574 ( \42825 , \42742 , \42743 );
buf \U$42575 ( \42826 , \42825 );
xnor \U$42576 ( \42827 , \42137 , \42577 );
buf \U$42577 ( \42828 , \42827 );
xnor \U$42578 ( \42829 , \42132 , \42135 );
buf \U$42579 ( \42830 , \42829 );
nor \U$42580 ( \42831 , \41848 , \41800 );
and \U$42581 ( \42832 , \42831 , \41752 );
not \U$42582 ( \42833 , \41781 );
not \U$42583 ( \42834 , \41771 );
nand \U$42584 ( \42835 , \42834 , \41980 );
nor \U$42585 ( \42836 , \42835 , \41769 );
nand \U$42586 ( \42837 , \42836 , \41776 );
nor \U$42587 ( \42838 , \42833 , \42837 );
nand \U$42588 ( \42839 , \42832 , \42838 );
not \U$42589 ( \42840 , \42839 );
nand \U$42590 ( \42841 , \42580 , \41698 , \41699 , \42840 );
not \U$42591 ( \42842 , \42841 );
and \U$42592 ( \42843 , \42124 , \42117 );
not \U$42593 ( \42844 , \42124 );
and \U$42594 ( \42845 , \42844 , \42118 );
nor \U$42595 ( \42846 , \42843 , \42845 );
nand \U$42596 ( \42847 , \42842 , \42846 , \41692 , \41701 );
xnor \U$42597 ( \42848 , \42847 , \41707 );
buf \U$42598 ( \42849 , \42848 );
nand \U$42599 ( \42850 , \42580 , \41699 , \42840 );
not \U$42600 ( \42851 , \42850 );
nand \U$42601 ( \42852 , \42851 , \42846 , \41692 , \41698 );
xnor \U$42602 ( \42853 , \42852 , \41701 );
buf \U$42603 ( \42854 , \42853 );
nand \U$42604 ( \42855 , \42580 , \42840 );
not \U$42605 ( \42856 , \42855 );
nand \U$42606 ( \42857 , \42856 , \41692 , \41698 , \41699 );
xnor \U$42607 ( \42858 , \42857 , \42846 );
buf \U$42608 ( \42859 , \42858 );
xnor \U$42609 ( \42860 , \42841 , \41692 );
buf \U$42610 ( \42861 , \42860 );
and \U$42611 ( \42862 , \42850 , \41697 );
not \U$42612 ( \42863 , \42850 );
and \U$42613 ( \42864 , \42863 , \41698 );
nor \U$42614 ( \42865 , \42862 , \42864 );
buf \U$42615 ( \42866 , \42865 );
xnor \U$42616 ( \42867 , \42855 , \41699 );
buf \U$42617 ( \42868 , \42867 );
not \U$42618 ( \42869 , \42100 );
not \U$42619 ( \42870 , \42027 );
buf \U$42620 ( \42871 , \42025 );
not \U$42621 ( \42872 , \42871 );
nand \U$42622 ( \42873 , \42870 , \42872 , \42832 , \42838 );
nor \U$42623 ( \42874 , \42869 , \42873 );
buf \U$42624 ( \42875 , \41663 );
buf \U$42625 ( \42876 , \41675 );
buf \U$42626 ( \42877 , \41793 );
not \U$42627 ( \42878 , \42877 );
nand \U$42628 ( \42879 , \42874 , \42875 , \42876 , \42878 );
not \U$42629 ( \42880 , \42879 );
buf \U$42630 ( \42881 , \42041 );
buf \U$42631 ( \42882 , \41676 );
buf \U$42632 ( \42883 , \41674 );
and \U$42633 ( \42884 , \42880 , \42881 , \42882 , \42883 );
nand \U$42634 ( \42885 , \42884 , \42114 );
not \U$42635 ( \42886 , \42885 );
buf \U$42636 ( \42887 , \42113 );
nand \U$42637 ( \42888 , \42886 , \42887 );
not \U$42638 ( \42889 , \42888 );
not \U$42639 ( \42890 , \41996 );
buf \U$42640 ( \42891 , \41997 );
buf \U$42641 ( \42892 , \42010 );
nand \U$42642 ( \42893 , \42889 , \42890 , \42891 , \42892 );
buf \U$42643 ( \42894 , \41998 );
not \U$42644 ( \42895 , \42894 );
and \U$42645 ( \42896 , \42893 , \42895 );
not \U$42646 ( \42897 , \42893 );
and \U$42647 ( \42898 , \42897 , \42894 );
nor \U$42648 ( \42899 , \42896 , \42898 );
buf \U$42649 ( \42900 , \42899 );
not \U$42650 ( \42901 , \42892 );
not \U$42651 ( \42902 , \42885 );
nand \U$42652 ( \42903 , \42902 , \42887 , \42890 , \42891 );
not \U$42653 ( \42904 , \42903 );
or \U$42654 ( \42905 , \42901 , \42904 );
or \U$42655 ( \42906 , \42892 , \42903 );
nand \U$42656 ( \42907 , \42905 , \42906 );
buf \U$42657 ( \42908 , \42907 );
nand \U$42658 ( \42909 , \42884 , \42891 , \42114 , \42887 );
and \U$42659 ( \42910 , \42909 , \41996 );
not \U$42660 ( \42911 , \42909 );
and \U$42661 ( \42912 , \42911 , \42890 );
nor \U$42662 ( \42913 , \42910 , \42912 );
buf \U$42663 ( \42914 , \42913 );
not \U$42664 ( \42915 , \42891 );
and \U$42665 ( \42916 , \42888 , \42915 );
not \U$42666 ( \42917 , \42888 );
and \U$42667 ( \42918 , \42917 , \42891 );
nor \U$42668 ( \42919 , \42916 , \42918 );
buf \U$42669 ( \42920 , \42919 );
not \U$42670 ( \42921 , \42887 );
and \U$42671 ( \42922 , \42885 , \42921 );
not \U$42672 ( \42923 , \42885 );
and \U$42673 ( \42924 , \42923 , \42887 );
nor \U$42674 ( \42925 , \42922 , \42924 );
buf \U$42675 ( \42926 , \42925 );
and \U$42676 ( \42927 , \42884 , \42114 );
not \U$42677 ( \42928 , \42884 );
not \U$42678 ( \42929 , \42114 );
and \U$42679 ( \42930 , \42928 , \42929 );
nor \U$42680 ( \42931 , \42927 , \42930 );
buf \U$42681 ( \42932 , \42931 );
not \U$42682 ( \42933 , \42879 );
nand \U$42683 ( \42934 , \42933 , \42883 , \42882 );
not \U$42684 ( \42935 , \42881 );
and \U$42685 ( \42936 , \42934 , \42935 );
not \U$42686 ( \42937 , \42934 );
and \U$42687 ( \42938 , \42937 , \42881 );
nor \U$42688 ( \42939 , \42936 , \42938 );
buf \U$42689 ( \42940 , \42939 );
nand \U$42690 ( \42941 , \42882 , \42880 );
not \U$42691 ( \42942 , \42883 );
and \U$42692 ( \42943 , \42941 , \42942 );
not \U$42693 ( \42944 , \42941 );
and \U$42694 ( \42945 , \42944 , \42883 );
nor \U$42695 ( \42946 , \42943 , \42945 );
buf \U$42696 ( \42947 , \42946 );
not \U$42697 ( \42948 , \42882 );
and \U$42698 ( \42949 , \42879 , \42948 );
not \U$42699 ( \42950 , \42879 );
and \U$42700 ( \42951 , \42950 , \42882 );
nor \U$42701 ( \42952 , \42949 , \42951 );
buf \U$42702 ( \42953 , \42952 );
not \U$42703 ( \42954 , \42875 );
nand \U$42704 ( \42955 , \42874 , \42876 );
nor \U$42705 ( \42956 , \42954 , \42955 );
and \U$42706 ( \42957 , \42956 , \42878 );
not \U$42707 ( \42958 , \42956 );
and \U$42708 ( \42959 , \42958 , \42877 );
nor \U$42709 ( \42960 , \42957 , \42959 );
buf \U$42710 ( \42961 , \42960 );
and \U$42711 ( \42962 , \42955 , \42954 );
not \U$42712 ( \42963 , \42955 );
and \U$42713 ( \42964 , \42963 , \42875 );
nor \U$42714 ( \42965 , \42962 , \42964 );
buf \U$42715 ( \42966 , \42965 );
xor \U$42716 ( \42967 , \42874 , \42876 );
buf \U$42717 ( \42968 , \42967 );
buf \U$42718 ( \42969 , \42096 );
not \U$42719 ( \42970 , \42969 );
nor \U$42720 ( \42971 , \42873 , \42970 );
nand \U$42721 ( \42972 , \42971 , \42091 );
not \U$42722 ( \42973 , \42972 );
not \U$42723 ( \42974 , \42074 );
not \U$42724 ( \42975 , \42974 );
nand \U$42725 ( \42976 , \42973 , \42975 , \42097 , \42077 );
not \U$42726 ( \42977 , \42976 );
buf \U$42727 ( \42978 , \42066 );
not \U$42728 ( \42979 , \42978 );
nand \U$42729 ( \42980 , \42977 , \42979 , \42095 , \42075 );
and \U$42730 ( \42981 , \42980 , \42072 );
not \U$42731 ( \42982 , \42980 );
not \U$42732 ( \42983 , \42072 );
and \U$42733 ( \42984 , \42982 , \42983 );
nor \U$42734 ( \42985 , \42981 , \42984 );
buf \U$42735 ( \42986 , \42985 );
nand \U$42736 ( \42987 , \42971 , \42091 , \42074 , \42077 );
not \U$42737 ( \42988 , \42987 );
nand \U$42738 ( \42989 , \42988 , \42979 , \42095 , \42097 );
xnor \U$42739 ( \42990 , \42989 , \42075 );
buf \U$42740 ( \42991 , \42990 );
not \U$42741 ( \42992 , \42873 );
nand \U$42742 ( \42993 , \42992 , \42091 , \42969 , \42077 );
not \U$42743 ( \42994 , \42993 );
nand \U$42744 ( \42995 , \42994 , \42095 , \42097 , \42074 );
and \U$42745 ( \42996 , \42995 , \42978 );
not \U$42746 ( \42997 , \42995 );
and \U$42747 ( \42998 , \42997 , \42979 );
nor \U$42748 ( \42999 , \42996 , \42998 );
buf \U$42749 ( \43000 , \42999 );
xnor \U$42750 ( \43001 , \42976 , \42095 );
buf \U$42751 ( \43002 , \43001 );
xnor \U$42752 ( \43003 , \42097 , \42987 );
buf \U$42753 ( \43004 , \43003 );
and \U$42754 ( \43005 , \42993 , \42974 );
not \U$42755 ( \43006 , \42993 );
and \U$42756 ( \43007 , \43006 , \42074 );
nor \U$42757 ( \43008 , \43005 , \43007 );
buf \U$42758 ( \43009 , \43008 );
not \U$42759 ( \43010 , \42077 );
not \U$42760 ( \43011 , \42972 );
or \U$42761 ( \43012 , \43010 , \43011 );
or \U$42762 ( \43013 , \42077 , \42972 );
nand \U$42763 ( \43014 , \43012 , \43013 );
buf \U$42764 ( \43015 , \43014 );
xor \U$42765 ( \43016 , \42971 , \42091 );
buf \U$42766 ( \43017 , \43016 );
and \U$42767 ( \43018 , \42873 , \42970 );
not \U$42768 ( \43019 , \42873 );
and \U$42769 ( \43020 , \43019 , \42969 );
nor \U$42770 ( \43021 , \43018 , \43020 );
buf \U$42771 ( \43022 , \43021 );
nor \U$42772 ( \43023 , \42839 , \42027 );
not \U$42773 ( \43024 , \42871 );
and \U$42774 ( \43025 , \43023 , \43024 );
not \U$42775 ( \43026 , \43023 );
and \U$42776 ( \43027 , \43026 , \42871 );
nor \U$42777 ( \43028 , \43025 , \43027 );
buf \U$42778 ( \43029 , \43028 );
xor \U$42779 ( \43030 , \42839 , \42027 );
buf \U$42780 ( \43031 , \43030 );
not \U$42781 ( \43032 , \41840 );
buf \U$42782 ( \43033 , \42838 );
nand \U$42783 ( \43034 , \43033 , \41829 , \41821 );
nor \U$42784 ( \43035 , \43034 , \41831 );
and \U$42785 ( \43036 , \43032 , \43035 );
nand \U$42786 ( \43037 , \43036 , \41847 );
not \U$42787 ( \43038 , \43037 );
buf \U$42788 ( \43039 , \42571 );
buf \U$42789 ( \43040 , \41801 );
nand \U$42790 ( \43041 , \43038 , \43039 , \43040 , \41813 );
not \U$42791 ( \43042 , \41816 );
and \U$42792 ( \43043 , \43041 , \43042 );
not \U$42793 ( \43044 , \43041 );
and \U$42794 ( \43045 , \43044 , \41816 );
nor \U$42795 ( \43046 , \43043 , \43045 );
buf \U$42796 ( \43047 , \43046 );
nand \U$42797 ( \43048 , \43036 , \43040 , \41847 , \43039 );
xnor \U$42798 ( \43049 , \43048 , \41813 );
buf \U$42799 ( \43050 , \43049 );
nand \U$42800 ( \43051 , \43036 , \43040 , \41847 );
not \U$42801 ( \43052 , \43039 );
and \U$42802 ( \43053 , \43051 , \43052 );
not \U$42803 ( \43054 , \43051 );
and \U$42804 ( \43055 , \43054 , \43039 );
nor \U$42805 ( \43056 , \43053 , \43055 );
buf \U$42806 ( \43057 , \43056 );
not \U$42807 ( \43058 , \43040 );
and \U$42808 ( \43059 , \43037 , \43058 );
not \U$42809 ( \43060 , \43037 );
and \U$42810 ( \43061 , \43060 , \43040 );
nor \U$42811 ( \43062 , \43059 , \43061 );
buf \U$42812 ( \43063 , \43062 );
xor \U$42813 ( \43064 , \43036 , \41847 );
buf \U$42814 ( \43065 , \43064 );
and \U$42815 ( \43066 , \43035 , \43032 );
not \U$42816 ( \43067 , \43035 );
and \U$42817 ( \43068 , \43067 , \41840 );
nor \U$42818 ( \43069 , \43066 , \43068 );
buf \U$42819 ( \43070 , \43069 );
xor \U$42820 ( \43071 , \43034 , \41831 );
buf \U$42821 ( \43072 , \43071 );
nand \U$42822 ( \43073 , \43033 , \41829 );
xnor \U$42823 ( \43074 , \43073 , \41821 );
buf \U$42824 ( \43075 , \43074 );
xor \U$42825 ( \43076 , \43033 , \41829 );
buf \U$42826 ( \43077 , \43076 );
not \U$42827 ( \43078 , \42837 );
not \U$42828 ( \43079 , \41781 );
or \U$42829 ( \43080 , \43078 , \43079 );
or \U$42830 ( \43081 , \41781 , \42837 );
nand \U$42831 ( \43082 , \43080 , \43081 );
buf \U$42832 ( \43083 , \43082 );
xor \U$42833 ( \43084 , \42836 , \41776 );
buf \U$42834 ( \43085 , \43084 );
not \U$42835 ( \43086 , \41769 );
not \U$42836 ( \43087 , \42835 );
not \U$42837 ( \43088 , \43087 );
or \U$42838 ( \43089 , \43086 , \43088 );
or \U$42839 ( \43090 , \41769 , \43087 );
nand \U$42840 ( \43091 , \43089 , \43090 );
buf \U$42841 ( \43092 , \43091 );
not \U$42842 ( \43093 , \41771 );
not \U$42843 ( \43094 , \41980 );
or \U$42844 ( \43095 , \43093 , \43094 );
or \U$42845 ( \43096 , \41771 , \41980 );
nand \U$42846 ( \43097 , \43095 , \43096 );
buf \U$42847 ( \43098 , \43097 );
not \U$42848 ( \43099 , \41979 );
not \U$42849 ( \43100 , \41978 );
not \U$42850 ( \43101 , \43100 );
or \U$42851 ( \43102 , \43099 , \43101 );
or \U$42852 ( \43103 , \41979 , \43100 );
nand \U$42853 ( \43104 , \43102 , \43103 );
buf \U$42854 ( \43105 , \43104 );
not \U$42855 ( \43106 , \41879 );
buf \U$42856 ( \43107 , \41864 );
nand \U$42857 ( \43108 , \41977 , \43107 );
not \U$42858 ( \43109 , \41893 );
nor \U$42859 ( \43110 , \43108 , \43109 );
nand \U$42860 ( \43111 , \43106 , \43110 );
not \U$42861 ( \43112 , \43111 );
buf \U$42862 ( \43113 , \41878 );
nand \U$42863 ( \43114 , \43112 , \43113 );
not \U$42864 ( \43115 , \43114 );
buf \U$42865 ( \43116 , \41899 );
nand \U$42866 ( \43117 , \43115 , \43116 );
not \U$42867 ( \43118 , \43117 );
nand \U$42868 ( \43119 , \43118 , \41906 );
xor \U$42869 ( \43120 , \43119 , \41880 );
buf \U$42870 ( \43121 , \43120 );
xnor \U$42871 ( \43122 , \43117 , \41906 );
buf \U$42872 ( \43123 , \43122 );
xnor \U$42873 ( \43124 , \43114 , \43116 );
buf \U$42874 ( \43125 , \43124 );
xnor \U$42875 ( \43126 , \43111 , \43113 );
buf \U$42876 ( \43127 , \43126 );
and \U$42877 ( \43128 , \43110 , \43106 );
not \U$42878 ( \43129 , \43110 );
and \U$42879 ( \43130 , \43129 , \41879 );
nor \U$42880 ( \43131 , \43128 , \43130 );
buf \U$42881 ( \43132 , \43131 );
and \U$42882 ( \43133 , \43108 , \43109 );
not \U$42883 ( \43134 , \43108 );
and \U$42884 ( \43135 , \43134 , \41893 );
nor \U$42885 ( \43136 , \43133 , \43135 );
buf \U$42886 ( \43137 , \43136 );
xor \U$42887 ( \43138 , \41977 , \43107 );
buf \U$42888 ( \43139 , \43138 );
xor \U$42889 ( \43140 , \41975 , \41976 );
buf \U$42890 ( \43141 , \43140 );
xor \U$42891 ( \43142 , \41973 , \41974 );
buf \U$42892 ( \43143 , \43142 );
xor \U$42893 ( \43144 , \41971 , \41972 );
buf \U$42894 ( \43145 , \43144 );
xor \U$42895 ( \43146 , \41969 , \41970 );
buf \U$42896 ( \43147 , \43146 );
xor \U$42897 ( \43148 , \41963 , \41968 );
buf \U$42898 ( \43149 , \43148 );
xor \U$42899 ( \43150 , \41957 , \41962 );
buf \U$42900 ( \43151 , \43150 );
and \U$42901 ( \43152 , \41956 , \41948 );
not \U$42902 ( \43153 , \41956 );
and \U$42903 ( \43154 , \43153 , \41947 );
nor \U$42904 ( \43155 , \43152 , \43154 );
buf \U$42905 ( \43156 , \43155 );
endmodule

