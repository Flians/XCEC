//
// Conformal-LEC Version 20.10-d213 (02-Sep-2020)
//
module top(RIae78da0_130,RIae78b48_125,RIae78c38_127,RIae78bc0_126,RIae78cb0_128,RIae78e90_132,RIae78ff8_135,RIae78a58_123,RIae76b68_57,
        RIae78f80_134,RIae78f08_133,RIae76988_53,RIae79070_136,RIae790e8_137,RIae76a78_55,RIae767a8_49,RIae76898_51,RIae79160_138,RIae792c8_141,
        RIae76208_37,RIae762f8_39,RIae79250_140,RIae791d8_139,RIae76118_35,RIae76028_33,RIae793b8_143,RIae79340_142,RIae765c8_45,RIae766b8_47,
        RIae764d8_43,RIae79610_148,RIae799d0_156,RIae763e8_41,RIae79688_149,RIae79598_147,RIae753f8_7,RIae75308_5,RIae79ac0_158,RIae79b38_159,
        RIae75128_1,RIae75218_3,RIae79520_146,RIae79a48_157,RIae756c8_13,RIae757b8_15,RIae79430_144,RIae794a8_145,RIae755d8_11,RIae754e8_9,
        RIae75e48_29,RIae75c68_25,RIae75d58_27,RIae797f0_152,RIae79868_153,RIae798e0_154,RIae79958_155,RIae75f38_31,RIae79700_150,RIae79778_151,
        RIae75998_19,RIae758a8_17,RIae79c28_161,RIae79bb0_160,RIae75a88_21,RIae75b78_23,RIae79ca0_162,RIae79d18_163,RIae78698_115,RIae78788_117,
        RIae79d90_164,RIae79e08_165,RIae78878_119,RIae79ef8_167,RIae79e80_166,RIae78968_121,RIae77e28_97,RIae77d38_95,RIae79f70_168,RIae79fe8_169,
        RIae7a2b8_175,RIae7a678_183,RIae77c48_93,RIae77b58_91,RIae7a240_174,RIae7a1c8_173,RIae783c8_109,RIae78530_112,RIae785a8_113,RIae781e8_105,
        RIae78008_101,RIae7a3a8_177,RIae7a330_176,RIae77f18_99,RIae7a510_180,RIae7a600_182,RIae782d8_107,RIae780f8_103,RIae7a588_181,RIae7a498_179,
        RIae772e8_73,RIae771f8_71,RIae7a150_172,RIae7a420_178,RIae77018_67,RIae77180_70,RIae7a060_170,RIae7a0d8_171,RIae76c58_59,RIae76d48_61,
        RIae7a7e0_186,RIae7a948_189,RIae76e38_63,RIae76f28_65,RIae77888_85,RIae7a6f0_184,RIae7a768_185,RIae77798_83,RIae7a8d0_188,RIae7a858_187,
        RIae77a68_89,RIae77978_87,RIae7aa38_191,RIae7a9c0_190,RIae773d8_75,RIae77720_82,RIae774c8_77,RIae7aab0_192,RIae775b8_79,RIae78e18_131,
        RIae78d28_129,RIae78ad0_124,RIae76be0_58,RIae76820_50,RIae76910_52,RIae76a00_54,RIae76af0_56,RIae76280_38,RIae76370_40,RIae760a0_34,
        RIae76190_36,RIae76640_46,RIae76460_42,RIae76550_44,RIae76730_48,RIae75470_8,RIae75380_6,RIae751a0_2,RIae75290_4,RIae75740_14,
        RIae75830_16,RIae75650_12,RIae75560_10,RIae75ce0_26,RIae75dd0_28,RIae75ec0_30,RIae75fb0_32,RIae75920_18,RIae75a10_20,RIae75b00_22,
        RIae75bf0_24,RIae78710_116,RIae78800_118,RIae77bd0_92,RIae77db0_96,RIae77ea0_98,RIae789e0_122,RIae77cc0_94,RIae788f0_120,RIae78440_110,
        RIae784b8_111,RIae78620_114,RIae78260_106,RIae78080_102,RIae77f90_100,RIae78170_104,RIae78350_108,RIae77360_74,RIae77270_72,RIae77090_68,
        RIae77108_69,RIae76cd0_60,RIae76dc0_62,RIae76eb0_64,RIae76fa0_66,RIae77900_86,RIae77810_84,RIae77ae0_90,RIae779f0_88,RIae77450_76,
        RIae776a8_81,RIae77540_78,RIae77630_80,RIae7c8b0_256,RIae7bfc8_237,RIae7c298_243,RIae7c838_255,RIae7b9b0_224,RIae7ab28_193,RIae7b398_211,
        RIae7c658_251,RIae7b578_215,RIae7b6e0_218,RIae7b2a8_209,RIae7bf50_236,RIae7b848_221,RIae7b938_223,RIae7bb90_228,RIae7afd8_203,RIae7c7c0_254,
        RIae7bc80_230,RIae7b8c0_222,RIae7b500_214,RIae7b410_212,RIae7c400_246,RIae7be60_234,RIae7c130_240,RIae7c310_244,RIae7c568_249,RIae7aba0_194,
        RIae7c6d0_252,RIae7ad80_198,RIae7b140_206,RIae7b050_204,RIae7c0b8_239,RIae7bc08_229,RIae7c748_253,RIae7c388_245,RIae7b488_213,RIae7b5f0_216,
        RIae7ac90_196,RIae7c040_238,RIae7c5e0_250,RIae7c478_247,RIae7b320_210,RIae7adf8_199,RIae7af60_202,RIae7b758_219,RIae7bcf8_231,RIae7b668_217,
        RIae7ad08_197,RIae7ac18_195,RIae7bd70_232,RIae7b7d0_220,RIae7aee8_201,RIae7c1a8_241,RIae7b1b8_207,RIae7ae70_200,RIae7c4f0_248,RIae7bde8_233,
        RIae7c220_242,RIae7bed8_235,RIae7b0c8_205,RIae7bb18_227,RIae7ba28_225,RIae7baa0_226,RIae7b230_208,R_101_77c8620,R_102_af8fd30,R_103_af901c8,
        R_104_af9a140,R_105_af99768,R_106_af8be30,R_107_77c1150,R_108_af8ddb0,R_109_af8f010,R_10a_af996c0,R_10b_77c34c0,R_10c_77c28f0,R_10d_af8d090,
        R_10e_77ca5a0,R_10f_77ce4a0,R_110_77cd780,R_111_af8f2b0,R_112_77c6550,R_113_af98ee0,R_114_77c2068,R_115_af99ea0,R_116_77c0eb0,R_117_77cc280,
        R_118_77bf860,R_119_77c9f10,R_11a_af8bf80,R_11b_77bf320,R_11c_77c4fa8,R_11d_af99ab0,R_11e_77ca258,R_11f_af92880,R_120_af91c08,R_121_af92298,
        R_122_af99ca8,R_123_af990d8,R_124_77c5638,R_125_af8e6e0,R_126_77c3aa8,R_127_77c8d58,R_128_77c1fc0,R_129_77c6748,R_12a_77c3370,R_12b_af99d50,
        R_12c_77c5248,R_12d_77ca840,R_12e_af8eec0,R_12f_77c1498,R_130_77c5398,R_131_77c0820,R_132_af8d480,R_133_77ce890,R_134_af97c80,R_135_77c65f8,
        R_136_af8d678,R_137_77c3e98,R_138_af8e0f8,R_139_af99378,R_13a_77c7078,R_13b_77ce740,R_13c_af97fc8,R_13d_77c62b0,R_13e_77c27a0,R_13f_af979e0,
        R_140_77c25a8,R_141_af921f0,R_142_af8b7a0,R_143_77bfcf8,R_144_af92148,R_145_77c1c78,R_146_77cb560,R_147_af99960,R_148_af92490,R_149_77c9298,
        R_14a_77cb170,R_14b_af98268,R_14c_77bf9b0,R_14d_af91b60,R_14e_af8f208,R_14f_77c7a50,R_150_af99030,R_151_77c67f0,R_152_af8c370,R_153_77c8818,
        R_154_77c6d30,R_155_af98c40,R_156_77c9538,R_157_af96f60,R_158_af96d68,R_159_af8d870,R_15a_af8e830,R_15b_77ccbb0,R_15c_af8c610,R_15d_77c6898,
        R_15e_af8cb50,R_15f_af92538,R_160_af975f0,R_161_77c71c8,R_162_af8d720,R_163_77cb608,R_164_af8b650,R_165_af988f8,R_166_77c41e0,R_167_af8e398,
        R_168_af974a0,R_169_af8d330,R_16a_af8c0d0,R_16b_77cc520,R_16c_77cb8a8,R_16d_77ccda8,R_16e_af973f8,R_16f_77cd6d8,R_170_af99ff0,R_171_77c54e8,
        R_172_77c3808,R_173_77c0580,R_174_af99618,R_175_77cd198,R_176_77c0628,R_177_af97698);
input RIae78da0_130,RIae78b48_125,RIae78c38_127,RIae78bc0_126,RIae78cb0_128,RIae78e90_132,RIae78ff8_135,RIae78a58_123,RIae76b68_57,
        RIae78f80_134,RIae78f08_133,RIae76988_53,RIae79070_136,RIae790e8_137,RIae76a78_55,RIae767a8_49,RIae76898_51,RIae79160_138,RIae792c8_141,
        RIae76208_37,RIae762f8_39,RIae79250_140,RIae791d8_139,RIae76118_35,RIae76028_33,RIae793b8_143,RIae79340_142,RIae765c8_45,RIae766b8_47,
        RIae764d8_43,RIae79610_148,RIae799d0_156,RIae763e8_41,RIae79688_149,RIae79598_147,RIae753f8_7,RIae75308_5,RIae79ac0_158,RIae79b38_159,
        RIae75128_1,RIae75218_3,RIae79520_146,RIae79a48_157,RIae756c8_13,RIae757b8_15,RIae79430_144,RIae794a8_145,RIae755d8_11,RIae754e8_9,
        RIae75e48_29,RIae75c68_25,RIae75d58_27,RIae797f0_152,RIae79868_153,RIae798e0_154,RIae79958_155,RIae75f38_31,RIae79700_150,RIae79778_151,
        RIae75998_19,RIae758a8_17,RIae79c28_161,RIae79bb0_160,RIae75a88_21,RIae75b78_23,RIae79ca0_162,RIae79d18_163,RIae78698_115,RIae78788_117,
        RIae79d90_164,RIae79e08_165,RIae78878_119,RIae79ef8_167,RIae79e80_166,RIae78968_121,RIae77e28_97,RIae77d38_95,RIae79f70_168,RIae79fe8_169,
        RIae7a2b8_175,RIae7a678_183,RIae77c48_93,RIae77b58_91,RIae7a240_174,RIae7a1c8_173,RIae783c8_109,RIae78530_112,RIae785a8_113,RIae781e8_105,
        RIae78008_101,RIae7a3a8_177,RIae7a330_176,RIae77f18_99,RIae7a510_180,RIae7a600_182,RIae782d8_107,RIae780f8_103,RIae7a588_181,RIae7a498_179,
        RIae772e8_73,RIae771f8_71,RIae7a150_172,RIae7a420_178,RIae77018_67,RIae77180_70,RIae7a060_170,RIae7a0d8_171,RIae76c58_59,RIae76d48_61,
        RIae7a7e0_186,RIae7a948_189,RIae76e38_63,RIae76f28_65,RIae77888_85,RIae7a6f0_184,RIae7a768_185,RIae77798_83,RIae7a8d0_188,RIae7a858_187,
        RIae77a68_89,RIae77978_87,RIae7aa38_191,RIae7a9c0_190,RIae773d8_75,RIae77720_82,RIae774c8_77,RIae7aab0_192,RIae775b8_79,RIae78e18_131,
        RIae78d28_129,RIae78ad0_124,RIae76be0_58,RIae76820_50,RIae76910_52,RIae76a00_54,RIae76af0_56,RIae76280_38,RIae76370_40,RIae760a0_34,
        RIae76190_36,RIae76640_46,RIae76460_42,RIae76550_44,RIae76730_48,RIae75470_8,RIae75380_6,RIae751a0_2,RIae75290_4,RIae75740_14,
        RIae75830_16,RIae75650_12,RIae75560_10,RIae75ce0_26,RIae75dd0_28,RIae75ec0_30,RIae75fb0_32,RIae75920_18,RIae75a10_20,RIae75b00_22,
        RIae75bf0_24,RIae78710_116,RIae78800_118,RIae77bd0_92,RIae77db0_96,RIae77ea0_98,RIae789e0_122,RIae77cc0_94,RIae788f0_120,RIae78440_110,
        RIae784b8_111,RIae78620_114,RIae78260_106,RIae78080_102,RIae77f90_100,RIae78170_104,RIae78350_108,RIae77360_74,RIae77270_72,RIae77090_68,
        RIae77108_69,RIae76cd0_60,RIae76dc0_62,RIae76eb0_64,RIae76fa0_66,RIae77900_86,RIae77810_84,RIae77ae0_90,RIae779f0_88,RIae77450_76,
        RIae776a8_81,RIae77540_78,RIae77630_80,RIae7c8b0_256,RIae7bfc8_237,RIae7c298_243,RIae7c838_255,RIae7b9b0_224,RIae7ab28_193,RIae7b398_211,
        RIae7c658_251,RIae7b578_215,RIae7b6e0_218,RIae7b2a8_209,RIae7bf50_236,RIae7b848_221,RIae7b938_223,RIae7bb90_228,RIae7afd8_203,RIae7c7c0_254,
        RIae7bc80_230,RIae7b8c0_222,RIae7b500_214,RIae7b410_212,RIae7c400_246,RIae7be60_234,RIae7c130_240,RIae7c310_244,RIae7c568_249,RIae7aba0_194,
        RIae7c6d0_252,RIae7ad80_198,RIae7b140_206,RIae7b050_204,RIae7c0b8_239,RIae7bc08_229,RIae7c748_253,RIae7c388_245,RIae7b488_213,RIae7b5f0_216,
        RIae7ac90_196,RIae7c040_238,RIae7c5e0_250,RIae7c478_247,RIae7b320_210,RIae7adf8_199,RIae7af60_202,RIae7b758_219,RIae7bcf8_231,RIae7b668_217,
        RIae7ad08_197,RIae7ac18_195,RIae7bd70_232,RIae7b7d0_220,RIae7aee8_201,RIae7c1a8_241,RIae7b1b8_207,RIae7ae70_200,RIae7c4f0_248,RIae7bde8_233,
        RIae7c220_242,RIae7bed8_235,RIae7b0c8_205,RIae7bb18_227,RIae7ba28_225,RIae7baa0_226,RIae7b230_208;
output R_101_77c8620,R_102_af8fd30,R_103_af901c8,R_104_af9a140,R_105_af99768,R_106_af8be30,R_107_77c1150,R_108_af8ddb0,R_109_af8f010,
        R_10a_af996c0,R_10b_77c34c0,R_10c_77c28f0,R_10d_af8d090,R_10e_77ca5a0,R_10f_77ce4a0,R_110_77cd780,R_111_af8f2b0,R_112_77c6550,R_113_af98ee0,
        R_114_77c2068,R_115_af99ea0,R_116_77c0eb0,R_117_77cc280,R_118_77bf860,R_119_77c9f10,R_11a_af8bf80,R_11b_77bf320,R_11c_77c4fa8,R_11d_af99ab0,
        R_11e_77ca258,R_11f_af92880,R_120_af91c08,R_121_af92298,R_122_af99ca8,R_123_af990d8,R_124_77c5638,R_125_af8e6e0,R_126_77c3aa8,R_127_77c8d58,
        R_128_77c1fc0,R_129_77c6748,R_12a_77c3370,R_12b_af99d50,R_12c_77c5248,R_12d_77ca840,R_12e_af8eec0,R_12f_77c1498,R_130_77c5398,R_131_77c0820,
        R_132_af8d480,R_133_77ce890,R_134_af97c80,R_135_77c65f8,R_136_af8d678,R_137_77c3e98,R_138_af8e0f8,R_139_af99378,R_13a_77c7078,R_13b_77ce740,
        R_13c_af97fc8,R_13d_77c62b0,R_13e_77c27a0,R_13f_af979e0,R_140_77c25a8,R_141_af921f0,R_142_af8b7a0,R_143_77bfcf8,R_144_af92148,R_145_77c1c78,
        R_146_77cb560,R_147_af99960,R_148_af92490,R_149_77c9298,R_14a_77cb170,R_14b_af98268,R_14c_77bf9b0,R_14d_af91b60,R_14e_af8f208,R_14f_77c7a50,
        R_150_af99030,R_151_77c67f0,R_152_af8c370,R_153_77c8818,R_154_77c6d30,R_155_af98c40,R_156_77c9538,R_157_af96f60,R_158_af96d68,R_159_af8d870,
        R_15a_af8e830,R_15b_77ccbb0,R_15c_af8c610,R_15d_77c6898,R_15e_af8cb50,R_15f_af92538,R_160_af975f0,R_161_77c71c8,R_162_af8d720,R_163_77cb608,
        R_164_af8b650,R_165_af988f8,R_166_77c41e0,R_167_af8e398,R_168_af974a0,R_169_af8d330,R_16a_af8c0d0,R_16b_77cc520,R_16c_77cb8a8,R_16d_77ccda8,
        R_16e_af973f8,R_16f_77cd6d8,R_170_af99ff0,R_171_77c54e8,R_172_77c3808,R_173_77c0580,R_174_af99618,R_175_77cd198,R_176_77c0628,R_177_af97698;

wire \376_ZERO , \377_ONE , \378 , \379 , \380 , \381 , \382 , \383 , \384 ,
         \385 , \386 , \387 , \388 , \389 , \390 , \391 , \392 , \393 , \394 ,
         \395 , \396 , \397 , \398 , \399 , \400 , \401 , \402 , \403 , \404 ,
         \405 , \406 , \407 , \408 , \409 , \410 , \411 , \412 , \413 , \414 ,
         \415 , \416 , \417 , \418 , \419 , \420 , \421 , \422 , \423 , \424 ,
         \425 , \426 , \427 , \428 , \429 , \430 , \431 , \432 , \433 , \434 ,
         \435 , \436 , \437 , \438 , \439 , \440 , \441 , \442 , \443 , \444 ,
         \445 , \446 , \447 , \448 , \449 , \450 , \451 , \452 , \453 , \454 ,
         \455 , \456 , \457 , \458 , \459 , \460 , \461 , \462 , \463 , \464 ,
         \465 , \466 , \467 , \468 , \469 , \470 , \471 , \472 , \473 , \474 ,
         \475 , \476 , \477 , \478 , \479 , \480 , \481 , \482 , \483 , \484 ,
         \485 , \486 , \487 , \488 , \489 , \490 , \491 , \492 , \493 , \494 ,
         \495 , \496 , \497 , \498 , \499 , \500 , \501 , \502 , \503 , \504 ,
         \505 , \506 , \507 , \508 , \509 , \510 , \511 , \512 , \513 , \514 ,
         \515 , \516 , \517 , \518 , \519 , \520 , \521 , \522 , \523 , \524 ,
         \525 , \526 , \527 , \528 , \529 , \530 , \531 , \532 , \533 , \534 ,
         \535 , \536 , \537 , \538 , \539 , \540 , \541 , \542 , \543 , \544 ,
         \545 , \546 , \547 , \548 , \549 , \550 , \551 , \552 , \553 , \554 ,
         \555 , \556 , \557 , \558 , \559 , \560 , \561 , \562 , \563 , \564 ,
         \565 , \566 , \567 , \568 , \569 , \570 , \571 , \572 , \573 , \574 ,
         \575 , \576 , \577 , \578 , \579 , \580 , \581 , \582 , \583 , \584 ,
         \585 , \586 , \587 , \588 , \589 , \590 , \591 , \592 , \593 , \594 ,
         \595 , \596 , \597 , \598 , \599 , \600 , \601 , \602 , \603 , \604 ,
         \605 , \606 , \607 , \608 , \609 , \610 , \611 , \612 , \613 , \614 ,
         \615 , \616 , \617 , \618 , \619 , \620 , \621 , \622 , \623 , \624 ,
         \625 , \626 , \627 , \628 , \629 , \630 , \631 , \632 , \633 , \634 ,
         \635 , \636 , \637 , \638 , \639 , \640 , \641 , \642 , \643 , \644 ,
         \645 , \646 , \647 , \648 , \649 , \650 , \651 , \652 , \653 , \654 ,
         \655 , \656 , \657 , \658 , \659 , \660 , \661 , \662 , \663 , \664 ,
         \665 , \666 , \667 , \668 , \669 , \670 , \671 , \672 , \673 , \674 ,
         \675 , \676 , \677 , \678 , \679 , \680 , \681 , \682 , \683 , \684 ,
         \685 , \686 , \687 , \688 , \689 , \690 , \691 , \692 , \693 , \694 ,
         \695 , \696 , \697 , \698 , \699 , \700 , \701 , \702 , \703 , \704 ,
         \705 , \706 , \707 , \708 , \709 , \710 , \711 , \712 , \713 , \714 ,
         \715 , \716 , \717 , \718 , \719 , \720 , \721 , \722 , \723 , \724 ,
         \725 , \726 , \727 , \728 , \729 , \730 , \731 , \732 , \733 , \734 ,
         \735 , \736 , \737 , \738 , \739 , \740 , \741 , \742 , \743 , \744 ,
         \745 , \746 , \747 , \748 , \749 , \750 , \751 , \752 , \753 , \754 ,
         \755 , \756 , \757 , \758 , \759 , \760 , \761 , \762 , \763 , \764 ,
         \765 , \766 , \767 , \768 , \769 , \770 , \771 , \772 , \773 , \774 ,
         \775 , \776 , \777 , \778 , \779 , \780 , \781 , \782 , \783 , \784 ,
         \785 , \786 , \787 , \788 , \789 , \790 , \791 , \792 , \793 , \794 ,
         \795 , \796 , \797 , \798 , \799 , \800 , \801 , \802 , \803 , \804 ,
         \805 , \806 , \807 , \808 , \809 , \810 , \811 , \812 , \813 , \814 ,
         \815 , \816 , \817 , \818 , \819 , \820 , \821 , \822 , \823 , \824 ,
         \825 , \826 , \827 , \828 , \829 , \830 , \831 , \832 , \833 , \834 ,
         \835 , \836 , \837 , \838 , \839 , \840 , \841 , \842 , \843 , \844 ,
         \845 , \846 , \847 , \848 , \849 , \850 , \851 , \852 , \853 , \854 ,
         \855 , \856 , \857 , \858 , \859 , \860 , \861 , \862 , \863 , \864 ,
         \865 , \866 , \867 , \868 , \869 , \870 , \871 , \872 , \873 , \874 ,
         \875 , \876 , \877 , \878 , \879 , \880 , \881 , \882 , \883 , \884 ,
         \885 , \886 , \887 , \888 , \889 , \890 , \891 , \892 , \893 , \894 ,
         \895 , \896 , \897 , \898 , \899 , \900 , \901 , \902 , \903 , \904 ,
         \905 , \906 , \907 , \908 , \909 , \910 , \911 , \912 , \913 , \914 ,
         \915 , \916 , \917 , \918 , \919 , \920 , \921 , \922 , \923 , \924 ,
         \925 , \926 , \927 , \928 , \929 , \930 , \931 , \932 , \933 , \934 ,
         \935 , \936 , \937 , \938 , \939 , \940 , \941 , \942 , \943 , \944 ,
         \945 , \946 , \947 , \948 , \949 , \950 , \951 , \952 , \953 , \954 ,
         \955 , \956 , \957 , \958 , \959 , \960 , \961 , \962 , \963 , \964 ,
         \965 , \966 , \967 , \968 , \969 , \970 , \971 , \972 , \973 , \974 ,
         \975 , \976 , \977 , \978 , \979 , \980 , \981 , \982 , \983 , \984 ,
         \985 , \986 , \987 , \988 , \989 , \990 , \991 , \992 , \993 , \994 ,
         \995 , \996 , \997 , \998 , \999 , \1000 , \1001 , \1002 , \1003 , \1004 ,
         \1005 , \1006 , \1007 , \1008 , \1009 , \1010 , \1011 , \1012 , \1013 , \1014 ,
         \1015 , \1016 , \1017 , \1018 , \1019 , \1020 , \1021 , \1022 , \1023 , \1024 ,
         \1025 , \1026 , \1027 , \1028 , \1029 , \1030 , \1031 , \1032 , \1033 , \1034 ,
         \1035 , \1036 , \1037 , \1038 , \1039 , \1040 , \1041 , \1042 , \1043 , \1044 ,
         \1045 , \1046 , \1047 , \1048 , \1049 , \1050 , \1051 , \1052 , \1053 , \1054 ,
         \1055 , \1056 , \1057 , \1058 , \1059 , \1060 , \1061 , \1062 , \1063 , \1064 ,
         \1065 , \1066 , \1067 , \1068 , \1069 , \1070 , \1071 , \1072 , \1073 , \1074 ,
         \1075 , \1076 , \1077 , \1078 , \1079 , \1080 , \1081 , \1082 , \1083 , \1084 ,
         \1085 , \1086 , \1087 , \1088 , \1089 , \1090 , \1091 , \1092 , \1093 , \1094 ,
         \1095 , \1096 , \1097 , \1098 , \1099 , \1100 , \1101 , \1102 , \1103 , \1104 ,
         \1105 , \1106 , \1107 , \1108 , \1109 , \1110 , \1111 , \1112 , \1113 , \1114 ,
         \1115 , \1116 , \1117 , \1118 , \1119 , \1120 , \1121 , \1122 , \1123 , \1124 ,
         \1125 , \1126 , \1127 , \1128 , \1129 , \1130 , \1131 , \1132 , \1133 , \1134 ,
         \1135 , \1136 , \1137 , \1138 , \1139 , \1140 , \1141 , \1142 , \1143 , \1144 ,
         \1145 , \1146 , \1147 , \1148 , \1149 , \1150 , \1151 , \1152 , \1153 , \1154 ,
         \1155 , \1156 , \1157 , \1158 , \1159 , \1160 , \1161 , \1162 , \1163 , \1164 ,
         \1165 , \1166 , \1167 , \1168 , \1169 , \1170 , \1171 , \1172 , \1173 , \1174 ,
         \1175 , \1176 , \1177 , \1178 , \1179 , \1180 , \1181 , \1182 , \1183 , \1184 ,
         \1185 , \1186 , \1187 , \1188 , \1189 , \1190 , \1191 , \1192 , \1193 , \1194 ,
         \1195 , \1196 , \1197 , \1198 , \1199 , \1200 , \1201 , \1202 , \1203 , \1204 ,
         \1205 , \1206 , \1207 , \1208 , \1209 , \1210 , \1211 , \1212 , \1213 , \1214 ,
         \1215 , \1216 , \1217 , \1218 , \1219 , \1220 , \1221 , \1222 , \1223 , \1224 ,
         \1225 , \1226 , \1227 , \1228 , \1229 , \1230 , \1231 , \1232 , \1233 , \1234 ,
         \1235 , \1236 , \1237 , \1238 , \1239 , \1240 , \1241 , \1242 , \1243 , \1244 ,
         \1245 , \1246 , \1247 , \1248 , \1249 , \1250 , \1251 , \1252 , \1253 , \1254 ,
         \1255 , \1256 , \1257 , \1258 , \1259 , \1260 , \1261 , \1262 , \1263 , \1264 ,
         \1265 , \1266 , \1267 , \1268 , \1269 , \1270 , \1271 , \1272 , \1273 , \1274 ,
         \1275 , \1276 , \1277 , \1278 , \1279 , \1280 , \1281 , \1282 , \1283 , \1284 ,
         \1285 , \1286 , \1287 , \1288 , \1289 , \1290 , \1291 , \1292 , \1293 , \1294 ,
         \1295 , \1296 , \1297 , \1298 , \1299 , \1300 , \1301 , \1302 , \1303 , \1304 ,
         \1305 , \1306 , \1307 , \1308 , \1309 , \1310 , \1311 , \1312 , \1313 , \1314 ,
         \1315 , \1316 , \1317 , \1318 , \1319 , \1320 , \1321 , \1322 , \1323 , \1324 ,
         \1325 , \1326 , \1327 , \1328 , \1329 , \1330 , \1331 , \1332 , \1333 , \1334 ,
         \1335 , \1336 , \1337 , \1338 , \1339 , \1340 , \1341 , \1342 , \1343 , \1344 ,
         \1345 , \1346 , \1347 , \1348 , \1349 , \1350 , \1351 , \1352 , \1353 , \1354 ,
         \1355 , \1356 , \1357 , \1358 , \1359 , \1360 , \1361 , \1362 , \1363 , \1364 ,
         \1365 , \1366 , \1367 , \1368 , \1369 , \1370 , \1371 , \1372 , \1373 , \1374 ,
         \1375 , \1376 , \1377 , \1378 , \1379 , \1380 , \1381 , \1382 , \1383 , \1384 ,
         \1385 , \1386 , \1387 , \1388 , \1389 , \1390 , \1391 , \1392 , \1393 , \1394 ,
         \1395 , \1396 , \1397 , \1398 , \1399 , \1400 , \1401 , \1402 , \1403 , \1404 ,
         \1405 , \1406 , \1407 , \1408 , \1409 , \1410 , \1411 , \1412 , \1413 , \1414 ,
         \1415 , \1416 , \1417 , \1418 , \1419 , \1420 , \1421 , \1422 , \1423 , \1424 ,
         \1425 , \1426 , \1427 , \1428 , \1429 , \1430 , \1431 , \1432 , \1433 , \1434 ,
         \1435 , \1436 , \1437 , \1438 , \1439 , \1440 , \1441 , \1442 , \1443 , \1444 ,
         \1445 , \1446 , \1447 , \1448 , \1449 , \1450 , \1451 , \1452 , \1453 , \1454 ,
         \1455 , \1456 , \1457 , \1458 , \1459 , \1460 , \1461 , \1462 , \1463 , \1464 ,
         \1465 , \1466 , \1467 , \1468 , \1469 , \1470 , \1471 , \1472 , \1473 , \1474 ,
         \1475 , \1476 , \1477 , \1478 , \1479 , \1480 , \1481 , \1482 , \1483 , \1484 ,
         \1485 , \1486 , \1487 , \1488 , \1489 , \1490 , \1491 , \1492 , \1493 , \1494 ,
         \1495 , \1496 , \1497 , \1498 , \1499 , \1500 , \1501 , \1502 , \1503 , \1504 ,
         \1505 , \1506 , \1507 , \1508 , \1509 , \1510 , \1511 , \1512 , \1513 , \1514 ,
         \1515 , \1516 , \1517 , \1518 , \1519 , \1520 , \1521 , \1522 , \1523 , \1524 ,
         \1525 , \1526 , \1527 , \1528 , \1529 , \1530 , \1531 , \1532 , \1533 , \1534 ,
         \1535 , \1536 , \1537 , \1538 , \1539 , \1540 , \1541 , \1542 , \1543 , \1544 ,
         \1545 , \1546 , \1547 , \1548 , \1549 , \1550 , \1551 , \1552 , \1553 , \1554 ,
         \1555 , \1556 , \1557 , \1558 , \1559 , \1560 , \1561 , \1562 , \1563 , \1564 ,
         \1565 , \1566 , \1567 , \1568 , \1569 , \1570 , \1571 , \1572 , \1573 , \1574 ,
         \1575 , \1576 , \1577 , \1578 , \1579 , \1580 , \1581 , \1582 , \1583 , \1584 ,
         \1585 , \1586 , \1587 , \1588 , \1589 , \1590 , \1591 , \1592 , \1593 , \1594 ,
         \1595 , \1596 , \1597 , \1598 , \1599 , \1600 , \1601 , \1602 , \1603 , \1604 ,
         \1605 , \1606 , \1607 , \1608 , \1609 , \1610 , \1611 , \1612 , \1613 , \1614 ,
         \1615 , \1616 , \1617 , \1618 , \1619 , \1620 , \1621 , \1622 , \1623 , \1624 ,
         \1625 , \1626 , \1627 , \1628 , \1629 , \1630 , \1631 , \1632 , \1633 , \1634 ,
         \1635 , \1636 , \1637 , \1638 , \1639 , \1640 , \1641 , \1642 , \1643 , \1644 ,
         \1645 , \1646 , \1647 , \1648 , \1649 , \1650 , \1651 , \1652 , \1653 , \1654 ,
         \1655 , \1656 , \1657 , \1658 , \1659 , \1660 , \1661 , \1662 , \1663 , \1664 ,
         \1665 , \1666 , \1667 , \1668 , \1669 , \1670 , \1671 , \1672 , \1673 , \1674 ,
         \1675 , \1676 , \1677 , \1678 , \1679 , \1680 , \1681 , \1682 , \1683 , \1684 ,
         \1685 , \1686 , \1687 , \1688 , \1689 , \1690 , \1691 , \1692 , \1693 , \1694 ,
         \1695 , \1696 , \1697 , \1698 , \1699 , \1700 , \1701 , \1702 , \1703 , \1704 ,
         \1705 , \1706 , \1707 , \1708 , \1709 , \1710 , \1711 , \1712 , \1713 , \1714 ,
         \1715 , \1716 , \1717 , \1718 , \1719 , \1720 , \1721 , \1722 , \1723 , \1724 ,
         \1725 , \1726 , \1727 , \1728 , \1729 , \1730 , \1731 , \1732 , \1733 , \1734 ,
         \1735 , \1736 , \1737 , \1738 , \1739 , \1740 , \1741 , \1742 , \1743 , \1744 ,
         \1745 , \1746 , \1747 , \1748 , \1749 , \1750 , \1751 , \1752 , \1753 , \1754 ,
         \1755 , \1756 , \1757 , \1758 , \1759 , \1760 , \1761 , \1762 , \1763 , \1764 ,
         \1765 , \1766 , \1767 , \1768 , \1769 , \1770 , \1771 , \1772 , \1773 , \1774 ,
         \1775 , \1776 , \1777 , \1778 , \1779 , \1780 , \1781 , \1782 , \1783 , \1784 ,
         \1785 , \1786 , \1787 , \1788 , \1789 , \1790 , \1791 , \1792 , \1793 , \1794 ,
         \1795 , \1796 , \1797 , \1798 , \1799 , \1800 , \1801 , \1802 , \1803 , \1804 ,
         \1805 , \1806 , \1807 , \1808 , \1809 , \1810 , \1811 , \1812 , \1813 , \1814 ,
         \1815 , \1816 , \1817 , \1818 , \1819 , \1820 , \1821 , \1822 , \1823 , \1824 ,
         \1825 , \1826 , \1827 , \1828 , \1829 , \1830 , \1831 , \1832 , \1833 , \1834 ,
         \1835 , \1836 , \1837 , \1838 , \1839 , \1840 , \1841 , \1842 , \1843 , \1844 ,
         \1845 , \1846 , \1847 , \1848 , \1849 , \1850 , \1851 , \1852 , \1853 , \1854 ,
         \1855 , \1856 , \1857 , \1858 , \1859 , \1860 , \1861 , \1862 , \1863 , \1864 ,
         \1865 , \1866 , \1867 , \1868 , \1869 , \1870 , \1871 , \1872 , \1873 , \1874 ,
         \1875 , \1876 , \1877 , \1878 , \1879 , \1880 , \1881 , \1882 , \1883 , \1884 ,
         \1885 , \1886 , \1887 , \1888 , \1889 , \1890 , \1891 , \1892 , \1893 , \1894 ,
         \1895 , \1896 , \1897 , \1898 , \1899 , \1900 , \1901 , \1902 , \1903 , \1904 ,
         \1905 , \1906 , \1907 , \1908 , \1909 , \1910 , \1911 , \1912 , \1913 , \1914 ,
         \1915 , \1916 , \1917 , \1918 , \1919 , \1920 , \1921 , \1922 , \1923 , \1924 ,
         \1925 , \1926 , \1927 , \1928 , \1929 , \1930 , \1931 , \1932 , \1933 , \1934 ,
         \1935 , \1936 , \1937 , \1938 , \1939 , \1940 , \1941 , \1942 , \1943 , \1944 ,
         \1945 , \1946 , \1947 , \1948 , \1949 , \1950 , \1951 , \1952 , \1953 , \1954 ,
         \1955 , \1956 , \1957 , \1958 , \1959 , \1960 , \1961 , \1962 , \1963 , \1964 ,
         \1965 , \1966 , \1967 , \1968 , \1969 , \1970 , \1971 , \1972 , \1973 , \1974 ,
         \1975 , \1976 , \1977 , \1978 , \1979 , \1980 , \1981 , \1982 , \1983 , \1984 ,
         \1985 , \1986 , \1987 , \1988 , \1989 , \1990 , \1991 , \1992 , \1993 , \1994 ,
         \1995 , \1996 , \1997 , \1998 , \1999 , \2000 , \2001 , \2002 , \2003 , \2004 ,
         \2005 , \2006 , \2007 , \2008 , \2009 , \2010 , \2011 , \2012 , \2013 , \2014 ,
         \2015 , \2016 , \2017 , \2018 , \2019 , \2020 , \2021 , \2022 , \2023 , \2024 ,
         \2025 , \2026 , \2027 , \2028 , \2029 , \2030 , \2031 , \2032 , \2033 , \2034 ,
         \2035 , \2036 , \2037 , \2038 , \2039 , \2040 , \2041 , \2042 , \2043 , \2044 ,
         \2045 , \2046 , \2047 , \2048 , \2049 , \2050 , \2051 , \2052 , \2053 , \2054 ,
         \2055 , \2056 , \2057 , \2058 , \2059 , \2060 , \2061 , \2062 , \2063 , \2064 ,
         \2065 , \2066 , \2067 , \2068 , \2069 , \2070 , \2071 , \2072 , \2073 , \2074 ,
         \2075 , \2076 , \2077 , \2078 , \2079 , \2080 , \2081 , \2082 , \2083 , \2084 ,
         \2085 , \2086 , \2087 , \2088 , \2089 , \2090 , \2091 , \2092 , \2093 , \2094 ,
         \2095 , \2096 , \2097 , \2098 , \2099 , \2100 , \2101 , \2102 , \2103 , \2104 ,
         \2105 , \2106 , \2107 , \2108 , \2109 , \2110 , \2111 , \2112 , \2113 , \2114 ,
         \2115 , \2116 , \2117 , \2118 , \2119 , \2120 , \2121 , \2122 , \2123 , \2124 ,
         \2125 , \2126 , \2127 , \2128 , \2129 , \2130 , \2131 , \2132 , \2133 , \2134 ,
         \2135 , \2136 , \2137 , \2138 , \2139 , \2140 , \2141 , \2142 , \2143 , \2144 ,
         \2145 , \2146 , \2147 , \2148 , \2149 , \2150 , \2151 , \2152 , \2153 , \2154 ,
         \2155 , \2156 , \2157 , \2158 , \2159 , \2160 , \2161 , \2162 , \2163 , \2164 ,
         \2165 , \2166 , \2167 , \2168 , \2169 , \2170 , \2171 , \2172 , \2173 , \2174 ,
         \2175 , \2176 , \2177 , \2178 , \2179 , \2180 , \2181 , \2182 , \2183 , \2184 ,
         \2185 , \2186 , \2187 , \2188 , \2189 , \2190 , \2191 , \2192 , \2193 , \2194 ,
         \2195 , \2196 , \2197 , \2198 , \2199 , \2200 , \2201 , \2202 , \2203 , \2204 ,
         \2205 , \2206 , \2207 , \2208 , \2209 , \2210 , \2211 , \2212 , \2213 , \2214 ,
         \2215 , \2216 , \2217 , \2218 , \2219 , \2220 , \2221 , \2222 , \2223 , \2224 ,
         \2225 , \2226 , \2227 , \2228 , \2229 , \2230 , \2231 , \2232 , \2233 , \2234 ,
         \2235 , \2236 , \2237 , \2238 , \2239 , \2240 , \2241 , \2242 , \2243 , \2244 ,
         \2245 , \2246 , \2247 , \2248 , \2249 , \2250 , \2251 , \2252 , \2253 , \2254 ,
         \2255 , \2256 , \2257 , \2258 , \2259 , \2260 , \2261 , \2262 , \2263 , \2264 ,
         \2265 , \2266 , \2267 , \2268 , \2269 , \2270 , \2271 , \2272 , \2273 , \2274 ,
         \2275 , \2276 , \2277 , \2278 , \2279 , \2280 , \2281 , \2282 , \2283 , \2284 ,
         \2285 , \2286 , \2287 , \2288 , \2289 , \2290 , \2291 , \2292 , \2293 , \2294 ,
         \2295 , \2296 , \2297 , \2298 , \2299 , \2300 , \2301 , \2302 , \2303 , \2304 ,
         \2305 , \2306 , \2307 , \2308 , \2309 , \2310 , \2311 , \2312 , \2313 , \2314 ,
         \2315 , \2316 , \2317 , \2318 , \2319 , \2320 , \2321 , \2322 , \2323 , \2324 ,
         \2325 , \2326 , \2327 , \2328 , \2329 , \2330 , \2331 , \2332 , \2333 , \2334 ,
         \2335 , \2336 , \2337 , \2338 , \2339 , \2340 , \2341 , \2342 , \2343 , \2344 ,
         \2345 , \2346 , \2347 , \2348 , \2349 , \2350 , \2351 , \2352 , \2353 , \2354 ,
         \2355 , \2356 , \2357 , \2358 , \2359 , \2360 , \2361 , \2362 , \2363 , \2364 ,
         \2365 , \2366 , \2367 , \2368 , \2369 , \2370 , \2371 , \2372 , \2373 , \2374 ,
         \2375 , \2376 , \2377 , \2378 , \2379 , \2380 , \2381 , \2382 , \2383 , \2384 ,
         \2385 , \2386 , \2387 , \2388 , \2389 , \2390 , \2391 , \2392 , \2393 , \2394 ,
         \2395 , \2396 , \2397 , \2398 , \2399 , \2400 , \2401 , \2402 , \2403 , \2404 ,
         \2405 , \2406 , \2407 , \2408 , \2409 , \2410 , \2411 , \2412 , \2413 , \2414 ,
         \2415 , \2416 , \2417 , \2418 , \2419 , \2420 , \2421 , \2422 , \2423 , \2424 ,
         \2425 , \2426 , \2427 , \2428 , \2429 , \2430 , \2431 , \2432 , \2433 , \2434 ,
         \2435 , \2436 , \2437 , \2438 , \2439 , \2440 , \2441 , \2442 , \2443 , \2444 ,
         \2445 , \2446 , \2447 , \2448 , \2449 , \2450 , \2451 , \2452 , \2453 , \2454 ,
         \2455 , \2456 , \2457 , \2458 , \2459 , \2460 , \2461 , \2462 , \2463 , \2464 ,
         \2465 , \2466 , \2467 , \2468 , \2469 , \2470 , \2471 , \2472 , \2473 , \2474 ,
         \2475 , \2476 , \2477 , \2478 , \2479 , \2480 , \2481 , \2482 , \2483 , \2484 ,
         \2485 , \2486 , \2487 , \2488 , \2489 , \2490 , \2491 , \2492 , \2493 , \2494 ,
         \2495 , \2496 , \2497 , \2498 , \2499 , \2500 , \2501 , \2502 , \2503 , \2504 ,
         \2505 , \2506 , \2507 , \2508 , \2509 , \2510 , \2511 , \2512 , \2513 , \2514 ,
         \2515 , \2516 , \2517 , \2518 , \2519 , \2520 , \2521 , \2522 , \2523 , \2524 ,
         \2525 , \2526 , \2527 , \2528 , \2529 , \2530 , \2531 , \2532 , \2533 , \2534 ,
         \2535 , \2536 , \2537 , \2538 , \2539 , \2540 , \2541 , \2542 , \2543 , \2544 ,
         \2545 , \2546 , \2547 , \2548 , \2549 , \2550 , \2551 , \2552 , \2553 , \2554 ,
         \2555 , \2556 , \2557 , \2558 , \2559 , \2560 , \2561 , \2562 , \2563 , \2564 ,
         \2565 , \2566 , \2567 , \2568 , \2569 , \2570 , \2571 , \2572 , \2573 , \2574 ,
         \2575 , \2576 , \2577 , \2578 , \2579 , \2580 , \2581 , \2582 , \2583 , \2584 ,
         \2585 , \2586 , \2587 , \2588 , \2589 , \2590 , \2591 , \2592 , \2593 , \2594 ,
         \2595 , \2596 , \2597 , \2598 , \2599 , \2600 , \2601 , \2602 , \2603 , \2604 ,
         \2605 , \2606 , \2607 , \2608 , \2609 , \2610 , \2611 , \2612 , \2613 , \2614 ,
         \2615 , \2616 , \2617 , \2618 , \2619 , \2620 , \2621 , \2622 , \2623 , \2624 ,
         \2625 , \2626 , \2627 , \2628 , \2629 , \2630 , \2631 , \2632 , \2633 , \2634 ,
         \2635 , \2636 , \2637 , \2638 , \2639 , \2640 , \2641 , \2642 , \2643 , \2644 ,
         \2645 , \2646 , \2647 , \2648 , \2649 , \2650 , \2651 , \2652 , \2653 , \2654 ,
         \2655 , \2656 , \2657 , \2658 , \2659 , \2660 , \2661 , \2662 , \2663 , \2664 ,
         \2665 , \2666 , \2667 , \2668 , \2669 , \2670 , \2671 , \2672 , \2673 , \2674 ,
         \2675 , \2676 , \2677 , \2678 , \2679 , \2680 , \2681 , \2682 , \2683 , \2684 ,
         \2685 , \2686 , \2687 , \2688 , \2689 , \2690 , \2691 , \2692 , \2693 , \2694 ,
         \2695 , \2696 , \2697 , \2698 , \2699 , \2700 , \2701 , \2702 , \2703 , \2704 ,
         \2705 , \2706 , \2707 , \2708 , \2709 , \2710 , \2711 , \2712 , \2713 , \2714 ,
         \2715 , \2716 , \2717 , \2718 , \2719 , \2720 , \2721 , \2722 , \2723 , \2724 ,
         \2725 , \2726 , \2727 , \2728 , \2729 , \2730 , \2731 , \2732 , \2733 , \2734 ,
         \2735 , \2736 , \2737 , \2738 , \2739 , \2740 , \2741 , \2742 , \2743 , \2744 ,
         \2745 , \2746 , \2747 , \2748 , \2749 , \2750 , \2751 , \2752 , \2753 , \2754 ,
         \2755 , \2756 , \2757 , \2758 , \2759 , \2760 , \2761 , \2762 , \2763 , \2764 ,
         \2765 , \2766 , \2767 , \2768 , \2769 , \2770 , \2771 , \2772 , \2773 , \2774 ,
         \2775 , \2776 , \2777 , \2778 , \2779 , \2780 , \2781 , \2782 , \2783 , \2784 ,
         \2785 , \2786 , \2787 , \2788 , \2789 , \2790 , \2791 , \2792 , \2793 , \2794 ,
         \2795 , \2796 , \2797 , \2798 , \2799 , \2800 , \2801 , \2802 , \2803 , \2804 ,
         \2805 , \2806 , \2807 , \2808 , \2809 , \2810 , \2811 , \2812 , \2813 , \2814 ,
         \2815 , \2816 , \2817 , \2818 , \2819 , \2820 , \2821 , \2822 , \2823 , \2824 ,
         \2825 , \2826 , \2827 , \2828 , \2829 , \2830 , \2831 , \2832 , \2833 , \2834 ,
         \2835 , \2836 , \2837 , \2838 , \2839 , \2840 , \2841 , \2842 , \2843 , \2844 ,
         \2845 , \2846 , \2847 , \2848 , \2849 , \2850 , \2851 , \2852 , \2853 , \2854 ,
         \2855 , \2856 , \2857 , \2858 , \2859 , \2860 , \2861 , \2862 , \2863 , \2864 ,
         \2865 , \2866 , \2867 , \2868 , \2869 , \2870 , \2871 , \2872 , \2873 , \2874 ,
         \2875 , \2876 , \2877 , \2878 , \2879 , \2880 , \2881 , \2882 , \2883 , \2884 ,
         \2885 , \2886 , \2887 , \2888 , \2889 , \2890 , \2891 , \2892 , \2893 , \2894 ,
         \2895 , \2896 , \2897 , \2898 , \2899 , \2900 , \2901 , \2902 , \2903 , \2904 ,
         \2905 , \2906 , \2907 , \2908 , \2909 , \2910 , \2911 , \2912 , \2913 , \2914 ,
         \2915 , \2916 , \2917 , \2918 , \2919 , \2920 , \2921 , \2922 , \2923 , \2924 ,
         \2925 , \2926 , \2927 , \2928 , \2929 , \2930 , \2931 , \2932 , \2933 , \2934 ,
         \2935 , \2936 , \2937 , \2938 , \2939 , \2940 , \2941 , \2942 , \2943 , \2944 ,
         \2945 , \2946 , \2947 , \2948 , \2949 , \2950 , \2951 , \2952 , \2953 , \2954 ,
         \2955 , \2956 , \2957 , \2958 , \2959 , \2960 , \2961 , \2962 , \2963 , \2964 ,
         \2965 , \2966 , \2967 , \2968 , \2969 , \2970 , \2971 , \2972 , \2973 , \2974 ,
         \2975 , \2976 , \2977 , \2978 , \2979 , \2980 , \2981 , \2982 , \2983 , \2984 ,
         \2985 , \2986 , \2987 , \2988 , \2989 , \2990 , \2991 , \2992 , \2993 , \2994 ,
         \2995 , \2996 , \2997 , \2998 , \2999 , \3000 , \3001 , \3002 , \3003 , \3004 ,
         \3005 , \3006 , \3007 , \3008 , \3009 , \3010 , \3011 , \3012 , \3013 , \3014 ,
         \3015 , \3016 , \3017 , \3018 , \3019 , \3020 , \3021 , \3022 , \3023 , \3024 ,
         \3025 , \3026 , \3027 , \3028 , \3029 , \3030 , \3031 , \3032 , \3033 , \3034 ,
         \3035 , \3036 , \3037 , \3038 , \3039 , \3040 , \3041 , \3042 , \3043 , \3044 ,
         \3045 , \3046 , \3047 , \3048 , \3049 , \3050 , \3051 , \3052 , \3053 , \3054 ,
         \3055 , \3056 , \3057 , \3058 , \3059 , \3060 , \3061 , \3062 , \3063 , \3064 ,
         \3065 , \3066 , \3067 , \3068 , \3069 , \3070 , \3071 , \3072 , \3073 , \3074 ,
         \3075 , \3076 , \3077 , \3078 , \3079 , \3080 , \3081 , \3082 , \3083 , \3084 ,
         \3085 , \3086 , \3087 , \3088 , \3089 , \3090 , \3091 , \3092 , \3093 , \3094 ,
         \3095 , \3096 , \3097 , \3098 , \3099 , \3100 , \3101 , \3102 , \3103 , \3104 ,
         \3105 , \3106 , \3107 , \3108 , \3109 , \3110 , \3111 , \3112 , \3113 , \3114 ,
         \3115 , \3116 , \3117 , \3118 , \3119 , \3120 , \3121 , \3122 , \3123 , \3124 ,
         \3125 , \3126 , \3127 , \3128 , \3129 , \3130 , \3131 , \3132 , \3133 , \3134 ,
         \3135 , \3136 , \3137 , \3138 , \3139 , \3140 , \3141 , \3142 , \3143 , \3144 ,
         \3145 , \3146 , \3147 , \3148 , \3149 , \3150 , \3151 , \3152 , \3153 , \3154 ,
         \3155 , \3156 , \3157 , \3158 , \3159 , \3160 , \3161 , \3162 , \3163 , \3164 ,
         \3165 , \3166 , \3167 , \3168 , \3169 , \3170 , \3171 , \3172 , \3173 , \3174 ,
         \3175 , \3176 , \3177 , \3178 , \3179 , \3180 , \3181 , \3182 , \3183 , \3184 ,
         \3185 , \3186 , \3187 , \3188 , \3189 , \3190 , \3191 , \3192 , \3193 , \3194 ,
         \3195 , \3196 , \3197 , \3198 , \3199 , \3200 , \3201 , \3202 , \3203 , \3204 ,
         \3205 , \3206 , \3207 , \3208 , \3209 , \3210 , \3211 , \3212 , \3213 , \3214 ,
         \3215 , \3216 , \3217 , \3218 , \3219 , \3220 , \3221 , \3222 , \3223 , \3224 ,
         \3225 , \3226 , \3227 , \3228 , \3229 , \3230 , \3231 , \3232 , \3233 , \3234 ,
         \3235 , \3236 , \3237 , \3238 , \3239 , \3240 , \3241 , \3242 , \3243 , \3244 ,
         \3245 , \3246 , \3247 , \3248 , \3249 , \3250 , \3251 , \3252 , \3253 , \3254 ,
         \3255 , \3256 , \3257 , \3258 , \3259 , \3260 , \3261 , \3262 , \3263 , \3264 ,
         \3265 , \3266 , \3267 , \3268 , \3269 , \3270 , \3271 , \3272 , \3273 , \3274 ,
         \3275 , \3276 , \3277 , \3278 , \3279 , \3280 , \3281 , \3282 , \3283 , \3284 ,
         \3285 , \3286 , \3287 , \3288 , \3289 , \3290 , \3291 , \3292 , \3293 , \3294 ,
         \3295 , \3296 , \3297 , \3298 , \3299 , \3300 , \3301 , \3302 , \3303 , \3304 ,
         \3305 , \3306 , \3307 , \3308 , \3309 , \3310 , \3311 , \3312 , \3313 , \3314 ,
         \3315 , \3316 , \3317 , \3318 , \3319 , \3320 , \3321 , \3322 , \3323 , \3324 ,
         \3325 , \3326 , \3327 , \3328 , \3329 , \3330 , \3331 , \3332 , \3333 , \3334 ,
         \3335 , \3336 , \3337 , \3338 , \3339 , \3340 , \3341 , \3342 , \3343 , \3344 ,
         \3345 , \3346 , \3347 , \3348 , \3349 , \3350 , \3351 , \3352 , \3353 , \3354 ,
         \3355 , \3356 , \3357 , \3358 , \3359 , \3360 , \3361 , \3362 , \3363 , \3364 ,
         \3365 , \3366 , \3367 , \3368 , \3369 , \3370 , \3371 , \3372 , \3373 , \3374 ,
         \3375 , \3376 , \3377 , \3378 , \3379 , \3380 , \3381 , \3382 , \3383 , \3384 ,
         \3385 , \3386 , \3387 , \3388 , \3389 , \3390 , \3391 , \3392 , \3393 , \3394 ,
         \3395 , \3396 , \3397 , \3398 , \3399 , \3400 , \3401 , \3402 , \3403 , \3404 ,
         \3405 , \3406 , \3407 , \3408 , \3409 , \3410 , \3411 , \3412 , \3413 , \3414 ,
         \3415 , \3416 , \3417 , \3418 , \3419 , \3420 , \3421 , \3422 , \3423 , \3424 ,
         \3425 , \3426 , \3427 , \3428 , \3429 , \3430 , \3431 , \3432 , \3433 , \3434 ,
         \3435 , \3436 , \3437 , \3438 , \3439 , \3440 , \3441 , \3442 , \3443 , \3444 ,
         \3445 , \3446 , \3447 , \3448 , \3449 , \3450 , \3451 , \3452 , \3453 , \3454 ,
         \3455 , \3456 , \3457 , \3458 , \3459 , \3460 , \3461 , \3462 , \3463 , \3464 ,
         \3465 , \3466 , \3467 , \3468 , \3469 , \3470 , \3471 , \3472 , \3473 , \3474 ,
         \3475 , \3476 , \3477 , \3478 , \3479 , \3480 , \3481 , \3482 , \3483 , \3484 ,
         \3485 , \3486 , \3487 , \3488 , \3489 , \3490 , \3491 , \3492 , \3493 , \3494 ,
         \3495 , \3496 , \3497 , \3498 , \3499 , \3500 , \3501 , \3502 , \3503 , \3504 ,
         \3505 , \3506 , \3507 , \3508 , \3509 , \3510 , \3511 , \3512 , \3513 , \3514 ,
         \3515 , \3516 , \3517 , \3518 , \3519 , \3520 , \3521 , \3522 , \3523 , \3524 ,
         \3525 , \3526 , \3527 , \3528 , \3529 , \3530 , \3531 , \3532 , \3533 , \3534 ,
         \3535 , \3536 , \3537 , \3538 , \3539 , \3540 , \3541 , \3542 , \3543 , \3544 ,
         \3545 , \3546 , \3547 , \3548 , \3549 , \3550 , \3551 , \3552 , \3553 , \3554 ,
         \3555 , \3556 , \3557 , \3558 , \3559 , \3560 , \3561 , \3562 , \3563 , \3564 ,
         \3565 , \3566 , \3567 , \3568 , \3569 , \3570 , \3571 , \3572 , \3573 , \3574 ,
         \3575 , \3576 , \3577 , \3578 , \3579 , \3580 , \3581 , \3582 , \3583 , \3584 ,
         \3585 , \3586 , \3587 , \3588 , \3589 , \3590 , \3591 , \3592 , \3593 , \3594 ,
         \3595 , \3596 , \3597 , \3598 , \3599 , \3600 , \3601 , \3602 , \3603 , \3604 ,
         \3605 , \3606 , \3607 , \3608 , \3609 , \3610 , \3611 , \3612 , \3613 , \3614 ,
         \3615 , \3616 , \3617 , \3618 , \3619 , \3620 , \3621 , \3622 , \3623 , \3624 ,
         \3625 , \3626 , \3627 , \3628 , \3629 , \3630 , \3631 , \3632 , \3633 , \3634 ,
         \3635 , \3636 , \3637 , \3638 , \3639 , \3640 , \3641 , \3642 , \3643 , \3644 ,
         \3645 , \3646 , \3647 , \3648 , \3649 , \3650 , \3651 , \3652 , \3653 , \3654 ,
         \3655 , \3656 , \3657 , \3658 , \3659 , \3660 , \3661 , \3662 , \3663 , \3664 ,
         \3665 , \3666 , \3667 , \3668 , \3669 , \3670 , \3671 , \3672 , \3673 , \3674 ,
         \3675 , \3676 , \3677 , \3678 , \3679 , \3680 , \3681 , \3682 , \3683 , \3684 ,
         \3685 , \3686 , \3687 , \3688 , \3689 , \3690 , \3691 , \3692 , \3693 , \3694 ,
         \3695 , \3696 , \3697 , \3698 , \3699 , \3700 , \3701 , \3702 , \3703 , \3704 ,
         \3705 , \3706 , \3707 , \3708 , \3709 , \3710 , \3711 , \3712 , \3713 , \3714 ,
         \3715 , \3716 , \3717 , \3718 , \3719 , \3720 , \3721 , \3722 , \3723 , \3724 ,
         \3725 , \3726 , \3727 , \3728 , \3729 , \3730 , \3731 , \3732 , \3733 , \3734 ,
         \3735 , \3736 , \3737 , \3738 , \3739 , \3740 , \3741 , \3742 , \3743 , \3744 ,
         \3745 , \3746 , \3747 , \3748 , \3749 , \3750 , \3751 , \3752 , \3753 , \3754 ,
         \3755 , \3756 , \3757 , \3758 , \3759 , \3760 , \3761 , \3762 , \3763 , \3764 ,
         \3765 , \3766 , \3767 , \3768 , \3769 , \3770 , \3771 , \3772 , \3773 , \3774 ,
         \3775 , \3776 , \3777 , \3778 , \3779 , \3780 , \3781 , \3782 , \3783 , \3784 ,
         \3785 , \3786 , \3787 , \3788 , \3789 , \3790 , \3791 , \3792 , \3793 , \3794 ,
         \3795 , \3796 , \3797 , \3798 , \3799 , \3800 , \3801 , \3802 , \3803 , \3804 ,
         \3805 , \3806 , \3807 , \3808 , \3809 , \3810 , \3811 , \3812 , \3813 , \3814 ,
         \3815 , \3816 , \3817 , \3818 , \3819 , \3820 , \3821 , \3822 , \3823 , \3824 ,
         \3825 , \3826 , \3827 , \3828 , \3829 , \3830 , \3831 , \3832 , \3833 , \3834 ,
         \3835 , \3836 , \3837 , \3838 , \3839 , \3840 , \3841 , \3842 , \3843 , \3844 ,
         \3845 , \3846 , \3847 , \3848 , \3849 , \3850 , \3851 , \3852 , \3853 , \3854 ,
         \3855 , \3856 , \3857 , \3858 , \3859 , \3860 , \3861 , \3862 , \3863 , \3864 ,
         \3865 , \3866 , \3867 , \3868 , \3869 , \3870 , \3871 , \3872 , \3873 , \3874 ,
         \3875 , \3876 , \3877 , \3878 , \3879 , \3880 , \3881 , \3882 , \3883 , \3884 ,
         \3885 , \3886 , \3887 , \3888 , \3889 , \3890 , \3891 , \3892 , \3893 , \3894 ,
         \3895 , \3896 , \3897 , \3898 , \3899 , \3900 , \3901 , \3902 , \3903 , \3904 ,
         \3905 , \3906 , \3907 , \3908 , \3909 , \3910 , \3911 , \3912 , \3913 , \3914 ,
         \3915 , \3916 , \3917 , \3918 , \3919 , \3920 , \3921 , \3922 , \3923 , \3924 ,
         \3925 , \3926 , \3927 , \3928 , \3929 , \3930 , \3931 , \3932 , \3933 , \3934 ,
         \3935 , \3936 , \3937 , \3938 , \3939 , \3940 , \3941 , \3942 , \3943 , \3944 ,
         \3945 , \3946 , \3947 , \3948 , \3949 , \3950 , \3951 , \3952 , \3953 , \3954 ,
         \3955 , \3956 , \3957 , \3958 , \3959 , \3960 , \3961 , \3962 , \3963 , \3964 ,
         \3965 , \3966 , \3967 , \3968 , \3969 , \3970 , \3971 , \3972 , \3973 , \3974 ,
         \3975 , \3976 , \3977 , \3978 , \3979 , \3980 , \3981 , \3982 , \3983 , \3984 ,
         \3985 , \3986 , \3987 , \3988 , \3989 , \3990 , \3991 , \3992 , \3993 , \3994 ,
         \3995 , \3996 , \3997 , \3998 , \3999 , \4000 , \4001 , \4002 , \4003 , \4004 ,
         \4005 , \4006 , \4007 , \4008 , \4009 , \4010 , \4011 , \4012 , \4013 , \4014 ,
         \4015 , \4016 , \4017 , \4018 , \4019 , \4020 , \4021 , \4022 , \4023 , \4024 ,
         \4025 , \4026 , \4027 , \4028 , \4029 , \4030 , \4031 , \4032 , \4033 , \4034 ,
         \4035 , \4036 , \4037 , \4038 , \4039 , \4040 , \4041 , \4042 , \4043 , \4044 ,
         \4045 , \4046 , \4047 , \4048 , \4049 , \4050 , \4051 , \4052 , \4053 , \4054 ,
         \4055 , \4056 , \4057 , \4058 , \4059 , \4060 , \4061 , \4062 , \4063 , \4064 ,
         \4065 , \4066 , \4067 , \4068 , \4069 , \4070 , \4071 , \4072 , \4073 , \4074 ,
         \4075 , \4076 , \4077 , \4078 , \4079 , \4080 , \4081 , \4082 , \4083 , \4084 ,
         \4085 , \4086 , \4087 , \4088 , \4089 , \4090 , \4091 , \4092 , \4093 , \4094 ,
         \4095 , \4096 , \4097 , \4098 , \4099 , \4100 , \4101 , \4102 , \4103 , \4104 ,
         \4105 , \4106 , \4107 , \4108 , \4109 , \4110 , \4111 , \4112 , \4113 , \4114 ,
         \4115 , \4116 , \4117 , \4118 , \4119 , \4120 , \4121 , \4122 , \4123 , \4124 ,
         \4125 , \4126 , \4127 , \4128 , \4129 , \4130 , \4131 , \4132 , \4133 , \4134 ,
         \4135 , \4136 , \4137 , \4138 , \4139 , \4140 , \4141 , \4142 , \4143 , \4144 ,
         \4145 , \4146 , \4147 , \4148 , \4149 , \4150 , \4151 , \4152 , \4153 , \4154 ,
         \4155 , \4156 , \4157 , \4158 , \4159 , \4160 , \4161 , \4162 , \4163 , \4164 ,
         \4165 , \4166 , \4167 , \4168 , \4169 , \4170 , \4171 , \4172 , \4173 , \4174 ,
         \4175 , \4176 , \4177 , \4178 , \4179 , \4180 , \4181 , \4182 , \4183 , \4184 ,
         \4185 , \4186 , \4187 , \4188 , \4189 , \4190 , \4191 , \4192 , \4193 , \4194 ,
         \4195 , \4196 , \4197 , \4198 , \4199 , \4200 , \4201 , \4202 , \4203 , \4204 ,
         \4205 , \4206 , \4207 , \4208 , \4209 , \4210 , \4211 , \4212 , \4213 , \4214 ,
         \4215 , \4216 , \4217 , \4218 , \4219 , \4220 , \4221 , \4222 , \4223 , \4224 ,
         \4225 , \4226 , \4227 , \4228 , \4229 , \4230 , \4231 , \4232 , \4233 , \4234 ,
         \4235 , \4236 , \4237 , \4238 , \4239 , \4240 , \4241 , \4242 , \4243 , \4244 ,
         \4245 , \4246 , \4247 , \4248 , \4249 , \4250 , \4251 , \4252 , \4253 , \4254 ,
         \4255 , \4256 , \4257 , \4258 , \4259 , \4260 , \4261 , \4262 , \4263 , \4264 ,
         \4265 , \4266 , \4267 , \4268 , \4269 , \4270 , \4271 , \4272 , \4273 , \4274 ,
         \4275 , \4276 , \4277 , \4278 , \4279 , \4280 , \4281 , \4282 , \4283 , \4284 ,
         \4285 , \4286 , \4287 , \4288 , \4289 , \4290 , \4291 , \4292 , \4293 , \4294 ,
         \4295 , \4296 , \4297 , \4298 , \4299 , \4300 , \4301 , \4302 , \4303 , \4304 ,
         \4305 , \4306 , \4307 , \4308 , \4309 , \4310 , \4311 , \4312 , \4313 , \4314 ,
         \4315 , \4316 , \4317 , \4318 , \4319 , \4320 , \4321 , \4322 , \4323 , \4324 ,
         \4325 , \4326 , \4327 , \4328 , \4329 , \4330 , \4331 , \4332 , \4333 , \4334 ,
         \4335 , \4336 , \4337 , \4338 , \4339 , \4340 , \4341 , \4342 , \4343 , \4344 ,
         \4345 , \4346 , \4347 , \4348 , \4349 , \4350 , \4351 , \4352 , \4353 , \4354 ,
         \4355 , \4356 , \4357 , \4358 , \4359 , \4360 , \4361 , \4362 , \4363 , \4364 ,
         \4365 , \4366 , \4367 , \4368 , \4369 , \4370 , \4371 , \4372 , \4373 , \4374 ,
         \4375 , \4376 , \4377 , \4378 , \4379 , \4380 , \4381 , \4382 , \4383 , \4384 ,
         \4385 , \4386 , \4387 , \4388 , \4389 , \4390 , \4391 , \4392 , \4393 , \4394 ,
         \4395 , \4396 , \4397 , \4398 , \4399 , \4400 , \4401 , \4402 , \4403 , \4404 ,
         \4405 , \4406 , \4407 , \4408 , \4409 , \4410 , \4411 , \4412 , \4413 , \4414 ,
         \4415 , \4416 , \4417 , \4418 , \4419 , \4420 , \4421 , \4422 , \4423 , \4424 ,
         \4425 , \4426 , \4427 , \4428 , \4429 , \4430 , \4431 , \4432 , \4433 , \4434 ,
         \4435 , \4436 , \4437 , \4438 , \4439 , \4440 , \4441 , \4442 , \4443 , \4444 ,
         \4445 , \4446 , \4447 , \4448 , \4449 , \4450 , \4451 , \4452 , \4453 , \4454 ,
         \4455 , \4456 , \4457 , \4458 , \4459 , \4460 , \4461 , \4462 , \4463 , \4464 ,
         \4465 , \4466 , \4467 , \4468 , \4469 , \4470 , \4471 , \4472 , \4473 , \4474 ,
         \4475 , \4476 , \4477 , \4478 , \4479 , \4480 , \4481 , \4482 , \4483 , \4484 ,
         \4485 , \4486 , \4487 , \4488 , \4489 , \4490 , \4491 , \4492 , \4493 , \4494 ,
         \4495 , \4496 , \4497 , \4498 , \4499 , \4500 , \4501 , \4502 , \4503 , \4504 ,
         \4505 , \4506 , \4507 , \4508 , \4509 , \4510 , \4511 , \4512 , \4513 , \4514 ,
         \4515 , \4516 , \4517 , \4518 , \4519 , \4520 , \4521 , \4522 , \4523 , \4524 ,
         \4525 , \4526 , \4527 , \4528 , \4529 , \4530 , \4531 , \4532 , \4533 , \4534 ,
         \4535 , \4536 , \4537 , \4538 , \4539 , \4540 , \4541 , \4542 , \4543 , \4544 ,
         \4545 , \4546 , \4547 , \4548 , \4549 , \4550 , \4551 , \4552 , \4553 , \4554 ,
         \4555 , \4556 , \4557 , \4558 , \4559 , \4560 , \4561 , \4562 , \4563 , \4564 ,
         \4565 , \4566 , \4567 , \4568 , \4569 , \4570 , \4571 , \4572 , \4573 , \4574 ,
         \4575 , \4576 , \4577 , \4578 , \4579 , \4580 , \4581 , \4582 , \4583 , \4584 ,
         \4585 , \4586 , \4587 , \4588 , \4589 , \4590 , \4591 , \4592 , \4593 , \4594 ,
         \4595 , \4596 , \4597 , \4598 , \4599 , \4600 , \4601 , \4602 , \4603 , \4604 ,
         \4605 , \4606 , \4607 , \4608 , \4609 , \4610 , \4611 , \4612 , \4613 , \4614 ,
         \4615 , \4616 , \4617 , \4618 , \4619 , \4620 , \4621 , \4622 , \4623 , \4624 ,
         \4625 , \4626 , \4627 , \4628 , \4629 , \4630 , \4631 , \4632 , \4633 , \4634 ,
         \4635 , \4636 , \4637 , \4638 , \4639 , \4640 , \4641 , \4642 , \4643 , \4644 ,
         \4645 , \4646 , \4647 , \4648 , \4649 , \4650 , \4651 , \4652 , \4653 , \4654 ,
         \4655 , \4656 , \4657 , \4658 , \4659 , \4660 , \4661 , \4662 , \4663 , \4664 ,
         \4665 , \4666 , \4667 , \4668 , \4669 , \4670 , \4671 , \4672 , \4673 , \4674 ,
         \4675 , \4676 , \4677 , \4678 , \4679 , \4680 , \4681 , \4682 , \4683 , \4684 ,
         \4685 , \4686 , \4687 , \4688 , \4689 , \4690 , \4691 , \4692 , \4693 , \4694 ,
         \4695 , \4696 , \4697 , \4698 , \4699 , \4700 , \4701 , \4702 , \4703 , \4704 ,
         \4705 , \4706 , \4707 , \4708 , \4709 , \4710 , \4711 , \4712 , \4713 , \4714 ,
         \4715 , \4716 , \4717 , \4718 , \4719 , \4720 , \4721 , \4722 , \4723 , \4724 ,
         \4725 , \4726 , \4727 , \4728 , \4729 , \4730 , \4731 , \4732 , \4733 , \4734 ,
         \4735 , \4736 , \4737 , \4738 , \4739 , \4740 , \4741 , \4742 , \4743 , \4744 ,
         \4745 , \4746 , \4747 , \4748 , \4749 , \4750 , \4751 , \4752 , \4753 , \4754 ,
         \4755 , \4756 , \4757 , \4758 , \4759 , \4760 , \4761 , \4762 , \4763 , \4764 ,
         \4765 , \4766 , \4767 , \4768 , \4769 , \4770 , \4771 , \4772 , \4773 , \4774 ,
         \4775 , \4776 , \4777 , \4778 , \4779 , \4780 , \4781 , \4782 , \4783 , \4784 ,
         \4785 , \4786 , \4787 , \4788 , \4789 , \4790 , \4791 , \4792 , \4793 , \4794 ,
         \4795 , \4796 , \4797 , \4798 , \4799 , \4800 , \4801 , \4802 , \4803 , \4804 ,
         \4805 , \4806 , \4807 , \4808 , \4809 , \4810 , \4811 , \4812 , \4813 , \4814 ,
         \4815 , \4816 , \4817 , \4818 , \4819 , \4820 , \4821 , \4822 , \4823 , \4824 ,
         \4825 , \4826 , \4827 , \4828 , \4829 , \4830 , \4831 , \4832 , \4833 , \4834 ,
         \4835 , \4836 , \4837 , \4838 , \4839 , \4840 , \4841 , \4842 , \4843 , \4844 ,
         \4845 , \4846 , \4847 , \4848 , \4849 , \4850 , \4851 , \4852 , \4853 , \4854 ,
         \4855 , \4856 , \4857 , \4858 , \4859 , \4860 , \4861 , \4862 , \4863 , \4864 ,
         \4865 , \4866 , \4867 , \4868 , \4869 , \4870 , \4871 , \4872 , \4873 , \4874 ,
         \4875 , \4876 , \4877 , \4878 , \4879 , \4880 , \4881 , \4882 , \4883 , \4884 ,
         \4885 , \4886 , \4887 , \4888 , \4889 , \4890 , \4891 , \4892 , \4893 , \4894 ,
         \4895 , \4896 , \4897 , \4898 , \4899 , \4900 , \4901 , \4902 , \4903 , \4904 ,
         \4905 , \4906 , \4907 , \4908 , \4909 , \4910 , \4911 , \4912 , \4913 , \4914 ,
         \4915 , \4916 , \4917 , \4918 , \4919 , \4920 , \4921 , \4922 , \4923 , \4924 ,
         \4925 , \4926 , \4927 , \4928 , \4929 , \4930 , \4931 , \4932 , \4933 , \4934 ,
         \4935 , \4936 , \4937 , \4938 , \4939 , \4940 , \4941 , \4942 , \4943 , \4944 ,
         \4945 , \4946 , \4947 , \4948 , \4949 , \4950 , \4951 , \4952 , \4953 , \4954 ,
         \4955 , \4956 , \4957 , \4958 , \4959 , \4960 , \4961 , \4962 , \4963 , \4964 ,
         \4965 , \4966 , \4967 , \4968 , \4969 , \4970 , \4971 , \4972 , \4973 , \4974 ,
         \4975 , \4976 , \4977 , \4978 , \4979 , \4980 , \4981 , \4982 , \4983 , \4984 ,
         \4985 , \4986 , \4987 , \4988 , \4989 , \4990 , \4991 , \4992 , \4993 , \4994 ,
         \4995 , \4996 , \4997 , \4998 , \4999 , \5000 , \5001 , \5002 , \5003 , \5004 ,
         \5005 , \5006 , \5007 , \5008 , \5009 , \5010 , \5011 , \5012 , \5013 , \5014 ,
         \5015 , \5016 , \5017 , \5018 , \5019 , \5020 , \5021 , \5022 , \5023 , \5024 ,
         \5025 , \5026 , \5027 , \5028 , \5029 , \5030 , \5031 , \5032 , \5033 , \5034 ,
         \5035 , \5036 , \5037 , \5038 , \5039 , \5040 , \5041 , \5042 , \5043 , \5044 ,
         \5045 , \5046 , \5047 , \5048 , \5049 , \5050 , \5051 , \5052 , \5053 , \5054 ,
         \5055 , \5056 , \5057 , \5058 , \5059 , \5060 , \5061 , \5062 , \5063 , \5064 ,
         \5065 , \5066 , \5067 , \5068 , \5069 , \5070 , \5071 , \5072 , \5073 , \5074 ,
         \5075 , \5076 , \5077 , \5078 , \5079 , \5080 , \5081 , \5082 , \5083 , \5084 ,
         \5085 , \5086 , \5087 , \5088 , \5089 , \5090 , \5091 , \5092 , \5093 , \5094 ,
         \5095 , \5096 , \5097 , \5098 , \5099 , \5100 , \5101 , \5102 , \5103 , \5104 ,
         \5105 , \5106 , \5107 , \5108 , \5109 , \5110 , \5111 , \5112 , \5113 , \5114 ,
         \5115 , \5116 , \5117 , \5118 , \5119 , \5120 , \5121 , \5122 , \5123 , \5124 ,
         \5125 , \5126 , \5127 , \5128 , \5129 , \5130 , \5131 , \5132 , \5133 , \5134 ,
         \5135 , \5136 , \5137 , \5138 , \5139 , \5140 , \5141 , \5142 , \5143 , \5144 ,
         \5145 , \5146 , \5147 , \5148 , \5149 , \5150 , \5151 , \5152 , \5153 , \5154 ,
         \5155 , \5156 , \5157 , \5158 , \5159 , \5160 , \5161 , \5162 , \5163 , \5164 ,
         \5165 , \5166 , \5167 , \5168 , \5169 , \5170 , \5171 , \5172 , \5173 , \5174 ,
         \5175 , \5176 , \5177 , \5178 , \5179 , \5180 , \5181 , \5182 , \5183 , \5184 ,
         \5185 , \5186 , \5187 , \5188 , \5189 , \5190 , \5191 , \5192 , \5193 , \5194 ,
         \5195 , \5196 , \5197 , \5198 , \5199 , \5200 , \5201 , \5202 , \5203 , \5204 ,
         \5205 , \5206 , \5207 , \5208 , \5209 , \5210 , \5211 , \5212 , \5213 , \5214 ,
         \5215 , \5216 , \5217 , \5218 , \5219 , \5220 , \5221 , \5222 , \5223 , \5224 ,
         \5225 , \5226 , \5227 , \5228 , \5229 , \5230 , \5231 , \5232 , \5233 , \5234 ,
         \5235 , \5236 , \5237 , \5238 , \5239 , \5240 , \5241 , \5242 , \5243 , \5244 ,
         \5245 , \5246 , \5247 , \5248 , \5249 , \5250 , \5251 , \5252 , \5253 , \5254 ,
         \5255 , \5256 , \5257 , \5258 , \5259 , \5260 , \5261 , \5262 , \5263 , \5264 ,
         \5265 , \5266 , \5267 , \5268 , \5269 , \5270 , \5271 , \5272 , \5273 , \5274 ,
         \5275 , \5276 , \5277 , \5278 , \5279 , \5280 , \5281 , \5282 , \5283 , \5284 ,
         \5285 , \5286 , \5287 , \5288 , \5289 , \5290 , \5291 , \5292 , \5293 , \5294 ,
         \5295 , \5296 , \5297 , \5298 , \5299 , \5300 , \5301 , \5302 , \5303 , \5304 ,
         \5305 , \5306 , \5307 , \5308 , \5309 , \5310 , \5311 , \5312 , \5313 , \5314 ,
         \5315 , \5316 , \5317 , \5318 , \5319 , \5320 , \5321 , \5322 , \5323 , \5324 ,
         \5325 , \5326 , \5327 , \5328 , \5329 , \5330 , \5331 , \5332 , \5333 , \5334 ,
         \5335 , \5336 , \5337 , \5338 , \5339 , \5340 , \5341 , \5342 , \5343 , \5344 ,
         \5345 , \5346 , \5347 , \5348 , \5349 , \5350 , \5351 , \5352 , \5353 , \5354 ,
         \5355 , \5356 , \5357 , \5358 , \5359 , \5360 , \5361 , \5362 , \5363 , \5364 ,
         \5365 , \5366 , \5367 , \5368 , \5369 , \5370 , \5371 , \5372 , \5373 , \5374 ,
         \5375 , \5376 , \5377 , \5378 , \5379 , \5380 , \5381 , \5382 , \5383 , \5384 ,
         \5385 , \5386 , \5387 , \5388 , \5389 , \5390 , \5391 , \5392 , \5393 , \5394 ,
         \5395 , \5396 , \5397 , \5398 , \5399 , \5400 , \5401 , \5402 , \5403 , \5404 ,
         \5405 , \5406 , \5407 , \5408 , \5409 , \5410 , \5411 , \5412 , \5413 , \5414 ,
         \5415 , \5416 , \5417 , \5418 , \5419 , \5420 , \5421 , \5422 , \5423 , \5424 ,
         \5425 , \5426 , \5427 , \5428 , \5429 , \5430 , \5431 , \5432 , \5433 , \5434 ,
         \5435 , \5436 , \5437 , \5438 , \5439 , \5440 , \5441 , \5442 , \5443 , \5444 ,
         \5445 , \5446 , \5447 , \5448 , \5449 , \5450 , \5451 , \5452 , \5453 , \5454 ,
         \5455 , \5456 , \5457 , \5458 , \5459 , \5460 , \5461 , \5462 , \5463 , \5464 ,
         \5465 , \5466 , \5467 , \5468 , \5469 , \5470 , \5471 , \5472 , \5473 , \5474 ,
         \5475 , \5476 , \5477 , \5478 , \5479 , \5480 , \5481 , \5482 , \5483 , \5484 ,
         \5485 , \5486 , \5487 , \5488 , \5489 , \5490 , \5491 , \5492 , \5493 , \5494 ,
         \5495 , \5496 , \5497 , \5498 , \5499 , \5500 , \5501 , \5502 , \5503 , \5504 ,
         \5505 , \5506 , \5507 , \5508 , \5509 , \5510 , \5511 , \5512 , \5513 , \5514 ,
         \5515 , \5516 , \5517 , \5518 , \5519 , \5520 , \5521 , \5522 , \5523 , \5524 ,
         \5525 , \5526 , \5527 , \5528 , \5529 , \5530 , \5531 , \5532 , \5533 , \5534 ,
         \5535 , \5536 , \5537 , \5538 , \5539 , \5540 , \5541 , \5542 , \5543 , \5544 ,
         \5545 , \5546 , \5547 , \5548 , \5549 , \5550 , \5551 , \5552 , \5553 , \5554 ,
         \5555 , \5556 , \5557 , \5558 , \5559 , \5560 , \5561 , \5562 , \5563 , \5564 ,
         \5565 , \5566 , \5567 , \5568 , \5569 , \5570 , \5571 , \5572 , \5573 , \5574 ,
         \5575 , \5576 , \5577 , \5578 , \5579 , \5580 , \5581 , \5582 , \5583 , \5584 ,
         \5585 , \5586 , \5587 , \5588 , \5589 , \5590 , \5591 , \5592 , \5593 , \5594 ,
         \5595 , \5596 , \5597 , \5598 , \5599 , \5600 , \5601 , \5602 , \5603 , \5604 ,
         \5605 , \5606 , \5607 , \5608 , \5609 , \5610 , \5611 , \5612 , \5613 , \5614 ,
         \5615 , \5616 , \5617 , \5618 , \5619 , \5620 , \5621 , \5622 , \5623 , \5624 ,
         \5625 , \5626 , \5627 , \5628 , \5629 , \5630 , \5631 , \5632 , \5633 , \5634 ,
         \5635 , \5636 , \5637 , \5638 , \5639 , \5640 , \5641 , \5642 , \5643 , \5644 ,
         \5645 , \5646 , \5647 , \5648 , \5649 , \5650 , \5651 , \5652 , \5653 , \5654 ,
         \5655 , \5656 , \5657 , \5658 , \5659 , \5660 , \5661 , \5662 , \5663 , \5664 ,
         \5665 , \5666 , \5667 , \5668 , \5669 , \5670 , \5671 , \5672 , \5673 , \5674 ,
         \5675 , \5676 , \5677 , \5678 , \5679 , \5680 , \5681 , \5682 , \5683 , \5684 ,
         \5685 , \5686 , \5687 , \5688 , \5689 , \5690 , \5691 , \5692 , \5693 , \5694 ,
         \5695 , \5696 , \5697 , \5698 , \5699 , \5700 , \5701 , \5702 , \5703 , \5704 ,
         \5705 , \5706 , \5707 , \5708 , \5709 , \5710 , \5711 , \5712 , \5713 , \5714 ,
         \5715 , \5716 , \5717 , \5718 , \5719 , \5720 , \5721 , \5722 , \5723 , \5724 ,
         \5725 , \5726 , \5727 , \5728 , \5729 , \5730 , \5731 , \5732 , \5733 , \5734 ,
         \5735 , \5736 , \5737 , \5738 , \5739 , \5740 , \5741 , \5742 , \5743 , \5744 ,
         \5745 , \5746 , \5747 , \5748 , \5749 , \5750 , \5751 , \5752 , \5753 , \5754 ,
         \5755 , \5756 , \5757 , \5758 , \5759 , \5760 , \5761 , \5762 , \5763 , \5764 ,
         \5765 , \5766 , \5767 , \5768 , \5769 , \5770 , \5771 , \5772 , \5773 , \5774 ,
         \5775 , \5776 , \5777 , \5778 , \5779 , \5780 , \5781 , \5782 , \5783 , \5784 ,
         \5785 , \5786 , \5787 , \5788 , \5789 , \5790 , \5791 , \5792 , \5793 , \5794 ,
         \5795 , \5796 , \5797 , \5798 , \5799 , \5800 , \5801 , \5802 , \5803 , \5804 ,
         \5805 , \5806 , \5807 , \5808 , \5809 , \5810 , \5811 , \5812 , \5813 , \5814 ,
         \5815 , \5816 , \5817 , \5818 , \5819 , \5820 , \5821 , \5822 , \5823 , \5824 ,
         \5825 , \5826 , \5827 , \5828 , \5829 , \5830 , \5831 , \5832 , \5833 , \5834 ,
         \5835 , \5836 , \5837 , \5838 , \5839 , \5840 , \5841 , \5842 , \5843 , \5844 ,
         \5845 , \5846 , \5847 , \5848 , \5849 , \5850 , \5851 , \5852 , \5853 , \5854 ,
         \5855 , \5856 , \5857 , \5858 , \5859 , \5860 , \5861 , \5862 , \5863 , \5864 ,
         \5865 , \5866 , \5867 , \5868 , \5869 , \5870 , \5871 , \5872 , \5873 , \5874 ,
         \5875 , \5876 , \5877 , \5878 , \5879 , \5880 , \5881 , \5882 , \5883 , \5884 ,
         \5885 , \5886 , \5887 , \5888 , \5889 , \5890 , \5891 , \5892 , \5893 , \5894 ,
         \5895 , \5896 , \5897 , \5898 , \5899 , \5900 , \5901 , \5902 , \5903 , \5904 ,
         \5905 , \5906 , \5907 , \5908 , \5909 , \5910 , \5911 , \5912 , \5913 , \5914 ,
         \5915 , \5916 , \5917 , \5918 , \5919 , \5920 , \5921 , \5922 , \5923 , \5924 ,
         \5925 , \5926 , \5927 , \5928 , \5929 , \5930 , \5931 , \5932 , \5933 , \5934 ,
         \5935 , \5936 , \5937 , \5938 , \5939 , \5940 , \5941 , \5942 , \5943 , \5944 ,
         \5945 , \5946 , \5947 , \5948 , \5949 , \5950 , \5951 , \5952 , \5953 , \5954 ,
         \5955 , \5956 , \5957 , \5958 , \5959 , \5960 , \5961 , \5962 , \5963 , \5964 ,
         \5965 , \5966 , \5967 , \5968 , \5969 , \5970 , \5971 , \5972 , \5973 , \5974 ,
         \5975 , \5976 , \5977 , \5978 , \5979 , \5980 , \5981 , \5982 , \5983 , \5984 ,
         \5985 , \5986 , \5987 , \5988 , \5989 , \5990 , \5991 , \5992 , \5993 , \5994 ,
         \5995 , \5996 , \5997 , \5998 , \5999 , \6000 , \6001 , \6002 , \6003 , \6004 ,
         \6005 , \6006 , \6007 , \6008 , \6009 , \6010 , \6011 , \6012 , \6013 , \6014 ,
         \6015 , \6016 , \6017 , \6018 , \6019 , \6020 , \6021 , \6022 , \6023 , \6024 ,
         \6025 , \6026 , \6027 , \6028 , \6029 , \6030 , \6031 , \6032 , \6033 , \6034 ,
         \6035 , \6036 , \6037 , \6038 , \6039 , \6040 , \6041 , \6042 , \6043 , \6044 ,
         \6045 , \6046 , \6047 , \6048 , \6049 , \6050 , \6051 , \6052 , \6053 , \6054 ,
         \6055 , \6056 , \6057 , \6058 , \6059 , \6060 , \6061 , \6062 , \6063 , \6064 ,
         \6065 , \6066 , \6067 , \6068 , \6069 , \6070 , \6071 , \6072 , \6073 , \6074 ,
         \6075 , \6076 , \6077 , \6078 , \6079 , \6080 , \6081 , \6082 , \6083 , \6084 ,
         \6085 , \6086 , \6087 , \6088 , \6089 , \6090 , \6091 , \6092 , \6093 , \6094 ,
         \6095 , \6096 , \6097 , \6098 , \6099 , \6100 , \6101 , \6102 , \6103 , \6104 ,
         \6105 , \6106 , \6107 , \6108 , \6109 , \6110 , \6111 , \6112 , \6113 , \6114 ,
         \6115 , \6116 , \6117 , \6118 , \6119 , \6120 , \6121 , \6122 , \6123 , \6124 ,
         \6125 , \6126 , \6127 , \6128 , \6129 , \6130 , \6131 , \6132 , \6133 , \6134 ,
         \6135 , \6136 , \6137 , \6138 , \6139 , \6140 , \6141 , \6142 , \6143 , \6144 ,
         \6145 , \6146 , \6147 , \6148 , \6149 , \6150 , \6151 , \6152 , \6153 , \6154 ,
         \6155 , \6156 , \6157 , \6158 , \6159 , \6160 , \6161 , \6162 , \6163 , \6164 ,
         \6165 , \6166 , \6167 , \6168 , \6169 , \6170 , \6171 , \6172 , \6173 , \6174 ,
         \6175 , \6176 , \6177 , \6178 , \6179 , \6180 , \6181 , \6182 , \6183 , \6184 ,
         \6185 , \6186 , \6187 , \6188 , \6189 , \6190 , \6191 , \6192 , \6193 , \6194 ,
         \6195 , \6196 , \6197 , \6198 , \6199 , \6200 , \6201 , \6202 , \6203 , \6204 ,
         \6205 , \6206 , \6207 , \6208 , \6209 , \6210 , \6211 , \6212 , \6213 , \6214 ,
         \6215 , \6216 , \6217 , \6218 , \6219 , \6220 , \6221 , \6222 , \6223 , \6224 ,
         \6225 , \6226 , \6227 , \6228 , \6229 , \6230 , \6231 , \6232 , \6233 , \6234 ,
         \6235 , \6236 , \6237 , \6238 , \6239 , \6240 , \6241 , \6242 , \6243 , \6244 ,
         \6245 , \6246 , \6247 , \6248 , \6249 , \6250 , \6251 , \6252 , \6253 , \6254 ,
         \6255 , \6256 , \6257 , \6258 , \6259 , \6260 , \6261 , \6262 , \6263 , \6264 ,
         \6265 , \6266 , \6267 , \6268 , \6269 , \6270 , \6271 , \6272 , \6273 , \6274 ,
         \6275 , \6276 , \6277 , \6278 , \6279 , \6280 , \6281 , \6282 , \6283 , \6284 ,
         \6285 , \6286 , \6287 , \6288 , \6289 , \6290 , \6291 , \6292 , \6293 , \6294 ,
         \6295 , \6296 , \6297 , \6298 , \6299 , \6300 , \6301 , \6302 , \6303 , \6304 ,
         \6305 , \6306 , \6307 , \6308 , \6309 , \6310 , \6311 , \6312 , \6313 , \6314 ,
         \6315 , \6316 , \6317 , \6318 , \6319 , \6320 , \6321 , \6322 , \6323 , \6324 ,
         \6325 , \6326 , \6327 , \6328 , \6329 , \6330 , \6331 , \6332 , \6333 , \6334 ,
         \6335 , \6336 , \6337 , \6338 , \6339 , \6340 , \6341 , \6342 , \6343 , \6344 ,
         \6345 , \6346 , \6347 , \6348 , \6349 , \6350 , \6351 , \6352 , \6353 , \6354 ,
         \6355 , \6356 , \6357 , \6358 , \6359 , \6360 , \6361 , \6362 , \6363 , \6364 ,
         \6365 , \6366 , \6367 , \6368 , \6369 , \6370 , \6371 , \6372 , \6373 , \6374 ,
         \6375 , \6376 , \6377 , \6378 , \6379 , \6380 , \6381 , \6382 , \6383 , \6384 ,
         \6385 , \6386 , \6387 , \6388 , \6389 , \6390 , \6391 , \6392 , \6393 , \6394 ,
         \6395 , \6396 , \6397 , \6398 , \6399 , \6400 , \6401 , \6402 , \6403 , \6404 ,
         \6405 , \6406 , \6407 , \6408 , \6409 , \6410 , \6411 , \6412 , \6413 , \6414 ,
         \6415 , \6416 , \6417 , \6418 , \6419 , \6420 , \6421 , \6422 , \6423 , \6424 ,
         \6425 , \6426 , \6427 , \6428 , \6429 , \6430 , \6431 , \6432 , \6433 , \6434 ,
         \6435 , \6436 , \6437 , \6438 , \6439 , \6440 , \6441 , \6442 , \6443 , \6444 ,
         \6445 , \6446 , \6447 , \6448 , \6449 , \6450 , \6451 , \6452 , \6453 , \6454 ,
         \6455 , \6456 , \6457 , \6458 , \6459 , \6460 , \6461 , \6462 , \6463 , \6464 ,
         \6465 , \6466 , \6467 , \6468 , \6469 , \6470 , \6471 , \6472 , \6473 , \6474 ,
         \6475 , \6476 , \6477 , \6478 , \6479 , \6480 , \6481 , \6482 , \6483 , \6484 ,
         \6485 , \6486 , \6487 , \6488 , \6489 , \6490 , \6491 , \6492 , \6493 , \6494 ,
         \6495 , \6496 , \6497 , \6498 , \6499 , \6500 , \6501 , \6502 , \6503 , \6504 ,
         \6505 , \6506 , \6507 , \6508 , \6509 , \6510 , \6511 , \6512 , \6513 , \6514 ,
         \6515 , \6516 , \6517 , \6518 , \6519 , \6520 , \6521 , \6522 , \6523 , \6524 ,
         \6525 , \6526 , \6527 , \6528 , \6529 , \6530 , \6531 , \6532 , \6533 , \6534 ,
         \6535 , \6536 , \6537 , \6538 , \6539 , \6540 , \6541 , \6542 , \6543 , \6544 ,
         \6545 , \6546 , \6547 , \6548 , \6549 , \6550 , \6551 , \6552 , \6553 , \6554 ,
         \6555 , \6556 , \6557 , \6558 , \6559 , \6560 , \6561 , \6562 , \6563 , \6564 ,
         \6565 , \6566 , \6567 , \6568 , \6569 , \6570 , \6571 , \6572 , \6573 , \6574 ,
         \6575 , \6576 , \6577 , \6578 , \6579 , \6580 , \6581 , \6582 , \6583 , \6584 ,
         \6585 , \6586 , \6587 , \6588 , \6589 , \6590 , \6591 , \6592 , \6593 , \6594 ,
         \6595 , \6596 , \6597 , \6598 , \6599 , \6600 , \6601 , \6602 , \6603 , \6604 ,
         \6605 , \6606 , \6607 , \6608 , \6609 , \6610 , \6611 , \6612 , \6613 , \6614 ,
         \6615 , \6616 , \6617 , \6618 , \6619 , \6620 , \6621 , \6622 , \6623 , \6624 ,
         \6625 , \6626 , \6627 , \6628 , \6629 , \6630 , \6631 , \6632 , \6633 , \6634 ,
         \6635 , \6636 , \6637 , \6638 , \6639 , \6640 , \6641 , \6642 , \6643 , \6644 ,
         \6645 , \6646 , \6647 , \6648 , \6649 , \6650 , \6651 , \6652 , \6653 , \6654 ,
         \6655 , \6656 , \6657 , \6658 , \6659 , \6660 , \6661 , \6662 , \6663 , \6664 ,
         \6665 , \6666 , \6667 , \6668 , \6669 , \6670 , \6671 , \6672 , \6673 , \6674 ,
         \6675 , \6676 , \6677 , \6678 , \6679 , \6680 , \6681 , \6682 , \6683 , \6684 ,
         \6685 , \6686 , \6687 , \6688 , \6689 , \6690 , \6691 , \6692 , \6693 , \6694 ,
         \6695 , \6696 , \6697 , \6698 , \6699 , \6700 , \6701 , \6702 , \6703 , \6704 ,
         \6705 , \6706 , \6707 , \6708 , \6709 , \6710 , \6711 , \6712 , \6713 , \6714 ,
         \6715 , \6716 , \6717 , \6718 , \6719 , \6720 , \6721 , \6722 , \6723 , \6724 ,
         \6725 , \6726 , \6727 , \6728 , \6729 , \6730 , \6731 , \6732 , \6733 , \6734 ,
         \6735 , \6736 , \6737 , \6738 , \6739 , \6740 , \6741 , \6742 , \6743 , \6744 ,
         \6745 , \6746 , \6747 , \6748 , \6749 , \6750 , \6751 , \6752 , \6753 , \6754 ,
         \6755 , \6756 , \6757 , \6758 , \6759 , \6760 , \6761 , \6762 , \6763 , \6764 ,
         \6765 , \6766 , \6767 , \6768 , \6769 , \6770 , \6771 , \6772 , \6773 , \6774 ,
         \6775 , \6776 , \6777 , \6778 , \6779 , \6780 , \6781 , \6782 , \6783 , \6784 ,
         \6785 , \6786 , \6787 , \6788 , \6789 , \6790 , \6791 , \6792 , \6793 , \6794 ,
         \6795 , \6796 , \6797 , \6798 , \6799 , \6800 , \6801 , \6802 , \6803 , \6804 ,
         \6805 , \6806 , \6807 , \6808 , \6809 , \6810 , \6811 , \6812 , \6813 , \6814 ,
         \6815 , \6816 , \6817 , \6818 , \6819 , \6820 , \6821 , \6822 , \6823 , \6824 ,
         \6825 , \6826 , \6827 , \6828 , \6829 , \6830 , \6831 , \6832 , \6833 , \6834 ,
         \6835 , \6836 , \6837 , \6838 , \6839 , \6840 , \6841 , \6842 , \6843 , \6844 ,
         \6845 , \6846 , \6847 , \6848 , \6849 , \6850 , \6851 , \6852 , \6853 , \6854 ,
         \6855 , \6856 , \6857 , \6858 , \6859 , \6860 , \6861 , \6862 , \6863 , \6864 ,
         \6865 , \6866 , \6867 , \6868 , \6869 , \6870 , \6871 , \6872 , \6873 , \6874 ,
         \6875 , \6876 , \6877 , \6878 , \6879 , \6880 , \6881 , \6882 , \6883 , \6884 ,
         \6885 , \6886 , \6887 , \6888 , \6889 , \6890 , \6891 , \6892 , \6893 , \6894 ,
         \6895 , \6896 , \6897 , \6898 , \6899 , \6900 , \6901 , \6902 , \6903 , \6904 ,
         \6905 , \6906 , \6907 , \6908 , \6909 , \6910 , \6911 , \6912 , \6913 , \6914 ,
         \6915 , \6916 , \6917 , \6918 , \6919 , \6920 , \6921 , \6922 , \6923 , \6924 ,
         \6925 , \6926 , \6927 , \6928 , \6929 , \6930 , \6931 , \6932 , \6933 , \6934 ,
         \6935 , \6936 , \6937 , \6938 , \6939 , \6940 , \6941 , \6942 , \6943 , \6944 ,
         \6945 , \6946 , \6947 , \6948 , \6949 , \6950 , \6951 , \6952 , \6953 , \6954 ,
         \6955 , \6956 , \6957 , \6958 , \6959 , \6960 , \6961 , \6962 , \6963 , \6964 ,
         \6965 , \6966 , \6967 , \6968 , \6969 , \6970 , \6971 , \6972 , \6973 , \6974 ,
         \6975 , \6976 , \6977 , \6978 , \6979 , \6980 , \6981 , \6982 , \6983 , \6984 ,
         \6985 , \6986 , \6987 , \6988 , \6989 , \6990 , \6991 , \6992 , \6993 , \6994 ,
         \6995 , \6996 , \6997 , \6998 , \6999 , \7000 , \7001 , \7002 , \7003 , \7004 ,
         \7005 , \7006 , \7007 , \7008 , \7009 , \7010 , \7011 , \7012 , \7013 , \7014 ,
         \7015 , \7016 , \7017 , \7018 , \7019 , \7020 , \7021 , \7022 , \7023 , \7024 ,
         \7025 , \7026 , \7027 , \7028 , \7029 , \7030 , \7031 , \7032 , \7033 , \7034 ,
         \7035 , \7036 , \7037 , \7038 , \7039 , \7040 , \7041 , \7042 , \7043 , \7044 ,
         \7045 , \7046 , \7047 , \7048 , \7049 , \7050 , \7051 , \7052 , \7053 , \7054 ,
         \7055 , \7056 , \7057 , \7058 , \7059 , \7060 , \7061 , \7062 , \7063 , \7064 ,
         \7065 , \7066 , \7067 , \7068 , \7069 , \7070 , \7071 , \7072 , \7073 , \7074 ,
         \7075 , \7076 , \7077 , \7078 , \7079 , \7080 , \7081 , \7082 , \7083 , \7084 ,
         \7085 , \7086 , \7087 , \7088 , \7089 , \7090 , \7091 , \7092 , \7093 , \7094 ,
         \7095 , \7096 , \7097 , \7098 , \7099 , \7100 , \7101 , \7102 , \7103 , \7104 ,
         \7105 , \7106 , \7107 , \7108 , \7109 , \7110 , \7111 , \7112 , \7113 , \7114 ,
         \7115 , \7116 , \7117 , \7118 , \7119 , \7120 , \7121 , \7122 , \7123 , \7124 ,
         \7125 , \7126 , \7127 , \7128 , \7129 , \7130 , \7131 , \7132 , \7133 , \7134 ,
         \7135 , \7136 , \7137 , \7138 , \7139 , \7140 , \7141 , \7142 , \7143 , \7144 ,
         \7145 , \7146 , \7147 , \7148 , \7149 , \7150 , \7151 , \7152 , \7153 , \7154 ,
         \7155 , \7156 , \7157 , \7158 , \7159 , \7160 , \7161 , \7162 , \7163 , \7164 ,
         \7165 , \7166 , \7167 , \7168 , \7169 , \7170 , \7171 , \7172 , \7173 , \7174 ,
         \7175 , \7176 , \7177 , \7178 , \7179 , \7180 , \7181 , \7182 , \7183 , \7184 ,
         \7185 , \7186 , \7187 , \7188 , \7189 , \7190 , \7191 , \7192 , \7193 , \7194 ,
         \7195 , \7196 , \7197 , \7198 , \7199 , \7200 , \7201 , \7202 , \7203 , \7204 ,
         \7205 , \7206 , \7207 , \7208 , \7209 , \7210 , \7211 , \7212 , \7213 , \7214 ,
         \7215 , \7216 , \7217 , \7218 , \7219 , \7220 , \7221 , \7222 , \7223 , \7224 ,
         \7225 , \7226 , \7227 , \7228 , \7229 , \7230 , \7231 , \7232 , \7233 , \7234 ,
         \7235 , \7236 , \7237 , \7238 , \7239 , \7240 , \7241 , \7242 , \7243 , \7244 ,
         \7245 , \7246 , \7247 , \7248 , \7249 , \7250 , \7251 , \7252 , \7253 , \7254 ,
         \7255 , \7256 , \7257 , \7258 , \7259 , \7260 , \7261 , \7262 , \7263 , \7264 ,
         \7265 , \7266 , \7267 , \7268 , \7269 , \7270 , \7271 , \7272 , \7273 , \7274 ,
         \7275 , \7276 , \7277 , \7278 , \7279 , \7280 , \7281 , \7282 , \7283 , \7284 ,
         \7285 , \7286 , \7287 , \7288 , \7289 , \7290 , \7291 , \7292 , \7293 , \7294 ,
         \7295 , \7296 , \7297 , \7298 , \7299 , \7300 , \7301 , \7302 , \7303 , \7304 ,
         \7305 , \7306 , \7307 , \7308 , \7309 , \7310 , \7311 , \7312 , \7313 , \7314 ,
         \7315 , \7316 , \7317 , \7318 , \7319 , \7320 , \7321 , \7322 , \7323 , \7324 ,
         \7325 , \7326 , \7327 , \7328 , \7329 , \7330 , \7331 , \7332 , \7333 , \7334 ,
         \7335 , \7336 , \7337 , \7338 , \7339 , \7340 , \7341 , \7342 , \7343 , \7344 ,
         \7345 , \7346 , \7347 , \7348 , \7349 , \7350 , \7351 , \7352 , \7353 , \7354 ,
         \7355 , \7356 , \7357 , \7358 , \7359 , \7360 , \7361 , \7362 , \7363 , \7364 ,
         \7365 , \7366 , \7367 , \7368 , \7369 , \7370 , \7371 , \7372 , \7373 , \7374 ,
         \7375 , \7376 , \7377 , \7378 , \7379 , \7380 , \7381 , \7382 , \7383 , \7384 ,
         \7385 , \7386 , \7387 , \7388 , \7389 , \7390 , \7391 , \7392 , \7393 , \7394 ,
         \7395 , \7396 , \7397 , \7398 , \7399 , \7400 , \7401 , \7402 , \7403 , \7404 ,
         \7405 , \7406 , \7407 , \7408 , \7409 , \7410 , \7411 , \7412 , \7413 , \7414 ,
         \7415 , \7416 , \7417 , \7418 , \7419 , \7420 , \7421 , \7422 , \7423 , \7424 ,
         \7425 , \7426 , \7427 , \7428 , \7429 , \7430 , \7431 , \7432 , \7433 , \7434 ,
         \7435 , \7436 , \7437 , \7438 , \7439 , \7440 , \7441 , \7442 , \7443 , \7444 ,
         \7445 , \7446 , \7447 , \7448 , \7449 , \7450 , \7451 , \7452 , \7453 , \7454 ,
         \7455 , \7456 , \7457 , \7458 , \7459 , \7460 , \7461 , \7462 , \7463 , \7464 ,
         \7465 , \7466 , \7467 , \7468 , \7469 , \7470 , \7471 , \7472 , \7473 , \7474 ,
         \7475 , \7476 , \7477 , \7478 , \7479 , \7480 , \7481 , \7482 , \7483 , \7484 ,
         \7485 , \7486 , \7487 , \7488 , \7489 , \7490 , \7491 , \7492 , \7493 , \7494 ,
         \7495 , \7496 , \7497 , \7498 , \7499 , \7500 , \7501 , \7502 , \7503 , \7504 ,
         \7505 , \7506 , \7507 , \7508 , \7509 , \7510 , \7511 , \7512 , \7513 , \7514 ,
         \7515 , \7516 , \7517 , \7518 , \7519 , \7520 , \7521 , \7522 , \7523 , \7524 ,
         \7525 , \7526 , \7527 , \7528 , \7529 , \7530 , \7531 , \7532 , \7533 , \7534 ,
         \7535 , \7536 , \7537 , \7538 , \7539 , \7540 , \7541 , \7542 , \7543 , \7544 ,
         \7545 , \7546 , \7547 , \7548 , \7549 , \7550 , \7551 , \7552 , \7553 , \7554 ,
         \7555 , \7556 , \7557 , \7558 , \7559 , \7560 , \7561 , \7562 , \7563 , \7564 ,
         \7565 , \7566 , \7567 , \7568 , \7569 , \7570 , \7571 , \7572 , \7573 , \7574 ,
         \7575 , \7576 , \7577 , \7578 , \7579 , \7580 , \7581 , \7582 , \7583 , \7584 ,
         \7585 , \7586 , \7587 , \7588 , \7589 , \7590 , \7591 , \7592 , \7593 , \7594 ,
         \7595 , \7596 , \7597 , \7598 , \7599 , \7600 , \7601 , \7602 , \7603 , \7604 ,
         \7605 , \7606 , \7607 , \7608 , \7609 , \7610 , \7611 , \7612 , \7613 , \7614 ,
         \7615 , \7616 , \7617 , \7618 , \7619 , \7620 , \7621 , \7622 , \7623 , \7624 ,
         \7625 , \7626 , \7627 , \7628 , \7629 , \7630 , \7631 , \7632 , \7633 , \7634 ,
         \7635 , \7636 , \7637 , \7638 , \7639 , \7640 , \7641 , \7642 , \7643 , \7644 ,
         \7645 , \7646 , \7647 , \7648 , \7649 , \7650 , \7651 , \7652 , \7653 , \7654 ,
         \7655 , \7656 , \7657 , \7658 , \7659 , \7660 , \7661 , \7662 , \7663 , \7664 ,
         \7665 , \7666 , \7667 , \7668 , \7669 , \7670 , \7671 , \7672 , \7673 , \7674 ,
         \7675 , \7676 , \7677 , \7678 , \7679 , \7680 , \7681 , \7682 , \7683 , \7684 ,
         \7685 , \7686 , \7687 , \7688 , \7689 , \7690 , \7691 , \7692 , \7693 , \7694 ,
         \7695 , \7696 , \7697 , \7698 , \7699 , \7700 , \7701 , \7702 , \7703 , \7704 ,
         \7705 , \7706 , \7707 , \7708 , \7709 , \7710 , \7711 , \7712 , \7713 , \7714 ,
         \7715 , \7716 , \7717 , \7718 , \7719 , \7720 , \7721 , \7722 , \7723 , \7724 ,
         \7725 , \7726 , \7727 , \7728 , \7729 , \7730 , \7731 , \7732 , \7733 , \7734 ,
         \7735 , \7736 , \7737 , \7738 , \7739 , \7740 , \7741 , \7742 , \7743 , \7744 ,
         \7745 , \7746 , \7747 , \7748 , \7749 , \7750 , \7751 , \7752 , \7753 , \7754 ,
         \7755 , \7756 , \7757 , \7758 , \7759 , \7760 , \7761 , \7762 , \7763 , \7764 ,
         \7765 , \7766 , \7767 , \7768 , \7769 , \7770 , \7771 , \7772 , \7773 , \7774 ,
         \7775 , \7776 , \7777 , \7778 , \7779 , \7780 , \7781 , \7782 , \7783 , \7784 ,
         \7785 , \7786 , \7787 , \7788 , \7789 , \7790 , \7791 , \7792 , \7793 , \7794 ,
         \7795 , \7796 , \7797 , \7798 , \7799 , \7800 , \7801 , \7802 , \7803 , \7804 ,
         \7805 , \7806 , \7807 , \7808 , \7809 , \7810 , \7811 , \7812 , \7813 , \7814 ,
         \7815 , \7816 , \7817 , \7818 , \7819 , \7820 , \7821 , \7822 , \7823 , \7824 ,
         \7825 , \7826 , \7827 , \7828 , \7829 , \7830 , \7831 , \7832 , \7833 , \7834 ,
         \7835 , \7836 , \7837 , \7838 , \7839 , \7840 , \7841 , \7842 , \7843 , \7844 ,
         \7845 , \7846 , \7847 , \7848 , \7849 , \7850 , \7851 , \7852 , \7853 , \7854 ,
         \7855 , \7856 , \7857 , \7858 , \7859 , \7860 , \7861 , \7862 , \7863 , \7864 ,
         \7865 , \7866 , \7867 , \7868 , \7869 , \7870 , \7871 , \7872 , \7873 , \7874 ,
         \7875 , \7876 , \7877 , \7878 , \7879 , \7880 , \7881 , \7882 , \7883 , \7884 ,
         \7885 , \7886 , \7887 , \7888 , \7889 , \7890 , \7891 , \7892 , \7893 , \7894 ,
         \7895 , \7896 , \7897 , \7898 , \7899 , \7900 , \7901 , \7902 , \7903 , \7904 ,
         \7905 , \7906 , \7907 , \7908 , \7909 , \7910 , \7911 , \7912 , \7913 , \7914 ,
         \7915 , \7916 , \7917 , \7918 , \7919 , \7920 , \7921 , \7922 , \7923 , \7924 ,
         \7925 , \7926 , \7927 , \7928 , \7929 , \7930 , \7931 , \7932 , \7933 , \7934 ,
         \7935 , \7936 , \7937 , \7938 , \7939 , \7940 , \7941 , \7942 , \7943 , \7944 ,
         \7945 , \7946 , \7947 , \7948 , \7949 , \7950 , \7951 , \7952 , \7953 , \7954 ,
         \7955 , \7956 , \7957 , \7958 , \7959 , \7960 , \7961 , \7962 , \7963 , \7964 ,
         \7965 , \7966 , \7967 , \7968 , \7969 , \7970 , \7971 , \7972 , \7973 , \7974 ,
         \7975 , \7976 , \7977 , \7978 , \7979 , \7980 , \7981 , \7982 , \7983 , \7984 ,
         \7985 , \7986 , \7987 , \7988 , \7989 , \7990 , \7991 , \7992 , \7993 , \7994 ,
         \7995 , \7996 , \7997 , \7998 , \7999 , \8000 , \8001 , \8002 , \8003 , \8004 ,
         \8005 , \8006 , \8007 , \8008 , \8009 , \8010 , \8011 , \8012 , \8013 , \8014 ,
         \8015 , \8016 , \8017 , \8018 , \8019 , \8020 , \8021 , \8022 , \8023 , \8024 ,
         \8025 , \8026 , \8027 , \8028 , \8029 , \8030 , \8031 , \8032 , \8033 , \8034 ,
         \8035 , \8036 , \8037 , \8038 , \8039 , \8040 , \8041 , \8042 , \8043 , \8044 ,
         \8045 , \8046 , \8047 , \8048 , \8049 , \8050 , \8051 , \8052 , \8053 , \8054 ,
         \8055 , \8056 , \8057 , \8058 , \8059 , \8060 , \8061 , \8062 , \8063 , \8064 ,
         \8065 , \8066 , \8067 , \8068 , \8069 , \8070 , \8071 , \8072 , \8073 , \8074 ,
         \8075 , \8076 , \8077 , \8078 , \8079 , \8080 , \8081 , \8082 , \8083 , \8084 ,
         \8085 , \8086 , \8087 , \8088 , \8089 , \8090 , \8091 , \8092 , \8093 , \8094 ,
         \8095 , \8096 , \8097 , \8098 , \8099 , \8100 , \8101 , \8102 , \8103 , \8104 ,
         \8105 , \8106 , \8107 , \8108 , \8109 , \8110 , \8111 , \8112 , \8113 , \8114 ,
         \8115 , \8116 , \8117 , \8118 , \8119 , \8120 , \8121 , \8122 , \8123 , \8124 ,
         \8125 , \8126 , \8127 , \8128 , \8129 , \8130 , \8131 , \8132 , \8133 , \8134 ,
         \8135 , \8136 , \8137 , \8138 , \8139 , \8140 , \8141 , \8142 , \8143 , \8144 ,
         \8145 , \8146 , \8147 , \8148 , \8149 , \8150 , \8151 , \8152 , \8153 , \8154 ,
         \8155 , \8156 , \8157 , \8158 , \8159 , \8160 , \8161 , \8162 , \8163 , \8164 ,
         \8165 , \8166 , \8167 , \8168 , \8169 , \8170 , \8171 , \8172 , \8173 , \8174 ,
         \8175 , \8176 , \8177 , \8178 , \8179 , \8180 , \8181 , \8182 , \8183 , \8184 ,
         \8185 , \8186 , \8187 , \8188 , \8189 , \8190 , \8191 , \8192 , \8193 , \8194 ,
         \8195 , \8196 , \8197 , \8198 , \8199 , \8200 , \8201 , \8202 , \8203 , \8204 ,
         \8205 , \8206 , \8207 , \8208 , \8209 , \8210 , \8211 , \8212 , \8213 , \8214 ,
         \8215 , \8216 , \8217 , \8218 , \8219 , \8220 , \8221 , \8222 , \8223 , \8224 ,
         \8225 , \8226 , \8227 , \8228 , \8229 , \8230 , \8231 , \8232 , \8233 , \8234 ,
         \8235 , \8236 , \8237 , \8238 , \8239 , \8240 , \8241 , \8242 , \8243 , \8244 ,
         \8245 , \8246 , \8247 , \8248 , \8249 , \8250 , \8251 , \8252 , \8253 , \8254 ,
         \8255 , \8256 , \8257 , \8258 , \8259 , \8260 , \8261 , \8262 , \8263 , \8264 ,
         \8265 , \8266 , \8267 , \8268 , \8269 , \8270 , \8271 , \8272 , \8273 , \8274 ,
         \8275 , \8276 , \8277 , \8278 , \8279 , \8280 , \8281 , \8282 , \8283 , \8284 ,
         \8285 , \8286 , \8287 , \8288 , \8289 , \8290 , \8291 , \8292 , \8293 , \8294 ,
         \8295 , \8296 , \8297 , \8298 , \8299 , \8300 , \8301 , \8302 , \8303 , \8304 ,
         \8305 , \8306 , \8307 , \8308 , \8309 , \8310 , \8311 , \8312 , \8313 , \8314 ,
         \8315 , \8316 , \8317 , \8318 , \8319 , \8320 , \8321 , \8322 , \8323 , \8324 ,
         \8325 , \8326 , \8327 , \8328 , \8329 , \8330 , \8331 , \8332 , \8333 , \8334 ,
         \8335 , \8336 , \8337 , \8338 , \8339 , \8340 , \8341 , \8342 , \8343 , \8344 ,
         \8345 , \8346 , \8347 , \8348 , \8349 , \8350 , \8351 , \8352 , \8353 , \8354 ,
         \8355 , \8356 , \8357 , \8358 , \8359 , \8360 , \8361 , \8362 , \8363 , \8364 ,
         \8365 , \8366 , \8367 , \8368 , \8369 , \8370 , \8371 , \8372 , \8373 , \8374 ,
         \8375 , \8376 , \8377 , \8378 , \8379 , \8380 , \8381 , \8382 , \8383 , \8384 ,
         \8385 , \8386 , \8387 , \8388 , \8389 , \8390 , \8391 , \8392 , \8393 , \8394 ,
         \8395 , \8396 , \8397 , \8398 , \8399 , \8400 , \8401 , \8402 , \8403 , \8404 ,
         \8405 , \8406 , \8407 , \8408 , \8409 , \8410 , \8411 , \8412 , \8413 , \8414 ,
         \8415 , \8416 , \8417 , \8418 , \8419 , \8420 , \8421 , \8422 , \8423 , \8424 ,
         \8425 , \8426 , \8427 , \8428 , \8429 , \8430 , \8431 , \8432 , \8433 , \8434 ,
         \8435 , \8436 , \8437 , \8438 , \8439 , \8440 , \8441 , \8442 , \8443 , \8444 ,
         \8445 , \8446 , \8447 , \8448 , \8449 , \8450 , \8451 , \8452 , \8453 , \8454 ,
         \8455 , \8456 , \8457 , \8458 , \8459 , \8460 , \8461 , \8462 , \8463 , \8464 ,
         \8465 , \8466 , \8467 , \8468 , \8469 , \8470 , \8471 , \8472 , \8473 , \8474 ,
         \8475 , \8476 , \8477 , \8478 , \8479 , \8480 , \8481 , \8482 , \8483 , \8484 ,
         \8485 , \8486 , \8487 , \8488 , \8489 , \8490 , \8491 , \8492 , \8493 , \8494 ,
         \8495 , \8496 , \8497 , \8498 , \8499 , \8500 , \8501 , \8502 , \8503 , \8504 ,
         \8505 , \8506 , \8507 , \8508 , \8509 , \8510 , \8511 , \8512 , \8513 , \8514 ,
         \8515 , \8516 , \8517 , \8518 , \8519 , \8520 , \8521 , \8522 , \8523 , \8524 ,
         \8525 , \8526 , \8527 , \8528 , \8529 , \8530 , \8531 , \8532 , \8533 , \8534 ,
         \8535 , \8536 , \8537 , \8538 , \8539 , \8540 , \8541 , \8542 , \8543 , \8544 ,
         \8545 , \8546 , \8547 , \8548 , \8549 , \8550 , \8551 , \8552 , \8553 , \8554 ,
         \8555 , \8556 , \8557 , \8558 , \8559 , \8560 , \8561 , \8562 , \8563 , \8564 ,
         \8565 , \8566 , \8567 , \8568 , \8569 , \8570 , \8571 , \8572 , \8573 , \8574 ,
         \8575 , \8576 , \8577 , \8578 , \8579 , \8580 , \8581 , \8582 , \8583 , \8584 ,
         \8585 , \8586 , \8587 , \8588 , \8589 , \8590 , \8591 , \8592 , \8593 , \8594 ,
         \8595 , \8596 , \8597 , \8598 , \8599 , \8600 , \8601 , \8602 , \8603 , \8604 ,
         \8605 , \8606 , \8607 , \8608 , \8609 , \8610 , \8611 , \8612 , \8613 , \8614 ,
         \8615 , \8616 , \8617 , \8618 , \8619 , \8620 , \8621 , \8622 , \8623 , \8624 ,
         \8625 , \8626 , \8627 , \8628 , \8629 , \8630 , \8631 , \8632 , \8633 , \8634 ,
         \8635 , \8636 , \8637 , \8638 , \8639 , \8640 , \8641 , \8642 , \8643 , \8644 ,
         \8645 , \8646 , \8647 , \8648 , \8649 , \8650 , \8651 , \8652 , \8653 , \8654 ,
         \8655 , \8656 , \8657 , \8658 , \8659 , \8660 , \8661 , \8662 , \8663 , \8664 ,
         \8665 , \8666 , \8667 , \8668 , \8669 , \8670 , \8671 , \8672 , \8673 , \8674 ,
         \8675 , \8676 , \8677 , \8678 , \8679 , \8680 , \8681 , \8682 , \8683 , \8684 ,
         \8685 , \8686 , \8687 , \8688 , \8689 , \8690 , \8691 , \8692 , \8693 , \8694 ,
         \8695 , \8696 , \8697 , \8698 , \8699 , \8700 , \8701 , \8702 , \8703 , \8704 ,
         \8705 , \8706 , \8707 , \8708 , \8709 , \8710 , \8711 , \8712 , \8713 , \8714 ,
         \8715 , \8716 , \8717 , \8718 , \8719 , \8720 , \8721 , \8722 , \8723 , \8724 ,
         \8725 , \8726 , \8727 , \8728 , \8729 , \8730 , \8731 , \8732 , \8733 , \8734 ,
         \8735 , \8736 , \8737 , \8738 , \8739 , \8740 , \8741 , \8742 , \8743 , \8744 ,
         \8745 , \8746 , \8747 , \8748 , \8749 , \8750 , \8751 , \8752 , \8753 , \8754 ,
         \8755 , \8756 , \8757 , \8758 , \8759 , \8760 , \8761 , \8762 , \8763 , \8764 ,
         \8765 , \8766 , \8767 , \8768 , \8769 , \8770 , \8771 , \8772 , \8773 , \8774 ,
         \8775 , \8776 , \8777 , \8778 , \8779 , \8780 , \8781 , \8782 , \8783 , \8784 ,
         \8785 , \8786 , \8787 , \8788 , \8789 , \8790 , \8791 , \8792 , \8793 , \8794 ,
         \8795 , \8796 , \8797 , \8798 , \8799 , \8800 , \8801 , \8802 , \8803 , \8804 ,
         \8805 , \8806 , \8807 , \8808 , \8809 , \8810 , \8811 , \8812 , \8813 , \8814 ,
         \8815 , \8816 , \8817 , \8818 , \8819 , \8820 , \8821 , \8822 , \8823 , \8824 ,
         \8825 , \8826 , \8827 , \8828 , \8829 , \8830 , \8831 , \8832 , \8833 , \8834 ,
         \8835 , \8836 , \8837 , \8838 , \8839 , \8840 , \8841 , \8842 , \8843 , \8844 ,
         \8845 , \8846 , \8847 , \8848 , \8849 , \8850 , \8851 , \8852 , \8853 , \8854 ,
         \8855 , \8856 , \8857 , \8858 , \8859 , \8860 , \8861 , \8862 , \8863 , \8864 ,
         \8865 , \8866 , \8867 , \8868 , \8869 , \8870 , \8871 , \8872 , \8873 , \8874 ,
         \8875 , \8876 , \8877 , \8878 , \8879 , \8880 , \8881 , \8882 , \8883 , \8884 ,
         \8885 , \8886 , \8887 , \8888 , \8889 , \8890 , \8891 , \8892 , \8893 , \8894 ,
         \8895 , \8896 , \8897 , \8898 , \8899 , \8900 , \8901 , \8902 , \8903 , \8904 ,
         \8905 , \8906 , \8907 , \8908 , \8909 , \8910 , \8911 , \8912 , \8913 , \8914 ,
         \8915 , \8916 , \8917 , \8918 , \8919 , \8920 , \8921 , \8922 , \8923 , \8924 ,
         \8925 , \8926 , \8927 , \8928 , \8929 , \8930 , \8931 , \8932 , \8933 , \8934 ,
         \8935 , \8936 , \8937 , \8938 , \8939 , \8940 , \8941 , \8942 , \8943 , \8944 ,
         \8945 , \8946 , \8947 , \8948 , \8949 , \8950 , \8951 , \8952 , \8953 , \8954 ,
         \8955 , \8956 , \8957 , \8958 , \8959 , \8960 , \8961 , \8962 , \8963 , \8964 ,
         \8965 , \8966 , \8967 , \8968 , \8969 , \8970 , \8971 , \8972 , \8973 , \8974 ,
         \8975 , \8976 , \8977 , \8978 , \8979 , \8980 , \8981 , \8982 , \8983 , \8984 ,
         \8985 , \8986 , \8987 , \8988 , \8989 , \8990 , \8991 , \8992 , \8993 , \8994 ,
         \8995 , \8996 , \8997 , \8998 , \8999 , \9000 , \9001 , \9002 , \9003 , \9004 ,
         \9005 , \9006 , \9007 , \9008 , \9009 , \9010 , \9011 , \9012 , \9013 , \9014 ,
         \9015 , \9016 , \9017 , \9018 , \9019 , \9020 , \9021 , \9022 , \9023 , \9024 ,
         \9025 , \9026 , \9027 , \9028 , \9029 , \9030 , \9031 , \9032 , \9033 , \9034 ,
         \9035 , \9036 , \9037 , \9038 , \9039 , \9040 , \9041 , \9042 , \9043 , \9044 ,
         \9045 , \9046 , \9047 , \9048 , \9049 , \9050 , \9051 , \9052 , \9053 , \9054 ,
         \9055 , \9056 , \9057 , \9058 , \9059 , \9060 , \9061 , \9062 , \9063 , \9064 ,
         \9065 , \9066 , \9067 , \9068 , \9069 , \9070 , \9071 , \9072 , \9073 , \9074 ,
         \9075 , \9076 , \9077 , \9078 , \9079 , \9080 , \9081 , \9082 , \9083 , \9084 ,
         \9085 , \9086 , \9087 , \9088 , \9089 , \9090 , \9091 , \9092 , \9093 , \9094 ,
         \9095 , \9096 , \9097 , \9098 , \9099 , \9100 , \9101 , \9102 , \9103 , \9104 ,
         \9105 , \9106 , \9107 , \9108 , \9109 , \9110 , \9111 , \9112 , \9113 , \9114 ,
         \9115 , \9116 , \9117 , \9118 , \9119 , \9120 , \9121 , \9122 , \9123 , \9124 ,
         \9125 , \9126 , \9127 , \9128 , \9129 , \9130 , \9131 , \9132 , \9133 , \9134 ,
         \9135 , \9136 , \9137 , \9138 , \9139 , \9140 , \9141 , \9142 , \9143 , \9144 ,
         \9145 , \9146 , \9147 , \9148 , \9149 , \9150 , \9151 , \9152 , \9153 , \9154 ,
         \9155 , \9156 , \9157 , \9158 , \9159 , \9160 , \9161 , \9162 , \9163 , \9164 ,
         \9165 , \9166 , \9167 , \9168 , \9169 , \9170 , \9171 , \9172 , \9173 , \9174 ,
         \9175 , \9176 , \9177 , \9178 , \9179 , \9180 , \9181 , \9182 , \9183 , \9184 ,
         \9185 , \9186 , \9187 , \9188 , \9189 , \9190 , \9191 , \9192 , \9193 , \9194 ,
         \9195 , \9196 , \9197 , \9198 , \9199 , \9200 , \9201 , \9202 , \9203 , \9204 ,
         \9205 , \9206 , \9207 , \9208 , \9209 , \9210 , \9211 , \9212 , \9213 , \9214 ,
         \9215 , \9216 , \9217 , \9218 , \9219 , \9220 , \9221 , \9222 , \9223 , \9224 ,
         \9225 , \9226 , \9227 , \9228 , \9229 , \9230 , \9231 , \9232 , \9233 , \9234 ,
         \9235 , \9236 , \9237 , \9238 , \9239 , \9240 , \9241 , \9242 , \9243 , \9244 ,
         \9245 , \9246 , \9247 , \9248 , \9249 , \9250 , \9251 , \9252 , \9253 , \9254 ,
         \9255 , \9256 , \9257 , \9258 , \9259 , \9260 , \9261 , \9262 , \9263 , \9264 ,
         \9265 , \9266 , \9267 , \9268 , \9269 , \9270 , \9271 , \9272 , \9273 , \9274 ,
         \9275 , \9276 , \9277 , \9278 , \9279 , \9280 , \9281 , \9282 , \9283 , \9284 ,
         \9285 , \9286 , \9287 , \9288 , \9289 , \9290 , \9291 , \9292 , \9293 , \9294 ,
         \9295 , \9296 , \9297 , \9298 , \9299 , \9300 , \9301 , \9302 , \9303 , \9304 ,
         \9305 , \9306 , \9307 , \9308 , \9309 , \9310 , \9311 , \9312 , \9313 , \9314 ,
         \9315 , \9316 , \9317 , \9318 , \9319 , \9320 , \9321 , \9322 , \9323 , \9324 ,
         \9325 , \9326 , \9327 , \9328 , \9329 , \9330 , \9331 , \9332 , \9333 , \9334 ,
         \9335 , \9336 , \9337 , \9338 , \9339 , \9340 , \9341 , \9342 , \9343 , \9344 ,
         \9345 , \9346 , \9347 , \9348 , \9349 , \9350 , \9351 , \9352 , \9353 , \9354 ,
         \9355 , \9356 , \9357 , \9358 , \9359 , \9360 , \9361 , \9362 , \9363 , \9364 ,
         \9365 , \9366 , \9367 , \9368 , \9369 , \9370 , \9371 , \9372 , \9373 , \9374 ,
         \9375 , \9376 , \9377 , \9378 , \9379 , \9380 , \9381 , \9382 , \9383 , \9384 ,
         \9385 , \9386 , \9387 , \9388 , \9389 , \9390 , \9391 , \9392 , \9393 , \9394 ,
         \9395 , \9396 , \9397 , \9398 , \9399 , \9400 , \9401 , \9402 , \9403 , \9404 ,
         \9405 , \9406 , \9407 , \9408 , \9409 , \9410 , \9411 , \9412 , \9413 , \9414 ,
         \9415 , \9416 , \9417 , \9418 , \9419 , \9420 , \9421 , \9422 , \9423 , \9424 ,
         \9425 , \9426 , \9427 , \9428 , \9429 , \9430 , \9431 , \9432 , \9433 , \9434 ,
         \9435 , \9436 , \9437 , \9438 , \9439 , \9440 , \9441 , \9442 , \9443 , \9444 ,
         \9445 , \9446 , \9447 , \9448 , \9449 , \9450 , \9451 , \9452 , \9453 , \9454 ,
         \9455 , \9456 , \9457 , \9458 , \9459 , \9460 , \9461 , \9462 , \9463 , \9464 ,
         \9465 , \9466 , \9467 , \9468 , \9469 , \9470 , \9471 , \9472 , \9473 , \9474 ,
         \9475 , \9476 , \9477 , \9478 , \9479 , \9480 , \9481 , \9482 , \9483 , \9484 ,
         \9485 , \9486 , \9487 , \9488 , \9489 , \9490 , \9491 , \9492 , \9493 , \9494 ,
         \9495 , \9496 , \9497 , \9498 , \9499 , \9500 , \9501 , \9502 , \9503 , \9504 ,
         \9505 , \9506 , \9507 , \9508 , \9509 , \9510 , \9511 , \9512 , \9513 , \9514 ,
         \9515 , \9516 , \9517 , \9518 , \9519 , \9520 , \9521 , \9522 , \9523 , \9524 ,
         \9525 , \9526 , \9527 , \9528 , \9529 , \9530 , \9531 , \9532 , \9533 , \9534 ,
         \9535 , \9536 , \9537 , \9538 , \9539 , \9540 , \9541 , \9542 , \9543 , \9544 ,
         \9545 , \9546 , \9547 , \9548 , \9549 , \9550 , \9551 , \9552 , \9553 , \9554 ,
         \9555 , \9556 , \9557 , \9558 , \9559 , \9560 , \9561 , \9562 , \9563 , \9564 ,
         \9565 , \9566 , \9567 , \9568 , \9569 , \9570 , \9571 , \9572 , \9573 , \9574 ,
         \9575 , \9576 , \9577 , \9578 , \9579 , \9580 , \9581 , \9582 , \9583 , \9584 ,
         \9585 , \9586 , \9587 , \9588 , \9589 , \9590 , \9591 , \9592 , \9593 , \9594 ,
         \9595 , \9596 , \9597 , \9598 , \9599 , \9600 , \9601 , \9602 , \9603 , \9604 ,
         \9605 , \9606 , \9607 , \9608 , \9609 , \9610 , \9611 , \9612 , \9613 , \9614 ,
         \9615 , \9616 , \9617 , \9618 , \9619 , \9620 , \9621 , \9622 , \9623 , \9624 ,
         \9625 , \9626 , \9627 , \9628 , \9629 , \9630 , \9631 , \9632 , \9633 , \9634 ,
         \9635 , \9636 , \9637 , \9638 , \9639 , \9640 , \9641 , \9642 , \9643 , \9644 ,
         \9645 , \9646 , \9647 , \9648 , \9649 , \9650 , \9651 , \9652 , \9653 , \9654 ,
         \9655 , \9656 , \9657 , \9658 , \9659 , \9660 , \9661 , \9662 , \9663 , \9664 ,
         \9665 , \9666 , \9667 , \9668 , \9669 , \9670 , \9671 , \9672 , \9673 , \9674 ,
         \9675 , \9676 , \9677 , \9678 , \9679 , \9680 , \9681 , \9682 , \9683 , \9684 ,
         \9685 , \9686 , \9687 , \9688 , \9689 , \9690 , \9691 , \9692 , \9693 , \9694 ,
         \9695 , \9696 , \9697 , \9698 , \9699 , \9700 , \9701 , \9702 , \9703 , \9704 ,
         \9705 , \9706 , \9707 , \9708 , \9709 , \9710 , \9711 , \9712 , \9713 , \9714 ,
         \9715 , \9716 , \9717 , \9718 , \9719 , \9720 , \9721 , \9722 , \9723 , \9724 ,
         \9725 , \9726 , \9727 , \9728 , \9729 , \9730 , \9731 , \9732 , \9733 , \9734 ,
         \9735 , \9736 , \9737 , \9738 , \9739 , \9740 , \9741 , \9742 , \9743 , \9744 ,
         \9745 , \9746 , \9747 , \9748 , \9749 , \9750 , \9751 , \9752 , \9753 , \9754 ,
         \9755 , \9756 , \9757 , \9758 , \9759 , \9760 , \9761 , \9762 , \9763 , \9764 ,
         \9765 , \9766 , \9767 , \9768 , \9769 , \9770 , \9771 , \9772 , \9773 , \9774 ,
         \9775 , \9776 , \9777 , \9778 , \9779 , \9780 , \9781 , \9782 , \9783 , \9784 ,
         \9785 , \9786 , \9787 , \9788 , \9789 , \9790 , \9791 , \9792 , \9793 , \9794 ,
         \9795 , \9796 , \9797 , \9798 , \9799 , \9800 , \9801 , \9802 , \9803 , \9804 ,
         \9805 , \9806 , \9807 , \9808 , \9809 , \9810 , \9811 , \9812 , \9813 , \9814 ,
         \9815 , \9816 , \9817 , \9818 , \9819 , \9820 , \9821 , \9822 , \9823 , \9824 ,
         \9825 , \9826 , \9827 , \9828 , \9829 , \9830 , \9831 , \9832 , \9833 , \9834 ,
         \9835 , \9836 , \9837 , \9838 , \9839 , \9840 , \9841 , \9842 , \9843 , \9844 ,
         \9845 , \9846 , \9847 , \9848 , \9849 , \9850 , \9851 , \9852 , \9853 , \9854 ,
         \9855 , \9856 , \9857 , \9858 , \9859 , \9860 , \9861 , \9862 , \9863 , \9864 ,
         \9865 , \9866 , \9867 , \9868 , \9869 , \9870 , \9871 , \9872 , \9873 , \9874 ,
         \9875 , \9876 , \9877 , \9878 , \9879 , \9880 , \9881 , \9882 , \9883 , \9884 ,
         \9885 , \9886 , \9887 , \9888 , \9889 , \9890 , \9891 , \9892 , \9893 , \9894 ,
         \9895 , \9896 , \9897 , \9898 , \9899 , \9900 , \9901 , \9902 , \9903 , \9904 ,
         \9905 , \9906 , \9907 , \9908 , \9909 , \9910 , \9911 , \9912 , \9913 , \9914 ,
         \9915 , \9916 , \9917 , \9918 , \9919 , \9920 , \9921 , \9922 , \9923 , \9924 ,
         \9925 , \9926 , \9927 , \9928 , \9929 , \9930 , \9931 , \9932 , \9933 , \9934 ,
         \9935 , \9936 , \9937 , \9938 , \9939 , \9940 , \9941 , \9942 , \9943 , \9944 ,
         \9945 , \9946 , \9947 , \9948 , \9949 , \9950 , \9951 , \9952 , \9953 , \9954 ,
         \9955 , \9956 , \9957 , \9958 , \9959 , \9960 , \9961 , \9962 , \9963 , \9964 ,
         \9965 , \9966 , \9967 , \9968 , \9969 , \9970 , \9971 , \9972 , \9973 , \9974 ,
         \9975 , \9976 , \9977 , \9978 , \9979 , \9980 , \9981 , \9982 , \9983 , \9984 ,
         \9985 , \9986 , \9987 , \9988 , \9989 , \9990 , \9991 , \9992 , \9993 , \9994 ,
         \9995 , \9996 , \9997 , \9998 , \9999 , \10000 , \10001 , \10002 , \10003 , \10004 ,
         \10005 , \10006 , \10007 , \10008 , \10009 , \10010 , \10011 , \10012 , \10013 , \10014 ,
         \10015 , \10016 , \10017 , \10018 , \10019 , \10020 , \10021 , \10022 , \10023 , \10024 ,
         \10025 , \10026 , \10027 , \10028 , \10029 , \10030 , \10031 , \10032 , \10033 , \10034 ,
         \10035 , \10036 , \10037 , \10038 , \10039 , \10040 , \10041 , \10042 , \10043 , \10044 ,
         \10045 , \10046 , \10047 , \10048 , \10049 , \10050 , \10051 , \10052 , \10053 , \10054 ,
         \10055 , \10056 , \10057 , \10058 , \10059 , \10060 , \10061 , \10062 , \10063 , \10064 ,
         \10065 , \10066 , \10067 , \10068 , \10069 , \10070 , \10071 , \10072 , \10073 , \10074 ,
         \10075 , \10076 , \10077 , \10078 , \10079 , \10080 , \10081 , \10082 , \10083 , \10084 ,
         \10085 , \10086 , \10087 , \10088 , \10089 , \10090 , \10091 , \10092 , \10093 , \10094 ,
         \10095 , \10096 , \10097 , \10098 , \10099 , \10100 , \10101 , \10102 , \10103 , \10104 ,
         \10105 , \10106 , \10107 , \10108 , \10109 , \10110 , \10111 , \10112 , \10113 , \10114 ,
         \10115 , \10116 , \10117 , \10118 , \10119 , \10120 , \10121 , \10122 , \10123 , \10124 ,
         \10125 , \10126 , \10127 , \10128 , \10129 , \10130 , \10131 , \10132 , \10133 , \10134 ,
         \10135 , \10136 , \10137 , \10138 , \10139 , \10140 , \10141 , \10142 , \10143 , \10144 ,
         \10145 , \10146 , \10147 , \10148 , \10149 , \10150 , \10151 , \10152 , \10153 , \10154 ,
         \10155 , \10156 , \10157 , \10158 , \10159 , \10160 , \10161 , \10162 , \10163 , \10164 ,
         \10165 , \10166 , \10167 , \10168 , \10169 , \10170 , \10171 , \10172 , \10173 , \10174 ,
         \10175 , \10176 , \10177 , \10178 , \10179 , \10180 , \10181 , \10182 , \10183 , \10184 ,
         \10185 , \10186 , \10187 , \10188 , \10189 , \10190 , \10191 , \10192 , \10193 , \10194 ,
         \10195 , \10196 , \10197 , \10198 , \10199 , \10200 , \10201 , \10202 , \10203 , \10204 ,
         \10205 , \10206 , \10207 , \10208 , \10209 , \10210 , \10211 , \10212 , \10213 , \10214 ,
         \10215 , \10216 , \10217 , \10218 , \10219 , \10220 , \10221 , \10222 , \10223 , \10224 ,
         \10225 , \10226 , \10227 , \10228 , \10229 , \10230 , \10231 , \10232 , \10233 , \10234 ,
         \10235 , \10236 , \10237 , \10238 , \10239 , \10240 , \10241 , \10242 , \10243 , \10244 ,
         \10245 , \10246 , \10247 , \10248 , \10249 , \10250 , \10251 , \10252 , \10253 , \10254 ,
         \10255 , \10256 , \10257 , \10258 , \10259 , \10260 , \10261 , \10262 , \10263 , \10264 ,
         \10265 , \10266 , \10267 , \10268 , \10269 , \10270 , \10271 , \10272 , \10273 , \10274 ,
         \10275 , \10276 , \10277 , \10278 , \10279 , \10280 , \10281 , \10282 , \10283 , \10284 ,
         \10285 , \10286 , \10287 , \10288 , \10289 , \10290 , \10291 , \10292 , \10293 , \10294 ,
         \10295 , \10296 , \10297 , \10298 , \10299 , \10300 , \10301 , \10302 , \10303 , \10304 ,
         \10305 , \10306 , \10307 , \10308 , \10309 , \10310 , \10311 , \10312 , \10313 , \10314 ,
         \10315 , \10316 , \10317 , \10318 , \10319 , \10320 , \10321 , \10322 , \10323 , \10324 ,
         \10325 , \10326 , \10327 , \10328 , \10329 , \10330 , \10331 , \10332 , \10333 , \10334 ,
         \10335 , \10336 , \10337 , \10338 , \10339 , \10340 , \10341 , \10342 , \10343 , \10344 ,
         \10345 , \10346 , \10347 , \10348 , \10349 , \10350 , \10351 , \10352 , \10353 , \10354 ,
         \10355 , \10356 , \10357 , \10358 , \10359 , \10360 , \10361 , \10362 , \10363 , \10364 ,
         \10365 , \10366 , \10367 , \10368 , \10369 , \10370 , \10371 , \10372 , \10373 , \10374 ,
         \10375 , \10376 , \10377 , \10378 , \10379 , \10380 , \10381 , \10382 , \10383 , \10384 ,
         \10385 , \10386 , \10387 , \10388 , \10389 , \10390 , \10391 , \10392 , \10393 , \10394 ,
         \10395 , \10396 , \10397 , \10398 , \10399 , \10400 , \10401 , \10402 , \10403 , \10404 ,
         \10405 , \10406 , \10407 , \10408 , \10409 , \10410 , \10411 , \10412 , \10413 , \10414 ,
         \10415 , \10416 , \10417 , \10418 , \10419 , \10420 , \10421 , \10422 , \10423 , \10424 ,
         \10425 , \10426 , \10427 , \10428 , \10429 , \10430 , \10431 , \10432 , \10433 , \10434 ,
         \10435 , \10436 , \10437 , \10438 , \10439 , \10440 , \10441 , \10442 , \10443 , \10444 ,
         \10445 , \10446 , \10447 , \10448 , \10449 , \10450 , \10451 , \10452 , \10453 , \10454 ,
         \10455 , \10456 , \10457 , \10458 , \10459 , \10460 , \10461 , \10462 , \10463 , \10464 ,
         \10465 , \10466 , \10467 , \10468 , \10469 , \10470 , \10471 , \10472 , \10473 , \10474 ,
         \10475 , \10476 , \10477 , \10478 , \10479 , \10480 , \10481 , \10482 , \10483 , \10484 ,
         \10485 , \10486 , \10487 , \10488 , \10489 , \10490 , \10491 , \10492 , \10493 , \10494 ,
         \10495 , \10496 , \10497 , \10498 , \10499 , \10500 , \10501 , \10502 , \10503 , \10504 ,
         \10505 , \10506 , \10507 , \10508 , \10509 , \10510 , \10511 , \10512 , \10513 , \10514 ,
         \10515 , \10516 , \10517 , \10518 , \10519 , \10520 , \10521 , \10522 , \10523 , \10524 ,
         \10525 , \10526 , \10527 , \10528 , \10529 , \10530 , \10531 , \10532 , \10533 , \10534 ,
         \10535 , \10536 , \10537 , \10538 , \10539 , \10540 , \10541 , \10542 , \10543 , \10544 ,
         \10545 , \10546 , \10547 , \10548 , \10549 , \10550 , \10551 , \10552 , \10553 , \10554 ,
         \10555 , \10556 , \10557 , \10558 , \10559 , \10560 , \10561 , \10562 , \10563 , \10564 ,
         \10565 , \10566 , \10567 , \10568 , \10569 , \10570 , \10571 , \10572 , \10573 , \10574 ,
         \10575 , \10576 , \10577 , \10578 , \10579 , \10580 , \10581 , \10582 , \10583 , \10584 ,
         \10585 , \10586 , \10587 , \10588 , \10589 , \10590 , \10591 , \10592 , \10593 , \10594 ,
         \10595 , \10596 , \10597 , \10598 , \10599 , \10600 , \10601 , \10602 , \10603 , \10604 ,
         \10605 , \10606 , \10607 , \10608 , \10609 , \10610 , \10611 , \10612 , \10613 , \10614 ,
         \10615 , \10616 , \10617 , \10618 , \10619 , \10620 , \10621 , \10622 , \10623 , \10624 ,
         \10625 , \10626 , \10627 , \10628 , \10629 , \10630 , \10631 , \10632 , \10633 , \10634 ,
         \10635 , \10636 , \10637 , \10638 , \10639 , \10640 , \10641 , \10642 , \10643 , \10644 ,
         \10645 , \10646 , \10647 , \10648 , \10649 , \10650 , \10651 , \10652 , \10653 , \10654 ,
         \10655 , \10656 , \10657 , \10658 , \10659 , \10660 , \10661 , \10662 , \10663 , \10664 ,
         \10665 , \10666 , \10667 , \10668 , \10669 , \10670 , \10671 , \10672 , \10673 , \10674 ,
         \10675 , \10676 , \10677 , \10678 , \10679 , \10680 , \10681 , \10682 , \10683 , \10684 ,
         \10685 , \10686 , \10687 , \10688 , \10689 , \10690 , \10691 , \10692 , \10693 , \10694 ,
         \10695 , \10696 , \10697 , \10698 , \10699 , \10700 , \10701 , \10702 , \10703 , \10704 ,
         \10705 , \10706 , \10707 , \10708 , \10709 , \10710 , \10711 , \10712 , \10713 , \10714 ,
         \10715 , \10716 , \10717 , \10718 , \10719 , \10720 , \10721 , \10722 , \10723 , \10724 ,
         \10725 , \10726 , \10727 , \10728 , \10729 , \10730 , \10731 , \10732 , \10733 , \10734 ,
         \10735 , \10736 , \10737 , \10738 , \10739 , \10740 , \10741 , \10742 , \10743 , \10744 ,
         \10745 , \10746 , \10747 , \10748 , \10749 , \10750 , \10751 , \10752 , \10753 , \10754 ,
         \10755 , \10756 , \10757 , \10758 , \10759 , \10760 , \10761 , \10762 , \10763 , \10764 ,
         \10765 , \10766 , \10767 , \10768 , \10769 , \10770 , \10771 , \10772 , \10773 , \10774 ,
         \10775 , \10776 , \10777 , \10778 , \10779 , \10780 , \10781 , \10782 , \10783 , \10784 ,
         \10785 , \10786 , \10787 , \10788 , \10789 , \10790 , \10791 , \10792 , \10793 , \10794 ,
         \10795 , \10796 , \10797 , \10798 , \10799 , \10800 , \10801 , \10802 , \10803 , \10804 ,
         \10805 , \10806 , \10807 , \10808 , \10809 , \10810 , \10811 , \10812 , \10813 , \10814 ,
         \10815 , \10816 , \10817 , \10818 , \10819 , \10820 , \10821 , \10822 , \10823 , \10824 ,
         \10825 , \10826 , \10827 , \10828 , \10829 , \10830 , \10831 , \10832 , \10833 , \10834 ,
         \10835 , \10836 , \10837 , \10838 , \10839 , \10840 , \10841 , \10842 , \10843 , \10844 ,
         \10845 , \10846 , \10847 , \10848 , \10849 , \10850 , \10851 , \10852 , \10853 , \10854 ,
         \10855 , \10856 , \10857 , \10858 , \10859 , \10860 , \10861 , \10862 , \10863 , \10864 ,
         \10865 , \10866 , \10867 , \10868 , \10869 , \10870 , \10871 , \10872 , \10873 , \10874 ,
         \10875 , \10876 , \10877 , \10878 , \10879 , \10880 , \10881 , \10882 , \10883 , \10884 ,
         \10885 , \10886 , \10887 , \10888 , \10889 , \10890 , \10891 , \10892 , \10893 , \10894 ,
         \10895 , \10896 , \10897 , \10898 , \10899 , \10900 , \10901 , \10902 , \10903 , \10904 ,
         \10905 , \10906 , \10907 , \10908 , \10909 , \10910 , \10911 , \10912 , \10913 , \10914 ,
         \10915 , \10916 , \10917 , \10918 , \10919 , \10920 , \10921 , \10922 , \10923 , \10924 ,
         \10925 , \10926 , \10927 , \10928 , \10929 , \10930 , \10931 , \10932 , \10933 , \10934 ,
         \10935 , \10936 , \10937 , \10938 , \10939 , \10940 , \10941 , \10942 , \10943 , \10944 ,
         \10945 , \10946 , \10947 , \10948 , \10949 , \10950 , \10951 , \10952 , \10953 , \10954 ,
         \10955 , \10956 , \10957 , \10958 , \10959 , \10960 , \10961 , \10962 , \10963 , \10964 ,
         \10965 , \10966 , \10967 , \10968 , \10969 , \10970 , \10971 , \10972 , \10973 , \10974 ,
         \10975 , \10976 , \10977 , \10978 , \10979 , \10980 , \10981 , \10982 , \10983 , \10984 ,
         \10985 , \10986 , \10987 , \10988 , \10989 , \10990 , \10991 , \10992 , \10993 , \10994 ,
         \10995 , \10996 , \10997 , \10998 , \10999 , \11000 , \11001 , \11002 , \11003 , \11004 ,
         \11005 , \11006 , \11007 , \11008 , \11009 , \11010 , \11011 , \11012 , \11013 , \11014 ,
         \11015 , \11016 , \11017 , \11018 , \11019 , \11020 , \11021 , \11022 , \11023 , \11024 ,
         \11025 , \11026 , \11027 , \11028 , \11029 , \11030 , \11031 , \11032 , \11033 , \11034 ,
         \11035 , \11036 , \11037 , \11038 , \11039 , \11040 , \11041 , \11042 , \11043 , \11044 ,
         \11045 , \11046 , \11047 , \11048 , \11049 , \11050 , \11051 , \11052 , \11053 , \11054 ,
         \11055 , \11056 , \11057 , \11058 , \11059 , \11060 , \11061 , \11062 , \11063 , \11064 ,
         \11065 , \11066 , \11067 , \11068 , \11069 , \11070 , \11071 , \11072 , \11073 , \11074 ,
         \11075 , \11076 , \11077 , \11078 , \11079 , \11080 , \11081 , \11082 , \11083 , \11084 ,
         \11085 , \11086 , \11087 , \11088 , \11089 , \11090 , \11091 , \11092 , \11093 , \11094 ,
         \11095 , \11096 , \11097 , \11098 , \11099 , \11100 , \11101 , \11102 , \11103 , \11104 ,
         \11105 , \11106 , \11107 , \11108 , \11109 , \11110 , \11111 , \11112 , \11113 , \11114 ,
         \11115 , \11116 , \11117 , \11118 , \11119 , \11120 , \11121 , \11122 , \11123 , \11124 ,
         \11125 , \11126 , \11127 , \11128 , \11129 , \11130 , \11131 , \11132 , \11133 , \11134 ,
         \11135 , \11136 , \11137 , \11138 , \11139 , \11140 , \11141 , \11142 , \11143 , \11144 ,
         \11145 , \11146 , \11147 , \11148 , \11149 , \11150 , \11151 , \11152 , \11153 , \11154 ,
         \11155 , \11156 , \11157 , \11158 , \11159 , \11160 , \11161 , \11162 , \11163 , \11164 ,
         \11165 , \11166 , \11167 , \11168 , \11169 , \11170 , \11171 , \11172 , \11173 , \11174 ,
         \11175 , \11176 , \11177 , \11178 , \11179 , \11180 , \11181 , \11182 , \11183 , \11184 ,
         \11185 , \11186 , \11187 , \11188 , \11189 , \11190 , \11191 , \11192 , \11193 , \11194 ,
         \11195 , \11196 , \11197 , \11198 , \11199 , \11200 , \11201 , \11202 , \11203 , \11204 ,
         \11205 , \11206 , \11207 , \11208 , \11209 , \11210 , \11211 , \11212 , \11213 , \11214 ,
         \11215 , \11216 , \11217 , \11218 , \11219 , \11220 , \11221 , \11222 , \11223 , \11224 ,
         \11225 , \11226 , \11227 , \11228 , \11229 , \11230 , \11231 , \11232 , \11233 , \11234 ,
         \11235 , \11236 , \11237 , \11238 , \11239 , \11240 , \11241 , \11242 , \11243 , \11244 ,
         \11245 , \11246 , \11247 , \11248 , \11249 , \11250 , \11251 , \11252 , \11253 , \11254 ,
         \11255 , \11256 , \11257 , \11258 , \11259 , \11260 , \11261 , \11262 , \11263 , \11264 ,
         \11265 , \11266 , \11267 , \11268 , \11269 , \11270 , \11271 , \11272 , \11273 , \11274 ,
         \11275 , \11276 , \11277 , \11278 , \11279 , \11280 , \11281 , \11282 , \11283 , \11284 ,
         \11285 , \11286 , \11287 , \11288 , \11289 , \11290 , \11291 , \11292 , \11293 , \11294 ,
         \11295 , \11296 , \11297 , \11298 , \11299 , \11300 , \11301 , \11302 , \11303 , \11304 ,
         \11305 , \11306 , \11307 , \11308 , \11309 , \11310 , \11311 , \11312 , \11313 , \11314 ,
         \11315 , \11316 , \11317 , \11318 , \11319 , \11320 , \11321 , \11322 , \11323 , \11324 ,
         \11325 , \11326 , \11327 , \11328 , \11329 , \11330 , \11331 , \11332 , \11333 , \11334 ,
         \11335 , \11336 , \11337 , \11338 , \11339 , \11340 , \11341 , \11342 , \11343 , \11344 ,
         \11345 , \11346 , \11347 , \11348 , \11349 , \11350 , \11351 , \11352 , \11353 , \11354 ,
         \11355 , \11356 , \11357 , \11358 , \11359 , \11360 , \11361 , \11362 , \11363 , \11364 ,
         \11365 , \11366 , \11367 , \11368 , \11369 , \11370 , \11371 , \11372 , \11373 , \11374 ,
         \11375 , \11376 , \11377 , \11378 , \11379 , \11380 , \11381 , \11382 , \11383 , \11384 ,
         \11385 , \11386 , \11387 , \11388 , \11389 , \11390 , \11391 , \11392 , \11393 , \11394 ,
         \11395 , \11396 , \11397 , \11398 , \11399 , \11400 , \11401 , \11402 , \11403 , \11404 ,
         \11405 , \11406 , \11407 , \11408 , \11409 , \11410 , \11411 , \11412 , \11413 , \11414 ,
         \11415 , \11416 , \11417 , \11418 , \11419 , \11420 , \11421 , \11422 , \11423 , \11424 ,
         \11425 , \11426 , \11427 , \11428 , \11429 , \11430 , \11431 , \11432 , \11433 , \11434 ,
         \11435 , \11436 , \11437 , \11438 , \11439 , \11440 , \11441 , \11442 , \11443 , \11444 ,
         \11445 , \11446 , \11447 , \11448 , \11449 , \11450 , \11451 , \11452 , \11453 , \11454 ,
         \11455 , \11456 , \11457 , \11458 , \11459 , \11460 , \11461 , \11462 , \11463 , \11464 ,
         \11465 , \11466 , \11467 , \11468 , \11469 , \11470 , \11471 , \11472 , \11473 , \11474 ,
         \11475 , \11476 , \11477 , \11478 , \11479 , \11480 , \11481 , \11482 , \11483 , \11484 ,
         \11485 , \11486 , \11487 , \11488 , \11489 , \11490 , \11491 , \11492 , \11493 , \11494 ,
         \11495 , \11496 , \11497 , \11498 , \11499 , \11500 , \11501 , \11502 , \11503 , \11504 ,
         \11505 , \11506 , \11507 , \11508 , \11509 , \11510 , \11511 , \11512 , \11513 , \11514 ,
         \11515 , \11516 , \11517 , \11518 , \11519 , \11520 , \11521 , \11522 , \11523 , \11524 ,
         \11525 , \11526 , \11527 , \11528 , \11529 , \11530 , \11531 , \11532 , \11533 , \11534 ,
         \11535 , \11536 , \11537 , \11538 , \11539 , \11540 , \11541 , \11542 , \11543 , \11544 ,
         \11545 , \11546 , \11547 , \11548 , \11549 , \11550 , \11551 , \11552 , \11553 , \11554 ,
         \11555 , \11556 , \11557 , \11558 , \11559 , \11560 , \11561 , \11562 , \11563 , \11564 ,
         \11565 , \11566 , \11567 , \11568 , \11569 , \11570 , \11571 , \11572 , \11573 , \11574 ,
         \11575 , \11576 , \11577 , \11578 , \11579 , \11580 , \11581 , \11582 , \11583 , \11584 ,
         \11585 , \11586 , \11587 , \11588 , \11589 , \11590 , \11591 , \11592 , \11593 , \11594 ,
         \11595 , \11596 , \11597 , \11598 , \11599 , \11600 , \11601 , \11602 , \11603 , \11604 ,
         \11605 , \11606 , \11607 , \11608 , \11609 , \11610 , \11611 , \11612 , \11613 , \11614 ,
         \11615 , \11616 , \11617 , \11618 , \11619 , \11620 , \11621 , \11622 , \11623 , \11624 ,
         \11625 , \11626 , \11627 , \11628 , \11629 , \11630 , \11631 , \11632 , \11633 , \11634 ,
         \11635 , \11636 , \11637 , \11638 , \11639 , \11640 , \11641 , \11642 , \11643 , \11644 ,
         \11645 , \11646 , \11647 , \11648 , \11649 , \11650 , \11651 , \11652 , \11653 , \11654 ,
         \11655 , \11656 , \11657 , \11658 , \11659 , \11660 , \11661 , \11662 , \11663 , \11664 ,
         \11665 , \11666 , \11667 , \11668 , \11669 , \11670 , \11671 , \11672 , \11673 , \11674 ,
         \11675 , \11676 , \11677 , \11678 , \11679 , \11680 , \11681 , \11682 , \11683 , \11684 ,
         \11685 , \11686 , \11687 , \11688 , \11689 , \11690 , \11691 , \11692 , \11693 , \11694 ,
         \11695 , \11696 , \11697 , \11698 , \11699 , \11700 , \11701 , \11702 , \11703 , \11704 ,
         \11705 , \11706 , \11707 , \11708 , \11709 , \11710 , \11711 , \11712 , \11713 , \11714 ,
         \11715 , \11716 , \11717 , \11718 , \11719 , \11720 , \11721 , \11722 , \11723 , \11724 ,
         \11725 , \11726 , \11727 , \11728 , \11729 , \11730 , \11731 , \11732 , \11733 , \11734 ,
         \11735 , \11736 , \11737 , \11738 , \11739 , \11740 , \11741 , \11742 , \11743 , \11744 ,
         \11745 , \11746 , \11747 , \11748 , \11749 , \11750 , \11751 , \11752 , \11753 , \11754 ,
         \11755 , \11756 , \11757 , \11758 , \11759 , \11760 , \11761 , \11762 , \11763 , \11764 ,
         \11765 , \11766 , \11767 , \11768 , \11769 , \11770 , \11771 , \11772 , \11773 , \11774 ,
         \11775 , \11776 , \11777 , \11778 , \11779 , \11780 , \11781 , \11782 , \11783 , \11784 ,
         \11785 , \11786 , \11787 , \11788 , \11789 , \11790 , \11791 , \11792 , \11793 , \11794 ,
         \11795 , \11796 , \11797 , \11798 , \11799 , \11800 , \11801 , \11802 , \11803 , \11804 ,
         \11805 , \11806 , \11807 , \11808 , \11809 , \11810 , \11811 , \11812 , \11813 , \11814 ,
         \11815 , \11816 , \11817 , \11818 , \11819 , \11820 , \11821 , \11822 , \11823 , \11824 ,
         \11825 , \11826 , \11827 , \11828 , \11829 , \11830 , \11831 , \11832 , \11833 , \11834 ,
         \11835 , \11836 , \11837 , \11838 , \11839 , \11840 , \11841 , \11842 , \11843 , \11844 ,
         \11845 , \11846 , \11847 , \11848 , \11849 , \11850 , \11851 , \11852 , \11853 , \11854 ,
         \11855 , \11856 , \11857 , \11858 , \11859 , \11860 , \11861 , \11862 , \11863 , \11864 ,
         \11865 , \11866 , \11867 , \11868 , \11869 , \11870 , \11871 , \11872 , \11873 , \11874 ,
         \11875 , \11876 , \11877 , \11878 , \11879 , \11880 , \11881 , \11882 , \11883 , \11884 ,
         \11885 , \11886 , \11887 , \11888 , \11889 , \11890 , \11891 , \11892 , \11893 , \11894 ,
         \11895 , \11896 , \11897 , \11898 , \11899 , \11900 , \11901 , \11902 , \11903 , \11904 ,
         \11905 , \11906 , \11907 , \11908 , \11909 , \11910 , \11911 , \11912 , \11913 , \11914 ,
         \11915 , \11916 , \11917 , \11918 , \11919 , \11920 , \11921 , \11922 , \11923 , \11924 ,
         \11925 , \11926 , \11927 , \11928 , \11929 , \11930 , \11931 , \11932 , \11933 , \11934 ,
         \11935 , \11936 , \11937 , \11938 , \11939 , \11940 , \11941 , \11942 , \11943 , \11944 ,
         \11945 , \11946 , \11947 , \11948 , \11949 , \11950 , \11951 , \11952 , \11953 , \11954 ,
         \11955 , \11956 , \11957 , \11958 , \11959 , \11960 , \11961 , \11962 , \11963 , \11964 ,
         \11965 , \11966 , \11967 , \11968 , \11969 , \11970 , \11971 , \11972 , \11973 , \11974 ,
         \11975 , \11976 , \11977 , \11978 , \11979 , \11980 , \11981 , \11982 , \11983 , \11984 ,
         \11985 , \11986 , \11987 , \11988 , \11989 , \11990 , \11991 , \11992 , \11993 , \11994 ,
         \11995 , \11996 , \11997 , \11998 , \11999 , \12000 , \12001 , \12002 , \12003 , \12004 ,
         \12005 , \12006 , \12007 , \12008 , \12009 , \12010 , \12011 , \12012 , \12013 , \12014 ,
         \12015 , \12016 , \12017 , \12018 , \12019 , \12020 , \12021 , \12022 , \12023 , \12024 ,
         \12025 , \12026 , \12027 , \12028 , \12029 , \12030 , \12031 , \12032 , \12033 , \12034 ,
         \12035 , \12036 , \12037 , \12038 , \12039 , \12040 , \12041 , \12042 , \12043 , \12044 ,
         \12045 , \12046 , \12047 , \12048 , \12049 , \12050 , \12051 , \12052 , \12053 , \12054 ,
         \12055 , \12056 , \12057 , \12058 , \12059 , \12060 , \12061 , \12062 , \12063 , \12064 ,
         \12065 , \12066 , \12067 , \12068 , \12069 , \12070 , \12071 , \12072 , \12073 , \12074 ,
         \12075 , \12076 , \12077 , \12078 , \12079 , \12080 , \12081 , \12082 , \12083 , \12084 ,
         \12085 , \12086 , \12087 , \12088 , \12089 , \12090 , \12091 , \12092 , \12093 , \12094 ,
         \12095 , \12096 , \12097 , \12098 , \12099 , \12100 , \12101 , \12102 , \12103 , \12104 ,
         \12105 , \12106 , \12107 , \12108 , \12109 , \12110 , \12111 , \12112 , \12113 , \12114 ,
         \12115 , \12116 , \12117 , \12118 , \12119 , \12120 , \12121 , \12122 , \12123 , \12124 ,
         \12125 , \12126 , \12127 , \12128 , \12129 , \12130 , \12131 , \12132 , \12133 , \12134 ,
         \12135 , \12136 , \12137 , \12138 , \12139 , \12140 , \12141 , \12142 , \12143 , \12144 ,
         \12145 , \12146 , \12147 , \12148 , \12149 , \12150 , \12151 , \12152 , \12153 , \12154 ,
         \12155 , \12156 , \12157 , \12158 , \12159 , \12160 , \12161 , \12162 , \12163 , \12164 ,
         \12165 , \12166 , \12167 , \12168 , \12169 , \12170 , \12171 , \12172 , \12173 , \12174 ,
         \12175 , \12176 , \12177 , \12178 , \12179 , \12180 , \12181 , \12182 , \12183 , \12184 ,
         \12185 , \12186 , \12187 , \12188 , \12189 , \12190 , \12191 , \12192 , \12193 , \12194 ,
         \12195 , \12196 , \12197 , \12198 , \12199 , \12200 , \12201 , \12202 , \12203 , \12204 ,
         \12205 , \12206 , \12207 , \12208 , \12209 , \12210 , \12211 , \12212 , \12213 , \12214 ,
         \12215 , \12216 , \12217 , \12218 , \12219 , \12220 , \12221 , \12222 , \12223 , \12224 ,
         \12225 , \12226 , \12227 , \12228 , \12229 , \12230 , \12231 , \12232 , \12233 , \12234 ,
         \12235 , \12236 , \12237 , \12238 , \12239 , \12240 , \12241 , \12242 , \12243 , \12244 ,
         \12245 , \12246 , \12247 , \12248 , \12249 , \12250 , \12251 , \12252 , \12253 , \12254 ,
         \12255 , \12256 , \12257 , \12258 , \12259 , \12260 , \12261 , \12262 , \12263 , \12264 ,
         \12265 , \12266 , \12267 , \12268 , \12269 , \12270 , \12271 , \12272 , \12273 , \12274 ,
         \12275 , \12276 , \12277 , \12278 , \12279 , \12280 , \12281 , \12282 , \12283 , \12284 ,
         \12285 , \12286 , \12287 , \12288 , \12289 , \12290 , \12291 , \12292 , \12293 , \12294 ,
         \12295 , \12296 , \12297 , \12298 , \12299 , \12300 , \12301 , \12302 , \12303 , \12304 ,
         \12305 , \12306 , \12307 , \12308 , \12309 , \12310 , \12311 , \12312 , \12313 , \12314 ,
         \12315 , \12316 , \12317 , \12318 , \12319 , \12320 , \12321 , \12322 , \12323 , \12324 ,
         \12325 , \12326 , \12327 , \12328 , \12329 , \12330 , \12331 , \12332 , \12333 , \12334 ,
         \12335 , \12336 , \12337 , \12338 , \12339 , \12340 , \12341 , \12342 , \12343 , \12344 ,
         \12345 , \12346 , \12347 , \12348 , \12349 , \12350 , \12351 , \12352 , \12353 , \12354 ,
         \12355 , \12356 , \12357 , \12358 , \12359 , \12360 , \12361 , \12362 , \12363 , \12364 ,
         \12365 , \12366 , \12367 , \12368 , \12369 , \12370 , \12371 , \12372 , \12373 , \12374 ,
         \12375 , \12376 , \12377 , \12378 , \12379 , \12380 , \12381 , \12382 , \12383 , \12384 ,
         \12385 , \12386 , \12387 , \12388 , \12389 , \12390 , \12391 , \12392 , \12393 , \12394 ,
         \12395 , \12396 , \12397 , \12398 , \12399 , \12400 , \12401 , \12402 , \12403 , \12404 ,
         \12405 , \12406 , \12407 , \12408 , \12409 , \12410 , \12411 , \12412 , \12413 , \12414 ,
         \12415 , \12416 , \12417 , \12418 , \12419 , \12420 , \12421 , \12422 , \12423 , \12424 ,
         \12425 , \12426 , \12427 , \12428 , \12429 , \12430 , \12431 , \12432 , \12433 , \12434 ,
         \12435 , \12436 , \12437 , \12438 , \12439 , \12440 , \12441 , \12442 , \12443 , \12444 ,
         \12445 , \12446 , \12447 , \12448 , \12449 , \12450 , \12451 , \12452 , \12453 , \12454 ,
         \12455 , \12456 , \12457 , \12458 , \12459 , \12460 , \12461 , \12462 , \12463 , \12464 ,
         \12465 , \12466 , \12467 , \12468 , \12469 , \12470 , \12471 , \12472 , \12473 , \12474 ,
         \12475 , \12476 , \12477 , \12478 , \12479 , \12480 , \12481 , \12482 , \12483 , \12484 ,
         \12485 , \12486 , \12487 , \12488 , \12489 , \12490 , \12491 , \12492 , \12493 , \12494 ,
         \12495 , \12496 , \12497 , \12498 , \12499 , \12500 , \12501 , \12502 , \12503 , \12504 ,
         \12505 , \12506 , \12507 , \12508 , \12509 , \12510 , \12511 , \12512 , \12513 , \12514 ,
         \12515 , \12516 , \12517 , \12518 , \12519 , \12520 , \12521 , \12522 , \12523 , \12524 ,
         \12525 , \12526 , \12527 , \12528 , \12529 , \12530 , \12531 , \12532 , \12533 , \12534 ,
         \12535 , \12536 , \12537 , \12538 , \12539 , \12540 , \12541 , \12542 , \12543 , \12544 ,
         \12545 , \12546 , \12547 , \12548 , \12549 , \12550 , \12551 , \12552 , \12553 , \12554 ,
         \12555 , \12556 , \12557 , \12558 , \12559 , \12560 , \12561 , \12562 , \12563 , \12564 ,
         \12565 , \12566 , \12567 , \12568 , \12569 , \12570 , \12571 , \12572 , \12573 , \12574 ,
         \12575 , \12576 , \12577 , \12578 , \12579 , \12580 , \12581 , \12582 , \12583 , \12584 ,
         \12585 , \12586 , \12587 , \12588 , \12589 , \12590 , \12591 , \12592 , \12593 , \12594 ,
         \12595 , \12596 , \12597 , \12598 , \12599 , \12600 , \12601 , \12602 , \12603 , \12604 ,
         \12605 , \12606 , \12607 , \12608 , \12609 , \12610 , \12611 , \12612 , \12613 , \12614 ,
         \12615 , \12616 , \12617 , \12618 , \12619 , \12620 , \12621 , \12622 , \12623 , \12624 ,
         \12625 , \12626 , \12627 , \12628 , \12629 , \12630 , \12631 , \12632 , \12633 , \12634 ,
         \12635 , \12636 , \12637 , \12638 , \12639 , \12640 , \12641 , \12642 , \12643 , \12644 ,
         \12645 , \12646 , \12647 , \12648 , \12649 , \12650 , \12651 , \12652 , \12653 , \12654 ,
         \12655 , \12656 , \12657 , \12658 , \12659 , \12660 , \12661 , \12662 , \12663 , \12664 ,
         \12665 , \12666 , \12667 , \12668 , \12669 , \12670 , \12671 , \12672 , \12673 , \12674 ,
         \12675 , \12676 , \12677 , \12678 , \12679 , \12680 , \12681 , \12682 , \12683 , \12684 ,
         \12685 , \12686 , \12687 , \12688 , \12689 , \12690 , \12691 , \12692 , \12693 , \12694 ,
         \12695 , \12696 , \12697 , \12698 , \12699 , \12700 , \12701 , \12702 , \12703 , \12704 ,
         \12705 , \12706 , \12707 , \12708 , \12709 , \12710 , \12711 , \12712 , \12713 , \12714 ,
         \12715 , \12716 , \12717 , \12718 , \12719 , \12720 , \12721 , \12722 , \12723 , \12724 ,
         \12725 , \12726 , \12727 , \12728 , \12729 , \12730 , \12731 , \12732 , \12733 , \12734 ,
         \12735 , \12736 , \12737 , \12738 , \12739 , \12740 , \12741 , \12742 , \12743 , \12744 ,
         \12745 , \12746 , \12747 , \12748 , \12749 , \12750 , \12751 , \12752 , \12753 , \12754 ,
         \12755 , \12756 , \12757 , \12758 , \12759 , \12760 , \12761 , \12762 , \12763 , \12764 ,
         \12765 , \12766 , \12767 , \12768 , \12769 , \12770 , \12771 , \12772 , \12773 , \12774 ,
         \12775 , \12776 , \12777 , \12778 , \12779 , \12780 , \12781 , \12782 , \12783 , \12784 ,
         \12785 , \12786 , \12787 , \12788 , \12789 , \12790 , \12791 , \12792 , \12793 , \12794 ,
         \12795 , \12796 , \12797 , \12798 , \12799 , \12800 , \12801 , \12802 , \12803 , \12804 ,
         \12805 , \12806 , \12807 , \12808 , \12809 , \12810 , \12811 , \12812 , \12813 , \12814 ,
         \12815 , \12816 , \12817 , \12818 , \12819 , \12820 , \12821 , \12822 , \12823 , \12824 ,
         \12825 , \12826 , \12827 , \12828 , \12829 , \12830 , \12831 , \12832 , \12833 , \12834 ,
         \12835 , \12836 , \12837 , \12838 , \12839 , \12840 , \12841 , \12842 , \12843 , \12844 ,
         \12845 , \12846 , \12847 , \12848 , \12849 , \12850 , \12851 , \12852 , \12853 , \12854 ,
         \12855 , \12856 , \12857 , \12858 , \12859 , \12860 , \12861 , \12862 , \12863 , \12864 ,
         \12865 , \12866 , \12867 , \12868 , \12869 , \12870 , \12871 , \12872 , \12873 , \12874 ,
         \12875 , \12876 , \12877 , \12878 , \12879 , \12880 , \12881 , \12882 , \12883 , \12884 ,
         \12885 , \12886 , \12887 , \12888 , \12889 , \12890 , \12891 , \12892 , \12893 , \12894 ,
         \12895 , \12896 , \12897 , \12898 , \12899 , \12900 , \12901 , \12902 , \12903 , \12904 ,
         \12905 , \12906 , \12907 , \12908 , \12909 , \12910 , \12911 , \12912 , \12913 , \12914 ,
         \12915 , \12916 , \12917 , \12918 , \12919 , \12920 , \12921 , \12922 , \12923 , \12924 ,
         \12925 , \12926 , \12927 , \12928 , \12929 , \12930 , \12931 , \12932 , \12933 , \12934 ,
         \12935 , \12936 , \12937 , \12938 , \12939 , \12940 , \12941 , \12942 , \12943 , \12944 ,
         \12945 , \12946 , \12947 , \12948 , \12949 , \12950 , \12951 , \12952 , \12953 , \12954 ,
         \12955 , \12956 , \12957 , \12958 , \12959 , \12960 , \12961 , \12962 , \12963 , \12964 ,
         \12965 , \12966 , \12967 , \12968 , \12969 , \12970 , \12971 , \12972 , \12973 , \12974 ,
         \12975 , \12976 , \12977 , \12978 , \12979 , \12980 , \12981 , \12982 , \12983 , \12984 ,
         \12985 , \12986 , \12987 , \12988 , \12989 , \12990 , \12991 , \12992 , \12993 , \12994 ,
         \12995 , \12996 , \12997 , \12998 , \12999 , \13000 , \13001 , \13002 , \13003 , \13004 ,
         \13005 , \13006 , \13007 , \13008 , \13009 , \13010 , \13011 , \13012 , \13013 , \13014 ,
         \13015 , \13016 , \13017 , \13018 , \13019 , \13020 , \13021 , \13022 , \13023 , \13024 ,
         \13025 , \13026 , \13027 , \13028 , \13029 , \13030 , \13031 , \13032 , \13033 , \13034 ,
         \13035 , \13036 , \13037 , \13038 , \13039 , \13040 , \13041 , \13042 , \13043 , \13044 ,
         \13045 , \13046 , \13047 , \13048 , \13049 , \13050 , \13051 , \13052 , \13053 , \13054 ,
         \13055 , \13056 , \13057 , \13058 , \13059 , \13060 , \13061 , \13062 , \13063 , \13064 ,
         \13065 , \13066 , \13067 , \13068 , \13069 , \13070 , \13071 , \13072 , \13073 , \13074 ,
         \13075 , \13076 , \13077 , \13078 , \13079 , \13080 , \13081 , \13082 , \13083 , \13084 ,
         \13085 , \13086 , \13087 , \13088 , \13089 , \13090 , \13091 , \13092 , \13093 , \13094 ,
         \13095 , \13096 , \13097 , \13098 , \13099 , \13100 , \13101 , \13102 , \13103 , \13104 ,
         \13105 , \13106 , \13107 , \13108 , \13109 , \13110 , \13111 , \13112 , \13113 , \13114 ,
         \13115 , \13116 , \13117 , \13118 , \13119 , \13120 , \13121 , \13122 , \13123 , \13124 ,
         \13125 , \13126 , \13127 , \13128 , \13129 , \13130 , \13131 , \13132 , \13133 , \13134 ,
         \13135 , \13136 , \13137 , \13138 , \13139 , \13140 , \13141 , \13142 , \13143 , \13144 ,
         \13145 , \13146 , \13147 , \13148 , \13149 , \13150 , \13151 , \13152 , \13153 , \13154 ,
         \13155 , \13156 , \13157 , \13158 , \13159 , \13160 , \13161 , \13162 , \13163 , \13164 ,
         \13165 , \13166 , \13167 , \13168 , \13169 , \13170 , \13171 , \13172 , \13173 , \13174 ,
         \13175 , \13176 , \13177 , \13178 , \13179 , \13180 , \13181 , \13182 , \13183 , \13184 ,
         \13185 , \13186 , \13187 , \13188 , \13189 , \13190 , \13191 , \13192 , \13193 , \13194 ,
         \13195 , \13196 , \13197 , \13198 , \13199 , \13200 , \13201 , \13202 , \13203 , \13204 ,
         \13205 , \13206 , \13207 , \13208 , \13209 , \13210 , \13211 , \13212 , \13213 , \13214 ,
         \13215 , \13216 , \13217 , \13218 , \13219 , \13220 , \13221 , \13222 , \13223 , \13224 ,
         \13225 , \13226 , \13227 , \13228 , \13229 , \13230 , \13231 , \13232 , \13233 , \13234 ,
         \13235 , \13236 , \13237 , \13238 , \13239 , \13240 , \13241 , \13242 , \13243 , \13244 ,
         \13245 , \13246 , \13247 , \13248 , \13249 , \13250 , \13251 , \13252 , \13253 , \13254 ,
         \13255 , \13256 , \13257 , \13258 , \13259 , \13260 , \13261 , \13262 , \13263 , \13264 ,
         \13265 , \13266 , \13267 , \13268 , \13269 , \13270 , \13271 , \13272 , \13273 , \13274 ,
         \13275 , \13276 , \13277 , \13278 , \13279 , \13280 , \13281 , \13282 , \13283 , \13284 ,
         \13285 , \13286 , \13287 , \13288 , \13289 , \13290 , \13291 , \13292 , \13293 , \13294 ,
         \13295 , \13296 , \13297 , \13298 , \13299 , \13300 , \13301 , \13302 , \13303 , \13304 ,
         \13305 , \13306 , \13307 , \13308 , \13309 , \13310 , \13311 , \13312 , \13313 , \13314 ,
         \13315 , \13316 , \13317 , \13318 , \13319 , \13320 , \13321 , \13322 , \13323 , \13324 ,
         \13325 , \13326 , \13327 , \13328 , \13329 , \13330 , \13331 , \13332 , \13333 , \13334 ,
         \13335 , \13336 , \13337 , \13338 , \13339 , \13340 , \13341 , \13342 , \13343 , \13344 ,
         \13345 , \13346 , \13347 , \13348 , \13349 , \13350 , \13351 , \13352 , \13353 , \13354 ,
         \13355 , \13356 , \13357 , \13358 , \13359 , \13360 , \13361 , \13362 , \13363 , \13364 ,
         \13365 , \13366 , \13367 , \13368 , \13369 , \13370 , \13371 , \13372 , \13373 , \13374 ,
         \13375 , \13376 , \13377 , \13378 , \13379 , \13380 , \13381 , \13382 , \13383 , \13384 ,
         \13385 , \13386 , \13387 , \13388 , \13389 , \13390 , \13391 , \13392 , \13393 , \13394 ,
         \13395 , \13396 , \13397 , \13398 , \13399 , \13400 , \13401 , \13402 , \13403 , \13404 ,
         \13405 , \13406 , \13407 , \13408 , \13409 , \13410 , \13411 , \13412 , \13413 , \13414 ,
         \13415 , \13416 , \13417 , \13418 , \13419 , \13420 , \13421 , \13422 , \13423 , \13424 ,
         \13425 , \13426 , \13427 , \13428 , \13429 , \13430 , \13431 , \13432 , \13433 , \13434 ,
         \13435 , \13436 , \13437 , \13438 , \13439 , \13440 , \13441 , \13442 , \13443 , \13444 ,
         \13445 , \13446 , \13447 , \13448 , \13449 , \13450 , \13451 , \13452 , \13453 , \13454 ,
         \13455 , \13456 , \13457 , \13458 , \13459 , \13460 , \13461 , \13462 , \13463 , \13464 ,
         \13465 , \13466 , \13467 , \13468 , \13469 , \13470 , \13471 , \13472 , \13473 , \13474 ,
         \13475 , \13476 , \13477 , \13478 , \13479 , \13480 , \13481 , \13482 , \13483 , \13484 ,
         \13485 , \13486 , \13487 , \13488 , \13489 , \13490 , \13491 , \13492 , \13493 , \13494 ,
         \13495 , \13496 , \13497 , \13498 , \13499 , \13500 , \13501 , \13502 , \13503 , \13504 ,
         \13505 , \13506 , \13507 , \13508 , \13509 , \13510 , \13511 , \13512 , \13513 , \13514 ,
         \13515 , \13516 , \13517 , \13518 , \13519 , \13520 , \13521 , \13522 , \13523 , \13524 ,
         \13525 , \13526 , \13527 , \13528 , \13529 , \13530 , \13531 , \13532 , \13533 , \13534 ,
         \13535 , \13536 , \13537 , \13538 , \13539 , \13540 , \13541 , \13542 , \13543 , \13544 ,
         \13545 , \13546 , \13547 , \13548 , \13549 , \13550 , \13551 , \13552 , \13553 , \13554 ,
         \13555 , \13556 , \13557 , \13558 , \13559 , \13560 , \13561 , \13562 , \13563 , \13564 ,
         \13565 , \13566 , \13567 , \13568 , \13569 , \13570 , \13571 , \13572 , \13573 , \13574 ,
         \13575 , \13576 , \13577 , \13578 , \13579 , \13580 , \13581 , \13582 , \13583 , \13584 ,
         \13585 , \13586 , \13587 , \13588 , \13589 , \13590 , \13591 , \13592 , \13593 , \13594 ,
         \13595 , \13596 , \13597 , \13598 , \13599 , \13600 , \13601 , \13602 , \13603 , \13604 ,
         \13605 , \13606 , \13607 , \13608 , \13609 , \13610 , \13611 , \13612 , \13613 , \13614 ,
         \13615 , \13616 , \13617 , \13618 , \13619 , \13620 , \13621 , \13622 , \13623 , \13624 ,
         \13625 , \13626 , \13627 , \13628 , \13629 , \13630 , \13631 , \13632 , \13633 , \13634 ,
         \13635 , \13636 , \13637 , \13638 , \13639 , \13640 , \13641 , \13642 , \13643 , \13644 ,
         \13645 , \13646 , \13647 , \13648 , \13649 , \13650 , \13651 , \13652 , \13653 , \13654 ,
         \13655 , \13656 , \13657 , \13658 , \13659 , \13660 , \13661 , \13662 , \13663 , \13664 ,
         \13665 , \13666 , \13667 , \13668 , \13669 , \13670 , \13671 , \13672 , \13673 , \13674 ,
         \13675 , \13676 , \13677 , \13678 , \13679 , \13680 , \13681 , \13682 , \13683 , \13684 ,
         \13685 , \13686 , \13687 , \13688 , \13689 , \13690 , \13691 , \13692 , \13693 , \13694 ,
         \13695 , \13696 , \13697 , \13698 , \13699 , \13700 , \13701 , \13702 , \13703 , \13704 ,
         \13705 , \13706 , \13707 , \13708 , \13709 , \13710 , \13711 , \13712 , \13713 , \13714 ,
         \13715 , \13716 , \13717 , \13718 , \13719 , \13720 , \13721 , \13722 , \13723 , \13724 ,
         \13725 , \13726 , \13727 , \13728 , \13729 , \13730 , \13731 , \13732 , \13733 , \13734 ,
         \13735 , \13736 , \13737 , \13738 , \13739 , \13740 , \13741 , \13742 , \13743 , \13744 ,
         \13745 , \13746 , \13747 , \13748 , \13749 , \13750 , \13751 , \13752 , \13753 , \13754 ,
         \13755 , \13756 , \13757 , \13758 , \13759 , \13760 , \13761 , \13762 , \13763 , \13764 ,
         \13765 , \13766 , \13767 , \13768 , \13769 , \13770 , \13771 , \13772 , \13773 , \13774 ,
         \13775 , \13776 , \13777 , \13778 , \13779 , \13780 , \13781 , \13782 , \13783 , \13784 ,
         \13785 , \13786 , \13787 , \13788 , \13789 , \13790 , \13791 , \13792 , \13793 , \13794 ,
         \13795 , \13796 , \13797 , \13798 , \13799 , \13800 , \13801 , \13802 , \13803 , \13804 ,
         \13805 , \13806 , \13807 , \13808 , \13809 , \13810 , \13811 , \13812 , \13813 , \13814 ,
         \13815 , \13816 , \13817 , \13818 , \13819 , \13820 , \13821 , \13822 , \13823 , \13824 ,
         \13825 , \13826 , \13827 , \13828 , \13829 , \13830 , \13831 , \13832 , \13833 , \13834 ,
         \13835 , \13836 , \13837 , \13838 , \13839 , \13840 , \13841 , \13842 , \13843 , \13844 ,
         \13845 , \13846 , \13847 , \13848 , \13849 , \13850 , \13851 , \13852 , \13853 , \13854 ,
         \13855 , \13856 , \13857 , \13858 , \13859 , \13860 , \13861 , \13862 , \13863 , \13864 ,
         \13865 , \13866 , \13867 , \13868 , \13869 , \13870 , \13871 , \13872 , \13873 , \13874 ,
         \13875 , \13876 , \13877 , \13878 , \13879 , \13880 , \13881 , \13882 , \13883 , \13884 ,
         \13885 , \13886 , \13887 , \13888 , \13889 , \13890 , \13891 , \13892 , \13893 , \13894 ,
         \13895 , \13896 , \13897 , \13898 , \13899 , \13900 , \13901 , \13902 , \13903 , \13904 ,
         \13905 , \13906 , \13907 , \13908 , \13909 , \13910 , \13911 , \13912 , \13913 , \13914 ,
         \13915 , \13916 , \13917 , \13918 , \13919 , \13920 , \13921 , \13922 , \13923 , \13924 ,
         \13925 , \13926 , \13927 , \13928 , \13929 , \13930 , \13931 , \13932 , \13933 , \13934 ,
         \13935 , \13936 , \13937 , \13938 , \13939 , \13940 , \13941 , \13942 , \13943 , \13944 ,
         \13945 , \13946 , \13947 , \13948 , \13949 , \13950 , \13951 , \13952 , \13953 , \13954 ,
         \13955 , \13956 , \13957 , \13958 , \13959 , \13960 , \13961 , \13962 , \13963 , \13964 ,
         \13965 , \13966 , \13967 , \13968 , \13969 , \13970 , \13971 , \13972 , \13973 , \13974 ,
         \13975 , \13976 , \13977 , \13978 , \13979 , \13980 , \13981 , \13982 , \13983 , \13984 ,
         \13985 , \13986 , \13987 , \13988 , \13989 , \13990 , \13991 , \13992 , \13993 , \13994 ,
         \13995 , \13996 , \13997 , \13998 , \13999 , \14000 , \14001 , \14002 , \14003 , \14004 ,
         \14005 , \14006 , \14007 , \14008 , \14009 , \14010 , \14011 , \14012 , \14013 , \14014 ,
         \14015 , \14016 , \14017 , \14018 , \14019 , \14020 , \14021 , \14022 , \14023 , \14024 ,
         \14025 , \14026 , \14027 , \14028 , \14029 , \14030 , \14031 , \14032 , \14033 , \14034 ,
         \14035 , \14036 , \14037 , \14038 , \14039 , \14040 , \14041 , \14042 , \14043 , \14044 ,
         \14045 , \14046 , \14047 , \14048 , \14049 , \14050 , \14051 , \14052 , \14053 , \14054 ,
         \14055 , \14056 , \14057 , \14058 , \14059 , \14060 , \14061 , \14062 , \14063 , \14064 ,
         \14065 , \14066 , \14067 , \14068 , \14069 , \14070 , \14071 , \14072 , \14073 , \14074 ,
         \14075 , \14076 , \14077 , \14078 , \14079 , \14080 , \14081 , \14082 , \14083 , \14084 ,
         \14085 , \14086 , \14087 , \14088 , \14089 , \14090 , \14091 , \14092 , \14093 , \14094 ,
         \14095 , \14096 , \14097 , \14098 , \14099 , \14100 , \14101 , \14102 , \14103 , \14104 ,
         \14105 , \14106 , \14107 , \14108 , \14109 , \14110 , \14111 , \14112 , \14113 , \14114 ,
         \14115 , \14116 , \14117 , \14118 , \14119 , \14120 , \14121 , \14122 , \14123 , \14124 ,
         \14125 , \14126 , \14127 , \14128 , \14129 , \14130 , \14131 , \14132 , \14133 , \14134 ,
         \14135 , \14136 , \14137 , \14138 , \14139 , \14140 , \14141 , \14142 , \14143 , \14144 ,
         \14145 , \14146 , \14147 , \14148 , \14149 , \14150 , \14151 , \14152 , \14153 , \14154 ,
         \14155 , \14156 , \14157 , \14158 , \14159 , \14160 , \14161 , \14162 , \14163 , \14164 ,
         \14165 , \14166 , \14167 , \14168 , \14169 , \14170 , \14171 , \14172 , \14173 , \14174 ,
         \14175 , \14176 , \14177 , \14178 , \14179 , \14180 , \14181 , \14182 , \14183 , \14184 ,
         \14185 , \14186 , \14187 , \14188 , \14189 , \14190 , \14191 , \14192 , \14193 , \14194 ,
         \14195 , \14196 , \14197 , \14198 , \14199 , \14200 , \14201 , \14202 , \14203 , \14204 ,
         \14205 , \14206 , \14207 , \14208 , \14209 , \14210 , \14211 , \14212 , \14213 , \14214 ,
         \14215 , \14216 , \14217 , \14218 , \14219 , \14220 , \14221 , \14222 , \14223 , \14224 ,
         \14225 , \14226 , \14227 , \14228 , \14229 , \14230 , \14231 , \14232 , \14233 , \14234 ,
         \14235 , \14236 , \14237 , \14238 , \14239 , \14240 , \14241 , \14242 , \14243 , \14244 ,
         \14245 , \14246 , \14247 , \14248 , \14249 , \14250 , \14251 , \14252 , \14253 , \14254 ,
         \14255 , \14256 , \14257 , \14258 , \14259 , \14260 , \14261 , \14262 , \14263 , \14264 ,
         \14265 , \14266 , \14267 , \14268 , \14269 , \14270 , \14271 , \14272 , \14273 , \14274 ,
         \14275 , \14276 , \14277 , \14278 , \14279 , \14280 , \14281 , \14282 , \14283 , \14284 ,
         \14285 , \14286 , \14287 , \14288 , \14289 , \14290 , \14291 , \14292 , \14293 , \14294 ,
         \14295 , \14296 , \14297 , \14298 , \14299 , \14300 , \14301 , \14302 , \14303 , \14304 ,
         \14305 , \14306 , \14307 , \14308 , \14309 , \14310 , \14311 , \14312 , \14313 , \14314 ,
         \14315 , \14316 , \14317 , \14318 , \14319 , \14320 , \14321 , \14322 , \14323 , \14324 ,
         \14325 , \14326 , \14327 , \14328 , \14329 , \14330 , \14331 , \14332 , \14333 , \14334 ,
         \14335 , \14336 , \14337 , \14338 , \14339 , \14340 , \14341 , \14342 , \14343 , \14344 ,
         \14345 , \14346 , \14347 , \14348 , \14349 , \14350 , \14351 , \14352 , \14353 , \14354 ,
         \14355 , \14356 , \14357 , \14358 , \14359 , \14360 , \14361 , \14362 , \14363 , \14364 ,
         \14365 , \14366 , \14367 , \14368 , \14369 , \14370 , \14371 , \14372 , \14373 , \14374 ,
         \14375 , \14376 , \14377 , \14378 , \14379 , \14380 , \14381 , \14382 , \14383 , \14384 ,
         \14385 , \14386 , \14387 , \14388 , \14389 , \14390 , \14391 , \14392 , \14393 , \14394 ,
         \14395 , \14396 , \14397 , \14398 , \14399 , \14400 , \14401 , \14402 , \14403 , \14404 ,
         \14405 , \14406 , \14407 , \14408 , \14409 , \14410 , \14411 , \14412 , \14413 , \14414 ,
         \14415 , \14416 , \14417 , \14418 , \14419 , \14420 , \14421 , \14422 , \14423 , \14424 ,
         \14425 , \14426 , \14427 , \14428 , \14429 , \14430 , \14431 , \14432 , \14433 , \14434 ,
         \14435 , \14436 , \14437 , \14438 , \14439 , \14440 , \14441 , \14442 , \14443 , \14444 ,
         \14445 , \14446 , \14447 , \14448 , \14449 , \14450 , \14451 , \14452 , \14453 , \14454 ,
         \14455 , \14456 , \14457 , \14458 , \14459 , \14460 , \14461 , \14462 , \14463 , \14464 ,
         \14465 , \14466 , \14467 , \14468 , \14469 , \14470 , \14471 , \14472 , \14473 , \14474 ,
         \14475 , \14476 , \14477 , \14478 , \14479 , \14480 , \14481 , \14482 , \14483 , \14484 ,
         \14485 , \14486 , \14487 , \14488 , \14489 , \14490 , \14491 , \14492 , \14493 , \14494 ,
         \14495 , \14496 , \14497 , \14498 , \14499 , \14500 , \14501 , \14502 , \14503 , \14504 ,
         \14505 , \14506 , \14507 , \14508 , \14509 , \14510 , \14511 , \14512 , \14513 , \14514 ,
         \14515 , \14516 , \14517 , \14518 , \14519 , \14520 , \14521 , \14522 , \14523 , \14524 ,
         \14525 , \14526 , \14527 , \14528 , \14529 , \14530 , \14531 , \14532 , \14533 , \14534 ,
         \14535 , \14536 , \14537 , \14538 , \14539 , \14540 , \14541 , \14542 , \14543 , \14544 ,
         \14545 , \14546 , \14547 , \14548 , \14549 , \14550 , \14551 , \14552 , \14553 , \14554 ,
         \14555 , \14556 , \14557 , \14558 , \14559 , \14560 , \14561 , \14562 , \14563 , \14564 ,
         \14565 , \14566 , \14567 , \14568 , \14569 , \14570 , \14571 , \14572 , \14573 , \14574 ,
         \14575 , \14576 , \14577 , \14578 , \14579 , \14580 , \14581 , \14582 , \14583 , \14584 ,
         \14585 , \14586 , \14587 , \14588 , \14589 , \14590 , \14591 , \14592 , \14593 , \14594 ,
         \14595 , \14596 , \14597 , \14598 , \14599 , \14600 , \14601 , \14602 , \14603 , \14604 ,
         \14605 , \14606 , \14607 , \14608 , \14609 , \14610 , \14611 , \14612 , \14613 , \14614 ,
         \14615 , \14616 , \14617 , \14618 , \14619 , \14620 , \14621 , \14622 , \14623 , \14624 ,
         \14625 , \14626 , \14627 , \14628 , \14629 , \14630 , \14631 , \14632 , \14633 , \14634 ,
         \14635 , \14636 , \14637 , \14638 , \14639 , \14640 , \14641 , \14642 , \14643 , \14644 ,
         \14645 , \14646 , \14647 , \14648 , \14649 , \14650 , \14651 , \14652 , \14653 , \14654 ,
         \14655 , \14656 , \14657 , \14658 , \14659 , \14660 , \14661 , \14662 , \14663 , \14664 ,
         \14665 , \14666 , \14667 , \14668 , \14669 , \14670 , \14671 , \14672 , \14673 , \14674 ,
         \14675 , \14676 , \14677 , \14678 , \14679 , \14680 , \14681 , \14682 , \14683 , \14684 ,
         \14685 , \14686 , \14687 , \14688 , \14689 , \14690 , \14691 , \14692 , \14693 , \14694 ,
         \14695 , \14696 , \14697 , \14698 , \14699 , \14700 , \14701 , \14702 , \14703 , \14704 ,
         \14705 , \14706 , \14707 , \14708 , \14709 , \14710 , \14711 , \14712 , \14713 , \14714 ,
         \14715 , \14716 , \14717 , \14718 , \14719 , \14720 , \14721 , \14722 , \14723 , \14724 ,
         \14725 , \14726 , \14727 , \14728 , \14729 , \14730 , \14731 , \14732 , \14733 , \14734 ,
         \14735 , \14736 , \14737 , \14738 , \14739 , \14740 , \14741 , \14742 , \14743 , \14744 ,
         \14745 , \14746 , \14747 , \14748 , \14749 , \14750 , \14751 , \14752 , \14753 , \14754 ,
         \14755 , \14756 , \14757 , \14758 , \14759 , \14760 , \14761 , \14762 , \14763 , \14764 ,
         \14765 , \14766 , \14767 , \14768 , \14769 , \14770 , \14771 , \14772 , \14773 , \14774 ,
         \14775 , \14776 , \14777 , \14778 , \14779 , \14780 , \14781 , \14782 , \14783 , \14784 ,
         \14785 , \14786 , \14787 , \14788 , \14789 , \14790 , \14791 , \14792 , \14793 , \14794 ,
         \14795 , \14796 , \14797 , \14798 , \14799 , \14800 , \14801 , \14802 , \14803 , \14804 ,
         \14805 , \14806 , \14807 , \14808 , \14809 , \14810 , \14811 , \14812 , \14813 , \14814 ,
         \14815 , \14816 , \14817 , \14818 , \14819 , \14820 , \14821 , \14822 , \14823 , \14824 ,
         \14825 , \14826 , \14827 , \14828 , \14829 , \14830 , \14831 , \14832 , \14833 , \14834 ,
         \14835 , \14836 , \14837 , \14838 , \14839 , \14840 , \14841 , \14842 , \14843 , \14844 ,
         \14845 , \14846 , \14847 , \14848 , \14849 , \14850 , \14851 , \14852 , \14853 , \14854 ,
         \14855 , \14856 , \14857 , \14858 , \14859 , \14860 , \14861 , \14862 , \14863 , \14864 ,
         \14865 , \14866 , \14867 , \14868 , \14869 , \14870 , \14871 , \14872 , \14873 , \14874 ,
         \14875 , \14876 , \14877 , \14878 , \14879 , \14880 , \14881 , \14882 , \14883 , \14884 ,
         \14885 , \14886 , \14887 , \14888 , \14889 , \14890 , \14891 , \14892 , \14893 , \14894 ,
         \14895 , \14896 , \14897 , \14898 , \14899 , \14900 , \14901 , \14902 , \14903 , \14904 ,
         \14905 , \14906 , \14907 , \14908 , \14909 , \14910 , \14911 , \14912 , \14913 , \14914 ,
         \14915 , \14916 , \14917 , \14918 , \14919 , \14920 , \14921 , \14922 , \14923 , \14924 ,
         \14925 , \14926 , \14927 , \14928 , \14929 , \14930 , \14931 , \14932 , \14933 , \14934 ,
         \14935 , \14936 , \14937 , \14938 , \14939 , \14940 , \14941 , \14942 , \14943 , \14944 ,
         \14945 , \14946 , \14947 , \14948 , \14949 , \14950 , \14951 , \14952 , \14953 , \14954 ,
         \14955 , \14956 , \14957 , \14958 , \14959 , \14960 , \14961 , \14962 , \14963 , \14964 ,
         \14965 , \14966 , \14967 , \14968 , \14969 , \14970 , \14971 , \14972 , \14973 , \14974 ,
         \14975 , \14976 , \14977 , \14978 , \14979 , \14980 , \14981 , \14982 , \14983 , \14984 ,
         \14985 , \14986 , \14987 , \14988 , \14989 , \14990 , \14991 , \14992 , \14993 , \14994 ,
         \14995 , \14996 , \14997 , \14998 , \14999 , \15000 , \15001 , \15002 , \15003 , \15004 ,
         \15005 , \15006 , \15007 , \15008 , \15009 , \15010 , \15011 , \15012 , \15013 , \15014 ,
         \15015 , \15016 , \15017 , \15018 , \15019 , \15020 , \15021 , \15022 , \15023 , \15024 ,
         \15025 , \15026 , \15027 , \15028 , \15029 , \15030 , \15031 , \15032 , \15033 , \15034 ,
         \15035 , \15036 , \15037 , \15038 , \15039 , \15040 , \15041 , \15042 , \15043 , \15044 ,
         \15045 , \15046 , \15047 , \15048 , \15049 , \15050 , \15051 , \15052 , \15053 , \15054 ,
         \15055 , \15056 , \15057 , \15058 , \15059 , \15060 , \15061 , \15062 , \15063 , \15064 ,
         \15065 , \15066 , \15067 , \15068 , \15069 , \15070 , \15071 , \15072 , \15073 , \15074 ,
         \15075 , \15076 , \15077 , \15078 , \15079 , \15080 , \15081 , \15082 , \15083 , \15084 ,
         \15085 , \15086 , \15087 , \15088 , \15089 , \15090 , \15091 , \15092 , \15093 , \15094 ,
         \15095 , \15096 , \15097 , \15098 , \15099 , \15100 , \15101 , \15102 , \15103 , \15104 ,
         \15105 , \15106 , \15107 , \15108 , \15109 , \15110 , \15111 , \15112 , \15113 , \15114 ,
         \15115 , \15116 , \15117 , \15118 , \15119 , \15120 , \15121 , \15122 , \15123 , \15124 ,
         \15125 , \15126 , \15127 , \15128 , \15129 , \15130 , \15131 , \15132 , \15133 , \15134 ,
         \15135 , \15136 , \15137 , \15138 , \15139 , \15140 , \15141 , \15142 , \15143 , \15144 ,
         \15145 , \15146 , \15147 , \15148 , \15149 , \15150 , \15151 , \15152 , \15153 , \15154 ,
         \15155 , \15156 , \15157 , \15158 , \15159 , \15160 , \15161 , \15162 , \15163 , \15164 ,
         \15165 , \15166 , \15167 , \15168 , \15169 , \15170 , \15171 , \15172 , \15173 , \15174 ,
         \15175 , \15176 , \15177 , \15178 , \15179 , \15180 , \15181 , \15182 , \15183 , \15184 ,
         \15185 , \15186 , \15187 , \15188 , \15189 , \15190 , \15191 , \15192 , \15193 , \15194 ,
         \15195 , \15196 , \15197 , \15198 , \15199 , \15200 , \15201 , \15202 , \15203 , \15204 ,
         \15205 , \15206 , \15207 , \15208 , \15209 , \15210 , \15211 , \15212 , \15213 , \15214 ,
         \15215 , \15216 , \15217 , \15218 , \15219 , \15220 , \15221 , \15222 , \15223 , \15224 ,
         \15225 , \15226 , \15227 , \15228 , \15229 , \15230 , \15231 , \15232 , \15233 , \15234 ,
         \15235 , \15236 , \15237 , \15238 , \15239 , \15240 , \15241 , \15242 , \15243 , \15244 ,
         \15245 , \15246 , \15247 , \15248 , \15249 , \15250 , \15251 , \15252 , \15253 , \15254 ,
         \15255 , \15256 , \15257 , \15258 , \15259 , \15260 , \15261 , \15262 , \15263 , \15264 ,
         \15265 , \15266 , \15267 , \15268 , \15269 , \15270 , \15271 , \15272 , \15273 , \15274 ,
         \15275 , \15276 , \15277 , \15278 , \15279 , \15280 , \15281 , \15282 , \15283 , \15284 ,
         \15285 , \15286 , \15287 , \15288 , \15289 , \15290 , \15291 , \15292 , \15293 , \15294 ,
         \15295 , \15296 , \15297 , \15298 , \15299 , \15300 , \15301 , \15302 , \15303 , \15304 ,
         \15305 , \15306 , \15307 , \15308 , \15309 , \15310 , \15311 , \15312 , \15313 , \15314 ,
         \15315 , \15316 , \15317 , \15318 , \15319 , \15320 , \15321 , \15322 , \15323 , \15324 ,
         \15325 , \15326 , \15327 , \15328 , \15329 , \15330 , \15331 , \15332 , \15333 , \15334 ,
         \15335 , \15336 , \15337 , \15338 , \15339 , \15340 , \15341 , \15342 , \15343 , \15344 ,
         \15345 , \15346 , \15347 , \15348 , \15349 , \15350 , \15351 , \15352 , \15353 , \15354 ,
         \15355 , \15356 , \15357 , \15358 , \15359 , \15360 , \15361 , \15362 , \15363 , \15364 ,
         \15365 , \15366 , \15367 , \15368 , \15369 , \15370 , \15371 , \15372 , \15373 , \15374 ,
         \15375 , \15376 , \15377 , \15378 , \15379 , \15380 , \15381 , \15382 , \15383 , \15384 ,
         \15385 , \15386 , \15387 , \15388 , \15389 , \15390 , \15391 , \15392 , \15393 , \15394 ,
         \15395 , \15396 , \15397 , \15398 , \15399 , \15400 , \15401 , \15402 , \15403 , \15404 ,
         \15405 , \15406 , \15407 , \15408 , \15409 , \15410 , \15411 , \15412 , \15413 , \15414 ,
         \15415 , \15416 , \15417 , \15418 , \15419 , \15420 , \15421 , \15422 , \15423 , \15424 ,
         \15425 , \15426 , \15427 , \15428 , \15429 , \15430 , \15431 , \15432 , \15433 , \15434 ,
         \15435 , \15436 , \15437 , \15438 , \15439 , \15440 , \15441 , \15442 , \15443 , \15444 ,
         \15445 , \15446 , \15447 , \15448 , \15449 , \15450 , \15451 , \15452 , \15453 , \15454 ,
         \15455 , \15456 , \15457 , \15458 , \15459 , \15460 , \15461 , \15462 , \15463 , \15464 ,
         \15465 , \15466 , \15467 , \15468 , \15469 , \15470 , \15471 , \15472 , \15473 , \15474 ,
         \15475 , \15476 , \15477 , \15478 , \15479 , \15480 , \15481 , \15482 , \15483 , \15484 ,
         \15485 , \15486 , \15487 , \15488 , \15489 , \15490 , \15491 , \15492 , \15493 , \15494 ,
         \15495 , \15496 , \15497 , \15498 , \15499 , \15500 , \15501 , \15502 , \15503 , \15504 ,
         \15505 , \15506 , \15507 , \15508 , \15509 , \15510 , \15511 , \15512 , \15513 , \15514 ,
         \15515 , \15516 , \15517 , \15518 , \15519 , \15520 , \15521 , \15522 , \15523 , \15524 ,
         \15525 , \15526 , \15527 , \15528 , \15529 , \15530 , \15531 , \15532 , \15533 , \15534 ,
         \15535 , \15536 , \15537 , \15538 , \15539 , \15540 , \15541 , \15542 , \15543 , \15544 ,
         \15545 , \15546 , \15547 , \15548 , \15549 , \15550 , \15551 , \15552 , \15553 , \15554 ,
         \15555 , \15556 , \15557 , \15558 , \15559 , \15560 , \15561 , \15562 , \15563 , \15564 ,
         \15565 , \15566 , \15567 , \15568 , \15569 , \15570 , \15571 , \15572 , \15573 , \15574 ,
         \15575 , \15576 , \15577 , \15578 , \15579 , \15580 , \15581 , \15582 , \15583 , \15584 ,
         \15585 , \15586 , \15587 , \15588 , \15589 , \15590 , \15591 , \15592 , \15593 , \15594 ,
         \15595 , \15596 , \15597 , \15598 , \15599 , \15600 , \15601 , \15602 , \15603 , \15604 ,
         \15605 , \15606 , \15607 , \15608 , \15609 , \15610 , \15611 , \15612 , \15613 , \15614 ,
         \15615 , \15616 , \15617 , \15618 , \15619 , \15620 , \15621 , \15622 , \15623 , \15624 ,
         \15625 , \15626 , \15627 , \15628 , \15629 , \15630 , \15631 , \15632 , \15633 , \15634 ,
         \15635 , \15636 , \15637 , \15638 , \15639 , \15640 , \15641 , \15642 , \15643 , \15644 ,
         \15645 , \15646 , \15647 , \15648 , \15649 , \15650 , \15651 , \15652 , \15653 , \15654 ,
         \15655 , \15656 , \15657 , \15658 , \15659 , \15660 , \15661 , \15662 , \15663 , \15664 ,
         \15665 , \15666 , \15667 , \15668 , \15669 , \15670 , \15671 , \15672 , \15673 , \15674 ,
         \15675 , \15676 , \15677 , \15678 , \15679 , \15680 , \15681 , \15682 , \15683 , \15684 ,
         \15685 , \15686 , \15687 , \15688 , \15689 , \15690 , \15691 , \15692 , \15693 , \15694 ,
         \15695 , \15696 , \15697 , \15698 , \15699 , \15700 , \15701 , \15702 , \15703 , \15704 ,
         \15705 , \15706 , \15707 , \15708 , \15709 , \15710 , \15711 , \15712 , \15713 , \15714 ,
         \15715 , \15716 , \15717 , \15718 , \15719 , \15720 , \15721 , \15722 , \15723 , \15724 ,
         \15725 , \15726 , \15727 , \15728 , \15729 , \15730 , \15731 , \15732 , \15733 , \15734 ,
         \15735 , \15736 , \15737 , \15738 , \15739 , \15740 , \15741 , \15742 , \15743 , \15744 ,
         \15745 , \15746 , \15747 , \15748 , \15749 , \15750 , \15751 , \15752 , \15753 , \15754 ,
         \15755 , \15756 , \15757 , \15758 , \15759 , \15760 , \15761 , \15762 , \15763 , \15764 ,
         \15765 , \15766 , \15767 , \15768 , \15769 , \15770 , \15771 , \15772 , \15773 , \15774 ,
         \15775 , \15776 , \15777 , \15778 , \15779 , \15780 , \15781 , \15782 , \15783 , \15784 ,
         \15785 , \15786 , \15787 , \15788 , \15789 , \15790 , \15791 , \15792 , \15793 , \15794 ,
         \15795 , \15796 , \15797 , \15798 , \15799 , \15800 , \15801 , \15802 , \15803 , \15804 ,
         \15805 , \15806 , \15807 , \15808 , \15809 , \15810 , \15811 , \15812 , \15813 , \15814 ,
         \15815 , \15816 , \15817 , \15818 , \15819 , \15820 , \15821 , \15822 , \15823 , \15824 ,
         \15825 , \15826 , \15827 , \15828 , \15829 , \15830 , \15831 , \15832 , \15833 , \15834 ,
         \15835 , \15836 , \15837 , \15838 , \15839 , \15840 , \15841 , \15842 , \15843 , \15844 ,
         \15845 , \15846 , \15847 , \15848 , \15849 , \15850 , \15851 , \15852 , \15853 , \15854 ,
         \15855 , \15856 , \15857 , \15858 , \15859 , \15860 , \15861 , \15862 , \15863 , \15864 ,
         \15865 , \15866 , \15867 , \15868 , \15869 , \15870 , \15871 , \15872 , \15873 , \15874 ,
         \15875 , \15876 , \15877 , \15878 , \15879 , \15880 , \15881 , \15882 , \15883 , \15884 ,
         \15885 , \15886 , \15887 , \15888 , \15889 , \15890 , \15891 , \15892 , \15893 , \15894 ,
         \15895 , \15896 , \15897 , \15898 , \15899 , \15900 , \15901 , \15902 , \15903 , \15904 ,
         \15905 , \15906 , \15907 , \15908 , \15909 , \15910 , \15911 , \15912 , \15913 , \15914 ,
         \15915 , \15916 , \15917 , \15918 , \15919 , \15920 , \15921 , \15922 , \15923 , \15924 ,
         \15925 , \15926 , \15927 , \15928 , \15929 , \15930 , \15931 , \15932 , \15933 , \15934 ,
         \15935 , \15936 , \15937 , \15938 , \15939 , \15940 , \15941 , \15942 , \15943 , \15944 ,
         \15945 , \15946 , \15947 , \15948 , \15949 , \15950 , \15951 , \15952 , \15953 , \15954 ,
         \15955 , \15956 , \15957 , \15958 , \15959 , \15960 , \15961 , \15962 , \15963 , \15964 ,
         \15965 , \15966 , \15967 , \15968 , \15969 , \15970 , \15971 , \15972 , \15973 , \15974 ,
         \15975 , \15976 , \15977 , \15978 , \15979 , \15980 , \15981 , \15982 , \15983 , \15984 ,
         \15985 , \15986 , \15987 , \15988 , \15989 , \15990 , \15991 , \15992 , \15993 , \15994 ,
         \15995 , \15996 , \15997 , \15998 , \15999 , \16000 , \16001 , \16002 , \16003 , \16004 ,
         \16005 , \16006 , \16007 , \16008 , \16009 , \16010 , \16011 , \16012 , \16013 , \16014 ,
         \16015 , \16016 , \16017 , \16018 , \16019 , \16020 , \16021 , \16022 , \16023 , \16024 ,
         \16025 , \16026 , \16027 , \16028 , \16029 , \16030 , \16031 , \16032 , \16033 , \16034 ,
         \16035 , \16036 , \16037 , \16038 , \16039 , \16040 , \16041 , \16042 , \16043 , \16044 ,
         \16045 , \16046 , \16047 , \16048 , \16049 , \16050 , \16051 , \16052 , \16053 , \16054 ,
         \16055 , \16056 , \16057 , \16058 , \16059 , \16060 , \16061 , \16062 , \16063 , \16064 ,
         \16065 , \16066 , \16067 , \16068 , \16069 , \16070 , \16071 , \16072 , \16073 , \16074 ,
         \16075 , \16076 , \16077 , \16078 , \16079 , \16080 , \16081 , \16082 , \16083 , \16084 ,
         \16085 , \16086 , \16087 , \16088 , \16089 , \16090 , \16091 , \16092 , \16093 , \16094 ,
         \16095 , \16096 , \16097 , \16098 , \16099 , \16100 , \16101 , \16102 , \16103 , \16104 ,
         \16105 , \16106 , \16107 , \16108 , \16109 , \16110 , \16111 , \16112 , \16113 , \16114 ,
         \16115 , \16116 , \16117 , \16118 , \16119 , \16120 , \16121 , \16122 , \16123 , \16124 ,
         \16125 , \16126 , \16127 , \16128 , \16129 , \16130 , \16131 , \16132 , \16133 , \16134 ,
         \16135 , \16136 , \16137 , \16138 , \16139 , \16140 , \16141 , \16142 , \16143 , \16144 ,
         \16145 , \16146 , \16147 , \16148 , \16149 , \16150 , \16151 , \16152 , \16153 , \16154 ,
         \16155 , \16156 , \16157 , \16158 , \16159 , \16160 , \16161 , \16162 , \16163 , \16164 ,
         \16165 , \16166 , \16167 , \16168 , \16169 , \16170 , \16171 , \16172 , \16173 , \16174 ,
         \16175 , \16176 , \16177 , \16178 , \16179 , \16180 , \16181 , \16182 , \16183 , \16184 ,
         \16185 , \16186 , \16187 , \16188 , \16189 , \16190 , \16191 , \16192 , \16193 , \16194 ,
         \16195 , \16196 , \16197 , \16198 , \16199 , \16200 , \16201 , \16202 , \16203 , \16204 ,
         \16205 , \16206 , \16207 , \16208 , \16209 , \16210 , \16211 , \16212 , \16213 , \16214 ,
         \16215 , \16216 , \16217 , \16218 , \16219 , \16220 , \16221 , \16222 , \16223 , \16224 ,
         \16225 , \16226 , \16227 , \16228 , \16229 , \16230 , \16231 , \16232 , \16233 , \16234 ,
         \16235 , \16236 , \16237 , \16238 , \16239 , \16240 , \16241 , \16242 , \16243 , \16244 ,
         \16245 , \16246 , \16247 , \16248 , \16249 , \16250 , \16251 , \16252 , \16253 , \16254 ,
         \16255 , \16256 , \16257 , \16258 , \16259 , \16260 , \16261 , \16262 , \16263 , \16264 ,
         \16265 , \16266 , \16267 , \16268 , \16269 , \16270 , \16271 , \16272 , \16273 , \16274 ,
         \16275 , \16276 , \16277 , \16278 , \16279 , \16280 , \16281 , \16282 , \16283 , \16284 ,
         \16285 , \16286 , \16287 , \16288 , \16289 , \16290 , \16291 , \16292 , \16293 , \16294 ,
         \16295 , \16296 , \16297 , \16298 , \16299 , \16300 , \16301 , \16302 , \16303 , \16304 ,
         \16305 , \16306 , \16307 , \16308 , \16309 , \16310 , \16311 , \16312 , \16313 , \16314 ,
         \16315 , \16316 , \16317 , \16318 , \16319 , \16320 , \16321 , \16322 , \16323 , \16324 ,
         \16325 , \16326 , \16327 , \16328 , \16329 , \16330 , \16331 , \16332 , \16333 , \16334 ,
         \16335 , \16336 , \16337 , \16338 , \16339 , \16340 , \16341 , \16342 , \16343 , \16344 ,
         \16345 , \16346 , \16347 , \16348 , \16349 , \16350 , \16351 , \16352 , \16353 , \16354 ,
         \16355 , \16356 , \16357 , \16358 , \16359 , \16360 , \16361 , \16362 , \16363 , \16364 ,
         \16365 , \16366 , \16367 , \16368 , \16369 , \16370 , \16371 , \16372 , \16373 , \16374 ,
         \16375 , \16376 , \16377 , \16378 , \16379 , \16380 , \16381 , \16382 , \16383 , \16384 ,
         \16385 , \16386 , \16387 , \16388 , \16389 , \16390 , \16391 , \16392 , \16393 , \16394 ,
         \16395 , \16396 , \16397 , \16398 , \16399 , \16400 , \16401 , \16402 , \16403 , \16404 ,
         \16405 , \16406 , \16407 , \16408 , \16409 , \16410 , \16411 , \16412 , \16413 , \16414 ,
         \16415 , \16416 , \16417 , \16418 , \16419 , \16420 , \16421 , \16422 , \16423 , \16424 ,
         \16425 , \16426 , \16427 , \16428 , \16429 , \16430 , \16431 , \16432 , \16433 , \16434 ,
         \16435 , \16436 , \16437 , \16438 , \16439 , \16440 , \16441 , \16442 , \16443 , \16444 ,
         \16445 , \16446 , \16447 , \16448 , \16449 , \16450 , \16451 , \16452 , \16453 , \16454 ,
         \16455 , \16456 , \16457 , \16458 , \16459 , \16460 , \16461 , \16462 , \16463 , \16464 ,
         \16465 , \16466 , \16467 , \16468 , \16469 , \16470 , \16471 , \16472 , \16473 , \16474 ,
         \16475 , \16476 , \16477 , \16478 , \16479 , \16480 , \16481 , \16482 , \16483 , \16484 ,
         \16485 , \16486 , \16487 , \16488 , \16489 , \16490 , \16491 , \16492 , \16493 , \16494 ,
         \16495 , \16496 , \16497 , \16498 , \16499 , \16500 , \16501 , \16502 , \16503 , \16504 ,
         \16505 , \16506 , \16507 , \16508 , \16509 , \16510 , \16511 , \16512 , \16513 , \16514 ,
         \16515 , \16516 , \16517 , \16518 , \16519 , \16520 , \16521 , \16522 , \16523 , \16524 ,
         \16525 , \16526 , \16527 , \16528 , \16529 , \16530 , \16531 , \16532 , \16533 , \16534 ,
         \16535 , \16536 , \16537 , \16538 , \16539 , \16540 , \16541 , \16542 , \16543 , \16544 ,
         \16545 , \16546 , \16547 , \16548 , \16549 , \16550 , \16551 , \16552 , \16553 , \16554 ,
         \16555 , \16556 , \16557 , \16558 , \16559 , \16560 , \16561 , \16562 , \16563 , \16564 ,
         \16565 , \16566 , \16567 , \16568 , \16569 , \16570 , \16571 , \16572 , \16573 , \16574 ,
         \16575 , \16576 , \16577 , \16578 , \16579 , \16580 , \16581 , \16582 , \16583 , \16584 ,
         \16585 , \16586 , \16587 , \16588 , \16589 , \16590 , \16591 , \16592 , \16593 , \16594 ,
         \16595 , \16596 , \16597 , \16598 , \16599 , \16600 , \16601 , \16602 , \16603 , \16604 ,
         \16605 , \16606 , \16607 , \16608 , \16609 , \16610 , \16611 , \16612 , \16613 , \16614 ,
         \16615 , \16616 , \16617 , \16618 , \16619 , \16620 , \16621 , \16622 , \16623 , \16624 ,
         \16625 , \16626 , \16627 , \16628 , \16629 , \16630 , \16631 , \16632 , \16633 , \16634 ,
         \16635 , \16636 , \16637 , \16638 , \16639 , \16640 , \16641 , \16642 , \16643 , \16644 ,
         \16645 , \16646 , \16647 , \16648 , \16649 , \16650 , \16651 , \16652 , \16653 , \16654 ,
         \16655 , \16656 , \16657 , \16658 , \16659 , \16660 , \16661 , \16662 , \16663 , \16664 ,
         \16665 , \16666 , \16667 , \16668 , \16669 , \16670 , \16671 , \16672 , \16673 , \16674 ,
         \16675 , \16676 , \16677 , \16678 , \16679 , \16680 , \16681 , \16682 , \16683 , \16684 ,
         \16685 , \16686 , \16687 , \16688 , \16689 , \16690 , \16691 , \16692 , \16693 , \16694 ,
         \16695 , \16696 , \16697 , \16698 , \16699 , \16700 , \16701 , \16702 , \16703 , \16704 ,
         \16705 , \16706 , \16707 , \16708 , \16709 , \16710 , \16711 , \16712 , \16713 , \16714 ,
         \16715 , \16716 , \16717 , \16718 , \16719 , \16720 , \16721 , \16722 , \16723 , \16724 ,
         \16725 , \16726 , \16727 , \16728 , \16729 , \16730 , \16731 , \16732 , \16733 , \16734 ,
         \16735 , \16736 , \16737 , \16738 , \16739 , \16740 , \16741 , \16742 , \16743 , \16744 ,
         \16745 , \16746 , \16747 , \16748 , \16749 , \16750 , \16751 , \16752 , \16753 , \16754 ,
         \16755 , \16756 , \16757 , \16758 , \16759 , \16760 , \16761 , \16762 , \16763 , \16764 ,
         \16765 , \16766 , \16767 , \16768 , \16769 , \16770 , \16771 , \16772 , \16773 , \16774 ,
         \16775 , \16776 , \16777 , \16778 , \16779 , \16780 , \16781 , \16782 , \16783 , \16784 ,
         \16785 , \16786 , \16787 , \16788 , \16789 , \16790 , \16791 , \16792 , \16793 , \16794 ,
         \16795 , \16796 , \16797 , \16798 , \16799 , \16800 , \16801 , \16802 , \16803 , \16804 ,
         \16805 , \16806 , \16807 , \16808 , \16809 , \16810 , \16811 , \16812 , \16813 , \16814 ,
         \16815 , \16816 , \16817 , \16818 , \16819 , \16820 , \16821 , \16822 , \16823 , \16824 ,
         \16825 , \16826 , \16827 , \16828 , \16829 , \16830 , \16831 , \16832 , \16833 , \16834 ,
         \16835 , \16836 , \16837 , \16838 , \16839 , \16840 , \16841 , \16842 , \16843 , \16844 ,
         \16845 , \16846 , \16847 , \16848 , \16849 , \16850 , \16851 , \16852 , \16853 , \16854 ,
         \16855 , \16856 , \16857 , \16858 , \16859 , \16860 , \16861 , \16862 , \16863 , \16864 ,
         \16865 , \16866 , \16867 , \16868 , \16869 , \16870 , \16871 , \16872 , \16873 , \16874 ,
         \16875 , \16876 , \16877 , \16878 , \16879 , \16880 , \16881 , \16882 , \16883 , \16884 ,
         \16885 , \16886 , \16887 , \16888 , \16889 , \16890 , \16891 , \16892 , \16893 , \16894 ,
         \16895 , \16896 , \16897 , \16898 , \16899 , \16900 , \16901 , \16902 , \16903 , \16904 ,
         \16905 , \16906 , \16907 , \16908 , \16909 , \16910 , \16911 , \16912 , \16913 , \16914 ,
         \16915 , \16916 , \16917 , \16918 , \16919 , \16920 , \16921 , \16922 , \16923 , \16924 ,
         \16925 , \16926 , \16927 , \16928 , \16929 , \16930 , \16931 , \16932 , \16933 , \16934 ,
         \16935 , \16936 , \16937 , \16938 , \16939 , \16940 , \16941 , \16942 , \16943 , \16944 ,
         \16945 , \16946 , \16947 , \16948 , \16949 , \16950 , \16951 , \16952 , \16953 , \16954 ,
         \16955 , \16956 , \16957 , \16958 , \16959 , \16960 , \16961 , \16962 , \16963 , \16964 ,
         \16965 , \16966 , \16967 , \16968 , \16969 , \16970 , \16971 , \16972 , \16973 , \16974 ,
         \16975 , \16976 , \16977 , \16978 , \16979 , \16980 , \16981 , \16982 , \16983 , \16984 ,
         \16985 , \16986 , \16987 , \16988 , \16989 , \16990 , \16991 , \16992 , \16993 , \16994 ,
         \16995 , \16996 , \16997 , \16998 , \16999 , \17000 , \17001 , \17002 , \17003 , \17004 ,
         \17005 , \17006 , \17007 , \17008 , \17009 , \17010 , \17011 , \17012 , \17013 , \17014 ,
         \17015 , \17016 , \17017 , \17018 , \17019 , \17020 , \17021 , \17022 , \17023 , \17024 ,
         \17025 , \17026 , \17027 , \17028 , \17029 , \17030 , \17031 , \17032 , \17033 , \17034 ,
         \17035 , \17036 , \17037 , \17038 , \17039 , \17040 , \17041 , \17042 , \17043 , \17044 ,
         \17045 , \17046 , \17047 , \17048 , \17049 , \17050 , \17051 , \17052 , \17053 , \17054 ,
         \17055 , \17056 , \17057 , \17058 , \17059 , \17060 , \17061 , \17062 , \17063 , \17064 ,
         \17065 , \17066 , \17067 , \17068 , \17069 , \17070 , \17071 , \17072 , \17073 , \17074 ,
         \17075 , \17076 , \17077 , \17078 , \17079 , \17080 , \17081 , \17082 , \17083 , \17084 ,
         \17085 , \17086 , \17087 , \17088 , \17089 , \17090 , \17091 , \17092 , \17093 , \17094 ,
         \17095 , \17096 , \17097 , \17098 , \17099 , \17100 , \17101 , \17102 , \17103 , \17104 ,
         \17105 , \17106 , \17107 , \17108 , \17109 , \17110 , \17111 , \17112 , \17113 , \17114 ,
         \17115 , \17116 , \17117 , \17118 , \17119 , \17120 , \17121 , \17122 , \17123 , \17124 ,
         \17125 , \17126 , \17127 , \17128 , \17129 , \17130 , \17131 , \17132 , \17133 , \17134 ,
         \17135 , \17136 , \17137 , \17138 , \17139 , \17140 , \17141 , \17142 , \17143 , \17144 ,
         \17145 , \17146 , \17147 , \17148 , \17149 , \17150 , \17151 , \17152 , \17153 , \17154 ,
         \17155 , \17156 , \17157 , \17158 , \17159 , \17160 , \17161 , \17162 , \17163 , \17164 ,
         \17165 , \17166 , \17167 , \17168 , \17169 , \17170 , \17171 , \17172 , \17173 , \17174 ,
         \17175 , \17176 , \17177 , \17178 , \17179 , \17180 , \17181 , \17182 , \17183 , \17184 ,
         \17185 , \17186 , \17187 , \17188 , \17189 , \17190 , \17191 , \17192 , \17193 , \17194 ,
         \17195 , \17196 , \17197 , \17198 , \17199 , \17200 , \17201 , \17202 , \17203 , \17204 ,
         \17205 , \17206 , \17207 , \17208 , \17209 , \17210 , \17211 , \17212 , \17213 , \17214 ,
         \17215 , \17216 , \17217 , \17218 , \17219 , \17220 , \17221 , \17222 , \17223 , \17224 ,
         \17225 , \17226 , \17227 , \17228 , \17229 , \17230 , \17231 , \17232 , \17233 , \17234 ,
         \17235 , \17236 , \17237 , \17238 , \17239 , \17240 , \17241 , \17242 , \17243 , \17244 ,
         \17245 , \17246 , \17247 , \17248 , \17249 , \17250 , \17251 , \17252 , \17253 , \17254 ,
         \17255 , \17256 , \17257 , \17258 , \17259 , \17260 , \17261 , \17262 , \17263 , \17264 ,
         \17265 , \17266 , \17267 , \17268 , \17269 , \17270 , \17271 , \17272 , \17273 , \17274 ,
         \17275 , \17276 , \17277 , \17278 , \17279 , \17280 , \17281 , \17282 , \17283 , \17284 ,
         \17285 , \17286 , \17287 , \17288 , \17289 , \17290 , \17291 , \17292 , \17293 , \17294 ,
         \17295 , \17296 , \17297 , \17298 , \17299 , \17300 , \17301 , \17302 , \17303 , \17304 ,
         \17305 , \17306 , \17307 , \17308 , \17309 , \17310 , \17311 , \17312 , \17313 , \17314 ,
         \17315 , \17316 , \17317 , \17318 , \17319 , \17320 , \17321 , \17322 , \17323 , \17324 ,
         \17325 , \17326 , \17327 , \17328 , \17329 , \17330 , \17331 , \17332 , \17333 , \17334 ,
         \17335 , \17336 , \17337 , \17338 , \17339 , \17340 , \17341 , \17342 , \17343 , \17344 ,
         \17345 , \17346 , \17347 , \17348 , \17349 , \17350 , \17351 , \17352 , \17353 , \17354 ,
         \17355 , \17356 , \17357 , \17358 , \17359 , \17360 , \17361 , \17362 , \17363 , \17364 ,
         \17365 , \17366 , \17367 , \17368 , \17369 , \17370 , \17371 , \17372 , \17373 , \17374 ,
         \17375 , \17376 , \17377 , \17378 , \17379 , \17380 , \17381 , \17382 , \17383 , \17384 ,
         \17385 , \17386 , \17387 , \17388 , \17389 , \17390 , \17391 , \17392 , \17393 , \17394 ,
         \17395 , \17396 , \17397 , \17398 , \17399 , \17400 , \17401 , \17402 , \17403 , \17404 ,
         \17405 , \17406 , \17407 , \17408 , \17409 , \17410 , \17411 , \17412 , \17413 , \17414 ,
         \17415 , \17416 , \17417 , \17418 , \17419 , \17420 , \17421 , \17422 , \17423 , \17424 ,
         \17425 , \17426 , \17427 , \17428 , \17429 , \17430 , \17431 , \17432 , \17433 , \17434 ,
         \17435 , \17436 , \17437 , \17438 , \17439 , \17440 , \17441 , \17442 , \17443 , \17444 ,
         \17445 , \17446 , \17447 , \17448 , \17449 , \17450 , \17451 , \17452 , \17453 , \17454 ,
         \17455 , \17456 , \17457 , \17458 , \17459 , \17460 , \17461 , \17462 , \17463 , \17464 ,
         \17465 , \17466 , \17467 , \17468 , \17469 , \17470 , \17471 , \17472 , \17473 , \17474 ,
         \17475 , \17476 , \17477 , \17478 , \17479 , \17480 , \17481 , \17482 , \17483 , \17484 ,
         \17485 , \17486 , \17487 , \17488 , \17489 , \17490 , \17491 , \17492 , \17493 , \17494 ,
         \17495 , \17496 , \17497 , \17498 , \17499 , \17500 , \17501 , \17502 , \17503 , \17504 ,
         \17505 , \17506 , \17507 , \17508 , \17509 , \17510 , \17511 , \17512 , \17513 , \17514 ,
         \17515 , \17516 , \17517 , \17518 , \17519 , \17520 , \17521 , \17522 , \17523 , \17524 ,
         \17525 , \17526 , \17527 , \17528 , \17529 , \17530 , \17531 , \17532 , \17533 , \17534 ,
         \17535 , \17536 , \17537 , \17538 , \17539 , \17540 , \17541 , \17542 , \17543 , \17544 ,
         \17545 , \17546 , \17547 , \17548 , \17549 , \17550 , \17551 , \17552 , \17553 , \17554 ,
         \17555 , \17556 , \17557 , \17558 , \17559 , \17560 , \17561 , \17562 , \17563 , \17564 ,
         \17565 , \17566 , \17567 , \17568 , \17569 , \17570 , \17571 , \17572 , \17573 , \17574 ,
         \17575 , \17576 , \17577 , \17578 , \17579 , \17580 , \17581 , \17582 , \17583 , \17584 ,
         \17585 , \17586 , \17587 , \17588 , \17589 , \17590 , \17591 , \17592 , \17593 , \17594 ,
         \17595 , \17596 , \17597 , \17598 , \17599 , \17600 , \17601 , \17602 , \17603 , \17604 ,
         \17605 , \17606 , \17607 , \17608 , \17609 , \17610 , \17611 , \17612 , \17613 , \17614 ,
         \17615 , \17616 , \17617 , \17618 , \17619 , \17620 , \17621 , \17622 , \17623 , \17624 ,
         \17625 , \17626 , \17627 , \17628 , \17629 , \17630 , \17631 , \17632 , \17633 , \17634 ,
         \17635 , \17636 , \17637 , \17638 , \17639 , \17640 , \17641 , \17642 , \17643 , \17644 ,
         \17645 , \17646 , \17647 , \17648 , \17649 , \17650 , \17651 , \17652 , \17653 , \17654 ,
         \17655 , \17656 , \17657 , \17658 , \17659 , \17660 , \17661 , \17662 , \17663 , \17664 ,
         \17665 , \17666 , \17667 , \17668 , \17669 , \17670 , \17671 , \17672 , \17673 , \17674 ,
         \17675 , \17676 , \17677 , \17678 , \17679 , \17680 , \17681 , \17682 , \17683 , \17684 ,
         \17685 , \17686 , \17687 , \17688 , \17689 , \17690 , \17691 , \17692 , \17693 , \17694 ,
         \17695 , \17696 , \17697 , \17698 , \17699 , \17700 , \17701 , \17702 , \17703 , \17704 ,
         \17705 , \17706 , \17707 , \17708 , \17709 , \17710 , \17711 , \17712 , \17713 , \17714 ,
         \17715 , \17716 , \17717 , \17718 , \17719 , \17720 , \17721 , \17722 , \17723 , \17724 ,
         \17725 , \17726 , \17727 , \17728 , \17729 , \17730 , \17731 , \17732 , \17733 , \17734 ,
         \17735 , \17736 , \17737 , \17738 , \17739 , \17740 , \17741 , \17742 , \17743 , \17744 ,
         \17745 , \17746 , \17747 , \17748 , \17749 , \17750 , \17751 , \17752 , \17753 , \17754 ,
         \17755 , \17756 , \17757 , \17758 , \17759 , \17760 , \17761 , \17762 , \17763 , \17764 ,
         \17765 , \17766 , \17767 , \17768 , \17769 , \17770 , \17771 , \17772 , \17773 , \17774 ,
         \17775 , \17776 , \17777 , \17778 , \17779 , \17780 , \17781 , \17782 , \17783 , \17784 ,
         \17785 , \17786 , \17787 , \17788 , \17789 , \17790 , \17791 , \17792 , \17793 , \17794 ,
         \17795 , \17796 , \17797 , \17798 , \17799 , \17800 , \17801 , \17802 , \17803 , \17804 ,
         \17805 , \17806 , \17807 , \17808 , \17809 , \17810 , \17811 , \17812 , \17813 , \17814 ,
         \17815 , \17816 , \17817 , \17818 , \17819 , \17820 , \17821 , \17822 , \17823 , \17824 ,
         \17825 , \17826 , \17827 , \17828 , \17829 , \17830 , \17831 , \17832 , \17833 , \17834 ,
         \17835 , \17836 , \17837 , \17838 , \17839 , \17840 , \17841 , \17842 , \17843 , \17844 ,
         \17845 , \17846 , \17847 , \17848 , \17849 , \17850 , \17851 , \17852 , \17853 , \17854 ,
         \17855 , \17856 , \17857 , \17858 , \17859 , \17860 , \17861 , \17862 , \17863 , \17864 ,
         \17865 , \17866 , \17867 , \17868 , \17869 , \17870 , \17871 , \17872 , \17873 , \17874 ,
         \17875 , \17876 , \17877 , \17878 , \17879 , \17880 , \17881 , \17882 , \17883 , \17884 ,
         \17885 , \17886 , \17887 , \17888 , \17889 , \17890 , \17891 , \17892 , \17893 , \17894 ,
         \17895 , \17896 , \17897 , \17898 , \17899 , \17900 , \17901 , \17902 , \17903 , \17904 ,
         \17905 , \17906 , \17907 , \17908 , \17909 , \17910 , \17911 , \17912 , \17913 , \17914 ,
         \17915 , \17916 , \17917 , \17918 , \17919 , \17920 , \17921 , \17922 , \17923 , \17924 ,
         \17925 , \17926 , \17927 , \17928 , \17929 , \17930 , \17931 , \17932 , \17933 , \17934 ,
         \17935 , \17936 , \17937 , \17938 , \17939 , \17940 , \17941 , \17942 , \17943 , \17944 ,
         \17945 , \17946 , \17947 , \17948 , \17949 , \17950 , \17951 , \17952 , \17953 , \17954 ,
         \17955 , \17956 , \17957 , \17958 , \17959 , \17960 , \17961 , \17962 , \17963 , \17964 ,
         \17965 , \17966 , \17967 , \17968 , \17969 , \17970 , \17971 , \17972 , \17973 , \17974 ,
         \17975 , \17976 , \17977 , \17978 , \17979 , \17980 , \17981 , \17982 , \17983 , \17984 ,
         \17985 , \17986 , \17987 , \17988 , \17989 , \17990 , \17991 , \17992 , \17993 , \17994 ,
         \17995 , \17996 , \17997 , \17998 , \17999 , \18000 , \18001 , \18002 , \18003 , \18004 ,
         \18005 , \18006 , \18007 , \18008 , \18009 , \18010 , \18011 , \18012 , \18013 , \18014 ,
         \18015 , \18016 , \18017 , \18018 , \18019 , \18020 , \18021 , \18022 , \18023 , \18024 ,
         \18025 , \18026 , \18027 , \18028 , \18029 , \18030 , \18031 , \18032 , \18033 , \18034 ,
         \18035 , \18036 , \18037 , \18038 , \18039 , \18040 , \18041 , \18042 , \18043 , \18044 ,
         \18045 , \18046 , \18047 , \18048 , \18049 , \18050 , \18051 , \18052 , \18053 , \18054 ,
         \18055 , \18056 , \18057 , \18058 , \18059 , \18060 , \18061 , \18062 , \18063 , \18064 ,
         \18065 , \18066 , \18067 , \18068 , \18069 , \18070 , \18071 , \18072 , \18073 , \18074 ,
         \18075 , \18076 , \18077 , \18078 , \18079 , \18080 , \18081 , \18082 , \18083 , \18084 ,
         \18085 , \18086 , \18087 , \18088 , \18089 , \18090 , \18091 , \18092 , \18093 , \18094 ,
         \18095 , \18096 , \18097 , \18098 , \18099 , \18100 , \18101 , \18102 , \18103 , \18104 ,
         \18105 , \18106 , \18107 , \18108 , \18109 , \18110 , \18111 , \18112 , \18113 , \18114 ,
         \18115 , \18116 , \18117 , \18118 , \18119 , \18120 , \18121 , \18122 , \18123 , \18124 ,
         \18125 , \18126 , \18127 , \18128 , \18129 , \18130 , \18131 , \18132 , \18133 , \18134 ,
         \18135 , \18136 , \18137 , \18138 , \18139 , \18140 , \18141 , \18142 , \18143 , \18144 ,
         \18145 , \18146 , \18147 , \18148 , \18149 , \18150 , \18151 , \18152 , \18153 , \18154 ,
         \18155 , \18156 , \18157 , \18158 , \18159 , \18160 , \18161 , \18162 , \18163 , \18164 ,
         \18165 , \18166 , \18167 , \18168 , \18169 , \18170 , \18171 , \18172 , \18173 , \18174 ,
         \18175 , \18176 , \18177 , \18178 , \18179 , \18180 , \18181 , \18182 , \18183 , \18184 ,
         \18185 , \18186 , \18187 , \18188 , \18189 , \18190 , \18191 , \18192 , \18193 , \18194 ,
         \18195 , \18196 , \18197 , \18198 , \18199 , \18200 , \18201 , \18202 , \18203 , \18204 ,
         \18205 , \18206 , \18207 , \18208 , \18209 , \18210 , \18211 , \18212 , \18213 , \18214 ,
         \18215 , \18216 , \18217 , \18218 , \18219 , \18220 , \18221 , \18222 , \18223 , \18224 ,
         \18225 , \18226 , \18227 , \18228 , \18229 , \18230 , \18231 , \18232 , \18233 , \18234 ,
         \18235 , \18236 , \18237 , \18238 , \18239 , \18240 , \18241 , \18242 , \18243 , \18244 ,
         \18245 , \18246 , \18247 , \18248 , \18249 , \18250 , \18251 , \18252 , \18253 , \18254 ,
         \18255 , \18256 , \18257 , \18258 , \18259 , \18260 , \18261 , \18262 , \18263 , \18264 ,
         \18265 , \18266 , \18267 , \18268 , \18269 , \18270 , \18271 , \18272 , \18273 , \18274 ,
         \18275 , \18276 , \18277 , \18278 , \18279 , \18280 , \18281 , \18282 , \18283 , \18284 ,
         \18285 , \18286 , \18287 , \18288 , \18289 , \18290 , \18291 , \18292 , \18293 , \18294 ,
         \18295 , \18296 , \18297 , \18298 , \18299 , \18300 , \18301 , \18302 , \18303 , \18304 ,
         \18305 , \18306 , \18307 , \18308 , \18309 , \18310 , \18311 , \18312 , \18313 , \18314 ,
         \18315 , \18316 , \18317 , \18318 , \18319 , \18320 , \18321 , \18322 , \18323 , \18324 ,
         \18325 , \18326 , \18327 , \18328 , \18329 , \18330 , \18331 , \18332 , \18333 , \18334 ,
         \18335 , \18336 , \18337 , \18338 , \18339 , \18340 , \18341 , \18342 , \18343 , \18344 ,
         \18345 , \18346 , \18347 , \18348 , \18349 , \18350 , \18351 , \18352 , \18353 , \18354 ,
         \18355 , \18356 , \18357 , \18358 , \18359 , \18360 , \18361 , \18362 , \18363 , \18364 ,
         \18365 , \18366 , \18367 , \18368 , \18369 , \18370 , \18371 , \18372 , \18373 , \18374 ,
         \18375 , \18376 , \18377 , \18378 , \18379 , \18380 , \18381 , \18382 , \18383 , \18384 ,
         \18385 , \18386 , \18387 , \18388 , \18389 , \18390 , \18391 , \18392 , \18393 , \18394 ,
         \18395 , \18396 , \18397 , \18398 , \18399 , \18400 , \18401 , \18402 , \18403 , \18404 ,
         \18405 , \18406 , \18407 , \18408 , \18409 , \18410 , \18411 , \18412 , \18413 , \18414 ,
         \18415 , \18416 , \18417 , \18418 , \18419 , \18420 , \18421 , \18422 , \18423 , \18424 ,
         \18425 , \18426 , \18427 , \18428 , \18429 , \18430 , \18431 , \18432 , \18433 , \18434 ,
         \18435 , \18436 , \18437 , \18438 , \18439 , \18440 , \18441 , \18442 , \18443 , \18444 ,
         \18445 , \18446 , \18447 , \18448 , \18449 , \18450 , \18451 , \18452 , \18453 , \18454 ,
         \18455 , \18456 , \18457 , \18458 , \18459 , \18460 , \18461 , \18462 , \18463 , \18464 ,
         \18465 , \18466 , \18467 , \18468 , \18469 , \18470 , \18471 , \18472 , \18473 , \18474 ,
         \18475 , \18476 , \18477 , \18478 , \18479 , \18480 , \18481 , \18482 , \18483 , \18484 ,
         \18485 , \18486 , \18487 , \18488 , \18489 , \18490 , \18491 , \18492 , \18493 , \18494 ,
         \18495 , \18496 , \18497 , \18498 , \18499 , \18500 , \18501 , \18502 , \18503 , \18504 ,
         \18505 , \18506 , \18507 , \18508 , \18509 , \18510 , \18511 , \18512 , \18513 , \18514 ,
         \18515 , \18516 , \18517 , \18518 , \18519 , \18520 , \18521 , \18522 , \18523 , \18524 ,
         \18525 , \18526 , \18527 , \18528 , \18529 , \18530 , \18531 , \18532 , \18533 , \18534 ,
         \18535 , \18536 , \18537 , \18538 , \18539 , \18540 , \18541 , \18542 , \18543 , \18544 ,
         \18545 , \18546 , \18547 , \18548 , \18549 , \18550 , \18551 , \18552 , \18553 , \18554 ,
         \18555 , \18556 , \18557 , \18558 , \18559 , \18560 , \18561 , \18562 , \18563 , \18564 ,
         \18565 , \18566 , \18567 , \18568 , \18569 , \18570 , \18571 , \18572 , \18573 , \18574 ,
         \18575 , \18576 , \18577 , \18578 , \18579 , \18580 , \18581 , \18582 , \18583 , \18584 ,
         \18585 , \18586 , \18587 , \18588 , \18589 , \18590 , \18591 , \18592 , \18593 , \18594 ,
         \18595 , \18596 , \18597 , \18598 , \18599 , \18600 , \18601 , \18602 , \18603 , \18604 ,
         \18605 , \18606 , \18607 , \18608 , \18609 , \18610 , \18611 , \18612 , \18613 , \18614 ,
         \18615 , \18616 , \18617 , \18618 , \18619 , \18620 , \18621 , \18622 , \18623 , \18624 ,
         \18625 , \18626 , \18627 , \18628 , \18629 , \18630 , \18631 , \18632 , \18633 , \18634 ,
         \18635 , \18636 , \18637 , \18638 , \18639 , \18640 , \18641 , \18642 , \18643 , \18644 ,
         \18645 , \18646 , \18647 , \18648 , \18649 , \18650 , \18651 , \18652 , \18653 , \18654 ,
         \18655 , \18656 , \18657 , \18658 , \18659 , \18660 , \18661 , \18662 , \18663 , \18664 ,
         \18665 , \18666 , \18667 , \18668 , \18669 , \18670 , \18671 , \18672 , \18673 , \18674 ,
         \18675 , \18676 , \18677 , \18678 , \18679 , \18680 , \18681 , \18682 , \18683 , \18684 ,
         \18685 , \18686 , \18687 , \18688 , \18689 , \18690 , \18691 , \18692 , \18693 , \18694 ,
         \18695 , \18696 , \18697 , \18698 , \18699 , \18700 , \18701 , \18702 , \18703 , \18704 ,
         \18705 , \18706 , \18707 , \18708 , \18709 , \18710 , \18711 , \18712 , \18713 , \18714 ,
         \18715 , \18716 , \18717 , \18718 , \18719 , \18720 , \18721 , \18722 , \18723 , \18724 ,
         \18725 , \18726 , \18727 , \18728 , \18729 , \18730 , \18731 , \18732 , \18733 , \18734 ,
         \18735 , \18736 , \18737 , \18738 , \18739 , \18740 , \18741 , \18742 , \18743 , \18744 ,
         \18745 , \18746 , \18747 , \18748 , \18749 , \18750 , \18751 , \18752 , \18753 , \18754 ,
         \18755 , \18756 , \18757 , \18758 , \18759 , \18760 , \18761 , \18762 , \18763 , \18764 ,
         \18765 , \18766 , \18767 , \18768 , \18769 , \18770 , \18771 , \18772 , \18773 , \18774 ,
         \18775 , \18776 , \18777 , \18778 , \18779 , \18780 , \18781 , \18782 , \18783 , \18784 ,
         \18785 , \18786 , \18787 , \18788 , \18789 , \18790 , \18791 , \18792 , \18793 , \18794 ,
         \18795 , \18796 , \18797 , \18798 , \18799 , \18800 , \18801 , \18802 , \18803 , \18804 ,
         \18805 , \18806 , \18807 , \18808 , \18809 , \18810 , \18811 , \18812 , \18813 , \18814 ,
         \18815 , \18816 , \18817 , \18818 , \18819 , \18820 , \18821 , \18822 , \18823 , \18824 ,
         \18825 , \18826 , \18827 , \18828 , \18829 , \18830 , \18831 , \18832 , \18833 , \18834 ,
         \18835 , \18836 , \18837 , \18838 , \18839 , \18840 , \18841 , \18842 , \18843 , \18844 ,
         \18845 , \18846 , \18847 , \18848 , \18849 , \18850 , \18851 , \18852 , \18853 , \18854 ,
         \18855 , \18856 , \18857 , \18858 , \18859 , \18860 , \18861 , \18862 , \18863 , \18864 ,
         \18865 , \18866 , \18867 , \18868 , \18869 , \18870 , \18871 , \18872 , \18873 , \18874 ,
         \18875 , \18876 , \18877 , \18878 , \18879 , \18880 , \18881 , \18882 , \18883 , \18884 ,
         \18885 , \18886 , \18887 , \18888 , \18889 , \18890 , \18891 , \18892 , \18893 , \18894 ,
         \18895 , \18896 , \18897 , \18898 , \18899 , \18900 , \18901 , \18902 , \18903 , \18904 ,
         \18905 , \18906 , \18907 , \18908 , \18909 , \18910 , \18911 , \18912 , \18913 , \18914 ,
         \18915 , \18916 , \18917 , \18918 , \18919 , \18920 , \18921 , \18922 , \18923 , \18924 ,
         \18925 , \18926 , \18927 , \18928 , \18929 , \18930 , \18931 , \18932 , \18933 , \18934 ,
         \18935 , \18936 , \18937 , \18938 , \18939 , \18940 , \18941 , \18942 , \18943 , \18944 ,
         \18945 , \18946 , \18947 , \18948 , \18949 , \18950 , \18951 , \18952 , \18953 , \18954 ,
         \18955 , \18956 , \18957 , \18958 , \18959 , \18960 , \18961 , \18962 , \18963 , \18964 ,
         \18965 , \18966 , \18967 , \18968 , \18969 , \18970 , \18971 , \18972 , \18973 , \18974 ,
         \18975 , \18976 , \18977 , \18978 , \18979 , \18980 , \18981 , \18982 , \18983 , \18984 ,
         \18985 , \18986 , \18987 , \18988 , \18989 , \18990 , \18991 , \18992 , \18993 , \18994 ,
         \18995 , \18996 , \18997 , \18998 , \18999 , \19000 , \19001 , \19002 , \19003 , \19004 ,
         \19005 , \19006 , \19007 , \19008 , \19009 , \19010 , \19011 , \19012 , \19013 , \19014 ,
         \19015 , \19016 , \19017 , \19018 , \19019 , \19020 , \19021 , \19022 , \19023 , \19024 ,
         \19025 , \19026 , \19027 , \19028 , \19029 , \19030 , \19031 , \19032 , \19033 , \19034 ,
         \19035 , \19036 , \19037 , \19038 , \19039 , \19040 , \19041 , \19042 , \19043 , \19044 ,
         \19045 , \19046 , \19047 , \19048 , \19049 , \19050 , \19051 , \19052 , \19053 , \19054 ,
         \19055 , \19056 , \19057 , \19058 , \19059 , \19060 , \19061 , \19062 , \19063 , \19064 ,
         \19065 , \19066 , \19067 , \19068 , \19069 , \19070 , \19071 , \19072 , \19073 , \19074 ,
         \19075 , \19076 , \19077 , \19078 , \19079 , \19080 , \19081 , \19082 , \19083 , \19084 ,
         \19085 , \19086 , \19087 , \19088 , \19089 , \19090 , \19091 , \19092 , \19093 , \19094 ,
         \19095 , \19096 , \19097 , \19098 , \19099 , \19100 , \19101 , \19102 , \19103 , \19104 ,
         \19105 , \19106 , \19107 , \19108 , \19109 , \19110 , \19111 , \19112 , \19113 , \19114 ,
         \19115 , \19116 , \19117 , \19118 , \19119 , \19120 , \19121 , \19122 , \19123 , \19124 ,
         \19125 , \19126 , \19127 , \19128 , \19129 , \19130 , \19131 , \19132 , \19133 , \19134 ,
         \19135 , \19136 , \19137 , \19138 , \19139 , \19140 , \19141 , \19142 , \19143 , \19144 ,
         \19145 , \19146 , \19147 , \19148 , \19149 , \19150 , \19151 , \19152 , \19153 , \19154 ,
         \19155 , \19156 , \19157 , \19158 , \19159 , \19160 , \19161 , \19162 , \19163 , \19164 ,
         \19165 , \19166 , \19167 , \19168 , \19169 , \19170 , \19171 , \19172 , \19173 , \19174 ,
         \19175 , \19176 , \19177 , \19178 , \19179 , \19180 , \19181 , \19182 , \19183 , \19184 ,
         \19185 , \19186 , \19187 , \19188 , \19189 , \19190 , \19191 , \19192 , \19193 , \19194 ,
         \19195 , \19196 , \19197 , \19198 , \19199 , \19200 , \19201 , \19202 , \19203 , \19204 ,
         \19205 , \19206 , \19207 , \19208 , \19209 , \19210 , \19211 , \19212 , \19213 , \19214 ,
         \19215 , \19216 , \19217 , \19218 , \19219 , \19220 , \19221 , \19222 , \19223 , \19224 ,
         \19225 , \19226 , \19227 , \19228 , \19229 , \19230 , \19231 , \19232 , \19233 , \19234 ,
         \19235 , \19236 , \19237 , \19238 , \19239 , \19240 , \19241 , \19242 , \19243 , \19244 ,
         \19245 , \19246 , \19247 , \19248 , \19249 , \19250 , \19251 , \19252 , \19253 , \19254 ,
         \19255 , \19256 , \19257 , \19258 , \19259 , \19260 , \19261 , \19262 , \19263 , \19264 ,
         \19265 , \19266 , \19267 , \19268 , \19269 , \19270 , \19271 , \19272 , \19273 , \19274 ,
         \19275 , \19276 , \19277 , \19278 , \19279 , \19280 , \19281 , \19282 , \19283 , \19284 ,
         \19285 , \19286 , \19287 , \19288 , \19289 , \19290 , \19291 , \19292 , \19293 , \19294 ,
         \19295 , \19296 , \19297 , \19298 , \19299 , \19300 , \19301 , \19302 , \19303 , \19304 ,
         \19305 , \19306 , \19307 , \19308 , \19309 , \19310 , \19311 , \19312 , \19313 , \19314 ,
         \19315 , \19316 , \19317 , \19318 , \19319 , \19320 , \19321 , \19322 , \19323 , \19324 ,
         \19325 , \19326 , \19327 , \19328 , \19329 , \19330 , \19331 , \19332 , \19333 , \19334 ,
         \19335 , \19336 , \19337 , \19338 , \19339 , \19340 , \19341 , \19342 , \19343 , \19344 ,
         \19345 , \19346 , \19347 , \19348 , \19349 , \19350 , \19351 , \19352 , \19353 , \19354 ,
         \19355 , \19356 , \19357 , \19358 , \19359 , \19360 , \19361 , \19362 , \19363 , \19364 ,
         \19365 , \19366 , \19367 , \19368 , \19369 , \19370 , \19371 , \19372 , \19373 , \19374 ,
         \19375 , \19376 , \19377 , \19378 , \19379 , \19380 , \19381 , \19382 , \19383 , \19384 ,
         \19385 , \19386 , \19387 , \19388 , \19389 , \19390 , \19391 , \19392 , \19393 , \19394 ,
         \19395 , \19396 , \19397 , \19398 , \19399 , \19400 , \19401 , \19402 , \19403 , \19404 ,
         \19405 , \19406 , \19407 , \19408 , \19409 , \19410 , \19411 , \19412 , \19413 , \19414 ,
         \19415 , \19416 , \19417 , \19418 , \19419 , \19420 , \19421 , \19422 , \19423 , \19424 ,
         \19425 , \19426 , \19427 , \19428 , \19429 , \19430 , \19431 , \19432 , \19433 , \19434 ,
         \19435 , \19436 , \19437 , \19438 , \19439 , \19440 , \19441 , \19442 , \19443 , \19444 ,
         \19445 , \19446 , \19447 , \19448 , \19449 , \19450 , \19451 , \19452 , \19453 , \19454 ,
         \19455 , \19456 , \19457 , \19458 , \19459 , \19460 , \19461 , \19462 , \19463 , \19464 ,
         \19465 , \19466 , \19467 , \19468 , \19469 , \19470 , \19471 , \19472 , \19473 , \19474 ,
         \19475 , \19476 , \19477 , \19478 , \19479 , \19480 , \19481 , \19482 , \19483 , \19484 ,
         \19485 , \19486 , \19487 , \19488 , \19489 , \19490 , \19491 , \19492 , \19493 , \19494 ,
         \19495 , \19496 , \19497 , \19498 , \19499 , \19500 , \19501 , \19502 , \19503 , \19504 ,
         \19505 , \19506 , \19507 , \19508 , \19509 , \19510 , \19511 , \19512 , \19513 , \19514 ,
         \19515 , \19516 , \19517 , \19518 , \19519 , \19520 , \19521 , \19522 , \19523 , \19524 ,
         \19525 , \19526 , \19527 , \19528 , \19529 , \19530 , \19531 , \19532 , \19533 , \19534 ,
         \19535 , \19536 , \19537 , \19538 , \19539 , \19540 , \19541 , \19542 , \19543 , \19544 ,
         \19545 , \19546 , \19547 , \19548 , \19549 , \19550 , \19551 , \19552 , \19553 , \19554 ,
         \19555 , \19556 , \19557 , \19558 , \19559 , \19560 , \19561 , \19562 , \19563 , \19564 ,
         \19565 , \19566 , \19567 , \19568 , \19569 , \19570 , \19571 , \19572 , \19573 , \19574 ,
         \19575 , \19576 , \19577 , \19578 , \19579 , \19580 , \19581 , \19582 , \19583 , \19584 ,
         \19585 , \19586 , \19587 , \19588 , \19589 , \19590 , \19591 , \19592 , \19593 , \19594 ,
         \19595 , \19596 , \19597 , \19598 , \19599 , \19600 , \19601 , \19602 , \19603 , \19604 ,
         \19605 , \19606 , \19607 , \19608 , \19609 , \19610 , \19611 , \19612 , \19613 , \19614 ,
         \19615 , \19616 , \19617 , \19618 , \19619 , \19620 , \19621 , \19622 , \19623 , \19624 ,
         \19625 , \19626 , \19627 , \19628 , \19629 , \19630 , \19631 , \19632 , \19633 , \19634 ,
         \19635 , \19636 , \19637 , \19638 , \19639 , \19640 , \19641 , \19642 , \19643 , \19644 ,
         \19645 , \19646 , \19647 , \19648 , \19649 , \19650 , \19651 , \19652 , \19653 , \19654 ,
         \19655 , \19656 , \19657 , \19658 , \19659 , \19660 , \19661 , \19662 , \19663 , \19664 ,
         \19665 , \19666 , \19667 , \19668 , \19669 , \19670 , \19671 , \19672 , \19673 , \19674 ,
         \19675 , \19676 , \19677 , \19678 , \19679 , \19680 , \19681 , \19682 , \19683 , \19684 ,
         \19685 , \19686 , \19687 , \19688 , \19689 , \19690 , \19691 , \19692 , \19693 , \19694 ,
         \19695 , \19696 , \19697 , \19698 , \19699 , \19700 , \19701 , \19702 , \19703 , \19704 ,
         \19705 , \19706 , \19707 , \19708 , \19709 , \19710 , \19711 , \19712 , \19713 , \19714 ,
         \19715 , \19716 , \19717 , \19718 , \19719 , \19720 , \19721 , \19722 , \19723 , \19724 ,
         \19725 , \19726 , \19727 , \19728 , \19729 , \19730 , \19731 , \19732 , \19733 , \19734 ,
         \19735 , \19736 , \19737 , \19738 , \19739 , \19740 , \19741 , \19742 , \19743 , \19744 ,
         \19745 , \19746 , \19747 , \19748 , \19749 , \19750 , \19751 , \19752 , \19753 , \19754 ,
         \19755 , \19756 , \19757 , \19758 , \19759 , \19760 , \19761 , \19762 , \19763 , \19764 ,
         \19765 , \19766 , \19767 , \19768 , \19769 , \19770 , \19771 , \19772 , \19773 , \19774 ,
         \19775 , \19776 , \19777 , \19778 , \19779 , \19780 , \19781 , \19782 , \19783 , \19784 ,
         \19785 , \19786 , \19787 , \19788 , \19789 , \19790 , \19791 , \19792 , \19793 , \19794 ,
         \19795 , \19796 , \19797 , \19798 , \19799 , \19800 , \19801 , \19802 , \19803 , \19804 ,
         \19805 , \19806 , \19807 , \19808 , \19809 , \19810 , \19811 , \19812 , \19813 , \19814 ,
         \19815 , \19816 , \19817 , \19818 , \19819 , \19820 , \19821 , \19822 , \19823 , \19824 ,
         \19825 , \19826 , \19827 , \19828 , \19829 , \19830 , \19831 , \19832 , \19833 , \19834 ,
         \19835 , \19836 , \19837 , \19838 , \19839 , \19840 , \19841 , \19842 , \19843 , \19844 ,
         \19845 , \19846 , \19847 , \19848 , \19849 , \19850 , \19851 , \19852 , \19853 , \19854 ,
         \19855 , \19856 , \19857 , \19858 , \19859 , \19860 , \19861 , \19862 , \19863 , \19864 ,
         \19865 , \19866 , \19867 , \19868 , \19869 , \19870 , \19871 , \19872 , \19873 , \19874 ,
         \19875 , \19876 , \19877 , \19878 , \19879 , \19880 , \19881 , \19882 , \19883 , \19884 ,
         \19885 , \19886 , \19887 , \19888 , \19889 , \19890 , \19891 , \19892 , \19893 , \19894 ,
         \19895 , \19896 , \19897 , \19898 , \19899 , \19900 , \19901 , \19902 , \19903 , \19904 ,
         \19905 , \19906 , \19907 , \19908 , \19909 , \19910 , \19911 , \19912 , \19913 , \19914 ,
         \19915 , \19916 , \19917 , \19918 , \19919 , \19920 , \19921 , \19922 , \19923 , \19924 ,
         \19925 , \19926 , \19927 , \19928 , \19929 , \19930 , \19931 , \19932 , \19933 , \19934 ,
         \19935 , \19936 , \19937 , \19938 , \19939 , \19940 , \19941 , \19942 , \19943 , \19944 ,
         \19945 , \19946 , \19947 , \19948 , \19949 , \19950 , \19951 , \19952 , \19953 , \19954 ,
         \19955 , \19956 , \19957 , \19958 , \19959 , \19960 , \19961 , \19962 , \19963 , \19964 ,
         \19965 , \19966 , \19967 , \19968 , \19969 , \19970 , \19971 , \19972 , \19973 , \19974 ,
         \19975 , \19976 , \19977 , \19978 , \19979 , \19980 , \19981 , \19982 , \19983 , \19984 ,
         \19985 , \19986 , \19987 , \19988 , \19989 , \19990 , \19991 , \19992 , \19993 , \19994 ,
         \19995 , \19996 , \19997 , \19998 , \19999 , \20000 , \20001 , \20002 , \20003 , \20004 ,
         \20005 , \20006 , \20007 , \20008 , \20009 , \20010 , \20011 , \20012 , \20013 , \20014 ,
         \20015 , \20016 , \20017 , \20018 , \20019 , \20020 , \20021 , \20022 , \20023 , \20024 ,
         \20025 , \20026 , \20027 , \20028 , \20029 , \20030 , \20031 , \20032 , \20033 , \20034 ,
         \20035 , \20036 , \20037 , \20038 , \20039 , \20040 , \20041 , \20042 , \20043 , \20044 ,
         \20045 , \20046 , \20047 , \20048 , \20049 , \20050 , \20051 , \20052 , \20053 , \20054 ,
         \20055 , \20056 , \20057 , \20058 , \20059 , \20060 , \20061 , \20062 , \20063 , \20064 ,
         \20065 , \20066 , \20067 , \20068 , \20069 , \20070 , \20071 , \20072 , \20073 , \20074 ,
         \20075 , \20076 , \20077 , \20078 , \20079 , \20080 , \20081 , \20082 , \20083 , \20084 ,
         \20085 , \20086 , \20087 , \20088 , \20089 , \20090 , \20091 , \20092 , \20093 , \20094 ,
         \20095 , \20096 , \20097 , \20098 , \20099 , \20100 , \20101 , \20102 , \20103 , \20104 ,
         \20105 , \20106 , \20107 , \20108 , \20109 , \20110 , \20111 , \20112 , \20113 , \20114 ,
         \20115 , \20116 , \20117 , \20118 , \20119 , \20120 , \20121 , \20122 , \20123 , \20124 ,
         \20125 , \20126 , \20127 , \20128 , \20129 , \20130 , \20131 , \20132 , \20133 , \20134 ,
         \20135 , \20136 , \20137 , \20138 , \20139 , \20140 , \20141 , \20142 , \20143 , \20144 ,
         \20145 , \20146 , \20147 , \20148 , \20149 , \20150 , \20151 , \20152 , \20153 , \20154 ,
         \20155 , \20156 , \20157 , \20158 , \20159 , \20160 , \20161 , \20162 , \20163 , \20164 ,
         \20165 , \20166 , \20167 , \20168 , \20169 , \20170 , \20171 , \20172 , \20173 , \20174 ,
         \20175 , \20176 , \20177 , \20178 , \20179 , \20180 , \20181 , \20182 , \20183 , \20184 ,
         \20185 , \20186 , \20187 , \20188 , \20189 , \20190 , \20191 , \20192 , \20193 , \20194 ,
         \20195 , \20196 , \20197 , \20198 , \20199 , \20200 , \20201 , \20202 , \20203 , \20204 ,
         \20205 , \20206 , \20207 , \20208 , \20209 , \20210 , \20211 , \20212 , \20213 , \20214 ,
         \20215 , \20216 , \20217 , \20218 , \20219 , \20220 , \20221 , \20222 , \20223 , \20224 ,
         \20225 , \20226 , \20227 , \20228 , \20229 , \20230 , \20231 , \20232 , \20233 , \20234 ,
         \20235 , \20236 , \20237 , \20238 , \20239 , \20240 , \20241 , \20242 , \20243 , \20244 ,
         \20245 , \20246 , \20247 , \20248 , \20249 , \20250 , \20251 , \20252 , \20253 , \20254 ,
         \20255 , \20256 , \20257 , \20258 , \20259 , \20260 , \20261 , \20262 , \20263 , \20264 ,
         \20265 , \20266 , \20267 , \20268 , \20269 , \20270 , \20271 , \20272 , \20273 , \20274 ,
         \20275 , \20276 , \20277 , \20278 , \20279 , \20280 , \20281 , \20282 , \20283 , \20284 ,
         \20285 , \20286 , \20287 , \20288 , \20289 , \20290 , \20291 , \20292 , \20293 , \20294 ,
         \20295 , \20296 , \20297 , \20298 , \20299 , \20300 , \20301 , \20302 , \20303 , \20304 ,
         \20305 , \20306 , \20307 , \20308 , \20309 , \20310 , \20311 , \20312 , \20313 , \20314 ,
         \20315 , \20316 , \20317 , \20318 , \20319 , \20320 , \20321 , \20322 , \20323 , \20324 ,
         \20325 , \20326 , \20327 , \20328 , \20329 , \20330 , \20331 , \20332 , \20333 , \20334 ,
         \20335 , \20336 , \20337 , \20338 , \20339 , \20340 , \20341 , \20342 , \20343 , \20344 ,
         \20345 , \20346 , \20347 , \20348 , \20349 , \20350 , \20351 , \20352 , \20353 , \20354 ,
         \20355 , \20356 , \20357 , \20358 , \20359 , \20360 , \20361 , \20362 , \20363 , \20364 ,
         \20365 , \20366 , \20367 , \20368 , \20369 , \20370 , \20371 , \20372 , \20373 , \20374 ,
         \20375 , \20376 , \20377 , \20378 , \20379 , \20380 , \20381 , \20382 , \20383 , \20384 ,
         \20385 , \20386 , \20387 , \20388 , \20389 , \20390 , \20391 , \20392 , \20393 , \20394 ,
         \20395 , \20396 , \20397 , \20398 , \20399 , \20400 , \20401 , \20402 , \20403 , \20404 ,
         \20405 , \20406 , \20407 , \20408 , \20409 , \20410 , \20411 , \20412 , \20413 , \20414 ,
         \20415 , \20416 , \20417 , \20418 , \20419 , \20420 , \20421 , \20422 , \20423 , \20424 ,
         \20425 , \20426 , \20427 , \20428 , \20429 , \20430 , \20431 , \20432 , \20433 , \20434 ,
         \20435 , \20436 , \20437 , \20438 , \20439 , \20440 , \20441 , \20442 , \20443 , \20444 ,
         \20445 , \20446 , \20447 , \20448 , \20449 , \20450 , \20451 , \20452 , \20453 , \20454 ,
         \20455 , \20456 , \20457 , \20458 , \20459 , \20460 , \20461 , \20462 , \20463 , \20464 ,
         \20465 , \20466 , \20467 , \20468 , \20469 , \20470 , \20471 , \20472 , \20473 , \20474 ,
         \20475 , \20476 , \20477 , \20478 , \20479 , \20480 , \20481 , \20482 , \20483 , \20484 ,
         \20485 , \20486 , \20487 , \20488 , \20489 , \20490 , \20491 , \20492 , \20493 , \20494 ,
         \20495 , \20496 , \20497 , \20498 , \20499 , \20500 , \20501 , \20502 , \20503 , \20504 ,
         \20505 , \20506 , \20507 , \20508 , \20509 , \20510 , \20511 , \20512 , \20513 , \20514 ,
         \20515 , \20516 , \20517 , \20518 , \20519 , \20520 , \20521 , \20522 , \20523 , \20524 ,
         \20525 , \20526 , \20527 , \20528 , \20529 , \20530 , \20531 , \20532 , \20533 , \20534 ,
         \20535 , \20536 , \20537 , \20538 , \20539 , \20540 , \20541 , \20542 , \20543 , \20544 ,
         \20545 , \20546 , \20547 , \20548 , \20549 , \20550 , \20551 , \20552 , \20553 , \20554 ,
         \20555 , \20556 , \20557 , \20558 , \20559 , \20560 , \20561 , \20562 , \20563 , \20564 ,
         \20565 , \20566 , \20567 , \20568 , \20569 , \20570 , \20571 , \20572 , \20573 , \20574 ,
         \20575 , \20576 , \20577 , \20578 , \20579 , \20580 , \20581 , \20582 , \20583 , \20584 ,
         \20585 , \20586 , \20587 , \20588 , \20589 , \20590 , \20591 , \20592 , \20593 , \20594 ,
         \20595 , \20596 , \20597 , \20598 , \20599 , \20600 , \20601 , \20602 , \20603 , \20604 ,
         \20605 , \20606 , \20607 , \20608 , \20609 , \20610 , \20611 , \20612 , \20613 , \20614 ,
         \20615 , \20616 , \20617 , \20618 , \20619 , \20620 , \20621 , \20622 , \20623 , \20624 ,
         \20625 , \20626 , \20627 , \20628 , \20629 , \20630 , \20631 , \20632 , \20633 , \20634 ,
         \20635 , \20636 , \20637 , \20638 , \20639 , \20640 , \20641 , \20642 , \20643 , \20644 ,
         \20645 , \20646 , \20647 , \20648 , \20649 , \20650 , \20651 , \20652 , \20653 , \20654 ,
         \20655 , \20656 , \20657 , \20658 , \20659 , \20660 , \20661 , \20662 , \20663 , \20664 ,
         \20665 , \20666 , \20667 , \20668 , \20669 , \20670 , \20671 , \20672 , \20673 , \20674 ,
         \20675 , \20676 , \20677 , \20678 , \20679 , \20680 , \20681 , \20682 , \20683 , \20684 ,
         \20685 , \20686 , \20687 , \20688 , \20689 , \20690 , \20691 , \20692 , \20693 , \20694 ,
         \20695 , \20696 , \20697 , \20698 , \20699 , \20700 , \20701 , \20702 , \20703 , \20704 ,
         \20705 , \20706 , \20707 , \20708 , \20709 , \20710 , \20711 , \20712 , \20713 , \20714 ,
         \20715 , \20716 , \20717 , \20718 , \20719 , \20720 , \20721 , \20722 , \20723 , \20724 ,
         \20725 , \20726 , \20727 , \20728 , \20729 , \20730 , \20731 , \20732 , \20733 , \20734 ,
         \20735 , \20736 , \20737 , \20738 , \20739 , \20740 , \20741 , \20742 , \20743 , \20744 ,
         \20745 , \20746 , \20747 , \20748 , \20749 , \20750 , \20751 , \20752 , \20753 , \20754 ,
         \20755 , \20756 , \20757 , \20758 , \20759 , \20760 , \20761 , \20762 , \20763 , \20764 ,
         \20765 , \20766 , \20767 , \20768 , \20769 , \20770 , \20771 , \20772 , \20773 , \20774 ,
         \20775 , \20776 , \20777 , \20778 , \20779 , \20780 , \20781 , \20782 , \20783 , \20784 ,
         \20785 , \20786 , \20787 , \20788 , \20789 , \20790 , \20791 , \20792 , \20793 , \20794 ,
         \20795 , \20796 , \20797 , \20798 , \20799 , \20800 , \20801 , \20802 , \20803 , \20804 ,
         \20805 , \20806 , \20807 , \20808 , \20809 , \20810 , \20811 , \20812 , \20813 , \20814 ,
         \20815 , \20816 , \20817 , \20818 , \20819 , \20820 , \20821 , \20822 , \20823 , \20824 ,
         \20825 , \20826 , \20827 , \20828 , \20829 , \20830 , \20831 , \20832 , \20833 , \20834 ,
         \20835 , \20836 , \20837 , \20838 , \20839 , \20840 , \20841 , \20842 , \20843 , \20844 ,
         \20845 , \20846 , \20847 , \20848 , \20849 , \20850 , \20851 , \20852 , \20853 , \20854 ,
         \20855 , \20856 , \20857 , \20858 , \20859 , \20860 , \20861 , \20862 , \20863 , \20864 ,
         \20865 , \20866 , \20867 , \20868 , \20869 , \20870 , \20871 , \20872 , \20873 , \20874 ,
         \20875 , \20876 , \20877 , \20878 , \20879 , \20880 , \20881 , \20882 , \20883 , \20884 ,
         \20885 , \20886 , \20887 , \20888 , \20889 , \20890 , \20891 , \20892 , \20893 , \20894 ,
         \20895 , \20896 , \20897 , \20898 , \20899 , \20900 , \20901 , \20902 , \20903 , \20904 ,
         \20905 , \20906 , \20907 , \20908 , \20909 , \20910 , \20911 , \20912 , \20913 , \20914 ,
         \20915 , \20916 , \20917 , \20918 , \20919 , \20920 , \20921 , \20922 , \20923 , \20924 ,
         \20925 , \20926 , \20927 , \20928 , \20929 , \20930 , \20931 , \20932 , \20933 , \20934 ,
         \20935 , \20936 , \20937 , \20938 , \20939 , \20940 , \20941 , \20942 , \20943 , \20944 ,
         \20945 , \20946 , \20947 , \20948 , \20949 , \20950 , \20951 , \20952 , \20953 , \20954 ,
         \20955 , \20956 , \20957 , \20958 , \20959 , \20960 , \20961 , \20962 , \20963 , \20964 ,
         \20965 , \20966 , \20967 , \20968 , \20969 , \20970 , \20971 , \20972 , \20973 , \20974 ,
         \20975 , \20976 , \20977 , \20978 , \20979 , \20980 , \20981 , \20982 , \20983 , \20984 ,
         \20985 , \20986 , \20987 , \20988 , \20989 , \20990 , \20991 , \20992 , \20993 , \20994 ,
         \20995 , \20996 , \20997 , \20998 , \20999 , \21000 , \21001 , \21002 , \21003 , \21004 ,
         \21005 , \21006 , \21007 , \21008 , \21009 , \21010 , \21011 , \21012 , \21013 , \21014 ,
         \21015 , \21016 , \21017 , \21018 , \21019 , \21020 , \21021 , \21022 , \21023 , \21024 ,
         \21025 , \21026 , \21027 , \21028 , \21029 , \21030 , \21031 , \21032 , \21033 , \21034 ,
         \21035 , \21036 , \21037 , \21038 , \21039 , \21040 , \21041 , \21042 , \21043 , \21044 ,
         \21045 , \21046 , \21047 , \21048 , \21049 , \21050 , \21051 , \21052 , \21053 , \21054 ,
         \21055 , \21056 , \21057 , \21058 , \21059 , \21060 , \21061 , \21062 , \21063 , \21064 ,
         \21065 , \21066 , \21067 , \21068 , \21069 , \21070 , \21071 , \21072 , \21073 , \21074 ,
         \21075 , \21076 , \21077 , \21078 , \21079 , \21080 , \21081 , \21082 , \21083 , \21084 ,
         \21085 , \21086 , \21087 , \21088 , \21089 , \21090 , \21091 , \21092 , \21093 , \21094 ,
         \21095 , \21096 , \21097 , \21098 , \21099 , \21100 , \21101 , \21102 , \21103 , \21104 ,
         \21105 , \21106 , \21107 , \21108 , \21109 , \21110 , \21111 , \21112 , \21113 , \21114 ,
         \21115 , \21116 , \21117 , \21118 , \21119 , \21120 , \21121 , \21122 , \21123 , \21124 ,
         \21125 , \21126 , \21127 , \21128 , \21129 , \21130 , \21131 , \21132 , \21133 , \21134 ,
         \21135 , \21136 , \21137 , \21138 , \21139 , \21140 , \21141 , \21142 , \21143 , \21144 ,
         \21145 , \21146 , \21147 , \21148 , \21149 , \21150 , \21151 , \21152 , \21153 , \21154 ,
         \21155 , \21156 , \21157 , \21158 , \21159 , \21160 , \21161 , \21162 , \21163 , \21164 ,
         \21165 , \21166 , \21167 , \21168 , \21169 , \21170 , \21171 , \21172 , \21173 , \21174 ,
         \21175 , \21176 , \21177 , \21178 , \21179 , \21180 , \21181 , \21182 , \21183 , \21184 ,
         \21185 , \21186 , \21187 , \21188 , \21189 , \21190 , \21191 , \21192 , \21193 , \21194 ,
         \21195 , \21196 , \21197 , \21198 , \21199 , \21200 , \21201 , \21202 , \21203 , \21204 ,
         \21205 , \21206 , \21207 , \21208 , \21209 , \21210 , \21211 , \21212 , \21213 , \21214 ,
         \21215 , \21216 , \21217 , \21218 , \21219 , \21220 , \21221 , \21222 , \21223 , \21224 ,
         \21225 , \21226 , \21227 , \21228 , \21229 , \21230 , \21231 , \21232 , \21233 , \21234 ,
         \21235 , \21236 , \21237 , \21238 , \21239 , \21240 , \21241 , \21242 , \21243 , \21244 ,
         \21245 , \21246 , \21247 , \21248 , \21249 , \21250 , \21251 , \21252 , \21253 , \21254 ,
         \21255 , \21256 , \21257 , \21258 , \21259 , \21260 , \21261 , \21262 , \21263 , \21264 ,
         \21265 , \21266 , \21267 , \21268 , \21269 , \21270 , \21271 , \21272 , \21273 , \21274 ,
         \21275 , \21276 , \21277 , \21278 , \21279 , \21280 , \21281 , \21282 , \21283 , \21284 ,
         \21285 , \21286 , \21287 , \21288 , \21289 , \21290 , \21291 , \21292 , \21293 , \21294 ,
         \21295 , \21296 , \21297 , \21298 , \21299 , \21300 , \21301 , \21302 , \21303 , \21304 ,
         \21305 , \21306 , \21307 , \21308 , \21309 , \21310 , \21311 , \21312 , \21313 , \21314 ,
         \21315 , \21316 , \21317 , \21318 , \21319 , \21320 , \21321 , \21322 , \21323 , \21324 ,
         \21325 , \21326 , \21327 , \21328 , \21329 , \21330 , \21331 , \21332 , \21333 , \21334 ,
         \21335 , \21336 , \21337 , \21338 , \21339 , \21340 , \21341 , \21342 , \21343 , \21344 ,
         \21345 , \21346 , \21347 , \21348 , \21349 , \21350 , \21351 , \21352 , \21353 , \21354 ,
         \21355 , \21356 , \21357 , \21358 , \21359 , \21360 , \21361 , \21362 , \21363 , \21364 ,
         \21365 , \21366 , \21367 , \21368 , \21369 , \21370 , \21371 , \21372 , \21373 , \21374 ,
         \21375 , \21376 , \21377 , \21378 , \21379 , \21380 , \21381 , \21382 , \21383 , \21384 ,
         \21385 , \21386 , \21387 , \21388 , \21389 , \21390 , \21391 , \21392 , \21393 , \21394 ,
         \21395 , \21396 , \21397 , \21398 , \21399 , \21400 , \21401 , \21402 , \21403 , \21404 ,
         \21405 , \21406 , \21407 , \21408 , \21409 , \21410 , \21411 , \21412 , \21413 , \21414 ,
         \21415 , \21416 , \21417 , \21418 , \21419 , \21420 , \21421 , \21422 , \21423 , \21424 ,
         \21425 , \21426 , \21427 , \21428 , \21429 , \21430 , \21431 , \21432 , \21433 , \21434 ,
         \21435 , \21436 , \21437 , \21438 , \21439 , \21440 , \21441 , \21442 , \21443 , \21444 ,
         \21445 , \21446 , \21447 , \21448 , \21449 , \21450 , \21451 , \21452 , \21453 , \21454 ,
         \21455 , \21456 , \21457 , \21458 , \21459 , \21460 , \21461 , \21462 , \21463 , \21464 ,
         \21465 , \21466 , \21467 , \21468 , \21469 , \21470 , \21471 , \21472 , \21473 , \21474 ,
         \21475 , \21476 , \21477 , \21478 , \21479 , \21480 , \21481 , \21482 , \21483 , \21484 ,
         \21485 , \21486 , \21487 , \21488 , \21489 , \21490 , \21491 , \21492 , \21493 , \21494 ,
         \21495 , \21496 , \21497 , \21498 , \21499 , \21500 , \21501 , \21502 , \21503 , \21504 ,
         \21505 , \21506 , \21507 , \21508 , \21509 , \21510 , \21511 , \21512 , \21513 , \21514 ,
         \21515 , \21516 , \21517 , \21518 , \21519 , \21520 , \21521 , \21522 , \21523 , \21524 ,
         \21525 , \21526 , \21527 , \21528 , \21529 , \21530 , \21531 , \21532 , \21533 , \21534 ,
         \21535 , \21536 , \21537 , \21538 , \21539 , \21540 , \21541 , \21542 , \21543 , \21544 ,
         \21545 , \21546 , \21547 , \21548 , \21549 , \21550 , \21551 , \21552 , \21553 , \21554 ,
         \21555 , \21556 , \21557 , \21558 , \21559 , \21560 , \21561 , \21562 , \21563 , \21564 ,
         \21565 , \21566 , \21567 , \21568 , \21569 , \21570 , \21571 , \21572 , \21573 , \21574 ,
         \21575 , \21576 , \21577 , \21578 , \21579 , \21580 , \21581 , \21582 , \21583 , \21584 ,
         \21585 , \21586 , \21587 , \21588 , \21589 , \21590 , \21591 , \21592 , \21593 , \21594 ,
         \21595 , \21596 , \21597 , \21598 , \21599 , \21600 , \21601 , \21602 , \21603 , \21604 ,
         \21605 , \21606 , \21607 , \21608 , \21609 , \21610 , \21611 , \21612 , \21613 , \21614 ,
         \21615 , \21616 , \21617 , \21618 , \21619 , \21620 , \21621 , \21622 , \21623 , \21624 ,
         \21625 , \21626 , \21627 , \21628 , \21629 , \21630 , \21631 , \21632 , \21633 , \21634 ,
         \21635 , \21636 , \21637 , \21638 , \21639 , \21640 , \21641 , \21642 , \21643 , \21644 ,
         \21645 , \21646 , \21647 , \21648 , \21649 , \21650 , \21651 , \21652 , \21653 , \21654 ,
         \21655 , \21656 , \21657 , \21658 , \21659 , \21660 , \21661 , \21662 , \21663 , \21664 ,
         \21665 , \21666 , \21667 , \21668 , \21669 , \21670 , \21671 , \21672 , \21673 , \21674 ,
         \21675 , \21676 , \21677 , \21678 , \21679 , \21680 , \21681 , \21682 , \21683 , \21684 ,
         \21685 , \21686 , \21687 , \21688 , \21689 , \21690 , \21691 , \21692 , \21693 , \21694 ,
         \21695 , \21696 , \21697 , \21698 , \21699 , \21700 , \21701 , \21702 , \21703 , \21704 ,
         \21705 , \21706 , \21707 , \21708 , \21709 , \21710 , \21711 , \21712 , \21713 , \21714 ,
         \21715 , \21716 , \21717 , \21718 , \21719 , \21720 , \21721 , \21722 , \21723 , \21724 ,
         \21725 , \21726 , \21727 , \21728 , \21729 , \21730 , \21731 , \21732 , \21733 , \21734 ,
         \21735 , \21736 , \21737 , \21738 , \21739 , \21740 , \21741 , \21742 , \21743 , \21744 ,
         \21745 , \21746 , \21747 , \21748 , \21749 , \21750 , \21751 , \21752 , \21753 , \21754 ,
         \21755 , \21756 , \21757 , \21758 , \21759 , \21760 , \21761 , \21762 , \21763 , \21764 ,
         \21765 , \21766 , \21767 , \21768 , \21769 , \21770 , \21771 , \21772 , \21773 , \21774 ,
         \21775 , \21776 , \21777 , \21778 , \21779 , \21780 , \21781 , \21782 , \21783 , \21784 ,
         \21785 , \21786 , \21787 , \21788 , \21789 , \21790 , \21791 , \21792 , \21793 , \21794 ,
         \21795 , \21796 , \21797 , \21798 , \21799 , \21800 , \21801 , \21802 , \21803 , \21804 ,
         \21805 , \21806 , \21807 , \21808 , \21809 , \21810 , \21811 , \21812 , \21813 , \21814 ,
         \21815 , \21816 , \21817 , \21818 , \21819 , \21820 , \21821 , \21822 , \21823 , \21824 ,
         \21825 , \21826 , \21827 , \21828 , \21829 , \21830 , \21831 , \21832 , \21833 , \21834 ,
         \21835 , \21836 , \21837 , \21838 , \21839 , \21840 , \21841 , \21842 , \21843 , \21844 ,
         \21845 , \21846 , \21847 , \21848 , \21849 , \21850 , \21851 , \21852 , \21853 , \21854 ,
         \21855 , \21856 , \21857 , \21858 , \21859 , \21860 , \21861 , \21862 , \21863 , \21864 ,
         \21865 , \21866 , \21867 , \21868 , \21869 , \21870 , \21871 , \21872 , \21873 , \21874 ,
         \21875 , \21876 , \21877 , \21878 , \21879 , \21880 , \21881 , \21882 , \21883 , \21884 ,
         \21885 , \21886 , \21887 , \21888 , \21889 , \21890 , \21891 , \21892 , \21893 , \21894 ,
         \21895 , \21896 , \21897 , \21898 , \21899 , \21900 , \21901 , \21902 , \21903 , \21904 ,
         \21905 , \21906 , \21907 , \21908 , \21909 , \21910 , \21911 , \21912 , \21913 , \21914 ,
         \21915 , \21916 , \21917 , \21918 , \21919 , \21920 , \21921 , \21922 , \21923 , \21924 ,
         \21925 , \21926 , \21927 , \21928 , \21929 , \21930 , \21931 , \21932 , \21933 , \21934 ,
         \21935 , \21936 , \21937 , \21938 , \21939 , \21940 , \21941 , \21942 , \21943 , \21944 ,
         \21945 , \21946 , \21947 , \21948 , \21949 , \21950 , \21951 , \21952 , \21953 , \21954 ,
         \21955 , \21956 , \21957 , \21958 , \21959 , \21960 , \21961 , \21962 , \21963 , \21964 ,
         \21965 , \21966 , \21967 , \21968 , \21969 , \21970 , \21971 , \21972 , \21973 , \21974 ,
         \21975 , \21976 , \21977 , \21978 , \21979 , \21980 , \21981 , \21982 , \21983 , \21984 ,
         \21985 , \21986 , \21987 , \21988 , \21989 , \21990 , \21991 , \21992 , \21993 , \21994 ,
         \21995 , \21996 , \21997 , \21998 , \21999 , \22000 , \22001 , \22002 , \22003 , \22004 ,
         \22005 , \22006 , \22007 , \22008 , \22009 , \22010 , \22011 , \22012 , \22013 , \22014 ,
         \22015 , \22016 , \22017 , \22018 , \22019 , \22020 , \22021 , \22022 , \22023 , \22024 ,
         \22025 , \22026 , \22027 , \22028 , \22029 , \22030 , \22031 , \22032 , \22033 , \22034 ,
         \22035 , \22036 , \22037 , \22038 , \22039 , \22040 , \22041 , \22042 , \22043 , \22044 ,
         \22045 , \22046 , \22047 , \22048 , \22049 , \22050 , \22051 , \22052 , \22053 , \22054 ,
         \22055 , \22056 , \22057 , \22058 , \22059 , \22060 , \22061 , \22062 , \22063 , \22064 ,
         \22065 , \22066 , \22067 , \22068 , \22069 , \22070 , \22071 , \22072 , \22073 , \22074 ,
         \22075 , \22076 , \22077 , \22078 , \22079 , \22080 , \22081 , \22082 , \22083 , \22084 ,
         \22085 , \22086 , \22087 , \22088 , \22089 , \22090 , \22091 , \22092 , \22093 , \22094 ,
         \22095 , \22096 , \22097 , \22098 , \22099 , \22100 , \22101 , \22102 , \22103 , \22104 ,
         \22105 , \22106 , \22107 , \22108 , \22109 , \22110 , \22111 , \22112 , \22113 , \22114 ,
         \22115 , \22116 , \22117 , \22118 , \22119 , \22120 , \22121 , \22122 , \22123 , \22124 ,
         \22125 , \22126 , \22127 , \22128 , \22129 , \22130 , \22131 , \22132 , \22133 , \22134 ,
         \22135 , \22136 , \22137 , \22138 , \22139 , \22140 , \22141 , \22142 , \22143 , \22144 ,
         \22145 , \22146 , \22147 , \22148 , \22149 , \22150 , \22151 , \22152 , \22153 , \22154 ,
         \22155 , \22156 , \22157 , \22158 , \22159 , \22160 , \22161 , \22162 , \22163 , \22164 ,
         \22165 , \22166 , \22167 , \22168 , \22169 , \22170 , \22171 , \22172 , \22173 , \22174 ,
         \22175 , \22176 , \22177 , \22178 , \22179 , \22180 , \22181 , \22182 , \22183 , \22184 ,
         \22185 , \22186 , \22187 , \22188 , \22189 , \22190 , \22191 , \22192 , \22193 , \22194 ,
         \22195 , \22196 , \22197 , \22198 , \22199 , \22200 , \22201 , \22202 , \22203 , \22204 ,
         \22205 , \22206 , \22207 , \22208 , \22209 , \22210 , \22211 , \22212 , \22213 , \22214 ,
         \22215 , \22216 , \22217 , \22218 , \22219 , \22220 , \22221 , \22222 , \22223 , \22224 ,
         \22225 , \22226 , \22227 , \22228 , \22229 , \22230 , \22231 , \22232 , \22233 , \22234 ,
         \22235 , \22236 , \22237 , \22238 , \22239 , \22240 , \22241 , \22242 , \22243 , \22244 ,
         \22245 , \22246 , \22247 , \22248 , \22249 , \22250 , \22251 , \22252 , \22253 , \22254 ,
         \22255 , \22256 , \22257 , \22258 , \22259 , \22260 , \22261 , \22262 , \22263 , \22264 ,
         \22265 , \22266 , \22267 , \22268 , \22269 , \22270 , \22271 , \22272 , \22273 , \22274 ,
         \22275 , \22276 , \22277 , \22278 , \22279 , \22280 , \22281 , \22282 , \22283 , \22284 ,
         \22285 , \22286 , \22287 , \22288 , \22289 , \22290 , \22291 , \22292 , \22293 , \22294 ,
         \22295 , \22296 , \22297 , \22298 , \22299 , \22300 , \22301 , \22302 , \22303 , \22304 ,
         \22305 , \22306 , \22307 , \22308 , \22309 , \22310 , \22311 , \22312 , \22313 , \22314 ,
         \22315 , \22316 , \22317 , \22318 , \22319 , \22320 , \22321 , \22322 , \22323 , \22324 ,
         \22325 , \22326 , \22327 , \22328 , \22329 , \22330 , \22331 , \22332 , \22333 , \22334 ,
         \22335 , \22336 , \22337 , \22338 , \22339 , \22340 , \22341 , \22342 , \22343 , \22344 ,
         \22345 , \22346 , \22347 , \22348 , \22349 , \22350 , \22351 , \22352 , \22353 , \22354 ,
         \22355 , \22356 , \22357 , \22358 , \22359 , \22360 , \22361 , \22362 , \22363 , \22364 ,
         \22365 , \22366 , \22367 , \22368 , \22369 , \22370 , \22371 , \22372 , \22373 , \22374 ,
         \22375 , \22376 , \22377 , \22378 , \22379 , \22380 , \22381 , \22382 , \22383 , \22384 ,
         \22385 , \22386 , \22387 , \22388 , \22389 , \22390 , \22391 , \22392 , \22393 , \22394 ,
         \22395 , \22396 , \22397 , \22398 , \22399 , \22400 , \22401 , \22402 , \22403 , \22404 ,
         \22405 , \22406 , \22407 , \22408 , \22409 , \22410 , \22411 , \22412 , \22413 , \22414 ,
         \22415 , \22416 , \22417 , \22418 , \22419 , \22420 , \22421 , \22422 , \22423 , \22424 ,
         \22425 , \22426 , \22427 , \22428 , \22429 , \22430 , \22431 , \22432 , \22433 , \22434 ,
         \22435 , \22436 , \22437 , \22438 , \22439 , \22440 , \22441 , \22442 , \22443 , \22444 ,
         \22445 , \22446 , \22447 , \22448 , \22449 , \22450 , \22451 , \22452 , \22453 , \22454 ,
         \22455 , \22456 , \22457 , \22458 , \22459 , \22460 , \22461 , \22462 , \22463 , \22464 ,
         \22465 , \22466 , \22467 , \22468 , \22469 , \22470 , \22471 , \22472 , \22473 , \22474 ,
         \22475 , \22476 , \22477 , \22478 , \22479 , \22480 , \22481 , \22482 , \22483 , \22484 ,
         \22485 , \22486 , \22487 , \22488 , \22489 , \22490 , \22491 , \22492 , \22493 , \22494 ,
         \22495 , \22496 , \22497 , \22498 , \22499 , \22500 , \22501 , \22502 , \22503 , \22504 ,
         \22505 , \22506 , \22507 , \22508 , \22509 , \22510 , \22511 , \22512 , \22513 , \22514 ,
         \22515 , \22516 , \22517 , \22518 , \22519 , \22520 , \22521 , \22522 , \22523 , \22524 ,
         \22525 , \22526 , \22527 , \22528 , \22529 , \22530 , \22531 , \22532 , \22533 , \22534 ,
         \22535 , \22536 , \22537 , \22538 , \22539 , \22540 , \22541 , \22542 , \22543 , \22544 ,
         \22545 , \22546 , \22547 , \22548 , \22549 , \22550 , \22551 , \22552 , \22553 , \22554 ,
         \22555 , \22556 , \22557 , \22558 , \22559 , \22560 , \22561 , \22562 , \22563 , \22564 ,
         \22565 , \22566 , \22567 , \22568 , \22569 , \22570 , \22571 , \22572 , \22573 , \22574 ,
         \22575 , \22576 , \22577 , \22578 , \22579 , \22580 , \22581 , \22582 , \22583 , \22584 ,
         \22585 , \22586 , \22587 , \22588 , \22589 , \22590 , \22591 , \22592 , \22593 , \22594 ,
         \22595 , \22596 , \22597 , \22598 , \22599 , \22600 , \22601 , \22602 , \22603 , \22604 ,
         \22605 , \22606 , \22607 , \22608 , \22609 , \22610 , \22611 , \22612 , \22613 , \22614 ,
         \22615 , \22616 , \22617 , \22618 , \22619 , \22620 , \22621 , \22622 , \22623 , \22624 ,
         \22625 , \22626 , \22627 , \22628 , \22629 , \22630 , \22631 , \22632 , \22633 , \22634 ,
         \22635 , \22636 , \22637 , \22638 , \22639 , \22640 , \22641 , \22642 , \22643 , \22644 ,
         \22645 , \22646 , \22647 , \22648 , \22649 , \22650 , \22651 , \22652 , \22653 , \22654 ,
         \22655 , \22656 , \22657 , \22658 , \22659 , \22660 , \22661 , \22662 , \22663 , \22664 ,
         \22665 , \22666 , \22667 , \22668 , \22669 , \22670 , \22671 , \22672 , \22673 , \22674 ,
         \22675 , \22676 , \22677 , \22678 , \22679 , \22680 , \22681 , \22682 , \22683 , \22684 ,
         \22685 , \22686 , \22687 , \22688 , \22689 , \22690 , \22691 , \22692 , \22693 , \22694 ,
         \22695 , \22696 , \22697 , \22698 , \22699 , \22700 , \22701 , \22702 , \22703 , \22704 ,
         \22705 , \22706 , \22707 , \22708 , \22709 , \22710 , \22711 , \22712 , \22713 , \22714 ,
         \22715 , \22716 , \22717 , \22718 , \22719 , \22720 , \22721 , \22722 , \22723 , \22724 ,
         \22725 , \22726 , \22727 , \22728 , \22729 , \22730 , \22731 , \22732 , \22733 , \22734 ,
         \22735 , \22736 , \22737 , \22738 , \22739 , \22740 , \22741 , \22742 , \22743 , \22744 ,
         \22745 , \22746 , \22747 , \22748 , \22749 , \22750 , \22751 , \22752 , \22753 , \22754 ,
         \22755 , \22756 , \22757 , \22758 , \22759 , \22760 , \22761 , \22762 , \22763 , \22764 ,
         \22765 , \22766 , \22767 , \22768 , \22769 , \22770 , \22771 , \22772 , \22773 , \22774 ,
         \22775 , \22776 , \22777 , \22778 , \22779 , \22780 , \22781 , \22782 , \22783 , \22784 ,
         \22785 , \22786 , \22787 , \22788 , \22789 , \22790 , \22791 , \22792 , \22793 , \22794 ,
         \22795 , \22796 , \22797 , \22798 , \22799 , \22800 , \22801 , \22802 , \22803 , \22804 ,
         \22805 , \22806 , \22807 , \22808 , \22809 , \22810 , \22811 , \22812 , \22813 , \22814 ,
         \22815 , \22816 , \22817 , \22818 , \22819 , \22820 , \22821 , \22822 , \22823 , \22824 ,
         \22825 , \22826 , \22827 , \22828 , \22829 , \22830 , \22831 , \22832 , \22833 , \22834 ,
         \22835 , \22836 , \22837 , \22838 , \22839 , \22840 , \22841 , \22842 , \22843 , \22844 ,
         \22845 , \22846 , \22847 , \22848 , \22849 , \22850 , \22851 , \22852 , \22853 , \22854 ,
         \22855 , \22856 , \22857 , \22858 , \22859 , \22860 , \22861 , \22862 , \22863 , \22864 ,
         \22865 , \22866 , \22867 , \22868 , \22869 , \22870 , \22871 , \22872 , \22873 , \22874 ,
         \22875 , \22876 , \22877 , \22878 , \22879 , \22880 , \22881 , \22882 , \22883 , \22884 ,
         \22885 , \22886 , \22887 , \22888 , \22889 , \22890 , \22891 , \22892 , \22893 , \22894 ,
         \22895 , \22896 , \22897 , \22898 , \22899 , \22900 , \22901 , \22902 , \22903 , \22904 ,
         \22905 , \22906 , \22907 , \22908 , \22909 , \22910 , \22911 , \22912 , \22913 , \22914 ,
         \22915 , \22916 , \22917 , \22918 , \22919 , \22920 , \22921 , \22922 , \22923 , \22924 ,
         \22925 , \22926 , \22927 , \22928 , \22929 , \22930 , \22931 , \22932 , \22933 , \22934 ,
         \22935 , \22936 , \22937 , \22938 , \22939 , \22940 , \22941 , \22942 , \22943 , \22944 ,
         \22945 , \22946 , \22947 , \22948 , \22949 , \22950 , \22951 , \22952 , \22953 , \22954 ,
         \22955 , \22956 , \22957 , \22958 , \22959 , \22960 , \22961 , \22962 , \22963 , \22964 ,
         \22965 , \22966 , \22967 , \22968 , \22969 , \22970 , \22971 , \22972 , \22973 , \22974 ,
         \22975 , \22976 , \22977 , \22978 , \22979 , \22980 , \22981 , \22982 , \22983 , \22984 ,
         \22985 , \22986 , \22987 , \22988 , \22989 , \22990 , \22991 , \22992 , \22993 , \22994 ,
         \22995 , \22996 , \22997 , \22998 , \22999 , \23000 , \23001 , \23002 , \23003 , \23004 ,
         \23005 , \23006 , \23007 , \23008 , \23009 , \23010 , \23011 , \23012 , \23013 , \23014 ,
         \23015 , \23016 , \23017 , \23018 , \23019 , \23020 , \23021 , \23022 , \23023 , \23024 ,
         \23025 , \23026 , \23027 , \23028 , \23029 , \23030 , \23031 , \23032 , \23033 , \23034 ,
         \23035 , \23036 , \23037 , \23038 , \23039 , \23040 , \23041 , \23042 , \23043 , \23044 ,
         \23045 , \23046 , \23047 , \23048 , \23049 , \23050 , \23051 , \23052 , \23053 , \23054 ,
         \23055 , \23056 , \23057 , \23058 , \23059 , \23060 , \23061 , \23062 , \23063 , \23064 ,
         \23065 , \23066 , \23067 , \23068 , \23069 , \23070 , \23071 , \23072 , \23073 , \23074 ,
         \23075 , \23076 , \23077 , \23078 , \23079 , \23080 , \23081 , \23082 , \23083 , \23084 ,
         \23085 , \23086 , \23087 , \23088 , \23089 , \23090 , \23091 , \23092 , \23093 , \23094 ,
         \23095 , \23096 , \23097 , \23098 , \23099 , \23100 , \23101 , \23102 , \23103 , \23104 ,
         \23105 , \23106 , \23107 , \23108 , \23109 , \23110 , \23111 , \23112 , \23113 , \23114 ,
         \23115 , \23116 , \23117 , \23118 , \23119 , \23120 , \23121 , \23122 , \23123 , \23124 ,
         \23125 , \23126 , \23127 , \23128 , \23129 , \23130 , \23131 , \23132 , \23133 , \23134 ,
         \23135 , \23136 , \23137 , \23138 , \23139 , \23140 , \23141 , \23142 , \23143 , \23144 ,
         \23145 , \23146 , \23147 , \23148 , \23149 , \23150 , \23151 , \23152 , \23153 , \23154 ,
         \23155 , \23156 , \23157 , \23158 , \23159 , \23160 , \23161 , \23162 , \23163 , \23164 ,
         \23165 , \23166 , \23167 , \23168 , \23169 , \23170 , \23171 , \23172 , \23173 , \23174 ,
         \23175 , \23176 , \23177 , \23178 , \23179 , \23180 , \23181 , \23182 , \23183 , \23184 ,
         \23185 , \23186 , \23187 , \23188 , \23189 , \23190 , \23191 , \23192 , \23193 , \23194 ,
         \23195 , \23196 , \23197 , \23198 , \23199 , \23200 , \23201 , \23202 , \23203 , \23204 ,
         \23205 , \23206 , \23207 , \23208 , \23209 , \23210 , \23211 , \23212 , \23213 , \23214 ,
         \23215 , \23216 , \23217 , \23218 , \23219 , \23220 , \23221 , \23222 , \23223 , \23224 ,
         \23225 , \23226 , \23227 , \23228 , \23229 , \23230 , \23231 , \23232 , \23233 , \23234 ,
         \23235 , \23236 , \23237 , \23238 , \23239 , \23240 , \23241 , \23242 , \23243 , \23244 ,
         \23245 , \23246 , \23247 , \23248 , \23249 , \23250 , \23251 , \23252 , \23253 , \23254 ,
         \23255 , \23256 , \23257 , \23258 , \23259 , \23260 , \23261 , \23262 , \23263 , \23264 ,
         \23265 , \23266 , \23267 , \23268 , \23269 , \23270 , \23271 , \23272 , \23273 , \23274 ,
         \23275 , \23276 , \23277 , \23278 , \23279 , \23280 , \23281 , \23282 , \23283 , \23284 ,
         \23285 , \23286 , \23287 , \23288 , \23289 , \23290 , \23291 , \23292 , \23293 , \23294 ,
         \23295 , \23296 , \23297 , \23298 , \23299 , \23300 , \23301 , \23302 , \23303 , \23304 ,
         \23305 , \23306 , \23307 , \23308 , \23309 , \23310 , \23311 , \23312 , \23313 , \23314 ,
         \23315 , \23316 , \23317 , \23318 , \23319 , \23320 , \23321 , \23322 , \23323 , \23324 ,
         \23325 , \23326 , \23327 , \23328 , \23329 , \23330 , \23331 , \23332 , \23333 , \23334 ,
         \23335 , \23336 , \23337 , \23338 , \23339 , \23340 , \23341 , \23342 , \23343 , \23344 ,
         \23345 , \23346 , \23347 , \23348 , \23349 , \23350 , \23351 , \23352 , \23353 , \23354 ,
         \23355 , \23356 , \23357 , \23358 , \23359 , \23360 , \23361 , \23362 , \23363 , \23364 ,
         \23365 , \23366 , \23367 , \23368 , \23369 , \23370 , \23371 , \23372 , \23373 , \23374 ,
         \23375 , \23376 , \23377 , \23378 , \23379 , \23380 , \23381 , \23382 , \23383 , \23384 ,
         \23385 , \23386 , \23387 , \23388 , \23389 , \23390 , \23391 , \23392 , \23393 , \23394 ,
         \23395 , \23396 , \23397 , \23398 , \23399 , \23400 , \23401 , \23402 , \23403 , \23404 ,
         \23405 , \23406 , \23407 , \23408 , \23409 , \23410 , \23411 , \23412 , \23413 , \23414 ,
         \23415 , \23416 , \23417 , \23418 , \23419 , \23420 , \23421 , \23422 , \23423 , \23424 ,
         \23425 , \23426 , \23427 , \23428 , \23429 , \23430 , \23431 , \23432 , \23433 , \23434 ,
         \23435 , \23436 , \23437 , \23438 , \23439 , \23440 , \23441 , \23442 , \23443 , \23444 ,
         \23445 , \23446 , \23447 , \23448 , \23449 , \23450 , \23451 , \23452 , \23453 , \23454 ,
         \23455 , \23456 , \23457 , \23458 , \23459 , \23460 , \23461 , \23462 , \23463 , \23464 ,
         \23465 , \23466 , \23467 , \23468 , \23469 , \23470 , \23471 , \23472 , \23473 , \23474 ,
         \23475 , \23476 , \23477 , \23478 , \23479 , \23480 , \23481 , \23482 , \23483 , \23484 ,
         \23485 , \23486 , \23487 , \23488 , \23489 , \23490 , \23491 , \23492 , \23493 , \23494 ,
         \23495 , \23496 , \23497 , \23498 , \23499 , \23500 , \23501 , \23502 , \23503 , \23504 ,
         \23505 , \23506 , \23507 , \23508 , \23509 , \23510 , \23511 , \23512 , \23513 , \23514 ,
         \23515 , \23516 , \23517 , \23518 , \23519 , \23520 , \23521 , \23522 , \23523 , \23524 ,
         \23525 , \23526 , \23527 , \23528 , \23529 , \23530 , \23531 , \23532 , \23533 , \23534 ,
         \23535 , \23536 , \23537 , \23538 , \23539 , \23540 , \23541 , \23542 , \23543 , \23544 ,
         \23545 , \23546 , \23547 , \23548 , \23549 , \23550 , \23551 , \23552 , \23553 , \23554 ,
         \23555 , \23556 , \23557 , \23558 , \23559 , \23560 , \23561 , \23562 , \23563 , \23564 ,
         \23565 , \23566 , \23567 , \23568 , \23569 , \23570 , \23571 , \23572 , \23573 , \23574 ,
         \23575 , \23576 , \23577 , \23578 , \23579 , \23580 , \23581 , \23582 , \23583 , \23584 ,
         \23585 , \23586 , \23587 , \23588 , \23589 , \23590 , \23591 , \23592 , \23593 , \23594 ,
         \23595 , \23596 , \23597 , \23598 , \23599 , \23600 , \23601 , \23602 , \23603 , \23604 ,
         \23605 , \23606 , \23607 , \23608 , \23609 , \23610 , \23611 , \23612 , \23613 , \23614 ,
         \23615 , \23616 , \23617 , \23618 , \23619 , \23620 , \23621 , \23622 , \23623 , \23624 ,
         \23625 , \23626 , \23627 , \23628 , \23629 , \23630 , \23631 , \23632 , \23633 , \23634 ,
         \23635 , \23636 , \23637 , \23638 , \23639 , \23640 , \23641 , \23642 , \23643 , \23644 ,
         \23645 , \23646 , \23647 , \23648 , \23649 , \23650 , \23651 , \23652 , \23653 , \23654 ,
         \23655 , \23656 , \23657 , \23658 , \23659 , \23660 , \23661 , \23662 , \23663 , \23664 ,
         \23665 , \23666 , \23667 , \23668 , \23669 , \23670 , \23671 , \23672 , \23673 , \23674 ,
         \23675 , \23676 , \23677 , \23678 , \23679 , \23680 , \23681 , \23682 , \23683 , \23684 ,
         \23685 , \23686 , \23687 , \23688 , \23689 , \23690 , \23691 , \23692 , \23693 , \23694 ,
         \23695 , \23696 , \23697 , \23698 , \23699 , \23700 , \23701 , \23702 , \23703 , \23704 ,
         \23705 , \23706 , \23707 , \23708 , \23709 , \23710 , \23711 , \23712 , \23713 , \23714 ,
         \23715 , \23716 , \23717 , \23718 , \23719 , \23720 , \23721 , \23722 , \23723 , \23724 ,
         \23725 , \23726 , \23727 , \23728 , \23729 , \23730 , \23731 , \23732 , \23733 , \23734 ,
         \23735 , \23736 , \23737 , \23738 , \23739 , \23740 , \23741 , \23742 , \23743 , \23744 ,
         \23745 , \23746 , \23747 , \23748 , \23749 , \23750 , \23751 , \23752 , \23753 , \23754 ,
         \23755 , \23756 , \23757 , \23758 , \23759 , \23760 , \23761 , \23762 , \23763 , \23764 ,
         \23765 , \23766 , \23767 , \23768 , \23769 , \23770 , \23771 , \23772 , \23773 , \23774 ,
         \23775 , \23776 , \23777 , \23778 , \23779 , \23780 , \23781 , \23782 , \23783 , \23784 ,
         \23785 , \23786 , \23787 , \23788 , \23789 , \23790 , \23791 , \23792 , \23793 , \23794 ,
         \23795 , \23796 , \23797 , \23798 , \23799 , \23800 , \23801 , \23802 , \23803 , \23804 ,
         \23805 , \23806 , \23807 , \23808 , \23809 , \23810 , \23811 , \23812 , \23813 , \23814 ,
         \23815 , \23816 , \23817 , \23818 , \23819 , \23820 , \23821 , \23822 , \23823 , \23824 ,
         \23825 , \23826 , \23827 , \23828 , \23829 , \23830 , \23831 , \23832 , \23833 , \23834 ,
         \23835 , \23836 , \23837 , \23838 , \23839 , \23840 , \23841 , \23842 , \23843 , \23844 ,
         \23845 , \23846 , \23847 , \23848 , \23849 , \23850 , \23851 , \23852 , \23853 , \23854 ,
         \23855 , \23856 , \23857 , \23858 , \23859 , \23860 , \23861 , \23862 , \23863 , \23864 ,
         \23865 , \23866 , \23867 , \23868 , \23869 , \23870 , \23871 , \23872 , \23873 , \23874 ,
         \23875 , \23876 , \23877 , \23878 , \23879 , \23880 , \23881 , \23882 , \23883 , \23884 ,
         \23885 , \23886 , \23887 , \23888 , \23889 , \23890 , \23891 , \23892 , \23893 , \23894 ,
         \23895 , \23896 , \23897 , \23898 , \23899 , \23900 , \23901 , \23902 , \23903 , \23904 ,
         \23905 , \23906 , \23907 , \23908 , \23909 , \23910 , \23911 , \23912 , \23913 , \23914 ,
         \23915 , \23916 , \23917 , \23918 , \23919 , \23920 , \23921 , \23922 , \23923 , \23924 ,
         \23925 , \23926 , \23927 , \23928 , \23929 , \23930 , \23931 , \23932 , \23933 , \23934 ,
         \23935 , \23936 , \23937 , \23938 , \23939 , \23940 , \23941 , \23942 , \23943 , \23944 ,
         \23945 , \23946 , \23947 , \23948 , \23949 , \23950 , \23951 , \23952 , \23953 , \23954 ,
         \23955 , \23956 , \23957 , \23958 , \23959 , \23960 , \23961 , \23962 , \23963 , \23964 ,
         \23965 , \23966 , \23967 , \23968 , \23969 , \23970 , \23971 , \23972 , \23973 , \23974 ,
         \23975 , \23976 , \23977 , \23978 , \23979 , \23980 , \23981 , \23982 , \23983 , \23984 ,
         \23985 , \23986 , \23987 , \23988 , \23989 , \23990 , \23991 , \23992 , \23993 , \23994 ,
         \23995 , \23996 , \23997 , \23998 , \23999 , \24000 , \24001 , \24002 , \24003 , \24004 ,
         \24005 , \24006 , \24007 , \24008 , \24009 , \24010 , \24011 , \24012 , \24013 , \24014 ,
         \24015 , \24016 , \24017 , \24018 , \24019 , \24020 , \24021 , \24022 , \24023 , \24024 ,
         \24025 , \24026 , \24027 , \24028 , \24029 , \24030 , \24031 , \24032 , \24033 , \24034 ,
         \24035 , \24036 , \24037 , \24038 , \24039 , \24040 , \24041 , \24042 , \24043 , \24044 ,
         \24045 , \24046 , \24047 , \24048 , \24049 , \24050 , \24051 , \24052 , \24053 , \24054 ,
         \24055 , \24056 , \24057 , \24058 , \24059 , \24060 , \24061 , \24062 , \24063 , \24064 ,
         \24065 , \24066 , \24067 , \24068 , \24069 , \24070 , \24071 , \24072 , \24073 , \24074 ,
         \24075 , \24076 , \24077 , \24078 , \24079 , \24080 , \24081 , \24082 , \24083 , \24084 ,
         \24085 , \24086 , \24087 , \24088 , \24089 , \24090 , \24091 , \24092 , \24093 , \24094 ,
         \24095 , \24096 , \24097 , \24098 , \24099 , \24100 , \24101 , \24102 , \24103 , \24104 ,
         \24105 , \24106 , \24107 , \24108 , \24109 , \24110 , \24111 , \24112 , \24113 , \24114 ,
         \24115 , \24116 , \24117 , \24118 , \24119 , \24120 , \24121 , \24122 , \24123 , \24124 ,
         \24125 , \24126 , \24127 , \24128 , \24129 , \24130 , \24131 , \24132 , \24133 , \24134 ,
         \24135 , \24136 , \24137 , \24138 , \24139 , \24140 , \24141 , \24142 , \24143 , \24144 ,
         \24145 , \24146 , \24147 , \24148 , \24149 , \24150 , \24151 , \24152 , \24153 , \24154 ,
         \24155 , \24156 , \24157 , \24158 , \24159 , \24160 , \24161 , \24162 , \24163 , \24164 ,
         \24165 , \24166 , \24167 , \24168 , \24169 , \24170 , \24171 , \24172 , \24173 , \24174 ,
         \24175 , \24176 , \24177 , \24178 , \24179 , \24180 , \24181 , \24182 , \24183 , \24184 ,
         \24185 , \24186 , \24187 , \24188 , \24189 , \24190 , \24191 , \24192 , \24193 , \24194 ,
         \24195 , \24196 , \24197 , \24198 , \24199 , \24200 , \24201 , \24202 , \24203 , \24204 ,
         \24205 , \24206 , \24207 , \24208 , \24209 , \24210 , \24211 , \24212 , \24213 , \24214 ,
         \24215 , \24216 , \24217 , \24218 , \24219 , \24220 , \24221 , \24222 , \24223 , \24224 ,
         \24225 , \24226 , \24227 , \24228 , \24229 , \24230 , \24231 , \24232 , \24233 , \24234 ,
         \24235 , \24236 , \24237 , \24238 , \24239 , \24240 , \24241 , \24242 , \24243 , \24244 ,
         \24245 , \24246 , \24247 , \24248 , \24249 , \24250 , \24251 , \24252 , \24253 , \24254 ,
         \24255 , \24256 , \24257 , \24258 , \24259 , \24260 , \24261 , \24262 , \24263 , \24264 ,
         \24265 , \24266 , \24267 , \24268 , \24269 , \24270 , \24271 , \24272 , \24273 , \24274 ,
         \24275 , \24276 , \24277 , \24278 , \24279 , \24280 , \24281 , \24282 , \24283 , \24284 ,
         \24285 , \24286 , \24287 , \24288 , \24289 , \24290 , \24291 , \24292 , \24293 , \24294 ,
         \24295 , \24296 , \24297 , \24298 , \24299 , \24300 , \24301 , \24302 , \24303 , \24304 ,
         \24305 , \24306 , \24307 , \24308 , \24309 , \24310 , \24311 , \24312 , \24313 , \24314 ,
         \24315 , \24316 , \24317 , \24318 , \24319 , \24320 , \24321 , \24322 , \24323 , \24324 ,
         \24325 , \24326 , \24327 , \24328 , \24329 , \24330 , \24331 , \24332 , \24333 , \24334 ,
         \24335 , \24336 , \24337 , \24338 , \24339 , \24340 , \24341 , \24342 , \24343 , \24344 ,
         \24345 , \24346 , \24347 , \24348 , \24349 , \24350 , \24351 , \24352 , \24353 , \24354 ,
         \24355 , \24356 , \24357 , \24358 , \24359 , \24360 , \24361 , \24362 , \24363 , \24364 ,
         \24365 , \24366 , \24367 , \24368 , \24369 , \24370 , \24371 , \24372 , \24373 , \24374 ,
         \24375 , \24376 , \24377 , \24378 , \24379 , \24380 , \24381 , \24382 , \24383 , \24384 ,
         \24385 , \24386 , \24387 , \24388 , \24389 , \24390 , \24391 , \24392 , \24393 , \24394 ,
         \24395 , \24396 , \24397 , \24398 , \24399 , \24400 , \24401 , \24402 , \24403 , \24404 ,
         \24405 , \24406 , \24407 , \24408 , \24409 , \24410 , \24411 , \24412 , \24413 , \24414 ,
         \24415 , \24416 , \24417 , \24418 , \24419 , \24420 , \24421 , \24422 , \24423 , \24424 ,
         \24425 , \24426 , \24427 , \24428 , \24429 , \24430 , \24431 , \24432 , \24433 , \24434 ,
         \24435 , \24436 , \24437 , \24438 , \24439 , \24440 , \24441 , \24442 , \24443 , \24444 ,
         \24445 , \24446 , \24447 , \24448 , \24449 , \24450 , \24451 , \24452 , \24453 , \24454 ,
         \24455 , \24456 , \24457 , \24458 , \24459 , \24460 , \24461 , \24462 , \24463 , \24464 ,
         \24465 , \24466 , \24467 , \24468 , \24469 , \24470 , \24471 , \24472 , \24473 , \24474 ,
         \24475 , \24476 , \24477 , \24478 , \24479 , \24480 , \24481 , \24482 , \24483 , \24484 ,
         \24485 , \24486 , \24487 , \24488 , \24489 , \24490 , \24491 , \24492 , \24493 , \24494 ,
         \24495 , \24496 , \24497 , \24498 , \24499 , \24500 , \24501 , \24502 , \24503 , \24504 ,
         \24505 , \24506 , \24507 , \24508 , \24509 , \24510 , \24511 , \24512 , \24513 , \24514 ,
         \24515 , \24516 , \24517 , \24518 , \24519 , \24520 , \24521 , \24522 , \24523 , \24524 ,
         \24525 , \24526 , \24527 , \24528 , \24529 , \24530 , \24531 , \24532 , \24533 , \24534 ,
         \24535 , \24536 , \24537 , \24538 , \24539 , \24540 , \24541 , \24542 , \24543 , \24544 ,
         \24545 , \24546 , \24547 , \24548 , \24549 , \24550 , \24551 , \24552 , \24553 , \24554 ,
         \24555 , \24556 , \24557 , \24558 , \24559 , \24560 , \24561 , \24562 , \24563 , \24564 ,
         \24565 , \24566 , \24567 , \24568 , \24569 , \24570 , \24571 , \24572 , \24573 , \24574 ,
         \24575 , \24576 , \24577 , \24578 , \24579 , \24580 , \24581 , \24582 , \24583 , \24584 ,
         \24585 , \24586 , \24587 , \24588 , \24589 , \24590 , \24591 , \24592 , \24593 , \24594 ,
         \24595 , \24596 , \24597 , \24598 , \24599 , \24600 , \24601 , \24602 , \24603 , \24604 ,
         \24605 , \24606 , \24607 , \24608 , \24609 , \24610 , \24611 , \24612 , \24613 , \24614 ,
         \24615 , \24616 , \24617 , \24618 , \24619 , \24620 , \24621 , \24622 , \24623 , \24624 ,
         \24625 , \24626 , \24627 , \24628 , \24629 , \24630 , \24631 , \24632 , \24633 , \24634 ,
         \24635 , \24636 , \24637 , \24638 , \24639 , \24640 , \24641 , \24642 , \24643 , \24644 ,
         \24645 , \24646 , \24647 , \24648 , \24649 , \24650 , \24651 , \24652 , \24653 , \24654 ,
         \24655 , \24656 , \24657 , \24658 , \24659 , \24660 , \24661 , \24662 , \24663 , \24664 ,
         \24665 , \24666 , \24667 , \24668 , \24669 , \24670 , \24671 , \24672 , \24673 , \24674 ,
         \24675 , \24676 , \24677 , \24678 , \24679 , \24680 , \24681 , \24682 , \24683 , \24684 ,
         \24685 , \24686 , \24687 , \24688 , \24689 , \24690 , \24691 , \24692 , \24693 , \24694 ,
         \24695 , \24696 , \24697 , \24698 , \24699 , \24700 , \24701 , \24702 , \24703 , \24704 ,
         \24705 , \24706 , \24707 , \24708 , \24709 , \24710 , \24711 , \24712 , \24713 , \24714 ,
         \24715 , \24716 , \24717 , \24718 , \24719 , \24720 , \24721 , \24722 , \24723 , \24724 ,
         \24725 , \24726 , \24727 , \24728 , \24729 , \24730 , \24731 , \24732 , \24733 , \24734 ,
         \24735 , \24736 , \24737 , \24738 , \24739 , \24740 , \24741 , \24742 , \24743 , \24744 ,
         \24745 , \24746 , \24747 , \24748 , \24749 , \24750 , \24751 , \24752 , \24753 , \24754 ,
         \24755 , \24756 , \24757 , \24758 , \24759 , \24760 , \24761 , \24762 , \24763 , \24764 ,
         \24765 , \24766 , \24767 , \24768 , \24769 , \24770 , \24771 , \24772 , \24773 , \24774 ,
         \24775 , \24776 , \24777 , \24778 , \24779 , \24780 , \24781 , \24782 , \24783 , \24784 ,
         \24785 , \24786 , \24787 , \24788 , \24789 , \24790 , \24791 , \24792 , \24793 , \24794 ,
         \24795 , \24796 , \24797 , \24798 , \24799 , \24800 , \24801 , \24802 , \24803 , \24804 ,
         \24805 , \24806 , \24807 , \24808 , \24809 , \24810 , \24811 , \24812 , \24813 , \24814 ,
         \24815 , \24816 , \24817 , \24818 , \24819 , \24820 , \24821 , \24822 , \24823 , \24824 ,
         \24825 , \24826 , \24827 , \24828 , \24829 , \24830 , \24831 , \24832 , \24833 , \24834 ,
         \24835 , \24836 , \24837 , \24838 , \24839 , \24840 , \24841 , \24842 , \24843 , \24844 ,
         \24845 , \24846 , \24847 , \24848 , \24849 , \24850 , \24851 , \24852 , \24853 , \24854 ,
         \24855 , \24856 , \24857 , \24858 , \24859 , \24860 , \24861 , \24862 , \24863 , \24864 ,
         \24865 , \24866 , \24867 , \24868 , \24869 , \24870 , \24871 , \24872 , \24873 , \24874 ,
         \24875 , \24876 , \24877 , \24878 , \24879 , \24880 , \24881 , \24882 , \24883 , \24884 ,
         \24885 , \24886 , \24887 , \24888 , \24889 , \24890 , \24891 , \24892 , \24893 , \24894 ,
         \24895 , \24896 , \24897 , \24898 , \24899 , \24900 , \24901 , \24902 , \24903 , \24904 ,
         \24905 , \24906 , \24907 , \24908 , \24909 , \24910 , \24911 , \24912 , \24913 , \24914 ,
         \24915 , \24916 , \24917 , \24918 , \24919 , \24920 , \24921 , \24922 , \24923 , \24924 ,
         \24925 , \24926 , \24927 , \24928 , \24929 , \24930 , \24931 , \24932 , \24933 , \24934 ,
         \24935 , \24936 , \24937 , \24938 , \24939 , \24940 , \24941 , \24942 , \24943 , \24944 ,
         \24945 , \24946 , \24947 , \24948 , \24949 , \24950 , \24951 , \24952 , \24953 , \24954 ,
         \24955 , \24956 , \24957 , \24958 , \24959 , \24960 , \24961 , \24962 , \24963 , \24964 ,
         \24965 , \24966 , \24967 , \24968 , \24969 , \24970 , \24971 , \24972 , \24973 , \24974 ,
         \24975 , \24976 , \24977 , \24978 , \24979 , \24980 , \24981 , \24982 , \24983 , \24984 ,
         \24985 , \24986 , \24987 , \24988 , \24989 , \24990 , \24991 , \24992 , \24993 , \24994 ,
         \24995 , \24996 , \24997 , \24998 , \24999 , \25000 , \25001 , \25002 , \25003 , \25004 ,
         \25005 , \25006 , \25007 , \25008 , \25009 , \25010 , \25011 , \25012 , \25013 , \25014 ,
         \25015 , \25016 , \25017 , \25018 , \25019 , \25020 , \25021 , \25022 , \25023 , \25024 ,
         \25025 , \25026 , \25027 , \25028 , \25029 , \25030 , \25031 , \25032 , \25033 , \25034 ,
         \25035 , \25036 , \25037 , \25038 , \25039 , \25040 , \25041 , \25042 , \25043 , \25044 ,
         \25045 , \25046 , \25047 , \25048 , \25049 , \25050 , \25051 , \25052 , \25053 , \25054 ,
         \25055 , \25056 , \25057 , \25058 , \25059 , \25060 , \25061 , \25062 , \25063 , \25064 ,
         \25065 , \25066 , \25067 , \25068 , \25069 , \25070 , \25071 , \25072 , \25073 , \25074 ,
         \25075 , \25076 , \25077 , \25078 , \25079 , \25080 , \25081 , \25082 , \25083 , \25084 ,
         \25085 , \25086 , \25087 , \25088 , \25089 , \25090 , \25091 , \25092 , \25093 , \25094 ,
         \25095 , \25096 , \25097 , \25098 , \25099 , \25100 , \25101 , \25102 , \25103 , \25104 ,
         \25105 , \25106 , \25107 , \25108 , \25109 , \25110 , \25111 , \25112 , \25113 , \25114 ,
         \25115 , \25116 , \25117 , \25118 , \25119 , \25120 , \25121 , \25122 , \25123 , \25124 ,
         \25125 , \25126 , \25127 , \25128 , \25129 , \25130 , \25131 , \25132 , \25133 , \25134 ,
         \25135 , \25136 , \25137 , \25138 , \25139 , \25140 , \25141 , \25142 , \25143 , \25144 ,
         \25145 , \25146 , \25147 , \25148 , \25149 , \25150 , \25151 , \25152 , \25153 , \25154 ,
         \25155 , \25156 , \25157 , \25158 , \25159 , \25160 , \25161 , \25162 , \25163 , \25164 ,
         \25165 , \25166 , \25167 , \25168 , \25169 , \25170 , \25171 , \25172 , \25173 , \25174 ,
         \25175 , \25176 , \25177 , \25178 , \25179 , \25180 , \25181 , \25182 , \25183 , \25184 ,
         \25185 , \25186 , \25187 , \25188 , \25189 , \25190 , \25191 , \25192 , \25193 , \25194 ,
         \25195 , \25196 , \25197 , \25198 , \25199 , \25200 , \25201 , \25202 , \25203 , \25204 ,
         \25205 , \25206 , \25207 , \25208 , \25209 , \25210 , \25211 , \25212 , \25213 , \25214 ,
         \25215 , \25216 , \25217 , \25218 , \25219 , \25220 , \25221 , \25222 , \25223 , \25224 ,
         \25225 , \25226 , \25227 , \25228 , \25229 , \25230 , \25231 , \25232 , \25233 , \25234 ,
         \25235 , \25236 , \25237 , \25238 , \25239 , \25240 , \25241 , \25242 , \25243 , \25244 ,
         \25245 , \25246 , \25247 , \25248 , \25249 , \25250 , \25251 , \25252 , \25253 , \25254 ,
         \25255 , \25256 , \25257 , \25258 , \25259 , \25260 , \25261 , \25262 , \25263 , \25264 ,
         \25265 , \25266 , \25267 , \25268 , \25269 , \25270 , \25271 , \25272 , \25273 , \25274 ,
         \25275 , \25276 , \25277 , \25278 , \25279 , \25280 , \25281 , \25282 , \25283 , \25284 ,
         \25285 , \25286 , \25287 , \25288 , \25289 , \25290 , \25291 , \25292 , \25293 , \25294 ,
         \25295 , \25296 , \25297 , \25298 , \25299 , \25300 , \25301 , \25302 , \25303 , \25304 ,
         \25305 , \25306 , \25307 , \25308 , \25309 , \25310 , \25311 , \25312 , \25313 , \25314 ,
         \25315 , \25316 , \25317 , \25318 , \25319 , \25320 , \25321 , \25322 , \25323 , \25324 ,
         \25325 , \25326 , \25327 , \25328 , \25329 , \25330 , \25331 , \25332 , \25333 , \25334 ,
         \25335 , \25336 , \25337 , \25338 , \25339 , \25340 , \25341 , \25342 , \25343 , \25344 ,
         \25345 , \25346 , \25347 , \25348 , \25349 , \25350 , \25351 , \25352 , \25353 , \25354 ,
         \25355 , \25356 , \25357 , \25358 , \25359 , \25360 , \25361 , \25362 , \25363 , \25364 ,
         \25365 , \25366 , \25367 , \25368 , \25369 , \25370 , \25371 , \25372 , \25373 , \25374 ,
         \25375 , \25376 , \25377 , \25378 , \25379 , \25380 , \25381 , \25382 , \25383 , \25384 ,
         \25385 , \25386 , \25387 , \25388 , \25389 , \25390 , \25391 , \25392 , \25393 , \25394 ,
         \25395 , \25396 , \25397 , \25398 , \25399 , \25400 , \25401 , \25402 , \25403 , \25404 ,
         \25405 , \25406 , \25407 , \25408 , \25409 , \25410 , \25411 , \25412 , \25413 , \25414 ,
         \25415 , \25416 , \25417 , \25418 , \25419 , \25420 , \25421 , \25422 , \25423 , \25424 ,
         \25425 , \25426 , \25427 , \25428 , \25429 , \25430 , \25431 , \25432 , \25433 , \25434 ,
         \25435 , \25436 , \25437 , \25438 , \25439 , \25440 , \25441 , \25442 , \25443 , \25444 ,
         \25445 , \25446 , \25447 , \25448 , \25449 , \25450 , \25451 , \25452 , \25453 , \25454 ,
         \25455 , \25456 , \25457 , \25458 , \25459 , \25460 , \25461 , \25462 , \25463 , \25464 ,
         \25465 , \25466 , \25467 , \25468 , \25469 , \25470 , \25471 , \25472 , \25473 , \25474 ,
         \25475 , \25476 , \25477 , \25478 , \25479 , \25480 , \25481 , \25482 , \25483 , \25484 ,
         \25485 , \25486 , \25487 , \25488 , \25489 , \25490 , \25491 , \25492 , \25493 , \25494 ,
         \25495 , \25496 , \25497 , \25498 , \25499 , \25500 , \25501 , \25502 , \25503 , \25504 ,
         \25505 , \25506 , \25507 , \25508 , \25509 , \25510 , \25511 , \25512 , \25513 , \25514 ,
         \25515 , \25516 , \25517 , \25518 , \25519 , \25520 , \25521 , \25522 , \25523 , \25524 ,
         \25525 , \25526 , \25527 , \25528 , \25529 , \25530 , \25531 , \25532 , \25533 , \25534 ,
         \25535 , \25536 , \25537 , \25538 , \25539 , \25540 , \25541 , \25542 , \25543 , \25544 ,
         \25545 , \25546 , \25547 , \25548 , \25549 , \25550 , \25551 , \25552 , \25553 , \25554 ,
         \25555 , \25556 , \25557 , \25558 , \25559 , \25560 , \25561 , \25562 , \25563 , \25564 ,
         \25565 , \25566 , \25567 , \25568 , \25569 , \25570 , \25571 , \25572 , \25573 , \25574 ,
         \25575 , \25576 , \25577 , \25578 , \25579 , \25580 , \25581 , \25582 , \25583 , \25584 ,
         \25585 , \25586 , \25587 , \25588 , \25589 , \25590 , \25591 , \25592 , \25593 , \25594 ,
         \25595 , \25596 , \25597 , \25598 , \25599 , \25600 , \25601 , \25602 , \25603 , \25604 ,
         \25605 , \25606 , \25607 , \25608 , \25609 , \25610 , \25611 , \25612 , \25613 , \25614 ,
         \25615 , \25616 , \25617 , \25618 , \25619 , \25620 , \25621 , \25622 , \25623 , \25624 ,
         \25625 , \25626 , \25627 , \25628 , \25629 , \25630 , \25631 , \25632 , \25633 , \25634 ,
         \25635 , \25636 , \25637 , \25638 , \25639 , \25640 , \25641 , \25642 , \25643 , \25644 ,
         \25645 , \25646 , \25647 , \25648 , \25649 , \25650 , \25651 , \25652 , \25653 , \25654 ,
         \25655 , \25656 , \25657 , \25658 , \25659 , \25660 , \25661 , \25662 , \25663 , \25664 ,
         \25665 , \25666 , \25667 , \25668 , \25669 , \25670 , \25671 , \25672 , \25673 , \25674 ,
         \25675 , \25676 , \25677 , \25678 , \25679 , \25680 , \25681 , \25682 , \25683 , \25684 ,
         \25685 , \25686 , \25687 , \25688 , \25689 , \25690 , \25691 , \25692 , \25693 , \25694 ,
         \25695 , \25696 , \25697 , \25698 , \25699 , \25700 , \25701 , \25702 , \25703 , \25704 ,
         \25705 , \25706 , \25707 , \25708 , \25709 , \25710 , \25711 , \25712 , \25713 , \25714 ,
         \25715 , \25716 , \25717 , \25718 , \25719 , \25720 , \25721 , \25722 , \25723 , \25724 ,
         \25725 , \25726 , \25727 , \25728 , \25729 , \25730 , \25731 , \25732 , \25733 , \25734 ,
         \25735 , \25736 , \25737 , \25738 , \25739 , \25740 , \25741 , \25742 , \25743 , \25744 ,
         \25745 , \25746 , \25747 , \25748 , \25749 , \25750 , \25751 , \25752 , \25753 , \25754 ,
         \25755 , \25756 , \25757 , \25758 , \25759 , \25760 , \25761 , \25762 , \25763 , \25764 ,
         \25765 , \25766 , \25767 , \25768 , \25769 , \25770 , \25771 , \25772 , \25773 , \25774 ,
         \25775 , \25776 , \25777 , \25778 , \25779 , \25780 , \25781 , \25782 , \25783 , \25784 ,
         \25785 , \25786 , \25787 , \25788 , \25789 , \25790 , \25791 , \25792 , \25793 , \25794 ,
         \25795 , \25796 , \25797 , \25798 , \25799 , \25800 , \25801 , \25802 , \25803 , \25804 ,
         \25805 , \25806 , \25807 , \25808 , \25809 , \25810 , \25811 , \25812 , \25813 , \25814 ,
         \25815 , \25816 , \25817 , \25818 , \25819 , \25820 , \25821 , \25822 , \25823 , \25824 ,
         \25825 , \25826 , \25827 , \25828 , \25829 , \25830 , \25831 , \25832 , \25833 , \25834 ,
         \25835 , \25836 , \25837 , \25838 , \25839 , \25840 , \25841 , \25842 , \25843 , \25844 ,
         \25845 , \25846 , \25847 , \25848 , \25849 , \25850 , \25851 , \25852 , \25853 , \25854 ,
         \25855 , \25856 , \25857 , \25858 , \25859 , \25860 , \25861 , \25862 , \25863 , \25864 ,
         \25865 , \25866 , \25867 , \25868 , \25869 , \25870 , \25871 , \25872 , \25873 , \25874 ,
         \25875 , \25876 , \25877 , \25878 , \25879 , \25880 , \25881 , \25882 , \25883 , \25884 ,
         \25885 , \25886 , \25887 , \25888 , \25889 , \25890 , \25891 , \25892 , \25893 , \25894 ,
         \25895 , \25896 , \25897 , \25898 , \25899 , \25900 , \25901 , \25902 , \25903 , \25904 ,
         \25905 , \25906 , \25907 , \25908 , \25909 , \25910 , \25911 , \25912 , \25913 , \25914 ,
         \25915 , \25916 , \25917 , \25918 , \25919 , \25920 , \25921 , \25922 , \25923 , \25924 ,
         \25925 , \25926 , \25927 , \25928 , \25929 , \25930 , \25931 , \25932 , \25933 , \25934 ,
         \25935 , \25936 , \25937 , \25938 , \25939 , \25940 , \25941 , \25942 , \25943 , \25944 ,
         \25945 , \25946 , \25947 , \25948 , \25949 , \25950 , \25951 , \25952 , \25953 , \25954 ,
         \25955 , \25956 , \25957 , \25958 , \25959 , \25960 , \25961 , \25962 , \25963 , \25964 ,
         \25965 , \25966 , \25967 , \25968 , \25969 , \25970 , \25971 , \25972 , \25973 , \25974 ,
         \25975 , \25976 , \25977 , \25978 , \25979 , \25980 , \25981 , \25982 , \25983 , \25984 ,
         \25985 , \25986 , \25987 , \25988 , \25989 , \25990 , \25991 , \25992 , \25993 , \25994 ,
         \25995 , \25996 , \25997 , \25998 , \25999 , \26000 , \26001 , \26002 , \26003 , \26004 ,
         \26005 , \26006 , \26007 , \26008 , \26009 , \26010 , \26011 , \26012 , \26013 , \26014 ,
         \26015 , \26016 , \26017 , \26018 , \26019 , \26020 , \26021 , \26022 , \26023 , \26024 ,
         \26025 , \26026 , \26027 , \26028 , \26029 , \26030 , \26031 , \26032 , \26033 , \26034 ,
         \26035 , \26036 , \26037 , \26038 , \26039 , \26040 , \26041 , \26042 , \26043 , \26044 ,
         \26045 , \26046 , \26047 , \26048 , \26049 , \26050 , \26051 , \26052 , \26053 , \26054 ,
         \26055 , \26056 , \26057 , \26058 , \26059 , \26060 , \26061 , \26062 , \26063 , \26064 ,
         \26065 , \26066 , \26067 , \26068 , \26069 , \26070 , \26071 , \26072 , \26073 , \26074 ,
         \26075 , \26076 , \26077 , \26078 , \26079 , \26080 , \26081 , \26082 , \26083 , \26084 ,
         \26085 , \26086 , \26087 , \26088 , \26089 , \26090 , \26091 , \26092 , \26093 , \26094 ,
         \26095 , \26096 , \26097 , \26098 , \26099 , \26100 , \26101 , \26102 , \26103 , \26104 ,
         \26105 , \26106 , \26107 , \26108 , \26109 , \26110 , \26111 , \26112 , \26113 , \26114 ,
         \26115 , \26116 , \26117 , \26118 , \26119 , \26120 , \26121 , \26122 , \26123 , \26124 ,
         \26125 , \26126 , \26127 , \26128 , \26129 , \26130 , \26131 , \26132 , \26133 , \26134 ,
         \26135 , \26136 , \26137 , \26138 , \26139 , \26140 , \26141 , \26142 , \26143 , \26144 ,
         \26145 , \26146 , \26147 , \26148 , \26149 , \26150 , \26151 , \26152 , \26153 , \26154 ,
         \26155 , \26156 , \26157 , \26158 , \26159 , \26160 , \26161 , \26162 , \26163 , \26164 ,
         \26165 , \26166 , \26167 , \26168 , \26169 , \26170 , \26171 , \26172 , \26173 , \26174 ,
         \26175 , \26176 , \26177 , \26178 , \26179 , \26180 , \26181 , \26182 , \26183 , \26184 ,
         \26185 , \26186 , \26187 , \26188 , \26189 , \26190 , \26191 , \26192 , \26193 , \26194 ,
         \26195 , \26196 , \26197 , \26198 , \26199 , \26200 , \26201 , \26202 , \26203 , \26204 ,
         \26205 , \26206 , \26207 , \26208 , \26209 , \26210 , \26211 , \26212 , \26213 , \26214 ,
         \26215 , \26216 , \26217 , \26218 , \26219 , \26220 , \26221 , \26222 , \26223 , \26224 ,
         \26225 , \26226 , \26227 , \26228 , \26229 , \26230 , \26231 , \26232 , \26233 , \26234 ,
         \26235 , \26236 , \26237 , \26238 , \26239 , \26240 , \26241 , \26242 , \26243 , \26244 ,
         \26245 , \26246 , \26247 , \26248 , \26249 , \26250 , \26251 , \26252 , \26253 , \26254 ,
         \26255 , \26256 , \26257 , \26258 , \26259 , \26260 , \26261 , \26262 , \26263 , \26264 ,
         \26265 , \26266 , \26267 , \26268 , \26269 , \26270 , \26271 , \26272 , \26273 , \26274 ,
         \26275 , \26276 , \26277 , \26278 , \26279 , \26280 , \26281 , \26282 , \26283 , \26284 ,
         \26285 , \26286 , \26287 , \26288 , \26289 , \26290 , \26291 , \26292 , \26293 , \26294 ,
         \26295 , \26296 , \26297 , \26298 , \26299 , \26300 , \26301 , \26302 , \26303 , \26304 ,
         \26305 , \26306 , \26307 , \26308 , \26309 , \26310 , \26311 , \26312 , \26313 , \26314 ,
         \26315 , \26316 , \26317 , \26318 , \26319 , \26320 , \26321 , \26322 , \26323 , \26324 ,
         \26325 , \26326 , \26327 , \26328 , \26329 , \26330 , \26331 , \26332 , \26333 , \26334 ,
         \26335 , \26336 , \26337 , \26338 , \26339 , \26340 , \26341 , \26342 , \26343 , \26344 ,
         \26345 , \26346 , \26347 , \26348 , \26349 , \26350 , \26351 , \26352 , \26353 , \26354 ,
         \26355 , \26356 , \26357 , \26358 , \26359 , \26360 , \26361 , \26362 , \26363 , \26364 ,
         \26365 , \26366 , \26367 , \26368 , \26369 , \26370 , \26371 , \26372 , \26373 , \26374 ,
         \26375 , \26376 , \26377 , \26378 , \26379 , \26380 , \26381 , \26382 , \26383 , \26384 ,
         \26385 , \26386 , \26387 , \26388 , \26389 , \26390 , \26391 , \26392 , \26393 , \26394 ,
         \26395 , \26396 , \26397 , \26398 , \26399 , \26400 , \26401 , \26402 , \26403 , \26404 ,
         \26405 , \26406 , \26407 , \26408 , \26409 , \26410 , \26411 , \26412 , \26413 , \26414 ,
         \26415 , \26416 , \26417 , \26418 , \26419 , \26420 , \26421 , \26422 , \26423 , \26424 ,
         \26425 , \26426 , \26427 , \26428 , \26429 , \26430 , \26431 , \26432 , \26433 , \26434 ,
         \26435 , \26436 , \26437 , \26438 , \26439 , \26440 , \26441 , \26442 , \26443 , \26444 ,
         \26445 , \26446 , \26447 , \26448 , \26449 , \26450 , \26451 , \26452 , \26453 , \26454 ,
         \26455 , \26456 , \26457 , \26458 , \26459 , \26460 , \26461 , \26462 , \26463 , \26464 ,
         \26465 , \26466 , \26467 , \26468 , \26469 , \26470 , \26471 , \26472 , \26473 , \26474 ,
         \26475 , \26476 , \26477 , \26478 , \26479 , \26480 , \26481 , \26482 , \26483 , \26484 ,
         \26485 , \26486 , \26487 , \26488 , \26489 , \26490 , \26491 , \26492 , \26493 , \26494 ,
         \26495 , \26496 , \26497 , \26498 , \26499 , \26500 , \26501 , \26502 , \26503 , \26504 ,
         \26505 , \26506 , \26507 , \26508 , \26509 , \26510 , \26511 , \26512 , \26513 , \26514 ,
         \26515 , \26516 , \26517 , \26518 , \26519 , \26520 , \26521 , \26522 , \26523 , \26524 ,
         \26525 , \26526 , \26527 , \26528 , \26529 , \26530 , \26531 , \26532 , \26533 , \26534 ,
         \26535 , \26536 , \26537 , \26538 , \26539 , \26540 , \26541 , \26542 , \26543 , \26544 ,
         \26545 , \26546 , \26547 , \26548 , \26549 , \26550 , \26551 , \26552 , \26553 , \26554 ,
         \26555 , \26556 , \26557 , \26558 , \26559 , \26560 , \26561 , \26562 , \26563 , \26564 ,
         \26565 , \26566 , \26567 , \26568 , \26569 , \26570 , \26571 , \26572 , \26573 , \26574 ,
         \26575 , \26576 , \26577 , \26578 , \26579 , \26580 , \26581 , \26582 , \26583 , \26584 ,
         \26585 , \26586 , \26587 , \26588 , \26589 , \26590 , \26591 , \26592 , \26593 , \26594 ,
         \26595 , \26596 , \26597 , \26598 , \26599 , \26600 , \26601 , \26602 , \26603 , \26604 ,
         \26605 , \26606 , \26607 , \26608 , \26609 , \26610 , \26611 , \26612 , \26613 , \26614 ,
         \26615 , \26616 , \26617 , \26618 , \26619 , \26620 , \26621 , \26622 , \26623 , \26624 ,
         \26625 , \26626 , \26627 , \26628 , \26629 , \26630 , \26631 , \26632 , \26633 , \26634 ,
         \26635 , \26636 , \26637 , \26638 , \26639 , \26640 , \26641 , \26642 , \26643 , \26644 ,
         \26645 , \26646 , \26647 , \26648 , \26649 , \26650 , \26651 , \26652 , \26653 , \26654 ,
         \26655 , \26656 , \26657 , \26658 , \26659 , \26660 , \26661 , \26662 , \26663 , \26664 ,
         \26665 , \26666 , \26667 , \26668 , \26669 , \26670 , \26671 , \26672 , \26673 , \26674 ,
         \26675 , \26676 , \26677 , \26678 , \26679 , \26680 , \26681 , \26682 , \26683 , \26684 ,
         \26685 , \26686 , \26687 , \26688 , \26689 , \26690 , \26691 , \26692 , \26693 , \26694 ,
         \26695 , \26696 , \26697 , \26698 , \26699 , \26700 , \26701 , \26702 , \26703 , \26704 ,
         \26705 , \26706 , \26707 , \26708 , \26709 , \26710 , \26711 , \26712 , \26713 , \26714 ,
         \26715 , \26716 , \26717 , \26718 , \26719 , \26720 , \26721 , \26722 , \26723 , \26724 ,
         \26725 , \26726 , \26727 , \26728 , \26729 , \26730 , \26731 , \26732 , \26733 , \26734 ,
         \26735 , \26736 , \26737 , \26738 , \26739 , \26740 , \26741 , \26742 , \26743 , \26744 ,
         \26745 , \26746 , \26747 , \26748 , \26749 , \26750 , \26751 , \26752 , \26753 , \26754 ,
         \26755 , \26756 , \26757 , \26758 , \26759 , \26760 , \26761 , \26762 , \26763 , \26764 ,
         \26765 , \26766 , \26767 , \26768 , \26769 , \26770 , \26771 , \26772 , \26773 , \26774 ,
         \26775 , \26776 , \26777 , \26778 , \26779 , \26780 , \26781 , \26782 , \26783 , \26784 ,
         \26785 , \26786 , \26787 , \26788 , \26789 , \26790 , \26791 , \26792 , \26793 , \26794 ,
         \26795 , \26796 , \26797 , \26798 , \26799 , \26800 , \26801 , \26802 , \26803 , \26804 ,
         \26805 , \26806 , \26807 , \26808 , \26809 , \26810 , \26811 , \26812 , \26813 , \26814 ,
         \26815 , \26816 , \26817 , \26818 , \26819 , \26820 , \26821 , \26822 , \26823 , \26824 ,
         \26825 , \26826 , \26827 , \26828 , \26829 , \26830 , \26831 , \26832 , \26833 , \26834 ,
         \26835 , \26836 , \26837 , \26838 , \26839 , \26840 , \26841 , \26842 , \26843 , \26844 ,
         \26845 , \26846 , \26847 , \26848 , \26849 , \26850 , \26851 , \26852 , \26853 , \26854 ,
         \26855 , \26856 , \26857 , \26858 , \26859 , \26860 , \26861 , \26862 , \26863 , \26864 ,
         \26865 , \26866 , \26867 , \26868 , \26869 , \26870 , \26871 , \26872 , \26873 , \26874 ,
         \26875 , \26876 , \26877 , \26878 , \26879 , \26880 , \26881 , \26882 , \26883 , \26884 ,
         \26885 , \26886 , \26887 , \26888 , \26889 , \26890 , \26891 , \26892 , \26893 , \26894 ,
         \26895 , \26896 , \26897 , \26898 , \26899 , \26900 , \26901 , \26902 , \26903 , \26904 ,
         \26905 , \26906 , \26907 , \26908 , \26909 , \26910 , \26911 , \26912 , \26913 , \26914 ,
         \26915 , \26916 , \26917 , \26918 , \26919 , \26920 , \26921 , \26922 , \26923 , \26924 ,
         \26925 , \26926 , \26927 , \26928 , \26929 , \26930 , \26931 , \26932 , \26933 , \26934 ,
         \26935 , \26936 , \26937 , \26938 , \26939 , \26940 , \26941 , \26942 , \26943 , \26944 ,
         \26945 , \26946 , \26947 , \26948 , \26949 , \26950 , \26951 , \26952 , \26953 , \26954 ,
         \26955 , \26956 , \26957 , \26958 , \26959 , \26960 , \26961 , \26962 , \26963 , \26964 ,
         \26965 , \26966 , \26967 , \26968 , \26969 , \26970 , \26971 , \26972 , \26973 , \26974 ,
         \26975 , \26976 , \26977 , \26978 , \26979 , \26980 , \26981 , \26982 , \26983 , \26984 ,
         \26985 , \26986 , \26987 , \26988 , \26989 , \26990 , \26991 , \26992 , \26993 , \26994 ,
         \26995 , \26996 , \26997 , \26998 , \26999 , \27000 , \27001 , \27002 , \27003 , \27004 ,
         \27005 , \27006 , \27007 , \27008 , \27009 , \27010 , \27011 , \27012 , \27013 , \27014 ,
         \27015 , \27016 , \27017 , \27018 , \27019 , \27020 , \27021 , \27022 , \27023 , \27024 ,
         \27025 , \27026 , \27027 , \27028 , \27029 , \27030 , \27031 , \27032 , \27033 , \27034 ,
         \27035 , \27036 , \27037 , \27038 , \27039 , \27040 , \27041 , \27042 , \27043 , \27044 ,
         \27045 , \27046 , \27047 , \27048 , \27049 , \27050 , \27051 , \27052 , \27053 , \27054 ,
         \27055 , \27056 , \27057 , \27058 , \27059 , \27060 , \27061 , \27062 , \27063 , \27064 ,
         \27065 , \27066 , \27067 , \27068 , \27069 , \27070 , \27071 , \27072 , \27073 , \27074 ,
         \27075 , \27076 , \27077 , \27078 , \27079 , \27080 , \27081 , \27082 , \27083 , \27084 ,
         \27085 , \27086 , \27087 , \27088 , \27089 , \27090 , \27091 , \27092 , \27093 , \27094 ,
         \27095 , \27096 , \27097 , \27098 , \27099 , \27100 , \27101 , \27102 , \27103 , \27104 ,
         \27105 , \27106 , \27107 , \27108 , \27109 , \27110 , \27111 , \27112 , \27113 , \27114 ,
         \27115 , \27116 , \27117 , \27118 , \27119 , \27120 , \27121 , \27122 , \27123 , \27124 ,
         \27125 , \27126 , \27127 , \27128 , \27129 , \27130 , \27131 , \27132 , \27133 , \27134 ,
         \27135 , \27136 , \27137 , \27138 , \27139 , \27140 , \27141 , \27142 , \27143 , \27144 ,
         \27145 , \27146 , \27147 , \27148 , \27149 , \27150 , \27151 , \27152 , \27153 , \27154 ,
         \27155 , \27156 , \27157 , \27158 , \27159 , \27160 , \27161 , \27162 , \27163 , \27164 ,
         \27165 , \27166 , \27167 , \27168 , \27169 , \27170 , \27171 , \27172 , \27173 , \27174 ,
         \27175 , \27176 , \27177 , \27178 , \27179 , \27180 , \27181 , \27182 , \27183 , \27184 ,
         \27185 , \27186 , \27187 , \27188 , \27189 , \27190 , \27191 , \27192 , \27193 , \27194 ,
         \27195 , \27196 , \27197 , \27198 , \27199 , \27200 , \27201 , \27202 , \27203 , \27204 ,
         \27205 , \27206 , \27207 , \27208 , \27209 , \27210 , \27211 , \27212 , \27213 , \27214 ,
         \27215 , \27216 , \27217 , \27218 , \27219 , \27220 , \27221 , \27222 , \27223 , \27224 ,
         \27225 , \27226 , \27227 , \27228 , \27229 , \27230 , \27231 , \27232 , \27233 , \27234 ,
         \27235 , \27236 , \27237 , \27238 , \27239 , \27240 , \27241 , \27242 , \27243 , \27244 ,
         \27245 , \27246 , \27247 , \27248 , \27249 , \27250 , \27251 , \27252 , \27253 , \27254 ,
         \27255 , \27256 , \27257 , \27258 , \27259 , \27260 , \27261 , \27262 , \27263 , \27264 ,
         \27265 , \27266 , \27267 , \27268 , \27269 , \27270 , \27271 , \27272 , \27273 , \27274 ,
         \27275 , \27276 , \27277 , \27278 , \27279 , \27280 , \27281 , \27282 , \27283 , \27284 ,
         \27285 , \27286 , \27287 , \27288 , \27289 , \27290 , \27291 , \27292 , \27293 , \27294 ,
         \27295 , \27296 , \27297 , \27298 , \27299 , \27300 , \27301 , \27302 , \27303 , \27304 ,
         \27305 , \27306 , \27307 , \27308 , \27309 , \27310 , \27311 , \27312 , \27313 , \27314 ,
         \27315 , \27316 , \27317 , \27318 , \27319 , \27320 , \27321 , \27322 , \27323 , \27324 ,
         \27325 , \27326 , \27327 , \27328 , \27329 , \27330 , \27331 , \27332 , \27333 , \27334 ,
         \27335 , \27336 , \27337 , \27338 , \27339 , \27340 , \27341 , \27342 , \27343 , \27344 ,
         \27345 , \27346 , \27347 , \27348 , \27349 , \27350 , \27351 , \27352 , \27353 , \27354 ,
         \27355 , \27356 , \27357 , \27358 , \27359 , \27360 , \27361 , \27362 , \27363 , \27364 ,
         \27365 , \27366 , \27367 , \27368 , \27369 , \27370 , \27371 , \27372 , \27373 , \27374 ,
         \27375 , \27376 , \27377 , \27378 , \27379 , \27380 , \27381 , \27382 , \27383 , \27384 ,
         \27385 , \27386 , \27387 , \27388 , \27389 , \27390 , \27391 , \27392 , \27393 , \27394 ,
         \27395 , \27396 , \27397 , \27398 , \27399 , \27400 , \27401 , \27402 , \27403 , \27404 ,
         \27405 , \27406 , \27407 , \27408 , \27409 , \27410 , \27411 , \27412 , \27413 , \27414 ,
         \27415 , \27416 , \27417 , \27418 , \27419 , \27420 , \27421 , \27422 , \27423 , \27424 ,
         \27425 , \27426 , \27427 , \27428 , \27429 , \27430 , \27431 , \27432 , \27433 , \27434 ,
         \27435 , \27436 , \27437 , \27438 , \27439 , \27440 , \27441 , \27442 , \27443 , \27444 ,
         \27445 , \27446 , \27447 , \27448 , \27449 , \27450 , \27451 , \27452 , \27453 , \27454 ,
         \27455 , \27456 , \27457 , \27458 , \27459 , \27460 , \27461 , \27462 , \27463 , \27464 ,
         \27465 , \27466 , \27467 , \27468 , \27469 , \27470 , \27471 , \27472 , \27473 , \27474 ,
         \27475 , \27476 , \27477 , \27478 , \27479 , \27480 , \27481 , \27482 , \27483 , \27484 ,
         \27485 , \27486 , \27487 , \27488 , \27489 , \27490 , \27491 , \27492 , \27493 , \27494 ,
         \27495 , \27496 , \27497 , \27498 , \27499 , \27500 , \27501 , \27502 , \27503 , \27504 ,
         \27505 , \27506 , \27507 , \27508 , \27509 , \27510 , \27511 , \27512 , \27513 , \27514 ,
         \27515 , \27516 , \27517 , \27518 , \27519 , \27520 , \27521 , \27522 , \27523 , \27524 ,
         \27525 , \27526 , \27527 , \27528 , \27529 , \27530 , \27531 , \27532 , \27533 , \27534 ,
         \27535 , \27536 , \27537 , \27538 , \27539 , \27540 , \27541 , \27542 , \27543 , \27544 ,
         \27545 , \27546 , \27547 , \27548 , \27549 , \27550 , \27551 , \27552 , \27553 , \27554 ,
         \27555 , \27556 , \27557 , \27558 , \27559 , \27560 , \27561 , \27562 , \27563 , \27564 ,
         \27565 , \27566 , \27567 , \27568 , \27569 , \27570 , \27571 , \27572 , \27573 , \27574 ,
         \27575 , \27576 , \27577 , \27578 , \27579 , \27580 , \27581 , \27582 , \27583 , \27584 ,
         \27585 , \27586 , \27587 , \27588 , \27589 , \27590 , \27591 , \27592 , \27593 , \27594 ,
         \27595 , \27596 , \27597 , \27598 , \27599 , \27600 , \27601 , \27602 , \27603 , \27604 ,
         \27605 , \27606 , \27607 , \27608 , \27609 , \27610 , \27611 , \27612 , \27613 , \27614 ,
         \27615 , \27616 , \27617 , \27618 , \27619 , \27620 , \27621 , \27622 , \27623 , \27624 ,
         \27625 , \27626 , \27627 , \27628 , \27629 , \27630 , \27631 , \27632 , \27633 , \27634 ,
         \27635 , \27636 , \27637 , \27638 , \27639 , \27640 , \27641 , \27642 , \27643 , \27644 ,
         \27645 , \27646 , \27647 , \27648 , \27649 , \27650 , \27651 , \27652 , \27653 , \27654 ,
         \27655 , \27656 , \27657 , \27658 , \27659 , \27660 , \27661 , \27662 , \27663 , \27664 ,
         \27665 , \27666 , \27667 , \27668 , \27669 , \27670 , \27671 , \27672 , \27673 , \27674 ,
         \27675 , \27676 , \27677 , \27678 , \27679 , \27680 , \27681 , \27682 , \27683 , \27684 ,
         \27685 , \27686 , \27687 , \27688 , \27689 , \27690 , \27691 , \27692 , \27693 , \27694 ,
         \27695 , \27696 , \27697 , \27698 , \27699 , \27700 , \27701 , \27702 , \27703 , \27704 ,
         \27705 , \27706 , \27707 , \27708 , \27709 , \27710 , \27711 , \27712 , \27713 , \27714 ,
         \27715 , \27716 , \27717 , \27718 , \27719 , \27720 , \27721 , \27722 , \27723 , \27724 ,
         \27725 , \27726 , \27727 , \27728 , \27729 , \27730 , \27731 , \27732 , \27733 , \27734 ,
         \27735 , \27736 , \27737 , \27738 , \27739 , \27740 , \27741 , \27742 , \27743 , \27744 ,
         \27745 , \27746 , \27747 , \27748 , \27749 , \27750 , \27751 , \27752 , \27753 , \27754 ,
         \27755 , \27756 , \27757 , \27758 , \27759 , \27760 , \27761 , \27762 , \27763 , \27764 ,
         \27765 , \27766 , \27767 , \27768 , \27769 , \27770 , \27771 , \27772 , \27773 , \27774 ,
         \27775 , \27776 , \27777 , \27778 , \27779 , \27780 , \27781 , \27782 , \27783 , \27784 ,
         \27785 , \27786 , \27787 , \27788 , \27789 , \27790 , \27791 , \27792 , \27793 , \27794 ,
         \27795 , \27796 , \27797 , \27798 , \27799 , \27800 , \27801 , \27802 , \27803 , \27804 ,
         \27805 , \27806 , \27807 , \27808 , \27809 , \27810 , \27811 , \27812 , \27813 , \27814 ,
         \27815 , \27816 , \27817 , \27818 , \27819 , \27820 , \27821 , \27822 , \27823 , \27824 ,
         \27825 , \27826 , \27827 , \27828 , \27829 , \27830 , \27831 , \27832 , \27833 , \27834 ,
         \27835 , \27836 , \27837 , \27838 , \27839 , \27840 , \27841 , \27842 , \27843 , \27844 ,
         \27845 , \27846 , \27847 , \27848 , \27849 , \27850 , \27851 , \27852 , \27853 , \27854 ,
         \27855 , \27856 , \27857 , \27858 , \27859 , \27860 , \27861 , \27862 , \27863 , \27864 ,
         \27865 , \27866 , \27867 , \27868 , \27869 , \27870 , \27871 , \27872 , \27873 , \27874 ,
         \27875 , \27876 , \27877 , \27878 , \27879 , \27880 , \27881 , \27882 , \27883 , \27884 ,
         \27885 , \27886 , \27887 , \27888 , \27889 , \27890 , \27891 , \27892 , \27893 , \27894 ,
         \27895 , \27896 , \27897 , \27898 , \27899 , \27900 , \27901 , \27902 , \27903 , \27904 ,
         \27905 , \27906 , \27907 , \27908 , \27909 , \27910 , \27911 , \27912 , \27913 , \27914 ,
         \27915 , \27916 , \27917 , \27918 , \27919 , \27920 , \27921 , \27922 , \27923 , \27924 ,
         \27925 , \27926 , \27927 , \27928 , \27929 , \27930 , \27931 , \27932 , \27933 , \27934 ,
         \27935 , \27936 , \27937 , \27938 , \27939 , \27940 , \27941 , \27942 , \27943 , \27944 ,
         \27945 , \27946 , \27947 , \27948 , \27949 , \27950 , \27951 , \27952 , \27953 , \27954 ,
         \27955 , \27956 , \27957 , \27958 , \27959 , \27960 , \27961 , \27962 , \27963 , \27964 ,
         \27965 , \27966 , \27967 , \27968 , \27969 , \27970 , \27971 , \27972 , \27973 , \27974 ,
         \27975 , \27976 , \27977 , \27978 , \27979 , \27980 , \27981 , \27982 , \27983 , \27984 ,
         \27985 , \27986 , \27987 , \27988 , \27989 , \27990 , \27991 , \27992 , \27993 , \27994 ,
         \27995 , \27996 , \27997 , \27998 , \27999 , \28000 , \28001 , \28002 , \28003 , \28004 ,
         \28005 , \28006 , \28007 , \28008 , \28009 , \28010 , \28011 , \28012 , \28013 , \28014 ,
         \28015 , \28016 , \28017 , \28018 , \28019 , \28020 , \28021 , \28022 , \28023 , \28024 ,
         \28025 , \28026 , \28027 , \28028 , \28029 , \28030 , \28031 , \28032 , \28033 , \28034 ,
         \28035 , \28036 , \28037 , \28038 , \28039 , \28040 , \28041 , \28042 , \28043 , \28044 ,
         \28045 , \28046 , \28047 , \28048 , \28049 , \28050 , \28051 , \28052 , \28053 , \28054 ,
         \28055 , \28056 , \28057 , \28058 , \28059 , \28060 , \28061 , \28062 , \28063 , \28064 ,
         \28065 , \28066 , \28067 , \28068 , \28069 , \28070 , \28071 , \28072 , \28073 , \28074 ,
         \28075 , \28076 , \28077 , \28078 , \28079 , \28080 , \28081 , \28082 , \28083 , \28084 ,
         \28085 , \28086 , \28087 , \28088 , \28089 , \28090 , \28091 , \28092 , \28093 , \28094 ,
         \28095 , \28096 , \28097 , \28098 , \28099 , \28100 , \28101 , \28102 , \28103 , \28104 ,
         \28105 , \28106 , \28107 , \28108 , \28109 , \28110 , \28111 , \28112 , \28113 , \28114 ,
         \28115 , \28116 , \28117 , \28118 , \28119 , \28120 , \28121 , \28122 , \28123 , \28124 ,
         \28125 , \28126 , \28127 , \28128 , \28129 , \28130 , \28131 , \28132 , \28133 , \28134 ,
         \28135 , \28136 , \28137 , \28138 , \28139 , \28140 , \28141 , \28142 , \28143 , \28144 ,
         \28145 , \28146 , \28147 , \28148 , \28149 , \28150 , \28151 , \28152 , \28153 , \28154 ,
         \28155 , \28156 , \28157 , \28158 , \28159 , \28160 , \28161 , \28162 , \28163 , \28164 ,
         \28165 , \28166 , \28167 , \28168 , \28169 , \28170 , \28171 , \28172 , \28173 , \28174 ,
         \28175 , \28176 , \28177 , \28178 , \28179 , \28180 , \28181 , \28182 , \28183 , \28184 ,
         \28185 , \28186 , \28187 , \28188 , \28189 , \28190 , \28191 , \28192 , \28193 , \28194 ,
         \28195 , \28196 , \28197 , \28198 , \28199 , \28200 , \28201 , \28202 , \28203 , \28204 ,
         \28205 , \28206 , \28207 , \28208 , \28209 , \28210 , \28211 , \28212 , \28213 , \28214 ,
         \28215 , \28216 , \28217 , \28218 , \28219 , \28220 , \28221 , \28222 , \28223 , \28224 ,
         \28225 , \28226 , \28227 , \28228 , \28229 , \28230 , \28231 , \28232 , \28233 , \28234 ,
         \28235 , \28236 , \28237 , \28238 , \28239 , \28240 , \28241 , \28242 , \28243 , \28244 ,
         \28245 , \28246 , \28247 , \28248 , \28249 , \28250 , \28251 , \28252 , \28253 , \28254 ,
         \28255 , \28256 , \28257 , \28258 , \28259 , \28260 , \28261 , \28262 , \28263 , \28264 ,
         \28265 , \28266 , \28267 , \28268 , \28269 , \28270 , \28271 , \28272 , \28273 , \28274 ,
         \28275 , \28276 , \28277 , \28278 , \28279 , \28280 , \28281 , \28282 , \28283 , \28284 ,
         \28285 , \28286 , \28287 , \28288 , \28289 , \28290 , \28291 , \28292 , \28293 , \28294 ,
         \28295 , \28296 , \28297 , \28298 , \28299 , \28300 , \28301 , \28302 , \28303 , \28304 ,
         \28305 , \28306 , \28307 , \28308 , \28309 , \28310 , \28311 , \28312 , \28313 , \28314 ,
         \28315 , \28316 , \28317 , \28318 , \28319 , \28320 , \28321 , \28322 , \28323 , \28324 ,
         \28325 , \28326 , \28327 , \28328 , \28329 , \28330 , \28331 , \28332 , \28333 , \28334 ,
         \28335 , \28336 , \28337 , \28338 , \28339 , \28340 , \28341 , \28342 , \28343 , \28344 ,
         \28345 , \28346 , \28347 , \28348 , \28349 , \28350 , \28351 , \28352 , \28353 , \28354 ,
         \28355 , \28356 , \28357 , \28358 , \28359 , \28360 , \28361 , \28362 , \28363 , \28364 ,
         \28365 , \28366 , \28367 , \28368 , \28369 , \28370 , \28371 , \28372 , \28373 , \28374 ,
         \28375 , \28376 , \28377 , \28378 , \28379 , \28380 , \28381 , \28382 , \28383 , \28384 ,
         \28385 , \28386 , \28387 , \28388 , \28389 , \28390 , \28391 , \28392 , \28393 , \28394 ,
         \28395 , \28396 , \28397 , \28398 , \28399 , \28400 , \28401 , \28402 , \28403 , \28404 ,
         \28405 , \28406 , \28407 , \28408 , \28409 , \28410 , \28411 , \28412 , \28413 , \28414 ,
         \28415 , \28416 , \28417 , \28418 , \28419 , \28420 , \28421 , \28422 , \28423 , \28424 ,
         \28425 , \28426 , \28427 , \28428 , \28429 , \28430 , \28431 , \28432 , \28433 , \28434 ,
         \28435 , \28436 , \28437 , \28438 , \28439 , \28440 , \28441 , \28442 , \28443 , \28444 ,
         \28445 , \28446 , \28447 , \28448 , \28449 , \28450 , \28451 , \28452 , \28453 , \28454 ,
         \28455 , \28456 , \28457 , \28458 , \28459 , \28460 , \28461 , \28462 , \28463 , \28464 ,
         \28465 , \28466 , \28467 , \28468 , \28469 , \28470 , \28471 , \28472 , \28473 , \28474 ,
         \28475 , \28476 , \28477 , \28478 , \28479 , \28480 , \28481 , \28482 , \28483 , \28484 ,
         \28485 , \28486 , \28487 , \28488 , \28489 , \28490 , \28491 , \28492 , \28493 , \28494 ,
         \28495 , \28496 , \28497 , \28498 , \28499 , \28500 , \28501 , \28502 , \28503 , \28504 ,
         \28505 , \28506 , \28507 , \28508 , \28509 , \28510 , \28511 , \28512 , \28513 , \28514 ,
         \28515 , \28516 , \28517 , \28518 , \28519 , \28520 , \28521 , \28522 , \28523 , \28524 ,
         \28525 , \28526 , \28527 , \28528 , \28529 , \28530 , \28531 , \28532 , \28533 , \28534 ,
         \28535 , \28536 , \28537 , \28538 , \28539 , \28540 , \28541 , \28542 , \28543 , \28544 ,
         \28545 , \28546 , \28547 , \28548 , \28549 , \28550 , \28551 , \28552 , \28553 , \28554 ,
         \28555 , \28556 , \28557 , \28558 , \28559 , \28560 , \28561 , \28562 , \28563 , \28564 ,
         \28565 , \28566 , \28567 , \28568 , \28569 , \28570 , \28571 , \28572 , \28573 , \28574 ,
         \28575 , \28576 , \28577 , \28578 , \28579 , \28580 , \28581 , \28582 , \28583 , \28584 ,
         \28585 , \28586 , \28587 , \28588 , \28589 , \28590 , \28591 , \28592 , \28593 , \28594 ,
         \28595 , \28596 , \28597 , \28598 , \28599 , \28600 , \28601 , \28602 , \28603 , \28604 ,
         \28605 , \28606 , \28607 , \28608 , \28609 , \28610 , \28611 , \28612 , \28613 , \28614 ,
         \28615 , \28616 , \28617 , \28618 , \28619 , \28620 , \28621 , \28622 , \28623 , \28624 ,
         \28625 , \28626 , \28627 , \28628 , \28629 , \28630 , \28631 , \28632 , \28633 , \28634 ,
         \28635 , \28636 , \28637 , \28638 , \28639 , \28640 , \28641 , \28642 , \28643 , \28644 ,
         \28645 , \28646 , \28647 , \28648 , \28649 , \28650 , \28651 , \28652 , \28653 , \28654 ,
         \28655 , \28656 , \28657 , \28658 , \28659 , \28660 , \28661 , \28662 , \28663 , \28664 ,
         \28665 , \28666 , \28667 , \28668 , \28669 , \28670 , \28671 , \28672 , \28673 , \28674 ,
         \28675 , \28676 , \28677 , \28678 , \28679 , \28680 , \28681 , \28682 , \28683 , \28684 ,
         \28685 , \28686 , \28687 , \28688 , \28689 , \28690 , \28691 , \28692 , \28693 , \28694 ,
         \28695 , \28696 , \28697 , \28698 , \28699 , \28700 , \28701 , \28702 , \28703 , \28704 ,
         \28705 , \28706 , \28707 , \28708 , \28709 , \28710 , \28711 , \28712 , \28713 , \28714 ,
         \28715 , \28716 , \28717 , \28718 , \28719 , \28720 , \28721 , \28722 , \28723 , \28724 ,
         \28725 , \28726 , \28727 , \28728 , \28729 , \28730 , \28731 , \28732 , \28733 , \28734 ,
         \28735 , \28736 , \28737 , \28738 , \28739 , \28740 , \28741 , \28742 , \28743 , \28744 ,
         \28745 , \28746 , \28747 , \28748 , \28749 , \28750 , \28751 , \28752 , \28753 , \28754 ,
         \28755 , \28756 , \28757 , \28758 , \28759 , \28760 , \28761 , \28762 , \28763 , \28764 ,
         \28765 , \28766 , \28767 , \28768 , \28769 , \28770 , \28771 , \28772 , \28773 , \28774 ,
         \28775 , \28776 , \28777 , \28778 , \28779 , \28780 , \28781 , \28782 , \28783 , \28784 ,
         \28785 , \28786 , \28787 , \28788 , \28789 , \28790 , \28791 , \28792 , \28793 , \28794 ,
         \28795 , \28796 , \28797 , \28798 , \28799 , \28800 , \28801 , \28802 , \28803 , \28804 ,
         \28805 , \28806 , \28807 , \28808 , \28809 , \28810 , \28811 , \28812 , \28813 , \28814 ,
         \28815 , \28816 , \28817 , \28818 , \28819 , \28820 , \28821 , \28822 , \28823 , \28824 ,
         \28825 , \28826 , \28827 , \28828 , \28829 , \28830 , \28831 , \28832 , \28833 , \28834 ,
         \28835 , \28836 , \28837 , \28838 , \28839 , \28840 , \28841 , \28842 , \28843 , \28844 ,
         \28845 , \28846 , \28847 , \28848 , \28849 , \28850 , \28851 , \28852 , \28853 , \28854 ,
         \28855 , \28856 , \28857 , \28858 , \28859 , \28860 , \28861 , \28862 , \28863 , \28864 ,
         \28865 , \28866 , \28867 , \28868 , \28869 , \28870 , \28871 , \28872 , \28873 , \28874 ,
         \28875 , \28876 , \28877 , \28878 , \28879 , \28880 , \28881 , \28882 , \28883 , \28884 ,
         \28885 , \28886 , \28887 , \28888 , \28889 , \28890 , \28891 , \28892 , \28893 , \28894 ,
         \28895 , \28896 , \28897 , \28898 , \28899 , \28900 , \28901 , \28902 , \28903 , \28904 ,
         \28905 , \28906 , \28907 , \28908 , \28909 , \28910 , \28911 , \28912 , \28913 , \28914 ,
         \28915 , \28916 , \28917 , \28918 , \28919 , \28920 , \28921 , \28922 , \28923 , \28924 ,
         \28925 , \28926 , \28927 , \28928 , \28929 , \28930 , \28931 , \28932 , \28933 , \28934 ,
         \28935 , \28936 , \28937 , \28938 , \28939 , \28940 , \28941 , \28942 , \28943 , \28944 ,
         \28945 , \28946 , \28947 , \28948 , \28949 , \28950 , \28951 , \28952 , \28953 , \28954 ,
         \28955 , \28956 , \28957 , \28958 , \28959 , \28960 , \28961 , \28962 , \28963 , \28964 ,
         \28965 , \28966 , \28967 , \28968 , \28969 , \28970 , \28971 , \28972 , \28973 , \28974 ,
         \28975 , \28976 , \28977 , \28978 , \28979 , \28980 , \28981 , \28982 , \28983 , \28984 ,
         \28985 , \28986 , \28987 , \28988 , \28989 , \28990 , \28991 , \28992 , \28993 , \28994 ,
         \28995 , \28996 , \28997 , \28998 , \28999 , \29000 , \29001 , \29002 , \29003 , \29004 ,
         \29005 , \29006 , \29007 , \29008 , \29009 , \29010 , \29011 , \29012 , \29013 , \29014 ,
         \29015 , \29016 , \29017 , \29018 , \29019 , \29020 , \29021 , \29022 , \29023 , \29024 ,
         \29025 , \29026 , \29027 , \29028 , \29029 , \29030 , \29031 , \29032 , \29033 , \29034 ,
         \29035 , \29036 , \29037 , \29038 , \29039 , \29040 , \29041 , \29042 , \29043 , \29044 ,
         \29045 , \29046 , \29047 , \29048 , \29049 , \29050 , \29051 , \29052 , \29053 , \29054 ,
         \29055 , \29056 , \29057 , \29058 , \29059 , \29060 , \29061 , \29062 , \29063 , \29064 ,
         \29065 , \29066 , \29067 , \29068 , \29069 , \29070 , \29071 , \29072 , \29073 , \29074 ,
         \29075 , \29076 , \29077 , \29078 , \29079 , \29080 , \29081 , \29082 , \29083 , \29084 ,
         \29085 , \29086 , \29087 , \29088 , \29089 , \29090 , \29091 , \29092 , \29093 , \29094 ,
         \29095 , \29096 , \29097 , \29098 , \29099 , \29100 , \29101 , \29102 , \29103 , \29104 ,
         \29105 , \29106 , \29107 , \29108 , \29109 , \29110 , \29111 , \29112 , \29113 , \29114 ,
         \29115 , \29116 , \29117 , \29118 , \29119 , \29120 , \29121 , \29122 , \29123 , \29124 ,
         \29125 , \29126 , \29127 , \29128 , \29129 , \29130 , \29131 , \29132 , \29133 , \29134 ,
         \29135 , \29136 , \29137 , \29138 , \29139 , \29140 , \29141 , \29142 , \29143 , \29144 ,
         \29145 , \29146 , \29147 , \29148 , \29149 , \29150 , \29151 , \29152 , \29153 , \29154 ,
         \29155 , \29156 , \29157 , \29158 , \29159 , \29160 , \29161 , \29162 , \29163 , \29164 ,
         \29165 , \29166 , \29167 , \29168 , \29169 , \29170 , \29171 , \29172 , \29173 , \29174 ,
         \29175 , \29176 , \29177 , \29178 , \29179 , \29180 , \29181 , \29182 , \29183 , \29184 ,
         \29185 , \29186 , \29187 , \29188 , \29189 , \29190 , \29191 , \29192 , \29193 , \29194 ,
         \29195 , \29196 , \29197 , \29198 , \29199 , \29200 , \29201 , \29202 , \29203 , \29204 ,
         \29205 , \29206 , \29207 , \29208 , \29209 , \29210 , \29211 , \29212 , \29213 , \29214 ,
         \29215 , \29216 , \29217 , \29218 , \29219 , \29220 , \29221 , \29222 , \29223 , \29224 ,
         \29225 , \29226 , \29227 , \29228 , \29229 , \29230 , \29231 , \29232 , \29233 , \29234 ,
         \29235 , \29236 , \29237 , \29238 , \29239 , \29240 , \29241 , \29242 , \29243 , \29244 ,
         \29245 , \29246 , \29247 , \29248 , \29249 , \29250 , \29251 , \29252 , \29253 , \29254 ,
         \29255 , \29256 , \29257 , \29258 , \29259 , \29260 , \29261 , \29262 , \29263 , \29264 ,
         \29265 , \29266 , \29267 , \29268 , \29269 , \29270 , \29271 , \29272 , \29273 , \29274 ,
         \29275 , \29276 , \29277 , \29278 , \29279 , \29280 , \29281 , \29282 , \29283 , \29284 ,
         \29285 , \29286 , \29287 , \29288 , \29289 , \29290 , \29291 , \29292 , \29293 , \29294 ,
         \29295 , \29296 , \29297 , \29298 , \29299 , \29300 , \29301 , \29302 , \29303 , \29304 ,
         \29305 , \29306 , \29307 , \29308 , \29309 , \29310 , \29311 , \29312 , \29313 , \29314 ,
         \29315 , \29316 , \29317 , \29318 , \29319 , \29320 , \29321 , \29322 , \29323 , \29324 ,
         \29325 , \29326 , \29327 , \29328 , \29329 , \29330 , \29331 , \29332 , \29333 , \29334 ,
         \29335 , \29336 , \29337 , \29338 , \29339 , \29340 , \29341 , \29342 , \29343 , \29344 ,
         \29345 , \29346 , \29347 , \29348 , \29349 , \29350 , \29351 , \29352 , \29353 , \29354 ,
         \29355 , \29356 , \29357 , \29358 , \29359 , \29360 , \29361 , \29362 , \29363 , \29364 ,
         \29365 , \29366 , \29367 , \29368 , \29369 , \29370 , \29371 , \29372 , \29373 , \29374 ,
         \29375 , \29376 , \29377 , \29378 , \29379 , \29380 , \29381 , \29382 , \29383 , \29384 ,
         \29385 , \29386 , \29387 , \29388 , \29389 , \29390 , \29391 , \29392 , \29393 , \29394 ,
         \29395 , \29396 , \29397 , \29398 , \29399 , \29400 , \29401 , \29402 , \29403 , \29404 ,
         \29405 , \29406 , \29407 , \29408 , \29409 , \29410 , \29411 , \29412 , \29413 , \29414 ,
         \29415 , \29416 , \29417 , \29418 , \29419 , \29420 , \29421 , \29422 , \29423 , \29424 ,
         \29425 , \29426 , \29427 , \29428 , \29429 , \29430 , \29431 , \29432 , \29433 , \29434 ,
         \29435 , \29436 , \29437 , \29438 , \29439 , \29440 , \29441 , \29442 , \29443 , \29444 ,
         \29445 , \29446 , \29447 , \29448 , \29449 , \29450 , \29451 , \29452 , \29453 , \29454 ,
         \29455 , \29456 , \29457 , \29458 , \29459 , \29460 , \29461 , \29462 , \29463 , \29464 ,
         \29465 , \29466 , \29467 , \29468 , \29469 , \29470 , \29471 , \29472 , \29473 , \29474 ,
         \29475 , \29476 , \29477 , \29478 , \29479 , \29480 , \29481 , \29482 , \29483 , \29484 ,
         \29485 , \29486 , \29487 , \29488 , \29489 , \29490 , \29491 , \29492 , \29493 , \29494 ,
         \29495 , \29496 , \29497 , \29498 , \29499 , \29500 , \29501 , \29502 , \29503 , \29504 ,
         \29505 , \29506 , \29507 , \29508 , \29509 , \29510 , \29511 , \29512 , \29513 , \29514 ,
         \29515 , \29516 , \29517 , \29518 , \29519 , \29520 , \29521 , \29522 , \29523 , \29524 ,
         \29525 , \29526 , \29527 , \29528 , \29529 , \29530 , \29531 , \29532 , \29533 , \29534 ,
         \29535 , \29536 , \29537 , \29538 , \29539 , \29540 , \29541 , \29542 , \29543 , \29544 ,
         \29545 , \29546 , \29547 , \29548 , \29549 , \29550 , \29551 , \29552 , \29553 , \29554 ,
         \29555 , \29556 , \29557 , \29558 , \29559 , \29560 , \29561 , \29562 , \29563 , \29564 ,
         \29565 , \29566 , \29567 , \29568 , \29569 , \29570 , \29571 , \29572 , \29573 , \29574 ,
         \29575 , \29576 , \29577 , \29578 , \29579 , \29580 , \29581 , \29582 , \29583 , \29584 ,
         \29585 , \29586 , \29587 , \29588 , \29589 , \29590 , \29591 , \29592 , \29593 , \29594 ,
         \29595 , \29596 , \29597 , \29598 , \29599 , \29600 , \29601 , \29602 , \29603 , \29604 ,
         \29605 , \29606 , \29607 , \29608 , \29609 , \29610 , \29611 , \29612 , \29613 , \29614 ,
         \29615 , \29616 , \29617 , \29618 , \29619 , \29620 , \29621 , \29622 , \29623 , \29624 ,
         \29625 , \29626 , \29627 , \29628 , \29629 , \29630 , \29631 , \29632 , \29633 , \29634 ,
         \29635 , \29636 , \29637 , \29638 , \29639 , \29640 , \29641 , \29642 , \29643 , \29644 ,
         \29645 , \29646 , \29647 , \29648 , \29649 , \29650 , \29651 , \29652 , \29653 , \29654 ,
         \29655 , \29656 , \29657 , \29658 , \29659 , \29660 , \29661 , \29662 , \29663 , \29664 ,
         \29665 , \29666 , \29667 , \29668 , \29669 , \29670 , \29671 , \29672 , \29673 , \29674 ,
         \29675 , \29676 , \29677 , \29678 , \29679 , \29680 , \29681 , \29682 , \29683 , \29684 ,
         \29685 , \29686 , \29687 , \29688 , \29689 , \29690 , \29691 , \29692 , \29693 , \29694 ,
         \29695 , \29696 , \29697 , \29698 , \29699 , \29700 , \29701 , \29702 , \29703 , \29704 ,
         \29705 , \29706 , \29707 , \29708 , \29709 , \29710 , \29711 , \29712 , \29713 , \29714 ,
         \29715 , \29716 , \29717 , \29718 , \29719 , \29720 , \29721 , \29722 , \29723 , \29724 ,
         \29725 , \29726 , \29727 , \29728 , \29729 , \29730 , \29731 , \29732 , \29733 , \29734 ,
         \29735 , \29736 , \29737 , \29738 , \29739 , \29740 , \29741 , \29742 , \29743 , \29744 ,
         \29745 , \29746 , \29747 , \29748 , \29749 , \29750 , \29751 , \29752 , \29753 , \29754 ,
         \29755 , \29756 , \29757 , \29758 , \29759 , \29760 , \29761 , \29762 , \29763 , \29764 ,
         \29765 , \29766 , \29767 , \29768 , \29769 , \29770 , \29771 , \29772 , \29773 , \29774 ,
         \29775 , \29776 , \29777 , \29778 , \29779 , \29780 , \29781 , \29782 , \29783 , \29784 ,
         \29785 , \29786 , \29787 , \29788 , \29789 , \29790 , \29791 , \29792 , \29793 , \29794 ,
         \29795 , \29796 , \29797 , \29798 , \29799 , \29800 , \29801 , \29802 , \29803 , \29804 ,
         \29805 , \29806 , \29807 , \29808 , \29809 , \29810 , \29811 , \29812 , \29813 , \29814 ,
         \29815 , \29816 , \29817 , \29818 , \29819 , \29820 , \29821 , \29822 , \29823 , \29824 ,
         \29825 , \29826 , \29827 , \29828 , \29829 , \29830 , \29831 , \29832 , \29833 , \29834 ,
         \29835 , \29836 , \29837 , \29838 , \29839 , \29840 , \29841 , \29842 , \29843 , \29844 ,
         \29845 , \29846 , \29847 , \29848 , \29849 , \29850 , \29851 , \29852 , \29853 , \29854 ,
         \29855 , \29856 , \29857 , \29858 , \29859 , \29860 , \29861 , \29862 , \29863 , \29864 ,
         \29865 , \29866 , \29867 , \29868 , \29869 , \29870 , \29871 , \29872 , \29873 , \29874 ,
         \29875 , \29876 , \29877 , \29878 , \29879 , \29880 , \29881 , \29882 , \29883 , \29884 ,
         \29885 , \29886 , \29887 , \29888 , \29889 , \29890 , \29891 , \29892 , \29893 , \29894 ,
         \29895 , \29896 , \29897 , \29898 , \29899 , \29900 , \29901 , \29902 , \29903 , \29904 ,
         \29905 , \29906 , \29907 , \29908 , \29909 , \29910 , \29911 , \29912 , \29913 , \29914 ,
         \29915 , \29916 , \29917 , \29918 , \29919 , \29920 , \29921 , \29922 , \29923 , \29924 ,
         \29925 , \29926 , \29927 , \29928 , \29929 , \29930 , \29931 , \29932 , \29933 , \29934 ,
         \29935 , \29936 , \29937 , \29938 , \29939 , \29940 , \29941 , \29942 , \29943 , \29944 ,
         \29945 , \29946 , \29947 , \29948 , \29949 , \29950 , \29951 , \29952 , \29953 , \29954 ,
         \29955 , \29956 , \29957 , \29958 , \29959 , \29960 , \29961 , \29962 , \29963 , \29964 ,
         \29965 , \29966 , \29967 , \29968 , \29969 , \29970 , \29971 , \29972 , \29973 , \29974 ,
         \29975 , \29976 , \29977 , \29978 , \29979 , \29980 , \29981 , \29982 , \29983 , \29984 ,
         \29985 , \29986 , \29987 , \29988 , \29989 , \29990 , \29991 , \29992 , \29993 , \29994 ,
         \29995 , \29996 , \29997 , \29998 , \29999 , \30000 , \30001 , \30002 , \30003 , \30004 ,
         \30005 , \30006 , \30007 , \30008 , \30009 , \30010 , \30011 , \30012 , \30013 , \30014 ,
         \30015 , \30016 , \30017 , \30018 , \30019 , \30020 , \30021 , \30022 , \30023 , \30024 ,
         \30025 , \30026 , \30027 , \30028 , \30029 , \30030 , \30031 , \30032 , \30033 , \30034 ,
         \30035 , \30036 , \30037 , \30038 , \30039 , \30040 , \30041 , \30042 , \30043 , \30044 ,
         \30045 , \30046 , \30047 , \30048 , \30049 , \30050 , \30051 , \30052 , \30053 , \30054 ,
         \30055 , \30056 , \30057 , \30058 , \30059 , \30060 , \30061 , \30062 , \30063 , \30064 ,
         \30065 , \30066 , \30067 , \30068 , \30069 , \30070 , \30071 , \30072 , \30073 , \30074 ,
         \30075 , \30076 , \30077 , \30078 , \30079 , \30080 , \30081 , \30082 , \30083 , \30084 ,
         \30085 , \30086 , \30087 , \30088 , \30089 , \30090 , \30091 , \30092 , \30093 , \30094 ,
         \30095 , \30096 , \30097 , \30098 , \30099 , \30100 , \30101 , \30102 , \30103 , \30104 ,
         \30105 , \30106 , \30107 , \30108 , \30109 , \30110 , \30111 , \30112 , \30113 , \30114 ,
         \30115 , \30116 , \30117 , \30118 , \30119 , \30120 , \30121 , \30122 , \30123 , \30124 ,
         \30125 , \30126 , \30127 , \30128 , \30129 , \30130 , \30131 , \30132 , \30133 , \30134 ,
         \30135 , \30136 , \30137 , \30138 , \30139 , \30140 , \30141 , \30142 , \30143 , \30144 ,
         \30145 , \30146 , \30147 , \30148 , \30149 , \30150 , \30151 , \30152 , \30153 , \30154 ,
         \30155 , \30156 , \30157 , \30158 , \30159 , \30160 , \30161 , \30162 , \30163 , \30164 ,
         \30165 , \30166 , \30167 , \30168 , \30169 , \30170 , \30171 , \30172 , \30173 , \30174 ,
         \30175 , \30176 , \30177 , \30178 , \30179 , \30180 , \30181 , \30182 , \30183 , \30184 ,
         \30185 , \30186 , \30187 , \30188 , \30189 , \30190 , \30191 , \30192 , \30193 , \30194 ,
         \30195 , \30196 , \30197 , \30198 , \30199 , \30200 , \30201 , \30202 , \30203 , \30204 ,
         \30205 , \30206 , \30207 , \30208 , \30209 , \30210 , \30211 , \30212 , \30213 , \30214 ,
         \30215 , \30216 , \30217 , \30218 , \30219 , \30220 , \30221 , \30222 , \30223 , \30224 ,
         \30225 , \30226 , \30227 , \30228 , \30229 , \30230 , \30231 , \30232 , \30233 , \30234 ,
         \30235 , \30236 , \30237 , \30238 , \30239 , \30240 , \30241 , \30242 , \30243 , \30244 ,
         \30245 , \30246 , \30247 , \30248 , \30249 , \30250 , \30251 , \30252 , \30253 , \30254 ,
         \30255 , \30256 , \30257 , \30258 , \30259 , \30260 , \30261 , \30262 , \30263 , \30264 ,
         \30265 , \30266 , \30267 , \30268 , \30269 , \30270 , \30271 , \30272 , \30273 , \30274 ,
         \30275 , \30276 , \30277 , \30278 , \30279 , \30280 , \30281 , \30282 , \30283 , \30284 ,
         \30285 , \30286 , \30287 , \30288 , \30289 , \30290 , \30291 , \30292 , \30293 , \30294 ,
         \30295 , \30296 , \30297 , \30298 , \30299 , \30300 , \30301 , \30302 , \30303 , \30304 ,
         \30305 , \30306 , \30307 , \30308 , \30309 , \30310 , \30311 , \30312 , \30313 , \30314 ,
         \30315 , \30316 , \30317 , \30318 , \30319 , \30320 , \30321 , \30322 , \30323 , \30324 ,
         \30325 , \30326 , \30327 , \30328 , \30329 , \30330 , \30331 , \30332 , \30333 , \30334 ,
         \30335 , \30336 , \30337 , \30338 , \30339 , \30340 , \30341 , \30342 , \30343 , \30344 ,
         \30345 , \30346 , \30347 , \30348 , \30349 , \30350 , \30351 , \30352 , \30353 , \30354 ,
         \30355 , \30356 , \30357 , \30358 , \30359 , \30360 , \30361 , \30362 , \30363 , \30364 ,
         \30365 , \30366 , \30367 , \30368 , \30369 , \30370 , \30371 , \30372 , \30373 , \30374 ,
         \30375 , \30376 , \30377 , \30378 , \30379 , \30380 , \30381 , \30382 , \30383 , \30384 ,
         \30385 , \30386 , \30387 , \30388 , \30389 , \30390 , \30391 , \30392 , \30393 , \30394 ,
         \30395 , \30396 , \30397 , \30398 , \30399 , \30400 , \30401 , \30402 , \30403 , \30404 ,
         \30405 , \30406 , \30407 , \30408 , \30409 , \30410 , \30411 , \30412 , \30413 , \30414 ,
         \30415 , \30416 , \30417 , \30418 , \30419 , \30420 , \30421 , \30422 , \30423 , \30424 ,
         \30425 , \30426 , \30427 , \30428 , \30429 , \30430 , \30431 , \30432 , \30433 , \30434 ,
         \30435 , \30436 , \30437 , \30438 , \30439 , \30440 , \30441 , \30442 , \30443 , \30444 ,
         \30445 , \30446 , \30447 , \30448 , \30449 , \30450 , \30451 , \30452 , \30453 , \30454 ,
         \30455 , \30456 , \30457 , \30458 , \30459 , \30460 , \30461 , \30462 , \30463 , \30464 ,
         \30465 , \30466 , \30467 , \30468 , \30469 , \30470 , \30471 , \30472 , \30473 , \30474 ,
         \30475 , \30476 , \30477 , \30478 , \30479 , \30480 , \30481 , \30482 , \30483 , \30484 ,
         \30485 , \30486 , \30487 , \30488 , \30489 , \30490 , \30491 , \30492 , \30493 , \30494 ,
         \30495 , \30496 , \30497 , \30498 , \30499 , \30500 , \30501 , \30502 , \30503 , \30504 ,
         \30505 , \30506 , \30507 , \30508 , \30509 , \30510 , \30511 , \30512 , \30513 , \30514 ,
         \30515 , \30516 , \30517 , \30518 , \30519 , \30520 , \30521 , \30522 , \30523 , \30524 ,
         \30525 , \30526 , \30527 , \30528 , \30529 , \30530 , \30531 , \30532 , \30533 , \30534 ,
         \30535 , \30536 , \30537 , \30538 , \30539 , \30540 , \30541 , \30542 , \30543 , \30544 ,
         \30545 , \30546 , \30547 , \30548 , \30549 , \30550 , \30551 , \30552 , \30553 , \30554 ,
         \30555 , \30556 , \30557 , \30558 , \30559 , \30560 , \30561 , \30562 , \30563 , \30564 ,
         \30565 , \30566 , \30567 , \30568 , \30569 , \30570 , \30571 , \30572 , \30573 , \30574 ,
         \30575 , \30576 , \30577 , \30578 , \30579 , \30580 , \30581 , \30582 , \30583 , \30584 ,
         \30585 , \30586 , \30587 , \30588 , \30589 , \30590 , \30591 , \30592 , \30593 , \30594 ,
         \30595 , \30596 , \30597 , \30598 , \30599 , \30600 , \30601 , \30602 , \30603 , \30604 ,
         \30605 , \30606 , \30607 , \30608 , \30609 , \30610 , \30611 , \30612 , \30613 , \30614 ,
         \30615 , \30616 , \30617 , \30618 , \30619 , \30620 , \30621 , \30622 , \30623 , \30624 ,
         \30625 , \30626 , \30627 , \30628 , \30629 , \30630 , \30631 , \30632 , \30633 , \30634 ,
         \30635 , \30636 , \30637 , \30638 , \30639 , \30640 , \30641 , \30642 , \30643 , \30644 ,
         \30645 , \30646 , \30647 , \30648 , \30649 , \30650 , \30651 , \30652 , \30653 , \30654 ,
         \30655 , \30656 , \30657 , \30658 , \30659 , \30660 , \30661 , \30662 , \30663 , \30664 ,
         \30665 , \30666 , \30667 , \30668 , \30669 , \30670 , \30671 , \30672 , \30673 , \30674 ,
         \30675 , \30676 , \30677 , \30678 , \30679 , \30680 , \30681 , \30682 , \30683 , \30684 ,
         \30685 , \30686 , \30687 , \30688 , \30689 , \30690 , \30691 , \30692 , \30693 , \30694 ,
         \30695 , \30696 , \30697 , \30698 , \30699 , \30700 , \30701 , \30702 , \30703 , \30704 ,
         \30705 , \30706 , \30707 , \30708 , \30709 , \30710 , \30711 , \30712 , \30713 , \30714 ,
         \30715 , \30716 , \30717 , \30718 , \30719 , \30720 , \30721 , \30722 , \30723 , \30724 ,
         \30725 , \30726 , \30727 , \30728 , \30729 , \30730 , \30731 , \30732 , \30733 , \30734 ,
         \30735 , \30736 , \30737 , \30738 , \30739 , \30740 , \30741 , \30742 , \30743 , \30744 ,
         \30745 , \30746 , \30747 , \30748 , \30749 , \30750 , \30751 , \30752 , \30753 , \30754 ,
         \30755 , \30756 , \30757 , \30758 , \30759 , \30760 , \30761 , \30762 , \30763 , \30764 ,
         \30765 , \30766 , \30767 , \30768 , \30769 , \30770 , \30771 , \30772 , \30773 , \30774 ,
         \30775 , \30776 , \30777 , \30778 , \30779 , \30780 , \30781 , \30782 , \30783 , \30784 ,
         \30785 , \30786 , \30787 , \30788 , \30789 , \30790 , \30791 , \30792 , \30793 , \30794 ,
         \30795 , \30796 , \30797 , \30798 , \30799 , \30800 , \30801 , \30802 , \30803 , \30804 ,
         \30805 , \30806 , \30807 , \30808 , \30809 , \30810 , \30811 , \30812 , \30813 , \30814 ,
         \30815 , \30816 , \30817 , \30818 , \30819 , \30820 , \30821 , \30822 , \30823 , \30824 ,
         \30825 , \30826 , \30827 , \30828 , \30829 , \30830 , \30831 , \30832 , \30833 , \30834 ,
         \30835 , \30836 , \30837 , \30838 , \30839 , \30840 , \30841 , \30842 , \30843 , \30844 ,
         \30845 , \30846 , \30847 , \30848 , \30849 , \30850 , \30851 , \30852 , \30853 , \30854 ,
         \30855 , \30856 , \30857 , \30858 , \30859 , \30860 , \30861 , \30862 , \30863 , \30864 ,
         \30865 , \30866 , \30867 , \30868 , \30869 , \30870 , \30871 , \30872 , \30873 , \30874 ,
         \30875 , \30876 , \30877 , \30878 , \30879 , \30880 , \30881 , \30882 , \30883 , \30884 ,
         \30885 , \30886 , \30887 , \30888 , \30889 , \30890 , \30891 , \30892 , \30893 , \30894 ,
         \30895 , \30896 , \30897 , \30898 , \30899 , \30900 , \30901 , \30902 , \30903 , \30904 ,
         \30905 , \30906 , \30907 , \30908 , \30909 , \30910 , \30911 , \30912 , \30913 , \30914 ,
         \30915 , \30916 , \30917 , \30918 , \30919 , \30920 , \30921 , \30922 , \30923 , \30924 ,
         \30925 , \30926 , \30927 , \30928 , \30929 , \30930 , \30931 , \30932 , \30933 , \30934 ,
         \30935 , \30936 , \30937 , \30938 , \30939 , \30940 , \30941 , \30942 , \30943 , \30944 ,
         \30945 , \30946 , \30947 , \30948 , \30949 , \30950 , \30951 , \30952 , \30953 , \30954 ,
         \30955 , \30956 , \30957 , \30958 , \30959 , \30960 , \30961 , \30962 , \30963 , \30964 ,
         \30965 , \30966 , \30967 , \30968 , \30969 , \30970 , \30971 , \30972 , \30973 , \30974 ,
         \30975 , \30976 , \30977 , \30978 , \30979 , \30980 , \30981 , \30982 , \30983 , \30984 ,
         \30985 , \30986 , \30987 , \30988 , \30989 , \30990 , \30991 , \30992 , \30993 , \30994 ,
         \30995 , \30996 , \30997 , \30998 , \30999 , \31000 , \31001 , \31002 , \31003 , \31004 ,
         \31005 , \31006 , \31007 , \31008 , \31009 , \31010 , \31011 , \31012 , \31013 , \31014 ,
         \31015 , \31016 , \31017 , \31018 , \31019 , \31020 , \31021 , \31022 , \31023 , \31024 ,
         \31025 , \31026 , \31027 , \31028 , \31029 , \31030 , \31031 , \31032 , \31033 , \31034 ,
         \31035 , \31036 , \31037 , \31038 , \31039 , \31040 , \31041 , \31042 , \31043 , \31044 ,
         \31045 , \31046 , \31047 , \31048 , \31049 , \31050 , \31051 , \31052 , \31053 , \31054 ,
         \31055 , \31056 , \31057 , \31058 , \31059 , \31060 , \31061 , \31062 , \31063 , \31064 ,
         \31065 , \31066 , \31067 , \31068 , \31069 , \31070 , \31071 , \31072 , \31073 , \31074 ,
         \31075 , \31076 , \31077 , \31078 , \31079 , \31080 , \31081 , \31082 , \31083 , \31084 ,
         \31085 , \31086 , \31087 , \31088 , \31089 , \31090 , \31091 , \31092 , \31093 , \31094 ,
         \31095 , \31096 , \31097 , \31098 , \31099 , \31100 , \31101 , \31102 , \31103 , \31104 ,
         \31105 , \31106 , \31107 , \31108 , \31109 , \31110 , \31111 , \31112 , \31113 , \31114 ,
         \31115 , \31116 , \31117 , \31118 , \31119 , \31120 , \31121 , \31122 , \31123 , \31124 ,
         \31125 , \31126 , \31127 , \31128 , \31129 , \31130 , \31131 , \31132 , \31133 , \31134 ,
         \31135 , \31136 , \31137 , \31138 , \31139 , \31140 , \31141 , \31142 , \31143 , \31144 ,
         \31145 , \31146 , \31147 , \31148 , \31149 , \31150 , \31151 , \31152 , \31153 , \31154 ,
         \31155 , \31156 , \31157 , \31158 , \31159 , \31160 , \31161 , \31162 , \31163 , \31164 ,
         \31165 , \31166 , \31167 , \31168 , \31169 , \31170 , \31171 , \31172 , \31173 , \31174 ,
         \31175 , \31176 , \31177 , \31178 , \31179 , \31180 , \31181 , \31182 , \31183 , \31184 ,
         \31185 , \31186 , \31187 , \31188 , \31189 , \31190 , \31191 , \31192 , \31193 , \31194 ,
         \31195 , \31196 , \31197 , \31198 , \31199 , \31200 , \31201 , \31202 , \31203 , \31204 ,
         \31205 , \31206 , \31207 , \31208 , \31209 , \31210 , \31211 , \31212 , \31213 , \31214 ,
         \31215 , \31216 , \31217 , \31218 , \31219 , \31220 , \31221 , \31222 , \31223 , \31224 ,
         \31225 , \31226 , \31227 , \31228 , \31229 , \31230 , \31231 , \31232 , \31233 , \31234 ,
         \31235 , \31236 , \31237 , \31238 , \31239 , \31240 , \31241 , \31242 , \31243 , \31244 ,
         \31245 , \31246 , \31247 , \31248 , \31249 , \31250 , \31251 , \31252 , \31253 , \31254 ,
         \31255 , \31256 , \31257 , \31258 , \31259 , \31260 , \31261 , \31262 , \31263 , \31264 ,
         \31265 , \31266 , \31267 , \31268 , \31269 , \31270 , \31271 , \31272 , \31273 , \31274 ,
         \31275 , \31276 , \31277 , \31278 , \31279 , \31280 , \31281 , \31282 , \31283 , \31284 ,
         \31285 , \31286 , \31287 , \31288 , \31289 , \31290 , \31291 , \31292 , \31293 , \31294 ,
         \31295 , \31296 , \31297 , \31298 , \31299 , \31300 , \31301 , \31302 , \31303 , \31304 ,
         \31305 , \31306 , \31307 , \31308 , \31309 , \31310 , \31311 , \31312 , \31313 , \31314 ,
         \31315 , \31316 , \31317 , \31318 , \31319 , \31320 , \31321 , \31322 , \31323 , \31324 ,
         \31325 , \31326 , \31327 , \31328 , \31329 , \31330 , \31331 , \31332 , \31333 , \31334 ,
         \31335 , \31336 , \31337 , \31338 , \31339 , \31340 , \31341 , \31342 , \31343 , \31344 ,
         \31345 , \31346 , \31347 , \31348 , \31349 , \31350 , \31351 , \31352 , \31353 , \31354 ,
         \31355 , \31356 , \31357 , \31358 , \31359 , \31360 , \31361 , \31362 , \31363 , \31364 ,
         \31365 , \31366 , \31367 , \31368 , \31369 , \31370 , \31371 , \31372 , \31373 , \31374 ,
         \31375 , \31376 , \31377 , \31378 , \31379 , \31380 , \31381 , \31382 , \31383 , \31384 ,
         \31385 , \31386 , \31387 , \31388 , \31389 , \31390 , \31391 , \31392 , \31393 , \31394 ,
         \31395 , \31396 , \31397 , \31398 , \31399 , \31400 , \31401 , \31402 , \31403 , \31404 ,
         \31405 , \31406 , \31407 , \31408 , \31409 , \31410 , \31411 , \31412 , \31413 , \31414 ,
         \31415 , \31416 , \31417 , \31418 , \31419 , \31420 , \31421 , \31422 , \31423 , \31424 ,
         \31425 , \31426 , \31427 , \31428 , \31429 , \31430 , \31431 , \31432 , \31433 , \31434 ,
         \31435 , \31436 , \31437 , \31438 , \31439 , \31440 , \31441 , \31442 , \31443 , \31444 ,
         \31445 , \31446 , \31447 , \31448 , \31449 , \31450 , \31451 , \31452 , \31453 , \31454 ,
         \31455 , \31456 , \31457 , \31458 , \31459 , \31460 , \31461 , \31462 , \31463 , \31464 ,
         \31465 , \31466 , \31467 , \31468 , \31469 , \31470 , \31471 , \31472 , \31473 , \31474 ,
         \31475 , \31476 , \31477 , \31478 , \31479 , \31480 , \31481 , \31482 , \31483 , \31484 ,
         \31485 , \31486 , \31487 , \31488 , \31489 , \31490 , \31491 , \31492 , \31493 , \31494 ,
         \31495 , \31496 , \31497 , \31498 , \31499 , \31500 , \31501 , \31502 , \31503 , \31504 ,
         \31505 , \31506 , \31507 , \31508 , \31509 , \31510 , \31511 , \31512 , \31513 , \31514 ,
         \31515 , \31516 , \31517 , \31518 , \31519 , \31520 , \31521 , \31522 , \31523 , \31524 ,
         \31525 , \31526 , \31527 , \31528 , \31529 , \31530 , \31531 , \31532 , \31533 , \31534 ,
         \31535 , \31536 , \31537 , \31538 , \31539 , \31540 , \31541 , \31542 , \31543 , \31544 ,
         \31545 , \31546 , \31547 , \31548 , \31549 , \31550 , \31551 , \31552 , \31553 , \31554 ,
         \31555 , \31556 , \31557 , \31558 , \31559 , \31560 , \31561 , \31562 , \31563 , \31564 ,
         \31565 , \31566 , \31567 , \31568 , \31569 , \31570 , \31571 , \31572 , \31573 , \31574 ,
         \31575 , \31576 , \31577 , \31578 , \31579 , \31580 , \31581 , \31582 , \31583 , \31584 ,
         \31585 , \31586 , \31587 , \31588 , \31589 , \31590 , \31591 , \31592 , \31593 , \31594 ,
         \31595 , \31596 , \31597 , \31598 , \31599 , \31600 , \31601 , \31602 , \31603 , \31604 ,
         \31605 , \31606 , \31607 , \31608 , \31609 , \31610 , \31611 , \31612 , \31613 , \31614 ,
         \31615 , \31616 , \31617 , \31618 , \31619 , \31620 , \31621 , \31622 , \31623 , \31624 ,
         \31625 , \31626 , \31627 , \31628 , \31629 , \31630 , \31631 , \31632 , \31633 , \31634 ,
         \31635 , \31636 , \31637 , \31638 , \31639 , \31640 , \31641 , \31642 , \31643 , \31644 ,
         \31645 , \31646 , \31647 , \31648 , \31649 , \31650 , \31651 , \31652 , \31653 , \31654 ,
         \31655 , \31656 , \31657 , \31658 , \31659 , \31660 , \31661 , \31662 , \31663 , \31664 ,
         \31665 , \31666 , \31667 , \31668 , \31669 , \31670 , \31671 , \31672 , \31673 , \31674 ,
         \31675 , \31676 , \31677 , \31678 , \31679 , \31680 , \31681 , \31682 , \31683 , \31684 ,
         \31685 , \31686 , \31687 , \31688 , \31689 , \31690 , \31691 , \31692 , \31693 , \31694 ,
         \31695 , \31696 , \31697 , \31698 , \31699 , \31700 , \31701 , \31702 , \31703 , \31704 ,
         \31705 , \31706 , \31707 , \31708 , \31709 , \31710 , \31711 , \31712 , \31713 , \31714 ,
         \31715 , \31716 , \31717 , \31718 , \31719 , \31720 , \31721 , \31722 , \31723 , \31724 ,
         \31725 , \31726 , \31727 , \31728 , \31729 , \31730 , \31731 , \31732 , \31733 , \31734 ,
         \31735 , \31736 , \31737 , \31738 , \31739 , \31740 , \31741 , \31742 , \31743 , \31744 ,
         \31745 , \31746 , \31747 , \31748 , \31749 , \31750 , \31751 , \31752 , \31753 , \31754 ,
         \31755 , \31756 , \31757 , \31758 , \31759 , \31760 , \31761 , \31762 , \31763 , \31764 ,
         \31765 , \31766 , \31767 , \31768 , \31769 , \31770 , \31771 , \31772 , \31773 , \31774 ,
         \31775 , \31776 , \31777 , \31778 , \31779 , \31780 , \31781 , \31782 , \31783 , \31784 ,
         \31785 , \31786 , \31787 , \31788 , \31789 , \31790 , \31791 , \31792 , \31793 , \31794 ,
         \31795 , \31796 , \31797 , \31798 , \31799 , \31800 , \31801 , \31802 , \31803 , \31804 ,
         \31805 , \31806 , \31807 , \31808 , \31809 , \31810 , \31811 , \31812 , \31813 , \31814 ,
         \31815 , \31816 , \31817 , \31818 , \31819 , \31820 , \31821 , \31822 , \31823 , \31824 ,
         \31825 , \31826 , \31827 , \31828 , \31829 , \31830 , \31831 , \31832 , \31833 , \31834 ,
         \31835 , \31836 , \31837 , \31838 , \31839 , \31840 , \31841 , \31842 , \31843 , \31844 ,
         \31845 , \31846 , \31847 , \31848 , \31849 , \31850 , \31851 , \31852 , \31853 , \31854 ,
         \31855 , \31856 , \31857 , \31858 , \31859 , \31860 , \31861 , \31862 , \31863 , \31864 ,
         \31865 , \31866 , \31867 , \31868 , \31869 , \31870 , \31871 , \31872 , \31873 , \31874 ,
         \31875 , \31876 , \31877 , \31878 , \31879 , \31880 , \31881 , \31882 , \31883 , \31884 ,
         \31885 , \31886 , \31887 , \31888 , \31889 , \31890 , \31891 , \31892 , \31893 , \31894 ,
         \31895 , \31896 , \31897 , \31898 , \31899 , \31900 , \31901 , \31902 , \31903 , \31904 ,
         \31905 , \31906 , \31907 , \31908 , \31909 , \31910 , \31911 , \31912 , \31913 , \31914 ,
         \31915 , \31916 , \31917 , \31918 , \31919 , \31920 , \31921 , \31922 , \31923 , \31924 ,
         \31925 , \31926 , \31927 , \31928 , \31929 , \31930 , \31931 , \31932 , \31933 , \31934 ,
         \31935 , \31936 , \31937 , \31938 , \31939 , \31940 , \31941 , \31942 , \31943 , \31944 ,
         \31945 , \31946 , \31947 , \31948 , \31949 , \31950 , \31951 , \31952 , \31953 , \31954 ,
         \31955 , \31956 , \31957 , \31958 , \31959 , \31960 , \31961 , \31962 , \31963 , \31964 ,
         \31965 , \31966 , \31967 , \31968 , \31969 , \31970 , \31971 , \31972 , \31973 , \31974 ,
         \31975 , \31976 , \31977 , \31978 , \31979 , \31980 , \31981 , \31982 , \31983 , \31984 ,
         \31985 , \31986 , \31987 , \31988 , \31989 , \31990 , \31991 , \31992 , \31993 , \31994 ,
         \31995 , \31996 , \31997 , \31998 , \31999 , \32000 , \32001 , \32002 , \32003 , \32004 ,
         \32005 , \32006 , \32007 , \32008 , \32009 , \32010 , \32011 , \32012 , \32013 , \32014 ,
         \32015 , \32016 , \32017 , \32018 , \32019 , \32020 , \32021 , \32022 , \32023 , \32024 ,
         \32025 , \32026 , \32027 , \32028 , \32029 , \32030 , \32031 , \32032 , \32033 , \32034 ,
         \32035 , \32036 , \32037 , \32038 , \32039 , \32040 , \32041 , \32042 , \32043 , \32044 ,
         \32045 , \32046 , \32047 , \32048 , \32049 , \32050 , \32051 , \32052 , \32053 , \32054 ,
         \32055 , \32056 , \32057 , \32058 , \32059 , \32060 , \32061 , \32062 , \32063 , \32064 ,
         \32065 , \32066 , \32067 , \32068 , \32069 , \32070 , \32071 , \32072 , \32073 , \32074 ,
         \32075 , \32076 , \32077 , \32078 , \32079 , \32080 , \32081 , \32082 , \32083 , \32084 ,
         \32085 , \32086 , \32087 , \32088 , \32089 , \32090 , \32091 , \32092 , \32093 , \32094 ,
         \32095 , \32096 , \32097 , \32098 , \32099 , \32100 , \32101 , \32102 , \32103 , \32104 ,
         \32105 , \32106 , \32107 , \32108 , \32109 , \32110 , \32111 , \32112 , \32113 , \32114 ,
         \32115 , \32116 , \32117 , \32118 , \32119 , \32120 , \32121 , \32122 , \32123 , \32124 ,
         \32125 , \32126 , \32127 , \32128 , \32129 , \32130 , \32131 , \32132 , \32133 , \32134 ,
         \32135 , \32136 , \32137 , \32138 , \32139 , \32140 , \32141 , \32142 , \32143 , \32144 ,
         \32145 , \32146 , \32147 , \32148 , \32149 , \32150 , \32151 , \32152 , \32153 , \32154 ,
         \32155 , \32156 , \32157 , \32158 , \32159 , \32160 , \32161 , \32162 , \32163 , \32164 ,
         \32165 , \32166 , \32167 , \32168 , \32169 , \32170 , \32171 , \32172 , \32173 , \32174 ,
         \32175 , \32176 , \32177 , \32178 , \32179 , \32180 , \32181 , \32182 , \32183 , \32184 ,
         \32185 , \32186 , \32187 , \32188 , \32189 , \32190 , \32191 , \32192 , \32193 , \32194 ,
         \32195 , \32196 , \32197 , \32198 , \32199 , \32200 , \32201 , \32202 , \32203 , \32204 ,
         \32205 , \32206 , \32207 , \32208 , \32209 , \32210 , \32211 , \32212 , \32213 , \32214 ,
         \32215 , \32216 , \32217 , \32218 , \32219 , \32220 , \32221 , \32222 , \32223 , \32224 ,
         \32225 , \32226 , \32227 , \32228 , \32229 , \32230 , \32231 , \32232 , \32233 , \32234 ,
         \32235 , \32236 , \32237 , \32238 , \32239 , \32240 , \32241 , \32242 , \32243 , \32244 ,
         \32245 , \32246 , \32247 , \32248 , \32249 , \32250 , \32251 , \32252 , \32253 , \32254 ,
         \32255 , \32256 , \32257 , \32258 , \32259 , \32260 , \32261 , \32262 , \32263 , \32264 ,
         \32265 , \32266 , \32267 , \32268 , \32269 , \32270 , \32271 , \32272 , \32273 , \32274 ,
         \32275 , \32276 , \32277 , \32278 , \32279 , \32280 , \32281 , \32282 , \32283 , \32284 ,
         \32285 , \32286 , \32287 , \32288 , \32289 , \32290 , \32291 , \32292 , \32293 , \32294 ,
         \32295 , \32296 , \32297 , \32298 , \32299 , \32300 , \32301 , \32302 , \32303 , \32304 ,
         \32305 , \32306 , \32307 , \32308 , \32309 , \32310 , \32311 , \32312 , \32313 , \32314 ,
         \32315 , \32316 , \32317 , \32318 , \32319 , \32320 , \32321 , \32322 , \32323 , \32324 ,
         \32325 , \32326 , \32327 , \32328 , \32329 , \32330 , \32331 , \32332 , \32333 , \32334 ,
         \32335 , \32336 , \32337 , \32338 , \32339 , \32340 , \32341 , \32342 , \32343 , \32344 ,
         \32345 , \32346 , \32347 , \32348 , \32349 , \32350 , \32351 , \32352 , \32353 , \32354 ,
         \32355 , \32356 , \32357 , \32358 , \32359 , \32360 , \32361 , \32362 , \32363 , \32364 ,
         \32365 , \32366 , \32367 , \32368 , \32369 , \32370 , \32371 , \32372 , \32373 , \32374 ,
         \32375 , \32376 , \32377 , \32378 , \32379 , \32380 , \32381 , \32382 , \32383 , \32384 ,
         \32385 , \32386 , \32387 , \32388 , \32389 , \32390 , \32391 , \32392 , \32393 , \32394 ,
         \32395 , \32396 , \32397 , \32398 , \32399 , \32400 , \32401 , \32402 , \32403 , \32404 ,
         \32405 , \32406 , \32407 , \32408 , \32409 , \32410 , \32411 , \32412 , \32413 , \32414 ,
         \32415 , \32416 , \32417 , \32418 , \32419 , \32420 , \32421 , \32422 , \32423 , \32424 ,
         \32425 , \32426 , \32427 , \32428 , \32429 , \32430 , \32431 , \32432 , \32433 , \32434 ,
         \32435 , \32436 , \32437 , \32438 , \32439 , \32440 , \32441 , \32442 , \32443 , \32444 ,
         \32445 , \32446 , \32447 , \32448 , \32449 , \32450 , \32451 , \32452 , \32453 , \32454 ,
         \32455 , \32456 , \32457 , \32458 , \32459 , \32460 , \32461 , \32462 , \32463 , \32464 ,
         \32465 , \32466 , \32467 , \32468 , \32469 , \32470 , \32471 , \32472 , \32473 , \32474 ,
         \32475 , \32476 , \32477 , \32478 , \32479 , \32480 , \32481 , \32482 , \32483 , \32484 ,
         \32485 , \32486 , \32487 , \32488 , \32489 , \32490 , \32491 , \32492 , \32493 , \32494 ,
         \32495 , \32496 , \32497 , \32498 , \32499 , \32500 , \32501 , \32502 , \32503 , \32504 ,
         \32505 , \32506 , \32507 , \32508 , \32509 , \32510 , \32511 , \32512 , \32513 , \32514 ,
         \32515 , \32516 , \32517 , \32518 , \32519 , \32520 , \32521 , \32522 , \32523 , \32524 ,
         \32525 , \32526 , \32527 , \32528 , \32529 , \32530 , \32531 , \32532 , \32533 , \32534 ,
         \32535 , \32536 , \32537 , \32538 , \32539 , \32540 , \32541 , \32542 , \32543 , \32544 ,
         \32545 , \32546 , \32547 , \32548 , \32549 , \32550 , \32551 , \32552 , \32553 , \32554 ,
         \32555 , \32556 , \32557 , \32558 , \32559 , \32560 , \32561 , \32562 , \32563 , \32564 ,
         \32565 , \32566 , \32567 , \32568 , \32569 , \32570 , \32571 , \32572 , \32573 , \32574 ,
         \32575 , \32576 , \32577 , \32578 , \32579 , \32580 , \32581 , \32582 , \32583 , \32584 ,
         \32585 , \32586 , \32587 , \32588 , \32589 , \32590 , \32591 , \32592 , \32593 , \32594 ,
         \32595 , \32596 , \32597 , \32598 , \32599 , \32600 , \32601 , \32602 , \32603 , \32604 ,
         \32605 , \32606 , \32607 , \32608 , \32609 , \32610 , \32611 , \32612 , \32613 , \32614 ,
         \32615 , \32616 , \32617 , \32618 , \32619 , \32620 , \32621 , \32622 , \32623 , \32624 ,
         \32625 , \32626 , \32627 , \32628 , \32629 , \32630 , \32631 , \32632 , \32633 , \32634 ,
         \32635 , \32636 , \32637 , \32638 , \32639 , \32640 , \32641 , \32642 , \32643 , \32644 ,
         \32645 , \32646 , \32647 , \32648 , \32649 , \32650 , \32651 , \32652 , \32653 , \32654 ,
         \32655 , \32656 , \32657 , \32658 , \32659 , \32660 , \32661 , \32662 , \32663 , \32664 ,
         \32665 , \32666 , \32667 , \32668 , \32669 , \32670 , \32671 , \32672 , \32673 , \32674 ,
         \32675 , \32676 , \32677 , \32678 , \32679 , \32680 , \32681 , \32682 , \32683 , \32684 ,
         \32685 , \32686 , \32687 , \32688 , \32689 , \32690 , \32691 , \32692 , \32693 , \32694 ,
         \32695 , \32696 , \32697 , \32698 , \32699 , \32700 , \32701 , \32702 , \32703 , \32704 ,
         \32705 , \32706 , \32707 , \32708 , \32709 , \32710 , \32711 , \32712 , \32713 , \32714 ,
         \32715 , \32716 , \32717 , \32718 , \32719 , \32720 , \32721 , \32722 , \32723 , \32724 ,
         \32725 , \32726 , \32727 , \32728 , \32729 , \32730 , \32731 , \32732 , \32733 , \32734 ,
         \32735 , \32736 , \32737 , \32738 , \32739 , \32740 , \32741 , \32742 , \32743 , \32744 ,
         \32745 , \32746 , \32747 , \32748 , \32749 , \32750 , \32751 , \32752 , \32753 , \32754 ,
         \32755 , \32756 , \32757 , \32758 , \32759 , \32760 , \32761 , \32762 , \32763 , \32764 ,
         \32765 , \32766 , \32767 , \32768 , \32769 , \32770 , \32771 , \32772 , \32773 , \32774 ,
         \32775 , \32776 , \32777 , \32778 , \32779 , \32780 , \32781 , \32782 , \32783 , \32784 ,
         \32785 , \32786 , \32787 , \32788 , \32789 , \32790 , \32791 , \32792 , \32793 , \32794 ,
         \32795 , \32796 , \32797 , \32798 , \32799 , \32800 , \32801 , \32802 , \32803 , \32804 ,
         \32805 , \32806 , \32807 , \32808 , \32809 , \32810 , \32811 , \32812 , \32813 , \32814 ,
         \32815 , \32816 , \32817 , \32818 , \32819 , \32820 , \32821 , \32822 , \32823 , \32824 ,
         \32825 , \32826 , \32827 , \32828 , \32829 , \32830 , \32831 , \32832 , \32833 , \32834 ,
         \32835 , \32836 , \32837 , \32838 , \32839 , \32840 , \32841 , \32842 , \32843 , \32844 ,
         \32845 , \32846 , \32847 , \32848 , \32849 , \32850 , \32851 , \32852 , \32853 , \32854 ,
         \32855 , \32856 , \32857 , \32858 , \32859 , \32860 , \32861 , \32862 , \32863 , \32864 ,
         \32865 , \32866 , \32867 , \32868 , \32869 , \32870 , \32871 , \32872 , \32873 , \32874 ,
         \32875 , \32876 , \32877 , \32878 , \32879 , \32880 , \32881 , \32882 , \32883 , \32884 ,
         \32885 , \32886 , \32887 , \32888 , \32889 , \32890 , \32891 , \32892 , \32893 , \32894 ,
         \32895 , \32896 , \32897 , \32898 , \32899 , \32900 , \32901 , \32902 , \32903 , \32904 ,
         \32905 , \32906 , \32907 , \32908 , \32909 , \32910 , \32911 , \32912 , \32913 , \32914 ,
         \32915 , \32916 , \32917 , \32918 , \32919 , \32920 , \32921 , \32922 , \32923 , \32924 ,
         \32925 , \32926 , \32927 , \32928 , \32929 , \32930 , \32931 , \32932 , \32933 , \32934 ,
         \32935 , \32936 , \32937 , \32938 , \32939 , \32940 , \32941 , \32942 , \32943 , \32944 ,
         \32945 , \32946 , \32947 , \32948 , \32949 , \32950 , \32951 , \32952 , \32953 , \32954 ,
         \32955 , \32956 , \32957 , \32958 , \32959 , \32960 , \32961 , \32962 , \32963 , \32964 ,
         \32965 , \32966 , \32967 , \32968 , \32969 , \32970 , \32971 , \32972 , \32973 , \32974 ,
         \32975 , \32976 , \32977 , \32978 , \32979 , \32980 , \32981 , \32982 , \32983 , \32984 ,
         \32985 , \32986 , \32987 , \32988 , \32989 , \32990 , \32991 , \32992 , \32993 , \32994 ,
         \32995 , \32996 , \32997 , \32998 , \32999 , \33000 , \33001 , \33002 , \33003 , \33004 ,
         \33005 , \33006 , \33007 , \33008 , \33009 , \33010 , \33011 , \33012 , \33013 , \33014 ,
         \33015 , \33016 , \33017 , \33018 , \33019 , \33020 , \33021 , \33022 , \33023 , \33024 ,
         \33025 , \33026 , \33027 , \33028 , \33029 , \33030 , \33031 , \33032 , \33033 , \33034 ,
         \33035 , \33036 , \33037 , \33038 , \33039 , \33040 , \33041 , \33042 , \33043 , \33044 ,
         \33045 , \33046 , \33047 , \33048 , \33049 , \33050 , \33051 , \33052 , \33053 , \33054 ,
         \33055 , \33056 , \33057 , \33058 , \33059 , \33060 , \33061 , \33062 , \33063 , \33064 ,
         \33065 , \33066 , \33067 , \33068 , \33069 , \33070 , \33071 , \33072 , \33073 , \33074 ,
         \33075 , \33076 , \33077 , \33078 , \33079 , \33080 , \33081 , \33082 , \33083 , \33084 ,
         \33085 , \33086 , \33087 , \33088 , \33089 , \33090 , \33091 , \33092 , \33093 , \33094 ,
         \33095 , \33096 , \33097 , \33098 , \33099 , \33100 , \33101 , \33102 , \33103 , \33104 ,
         \33105 , \33106 , \33107 , \33108 , \33109 , \33110 , \33111 , \33112 , \33113 , \33114 ,
         \33115 , \33116 , \33117 , \33118 , \33119 , \33120 , \33121 , \33122 , \33123 , \33124 ,
         \33125 , \33126 , \33127 , \33128 , \33129 , \33130 , \33131 , \33132 , \33133 , \33134 ,
         \33135 , \33136 , \33137 , \33138 , \33139 , \33140 , \33141 , \33142 , \33143 , \33144 ,
         \33145 , \33146 , \33147 , \33148 , \33149 , \33150 , \33151 , \33152 , \33153 , \33154 ,
         \33155 , \33156 , \33157 , \33158 , \33159 , \33160 , \33161 , \33162 , \33163 , \33164 ,
         \33165 , \33166 , \33167 , \33168 , \33169 , \33170 , \33171 , \33172 , \33173 , \33174 ,
         \33175 , \33176 , \33177 , \33178 , \33179 , \33180 , \33181 , \33182 , \33183 , \33184 ,
         \33185 , \33186 , \33187 , \33188 , \33189 , \33190 , \33191 , \33192 , \33193 , \33194 ,
         \33195 , \33196 , \33197 , \33198 , \33199 , \33200 , \33201 , \33202 , \33203 , \33204 ,
         \33205 , \33206 , \33207 , \33208 , \33209 , \33210 , \33211 , \33212 , \33213 , \33214 ,
         \33215 , \33216 , \33217 , \33218 , \33219 , \33220 , \33221 , \33222 , \33223 , \33224 ,
         \33225 , \33226 , \33227 , \33228 , \33229 , \33230 , \33231 , \33232 , \33233 , \33234 ,
         \33235 , \33236 , \33237 , \33238 , \33239 , \33240 , \33241 , \33242 , \33243 , \33244 ,
         \33245 , \33246 , \33247 , \33248 , \33249 , \33250 , \33251 , \33252 , \33253 , \33254 ,
         \33255 , \33256 , \33257 , \33258 , \33259 , \33260 , \33261 , \33262 , \33263 , \33264 ,
         \33265 , \33266 , \33267 , \33268 , \33269 , \33270 , \33271 , \33272 , \33273 , \33274 ,
         \33275 , \33276 , \33277 , \33278 , \33279 , \33280 , \33281 , \33282 , \33283 , \33284 ,
         \33285 , \33286 , \33287 , \33288 , \33289 , \33290 , \33291 , \33292 , \33293 , \33294 ,
         \33295 , \33296 , \33297 , \33298 , \33299 , \33300 , \33301 , \33302 , \33303 , \33304 ,
         \33305 , \33306 , \33307 , \33308 , \33309 , \33310 , \33311 , \33312 , \33313 , \33314 ,
         \33315 , \33316 , \33317 , \33318 , \33319 , \33320 , \33321 , \33322 , \33323 , \33324 ,
         \33325 , \33326 , \33327 , \33328 , \33329 , \33330 , \33331 , \33332 , \33333 , \33334 ,
         \33335 , \33336 , \33337 , \33338 , \33339 , \33340 , \33341 , \33342 , \33343 , \33344 ,
         \33345 , \33346 , \33347 , \33348 , \33349 , \33350 , \33351 , \33352 , \33353 , \33354 ,
         \33355 , \33356 , \33357 , \33358 , \33359 , \33360 , \33361 , \33362 , \33363 , \33364 ,
         \33365 , \33366 , \33367 , \33368 , \33369 , \33370 , \33371 , \33372 , \33373 , \33374 ,
         \33375 , \33376 , \33377 , \33378 , \33379 , \33380 , \33381 , \33382 , \33383 , \33384 ,
         \33385 , \33386 , \33387 , \33388 , \33389 , \33390 , \33391 , \33392 , \33393 , \33394 ,
         \33395 , \33396 , \33397 , \33398 , \33399 , \33400 , \33401 , \33402 , \33403 , \33404 ,
         \33405 , \33406 , \33407 , \33408 , \33409 , \33410 , \33411 , \33412 , \33413 , \33414 ,
         \33415 , \33416 , \33417 , \33418 , \33419 , \33420 , \33421 , \33422 , \33423 , \33424 ,
         \33425 , \33426 , \33427 , \33428 , \33429 , \33430 , \33431 , \33432 , \33433 , \33434 ,
         \33435 , \33436 , \33437 , \33438 , \33439 , \33440 , \33441 , \33442 , \33443 , \33444 ,
         \33445 , \33446 , \33447 , \33448 , \33449 , \33450 , \33451 , \33452 , \33453 , \33454 ,
         \33455 , \33456 , \33457 , \33458 , \33459 , \33460 , \33461 , \33462 , \33463 , \33464 ,
         \33465 , \33466 , \33467 , \33468 , \33469 , \33470 , \33471 , \33472 , \33473 , \33474 ,
         \33475 , \33476 , \33477 , \33478 , \33479 , \33480 , \33481 , \33482 , \33483 , \33484 ,
         \33485 , \33486 , \33487 , \33488 , \33489 , \33490 , \33491 , \33492 , \33493 , \33494 ,
         \33495 , \33496 , \33497 , \33498 , \33499 , \33500 , \33501 , \33502 , \33503 , \33504 ,
         \33505 , \33506 , \33507 , \33508 , \33509 , \33510 , \33511 , \33512 , \33513 , \33514 ,
         \33515 , \33516 , \33517 , \33518 , \33519 , \33520 , \33521 , \33522 , \33523 , \33524 ,
         \33525 , \33526 , \33527 , \33528 , \33529 , \33530 , \33531 , \33532 , \33533 , \33534 ,
         \33535 , \33536 , \33537 , \33538 , \33539 , \33540 , \33541 , \33542 , \33543 , \33544 ,
         \33545 , \33546 , \33547 , \33548 , \33549 , \33550 , \33551 , \33552 , \33553 , \33554 ,
         \33555 , \33556 , \33557 , \33558 , \33559 , \33560 , \33561 , \33562 , \33563 , \33564 ,
         \33565 , \33566 , \33567 , \33568 , \33569 , \33570 , \33571 , \33572 , \33573 , \33574 ,
         \33575 , \33576 , \33577 , \33578 , \33579 , \33580 , \33581 , \33582 , \33583 , \33584 ,
         \33585 , \33586 , \33587 , \33588 , \33589 , \33590 , \33591 , \33592 , \33593 , \33594 ,
         \33595 , \33596 , \33597 , \33598 , \33599 , \33600 , \33601 , \33602 , \33603 , \33604 ,
         \33605 , \33606 , \33607 , \33608 , \33609 , \33610 , \33611 , \33612 , \33613 , \33614 ,
         \33615 , \33616 , \33617 , \33618 , \33619 , \33620 , \33621 , \33622 , \33623 , \33624 ,
         \33625 , \33626 , \33627 , \33628 , \33629 , \33630 , \33631 , \33632 , \33633 , \33634 ,
         \33635 , \33636 , \33637 , \33638 , \33639 , \33640 , \33641 , \33642 , \33643 , \33644 ,
         \33645 , \33646 , \33647 , \33648 , \33649 , \33650 , \33651 , \33652 , \33653 , \33654 ,
         \33655 , \33656 , \33657 , \33658 , \33659 , \33660 , \33661 , \33662 , \33663 , \33664 ,
         \33665 , \33666 , \33667 , \33668 , \33669 , \33670 , \33671 , \33672 , \33673 , \33674 ,
         \33675 , \33676 , \33677 , \33678 , \33679 , \33680 , \33681 , \33682 , \33683 , \33684 ,
         \33685 , \33686 , \33687 , \33688 , \33689 , \33690 , \33691 , \33692 , \33693 , \33694 ,
         \33695 , \33696 , \33697 , \33698 , \33699 , \33700 , \33701 , \33702 , \33703 , \33704 ,
         \33705 , \33706 , \33707 , \33708 , \33709 , \33710 , \33711 , \33712 , \33713 , \33714 ,
         \33715 , \33716 , \33717 , \33718 , \33719 , \33720 , \33721 , \33722 , \33723 , \33724 ,
         \33725 , \33726 , \33727 , \33728 , \33729 , \33730 , \33731 , \33732 , \33733 , \33734 ,
         \33735 , \33736 , \33737 , \33738 , \33739 , \33740 , \33741 , \33742 , \33743 , \33744 ,
         \33745 , \33746 , \33747 , \33748 , \33749 , \33750 , \33751 , \33752 , \33753 , \33754 ,
         \33755 , \33756 , \33757 , \33758 , \33759 , \33760 , \33761 , \33762 , \33763 , \33764 ,
         \33765 , \33766 , \33767 , \33768 , \33769 , \33770 , \33771 , \33772 , \33773 , \33774 ,
         \33775 , \33776 , \33777 , \33778 , \33779 , \33780 , \33781 , \33782 , \33783 , \33784 ,
         \33785 , \33786 , \33787 , \33788 , \33789 , \33790 , \33791 , \33792 , \33793 , \33794 ,
         \33795 , \33796 , \33797 , \33798 , \33799 , \33800 , \33801 , \33802 , \33803 , \33804 ,
         \33805 , \33806 , \33807 , \33808 , \33809 , \33810 , \33811 , \33812 , \33813 , \33814 ,
         \33815 , \33816 , \33817 , \33818 , \33819 , \33820 , \33821 , \33822 , \33823 , \33824 ,
         \33825 , \33826 , \33827 , \33828 , \33829 , \33830 , \33831 , \33832 , \33833 , \33834 ,
         \33835 , \33836 , \33837 , \33838 , \33839 , \33840 , \33841 , \33842 , \33843 , \33844 ,
         \33845 , \33846 , \33847 , \33848 , \33849 , \33850 , \33851 , \33852 , \33853 , \33854 ,
         \33855 , \33856 , \33857 , \33858 , \33859 , \33860 , \33861 , \33862 , \33863 , \33864 ,
         \33865 , \33866 , \33867 , \33868 , \33869 , \33870 , \33871 , \33872 , \33873 , \33874 ,
         \33875 , \33876 , \33877 , \33878 , \33879 , \33880 , \33881 , \33882 , \33883 , \33884 ,
         \33885 , \33886 , \33887 , \33888 , \33889 , \33890 , \33891 , \33892 , \33893 , \33894 ,
         \33895 , \33896 , \33897 , \33898 , \33899 , \33900 , \33901 , \33902 , \33903 , \33904 ,
         \33905 , \33906 , \33907 , \33908 , \33909 , \33910 , \33911 , \33912 , \33913 , \33914 ,
         \33915 , \33916 , \33917 , \33918 , \33919 , \33920 , \33921 , \33922 , \33923 , \33924 ,
         \33925 , \33926 , \33927 , \33928 , \33929 , \33930 , \33931 , \33932 , \33933 , \33934 ,
         \33935 , \33936 , \33937 , \33938 , \33939 , \33940 , \33941 , \33942 , \33943 , \33944 ,
         \33945 , \33946 , \33947 , \33948 , \33949 , \33950 , \33951 , \33952 , \33953 , \33954 ,
         \33955 , \33956 , \33957 , \33958 , \33959 , \33960 , \33961 , \33962 , \33963 , \33964 ,
         \33965 , \33966 , \33967 , \33968 , \33969 , \33970 , \33971 , \33972 , \33973 , \33974 ,
         \33975 , \33976 , \33977 , \33978 , \33979 , \33980 , \33981 , \33982 , \33983 , \33984 ,
         \33985 , \33986 , \33987 , \33988 , \33989 , \33990 , \33991 , \33992 , \33993 , \33994 ,
         \33995 , \33996 , \33997 , \33998 , \33999 , \34000 , \34001 , \34002 , \34003 , \34004 ,
         \34005 , \34006 , \34007 , \34008 , \34009 , \34010 , \34011 , \34012 , \34013 , \34014 ,
         \34015 , \34016 , \34017 , \34018 , \34019 , \34020 , \34021 , \34022 , \34023 , \34024 ,
         \34025 , \34026 , \34027 , \34028 , \34029 , \34030 , \34031 , \34032 , \34033 , \34034 ,
         \34035 , \34036 , \34037 , \34038 , \34039 , \34040 , \34041 , \34042 , \34043 , \34044 ,
         \34045 , \34046 , \34047 , \34048 , \34049 , \34050 , \34051 , \34052 , \34053 , \34054 ,
         \34055 , \34056 , \34057 , \34058 , \34059 , \34060 , \34061 , \34062 , \34063 , \34064 ,
         \34065 , \34066 , \34067 , \34068 , \34069 , \34070 , \34071 , \34072 , \34073 , \34074 ,
         \34075 , \34076 , \34077 , \34078 , \34079 , \34080 , \34081 , \34082 , \34083 , \34084 ,
         \34085 , \34086 , \34087 , \34088 , \34089 , \34090 , \34091 , \34092 , \34093 , \34094 ,
         \34095 , \34096 , \34097 , \34098 , \34099 , \34100 , \34101 , \34102 , \34103 , \34104 ,
         \34105 , \34106 , \34107 , \34108 , \34109 , \34110 , \34111 , \34112 , \34113 , \34114 ,
         \34115 , \34116 , \34117 , \34118 , \34119 , \34120 , \34121 , \34122 , \34123 , \34124 ,
         \34125 , \34126 , \34127 , \34128 , \34129 , \34130 , \34131 , \34132 , \34133 , \34134 ,
         \34135 , \34136 , \34137 , \34138 , \34139 , \34140 , \34141 , \34142 , \34143 , \34144 ,
         \34145 , \34146 , \34147 , \34148 , \34149 , \34150 , \34151 , \34152 , \34153 , \34154 ,
         \34155 , \34156 , \34157 , \34158 , \34159 , \34160 , \34161 , \34162 , \34163 , \34164 ,
         \34165 , \34166 , \34167 , \34168 , \34169 , \34170 , \34171 , \34172 , \34173 , \34174 ,
         \34175 , \34176 , \34177 , \34178 , \34179 , \34180 , \34181 , \34182 , \34183 , \34184 ,
         \34185 , \34186 , \34187 , \34188 , \34189 , \34190 , \34191 , \34192 , \34193 , \34194 ,
         \34195 , \34196 , \34197 , \34198 , \34199 , \34200 , \34201 , \34202 , \34203 , \34204 ,
         \34205 , \34206 , \34207 , \34208 , \34209 , \34210 , \34211 , \34212 , \34213 , \34214 ,
         \34215 , \34216 , \34217 , \34218 , \34219 , \34220 , \34221 , \34222 , \34223 , \34224 ,
         \34225 , \34226 , \34227 , \34228 , \34229 , \34230 , \34231 , \34232 , \34233 , \34234 ,
         \34235 , \34236 , \34237 , \34238 , \34239 , \34240 , \34241 , \34242 , \34243 , \34244 ,
         \34245 , \34246 , \34247 , \34248 , \34249 , \34250 , \34251 , \34252 , \34253 , \34254 ,
         \34255 , \34256 , \34257 , \34258 , \34259 , \34260 , \34261 , \34262 , \34263 , \34264 ,
         \34265 , \34266 , \34267 , \34268 , \34269 , \34270 , \34271 , \34272 , \34273 , \34274 ,
         \34275 , \34276 , \34277 , \34278 , \34279 , \34280 , \34281 , \34282 , \34283 , \34284 ,
         \34285 , \34286 , \34287 , \34288 , \34289 , \34290 , \34291 , \34292 , \34293 , \34294 ,
         \34295 , \34296 , \34297 , \34298 , \34299 , \34300 , \34301 , \34302 , \34303 , \34304 ,
         \34305 , \34306 , \34307 , \34308 , \34309 , \34310 , \34311 , \34312 , \34313 , \34314 ,
         \34315 , \34316 , \34317 , \34318 , \34319 , \34320 , \34321 , \34322 , \34323 , \34324 ,
         \34325 , \34326 , \34327 , \34328 , \34329 , \34330 , \34331 , \34332 , \34333 , \34334 ,
         \34335 , \34336 , \34337 , \34338 , \34339 , \34340 , \34341 , \34342 , \34343 , \34344 ,
         \34345 , \34346 , \34347 , \34348 , \34349 , \34350 , \34351 , \34352 , \34353 , \34354 ,
         \34355 , \34356 , \34357 , \34358 , \34359 , \34360 , \34361 , \34362 , \34363 , \34364 ,
         \34365 , \34366 , \34367 , \34368 , \34369 , \34370 , \34371 , \34372 , \34373 , \34374 ,
         \34375 , \34376 , \34377 , \34378 , \34379 , \34380 , \34381 , \34382 , \34383 , \34384 ,
         \34385 , \34386 , \34387 , \34388 , \34389 , \34390 , \34391 , \34392 , \34393 , \34394 ,
         \34395 , \34396 , \34397 , \34398 , \34399 , \34400 , \34401 , \34402 , \34403 , \34404 ,
         \34405 , \34406 , \34407 , \34408 , \34409 , \34410 , \34411 , \34412 , \34413 , \34414 ,
         \34415 , \34416 , \34417 , \34418 , \34419 , \34420 , \34421 , \34422 , \34423 , \34424 ,
         \34425 , \34426 , \34427 , \34428 , \34429 , \34430 , \34431 , \34432 , \34433 , \34434 ,
         \34435 , \34436 , \34437 , \34438 , \34439 , \34440 , \34441 , \34442 , \34443 , \34444 ,
         \34445 , \34446 , \34447 , \34448 , \34449 , \34450 , \34451 , \34452 , \34453 , \34454 ,
         \34455 , \34456 , \34457 , \34458 , \34459 , \34460 , \34461 , \34462 , \34463 , \34464 ,
         \34465 , \34466 , \34467 , \34468 , \34469 , \34470 , \34471 , \34472 , \34473 , \34474 ,
         \34475 , \34476 , \34477 , \34478 , \34479 , \34480 , \34481 , \34482 , \34483 , \34484 ,
         \34485 , \34486 , \34487 , \34488 , \34489 , \34490 , \34491 , \34492 , \34493 , \34494 ,
         \34495 , \34496 , \34497 , \34498 , \34499 , \34500 , \34501 , \34502 , \34503 , \34504 ,
         \34505 , \34506 , \34507 , \34508 , \34509 , \34510 , \34511 , \34512 , \34513 , \34514 ,
         \34515 , \34516 , \34517 , \34518 , \34519 , \34520 , \34521 , \34522 , \34523 , \34524 ,
         \34525 , \34526 , \34527 , \34528 , \34529 , \34530 , \34531 , \34532 , \34533 , \34534 ,
         \34535 , \34536 , \34537 , \34538 , \34539 , \34540 , \34541 , \34542 , \34543 , \34544 ,
         \34545 , \34546 , \34547 , \34548 , \34549 , \34550 , \34551 , \34552 , \34553 , \34554 ,
         \34555 , \34556 , \34557 , \34558 , \34559 , \34560 , \34561 , \34562 , \34563 , \34564 ,
         \34565 , \34566 , \34567 , \34568 , \34569 , \34570 , \34571 , \34572 , \34573 , \34574 ,
         \34575 , \34576 , \34577 , \34578 , \34579 , \34580 , \34581 , \34582 , \34583 , \34584 ,
         \34585 , \34586 , \34587 , \34588 , \34589 , \34590 , \34591 , \34592 , \34593 , \34594 ,
         \34595 , \34596 , \34597 , \34598 , \34599 , \34600 , \34601 , \34602 , \34603 , \34604 ,
         \34605 , \34606 , \34607 , \34608 , \34609 , \34610 , \34611 , \34612 , \34613 , \34614 ,
         \34615 , \34616 , \34617 , \34618 , \34619 , \34620 , \34621 , \34622 , \34623 , \34624 ,
         \34625 , \34626 , \34627 , \34628 , \34629 , \34630 , \34631 , \34632 , \34633 , \34634 ,
         \34635 , \34636 , \34637 , \34638 , \34639 , \34640 , \34641 , \34642 , \34643 , \34644 ,
         \34645 , \34646 , \34647 , \34648 , \34649 , \34650 , \34651 , \34652 , \34653 , \34654 ,
         \34655 , \34656 , \34657 , \34658 , \34659 , \34660 , \34661 , \34662 , \34663 , \34664 ,
         \34665 , \34666 , \34667 , \34668 , \34669 , \34670 , \34671 , \34672 , \34673 , \34674 ,
         \34675 , \34676 , \34677 , \34678 , \34679 , \34680 , \34681 , \34682 , \34683 , \34684 ,
         \34685 , \34686 , \34687 , \34688 , \34689 , \34690 , \34691 , \34692 , \34693 , \34694 ,
         \34695 , \34696 , \34697 , \34698 , \34699 , \34700 , \34701 , \34702 , \34703 , \34704 ,
         \34705 , \34706 , \34707 , \34708 , \34709 , \34710 , \34711 , \34712 , \34713 , \34714 ,
         \34715 , \34716 , \34717 , \34718 , \34719 , \34720 , \34721 , \34722 , \34723 , \34724 ,
         \34725 , \34726 , \34727 , \34728 , \34729 , \34730 , \34731 , \34732 , \34733 , \34734 ,
         \34735 , \34736 , \34737 , \34738 , \34739 , \34740 , \34741 , \34742 , \34743 , \34744 ,
         \34745 , \34746 , \34747 , \34748 , \34749 , \34750 , \34751 , \34752 , \34753 , \34754 ,
         \34755 , \34756 , \34757 , \34758 , \34759 , \34760 , \34761 , \34762 , \34763 , \34764 ,
         \34765 , \34766 , \34767 , \34768 , \34769 , \34770 , \34771 , \34772 , \34773 , \34774 ,
         \34775 , \34776 , \34777 , \34778 , \34779 , \34780 , \34781 , \34782 , \34783 , \34784 ,
         \34785 , \34786 , \34787 , \34788 , \34789 , \34790 , \34791 , \34792 , \34793 , \34794 ,
         \34795 , \34796 , \34797 , \34798 , \34799 , \34800 , \34801 , \34802 , \34803 , \34804 ,
         \34805 , \34806 , \34807 , \34808 , \34809 , \34810 , \34811 , \34812 , \34813 , \34814 ,
         \34815 , \34816 , \34817 , \34818 , \34819 , \34820 , \34821 , \34822 , \34823 , \34824 ,
         \34825 , \34826 , \34827 , \34828 , \34829 , \34830 , \34831 , \34832 , \34833 , \34834 ,
         \34835 , \34836 , \34837 , \34838 , \34839 , \34840 , \34841 , \34842 , \34843 , \34844 ,
         \34845 , \34846 , \34847 , \34848 , \34849 , \34850 , \34851 , \34852 , \34853 , \34854 ,
         \34855 , \34856 , \34857 , \34858 , \34859 , \34860 , \34861 , \34862 , \34863 , \34864 ,
         \34865 , \34866 , \34867 , \34868 , \34869 , \34870 , \34871 , \34872 , \34873 , \34874 ,
         \34875 , \34876 , \34877 , \34878 , \34879 , \34880 , \34881 , \34882 , \34883 , \34884 ,
         \34885 , \34886 , \34887 , \34888 , \34889 , \34890 , \34891 , \34892 , \34893 , \34894 ,
         \34895 , \34896 , \34897 , \34898 , \34899 , \34900 , \34901 , \34902 , \34903 , \34904 ,
         \34905 , \34906 , \34907 , \34908 , \34909 , \34910 , \34911 , \34912 , \34913 , \34914 ,
         \34915 , \34916 , \34917 , \34918 , \34919 , \34920 , \34921 , \34922 , \34923 , \34924 ,
         \34925 , \34926 , \34927 , \34928 , \34929 , \34930 , \34931 , \34932 , \34933 , \34934 ,
         \34935 , \34936 , \34937 , \34938 , \34939 , \34940 , \34941 , \34942 , \34943 , \34944 ,
         \34945 , \34946 , \34947 , \34948 , \34949 , \34950 , \34951 , \34952 , \34953 , \34954 ,
         \34955 , \34956 , \34957 , \34958 , \34959 , \34960 , \34961 , \34962 , \34963 , \34964 ,
         \34965 , \34966 , \34967 , \34968 , \34969 , \34970 , \34971 , \34972 , \34973 , \34974 ,
         \34975 , \34976 , \34977 , \34978 , \34979 , \34980 , \34981 , \34982 , \34983 , \34984 ,
         \34985 , \34986 , \34987 , \34988 , \34989 , \34990 , \34991 , \34992 , \34993 , \34994 ,
         \34995 , \34996 , \34997 , \34998 , \34999 , \35000 , \35001 , \35002 , \35003 , \35004 ,
         \35005 , \35006 , \35007 , \35008 , \35009 , \35010 , \35011 , \35012 , \35013 , \35014 ,
         \35015 , \35016 , \35017 , \35018 , \35019 , \35020 , \35021 , \35022 , \35023 , \35024 ,
         \35025 , \35026 , \35027 , \35028 , \35029 , \35030 , \35031 , \35032 , \35033 , \35034 ,
         \35035 , \35036 , \35037 , \35038 , \35039 , \35040 , \35041 , \35042 , \35043 , \35044 ,
         \35045 , \35046 , \35047 , \35048 , \35049 , \35050 , \35051 , \35052 , \35053 , \35054 ,
         \35055 , \35056 , \35057 , \35058 , \35059 , \35060 , \35061 , \35062 , \35063 , \35064 ,
         \35065 , \35066 , \35067 , \35068 , \35069 , \35070 , \35071 , \35072 , \35073 , \35074 ,
         \35075 , \35076 , \35077 , \35078 , \35079 , \35080 , \35081 , \35082 , \35083 , \35084 ,
         \35085 , \35086 , \35087 , \35088 , \35089 , \35090 , \35091 , \35092 , \35093 , \35094 ,
         \35095 , \35096 , \35097 , \35098 , \35099 , \35100 , \35101 , \35102 , \35103 , \35104 ,
         \35105 , \35106 , \35107 , \35108 , \35109 , \35110 , \35111 , \35112 , \35113 , \35114 ,
         \35115 , \35116 , \35117 , \35118 , \35119 , \35120 , \35121 , \35122 , \35123 , \35124 ,
         \35125 , \35126 , \35127 , \35128 , \35129 , \35130 , \35131 , \35132 , \35133 , \35134 ,
         \35135 , \35136 , \35137 , \35138 , \35139 , \35140 , \35141 , \35142 , \35143 , \35144 ,
         \35145 , \35146 , \35147 , \35148 , \35149 , \35150 , \35151 , \35152 , \35153 , \35154 ,
         \35155 , \35156 , \35157 , \35158 , \35159 , \35160 , \35161 , \35162 , \35163 , \35164 ,
         \35165 , \35166 , \35167 , \35168 , \35169 , \35170 , \35171 , \35172 , \35173 , \35174 ,
         \35175 , \35176 , \35177 , \35178 , \35179 , \35180 , \35181 , \35182 , \35183 , \35184 ,
         \35185 , \35186 , \35187 , \35188 , \35189 , \35190 , \35191 , \35192 , \35193 , \35194 ,
         \35195 , \35196 , \35197 , \35198 , \35199 , \35200 , \35201 , \35202 , \35203 , \35204 ,
         \35205 , \35206 , \35207 , \35208 , \35209 , \35210 , \35211 , \35212 , \35213 , \35214 ,
         \35215 , \35216 , \35217 , \35218 , \35219 , \35220 , \35221 , \35222 , \35223 , \35224 ,
         \35225 , \35226 , \35227 , \35228 , \35229 , \35230 , \35231 , \35232 , \35233 , \35234 ,
         \35235 , \35236 , \35237 , \35238 , \35239 , \35240 , \35241 , \35242 , \35243 , \35244 ,
         \35245 , \35246 , \35247 , \35248 , \35249 , \35250 , \35251 , \35252 , \35253 , \35254 ,
         \35255 , \35256 , \35257 , \35258 , \35259 , \35260 , \35261 , \35262 , \35263 , \35264 ,
         \35265 , \35266 , \35267 , \35268 , \35269 , \35270 , \35271 , \35272 , \35273 , \35274 ,
         \35275 , \35276 , \35277 , \35278 , \35279 , \35280 , \35281 , \35282 , \35283 , \35284 ,
         \35285 , \35286 , \35287 , \35288 , \35289 , \35290 , \35291 , \35292 , \35293 , \35294 ,
         \35295 , \35296 , \35297 , \35298 , \35299 , \35300 , \35301 , \35302 , \35303 , \35304 ,
         \35305 , \35306 , \35307 , \35308 , \35309 , \35310 , \35311 , \35312 , \35313 , \35314 ,
         \35315 , \35316 , \35317 , \35318 , \35319 , \35320 , \35321 , \35322 , \35323 , \35324 ,
         \35325 , \35326 , \35327 , \35328 , \35329 , \35330 , \35331 , \35332 , \35333 , \35334 ,
         \35335 , \35336 , \35337 , \35338 , \35339 , \35340 , \35341 , \35342 , \35343 , \35344 ,
         \35345 , \35346 , \35347 , \35348 , \35349 , \35350 , \35351 , \35352 , \35353 , \35354 ,
         \35355 , \35356 , \35357 , \35358 , \35359 , \35360 , \35361 , \35362 , \35363 , \35364 ,
         \35365 , \35366 , \35367 , \35368 , \35369 , \35370 , \35371 , \35372 , \35373 , \35374 ,
         \35375 , \35376 , \35377 , \35378 , \35379 , \35380 , \35381 , \35382 , \35383 , \35384 ,
         \35385 , \35386 , \35387 , \35388 , \35389 , \35390 , \35391 , \35392 , \35393 , \35394 ,
         \35395 , \35396 , \35397 , \35398 , \35399 , \35400 , \35401 , \35402 , \35403 , \35404 ,
         \35405 , \35406 , \35407 , \35408 , \35409 , \35410 , \35411 , \35412 , \35413 , \35414 ,
         \35415 , \35416 , \35417 , \35418 , \35419 , \35420 , \35421 , \35422 , \35423 , \35424 ,
         \35425 , \35426 , \35427 , \35428 , \35429 , \35430 , \35431 , \35432 , \35433 , \35434 ,
         \35435 , \35436 , \35437 , \35438 , \35439 , \35440 , \35441 , \35442 , \35443 , \35444 ,
         \35445 , \35446 , \35447 , \35448 , \35449 , \35450 , \35451 , \35452 , \35453 , \35454 ,
         \35455 , \35456 , \35457 , \35458 , \35459 , \35460 , \35461 , \35462 , \35463 , \35464 ,
         \35465 , \35466 , \35467 , \35468 , \35469 , \35470 , \35471 , \35472 , \35473 , \35474 ,
         \35475 , \35476 , \35477 , \35478 , \35479 , \35480 , \35481 , \35482 , \35483 , \35484 ,
         \35485 , \35486 , \35487 , \35488 , \35489 , \35490 , \35491 , \35492 , \35493 , \35494 ,
         \35495 , \35496 , \35497 , \35498 , \35499 , \35500 , \35501 , \35502 , \35503 , \35504 ,
         \35505 , \35506 , \35507 , \35508 , \35509 , \35510 , \35511 , \35512 , \35513 , \35514 ,
         \35515 , \35516 , \35517 , \35518 , \35519 , \35520 , \35521 , \35522 , \35523 , \35524 ,
         \35525 , \35526 , \35527 , \35528 , \35529 , \35530 , \35531 , \35532 , \35533 , \35534 ,
         \35535 , \35536 , \35537 , \35538 , \35539 , \35540 , \35541 , \35542 , \35543 , \35544 ,
         \35545 , \35546 , \35547 , \35548 , \35549 , \35550 , \35551 , \35552 , \35553 , \35554 ,
         \35555 , \35556 , \35557 , \35558 , \35559 , \35560 , \35561 , \35562 , \35563 , \35564 ,
         \35565 , \35566 , \35567 , \35568 , \35569 , \35570 , \35571 , \35572 , \35573 , \35574 ,
         \35575 , \35576 , \35577 , \35578 , \35579 , \35580 , \35581 , \35582 , \35583 , \35584 ,
         \35585 , \35586 , \35587 , \35588 , \35589 , \35590 , \35591 , \35592 , \35593 , \35594 ,
         \35595 , \35596 , \35597 , \35598 , \35599 , \35600 , \35601 , \35602 , \35603 , \35604 ,
         \35605 , \35606 , \35607 , \35608 , \35609 , \35610 , \35611 , \35612 , \35613 , \35614 ,
         \35615 , \35616 , \35617 , \35618 , \35619 , \35620 , \35621 , \35622 , \35623 , \35624 ,
         \35625 , \35626 , \35627 , \35628 , \35629 , \35630 , \35631 , \35632 , \35633 , \35634 ,
         \35635 , \35636 , \35637 , \35638 , \35639 , \35640 , \35641 , \35642 , \35643 , \35644 ,
         \35645 , \35646 , \35647 , \35648 , \35649 , \35650 , \35651 , \35652 , \35653 , \35654 ,
         \35655 , \35656 , \35657 , \35658 , \35659 , \35660 , \35661 , \35662 , \35663 , \35664 ,
         \35665 , \35666 , \35667 , \35668 , \35669 , \35670 , \35671 , \35672 , \35673 , \35674 ,
         \35675 , \35676 , \35677 , \35678 , \35679 , \35680 , \35681 , \35682 , \35683 , \35684 ,
         \35685 , \35686 , \35687 , \35688 , \35689 , \35690 , \35691 , \35692 , \35693 , \35694 ,
         \35695 , \35696 , \35697 , \35698 , \35699 , \35700 , \35701 , \35702 , \35703 , \35704 ,
         \35705 , \35706 , \35707 , \35708 , \35709 , \35710 , \35711 , \35712 , \35713 , \35714 ,
         \35715 , \35716 , \35717 , \35718 , \35719 , \35720 , \35721 , \35722 , \35723 , \35724 ,
         \35725 , \35726 , \35727 , \35728 , \35729 , \35730 , \35731 , \35732 , \35733 , \35734 ,
         \35735 , \35736 , \35737 , \35738 , \35739 , \35740 , \35741 , \35742 , \35743 , \35744 ,
         \35745 , \35746 , \35747 , \35748 , \35749 , \35750 , \35751 , \35752 , \35753 , \35754 ,
         \35755 , \35756 , \35757 , \35758 , \35759 , \35760 , \35761 , \35762 , \35763 , \35764 ,
         \35765 , \35766 , \35767 , \35768 , \35769 , \35770 , \35771 , \35772 , \35773 , \35774 ,
         \35775 , \35776 , \35777 , \35778 , \35779 , \35780 , \35781 , \35782 , \35783 , \35784 ,
         \35785 , \35786 , \35787 , \35788 , \35789 , \35790 , \35791 , \35792 , \35793 , \35794 ,
         \35795 , \35796 , \35797 , \35798 , \35799 , \35800 , \35801 , \35802 , \35803 , \35804 ,
         \35805 , \35806 , \35807 , \35808 , \35809 , \35810 , \35811 , \35812 , \35813 , \35814 ,
         \35815 , \35816 , \35817 , \35818 , \35819 , \35820 , \35821 , \35822 , \35823 , \35824 ,
         \35825 , \35826 , \35827 , \35828 , \35829 , \35830 , \35831 , \35832 , \35833 , \35834 ,
         \35835 , \35836 , \35837 , \35838 , \35839 , \35840 , \35841 , \35842 , \35843 , \35844 ,
         \35845 , \35846 , \35847 , \35848 , \35849 , \35850 , \35851 , \35852 , \35853 , \35854 ,
         \35855 , \35856 , \35857 , \35858 , \35859 , \35860 , \35861 , \35862 , \35863 , \35864 ,
         \35865 , \35866 , \35867 , \35868 , \35869 , \35870 , \35871 , \35872 , \35873 , \35874 ,
         \35875 , \35876 , \35877 , \35878 , \35879 , \35880 , \35881 , \35882 , \35883 , \35884 ,
         \35885 , \35886 , \35887 , \35888 , \35889 , \35890 , \35891 , \35892 , \35893 , \35894 ,
         \35895 , \35896 , \35897 , \35898 , \35899 , \35900 , \35901 , \35902 , \35903 , \35904 ,
         \35905 , \35906 , \35907 , \35908 , \35909 , \35910 , \35911 , \35912 , \35913 , \35914 ,
         \35915 , \35916 , \35917 , \35918 , \35919 , \35920 , \35921 , \35922 , \35923 , \35924 ,
         \35925 , \35926 , \35927 , \35928 , \35929 , \35930 , \35931 , \35932 , \35933 , \35934 ,
         \35935 , \35936 , \35937 , \35938 , \35939 , \35940 , \35941 , \35942 , \35943 , \35944 ,
         \35945 , \35946 , \35947 , \35948 , \35949 , \35950 , \35951 , \35952 , \35953 , \35954 ,
         \35955 , \35956 , \35957 , \35958 , \35959 , \35960 , \35961 , \35962 , \35963 , \35964 ,
         \35965 , \35966 , \35967 , \35968 , \35969 , \35970 , \35971 , \35972 , \35973 , \35974 ,
         \35975 , \35976 , \35977 , \35978 , \35979 , \35980 , \35981 , \35982 , \35983 , \35984 ,
         \35985 , \35986 , \35987 , \35988 , \35989 , \35990 , \35991 , \35992 , \35993 , \35994 ,
         \35995 , \35996 , \35997 , \35998 , \35999 , \36000 , \36001 , \36002 , \36003 , \36004 ,
         \36005 , \36006 , \36007 , \36008 , \36009 , \36010 , \36011 , \36012 , \36013 , \36014 ,
         \36015 , \36016 , \36017 , \36018 , \36019 , \36020 , \36021 , \36022 , \36023 , \36024 ,
         \36025 , \36026 , \36027 , \36028 , \36029 , \36030 , \36031 , \36032 , \36033 , \36034 ,
         \36035 , \36036 , \36037 , \36038 , \36039 , \36040 , \36041 , \36042 , \36043 , \36044 ,
         \36045 , \36046 , \36047 , \36048 , \36049 , \36050 , \36051 , \36052 , \36053 , \36054 ,
         \36055 , \36056 , \36057 , \36058 , \36059 , \36060 , \36061 , \36062 , \36063 , \36064 ,
         \36065 , \36066 , \36067 , \36068 , \36069 , \36070 , \36071 , \36072 , \36073 , \36074 ,
         \36075 , \36076 , \36077 , \36078 , \36079 , \36080 , \36081 , \36082 , \36083 , \36084 ,
         \36085 , \36086 , \36087 , \36088 , \36089 , \36090 , \36091 , \36092 , \36093 , \36094 ,
         \36095 , \36096 , \36097 , \36098 , \36099 , \36100 , \36101 , \36102 , \36103 , \36104 ,
         \36105 , \36106 , \36107 , \36108 , \36109 , \36110 , \36111 , \36112 , \36113 , \36114 ,
         \36115 , \36116 , \36117 , \36118 , \36119 , \36120 , \36121 , \36122 , \36123 , \36124 ,
         \36125 , \36126 , \36127 , \36128 , \36129 , \36130 , \36131 , \36132 , \36133 , \36134 ,
         \36135 , \36136 , \36137 , \36138 , \36139 , \36140 , \36141 , \36142 , \36143 , \36144 ,
         \36145 , \36146 , \36147 , \36148 , \36149 , \36150 , \36151 , \36152 , \36153 , \36154 ,
         \36155 , \36156 , \36157 , \36158 , \36159 , \36160 , \36161 , \36162 , \36163 , \36164 ,
         \36165 , \36166 , \36167 , \36168 , \36169 , \36170 , \36171 , \36172 , \36173 , \36174 ,
         \36175 , \36176 , \36177 , \36178 , \36179 , \36180 , \36181 , \36182 , \36183 , \36184 ,
         \36185 , \36186 , \36187 , \36188 , \36189 , \36190 , \36191 , \36192 , \36193 , \36194 ,
         \36195 , \36196 , \36197 , \36198 , \36199 , \36200 , \36201 , \36202 , \36203 , \36204 ,
         \36205 , \36206 , \36207 , \36208 , \36209 , \36210 , \36211 , \36212 , \36213 , \36214 ,
         \36215 , \36216 , \36217 , \36218 , \36219 , \36220 , \36221 , \36222 , \36223 , \36224 ,
         \36225 , \36226 , \36227 , \36228 , \36229 , \36230 , \36231 , \36232 , \36233 , \36234 ,
         \36235 , \36236 , \36237 , \36238 , \36239 , \36240 , \36241 , \36242 , \36243 , \36244 ,
         \36245 , \36246 , \36247 , \36248 , \36249 , \36250 , \36251 , \36252 , \36253 , \36254 ,
         \36255 , \36256 , \36257 , \36258 , \36259 , \36260 , \36261 , \36262 , \36263 , \36264 ,
         \36265 , \36266 , \36267 , \36268 , \36269 , \36270 , \36271 , \36272 , \36273 , \36274 ,
         \36275 , \36276 , \36277 , \36278 , \36279 , \36280 , \36281 , \36282 , \36283 , \36284 ,
         \36285 , \36286 , \36287 , \36288 , \36289 , \36290 , \36291 , \36292 , \36293 , \36294 ,
         \36295 , \36296 , \36297 , \36298 , \36299 , \36300 , \36301 , \36302 , \36303 , \36304 ,
         \36305 , \36306 , \36307 , \36308 , \36309 , \36310 , \36311 , \36312 , \36313 , \36314 ,
         \36315 , \36316 , \36317 , \36318 , \36319 , \36320 , \36321 , \36322 , \36323 , \36324 ,
         \36325 , \36326 , \36327 , \36328 , \36329 , \36330 , \36331 , \36332 , \36333 , \36334 ,
         \36335 , \36336 , \36337 , \36338 , \36339 , \36340 , \36341 , \36342 , \36343 , \36344 ,
         \36345 , \36346 , \36347 , \36348 , \36349 , \36350 , \36351 , \36352 , \36353 , \36354 ,
         \36355 , \36356 , \36357 , \36358 , \36359 , \36360 , \36361 , \36362 , \36363 , \36364 ,
         \36365 , \36366 , \36367 , \36368 , \36369 , \36370 , \36371 , \36372 , \36373 , \36374 ,
         \36375 , \36376 , \36377 , \36378 , \36379 , \36380 , \36381 , \36382 , \36383 , \36384 ,
         \36385 , \36386 , \36387 , \36388 , \36389 , \36390 , \36391 , \36392 , \36393 , \36394 ,
         \36395 , \36396 , \36397 , \36398 , \36399 , \36400 , \36401 , \36402 , \36403 , \36404 ,
         \36405 , \36406 , \36407 , \36408 , \36409 , \36410 , \36411 , \36412 , \36413 , \36414 ,
         \36415 , \36416 , \36417 , \36418 , \36419 , \36420 , \36421 , \36422 , \36423 , \36424 ,
         \36425 , \36426 , \36427 , \36428 , \36429 , \36430 , \36431 , \36432 , \36433 , \36434 ,
         \36435 , \36436 , \36437 , \36438 , \36439 , \36440 , \36441 , \36442 , \36443 , \36444 ,
         \36445 , \36446 , \36447 , \36448 , \36449 , \36450 , \36451 , \36452 , \36453 , \36454 ,
         \36455 , \36456 , \36457 , \36458 , \36459 , \36460 , \36461 , \36462 , \36463 , \36464 ,
         \36465 , \36466 , \36467 , \36468 , \36469 , \36470 , \36471 , \36472 , \36473 , \36474 ,
         \36475 , \36476 , \36477 , \36478 , \36479 , \36480 , \36481 , \36482 , \36483 , \36484 ,
         \36485 , \36486 , \36487 , \36488 , \36489 , \36490 , \36491 , \36492 , \36493 , \36494 ,
         \36495 , \36496 , \36497 , \36498 , \36499 , \36500 , \36501 , \36502 , \36503 , \36504 ,
         \36505 , \36506 , \36507 , \36508 , \36509 , \36510 , \36511 , \36512 , \36513 , \36514 ,
         \36515 , \36516 , \36517 , \36518 , \36519 , \36520 , \36521 , \36522 , \36523 , \36524 ,
         \36525 , \36526 , \36527 , \36528 , \36529 , \36530 , \36531 , \36532 , \36533 , \36534 ,
         \36535 , \36536 , \36537 , \36538 , \36539 , \36540 , \36541 , \36542 , \36543 , \36544 ,
         \36545 , \36546 , \36547 , \36548 , \36549 , \36550 , \36551 , \36552 , \36553 , \36554 ,
         \36555 , \36556 , \36557 , \36558 , \36559 , \36560 , \36561 , \36562 , \36563 , \36564 ,
         \36565 , \36566 , \36567 , \36568 , \36569 , \36570 , \36571 , \36572 , \36573 , \36574 ,
         \36575 , \36576 , \36577 , \36578 , \36579 , \36580 , \36581 , \36582 , \36583 , \36584 ,
         \36585 , \36586 , \36587 , \36588 , \36589 , \36590 , \36591 , \36592 , \36593 , \36594 ,
         \36595 , \36596 , \36597 , \36598 , \36599 , \36600 , \36601 , \36602 , \36603 , \36604 ,
         \36605 , \36606 , \36607 , \36608 , \36609 , \36610 , \36611 , \36612 , \36613 , \36614 ,
         \36615 , \36616 , \36617 , \36618 , \36619 , \36620 , \36621 , \36622 , \36623 , \36624 ,
         \36625 , \36626 , \36627 , \36628 , \36629 , \36630 , \36631 , \36632 , \36633 , \36634 ,
         \36635 , \36636 , \36637 , \36638 , \36639 , \36640 , \36641 , \36642 , \36643 , \36644 ,
         \36645 , \36646 , \36647 , \36648 , \36649 , \36650 , \36651 , \36652 , \36653 , \36654 ,
         \36655 , \36656 , \36657 , \36658 , \36659 , \36660 , \36661 , \36662 , \36663 , \36664 ,
         \36665 , \36666 , \36667 , \36668 , \36669 , \36670 , \36671 , \36672 , \36673 , \36674 ,
         \36675 , \36676 , \36677 , \36678 , \36679 , \36680 , \36681 , \36682 , \36683 , \36684 ,
         \36685 , \36686 , \36687 , \36688 , \36689 , \36690 , \36691 , \36692 , \36693 , \36694 ,
         \36695 , \36696 , \36697 , \36698 , \36699 , \36700 , \36701 , \36702 , \36703 , \36704 ,
         \36705 , \36706 , \36707 , \36708 , \36709 , \36710 , \36711 , \36712 , \36713 , \36714 ,
         \36715 , \36716 , \36717 , \36718 , \36719 , \36720 , \36721 , \36722 , \36723 , \36724 ,
         \36725 , \36726 , \36727 , \36728 , \36729 , \36730 , \36731 , \36732 , \36733 , \36734 ,
         \36735 , \36736 , \36737 , \36738 , \36739 , \36740 , \36741 , \36742 , \36743 , \36744 ,
         \36745 , \36746 , \36747 , \36748 , \36749 , \36750 , \36751 , \36752 , \36753 , \36754 ,
         \36755 , \36756 , \36757 , \36758 , \36759 , \36760 , \36761 , \36762 , \36763 , \36764 ,
         \36765 , \36766 , \36767 , \36768 , \36769 , \36770 , \36771 , \36772 , \36773 , \36774 ,
         \36775 , \36776 , \36777 , \36778 , \36779 , \36780 , \36781 , \36782 , \36783 , \36784 ,
         \36785 , \36786 , \36787 , \36788 , \36789 , \36790 , \36791 , \36792 , \36793 , \36794 ,
         \36795 , \36796 , \36797 , \36798 , \36799 , \36800 , \36801 , \36802 , \36803 , \36804 ,
         \36805 , \36806 , \36807 , \36808 , \36809 , \36810 , \36811 , \36812 , \36813 , \36814 ,
         \36815 , \36816 , \36817 , \36818 , \36819 , \36820 , \36821 , \36822 , \36823 , \36824 ,
         \36825 , \36826 , \36827 , \36828 , \36829 , \36830 , \36831 , \36832 , \36833 , \36834 ,
         \36835 , \36836 , \36837 , \36838 , \36839 , \36840 , \36841 , \36842 , \36843 , \36844 ,
         \36845 , \36846 , \36847 , \36848 , \36849 , \36850 , \36851 , \36852 , \36853 , \36854 ,
         \36855 , \36856 , \36857 , \36858 , \36859 , \36860 , \36861 , \36862 , \36863 , \36864 ,
         \36865 , \36866 , \36867 , \36868 , \36869 , \36870 , \36871 , \36872 , \36873 , \36874 ,
         \36875 , \36876 , \36877 , \36878 , \36879 , \36880 , \36881 , \36882 , \36883 , \36884 ,
         \36885 , \36886 , \36887 , \36888 , \36889 , \36890 , \36891 , \36892 , \36893 , \36894 ,
         \36895 , \36896 , \36897 , \36898 , \36899 , \36900 , \36901 , \36902 , \36903 , \36904 ,
         \36905 , \36906 , \36907 , \36908 , \36909 , \36910 , \36911 , \36912 , \36913 , \36914 ,
         \36915 , \36916 , \36917 , \36918 , \36919 , \36920 , \36921 , \36922 , \36923 , \36924 ,
         \36925 , \36926 , \36927 , \36928 , \36929 , \36930 , \36931 , \36932 , \36933 , \36934 ,
         \36935 , \36936 , \36937 , \36938 , \36939 , \36940 , \36941 , \36942 , \36943 , \36944 ,
         \36945 , \36946 , \36947 , \36948 , \36949 , \36950 , \36951 , \36952 , \36953 , \36954 ,
         \36955 , \36956 , \36957 , \36958 , \36959 , \36960 , \36961 , \36962 , \36963 , \36964 ,
         \36965 , \36966 , \36967 , \36968 , \36969 , \36970 , \36971 , \36972 , \36973 , \36974 ,
         \36975 , \36976 , \36977 , \36978 , \36979 , \36980 , \36981 , \36982 , \36983 , \36984 ,
         \36985 , \36986 , \36987 , \36988 , \36989 , \36990 , \36991 , \36992 , \36993 , \36994 ,
         \36995 , \36996 , \36997 , \36998 , \36999 , \37000 , \37001 , \37002 , \37003 , \37004 ,
         \37005 , \37006 , \37007 , \37008 , \37009 , \37010 , \37011 , \37012 , \37013 , \37014 ,
         \37015 , \37016 , \37017 , \37018 , \37019 , \37020 , \37021 , \37022 , \37023 , \37024 ,
         \37025 , \37026 , \37027 , \37028 , \37029 , \37030 , \37031 , \37032 , \37033 , \37034 ,
         \37035 , \37036 , \37037 , \37038 , \37039 , \37040 , \37041 , \37042 , \37043 , \37044 ,
         \37045 , \37046 , \37047 , \37048 , \37049 , \37050 , \37051 , \37052 , \37053 , \37054 ,
         \37055 , \37056 , \37057 , \37058 , \37059 , \37060 , \37061 , \37062 , \37063 , \37064 ,
         \37065 , \37066 , \37067 , \37068 , \37069 , \37070 , \37071 , \37072 , \37073 , \37074 ,
         \37075 , \37076 , \37077 , \37078 , \37079 , \37080 , \37081 , \37082 , \37083 , \37084 ,
         \37085 , \37086 , \37087 , \37088 , \37089 , \37090 , \37091 , \37092 , \37093 , \37094 ,
         \37095 , \37096 , \37097 , \37098 , \37099 , \37100 , \37101 , \37102 , \37103 , \37104 ,
         \37105 , \37106 , \37107 , \37108 , \37109 , \37110 , \37111 , \37112 , \37113 , \37114 ,
         \37115 , \37116 , \37117 , \37118 , \37119 , \37120 , \37121 , \37122 , \37123 , \37124 ,
         \37125 , \37126 , \37127 , \37128 , \37129 , \37130 , \37131 , \37132 , \37133 , \37134 ,
         \37135 , \37136 , \37137 , \37138 , \37139 , \37140 , \37141 , \37142 , \37143 , \37144 ,
         \37145 , \37146 , \37147 , \37148 , \37149 , \37150 , \37151 , \37152 , \37153 , \37154 ,
         \37155 , \37156 , \37157 , \37158 , \37159 , \37160 , \37161 , \37162 , \37163 , \37164 ,
         \37165 , \37166 , \37167 , \37168 , \37169 , \37170 , \37171 , \37172 , \37173 , \37174 ,
         \37175 , \37176 , \37177 , \37178 , \37179 , \37180 , \37181 , \37182 , \37183 , \37184 ,
         \37185 , \37186 , \37187 , \37188 , \37189 , \37190 , \37191 , \37192 , \37193 , \37194 ,
         \37195 , \37196 , \37197 , \37198 , \37199 , \37200 , \37201 , \37202 , \37203 , \37204 ,
         \37205 , \37206 , \37207 , \37208 , \37209 , \37210 , \37211 , \37212 , \37213 , \37214 ,
         \37215 , \37216 , \37217 , \37218 , \37219 , \37220 , \37221 , \37222 , \37223 , \37224 ,
         \37225 , \37226 , \37227 , \37228 , \37229 , \37230 , \37231 , \37232 , \37233 , \37234 ,
         \37235 , \37236 , \37237 , \37238 , \37239 , \37240 , \37241 , \37242 , \37243 , \37244 ,
         \37245 , \37246 , \37247 , \37248 , \37249 , \37250 , \37251 , \37252 , \37253 , \37254 ,
         \37255 , \37256 , \37257 , \37258 , \37259 , \37260 , \37261 , \37262 , \37263 , \37264 ,
         \37265 , \37266 , \37267 , \37268 , \37269 , \37270 , \37271 , \37272 , \37273 , \37274 ,
         \37275 , \37276 , \37277 , \37278 , \37279 , \37280 , \37281 , \37282 , \37283 , \37284 ,
         \37285 , \37286 , \37287 , \37288 , \37289 , \37290 , \37291 , \37292 , \37293 , \37294 ,
         \37295 , \37296 , \37297 , \37298 , \37299 , \37300 , \37301 , \37302 , \37303 , \37304 ,
         \37305 , \37306 , \37307 , \37308 , \37309 , \37310 , \37311 , \37312 , \37313 , \37314 ,
         \37315 , \37316 , \37317 , \37318 , \37319 , \37320 , \37321 , \37322 , \37323 , \37324 ,
         \37325 , \37326 , \37327 , \37328 , \37329 , \37330 , \37331 , \37332 , \37333 , \37334 ,
         \37335 , \37336 , \37337 , \37338 , \37339 , \37340 , \37341 , \37342 , \37343 , \37344 ,
         \37345 , \37346 , \37347 , \37348 , \37349 , \37350 , \37351 , \37352 , \37353 , \37354 ,
         \37355 , \37356 , \37357 , \37358 , \37359 , \37360 , \37361 , \37362 , \37363 , \37364 ,
         \37365 , \37366 , \37367 , \37368 , \37369 , \37370 , \37371 , \37372 , \37373 , \37374 ,
         \37375 , \37376 , \37377 , \37378 , \37379 , \37380 , \37381 , \37382 , \37383 , \37384 ,
         \37385 , \37386 , \37387 , \37388 , \37389 , \37390 , \37391 , \37392 , \37393 , \37394 ,
         \37395 , \37396 , \37397 , \37398 , \37399 , \37400 , \37401 , \37402 , \37403 , \37404 ,
         \37405 , \37406 , \37407 , \37408 , \37409 , \37410 , \37411 , \37412 , \37413 , \37414 ,
         \37415 , \37416 , \37417 , \37418 , \37419 , \37420 , \37421 , \37422 , \37423 , \37424 ,
         \37425 , \37426 , \37427 , \37428 , \37429 , \37430 , \37431 , \37432 , \37433 , \37434 ,
         \37435 , \37436 , \37437 , \37438 , \37439 , \37440 , \37441 , \37442 , \37443 , \37444 ,
         \37445 , \37446 , \37447 , \37448 , \37449 , \37450 , \37451 , \37452 , \37453 , \37454 ,
         \37455 , \37456 , \37457 , \37458 , \37459 , \37460 , \37461 , \37462 , \37463 , \37464 ,
         \37465 , \37466 , \37467 , \37468 , \37469 , \37470 , \37471 , \37472 , \37473 , \37474 ,
         \37475 , \37476 , \37477 , \37478 , \37479 , \37480 , \37481 , \37482 , \37483 , \37484 ,
         \37485 , \37486 , \37487 , \37488 , \37489 , \37490 , \37491 , \37492 , \37493 , \37494 ,
         \37495 , \37496 , \37497 , \37498 , \37499 , \37500 , \37501 , \37502 , \37503 , \37504 ,
         \37505 , \37506 , \37507 , \37508 , \37509 , \37510 , \37511 , \37512 , \37513 , \37514 ,
         \37515 , \37516 , \37517 , \37518 , \37519 , \37520 , \37521 , \37522 , \37523 , \37524 ,
         \37525 , \37526 , \37527 , \37528 , \37529 , \37530 , \37531 , \37532 , \37533 , \37534 ,
         \37535 , \37536 , \37537 , \37538 , \37539 , \37540 , \37541 , \37542 , \37543 , \37544 ,
         \37545 , \37546 , \37547 , \37548 , \37549 , \37550 , \37551 , \37552 , \37553 , \37554 ,
         \37555 , \37556 , \37557 , \37558 , \37559 , \37560 , \37561 , \37562 , \37563 , \37564 ,
         \37565 , \37566 , \37567 , \37568 , \37569 , \37570 , \37571 , \37572 , \37573 , \37574 ,
         \37575 , \37576 , \37577 , \37578 , \37579 , \37580 , \37581 , \37582 , \37583 , \37584 ,
         \37585 , \37586 , \37587 , \37588 , \37589 , \37590 , \37591 , \37592 , \37593 , \37594 ,
         \37595 , \37596 , \37597 , \37598 , \37599 , \37600 , \37601 , \37602 , \37603 , \37604 ,
         \37605 , \37606 , \37607 , \37608 , \37609 , \37610 , \37611 , \37612 , \37613 , \37614 ,
         \37615 , \37616 , \37617 , \37618 , \37619 , \37620 , \37621 , \37622 , \37623 , \37624 ,
         \37625 , \37626 , \37627 , \37628 , \37629 , \37630 , \37631 , \37632 , \37633 , \37634 ,
         \37635 , \37636 , \37637 , \37638 , \37639 , \37640 , \37641 , \37642 , \37643 , \37644 ,
         \37645 , \37646 , \37647 , \37648 , \37649 , \37650 , \37651 , \37652 , \37653 , \37654 ,
         \37655 , \37656 , \37657 , \37658 , \37659 , \37660 , \37661 , \37662 , \37663 , \37664 ,
         \37665 , \37666 , \37667 , \37668 , \37669 , \37670 , \37671 , \37672 , \37673 , \37674 ,
         \37675 , \37676 , \37677 , \37678 , \37679 , \37680 , \37681 , \37682 , \37683 , \37684 ,
         \37685 , \37686 , \37687 , \37688 , \37689 , \37690 , \37691 , \37692 , \37693 , \37694 ,
         \37695 , \37696 , \37697 , \37698 , \37699 , \37700 , \37701 , \37702 , \37703 , \37704 ,
         \37705 , \37706 , \37707 , \37708 , \37709 , \37710 , \37711 , \37712 , \37713 , \37714 ,
         \37715 , \37716 , \37717 , \37718 , \37719 , \37720 , \37721 , \37722 , \37723 , \37724 ,
         \37725 , \37726 , \37727 , \37728 , \37729 , \37730 , \37731 , \37732 , \37733 , \37734 ,
         \37735 , \37736 , \37737 , \37738 , \37739 , \37740 , \37741 , \37742 , \37743 , \37744 ,
         \37745 , \37746 , \37747 , \37748 , \37749 , \37750 , \37751 , \37752 , \37753 , \37754 ,
         \37755 , \37756 , \37757 , \37758 , \37759 , \37760 , \37761 , \37762 , \37763 , \37764 ,
         \37765 , \37766 , \37767 , \37768 , \37769 , \37770 , \37771 , \37772 , \37773 , \37774 ,
         \37775 , \37776 , \37777 , \37778 , \37779 , \37780 , \37781 , \37782 , \37783 , \37784 ,
         \37785 , \37786 , \37787 , \37788 , \37789 , \37790 , \37791 , \37792 , \37793 , \37794 ,
         \37795 , \37796 , \37797 , \37798 , \37799 , \37800 , \37801 , \37802 , \37803 , \37804 ,
         \37805 , \37806 , \37807 , \37808 , \37809 , \37810 , \37811 , \37812 , \37813 , \37814 ,
         \37815 , \37816 , \37817 , \37818 , \37819 , \37820 , \37821 , \37822 , \37823 , \37824 ,
         \37825 , \37826 , \37827 , \37828 , \37829 , \37830 , \37831 , \37832 , \37833 , \37834 ,
         \37835 , \37836 , \37837 , \37838 , \37839 , \37840 , \37841 , \37842 , \37843 , \37844 ,
         \37845 , \37846 , \37847 , \37848 , \37849 , \37850 , \37851 , \37852 , \37853 , \37854 ,
         \37855 , \37856 , \37857 , \37858 , \37859 , \37860 , \37861 , \37862 , \37863 , \37864 ,
         \37865 , \37866 , \37867 , \37868 , \37869 , \37870 , \37871 , \37872 , \37873 , \37874 ,
         \37875 , \37876 , \37877 , \37878 , \37879 , \37880 , \37881 , \37882 , \37883 , \37884 ,
         \37885 , \37886 , \37887 , \37888 , \37889 , \37890 , \37891 , \37892 , \37893 , \37894 ,
         \37895 , \37896 , \37897 , \37898 , \37899 , \37900 , \37901 , \37902 , \37903 , \37904 ,
         \37905 , \37906 , \37907 , \37908 , \37909 , \37910 , \37911 , \37912 , \37913 , \37914 ,
         \37915 , \37916 , \37917 , \37918 , \37919 , \37920 , \37921 , \37922 , \37923 , \37924 ,
         \37925 , \37926 , \37927 , \37928 , \37929 , \37930 , \37931 , \37932 , \37933 , \37934 ,
         \37935 , \37936 , \37937 , \37938 , \37939 , \37940 , \37941 , \37942 , \37943 , \37944 ,
         \37945 , \37946 , \37947 , \37948 , \37949 , \37950 , \37951 , \37952 , \37953 , \37954 ,
         \37955 , \37956 , \37957 , \37958 , \37959 , \37960 , \37961 , \37962 , \37963 , \37964 ,
         \37965 , \37966 , \37967 , \37968 , \37969 , \37970 , \37971 , \37972 , \37973 , \37974 ,
         \37975 , \37976 , \37977 , \37978 , \37979 , \37980 , \37981 , \37982 , \37983 , \37984 ,
         \37985 , \37986 , \37987 , \37988 , \37989 , \37990 , \37991 , \37992 , \37993 , \37994 ,
         \37995 , \37996 , \37997 , \37998 , \37999 , \38000 , \38001 , \38002 , \38003 , \38004 ,
         \38005 , \38006 , \38007 , \38008 , \38009 , \38010 , \38011 , \38012 , \38013 , \38014 ,
         \38015 , \38016 , \38017 , \38018 , \38019 , \38020 , \38021 , \38022 , \38023 , \38024 ,
         \38025 , \38026 , \38027 , \38028 , \38029 , \38030 , \38031 , \38032 , \38033 , \38034 ,
         \38035 , \38036 , \38037 , \38038 , \38039 , \38040 , \38041 , \38042 , \38043 , \38044 ,
         \38045 , \38046 , \38047 , \38048 , \38049 , \38050 , \38051 , \38052 , \38053 , \38054 ,
         \38055 , \38056 , \38057 , \38058 , \38059 , \38060 , \38061 , \38062 , \38063 , \38064 ,
         \38065 , \38066 , \38067 , \38068 , \38069 , \38070 , \38071 , \38072 , \38073 , \38074 ,
         \38075 , \38076 , \38077 , \38078 , \38079 , \38080 , \38081 , \38082 , \38083 , \38084 ,
         \38085 , \38086 , \38087 , \38088 , \38089 , \38090 , \38091 , \38092 , \38093 , \38094 ,
         \38095 , \38096 , \38097 , \38098 , \38099 , \38100 , \38101 , \38102 , \38103 , \38104 ,
         \38105 , \38106 , \38107 , \38108 , \38109 , \38110 , \38111 , \38112 , \38113 , \38114 ,
         \38115 , \38116 , \38117 , \38118 , \38119 , \38120 , \38121 , \38122 , \38123 , \38124 ,
         \38125 , \38126 , \38127 , \38128 , \38129 , \38130 , \38131 , \38132 , \38133 , \38134 ,
         \38135 , \38136 , \38137 , \38138 , \38139 , \38140 , \38141 , \38142 , \38143 , \38144 ,
         \38145 , \38146 , \38147 , \38148 , \38149 , \38150 , \38151 , \38152 , \38153 , \38154 ,
         \38155 , \38156 , \38157 , \38158 , \38159 , \38160 , \38161 , \38162 , \38163 , \38164 ,
         \38165 , \38166 , \38167 , \38168 , \38169 , \38170 , \38171 , \38172 , \38173 , \38174 ,
         \38175 , \38176 , \38177 , \38178 , \38179 , \38180 , \38181 , \38182 , \38183 , \38184 ,
         \38185 , \38186 , \38187 , \38188 , \38189 , \38190 , \38191 , \38192 , \38193 , \38194 ,
         \38195 , \38196 , \38197 , \38198 , \38199 , \38200 , \38201 , \38202 , \38203 , \38204 ,
         \38205 , \38206 , \38207 , \38208 , \38209 , \38210 , \38211 , \38212 , \38213 , \38214 ,
         \38215 , \38216 , \38217 , \38218 , \38219 , \38220 , \38221 , \38222 , \38223 , \38224 ,
         \38225 , \38226 , \38227 , \38228 , \38229 , \38230 , \38231 , \38232 , \38233 , \38234 ,
         \38235 , \38236 , \38237 , \38238 , \38239 , \38240 , \38241 , \38242 , \38243 , \38244 ,
         \38245 , \38246 , \38247 , \38248 , \38249 , \38250 , \38251 , \38252 , \38253 , \38254 ,
         \38255 , \38256 , \38257 , \38258 , \38259 , \38260 , \38261 , \38262 , \38263 , \38264 ,
         \38265 , \38266 , \38267 , \38268 , \38269 , \38270 , \38271 , \38272 , \38273 , \38274 ,
         \38275 , \38276 , \38277 , \38278 , \38279 , \38280 , \38281 , \38282 , \38283 , \38284 ,
         \38285 , \38286 , \38287 , \38288 , \38289 , \38290 , \38291 , \38292 , \38293 , \38294 ,
         \38295 , \38296 , \38297 , \38298 , \38299 , \38300 , \38301 , \38302 , \38303 , \38304 ,
         \38305 , \38306 , \38307 , \38308 , \38309 , \38310 , \38311 , \38312 , \38313 , \38314 ,
         \38315 , \38316 , \38317 , \38318 , \38319 , \38320 , \38321 , \38322 , \38323 , \38324 ,
         \38325 , \38326 , \38327 , \38328 , \38329 , \38330 , \38331 , \38332 , \38333 , \38334 ,
         \38335 , \38336 , \38337 , \38338 , \38339 , \38340 , \38341 , \38342 , \38343 , \38344 ,
         \38345 , \38346 , \38347 , \38348 , \38349 , \38350 , \38351 , \38352 , \38353 , \38354 ,
         \38355 , \38356 , \38357 , \38358 , \38359 , \38360 , \38361 , \38362 , \38363 , \38364 ,
         \38365 , \38366 , \38367 , \38368 , \38369 , \38370 , \38371 , \38372 , \38373 , \38374 ,
         \38375 , \38376 , \38377 , \38378 , \38379 , \38380 , \38381 , \38382 , \38383 , \38384 ,
         \38385 , \38386 , \38387 , \38388 , \38389 , \38390 , \38391 , \38392 , \38393 , \38394 ,
         \38395 , \38396 , \38397 , \38398 , \38399 , \38400 , \38401 , \38402 , \38403 , \38404 ,
         \38405 , \38406 , \38407 , \38408 , \38409 , \38410 , \38411 , \38412 , \38413 , \38414 ,
         \38415 , \38416 , \38417 , \38418 , \38419 , \38420 , \38421 , \38422 , \38423 , \38424 ,
         \38425 , \38426 , \38427 , \38428 , \38429 , \38430 , \38431 , \38432 , \38433 , \38434 ,
         \38435 , \38436 , \38437 , \38438 , \38439 , \38440 , \38441 , \38442 , \38443 , \38444 ,
         \38445 , \38446 , \38447 , \38448 , \38449 , \38450 , \38451 , \38452 , \38453 , \38454 ,
         \38455 , \38456 , \38457 , \38458 , \38459 , \38460 , \38461 , \38462 , \38463 , \38464 ,
         \38465 , \38466 , \38467 , \38468 , \38469 , \38470 , \38471 , \38472 , \38473 , \38474 ,
         \38475 , \38476 , \38477 , \38478 , \38479 , \38480 , \38481 , \38482 , \38483 , \38484 ,
         \38485 , \38486 , \38487 , \38488 , \38489 , \38490 , \38491 , \38492 , \38493 , \38494 ,
         \38495 , \38496 , \38497 , \38498 , \38499 , \38500 , \38501 , \38502 , \38503 , \38504 ,
         \38505 , \38506 , \38507 , \38508 , \38509 , \38510 , \38511 , \38512 , \38513 , \38514 ,
         \38515 , \38516 , \38517 , \38518 , \38519 , \38520 , \38521 , \38522 , \38523 , \38524 ,
         \38525 , \38526 , \38527 , \38528 , \38529 , \38530 , \38531 , \38532 , \38533 , \38534 ,
         \38535 , \38536 , \38537 , \38538 , \38539 , \38540 , \38541 , \38542 , \38543 , \38544 ,
         \38545 , \38546 , \38547 , \38548 , \38549 , \38550 , \38551 , \38552 , \38553 , \38554 ,
         \38555 , \38556 , \38557 , \38558 , \38559 , \38560 , \38561 , \38562 , \38563 , \38564 ,
         \38565 , \38566 , \38567 , \38568 , \38569 , \38570 , \38571 , \38572 , \38573 , \38574 ,
         \38575 , \38576 , \38577 , \38578 , \38579 , \38580 , \38581 , \38582 , \38583 , \38584 ,
         \38585 , \38586 , \38587 , \38588 , \38589 , \38590 , \38591 , \38592 , \38593 , \38594 ,
         \38595 , \38596 , \38597 , \38598 , \38599 , \38600 , \38601 , \38602 , \38603 , \38604 ,
         \38605 , \38606 , \38607 , \38608 , \38609 , \38610 , \38611 , \38612 , \38613 , \38614 ,
         \38615 , \38616 , \38617 , \38618 , \38619 , \38620 , \38621 , \38622 , \38623 , \38624 ,
         \38625 , \38626 , \38627 , \38628 , \38629 , \38630 , \38631 , \38632 , \38633 , \38634 ,
         \38635 , \38636 , \38637 , \38638 , \38639 , \38640 , \38641 , \38642 , \38643 , \38644 ,
         \38645 , \38646 , \38647 , \38648 , \38649 , \38650 , \38651 , \38652 , \38653 , \38654 ,
         \38655 , \38656 , \38657 , \38658 , \38659 , \38660 , \38661 , \38662 , \38663 , \38664 ,
         \38665 , \38666 , \38667 , \38668 , \38669 , \38670 , \38671 , \38672 , \38673 , \38674 ,
         \38675 , \38676 , \38677 , \38678 , \38679 , \38680 , \38681 , \38682 , \38683 , \38684 ,
         \38685 , \38686 , \38687 , \38688 , \38689 , \38690 , \38691 , \38692 , \38693 , \38694 ,
         \38695 , \38696 , \38697 , \38698 , \38699 , \38700 , \38701 , \38702 , \38703 , \38704 ,
         \38705 , \38706 , \38707 , \38708 , \38709 , \38710 , \38711 , \38712 , \38713 , \38714 ,
         \38715 , \38716 , \38717 , \38718 , \38719 , \38720 , \38721 , \38722 , \38723 , \38724 ,
         \38725 , \38726 , \38727 , \38728 , \38729 , \38730 , \38731 , \38732 , \38733 , \38734 ,
         \38735 , \38736 , \38737 , \38738 , \38739 , \38740 , \38741 , \38742 , \38743 , \38744 ,
         \38745 , \38746 , \38747 , \38748 , \38749 , \38750 , \38751 , \38752 , \38753 , \38754 ,
         \38755 , \38756 , \38757 , \38758 , \38759 , \38760 , \38761 , \38762 , \38763 , \38764 ,
         \38765 , \38766 , \38767 , \38768 , \38769 , \38770 , \38771 , \38772 , \38773 , \38774 ,
         \38775 , \38776 , \38777 , \38778 , \38779 , \38780 , \38781 , \38782 , \38783 , \38784 ,
         \38785 , \38786 , \38787 , \38788 , \38789 , \38790 , \38791 , \38792 , \38793 , \38794 ,
         \38795 , \38796 , \38797 , \38798 , \38799 , \38800 , \38801 , \38802 , \38803 , \38804 ,
         \38805 , \38806 , \38807 , \38808 , \38809 , \38810 , \38811 , \38812 , \38813 , \38814 ,
         \38815 , \38816 , \38817 , \38818 , \38819 , \38820 , \38821 , \38822 , \38823 , \38824 ,
         \38825 , \38826 , \38827 , \38828 , \38829 , \38830 , \38831 , \38832 , \38833 , \38834 ,
         \38835 , \38836 , \38837 , \38838 , \38839 , \38840 , \38841 , \38842 , \38843 , \38844 ,
         \38845 , \38846 , \38847 , \38848 , \38849 , \38850 , \38851 , \38852 , \38853 , \38854 ,
         \38855 , \38856 , \38857 , \38858 , \38859 , \38860 , \38861 , \38862 , \38863 , \38864 ,
         \38865 , \38866 , \38867 , \38868 , \38869 , \38870 , \38871 , \38872 , \38873 , \38874 ,
         \38875 , \38876 , \38877 , \38878 , \38879 , \38880 , \38881 , \38882 , \38883 , \38884 ,
         \38885 , \38886 , \38887 , \38888 , \38889 , \38890 , \38891 , \38892 , \38893 , \38894 ,
         \38895 , \38896 , \38897 , \38898 , \38899 , \38900 , \38901 , \38902 , \38903 , \38904 ,
         \38905 , \38906 , \38907 , \38908 , \38909 , \38910 , \38911 , \38912 , \38913 , \38914 ,
         \38915 , \38916 , \38917 , \38918 , \38919 , \38920 , \38921 , \38922 , \38923 , \38924 ,
         \38925 , \38926 , \38927 , \38928 , \38929 , \38930 , \38931 , \38932 , \38933 , \38934 ,
         \38935 , \38936 , \38937 , \38938 , \38939 , \38940 , \38941 , \38942 , \38943 , \38944 ,
         \38945 , \38946 , \38947 , \38948 , \38949 , \38950 , \38951 , \38952 , \38953 , \38954 ,
         \38955 , \38956 , \38957 , \38958 , \38959 , \38960 , \38961 , \38962 , \38963 , \38964 ,
         \38965 , \38966 , \38967 , \38968 , \38969 , \38970 , \38971 , \38972 , \38973 , \38974 ,
         \38975 , \38976 , \38977 , \38978 , \38979 , \38980 , \38981 , \38982 , \38983 , \38984 ,
         \38985 , \38986 , \38987 , \38988 , \38989 , \38990 , \38991 , \38992 , \38993 , \38994 ,
         \38995 , \38996 , \38997 , \38998 , \38999 , \39000 , \39001 , \39002 , \39003 , \39004 ,
         \39005 , \39006 , \39007 , \39008 , \39009 , \39010 , \39011 , \39012 , \39013 , \39014 ,
         \39015 , \39016 , \39017 , \39018 , \39019 , \39020 , \39021 , \39022 , \39023 , \39024 ,
         \39025 , \39026 , \39027 , \39028 , \39029 , \39030 , \39031 , \39032 , \39033 , \39034 ,
         \39035 , \39036 , \39037 , \39038 , \39039 , \39040 , \39041 , \39042 , \39043 , \39044 ,
         \39045 , \39046 , \39047 , \39048 , \39049 , \39050 , \39051 , \39052 , \39053 , \39054 ,
         \39055 , \39056 , \39057 , \39058 , \39059 , \39060 , \39061 , \39062 , \39063 , \39064 ,
         \39065 , \39066 , \39067 , \39068 , \39069 , \39070 , \39071 , \39072 , \39073 , \39074 ,
         \39075 , \39076 , \39077 , \39078 , \39079 , \39080 , \39081 , \39082 , \39083 , \39084 ,
         \39085 , \39086 , \39087 , \39088 , \39089 , \39090 , \39091 , \39092 , \39093 , \39094 ,
         \39095 , \39096 , \39097 , \39098 , \39099 , \39100 , \39101 , \39102 , \39103 , \39104 ,
         \39105 , \39106 , \39107 , \39108 , \39109 , \39110 , \39111 , \39112 , \39113 , \39114 ,
         \39115 , \39116 , \39117 , \39118 , \39119 , \39120 , \39121 , \39122 , \39123 , \39124 ,
         \39125 , \39126 , \39127 , \39128 , \39129 , \39130 , \39131 , \39132 , \39133 , \39134 ,
         \39135 , \39136 , \39137 , \39138 , \39139 , \39140 , \39141 , \39142 , \39143 , \39144 ,
         \39145 , \39146 , \39147 , \39148 , \39149 , \39150 , \39151 , \39152 , \39153 , \39154 ,
         \39155 , \39156 , \39157 , \39158 , \39159 , \39160 , \39161 , \39162 , \39163 , \39164 ,
         \39165 , \39166 , \39167 , \39168 , \39169 , \39170 , \39171 , \39172 , \39173 , \39174 ,
         \39175 , \39176 , \39177 , \39178 , \39179 , \39180 , \39181 , \39182 , \39183 , \39184 ,
         \39185 , \39186 , \39187 , \39188 , \39189 , \39190 , \39191 , \39192 , \39193 , \39194 ,
         \39195 , \39196 , \39197 , \39198 , \39199 , \39200 , \39201 , \39202 , \39203 , \39204 ,
         \39205 , \39206 , \39207 , \39208 , \39209 , \39210 , \39211 , \39212 , \39213 , \39214 ,
         \39215 , \39216 , \39217 , \39218 , \39219 , \39220 , \39221 , \39222 , \39223 , \39224 ,
         \39225 , \39226 , \39227 , \39228 , \39229 , \39230 , \39231 , \39232 , \39233 , \39234 ,
         \39235 , \39236 , \39237 , \39238 , \39239 , \39240 , \39241 , \39242 , \39243 , \39244 ,
         \39245 , \39246 , \39247 , \39248 , \39249 , \39250 , \39251 , \39252 , \39253 , \39254 ,
         \39255 , \39256 , \39257 , \39258 , \39259 , \39260 , \39261 , \39262 , \39263 , \39264 ,
         \39265 , \39266 , \39267 , \39268 , \39269 , \39270 , \39271 , \39272 , \39273 , \39274 ,
         \39275 , \39276 , \39277 , \39278 , \39279 , \39280 , \39281 , \39282 , \39283 , \39284 ,
         \39285 , \39286 , \39287 , \39288 , \39289 , \39290 , \39291 , \39292 , \39293 , \39294 ,
         \39295 , \39296 , \39297 , \39298 , \39299 , \39300 , \39301 , \39302 , \39303 , \39304 ,
         \39305 , \39306 , \39307 , \39308 , \39309 , \39310 , \39311 , \39312 , \39313 , \39314 ,
         \39315 , \39316 , \39317 , \39318 , \39319 , \39320 , \39321 , \39322 , \39323 , \39324 ,
         \39325 , \39326 , \39327 , \39328 , \39329 , \39330 , \39331 , \39332 , \39333 , \39334 ,
         \39335 , \39336 , \39337 , \39338 , \39339 , \39340 , \39341 , \39342 , \39343 , \39344 ,
         \39345 , \39346 , \39347 , \39348 , \39349 , \39350 , \39351 , \39352 , \39353 , \39354 ,
         \39355 , \39356 , \39357 , \39358 , \39359 , \39360 , \39361 , \39362 , \39363 , \39364 ,
         \39365 , \39366 , \39367 , \39368 , \39369 , \39370 , \39371 , \39372 , \39373 , \39374 ,
         \39375 , \39376 , \39377 , \39378 , \39379 , \39380 , \39381 , \39382 , \39383 , \39384 ,
         \39385 , \39386 , \39387 , \39388 , \39389 , \39390 , \39391 , \39392 , \39393 , \39394 ,
         \39395 , \39396 , \39397 , \39398 , \39399 , \39400 , \39401 , \39402 , \39403 , \39404 ,
         \39405 , \39406 , \39407 , \39408 , \39409 , \39410 , \39411 , \39412 , \39413 , \39414 ,
         \39415 , \39416 , \39417 , \39418 , \39419 , \39420 , \39421 , \39422 , \39423 , \39424 ,
         \39425 , \39426 , \39427 , \39428 , \39429 , \39430 , \39431 , \39432 , \39433 , \39434 ,
         \39435 , \39436 , \39437 , \39438 , \39439 , \39440 , \39441 , \39442 , \39443 , \39444 ,
         \39445 , \39446 , \39447 , \39448 , \39449 , \39450 , \39451 , \39452 , \39453 , \39454 ,
         \39455 , \39456 , \39457 , \39458 , \39459 , \39460 , \39461 , \39462 , \39463 , \39464 ,
         \39465 , \39466 , \39467 , \39468 , \39469 , \39470 , \39471 , \39472 , \39473 , \39474 ,
         \39475 , \39476 , \39477 , \39478 , \39479 , \39480 , \39481 , \39482 , \39483 , \39484 ,
         \39485 , \39486 , \39487 , \39488 , \39489 , \39490 , \39491 , \39492 , \39493 , \39494 ,
         \39495 , \39496 , \39497 , \39498 , \39499 , \39500 , \39501 , \39502 , \39503 , \39504 ,
         \39505 , \39506 , \39507 , \39508 , \39509 , \39510 , \39511 , \39512 , \39513 , \39514 ,
         \39515 , \39516 , \39517 , \39518 , \39519 , \39520 , \39521 , \39522 , \39523 , \39524 ,
         \39525 , \39526 , \39527 , \39528 , \39529 , \39530 , \39531 , \39532 , \39533 , \39534 ,
         \39535 , \39536 , \39537 , \39538 , \39539 , \39540 , \39541 , \39542 , \39543 , \39544 ,
         \39545 , \39546 , \39547 , \39548 , \39549 , \39550 , \39551 , \39552 , \39553 , \39554 ,
         \39555 , \39556 , \39557 , \39558 , \39559 , \39560 , \39561 , \39562 , \39563 , \39564 ,
         \39565 , \39566 , \39567 , \39568 , \39569 , \39570 , \39571 , \39572 , \39573 , \39574 ,
         \39575 , \39576 , \39577 , \39578 , \39579 , \39580 , \39581 , \39582 , \39583 , \39584 ,
         \39585 , \39586 , \39587 , \39588 , \39589 , \39590 , \39591 , \39592 , \39593 , \39594 ,
         \39595 , \39596 , \39597 , \39598 , \39599 , \39600 , \39601 , \39602 , \39603 , \39604 ,
         \39605 , \39606 , \39607 , \39608 , \39609 , \39610 , \39611 , \39612 , \39613 , \39614 ,
         \39615 , \39616 , \39617 , \39618 , \39619 , \39620 , \39621 , \39622 , \39623 , \39624 ,
         \39625 , \39626 , \39627 , \39628 , \39629 , \39630 , \39631 , \39632 , \39633 , \39634 ,
         \39635 , \39636 , \39637 , \39638 , \39639 , \39640 , \39641 , \39642 , \39643 , \39644 ,
         \39645 , \39646 , \39647 , \39648 , \39649 , \39650 , \39651 , \39652 , \39653 , \39654 ,
         \39655 , \39656 , \39657 , \39658 , \39659 , \39660 , \39661 , \39662 , \39663 , \39664 ,
         \39665 , \39666 , \39667 , \39668 , \39669 , \39670 , \39671 , \39672 , \39673 , \39674 ,
         \39675 , \39676 , \39677 , \39678 , \39679 , \39680 , \39681 , \39682 , \39683 , \39684 ,
         \39685 , \39686 , \39687 , \39688 , \39689 , \39690 , \39691 , \39692 , \39693 , \39694 ,
         \39695 , \39696 , \39697 , \39698 , \39699 , \39700 , \39701 , \39702 , \39703 , \39704 ,
         \39705 , \39706 , \39707 , \39708 , \39709 , \39710 , \39711 , \39712 , \39713 , \39714 ,
         \39715 , \39716 , \39717 , \39718 , \39719 , \39720 , \39721 , \39722 , \39723 , \39724 ,
         \39725 , \39726 , \39727 , \39728 , \39729 , \39730 , \39731 , \39732 , \39733 , \39734 ,
         \39735 , \39736 , \39737 , \39738 , \39739 , \39740 , \39741 , \39742 , \39743 , \39744 ,
         \39745 , \39746 , \39747 , \39748 , \39749 , \39750 , \39751 , \39752 , \39753 , \39754 ,
         \39755 , \39756 , \39757 , \39758 , \39759 , \39760 , \39761 , \39762 , \39763 , \39764 ,
         \39765 , \39766 , \39767 , \39768 , \39769 , \39770 , \39771 , \39772 , \39773 , \39774 ,
         \39775 , \39776 , \39777 , \39778 , \39779 , \39780 , \39781 , \39782 , \39783 , \39784 ,
         \39785 , \39786 , \39787 , \39788 , \39789 , \39790 , \39791 , \39792 , \39793 , \39794 ,
         \39795 , \39796 , \39797 , \39798 , \39799 , \39800 , \39801 , \39802 , \39803 , \39804 ,
         \39805 , \39806 , \39807 , \39808 , \39809 , \39810 , \39811 , \39812 , \39813 , \39814 ,
         \39815 , \39816 , \39817 , \39818 , \39819 , \39820 , \39821 , \39822 , \39823 , \39824 ,
         \39825 , \39826 , \39827 , \39828 , \39829 , \39830 , \39831 , \39832 , \39833 , \39834 ,
         \39835 , \39836 , \39837 , \39838 , \39839 , \39840 , \39841 , \39842 , \39843 , \39844 ,
         \39845 , \39846 , \39847 , \39848 , \39849 , \39850 , \39851 , \39852 , \39853 , \39854 ,
         \39855 , \39856 , \39857 , \39858 , \39859 , \39860 , \39861 , \39862 , \39863 , \39864 ,
         \39865 , \39866 , \39867 , \39868 , \39869 , \39870 , \39871 , \39872 , \39873 , \39874 ,
         \39875 , \39876 , \39877 , \39878 , \39879 , \39880 , \39881 , \39882 , \39883 , \39884 ,
         \39885 , \39886 , \39887 , \39888 , \39889 , \39890 , \39891 , \39892 , \39893 , \39894 ,
         \39895 , \39896 , \39897 , \39898 , \39899 , \39900 , \39901 , \39902 , \39903 , \39904 ,
         \39905 , \39906 , \39907 , \39908 , \39909 , \39910 , \39911 , \39912 , \39913 , \39914 ,
         \39915 , \39916 , \39917 , \39918 , \39919 , \39920 , \39921 , \39922 , \39923 , \39924 ,
         \39925 , \39926 , \39927 , \39928 , \39929 , \39930 , \39931 , \39932 , \39933 , \39934 ,
         \39935 , \39936 , \39937 , \39938 , \39939 , \39940 , \39941 , \39942 , \39943 , \39944 ,
         \39945 , \39946 , \39947 , \39948 , \39949 , \39950 , \39951 , \39952 , \39953 , \39954 ,
         \39955 , \39956 , \39957 , \39958 , \39959 , \39960 , \39961 , \39962 , \39963 , \39964 ,
         \39965 , \39966 , \39967 , \39968 , \39969 , \39970 , \39971 , \39972 , \39973 , \39974 ,
         \39975 , \39976 , \39977 , \39978 , \39979 , \39980 , \39981 , \39982 , \39983 , \39984 ,
         \39985 , \39986 , \39987 , \39988 , \39989 , \39990 , \39991 , \39992 , \39993 , \39994 ,
         \39995 , \39996 , \39997 , \39998 , \39999 , \40000 , \40001 , \40002 , \40003 , \40004 ,
         \40005 , \40006 , \40007 , \40008 , \40009 , \40010 , \40011 , \40012 , \40013 , \40014 ,
         \40015 , \40016 , \40017 , \40018 , \40019 , \40020 , \40021 , \40022 , \40023 , \40024 ,
         \40025 , \40026 , \40027 , \40028 , \40029 , \40030 , \40031 , \40032 , \40033 , \40034 ,
         \40035 , \40036 , \40037 , \40038 , \40039 , \40040 , \40041 , \40042 , \40043 , \40044 ,
         \40045 , \40046 , \40047 , \40048 , \40049 , \40050 , \40051 , \40052 , \40053 , \40054 ,
         \40055 , \40056 , \40057 , \40058 , \40059 , \40060 , \40061 , \40062 , \40063 , \40064 ,
         \40065 , \40066 , \40067 , \40068 , \40069 , \40070 , \40071 , \40072 , \40073 , \40074 ,
         \40075 , \40076 , \40077 , \40078 , \40079 , \40080 , \40081 , \40082 , \40083 , \40084 ,
         \40085 , \40086 , \40087 , \40088 , \40089 , \40090 , \40091 , \40092 , \40093 , \40094 ,
         \40095 , \40096 , \40097 , \40098 , \40099 , \40100 , \40101 , \40102 , \40103 , \40104 ,
         \40105 , \40106 , \40107 , \40108 , \40109 , \40110 , \40111 , \40112 , \40113 , \40114 ,
         \40115 , \40116 , \40117 , \40118 , \40119 , \40120 , \40121 , \40122 , \40123 , \40124 ,
         \40125 , \40126 , \40127 , \40128 , \40129 , \40130 , \40131 , \40132 , \40133 , \40134 ,
         \40135 , \40136 , \40137 , \40138 , \40139 , \40140 , \40141 , \40142 , \40143 , \40144 ,
         \40145 , \40146 , \40147 , \40148 , \40149 , \40150 , \40151 , \40152 , \40153 , \40154 ,
         \40155 , \40156 , \40157 , \40158 , \40159 , \40160 , \40161 , \40162 , \40163 , \40164 ,
         \40165 , \40166 , \40167 , \40168 , \40169 , \40170 , \40171 , \40172 , \40173 , \40174 ,
         \40175 , \40176 , \40177 , \40178 , \40179 , \40180 , \40181 , \40182 , \40183 , \40184 ,
         \40185 , \40186 , \40187 , \40188 , \40189 , \40190 , \40191 , \40192 , \40193 , \40194 ,
         \40195 , \40196 , \40197 , \40198 , \40199 , \40200 , \40201 , \40202 , \40203 , \40204 ,
         \40205 , \40206 , \40207 , \40208 , \40209 , \40210 , \40211 , \40212 , \40213 , \40214 ,
         \40215 , \40216 , \40217 , \40218 , \40219 , \40220 , \40221 , \40222 , \40223 , \40224 ,
         \40225 , \40226 , \40227 , \40228 , \40229 , \40230 , \40231 , \40232 , \40233 , \40234 ,
         \40235 , \40236 , \40237 , \40238 , \40239 , \40240 , \40241 , \40242 , \40243 , \40244 ,
         \40245 , \40246 , \40247 , \40248 , \40249 , \40250 , \40251 , \40252 , \40253 , \40254 ,
         \40255 , \40256 , \40257 , \40258 , \40259 , \40260 , \40261 , \40262 , \40263 , \40264 ,
         \40265 , \40266 , \40267 , \40268 , \40269 , \40270 , \40271 , \40272 , \40273 , \40274 ,
         \40275 , \40276 , \40277 , \40278 , \40279 , \40280 , \40281 , \40282 , \40283 , \40284 ,
         \40285 , \40286 , \40287 , \40288 , \40289 , \40290 , \40291 , \40292 , \40293 , \40294 ,
         \40295 , \40296 , \40297 , \40298 , \40299 , \40300 , \40301 , \40302 , \40303 , \40304 ,
         \40305 , \40306 , \40307 , \40308 , \40309 , \40310 , \40311 , \40312 , \40313 , \40314 ,
         \40315 , \40316 , \40317 , \40318 , \40319 , \40320 , \40321 , \40322 , \40323 , \40324 ,
         \40325 , \40326 , \40327 , \40328 , \40329 , \40330 , \40331 , \40332 , \40333 , \40334 ,
         \40335 , \40336 , \40337 , \40338 , \40339 , \40340 , \40341 , \40342 , \40343 , \40344 ,
         \40345 , \40346 , \40347 , \40348 , \40349 , \40350 , \40351 , \40352 , \40353 , \40354 ,
         \40355 , \40356 , \40357 , \40358 , \40359 , \40360 , \40361 , \40362 , \40363 , \40364 ,
         \40365 , \40366 , \40367 , \40368 , \40369 , \40370 , \40371 , \40372 , \40373 , \40374 ,
         \40375 , \40376 , \40377 , \40378 , \40379 , \40380 , \40381 , \40382 , \40383 , \40384 ,
         \40385 , \40386 , \40387 , \40388 , \40389 , \40390 , \40391 , \40392 , \40393 , \40394 ,
         \40395 , \40396 , \40397 , \40398 , \40399 , \40400 , \40401 , \40402 , \40403 , \40404 ,
         \40405 , \40406 , \40407 , \40408 , \40409 , \40410 , \40411 , \40412 , \40413 , \40414 ,
         \40415 , \40416 , \40417 , \40418 , \40419 , \40420 , \40421 , \40422 , \40423 , \40424 ,
         \40425 , \40426 , \40427 , \40428 , \40429 , \40430 , \40431 , \40432 , \40433 , \40434 ,
         \40435 , \40436 , \40437 , \40438 , \40439 , \40440 , \40441 , \40442 , \40443 , \40444 ,
         \40445 , \40446 , \40447 , \40448 , \40449 , \40450 , \40451 , \40452 , \40453 , \40454 ,
         \40455 , \40456 , \40457 , \40458 , \40459 , \40460 , \40461 , \40462 , \40463 , \40464 ,
         \40465 , \40466 , \40467 , \40468 , \40469 , \40470 , \40471 , \40472 , \40473 , \40474 ,
         \40475 , \40476 , \40477 , \40478 , \40479 , \40480 , \40481 , \40482 , \40483 , \40484 ,
         \40485 , \40486 , \40487 , \40488 , \40489 , \40490 , \40491 , \40492 , \40493 , \40494 ,
         \40495 , \40496 , \40497 , \40498 , \40499 , \40500 , \40501 , \40502 , \40503 , \40504 ,
         \40505 , \40506 , \40507 , \40508 , \40509 , \40510 , \40511 , \40512 , \40513 , \40514 ,
         \40515 , \40516 , \40517 , \40518 , \40519 , \40520 , \40521 , \40522 , \40523 , \40524 ,
         \40525 , \40526 , \40527 , \40528 , \40529 , \40530 , \40531 , \40532 , \40533 , \40534 ,
         \40535 , \40536 , \40537 , \40538 , \40539 , \40540 , \40541 , \40542 , \40543 , \40544 ,
         \40545 , \40546 , \40547 , \40548 , \40549 , \40550 , \40551 , \40552 , \40553 , \40554 ,
         \40555 , \40556 , \40557 , \40558 , \40559 , \40560 , \40561 , \40562 , \40563 , \40564 ,
         \40565 , \40566 , \40567 , \40568 , \40569 , \40570 , \40571 , \40572 , \40573 , \40574 ,
         \40575 , \40576 , \40577 , \40578 , \40579 , \40580 , \40581 , \40582 , \40583 , \40584 ,
         \40585 , \40586 , \40587 , \40588 , \40589 , \40590 , \40591 , \40592 , \40593 , \40594 ,
         \40595 , \40596 , \40597 , \40598 , \40599 , \40600 , \40601 , \40602 , \40603 , \40604 ,
         \40605 , \40606 , \40607 , \40608 , \40609 , \40610 , \40611 , \40612 , \40613 , \40614 ,
         \40615 , \40616 , \40617 , \40618 , \40619 , \40620 , \40621 , \40622 , \40623 , \40624 ,
         \40625 , \40626 , \40627 , \40628 , \40629 , \40630 , \40631 , \40632 , \40633 , \40634 ,
         \40635 , \40636 , \40637 , \40638 , \40639 , \40640 , \40641 , \40642 , \40643 , \40644 ,
         \40645 , \40646 , \40647 , \40648 , \40649 , \40650 , \40651 , \40652 , \40653 , \40654 ,
         \40655 , \40656 , \40657 , \40658 , \40659 , \40660 , \40661 , \40662 , \40663 , \40664 ,
         \40665 , \40666 , \40667 , \40668 , \40669 , \40670 , \40671 , \40672 , \40673 , \40674 ,
         \40675 , \40676 , \40677 , \40678 , \40679 , \40680 , \40681 , \40682 , \40683 , \40684 ,
         \40685 , \40686 , \40687 , \40688 , \40689 , \40690 , \40691 , \40692 , \40693 , \40694 ,
         \40695 , \40696 , \40697 , \40698 , \40699 , \40700 , \40701 , \40702 , \40703 , \40704 ,
         \40705 , \40706 , \40707 , \40708 , \40709 , \40710 , \40711 , \40712 , \40713 , \40714 ,
         \40715 , \40716 , \40717 , \40718 , \40719 , \40720 , \40721 , \40722 , \40723 , \40724 ,
         \40725 , \40726 , \40727 , \40728 , \40729 , \40730 , \40731 , \40732 , \40733 , \40734 ,
         \40735 , \40736 , \40737 , \40738 , \40739 , \40740 , \40741 , \40742 , \40743 , \40744 ,
         \40745 , \40746 , \40747 , \40748 , \40749 , \40750 , \40751 , \40752 , \40753 , \40754 ,
         \40755 , \40756 , \40757 , \40758 , \40759 , \40760 , \40761 , \40762 , \40763 , \40764 ,
         \40765 , \40766 , \40767 , \40768 , \40769 , \40770 , \40771 , \40772 , \40773 , \40774 ,
         \40775 , \40776 , \40777 , \40778 , \40779 , \40780 , \40781 , \40782 , \40783 , \40784 ,
         \40785 , \40786 , \40787 , \40788 , \40789 , \40790 , \40791 , \40792 , \40793 , \40794 ,
         \40795 , \40796 , \40797 , \40798 , \40799 , \40800 , \40801 , \40802 , \40803 , \40804 ,
         \40805 , \40806 , \40807 , \40808 , \40809 , \40810 , \40811 , \40812 , \40813 , \40814 ,
         \40815 , \40816 , \40817 , \40818 , \40819 , \40820 , \40821 , \40822 , \40823 , \40824 ,
         \40825 , \40826 , \40827 , \40828 , \40829 , \40830 , \40831 , \40832 , \40833 , \40834 ,
         \40835 , \40836 , \40837 , \40838 , \40839 , \40840 , \40841 , \40842 , \40843 , \40844 ,
         \40845 , \40846 , \40847 , \40848 , \40849 , \40850 , \40851 , \40852 , \40853 , \40854 ,
         \40855 , \40856 , \40857 , \40858 , \40859 , \40860 , \40861 , \40862 , \40863 , \40864 ,
         \40865 , \40866 , \40867 , \40868 , \40869 , \40870 , \40871 , \40872 , \40873 , \40874 ,
         \40875 , \40876 , \40877 , \40878 , \40879 , \40880 , \40881 , \40882 , \40883 , \40884 ,
         \40885 , \40886 , \40887 , \40888 , \40889 , \40890 , \40891 , \40892 , \40893 , \40894 ,
         \40895 , \40896 , \40897 , \40898 , \40899 , \40900 , \40901 , \40902 , \40903 , \40904 ,
         \40905 , \40906 , \40907 , \40908 , \40909 , \40910 , \40911 , \40912 , \40913 , \40914 ,
         \40915 , \40916 , \40917 , \40918 , \40919 , \40920 , \40921 , \40922 , \40923 , \40924 ,
         \40925 , \40926 , \40927 , \40928 , \40929 , \40930 , \40931 , \40932 , \40933 , \40934 ,
         \40935 , \40936 , \40937 , \40938 , \40939 , \40940 , \40941 , \40942 , \40943 , \40944 ,
         \40945 , \40946 , \40947 , \40948 , \40949 , \40950 , \40951 , \40952 , \40953 , \40954 ,
         \40955 , \40956 , \40957 , \40958 , \40959 , \40960 , \40961 , \40962 , \40963 , \40964 ,
         \40965 , \40966 , \40967 , \40968 , \40969 , \40970 , \40971 , \40972 , \40973 , \40974 ,
         \40975 , \40976 , \40977 , \40978 , \40979 , \40980 , \40981 , \40982 , \40983 , \40984 ,
         \40985 , \40986 , \40987 , \40988 , \40989 , \40990 , \40991 , \40992 , \40993 , \40994 ,
         \40995 , \40996 , \40997 , \40998 , \40999 , \41000 , \41001 , \41002 , \41003 , \41004 ,
         \41005 , \41006 , \41007 , \41008 , \41009 , \41010 , \41011 , \41012 , \41013 , \41014 ,
         \41015 , \41016 , \41017 , \41018 , \41019 , \41020 , \41021 , \41022 , \41023 , \41024 ,
         \41025 , \41026 , \41027 , \41028 , \41029 , \41030 , \41031 , \41032 , \41033 , \41034 ,
         \41035 , \41036 , \41037 , \41038 , \41039 , \41040 , \41041 , \41042 , \41043 , \41044 ,
         \41045 , \41046 , \41047 , \41048 , \41049 , \41050 , \41051 , \41052 , \41053 , \41054 ,
         \41055 , \41056 , \41057 , \41058 , \41059 , \41060 , \41061 , \41062 , \41063 , \41064 ,
         \41065 , \41066 , \41067 , \41068 , \41069 , \41070 , \41071 , \41072 , \41073 , \41074 ,
         \41075 , \41076 , \41077 , \41078 , \41079 , \41080 , \41081 , \41082 , \41083 , \41084 ,
         \41085 , \41086 , \41087 , \41088 , \41089 , \41090 , \41091 , \41092 , \41093 , \41094 ,
         \41095 , \41096 , \41097 , \41098 , \41099 , \41100 , \41101 , \41102 , \41103 , \41104 ,
         \41105 , \41106 , \41107 , \41108 , \41109 , \41110 , \41111 , \41112 , \41113 , \41114 ,
         \41115 , \41116 , \41117 , \41118 , \41119 , \41120 , \41121 , \41122 , \41123 , \41124 ,
         \41125 , \41126 , \41127 , \41128 , \41129 , \41130 , \41131 , \41132 , \41133 , \41134 ,
         \41135 , \41136 , \41137 , \41138 , \41139 , \41140 , \41141 , \41142 , \41143 , \41144 ,
         \41145 , \41146 , \41147 , \41148 , \41149 , \41150 , \41151 , \41152 , \41153 , \41154 ,
         \41155 , \41156 , \41157 , \41158 , \41159 , \41160 , \41161 , \41162 , \41163 , \41164 ,
         \41165 , \41166 , \41167 , \41168 , \41169 , \41170 , \41171 , \41172 , \41173 , \41174 ,
         \41175 , \41176 , \41177 , \41178 , \41179 , \41180 , \41181 , \41182 , \41183 , \41184 ,
         \41185 , \41186 , \41187 , \41188 , \41189 , \41190 , \41191 , \41192 , \41193 , \41194 ,
         \41195 , \41196 , \41197 , \41198 , \41199 , \41200 , \41201 , \41202 , \41203 , \41204 ,
         \41205 , \41206 , \41207 , \41208 , \41209 , \41210 , \41211 , \41212 , \41213 , \41214 ,
         \41215 , \41216 , \41217 , \41218 , \41219 , \41220 , \41221 , \41222 , \41223 , \41224 ,
         \41225 , \41226 , \41227 , \41228 , \41229 , \41230 , \41231 , \41232 , \41233 , \41234 ,
         \41235 , \41236 , \41237 , \41238 , \41239 , \41240 , \41241 , \41242 , \41243 , \41244 ,
         \41245 , \41246 , \41247 , \41248 , \41249 , \41250 , \41251 , \41252 , \41253 , \41254 ,
         \41255 , \41256 , \41257 , \41258 , \41259 , \41260 , \41261 , \41262 , \41263 , \41264 ,
         \41265 , \41266 , \41267 , \41268 , \41269 , \41270 , \41271 , \41272 , \41273 , \41274 ,
         \41275 , \41276 , \41277 , \41278 , \41279 , \41280 , \41281 , \41282 , \41283 , \41284 ,
         \41285 , \41286 , \41287 , \41288 , \41289 , \41290 , \41291 , \41292 , \41293 , \41294 ,
         \41295 , \41296 , \41297 , \41298 , \41299 , \41300 , \41301 , \41302 , \41303 , \41304 ,
         \41305 , \41306 , \41307 , \41308 , \41309 , \41310 , \41311 , \41312 , \41313 , \41314 ,
         \41315 , \41316 , \41317 , \41318 , \41319 , \41320 , \41321 , \41322 , \41323 , \41324 ,
         \41325 , \41326 , \41327 , \41328 , \41329 , \41330 , \41331 , \41332 , \41333 , \41334 ,
         \41335 , \41336 , \41337 , \41338 , \41339 , \41340 , \41341 , \41342 , \41343 , \41344 ,
         \41345 , \41346 , \41347 , \41348 , \41349 , \41350 , \41351 , \41352 , \41353 , \41354 ,
         \41355 , \41356 , \41357 , \41358 , \41359 , \41360 , \41361 , \41362 , \41363 , \41364 ,
         \41365 , \41366 , \41367 , \41368 , \41369 , \41370 , \41371 , \41372 , \41373 , \41374 ,
         \41375 , \41376 , \41377 , \41378 , \41379 , \41380 , \41381 , \41382 , \41383 , \41384 ,
         \41385 , \41386 , \41387 , \41388 , \41389 , \41390 , \41391 , \41392 , \41393 , \41394 ,
         \41395 , \41396 , \41397 , \41398 , \41399 , \41400 , \41401 , \41402 , \41403 , \41404 ,
         \41405 , \41406 , \41407 , \41408 , \41409 , \41410 , \41411 , \41412 , \41413 , \41414 ,
         \41415 , \41416 , \41417 , \41418 , \41419 , \41420 , \41421 , \41422 , \41423 , \41424 ,
         \41425 , \41426 , \41427 , \41428 , \41429 , \41430 , \41431 , \41432 , \41433 , \41434 ,
         \41435 , \41436 , \41437 , \41438 , \41439 , \41440 , \41441 , \41442 , \41443 , \41444 ,
         \41445 , \41446 , \41447 , \41448 , \41449 , \41450 , \41451 , \41452 , \41453 , \41454 ,
         \41455 , \41456 , \41457 , \41458 , \41459 , \41460 , \41461 , \41462 , \41463 , \41464 ,
         \41465 , \41466 , \41467 , \41468 , \41469 , \41470 , \41471 , \41472 , \41473 , \41474 ,
         \41475 , \41476 , \41477 , \41478 , \41479 , \41480 , \41481 , \41482 , \41483 , \41484 ,
         \41485 , \41486 , \41487 , \41488 , \41489 , \41490 , \41491 , \41492 , \41493 , \41494 ,
         \41495 , \41496 , \41497 , \41498 , \41499 , \41500 , \41501 , \41502 , \41503 , \41504 ,
         \41505 , \41506 , \41507 , \41508 , \41509 , \41510 , \41511 , \41512 , \41513 , \41514 ,
         \41515 , \41516 , \41517 , \41518 , \41519 , \41520 , \41521 , \41522 , \41523 , \41524 ,
         \41525 , \41526 , \41527 , \41528 , \41529 , \41530 , \41531 , \41532 , \41533 , \41534 ,
         \41535 , \41536 , \41537 , \41538 , \41539 , \41540 , \41541 , \41542 , \41543 , \41544 ,
         \41545 , \41546 , \41547 , \41548 , \41549 , \41550 , \41551 , \41552 , \41553 , \41554 ,
         \41555 , \41556 , \41557 , \41558 , \41559 , \41560 , \41561 , \41562 , \41563 , \41564 ,
         \41565 , \41566 , \41567 , \41568 , \41569 , \41570 , \41571 , \41572 , \41573 , \41574 ,
         \41575 , \41576 , \41577 , \41578 , \41579 , \41580 , \41581 , \41582 , \41583 , \41584 ,
         \41585 , \41586 , \41587 , \41588 , \41589 , \41590 , \41591 , \41592 , \41593 , \41594 ,
         \41595 , \41596 , \41597 , \41598 , \41599 , \41600 , \41601 , \41602 , \41603 , \41604 ,
         \41605 , \41606 , \41607 , \41608 , \41609 , \41610 , \41611 , \41612 , \41613 , \41614 ,
         \41615 , \41616 , \41617 , \41618 , \41619 , \41620 , \41621 , \41622 , \41623 , \41624 ,
         \41625 , \41626 , \41627 , \41628 , \41629 , \41630 , \41631 , \41632 , \41633 , \41634 ,
         \41635 , \41636 , \41637 , \41638 , \41639 , \41640 , \41641 , \41642 , \41643 , \41644 ,
         \41645 , \41646 , \41647 , \41648 , \41649 , \41650 , \41651 , \41652 , \41653 , \41654 ,
         \41655 , \41656 , \41657 , \41658 , \41659 , \41660 , \41661 , \41662 , \41663 , \41664 ,
         \41665 , \41666 , \41667 , \41668 , \41669 , \41670 , \41671 , \41672 , \41673 , \41674 ,
         \41675 , \41676 , \41677 , \41678 , \41679 , \41680 , \41681 , \41682 , \41683 , \41684 ,
         \41685 , \41686 , \41687 , \41688 , \41689 , \41690 , \41691 , \41692 , \41693 , \41694 ,
         \41695 , \41696 , \41697 , \41698 , \41699 , \41700 , \41701 , \41702 , \41703 , \41704 ,
         \41705 , \41706 , \41707 , \41708 , \41709 , \41710 , \41711 , \41712 , \41713 , \41714 ,
         \41715 , \41716 , \41717 , \41718 , \41719 , \41720 , \41721 , \41722 , \41723 , \41724 ,
         \41725 , \41726 , \41727 , \41728 , \41729 , \41730 , \41731 , \41732 , \41733 , \41734 ,
         \41735 , \41736 , \41737 , \41738 , \41739 , \41740 , \41741 , \41742 , \41743 , \41744 ,
         \41745 , \41746 , \41747 , \41748 , \41749 , \41750 , \41751 , \41752 , \41753 , \41754 ,
         \41755 , \41756 , \41757 , \41758 , \41759 , \41760 , \41761 , \41762 , \41763 , \41764 ,
         \41765 , \41766 , \41767 , \41768 , \41769 , \41770 , \41771 , \41772 , \41773 , \41774 ,
         \41775 , \41776 , \41777 , \41778 , \41779 , \41780 , \41781 , \41782 , \41783 , \41784 ,
         \41785 , \41786 , \41787 , \41788 , \41789 , \41790 , \41791 , \41792 , \41793 , \41794 ,
         \41795 , \41796 , \41797 , \41798 , \41799 , \41800 , \41801 , \41802 , \41803 , \41804 ,
         \41805 , \41806 , \41807 , \41808 , \41809 , \41810 , \41811 , \41812 , \41813 , \41814 ,
         \41815 , \41816 , \41817 , \41818 , \41819 , \41820 , \41821 , \41822 , \41823 , \41824 ,
         \41825 , \41826 , \41827 , \41828 , \41829 , \41830 , \41831 , \41832 , \41833 , \41834 ,
         \41835 , \41836 , \41837 , \41838 , \41839 , \41840 , \41841 , \41842 , \41843 , \41844 ,
         \41845 , \41846 , \41847 , \41848 , \41849 , \41850 , \41851 , \41852 , \41853 , \41854 ,
         \41855 , \41856 , \41857 , \41858 , \41859 , \41860 , \41861 , \41862 , \41863 , \41864 ,
         \41865 , \41866 , \41867 , \41868 , \41869 , \41870 , \41871 , \41872 , \41873 , \41874 ,
         \41875 , \41876 , \41877 , \41878 , \41879 , \41880 , \41881 , \41882 , \41883 , \41884 ,
         \41885 , \41886 , \41887 , \41888 , \41889 , \41890 , \41891 , \41892 , \41893 , \41894 ,
         \41895 , \41896 , \41897 , \41898 , \41899 , \41900 , \41901 , \41902 , \41903 , \41904 ,
         \41905 , \41906 , \41907 , \41908 , \41909 , \41910 , \41911 , \41912 , \41913 , \41914 ,
         \41915 , \41916 , \41917 , \41918 , \41919 , \41920 , \41921 , \41922 , \41923 , \41924 ,
         \41925 , \41926 , \41927 , \41928 , \41929 , \41930 , \41931 , \41932 , \41933 , \41934 ,
         \41935 , \41936 , \41937 , \41938 , \41939 , \41940 , \41941 , \41942 , \41943 , \41944 ,
         \41945 , \41946 , \41947 , \41948 , \41949 , \41950 , \41951 , \41952 , \41953 , \41954 ,
         \41955 , \41956 , \41957 , \41958 , \41959 , \41960 , \41961 , \41962 , \41963 , \41964 ,
         \41965 , \41966 , \41967 , \41968 , \41969 , \41970 , \41971 , \41972 , \41973 , \41974 ,
         \41975 , \41976 , \41977 , \41978 , \41979 , \41980 , \41981 , \41982 , \41983 , \41984 ,
         \41985 , \41986 , \41987 , \41988 , \41989 , \41990 , \41991 , \41992 , \41993 , \41994 ,
         \41995 , \41996 , \41997 , \41998 , \41999 , \42000 , \42001 , \42002 , \42003 , \42004 ,
         \42005 , \42006 , \42007 , \42008 , \42009 , \42010 , \42011 , \42012 , \42013 , \42014 ,
         \42015 , \42016 , \42017 , \42018 , \42019 , \42020 , \42021 , \42022 , \42023 , \42024 ,
         \42025 , \42026 , \42027 , \42028 , \42029 , \42030 , \42031 , \42032 , \42033 , \42034 ,
         \42035 , \42036 , \42037 , \42038 , \42039 , \42040 , \42041 , \42042 , \42043 , \42044 ,
         \42045 , \42046 , \42047 , \42048 , \42049 , \42050 , \42051 , \42052 , \42053 , \42054 ,
         \42055 , \42056 , \42057 , \42058 , \42059 , \42060 , \42061 , \42062 , \42063 , \42064 ,
         \42065 , \42066 , \42067 , \42068 , \42069 , \42070 , \42071 , \42072 , \42073 , \42074 ,
         \42075 , \42076 , \42077 , \42078 , \42079 , \42080 , \42081 , \42082 , \42083 , \42084 ,
         \42085 , \42086 , \42087 , \42088 , \42089 , \42090 , \42091 , \42092 , \42093 , \42094 ,
         \42095 , \42096 , \42097 , \42098 , \42099 , \42100 , \42101 , \42102 , \42103 , \42104 ,
         \42105 , \42106 , \42107 , \42108 , \42109 , \42110 , \42111 , \42112 , \42113 , \42114 ,
         \42115 , \42116 , \42117 , \42118 , \42119 , \42120 , \42121 , \42122 , \42123 , \42124 ,
         \42125 , \42126 , \42127 , \42128 , \42129 , \42130 , \42131 , \42132 , \42133 , \42134 ,
         \42135 , \42136 , \42137 , \42138 , \42139 , \42140 , \42141 , \42142 , \42143 , \42144 ,
         \42145 , \42146 , \42147 , \42148 , \42149 , \42150 , \42151 , \42152 , \42153 , \42154 ,
         \42155 , \42156 , \42157 , \42158 , \42159 , \42160 , \42161 , \42162 , \42163 , \42164 ,
         \42165 , \42166 , \42167 , \42168 , \42169 , \42170 , \42171 , \42172 , \42173 , \42174 ,
         \42175 , \42176 , \42177 , \42178 , \42179 , \42180 , \42181 , \42182 , \42183 , \42184 ,
         \42185 , \42186 , \42187 , \42188 , \42189 , \42190 , \42191 , \42192 , \42193 , \42194 ,
         \42195 , \42196 , \42197 , \42198 , \42199 , \42200 , \42201 , \42202 , \42203 , \42204 ,
         \42205 , \42206 , \42207 , \42208 , \42209 , \42210 , \42211 , \42212 , \42213 , \42214 ,
         \42215 , \42216 , \42217 , \42218 , \42219 , \42220 , \42221 , \42222 , \42223 , \42224 ,
         \42225 , \42226 , \42227 , \42228 , \42229 , \42230 , \42231 , \42232 , \42233 , \42234 ,
         \42235 , \42236 , \42237 , \42238 , \42239 , \42240 , \42241 , \42242 , \42243 , \42244 ,
         \42245 , \42246 , \42247 , \42248 , \42249 , \42250 , \42251 , \42252 , \42253 , \42254 ,
         \42255 , \42256 , \42257 , \42258 , \42259 , \42260 , \42261 , \42262 , \42263 , \42264 ,
         \42265 , \42266 , \42267 , \42268 , \42269 , \42270 , \42271 , \42272 , \42273 , \42274 ,
         \42275 , \42276 , \42277 , \42278 , \42279 , \42280 , \42281 , \42282 , \42283 , \42284 ,
         \42285 , \42286 , \42287 , \42288 , \42289 , \42290 , \42291 , \42292 , \42293 , \42294 ,
         \42295 , \42296 , \42297 , \42298 , \42299 , \42300 , \42301 , \42302 , \42303 , \42304 ,
         \42305 , \42306 , \42307 , \42308 , \42309 , \42310 , \42311 , \42312 , \42313 , \42314 ,
         \42315 , \42316 , \42317 , \42318 , \42319 , \42320 , \42321 , \42322 , \42323 , \42324 ,
         \42325 , \42326 , \42327 , \42328 , \42329 , \42330 , \42331 , \42332 , \42333 , \42334 ,
         \42335 , \42336 , \42337 , \42338 , \42339 , \42340 , \42341 , \42342 , \42343 , \42344 ,
         \42345 , \42346 , \42347 , \42348 , \42349 , \42350 , \42351 , \42352 , \42353 , \42354 ,
         \42355 , \42356 , \42357 , \42358 , \42359 , \42360 , \42361 , \42362 , \42363 , \42364 ,
         \42365 , \42366 , \42367 , \42368 , \42369 , \42370 , \42371 , \42372 , \42373 , \42374 ,
         \42375 , \42376 , \42377 , \42378 , \42379 , \42380 , \42381 , \42382 , \42383 , \42384 ,
         \42385 , \42386 , \42387 , \42388 , \42389 , \42390 , \42391 , \42392 , \42393 , \42394 ,
         \42395 , \42396 , \42397 , \42398 , \42399 , \42400 , \42401 , \42402 , \42403 , \42404 ,
         \42405 , \42406 , \42407 , \42408 , \42409 , \42410 , \42411 , \42412 , \42413 , \42414 ,
         \42415 , \42416 , \42417 , \42418 , \42419 , \42420 , \42421 , \42422 , \42423 , \42424 ,
         \42425 , \42426 , \42427 , \42428 , \42429 , \42430 , \42431 , \42432 , \42433 , \42434 ,
         \42435 , \42436 , \42437 , \42438 , \42439 , \42440 , \42441 , \42442 , \42443 , \42444 ,
         \42445 , \42446 , \42447 , \42448 , \42449 , \42450 , \42451 , \42452 , \42453 , \42454 ,
         \42455 , \42456 , \42457 , \42458 , \42459 , \42460 , \42461 , \42462 , \42463 , \42464 ,
         \42465 , \42466 , \42467 , \42468 , \42469 , \42470 , \42471 , \42472 , \42473 , \42474 ,
         \42475 , \42476 , \42477 , \42478 , \42479 , \42480 , \42481 , \42482 , \42483 , \42484 ,
         \42485 , \42486 , \42487 , \42488 , \42489 , \42490 , \42491 , \42492 , \42493 , \42494 ,
         \42495 , \42496 , \42497 , \42498 , \42499 , \42500 , \42501 , \42502 , \42503 , \42504 ,
         \42505 , \42506 , \42507 , \42508 , \42509 , \42510 , \42511 , \42512 , \42513 , \42514 ,
         \42515 , \42516 , \42517 , \42518 , \42519 , \42520 , \42521 , \42522 , \42523 , \42524 ,
         \42525 , \42526 , \42527 , \42528 , \42529 , \42530 , \42531 , \42532 , \42533 , \42534 ,
         \42535 , \42536 , \42537 , \42538 , \42539 , \42540 , \42541 , \42542 , \42543 , \42544 ,
         \42545 , \42546 , \42547 , \42548 , \42549 , \42550 , \42551 , \42552 , \42553 , \42554 ,
         \42555 , \42556 , \42557 , \42558 , \42559 , \42560 , \42561 , \42562 , \42563 , \42564 ,
         \42565 , \42566 , \42567 , \42568 , \42569 , \42570 , \42571 , \42572 , \42573 , \42574 ,
         \42575 , \42576 , \42577 , \42578 , \42579 , \42580 , \42581 , \42582 , \42583 , \42584 ,
         \42585 , \42586 , \42587 , \42588 , \42589 , \42590 , \42591 , \42592 , \42593 , \42594 ,
         \42595 , \42596 , \42597 , \42598 , \42599 , \42600 , \42601 , \42602 , \42603 , \42604 ,
         \42605 , \42606 , \42607 , \42608 , \42609 , \42610 , \42611 , \42612 , \42613 , \42614 ,
         \42615 , \42616 , \42617 , \42618 , \42619 , \42620 , \42621 , \42622 , \42623 , \42624 ,
         \42625 , \42626 , \42627 , \42628 , \42629 , \42630 , \42631 , \42632 , \42633 , \42634 ,
         \42635 , \42636 , \42637 , \42638 , \42639 , \42640 , \42641 , \42642 , \42643 , \42644 ,
         \42645 , \42646 , \42647 , \42648 , \42649 , \42650 , \42651 , \42652 , \42653 , \42654 ,
         \42655 , \42656 , \42657 , \42658 , \42659 , \42660 , \42661 , \42662 , \42663 , \42664 ,
         \42665 , \42666 , \42667 , \42668 , \42669 , \42670 , \42671 , \42672 , \42673 , \42674 ,
         \42675 , \42676 , \42677 , \42678 , \42679 , \42680 , \42681 , \42682 , \42683 , \42684 ,
         \42685 , \42686 , \42687 , \42688 , \42689 , \42690 , \42691 , \42692 , \42693 , \42694 ,
         \42695 , \42696 , \42697 , \42698 , \42699 , \42700 , \42701 , \42702 , \42703 , \42704 ,
         \42705 , \42706 , \42707 , \42708 , \42709 , \42710 , \42711 , \42712 , \42713 , \42714 ,
         \42715 , \42716 , \42717 , \42718 , \42719 , \42720 , \42721 , \42722 , \42723 , \42724 ,
         \42725 , \42726 , \42727 , \42728 , \42729 , \42730 , \42731 , \42732 , \42733 , \42734 ,
         \42735 , \42736 , \42737 , \42738 , \42739 , \42740 , \42741 , \42742 , \42743 , \42744 ,
         \42745 , \42746 , \42747 , \42748 , \42749 , \42750 , \42751 , \42752 , \42753 , \42754 ,
         \42755 , \42756 , \42757 , \42758 , \42759 , \42760 , \42761 , \42762 , \42763 , \42764 ,
         \42765 , \42766 , \42767 , \42768 , \42769 , \42770 , \42771 , \42772 , \42773 , \42774 ,
         \42775 , \42776 , \42777 , \42778 , \42779 , \42780 , \42781 , \42782 , \42783 , \42784 ,
         \42785 , \42786 , \42787 , \42788 , \42789 , \42790 , \42791 , \42792 , \42793 , \42794 ,
         \42795 , \42796 , \42797 , \42798 , \42799 , \42800 , \42801 , \42802 , \42803 , \42804 ,
         \42805 , \42806 , \42807 , \42808 , \42809 , \42810 , \42811 , \42812 , \42813 , \42814 ,
         \42815 , \42816 , \42817 , \42818 , \42819 , \42820 , \42821 , \42822 , \42823 , \42824 ,
         \42825 , \42826 , \42827 , \42828 , \42829 , \42830 , \42831 , \42832 , \42833 , \42834 ,
         \42835 , \42836 , \42837 , \42838 , \42839 , \42840 , \42841 , \42842 , \42843 , \42844 ,
         \42845 , \42846 , \42847 , \42848 , \42849 , \42850 , \42851 , \42852 , \42853 , \42854 ,
         \42855 , \42856 , \42857 , \42858 , \42859 , \42860 , \42861 , \42862 , \42863 , \42864 ,
         \42865 , \42866 , \42867 , \42868 , \42869 , \42870 , \42871 , \42872 , \42873 , \42874 ,
         \42875 , \42876 , \42877 , \42878 , \42879 , \42880 , \42881 , \42882 , \42883 , \42884 ,
         \42885 , \42886 , \42887 , \42888 , \42889 , \42890 , \42891 , \42892 , \42893 , \42894 ,
         \42895 , \42896 , \42897 , \42898 , \42899 , \42900 , \42901 , \42902 , \42903 , \42904 ,
         \42905 , \42906 , \42907 , \42908 , \42909 , \42910 , \42911 , \42912 , \42913 , \42914 ,
         \42915 , \42916 , \42917 , \42918 , \42919 , \42920 , \42921 , \42922 , \42923 , \42924 ,
         \42925 , \42926 , \42927 , \42928 , \42929 , \42930 , \42931 , \42932 , \42933 , \42934 ,
         \42935 , \42936 , \42937 , \42938 , \42939 , \42940 , \42941 , \42942 , \42943 , \42944 ,
         \42945 , \42946 , \42947 , \42948 , \42949 , \42950 , \42951 , \42952 , \42953 , \42954 ,
         \42955 , \42956 , \42957 , \42958 , \42959 , \42960 , \42961 , \42962 , \42963 , \42964 ,
         \42965 , \42966 , \42967 , \42968 , \42969 , \42970 , \42971 , \42972 , \42973 , \42974 ,
         \42975 , \42976 , \42977 , \42978 , \42979 , \42980 , \42981 , \42982 , \42983 , \42984 ,
         \42985 , \42986 , \42987 , \42988 , \42989 , \42990 , \42991 , \42992 , \42993 , \42994 ,
         \42995 , \42996 , \42997 , \42998 , \42999 , \43000 , \43001 , \43002 , \43003 , \43004 ,
         \43005 , \43006 , \43007 , \43008 , \43009 , \43010 , \43011 , \43012 , \43013 , \43014 ,
         \43015 , \43016 , \43017 , \43018 , \43019 , \43020 , \43021 , \43022 , \43023 , \43024 ,
         \43025 , \43026 , \43027 , \43028 , \43029 , \43030 , \43031 , \43032 , \43033 , \43034 ,
         \43035 , \43036 , \43037 , \43038 , \43039 , \43040 , \43041 , \43042 , \43043 , \43044 ,
         \43045 , \43046 , \43047 , \43048 , \43049 , \43050 , \43051 , \43052 , \43053 , \43054 ,
         \43055 , \43056 , \43057 , \43058 , \43059 , \43060 , \43061 , \43062 , \43063 , \43064 ,
         \43065 , \43066 , \43067 , \43068 , \43069 , \43070 , \43071 , \43072 , \43073 , \43074 ,
         \43075 , \43076 , \43077 , \43078 , \43079 , \43080 , \43081 , \43082 , \43083 , \43084 ,
         \43085 , \43086 , \43087 , \43088 , \43089 , \43090 , \43091 , \43092 , \43093 , \43094 ,
         \43095 , \43096 , \43097 , \43098 , \43099 , \43100 , \43101 , \43102 , \43103 , \43104 ,
         \43105 , \43106 , \43107 , \43108 , \43109 , \43110 , \43111 , \43112 , \43113 , \43114 ,
         \43115 , \43116 , \43117 , \43118 , \43119 , \43120 , \43121 , \43122 , \43123 , \43124 ,
         \43125 , \43126 , \43127 , \43128 , \43129 , \43130 , \43131 , \43132 , \43133 , \43134 ,
         \43135 , \43136 , \43137 , \43138 , \43139 , \43140 , \43141 , \43142 , \43143 , \43144 ,
         \43145 , \43146 , \43147 , \43148 , \43149 , \43150 , \43151 , \43152 , \43153 , \43154 ,
         \43155 , \43156 , \43157 , \43158 , \43159 , \43160 , \43161 , \43162 , \43163 , \43164 ,
         \43165 , \43166 , \43167 , \43168 , \43169 , \43170 , \43171 , \43172 , \43173 , \43174 ,
         \43175 , \43176 , \43177 , \43178 , \43179 , \43180 , \43181 , \43182 , \43183 , \43184 ,
         \43185 , \43186 , \43187 , \43188 , \43189 , \43190 , \43191 , \43192 , \43193 , \43194 ,
         \43195 , \43196 , \43197 , \43198 , \43199 , \43200 , \43201 , \43202 , \43203 , \43204 ,
         \43205 , \43206 , \43207 , \43208 , \43209 , \43210 , \43211 , \43212 , \43213 , \43214 ,
         \43215 , \43216 , \43217 , \43218 , \43219 , \43220 , \43221 , \43222 , \43223 , \43224 ,
         \43225 , \43226 , \43227 , \43228 , \43229 , \43230 , \43231 , \43232 , \43233 , \43234 ,
         \43235 , \43236 , \43237 , \43238 , \43239 , \43240 , \43241 , \43242 , \43243 , \43244 ,
         \43245 , \43246 , \43247 , \43248 , \43249 , \43250 , \43251 , \43252 , \43253 , \43254 ,
         \43255 , \43256 , \43257 , \43258 , \43259 , \43260 , \43261 , \43262 , \43263 , \43264 ,
         \43265 , \43266 , \43267 , \43268 , \43269 , \43270 , \43271 , \43272 , \43273 , \43274 ,
         \43275 , \43276 , \43277 , \43278 , \43279 , \43280 , \43281 , \43282 , \43283 , \43284 ,
         \43285 , \43286 , \43287 , \43288 , \43289 , \43290 , \43291 , \43292 , \43293 , \43294 ,
         \43295 , \43296 , \43297 , \43298 , \43299 , \43300 , \43301 , \43302 , \43303 , \43304 ,
         \43305 , \43306 , \43307 , \43308 , \43309 , \43310 , \43311 , \43312 , \43313 , \43314 ,
         \43315 , \43316 , \43317 , \43318 , \43319 , \43320 , \43321 , \43322 , \43323 , \43324 ,
         \43325 , \43326 , \43327 , \43328 , \43329 , \43330 , \43331 , \43332 , \43333 , \43334 ,
         \43335 , \43336 , \43337 , \43338 , \43339 , \43340 , \43341 , \43342 , \43343 , \43344 ,
         \43345 , \43346 , \43347 , \43348 , \43349 , \43350 , \43351 , \43352 , \43353 , \43354 ,
         \43355 , \43356 , \43357 , \43358 , \43359 , \43360 , \43361 , \43362 , \43363 , \43364 ,
         \43365 , \43366 , \43367 , \43368 , \43369 , \43370 , \43371 , \43372 , \43373 , \43374 ,
         \43375 , \43376 , \43377 , \43378 , \43379 , \43380 , \43381 , \43382 , \43383 , \43384 ,
         \43385 , \43386 , \43387 , \43388 , \43389 , \43390 , \43391 , \43392 , \43393 , \43394 ,
         \43395 , \43396 , \43397 , \43398 , \43399 , \43400 , \43401 , \43402 , \43403 , \43404 ,
         \43405 , \43406 , \43407 , \43408 , \43409 , \43410 , \43411 , \43412 , \43413 , \43414 ,
         \43415 , \43416 , \43417 , \43418 , \43419 , \43420 , \43421 , \43422 , \43423 , \43424 ,
         \43425 , \43426 , \43427 , \43428 , \43429 , \43430 , \43431 , \43432 , \43433 , \43434 ,
         \43435 , \43436 , \43437 , \43438 , \43439 , \43440 , \43441 , \43442 , \43443 , \43444 ,
         \43445 , \43446 , \43447 , \43448 , \43449 , \43450 , \43451 , \43452 , \43453 , \43454 ,
         \43455 , \43456 , \43457 , \43458 , \43459 , \43460 , \43461 , \43462 , \43463 , \43464 ,
         \43465 , \43466 , \43467 , \43468 , \43469 , \43470 , \43471 , \43472 , \43473 , \43474 ,
         \43475 , \43476 , \43477 , \43478 , \43479 , \43480 , \43481 , \43482 , \43483 , \43484 ,
         \43485 , \43486 , \43487 , \43488 , \43489 , \43490 , \43491 , \43492 , \43493 , \43494 ,
         \43495 , \43496 , \43497 , \43498 , \43499 , \43500 , \43501 , \43502 , \43503 , \43504 ,
         \43505 , \43506 , \43507 , \43508 , \43509 , \43510 , \43511 , \43512 , \43513 , \43514 ,
         \43515 , \43516 , \43517 , \43518 , \43519 , \43520 , \43521 , \43522 , \43523 , \43524 ,
         \43525 , \43526 , \43527 , \43528 , \43529 , \43530 , \43531 , \43532 , \43533 , \43534 ,
         \43535 , \43536 , \43537 , \43538 , \43539 , \43540 , \43541 , \43542 , \43543 , \43544 ,
         \43545 , \43546 , \43547 , \43548 , \43549 , \43550 , \43551 , \43552 , \43553 , \43554 ,
         \43555 , \43556 , \43557 , \43558 , \43559 , \43560 , \43561 , \43562 , \43563 , \43564 ,
         \43565 , \43566 , \43567 , \43568 , \43569 , \43570 , \43571 , \43572 , \43573 , \43574 ,
         \43575 , \43576 , \43577 , \43578 , \43579 , \43580 , \43581 , \43582 , \43583 , \43584 ,
         \43585 , \43586 , \43587 , \43588 , \43589 , \43590 , \43591 , \43592 , \43593 , \43594 ,
         \43595 , \43596 , \43597 , \43598 , \43599 , \43600 , \43601 , \43602 , \43603 , \43604 ,
         \43605 , \43606 , \43607 , \43608 , \43609 , \43610 , \43611 , \43612 , \43613 , \43614 ,
         \43615 , \43616 , \43617 , \43618 , \43619 , \43620 , \43621 , \43622 , \43623 , \43624 ,
         \43625 , \43626 , \43627 , \43628 , \43629 , \43630 , \43631 , \43632 , \43633 , \43634 ,
         \43635 , \43636 , \43637 , \43638 , \43639 , \43640 , \43641 , \43642 , \43643 , \43644 ,
         \43645 , \43646 , \43647 , \43648 , \43649 , \43650 , \43651 , \43652 , \43653 , \43654 ,
         \43655 , \43656 , \43657 , \43658 , \43659 , \43660 , \43661 , \43662 , \43663 , \43664 ,
         \43665 , \43666 , \43667 , \43668 , \43669 , \43670 , \43671 , \43672 , \43673 , \43674 ,
         \43675 , \43676 , \43677 , \43678 , \43679 , \43680 , \43681 , \43682 , \43683 , \43684 ,
         \43685 , \43686 , \43687 , \43688 , \43689 , \43690 , \43691 , \43692 , \43693 , \43694 ,
         \43695 , \43696 , \43697 , \43698 , \43699 , \43700 , \43701 , \43702 , \43703 , \43704 ,
         \43705 , \43706 , \43707 , \43708 , \43709 , \43710 , \43711 , \43712 , \43713 , \43714 ,
         \43715 , \43716 , \43717 , \43718 , \43719 , \43720 , \43721 , \43722 , \43723 , \43724 ,
         \43725 , \43726 , \43727 , \43728 , \43729 , \43730 , \43731 , \43732 , \43733 , \43734 ,
         \43735 , \43736 , \43737 , \43738 , \43739 , \43740 , \43741 , \43742 , \43743 , \43744 ,
         \43745 , \43746 , \43747 , \43748 , \43749 , \43750 , \43751 , \43752 , \43753 , \43754 ,
         \43755 , \43756 , \43757 , \43758 , \43759 , \43760 , \43761 , \43762 , \43763 , \43764 ,
         \43765 , \43766 , \43767 , \43768 , \43769 , \43770 , \43771 , \43772 , \43773 , \43774 ,
         \43775 , \43776 , \43777 , \43778 , \43779 , \43780 , \43781 , \43782 , \43783 , \43784 ,
         \43785 , \43786 , \43787 , \43788 , \43789 , \43790 , \43791 , \43792 , \43793 , \43794 ,
         \43795 , \43796 , \43797 , \43798 , \43799 , \43800 , \43801 , \43802 , \43803 , \43804 ,
         \43805 , \43806 , \43807 , \43808 , \43809 , \43810 , \43811 , \43812 , \43813 , \43814 ,
         \43815 , \43816 , \43817 , \43818 , \43819 , \43820 , \43821 , \43822 , \43823 , \43824 ,
         \43825 , \43826 , \43827 , \43828 , \43829 , \43830 , \43831 , \43832 , \43833 , \43834 ,
         \43835 , \43836 , \43837 , \43838 , \43839 , \43840 , \43841 , \43842 , \43843 , \43844 ,
         \43845 , \43846 , \43847 , \43848 , \43849 , \43850 , \43851 , \43852 , \43853 , \43854 ,
         \43855 , \43856 , \43857 , \43858 , \43859 , \43860 , \43861 , \43862 , \43863 , \43864 ,
         \43865 , \43866 , \43867 , \43868 , \43869 , \43870 , \43871 , \43872 , \43873 , \43874 ,
         \43875 , \43876 , \43877 , \43878 , \43879 , \43880 , \43881 , \43882 , \43883 , \43884 ,
         \43885 , \43886 , \43887 , \43888 , \43889 , \43890 , \43891 , \43892 , \43893 , \43894 ,
         \43895 , \43896 , \43897 , \43898 , \43899 , \43900 , \43901 , \43902 , \43903 , \43904 ,
         \43905 , \43906 , \43907 , \43908 , \43909 , \43910 , \43911 , \43912 , \43913 , \43914 ,
         \43915 , \43916 , \43917 , \43918 , \43919 , \43920 , \43921 , \43922 , \43923 , \43924 ,
         \43925 , \43926 , \43927 , \43928 , \43929 , \43930 , \43931 , \43932 , \43933 , \43934 ,
         \43935 , \43936 , \43937 , \43938 , \43939 , \43940 , \43941 , \43942 , \43943 , \43944 ,
         \43945 , \43946 , \43947 , \43948 , \43949 , \43950 , \43951 , \43952 , \43953 , \43954 ,
         \43955 , \43956 , \43957 , \43958 , \43959 , \43960 , \43961 , \43962 , \43963 , \43964 ,
         \43965 , \43966 , \43967 , \43968 , \43969 , \43970 , \43971 , \43972 , \43973 , \43974 ,
         \43975 , \43976 , \43977 , \43978 , \43979 , \43980 , \43981 , \43982 , \43983 , \43984 ,
         \43985 , \43986 , \43987 , \43988 , \43989 , \43990 , \43991 , \43992 , \43993 , \43994 ,
         \43995 , \43996 , \43997 , \43998 , \43999 , \44000 , \44001 , \44002 , \44003 , \44004 ,
         \44005 , \44006 , \44007 , \44008 , \44009 , \44010 , \44011 , \44012 , \44013 , \44014 ,
         \44015 , \44016 , \44017 , \44018 , \44019 , \44020 , \44021 , \44022 , \44023 , \44024 ,
         \44025 , \44026 , \44027 , \44028 , \44029 , \44030 , \44031 , \44032 , \44033 , \44034 ,
         \44035 , \44036 , \44037 , \44038 , \44039 , \44040 , \44041 , \44042 , \44043 , \44044 ,
         \44045 , \44046 , \44047 , \44048 , \44049 , \44050 , \44051 , \44052 , \44053 , \44054 ,
         \44055 , \44056 , \44057 , \44058 , \44059 , \44060 , \44061 , \44062 , \44063 , \44064 ,
         \44065 , \44066 , \44067 , \44068 , \44069 , \44070 , \44071 , \44072 , \44073 , \44074 ,
         \44075 , \44076 , \44077 , \44078 , \44079 , \44080 , \44081 , \44082 , \44083 , \44084 ,
         \44085 , \44086 , \44087 , \44088 , \44089 , \44090 , \44091 , \44092 , \44093 , \44094 ,
         \44095 , \44096 , \44097 , \44098 , \44099 , \44100 , \44101 , \44102 , \44103 , \44104 ,
         \44105 , \44106 , \44107 , \44108 , \44109 , \44110 , \44111 , \44112 , \44113 , \44114 ,
         \44115 , \44116 , \44117 , \44118 , \44119 , \44120 , \44121 , \44122 , \44123 , \44124 ,
         \44125 , \44126 , \44127 , \44128 , \44129 , \44130 , \44131 , \44132 , \44133 , \44134 ,
         \44135 , \44136 , \44137 , \44138 , \44139 , \44140 , \44141 , \44142 , \44143 , \44144 ,
         \44145 , \44146 , \44147 , \44148 , \44149 , \44150 , \44151 , \44152 , \44153 , \44154 ,
         \44155 , \44156 , \44157 , \44158 , \44159 , \44160 , \44161 , \44162 , \44163 , \44164 ,
         \44165 , \44166 , \44167 , \44168 , \44169 , \44170 , \44171 , \44172 , \44173 , \44174 ,
         \44175 , \44176 , \44177 , \44178 , \44179 , \44180 , \44181 , \44182 , \44183 , \44184 ,
         \44185 , \44186 , \44187 , \44188 , \44189 , \44190 , \44191 , \44192 , \44193 , \44194 ,
         \44195 , \44196 , \44197 , \44198 , \44199 , \44200 , \44201 , \44202 , \44203 , \44204 ,
         \44205 , \44206 , \44207 , \44208 , \44209 , \44210 , \44211 , \44212 , \44213 , \44214 ,
         \44215 , \44216 , \44217 , \44218 , \44219 , \44220 , \44221 , \44222 , \44223 , \44224 ,
         \44225 , \44226 , \44227 , \44228 , \44229 , \44230 , \44231 , \44232 , \44233 , \44234 ,
         \44235 , \44236 , \44237 , \44238 , \44239 , \44240 , \44241 , \44242 , \44243 , \44244 ,
         \44245 , \44246 , \44247 , \44248 , \44249 , \44250 , \44251 , \44252 , \44253 , \44254 ,
         \44255 , \44256 , \44257 , \44258 , \44259 , \44260 , \44261 , \44262 , \44263 , \44264 ,
         \44265 , \44266 , \44267 , \44268 , \44269 , \44270 , \44271 , \44272 , \44273 , \44274 ,
         \44275 , \44276 , \44277 , \44278 , \44279 , \44280 , \44281 , \44282 , \44283 , \44284 ,
         \44285 , \44286 , \44287 , \44288 , \44289 , \44290 , \44291 , \44292 , \44293 , \44294 ,
         \44295 , \44296 , \44297 , \44298 , \44299 , \44300 , \44301 , \44302 , \44303 , \44304 ,
         \44305 , \44306 , \44307 , \44308 , \44309 , \44310 , \44311 , \44312 , \44313 , \44314 ,
         \44315 , \44316 , \44317 , \44318 , \44319 , \44320 , \44321 , \44322 , \44323 , \44324 ,
         \44325 , \44326 , \44327 , \44328 , \44329 , \44330 , \44331 , \44332 , \44333 , \44334 ,
         \44335 , \44336 , \44337 , \44338 , \44339 , \44340 , \44341 , \44342 , \44343 , \44344 ,
         \44345 , \44346 , \44347 , \44348 , \44349 , \44350 , \44351 , \44352 , \44353 , \44354 ,
         \44355 , \44356 , \44357 , \44358 , \44359 , \44360 , \44361 , \44362 , \44363 , \44364 ,
         \44365 , \44366 , \44367 , \44368 , \44369 , \44370 , \44371 , \44372 , \44373 , \44374 ,
         \44375 , \44376 , \44377 , \44378 , \44379 , \44380 , \44381 , \44382 , \44383 , \44384 ,
         \44385 , \44386 , \44387 , \44388 , \44389 , \44390 , \44391 , \44392 , \44393 , \44394 ,
         \44395 , \44396 , \44397 , \44398 , \44399 , \44400 , \44401 , \44402 , \44403 , \44404 ,
         \44405 , \44406 , \44407 , \44408 , \44409 , \44410 , \44411 , \44412 , \44413 , \44414 ,
         \44415 , \44416 , \44417 , \44418 , \44419 , \44420 , \44421 , \44422 , \44423 , \44424 ,
         \44425 , \44426 , \44427 , \44428 , \44429 , \44430 , \44431 , \44432 , \44433 , \44434 ,
         \44435 , \44436 , \44437 , \44438 , \44439 , \44440 , \44441 , \44442 , \44443 , \44444 ,
         \44445 , \44446 , \44447 , \44448 , \44449 , \44450 , \44451 , \44452 , \44453 , \44454 ,
         \44455 , \44456 , \44457 , \44458 , \44459 , \44460 , \44461 , \44462 , \44463 , \44464 ,
         \44465 , \44466 , \44467 , \44468 , \44469 , \44470 , \44471 , \44472 , \44473 , \44474 ,
         \44475 , \44476 , \44477 , \44478 , \44479 , \44480 , \44481 , \44482 , \44483 , \44484 ,
         \44485 , \44486 , \44487 , \44488 , \44489 , \44490 , \44491 , \44492 , \44493 , \44494 ,
         \44495 , \44496 , \44497 , \44498 , \44499 , \44500 , \44501 , \44502 , \44503 , \44504 ,
         \44505 , \44506 , \44507 , \44508 , \44509 , \44510 , \44511 , \44512 , \44513 , \44514 ,
         \44515 , \44516 , \44517 , \44518 , \44519 , \44520 , \44521 , \44522 , \44523 , \44524 ,
         \44525 , \44526 , \44527 , \44528 , \44529 , \44530 , \44531 , \44532 , \44533 , \44534 ,
         \44535 , \44536 , \44537 , \44538 , \44539 , \44540 , \44541 , \44542 , \44543 , \44544 ,
         \44545 , \44546 , \44547 , \44548 , \44549 , \44550 , \44551 , \44552 , \44553 , \44554 ,
         \44555 , \44556 , \44557 , \44558 , \44559 , \44560 , \44561 , \44562 , \44563 , \44564 ,
         \44565 , \44566 , \44567 , \44568 , \44569 , \44570 , \44571 , \44572 , \44573 , \44574 ,
         \44575 , \44576 , \44577 , \44578 , \44579 , \44580 , \44581 , \44582 , \44583 , \44584 ,
         \44585 , \44586 , \44587 , \44588 , \44589 , \44590 , \44591 , \44592 , \44593 , \44594 ,
         \44595 , \44596 , \44597 , \44598 , \44599 , \44600 , \44601 , \44602 , \44603 , \44604 ,
         \44605 , \44606 , \44607 , \44608 , \44609 , \44610 , \44611 , \44612 , \44613 , \44614 ,
         \44615 , \44616 , \44617 , \44618 , \44619 , \44620 , \44621 , \44622 , \44623 , \44624 ,
         \44625 , \44626 , \44627 , \44628 , \44629 , \44630 , \44631 , \44632 , \44633 , \44634 ,
         \44635 , \44636 , \44637 , \44638 , \44639 , \44640 , \44641 , \44642 , \44643 , \44644 ,
         \44645 , \44646 , \44647 , \44648 , \44649 , \44650 , \44651 , \44652 , \44653 , \44654 ,
         \44655 , \44656 , \44657 , \44658 , \44659 , \44660 , \44661 , \44662 , \44663 , \44664 ,
         \44665 , \44666 , \44667 , \44668 , \44669 , \44670 , \44671 , \44672 , \44673 , \44674 ,
         \44675 , \44676 , \44677 , \44678 , \44679 , \44680 , \44681 , \44682 , \44683 , \44684 ,
         \44685 , \44686 , \44687 , \44688 , \44689 , \44690 , \44691 , \44692 , \44693 , \44694 ,
         \44695 , \44696 , \44697 , \44698 , \44699 , \44700 , \44701 , \44702 , \44703 , \44704 ,
         \44705 , \44706 , \44707 , \44708 , \44709 , \44710 , \44711 , \44712 , \44713 , \44714 ,
         \44715 , \44716 , \44717 , \44718 , \44719 , \44720 , \44721 , \44722 , \44723 , \44724 ,
         \44725 , \44726 , \44727 , \44728 , \44729 , \44730 , \44731 , \44732 , \44733 , \44734 ,
         \44735 , \44736 , \44737 , \44738 , \44739 , \44740 , \44741 , \44742 , \44743 , \44744 ,
         \44745 , \44746 , \44747 , \44748 , \44749 , \44750 , \44751 , \44752 , \44753 , \44754 ,
         \44755 , \44756 , \44757 , \44758 , \44759 , \44760 , \44761 , \44762 , \44763 , \44764 ,
         \44765 , \44766 , \44767 , \44768 , \44769 , \44770 , \44771 , \44772 , \44773 , \44774 ,
         \44775 , \44776 , \44777 , \44778 , \44779 , \44780 , \44781 , \44782 , \44783 , \44784 ,
         \44785 , \44786 , \44787 , \44788 , \44789 , \44790 , \44791 , \44792 , \44793 , \44794 ,
         \44795 , \44796 , \44797 , \44798 , \44799 , \44800 , \44801 , \44802 , \44803 , \44804 ,
         \44805 , \44806 , \44807 , \44808 , \44809 , \44810 , \44811 , \44812 , \44813 , \44814 ,
         \44815 , \44816 , \44817 , \44818 , \44819 , \44820 , \44821 , \44822 , \44823 , \44824 ,
         \44825 , \44826 , \44827 , \44828 , \44829 , \44830 , \44831 , \44832 , \44833 , \44834 ,
         \44835 , \44836 , \44837 , \44838 , \44839 , \44840 , \44841 , \44842 , \44843 , \44844 ,
         \44845 , \44846 , \44847 , \44848 , \44849 , \44850 , \44851 , \44852 , \44853 , \44854 ,
         \44855 , \44856 , \44857 , \44858 , \44859 , \44860 , \44861 , \44862 , \44863 , \44864 ,
         \44865 , \44866 , \44867 , \44868 , \44869 , \44870 , \44871 , \44872 , \44873 , \44874 ,
         \44875 , \44876 , \44877 , \44878 , \44879 , \44880 , \44881 , \44882 , \44883 , \44884 ,
         \44885 , \44886 , \44887 , \44888 , \44889 , \44890 , \44891 , \44892 , \44893 , \44894 ,
         \44895 , \44896 , \44897 , \44898 , \44899 , \44900 , \44901 , \44902 , \44903 , \44904 ,
         \44905 , \44906 , \44907 , \44908 , \44909 , \44910 , \44911 , \44912 , \44913 , \44914 ,
         \44915 , \44916 , \44917 , \44918 , \44919 , \44920 , \44921 , \44922 , \44923 , \44924 ,
         \44925 , \44926 , \44927 , \44928 , \44929 , \44930 , \44931 , \44932 , \44933 , \44934 ,
         \44935 , \44936 , \44937 , \44938 , \44939 , \44940 , \44941 , \44942 , \44943 , \44944 ,
         \44945 , \44946 , \44947 , \44948 , \44949 , \44950 , \44951 , \44952 , \44953 , \44954 ,
         \44955 , \44956 , \44957 , \44958 , \44959 , \44960 , \44961 , \44962 , \44963 , \44964 ,
         \44965 , \44966 , \44967 , \44968 , \44969 , \44970 , \44971 , \44972 , \44973 , \44974 ,
         \44975 , \44976 , \44977 , \44978 , \44979 , \44980 , \44981 , \44982 , \44983 , \44984 ,
         \44985 , \44986 , \44987 , \44988 , \44989 , \44990 , \44991 , \44992 , \44993 , \44994 ,
         \44995 , \44996 , \44997 , \44998 , \44999 , \45000 , \45001 , \45002 , \45003 , \45004 ,
         \45005 , \45006 , \45007 , \45008 , \45009 , \45010 , \45011 , \45012 , \45013 , \45014 ,
         \45015 , \45016 , \45017 , \45018 , \45019 , \45020 , \45021 , \45022 , \45023 , \45024 ,
         \45025 , \45026 , \45027 , \45028 , \45029 , \45030 , \45031 , \45032 , \45033 , \45034 ,
         \45035 , \45036 , \45037 , \45038 , \45039 , \45040 , \45041 , \45042 , \45043 , \45044 ,
         \45045 , \45046 , \45047 , \45048 , \45049 , \45050 , \45051 , \45052 , \45053 , \45054 ,
         \45055 , \45056 , \45057 , \45058 , \45059 , \45060 , \45061 , \45062 , \45063 , \45064 ,
         \45065 , \45066 , \45067 , \45068 , \45069 , \45070 , \45071 , \45072 , \45073 , \45074 ,
         \45075 , \45076 , \45077 , \45078 , \45079 , \45080 , \45081 , \45082 , \45083 , \45084 ,
         \45085 , \45086 , \45087 , \45088 , \45089 , \45090 , \45091 , \45092 , \45093 , \45094 ,
         \45095 , \45096 , \45097 , \45098 , \45099 , \45100 , \45101 , \45102 , \45103 , \45104 ,
         \45105 , \45106 , \45107 , \45108 , \45109 , \45110 , \45111 , \45112 , \45113 , \45114 ,
         \45115 , \45116 , \45117 , \45118 , \45119 , \45120 , \45121 , \45122 , \45123 , \45124 ,
         \45125 , \45126 , \45127 , \45128 , \45129 , \45130 , \45131 , \45132 , \45133 , \45134 ,
         \45135 , \45136 , \45137 , \45138 , \45139 , \45140 , \45141 , \45142 , \45143 , \45144 ,
         \45145 , \45146 , \45147 , \45148 , \45149 , \45150 , \45151 , \45152 , \45153 , \45154 ,
         \45155 , \45156 , \45157 , \45158 , \45159 , \45160 , \45161 , \45162 , \45163 , \45164 ,
         \45165 , \45166 , \45167 , \45168 , \45169 , \45170 , \45171 , \45172 , \45173 , \45174 ,
         \45175 , \45176 , \45177 , \45178 , \45179 , \45180 , \45181 , \45182 , \45183 , \45184 ,
         \45185 , \45186 , \45187 , \45188 , \45189 , \45190 , \45191 , \45192 , \45193 , \45194 ,
         \45195 , \45196 , \45197 , \45198 , \45199 , \45200 , \45201 , \45202 , \45203 , \45204 ,
         \45205 , \45206 , \45207 , \45208 , \45209 , \45210 , \45211 , \45212 , \45213 , \45214 ,
         \45215 , \45216 , \45217 , \45218 , \45219 , \45220 , \45221 , \45222 , \45223 , \45224 ,
         \45225 , \45226 , \45227 , \45228 , \45229 , \45230 , \45231 , \45232 , \45233 , \45234 ,
         \45235 , \45236 , \45237 , \45238 , \45239 , \45240 , \45241 , \45242 , \45243 , \45244 ,
         \45245 , \45246 , \45247 , \45248 , \45249 , \45250 , \45251 , \45252 , \45253 , \45254 ,
         \45255 , \45256 , \45257 , \45258 , \45259 , \45260 , \45261 , \45262 , \45263 , \45264 ,
         \45265 , \45266 , \45267 , \45268 , \45269 , \45270 , \45271 , \45272 , \45273 , \45274 ,
         \45275 , \45276 , \45277 , \45278 , \45279 , \45280 , \45281 , \45282 , \45283 , \45284 ,
         \45285 , \45286 , \45287 , \45288 , \45289 , \45290 , \45291 , \45292 , \45293 , \45294 ,
         \45295 , \45296 , \45297 , \45298 , \45299 , \45300 , \45301 , \45302 , \45303 , \45304 ,
         \45305 , \45306 , \45307 , \45308 , \45309 , \45310 , \45311 , \45312 , \45313 , \45314 ,
         \45315 , \45316 , \45317 , \45318 , \45319 , \45320 , \45321 , \45322 , \45323 , \45324 ,
         \45325 , \45326 , \45327 , \45328 , \45329 , \45330 , \45331 , \45332 , \45333 , \45334 ,
         \45335 , \45336 , \45337 , \45338 , \45339 , \45340 , \45341 , \45342 , \45343 , \45344 ,
         \45345 , \45346 , \45347 , \45348 , \45349 , \45350 , \45351 , \45352 , \45353 , \45354 ,
         \45355 , \45356 , \45357 , \45358 , \45359 , \45360 , \45361 , \45362 , \45363 , \45364 ,
         \45365 , \45366 , \45367 , \45368 , \45369 , \45370 , \45371 , \45372 , \45373 , \45374 ,
         \45375 , \45376 , \45377 , \45378 , \45379 , \45380 , \45381 , \45382 , \45383 , \45384 ,
         \45385 , \45386 , \45387 , \45388 , \45389 , \45390 , \45391 , \45392 , \45393 , \45394 ,
         \45395 , \45396 , \45397 , \45398 , \45399 , \45400 , \45401 , \45402 , \45403 , \45404 ,
         \45405 , \45406 , \45407 , \45408 , \45409 , \45410 , \45411 , \45412 , \45413 , \45414 ,
         \45415 , \45416 , \45417 , \45418 , \45419 , \45420 , \45421 , \45422 , \45423 , \45424 ,
         \45425 , \45426 , \45427 , \45428 , \45429 , \45430 , \45431 , \45432 , \45433 , \45434 ,
         \45435 , \45436 , \45437 , \45438 , \45439 , \45440 , \45441 , \45442 , \45443 , \45444 ,
         \45445 , \45446 , \45447 , \45448 , \45449 , \45450 , \45451 , \45452 , \45453 , \45454 ,
         \45455 , \45456 , \45457 , \45458 , \45459 , \45460 , \45461 , \45462 , \45463 , \45464 ,
         \45465 , \45466 , \45467 , \45468 , \45469 , \45470 , \45471 , \45472 , \45473 , \45474 ,
         \45475 , \45476 , \45477 , \45478 , \45479 , \45480 , \45481 , \45482 , \45483 , \45484 ,
         \45485 , \45486 , \45487 , \45488 , \45489 , \45490 , \45491 , \45492 , \45493 , \45494 ,
         \45495 , \45496 , \45497 , \45498 , \45499 , \45500 , \45501 , \45502 , \45503 , \45504 ,
         \45505 , \45506 , \45507 , \45508 , \45509 , \45510 , \45511 , \45512 , \45513 , \45514 ,
         \45515 , \45516 , \45517 , \45518 , \45519 , \45520 , \45521 , \45522 , \45523 , \45524 ,
         \45525 , \45526 , \45527 , \45528 , \45529 , \45530 , \45531 , \45532 , \45533 , \45534 ,
         \45535 , \45536 , \45537 , \45538 , \45539 , \45540 , \45541 , \45542 , \45543 , \45544 ,
         \45545 , \45546 , \45547 , \45548 , \45549 , \45550 , \45551 , \45552 , \45553 , \45554 ,
         \45555 , \45556 , \45557 , \45558 , \45559 , \45560 , \45561 , \45562 , \45563 , \45564 ,
         \45565 , \45566 , \45567 , \45568 , \45569 , \45570 , \45571 , \45572 , \45573 , \45574 ,
         \45575 , \45576 , \45577 , \45578 , \45579 , \45580 , \45581 , \45582 , \45583 , \45584 ,
         \45585 , \45586 , \45587 , \45588 , \45589 , \45590 , \45591 , \45592 , \45593 , \45594 ,
         \45595 , \45596 , \45597 , \45598 , \45599 , \45600 , \45601 , \45602 , \45603 , \45604 ,
         \45605 , \45606 , \45607 , \45608 , \45609 , \45610 , \45611 , \45612 , \45613 , \45614 ,
         \45615 , \45616 , \45617 , \45618 , \45619 , \45620 , \45621 , \45622 , \45623 , \45624 ,
         \45625 , \45626 , \45627 , \45628 , \45629 , \45630 , \45631 , \45632 , \45633 , \45634 ,
         \45635 , \45636 , \45637 , \45638 , \45639 , \45640 , \45641 , \45642 , \45643 , \45644 ,
         \45645 , \45646 , \45647 , \45648 , \45649 , \45650 , \45651 , \45652 , \45653 , \45654 ,
         \45655 , \45656 , \45657 , \45658 , \45659 , \45660 , \45661 , \45662 , \45663 , \45664 ,
         \45665 , \45666 , \45667 , \45668 , \45669 , \45670 , \45671 , \45672 , \45673 , \45674 ,
         \45675 , \45676 , \45677 , \45678 , \45679 , \45680 , \45681 , \45682 , \45683 , \45684 ,
         \45685 , \45686 , \45687 , \45688 , \45689 , \45690 , \45691 , \45692 , \45693 , \45694 ,
         \45695 , \45696 , \45697 , \45698 , \45699 , \45700 , \45701 , \45702 , \45703 , \45704 ,
         \45705 , \45706 , \45707 , \45708 , \45709 , \45710 , \45711 , \45712 , \45713 , \45714 ,
         \45715 , \45716 , \45717 , \45718 , \45719 , \45720 , \45721 , \45722 , \45723 , \45724 ,
         \45725 , \45726 , \45727 , \45728 , \45729 , \45730 , \45731 , \45732 , \45733 , \45734 ,
         \45735 , \45736 , \45737 , \45738 , \45739 , \45740 , \45741 , \45742 , \45743 , \45744 ,
         \45745 , \45746 , \45747 , \45748 , \45749 , \45750 , \45751 , \45752 , \45753 , \45754 ,
         \45755 , \45756 , \45757 , \45758 , \45759 , \45760 , \45761 , \45762 , \45763 , \45764 ,
         \45765 , \45766 , \45767 , \45768 , \45769 , \45770 , \45771 , \45772 , \45773 , \45774 ,
         \45775 , \45776 , \45777 , \45778 , \45779 , \45780 , \45781 , \45782 , \45783 , \45784 ,
         \45785 , \45786 , \45787 , \45788 , \45789 , \45790 , \45791 , \45792 , \45793 , \45794 ,
         \45795 , \45796 , \45797 , \45798 , \45799 , \45800 , \45801 , \45802 , \45803 , \45804 ,
         \45805 , \45806 , \45807 , \45808 , \45809 , \45810 , \45811 , \45812 , \45813 , \45814 ,
         \45815 , \45816 , \45817 , \45818 , \45819 , \45820 , \45821 , \45822 , \45823 , \45824 ,
         \45825 , \45826 , \45827 , \45828 , \45829 , \45830 , \45831 , \45832 , \45833 , \45834 ,
         \45835 , \45836 , \45837 , \45838 , \45839 , \45840 , \45841 , \45842 , \45843 , \45844 ,
         \45845 , \45846 , \45847 , \45848 , \45849 , \45850 , \45851 , \45852 , \45853 , \45854 ,
         \45855 , \45856 , \45857 , \45858 , \45859 , \45860 , \45861 , \45862 , \45863 , \45864 ,
         \45865 , \45866 , \45867 , \45868 , \45869 , \45870 , \45871 , \45872 , \45873 , \45874 ,
         \45875 , \45876 , \45877 , \45878 , \45879 , \45880 , \45881 , \45882 , \45883 , \45884 ,
         \45885 , \45886 , \45887 , \45888 , \45889 , \45890 , \45891 , \45892 , \45893 , \45894 ,
         \45895 , \45896 , \45897 , \45898 , \45899 , \45900 , \45901 , \45902 , \45903 , \45904 ,
         \45905 , \45906 , \45907 , \45908 , \45909 , \45910 , \45911 , \45912 , \45913 , \45914 ,
         \45915 , \45916 , \45917 , \45918 , \45919 , \45920 , \45921 , \45922 , \45923 , \45924 ,
         \45925 , \45926 , \45927 , \45928 , \45929 , \45930 , \45931 , \45932 , \45933 , \45934 ,
         \45935 , \45936 , \45937 , \45938 , \45939 , \45940 , \45941 , \45942 , \45943 , \45944 ,
         \45945 , \45946 , \45947 , \45948 , \45949 , \45950 , \45951 , \45952 , \45953 , \45954 ,
         \45955 , \45956 , \45957 , \45958 , \45959 , \45960 , \45961 , \45962 , \45963 , \45964 ,
         \45965 , \45966 , \45967 , \45968 , \45969 , \45970 , \45971 , \45972 , \45973 , \45974 ,
         \45975 , \45976 , \45977 , \45978 , \45979 , \45980 , \45981 , \45982 , \45983 , \45984 ,
         \45985 , \45986 , \45987 , \45988 , \45989 , \45990 , \45991 , \45992 , \45993 , \45994 ,
         \45995 , \45996 , \45997 , \45998 , \45999 , \46000 , \46001 , \46002 , \46003 , \46004 ,
         \46005 , \46006 , \46007 , \46008 , \46009 , \46010 , \46011 , \46012 , \46013 , \46014 ,
         \46015 , \46016 , \46017 , \46018 , \46019 , \46020 , \46021 , \46022 , \46023 , \46024 ,
         \46025 , \46026 , \46027 , \46028 , \46029 , \46030 , \46031 , \46032 , \46033 , \46034 ,
         \46035 , \46036 , \46037 , \46038 , \46039 , \46040 , \46041 , \46042 , \46043 , \46044 ,
         \46045 , \46046 , \46047 , \46048 , \46049 , \46050 , \46051 , \46052 , \46053 , \46054 ,
         \46055 , \46056 , \46057 , \46058 , \46059 , \46060 , \46061 , \46062 , \46063 , \46064 ,
         \46065 , \46066 , \46067 , \46068 , \46069 , \46070 , \46071 , \46072 , \46073 , \46074 ,
         \46075 , \46076 , \46077 , \46078 , \46079 , \46080 , \46081 , \46082 , \46083 , \46084 ,
         \46085 , \46086 , \46087 , \46088 , \46089 , \46090 , \46091 , \46092 , \46093 , \46094 ,
         \46095 , \46096 , \46097 , \46098 , \46099 , \46100 , \46101 , \46102 , \46103 , \46104 ,
         \46105 , \46106 , \46107 , \46108 , \46109 , \46110 , \46111 , \46112 , \46113 , \46114 ,
         \46115 , \46116 , \46117 , \46118 , \46119 , \46120 , \46121 , \46122 , \46123 , \46124 ,
         \46125 , \46126 , \46127 , \46128 , \46129 , \46130 , \46131 , \46132 , \46133 , \46134 ,
         \46135 , \46136 , \46137 , \46138 , \46139 , \46140 , \46141 , \46142 , \46143 , \46144 ,
         \46145 , \46146 , \46147 , \46148 , \46149 , \46150 , \46151 , \46152 , \46153 , \46154 ,
         \46155 , \46156 , \46157 , \46158 , \46159 , \46160 , \46161 , \46162 , \46163 , \46164 ,
         \46165 , \46166 , \46167 , \46168 , \46169 , \46170 , \46171 , \46172 , \46173 , \46174 ,
         \46175 , \46176 , \46177 , \46178 , \46179 , \46180 , \46181 , \46182 , \46183 , \46184 ,
         \46185 , \46186 , \46187 , \46188 , \46189 , \46190 , \46191 , \46192 , \46193 , \46194 ,
         \46195 , \46196 , \46197 , \46198 , \46199 , \46200 , \46201 , \46202 , \46203 , \46204 ,
         \46205 , \46206 , \46207 , \46208 , \46209 , \46210 , \46211 , \46212 , \46213 , \46214 ,
         \46215 , \46216 , \46217 , \46218 , \46219 , \46220 , \46221 , \46222 , \46223 , \46224 ,
         \46225 , \46226 , \46227 , \46228 , \46229 , \46230 , \46231 , \46232 , \46233 , \46234 ,
         \46235 , \46236 , \46237 , \46238 , \46239 , \46240 , \46241 , \46242 , \46243 , \46244 ,
         \46245 , \46246 , \46247 , \46248 , \46249 , \46250 , \46251 , \46252 , \46253 , \46254 ,
         \46255 , \46256 , \46257 , \46258 , \46259 , \46260 , \46261 , \46262 , \46263 , \46264 ,
         \46265 , \46266 , \46267 , \46268 , \46269 , \46270 , \46271 , \46272 , \46273 , \46274 ,
         \46275 , \46276 , \46277 , \46278 , \46279 , \46280 , \46281 , \46282 , \46283 , \46284 ,
         \46285 , \46286 , \46287 , \46288 , \46289 , \46290 , \46291 , \46292 , \46293 , \46294 ,
         \46295 , \46296 , \46297 , \46298 , \46299 , \46300 , \46301 , \46302 , \46303 , \46304 ,
         \46305 , \46306 , \46307 , \46308 , \46309 , \46310 , \46311 , \46312 , \46313 , \46314 ,
         \46315 , \46316 , \46317 , \46318 , \46319 , \46320 , \46321 , \46322 , \46323 , \46324 ,
         \46325 , \46326 , \46327 , \46328 , \46329 , \46330 , \46331 , \46332 , \46333 , \46334 ,
         \46335 , \46336 , \46337 , \46338 , \46339 , \46340 , \46341 , \46342 , \46343 , \46344 ,
         \46345 , \46346 , \46347 , \46348 , \46349 , \46350 , \46351 , \46352 , \46353 , \46354 ,
         \46355 , \46356 , \46357 , \46358 , \46359 , \46360 , \46361 , \46362 , \46363 , \46364 ,
         \46365 , \46366 , \46367 , \46368 , \46369 , \46370 , \46371 , \46372 , \46373 , \46374 ,
         \46375 , \46376 , \46377 , \46378 , \46379 , \46380 , \46381 , \46382 , \46383 , \46384 ,
         \46385 , \46386 , \46387 , \46388 , \46389 , \46390 , \46391 , \46392 , \46393 , \46394 ,
         \46395 , \46396 , \46397 , \46398 , \46399 , \46400 , \46401 , \46402 , \46403 , \46404 ,
         \46405 , \46406 , \46407 , \46408 , \46409 , \46410 , \46411 , \46412 , \46413 , \46414 ,
         \46415 , \46416 , \46417 , \46418 , \46419 , \46420 , \46421 , \46422 , \46423 , \46424 ,
         \46425 , \46426 , \46427 , \46428 , \46429 , \46430 , \46431 , \46432 , \46433 , \46434 ,
         \46435 , \46436 , \46437 , \46438 , \46439 , \46440 , \46441 , \46442 , \46443 , \46444 ,
         \46445 , \46446 , \46447 , \46448 , \46449 , \46450 , \46451 , \46452 , \46453 , \46454 ,
         \46455 , \46456 , \46457 , \46458 , \46459 , \46460 , \46461 , \46462 , \46463 , \46464 ,
         \46465 , \46466 , \46467 , \46468 , \46469 , \46470 , \46471 , \46472 , \46473 , \46474 ,
         \46475 , \46476 , \46477 , \46478 , \46479 , \46480 , \46481 , \46482 , \46483 , \46484 ,
         \46485 , \46486 , \46487 , \46488 , \46489 , \46490 , \46491 , \46492 , \46493 , \46494 ,
         \46495 , \46496 , \46497 , \46498 , \46499 , \46500 , \46501 , \46502 , \46503 , \46504 ,
         \46505 , \46506 , \46507 , \46508 , \46509 , \46510 , \46511 , \46512 , \46513 , \46514 ,
         \46515 , \46516 , \46517 , \46518 , \46519 , \46520 , \46521 , \46522 , \46523 , \46524 ,
         \46525 , \46526 , \46527 , \46528 , \46529 , \46530 , \46531 , \46532 , \46533 , \46534 ,
         \46535 , \46536 , \46537 , \46538 , \46539 , \46540 , \46541 , \46542 , \46543 , \46544 ,
         \46545 , \46546 , \46547 , \46548 , \46549 , \46550 , \46551 , \46552 , \46553 , \46554 ,
         \46555 , \46556 , \46557 , \46558 , \46559 , \46560 , \46561 , \46562 , \46563 , \46564 ,
         \46565 , \46566 , \46567 , \46568 , \46569 , \46570 , \46571 , \46572 , \46573 , \46574 ,
         \46575 , \46576 , \46577 , \46578 , \46579 , \46580 , \46581 , \46582 , \46583 , \46584 ,
         \46585 , \46586 , \46587 , \46588 , \46589 , \46590 , \46591 , \46592 , \46593 , \46594 ,
         \46595 , \46596 , \46597 , \46598 , \46599 , \46600 , \46601 , \46602 , \46603 , \46604 ,
         \46605 , \46606 , \46607 , \46608 , \46609 , \46610 , \46611 , \46612 , \46613 , \46614 ,
         \46615 , \46616 , \46617 , \46618 , \46619 , \46620 , \46621 , \46622 , \46623 , \46624 ,
         \46625 , \46626 , \46627 , \46628 , \46629 , \46630 , \46631 , \46632 , \46633 , \46634 ,
         \46635 , \46636 , \46637 , \46638 , \46639 , \46640 , \46641 , \46642 , \46643 , \46644 ,
         \46645 , \46646 , \46647 , \46648 , \46649 , \46650 , \46651 , \46652 , \46653 , \46654 ,
         \46655 , \46656 , \46657 , \46658 , \46659 , \46660 , \46661 , \46662 , \46663 , \46664 ,
         \46665 , \46666 , \46667 , \46668 , \46669 , \46670 , \46671 , \46672 , \46673 , \46674 ,
         \46675 , \46676 , \46677 , \46678 , \46679 , \46680 , \46681 , \46682 , \46683 , \46684 ,
         \46685 , \46686 , \46687 , \46688 , \46689 , \46690 , \46691 , \46692 , \46693 , \46694 ,
         \46695 , \46696 , \46697 , \46698 , \46699 , \46700 , \46701 , \46702 , \46703 , \46704 ,
         \46705 , \46706 , \46707 , \46708 , \46709 , \46710 , \46711 , \46712 , \46713 , \46714 ,
         \46715 , \46716 , \46717 , \46718 , \46719 , \46720 , \46721 , \46722 , \46723 , \46724 ,
         \46725 , \46726 , \46727 , \46728 , \46729 , \46730 , \46731 , \46732 , \46733 , \46734 ,
         \46735 , \46736 , \46737 , \46738 , \46739 , \46740 , \46741 , \46742 , \46743 , \46744 ,
         \46745 , \46746 , \46747 , \46748 , \46749 , \46750 , \46751 , \46752 , \46753 , \46754 ,
         \46755 , \46756 , \46757 , \46758 , \46759 , \46760 , \46761 , \46762 , \46763 , \46764 ,
         \46765 , \46766 , \46767 , \46768 , \46769 , \46770 , \46771 , \46772 , \46773 , \46774 ,
         \46775 , \46776 , \46777 , \46778 , \46779 , \46780 , \46781 , \46782 , \46783 , \46784 ,
         \46785 , \46786 , \46787 , \46788 , \46789 , \46790 , \46791 , \46792 , \46793 , \46794 ,
         \46795 , \46796 , \46797 , \46798 , \46799 , \46800 , \46801 , \46802 , \46803 , \46804 ,
         \46805 , \46806 , \46807 , \46808 , \46809 , \46810 , \46811 , \46812 , \46813 , \46814 ,
         \46815 , \46816 , \46817 , \46818 , \46819 , \46820 , \46821 , \46822 , \46823 , \46824 ,
         \46825 , \46826 , \46827 , \46828 , \46829 , \46830 , \46831 , \46832 , \46833 , \46834 ,
         \46835 , \46836 , \46837 , \46838 , \46839 , \46840 , \46841 , \46842 , \46843 , \46844 ,
         \46845 , \46846 , \46847 , \46848 , \46849 , \46850 , \46851 , \46852 , \46853 , \46854 ,
         \46855 , \46856 , \46857 , \46858 , \46859 , \46860 , \46861 , \46862 , \46863 , \46864 ,
         \46865 , \46866 , \46867 , \46868 , \46869 , \46870 , \46871 , \46872 , \46873 , \46874 ,
         \46875 , \46876 , \46877 , \46878 , \46879 , \46880 , \46881 , \46882 , \46883 , \46884 ,
         \46885 , \46886 , \46887 , \46888 , \46889 , \46890 , \46891 , \46892 , \46893 , \46894 ,
         \46895 , \46896 , \46897 , \46898 , \46899 , \46900 , \46901 , \46902 , \46903 , \46904 ,
         \46905 , \46906 , \46907 , \46908 , \46909 , \46910 , \46911 , \46912 , \46913 , \46914 ,
         \46915 , \46916 , \46917 , \46918 , \46919 , \46920 , \46921 , \46922 , \46923 , \46924 ,
         \46925 , \46926 , \46927 , \46928 , \46929 , \46930 , \46931 , \46932 , \46933 , \46934 ,
         \46935 , \46936 , \46937 , \46938 , \46939 , \46940 , \46941 , \46942 , \46943 , \46944 ,
         \46945 , \46946 , \46947 , \46948 , \46949 , \46950 , \46951 , \46952 , \46953 , \46954 ,
         \46955 , \46956 , \46957 , \46958 , \46959 , \46960 , \46961 , \46962 , \46963 , \46964 ,
         \46965 , \46966 , \46967 , \46968 , \46969 , \46970 , \46971 , \46972 , \46973 , \46974 ,
         \46975 , \46976 , \46977 , \46978 , \46979 , \46980 , \46981 , \46982 , \46983 , \46984 ,
         \46985 , \46986 , \46987 , \46988 , \46989 , \46990 , \46991 , \46992 , \46993 , \46994 ,
         \46995 , \46996 , \46997 , \46998 , \46999 , \47000 , \47001 , \47002 , \47003 , \47004 ,
         \47005 , \47006 , \47007 , \47008 , \47009 , \47010 , \47011 , \47012 , \47013 , \47014 ,
         \47015 , \47016 , \47017 , \47018 , \47019 , \47020 , \47021 , \47022 , \47023 , \47024 ,
         \47025 , \47026 , \47027 , \47028 , \47029 , \47030 , \47031 , \47032 , \47033 , \47034 ,
         \47035 , \47036 , \47037 , \47038 , \47039 , \47040 , \47041 , \47042 , \47043 , \47044 ,
         \47045 , \47046 , \47047 , \47048 , \47049 , \47050 , \47051 , \47052 , \47053 , \47054 ,
         \47055 , \47056 , \47057 , \47058 , \47059 , \47060 , \47061 , \47062 , \47063 , \47064 ,
         \47065 , \47066 , \47067 , \47068 , \47069 , \47070 , \47071 , \47072 , \47073 , \47074 ,
         \47075 , \47076 , \47077 , \47078 , \47079 , \47080 , \47081 , \47082 , \47083 , \47084 ,
         \47085 , \47086 , \47087 , \47088 , \47089 , \47090 , \47091 , \47092 , \47093 , \47094 ,
         \47095 , \47096 , \47097 , \47098 , \47099 , \47100 , \47101 , \47102 , \47103 , \47104 ,
         \47105 , \47106 , \47107 , \47108 , \47109 , \47110 , \47111 , \47112 , \47113 , \47114 ,
         \47115 , \47116 , \47117 , \47118 , \47119 , \47120 , \47121 , \47122 , \47123 , \47124 ,
         \47125 , \47126 , \47127 , \47128 , \47129 , \47130 , \47131 , \47132 , \47133 , \47134 ,
         \47135 , \47136 , \47137 , \47138 , \47139 , \47140 , \47141 , \47142 , \47143 , \47144 ,
         \47145 , \47146 , \47147 , \47148 , \47149 , \47150 , \47151 , \47152 , \47153 , \47154 ,
         \47155 , \47156 , \47157 , \47158 , \47159 , \47160 , \47161 , \47162 , \47163 , \47164 ,
         \47165 , \47166 , \47167 , \47168 , \47169 , \47170 , \47171 , \47172 , \47173 , \47174 ,
         \47175 , \47176 , \47177 , \47178 , \47179 , \47180 , \47181 , \47182 , \47183 , \47184 ,
         \47185 , \47186 , \47187 , \47188 , \47189 , \47190 , \47191 , \47192 , \47193 , \47194 ,
         \47195 , \47196 , \47197 , \47198 , \47199 , \47200 , \47201 , \47202 , \47203 , \47204 ,
         \47205 , \47206 , \47207 , \47208 , \47209 , \47210 , \47211 , \47212 , \47213 , \47214 ,
         \47215 , \47216 , \47217 , \47218 , \47219 , \47220 , \47221 , \47222 , \47223 , \47224 ,
         \47225 , \47226 , \47227 , \47228 , \47229 , \47230 , \47231 , \47232 , \47233 , \47234 ,
         \47235 , \47236 , \47237 , \47238 , \47239 , \47240 , \47241 , \47242 , \47243 , \47244 ,
         \47245 , \47246 , \47247 , \47248 , \47249 , \47250 , \47251 , \47252 , \47253 , \47254 ,
         \47255 , \47256 , \47257 , \47258 , \47259 , \47260 , \47261 , \47262 , \47263 , \47264 ,
         \47265 , \47266 , \47267 , \47268 , \47269 , \47270 , \47271 , \47272 , \47273 , \47274 ,
         \47275 , \47276 , \47277 , \47278 , \47279 , \47280 , \47281 , \47282 , \47283 , \47284 ,
         \47285 , \47286 , \47287 , \47288 , \47289 , \47290 , \47291 , \47292 , \47293 , \47294 ,
         \47295 , \47296 , \47297 , \47298 , \47299 , \47300 , \47301 , \47302 , \47303 , \47304 ,
         \47305 , \47306 , \47307 , \47308 , \47309 , \47310 , \47311 , \47312 , \47313 , \47314 ,
         \47315 , \47316 , \47317 , \47318 , \47319 , \47320 , \47321 , \47322 , \47323 , \47324 ,
         \47325 , \47326 , \47327 , \47328 , \47329 , \47330 , \47331 , \47332 , \47333 , \47334 ,
         \47335 , \47336 , \47337 , \47338 , \47339 , \47340 , \47341 , \47342 , \47343 , \47344 ,
         \47345 , \47346 , \47347 , \47348 , \47349 , \47350 , \47351 , \47352 , \47353 , \47354 ,
         \47355 , \47356 , \47357 , \47358 , \47359 , \47360 , \47361 , \47362 , \47363 , \47364 ,
         \47365 , \47366 , \47367 , \47368 , \47369 , \47370 , \47371 , \47372 , \47373 , \47374 ,
         \47375 , \47376 , \47377 , \47378 , \47379 , \47380 , \47381 , \47382 , \47383 , \47384 ,
         \47385 , \47386 , \47387 , \47388 , \47389 , \47390 , \47391 , \47392 , \47393 , \47394 ,
         \47395 , \47396 , \47397 , \47398 , \47399 , \47400 , \47401 , \47402 , \47403 , \47404 ,
         \47405 , \47406 , \47407 , \47408 , \47409 , \47410 , \47411 , \47412 , \47413 , \47414 ,
         \47415 , \47416 , \47417 , \47418 , \47419 , \47420 , \47421 , \47422 , \47423 , \47424 ,
         \47425 , \47426 , \47427 , \47428 , \47429 , \47430 , \47431 , \47432 , \47433 , \47434 ,
         \47435 , \47436 , \47437 , \47438 , \47439 , \47440 , \47441 , \47442 , \47443 , \47444 ,
         \47445 , \47446 , \47447 , \47448 , \47449 , \47450 , \47451 , \47452 , \47453 , \47454 ,
         \47455 , \47456 , \47457 , \47458 , \47459 , \47460 , \47461 , \47462 , \47463 , \47464 ,
         \47465 , \47466 , \47467 , \47468 , \47469 , \47470 , \47471 , \47472 , \47473 , \47474 ,
         \47475 , \47476 , \47477 , \47478 , \47479 , \47480 , \47481 , \47482 , \47483 , \47484 ,
         \47485 , \47486 , \47487 , \47488 , \47489 , \47490 , \47491 , \47492 , \47493 , \47494 ,
         \47495 , \47496 , \47497 , \47498 , \47499 , \47500 , \47501 , \47502 , \47503 , \47504 ,
         \47505 , \47506 , \47507 , \47508 , \47509 , \47510 , \47511 , \47512 , \47513 , \47514 ,
         \47515 , \47516 , \47517 , \47518 , \47519 , \47520 , \47521 , \47522 , \47523 , \47524 ,
         \47525 , \47526 , \47527 , \47528 , \47529 , \47530 , \47531 , \47532 , \47533 , \47534 ,
         \47535 , \47536 , \47537 , \47538 , \47539 , \47540 , \47541 , \47542 , \47543 , \47544 ,
         \47545 , \47546 , \47547 , \47548 , \47549 , \47550 , \47551 , \47552 , \47553 , \47554 ,
         \47555 , \47556 , \47557 , \47558 , \47559 , \47560 , \47561 , \47562 , \47563 , \47564 ,
         \47565 , \47566 , \47567 , \47568 , \47569 , \47570 , \47571 , \47572 , \47573 , \47574 ,
         \47575 , \47576 , \47577 , \47578 , \47579 , \47580 , \47581 , \47582 , \47583 , \47584 ,
         \47585 , \47586 , \47587 , \47588 , \47589 , \47590 , \47591 , \47592 , \47593 , \47594 ,
         \47595 , \47596 , \47597 , \47598 , \47599 , \47600 , \47601 , \47602 , \47603 , \47604 ,
         \47605 , \47606 , \47607 , \47608 , \47609 , \47610 , \47611 , \47612 , \47613 , \47614 ,
         \47615 , \47616 , \47617 , \47618 , \47619 , \47620 , \47621 , \47622 , \47623 , \47624 ,
         \47625 , \47626 , \47627 , \47628 , \47629 , \47630 , \47631 , \47632 , \47633 , \47634 ,
         \47635 , \47636 , \47637 , \47638 , \47639 , \47640 , \47641 , \47642 , \47643 , \47644 ,
         \47645 , \47646 , \47647 , \47648 , \47649 , \47650 , \47651 , \47652 , \47653 , \47654 ,
         \47655 , \47656 , \47657 , \47658 , \47659 , \47660 , \47661 , \47662 , \47663 , \47664 ,
         \47665 , \47666 , \47667 , \47668 , \47669 , \47670 , \47671 , \47672 , \47673 , \47674 ,
         \47675 , \47676 , \47677 , \47678 , \47679 , \47680 , \47681 , \47682 , \47683 , \47684 ,
         \47685 , \47686 , \47687 , \47688 , \47689 , \47690 , \47691 , \47692 , \47693 , \47694 ,
         \47695 , \47696 , \47697 , \47698 , \47699 , \47700 , \47701 , \47702 , \47703 , \47704 ,
         \47705 , \47706 , \47707 , \47708 , \47709 , \47710 , \47711 , \47712 , \47713 , \47714 ,
         \47715 , \47716 , \47717 , \47718 , \47719 , \47720 , \47721 , \47722 , \47723 , \47724 ,
         \47725 , \47726 , \47727 , \47728 , \47729 , \47730 , \47731 , \47732 , \47733 , \47734 ,
         \47735 , \47736 , \47737 , \47738 , \47739 , \47740 , \47741 , \47742 , \47743 , \47744 ,
         \47745 , \47746 , \47747 , \47748 , \47749 , \47750 , \47751 , \47752 , \47753 , \47754 ,
         \47755 , \47756 , \47757 , \47758 , \47759 , \47760 , \47761 , \47762 , \47763 , \47764 ,
         \47765 , \47766 , \47767 , \47768 , \47769 , \47770 , \47771 , \47772 , \47773 , \47774 ,
         \47775 , \47776 , \47777 , \47778 , \47779 , \47780 , \47781 , \47782 , \47783 , \47784 ,
         \47785 , \47786 , \47787 , \47788 , \47789 , \47790 , \47791 , \47792 , \47793 , \47794 ,
         \47795 , \47796 , \47797 , \47798 , \47799 , \47800 , \47801 , \47802 , \47803 , \47804 ,
         \47805 , \47806 , \47807 , \47808 , \47809 , \47810 , \47811 , \47812 , \47813 , \47814 ,
         \47815 , \47816 , \47817 , \47818 , \47819 , \47820 , \47821 , \47822 , \47823 , \47824 ,
         \47825 , \47826 , \47827 , \47828 , \47829 , \47830 , \47831 , \47832 , \47833 , \47834 ,
         \47835 , \47836 , \47837 , \47838 , \47839 , \47840 , \47841 , \47842 , \47843 , \47844 ,
         \47845 , \47846 , \47847 , \47848 , \47849 , \47850 , \47851 , \47852 , \47853 , \47854 ,
         \47855 , \47856 , \47857 , \47858 , \47859 , \47860 , \47861 , \47862 , \47863 , \47864 ,
         \47865 , \47866 , \47867 , \47868 , \47869 , \47870 , \47871 , \47872 , \47873 , \47874 ,
         \47875 , \47876 , \47877 , \47878 , \47879 , \47880 , \47881 , \47882 , \47883 , \47884 ,
         \47885 , \47886 , \47887 , \47888 , \47889 , \47890 , \47891 , \47892 , \47893 , \47894 ,
         \47895 , \47896 , \47897 , \47898 , \47899 , \47900 , \47901 , \47902 , \47903 , \47904 ,
         \47905 , \47906 , \47907 , \47908 , \47909 , \47910 , \47911 , \47912 , \47913 , \47914 ,
         \47915 , \47916 , \47917 , \47918 , \47919 , \47920 , \47921 , \47922 , \47923 , \47924 ,
         \47925 , \47926 , \47927 , \47928 , \47929 , \47930 , \47931 , \47932 , \47933 , \47934 ,
         \47935 , \47936 , \47937 , \47938 , \47939 , \47940 , \47941 , \47942 , \47943 , \47944 ,
         \47945 , \47946 , \47947 , \47948 , \47949 , \47950 , \47951 , \47952 , \47953 , \47954 ,
         \47955 , \47956 , \47957 , \47958 , \47959 , \47960 , \47961 , \47962 , \47963 , \47964 ,
         \47965 , \47966 , \47967 , \47968 , \47969 , \47970 , \47971 , \47972 , \47973 , \47974 ,
         \47975 , \47976 , \47977 , \47978 , \47979 , \47980 , \47981 , \47982 , \47983 , \47984 ,
         \47985 , \47986 , \47987 , \47988 , \47989 , \47990 , \47991 , \47992 , \47993 , \47994 ,
         \47995 , \47996 , \47997 , \47998 , \47999 , \48000 , \48001 , \48002 , \48003 , \48004 ,
         \48005 , \48006 , \48007 , \48008 , \48009 , \48010 , \48011 , \48012 , \48013 , \48014 ,
         \48015 , \48016 , \48017 , \48018 , \48019 , \48020 , \48021 , \48022 , \48023 , \48024 ,
         \48025 , \48026 , \48027 , \48028 , \48029 , \48030 , \48031 , \48032 , \48033 , \48034 ,
         \48035 , \48036 , \48037 , \48038 , \48039 , \48040 , \48041 , \48042 , \48043 , \48044 ,
         \48045 , \48046 , \48047 , \48048 , \48049 , \48050 , \48051 , \48052 , \48053 , \48054 ,
         \48055 , \48056 , \48057 , \48058 , \48059 , \48060 , \48061 , \48062 , \48063 , \48064 ,
         \48065 , \48066 , \48067 , \48068 , \48069 , \48070 , \48071 , \48072 , \48073 , \48074 ,
         \48075 , \48076 , \48077 , \48078 , \48079 , \48080 , \48081 , \48082 , \48083 , \48084 ,
         \48085 , \48086 , \48087 , \48088 , \48089 , \48090 , \48091 , \48092 , \48093 , \48094 ,
         \48095 , \48096 , \48097 , \48098 , \48099 , \48100 , \48101 , \48102 , \48103 , \48104 ,
         \48105 , \48106 , \48107 , \48108 , \48109 , \48110 , \48111 , \48112 , \48113 , \48114 ,
         \48115 , \48116 , \48117 , \48118 , \48119 , \48120 , \48121 , \48122 , \48123 , \48124 ,
         \48125 , \48126 , \48127 , \48128 , \48129 , \48130 , \48131 , \48132 , \48133 , \48134 ,
         \48135 , \48136 , \48137 , \48138 , \48139 , \48140 , \48141 , \48142 , \48143 , \48144 ,
         \48145 , \48146 , \48147 , \48148 , \48149 , \48150 , \48151 , \48152 , \48153 , \48154 ,
         \48155 , \48156 , \48157 , \48158 , \48159 , \48160 , \48161 , \48162 , \48163 , \48164 ,
         \48165 , \48166 , \48167 , \48168 , \48169 , \48170 , \48171 , \48172 , \48173 , \48174 ,
         \48175 , \48176 , \48177 , \48178 , \48179 , \48180 , \48181 , \48182 , \48183 , \48184 ,
         \48185 , \48186 , \48187 , \48188 , \48189 , \48190 , \48191 , \48192 , \48193 , \48194 ,
         \48195 , \48196 , \48197 , \48198 , \48199 , \48200 , \48201 , \48202 , \48203 , \48204 ,
         \48205 , \48206 , \48207 , \48208 , \48209 , \48210 , \48211 , \48212 , \48213 , \48214 ,
         \48215 , \48216 , \48217 , \48218 , \48219 , \48220 , \48221 , \48222 , \48223 , \48224 ,
         \48225 , \48226 , \48227 , \48228 , \48229 , \48230 , \48231 , \48232 , \48233 , \48234 ,
         \48235 , \48236 , \48237 , \48238 , \48239 , \48240 , \48241 , \48242 , \48243 , \48244 ,
         \48245 , \48246 , \48247 , \48248 , \48249 , \48250 , \48251 , \48252 , \48253 , \48254 ,
         \48255 , \48256 , \48257 , \48258 , \48259 , \48260 , \48261 , \48262 , \48263 , \48264 ,
         \48265 , \48266 , \48267 , \48268 , \48269 , \48270 , \48271 , \48272 , \48273 , \48274 ,
         \48275 , \48276 , \48277 , \48278 , \48279 , \48280 , \48281 , \48282 , \48283 , \48284 ,
         \48285 , \48286 , \48287 , \48288 , \48289 , \48290 , \48291 , \48292 , \48293 , \48294 ,
         \48295 , \48296 , \48297 , \48298 , \48299 , \48300 , \48301 , \48302 , \48303 , \48304 ,
         \48305 , \48306 , \48307 , \48308 , \48309 , \48310 , \48311 , \48312 , \48313 , \48314 ,
         \48315 , \48316 , \48317 , \48318 , \48319 , \48320 , \48321 , \48322 , \48323 , \48324 ,
         \48325 , \48326 , \48327 , \48328 , \48329 , \48330 , \48331 , \48332 , \48333 , \48334 ,
         \48335 , \48336 , \48337 , \48338 , \48339 , \48340 , \48341 , \48342 , \48343 , \48344 ,
         \48345 , \48346 , \48347 , \48348 , \48349 , \48350 , \48351 , \48352 , \48353 , \48354 ,
         \48355 , \48356 , \48357 , \48358 , \48359 , \48360 , \48361 , \48362 , \48363 , \48364 ,
         \48365 , \48366 , \48367 , \48368 , \48369 , \48370 , \48371 , \48372 , \48373 , \48374 ,
         \48375 , \48376 , \48377 , \48378 , \48379 , \48380 , \48381 , \48382 , \48383 , \48384 ,
         \48385 , \48386 , \48387 , \48388 , \48389 , \48390 , \48391 , \48392 , \48393 , \48394 ,
         \48395 , \48396 , \48397 , \48398 , \48399 , \48400 , \48401 , \48402 , \48403 , \48404 ,
         \48405 , \48406 , \48407 , \48408 , \48409 , \48410 , \48411 , \48412 , \48413 , \48414 ,
         \48415 , \48416 , \48417 , \48418 , \48419 , \48420 , \48421 , \48422 , \48423 , \48424 ,
         \48425 , \48426 , \48427 , \48428 , \48429 , \48430 , \48431 , \48432 , \48433 , \48434 ,
         \48435 , \48436 , \48437 , \48438 , \48439 , \48440 , \48441 , \48442 , \48443 , \48444 ,
         \48445 , \48446 , \48447 , \48448 , \48449 , \48450 , \48451 , \48452 , \48453 , \48454 ,
         \48455 , \48456 , \48457 , \48458 , \48459 , \48460 , \48461 , \48462 , \48463 , \48464 ,
         \48465 , \48466 , \48467 , \48468 , \48469 , \48470 , \48471 , \48472 , \48473 , \48474 ,
         \48475 , \48476 , \48477 , \48478 , \48479 , \48480 , \48481 , \48482 , \48483 , \48484 ,
         \48485 , \48486 , \48487 , \48488 , \48489 , \48490 , \48491 , \48492 , \48493 , \48494 ,
         \48495 , \48496 , \48497 , \48498 , \48499 , \48500 , \48501 , \48502 , \48503 , \48504 ,
         \48505 , \48506 , \48507 , \48508 , \48509 , \48510 , \48511 , \48512 , \48513 , \48514 ,
         \48515 , \48516 , \48517 , \48518 , \48519 , \48520 , \48521 , \48522 , \48523 , \48524 ,
         \48525 , \48526 , \48527 , \48528 , \48529 , \48530 , \48531 , \48532 , \48533 , \48534 ,
         \48535 , \48536 , \48537 , \48538 , \48539 , \48540 , \48541 , \48542 , \48543 , \48544 ,
         \48545 , \48546 , \48547 , \48548 , \48549 , \48550 , \48551 , \48552 , \48553 , \48554 ,
         \48555 , \48556 , \48557 , \48558 , \48559 , \48560 , \48561 , \48562 , \48563 , \48564 ,
         \48565 , \48566 , \48567 , \48568 , \48569 , \48570 , \48571 , \48572 , \48573 , \48574 ,
         \48575 , \48576 , \48577 , \48578 , \48579 , \48580 , \48581 , \48582 , \48583 , \48584 ,
         \48585 , \48586 , \48587 , \48588 , \48589 , \48590 , \48591 , \48592 , \48593 , \48594 ,
         \48595 , \48596 , \48597 , \48598 , \48599 , \48600 , \48601 , \48602 , \48603 , \48604 ,
         \48605 , \48606 , \48607 , \48608 , \48609 , \48610 , \48611 , \48612 , \48613 , \48614 ,
         \48615 , \48616 , \48617 , \48618 , \48619 , \48620 , \48621 , \48622 , \48623 , \48624 ,
         \48625 , \48626 , \48627 , \48628 , \48629 , \48630 , \48631 , \48632 , \48633 , \48634 ,
         \48635 , \48636 , \48637 , \48638 , \48639 , \48640 , \48641 , \48642 , \48643 , \48644 ,
         \48645 , \48646 , \48647 , \48648 , \48649 , \48650 , \48651 , \48652 , \48653 , \48654 ,
         \48655 , \48656 , \48657 , \48658 , \48659 , \48660 , \48661 , \48662 , \48663 , \48664 ,
         \48665 , \48666 , \48667 , \48668 , \48669 , \48670 , \48671 , \48672 , \48673 , \48674 ,
         \48675 , \48676 , \48677 , \48678 , \48679 , \48680 , \48681 , \48682 , \48683 , \48684 ,
         \48685 , \48686 , \48687 , \48688 , \48689 , \48690 , \48691 , \48692 , \48693 , \48694 ,
         \48695 , \48696 , \48697 , \48698 , \48699 , \48700 , \48701 , \48702 , \48703 , \48704 ,
         \48705 , \48706 , \48707 , \48708 , \48709 , \48710 , \48711 , \48712 , \48713 , \48714 ,
         \48715 , \48716 , \48717 , \48718 , \48719 , \48720 , \48721 , \48722 , \48723 , \48724 ,
         \48725 , \48726 , \48727 , \48728 , \48729 , \48730 , \48731 , \48732 , \48733 , \48734 ,
         \48735 , \48736 , \48737 , \48738 , \48739 , \48740 , \48741 , \48742 , \48743 , \48744 ,
         \48745 , \48746 , \48747 , \48748 , \48749 , \48750 , \48751 , \48752 , \48753 , \48754 ,
         \48755 , \48756 , \48757 , \48758 , \48759 , \48760 , \48761 , \48762 , \48763 , \48764 ,
         \48765 , \48766 , \48767 , \48768 , \48769 , \48770 , \48771 , \48772 , \48773 , \48774 ,
         \48775 , \48776 , \48777 , \48778 , \48779 , \48780 , \48781 , \48782 , \48783 , \48784 ,
         \48785 , \48786 , \48787 , \48788 , \48789 , \48790 , \48791 , \48792 , \48793 , \48794 ,
         \48795 , \48796 , \48797 , \48798 , \48799 , \48800 , \48801 , \48802 , \48803 , \48804 ,
         \48805 , \48806 , \48807 , \48808 , \48809 , \48810 , \48811 , \48812 , \48813 , \48814 ,
         \48815 , \48816 , \48817 , \48818 , \48819 , \48820 , \48821 , \48822 , \48823 , \48824 ,
         \48825 , \48826 , \48827 , \48828 , \48829 , \48830 , \48831 , \48832 , \48833 , \48834 ,
         \48835 , \48836 , \48837 , \48838 , \48839 , \48840 , \48841 , \48842 , \48843 , \48844 ,
         \48845 , \48846 , \48847 , \48848 , \48849 , \48850 , \48851 , \48852 , \48853 , \48854 ,
         \48855 , \48856 , \48857 , \48858 , \48859 , \48860 , \48861 , \48862 , \48863 , \48864 ,
         \48865 , \48866 , \48867 , \48868 , \48869 , \48870 , \48871 , \48872 , \48873 , \48874 ,
         \48875 , \48876 , \48877 , \48878 , \48879 , \48880 , \48881 , \48882 , \48883 , \48884 ,
         \48885 , \48886 , \48887 , \48888 , \48889 , \48890 , \48891 , \48892 , \48893 , \48894 ,
         \48895 , \48896 , \48897 , \48898 , \48899 , \48900 , \48901 , \48902 , \48903 , \48904 ,
         \48905 , \48906 , \48907 , \48908 , \48909 , \48910 , \48911 , \48912 , \48913 , \48914 ,
         \48915 , \48916 , \48917 , \48918 , \48919 , \48920 , \48921 , \48922 , \48923 , \48924 ,
         \48925 , \48926 , \48927 , \48928 , \48929 , \48930 , \48931 , \48932 , \48933 , \48934 ,
         \48935 , \48936 , \48937 , \48938 , \48939 , \48940 , \48941 , \48942 , \48943 , \48944 ,
         \48945 , \48946 , \48947 , \48948 , \48949 , \48950 , \48951 , \48952 , \48953 , \48954 ,
         \48955 , \48956 , \48957 , \48958 , \48959 , \48960 , \48961 , \48962 , \48963 , \48964 ,
         \48965 , \48966 , \48967 , \48968 , \48969 , \48970 , \48971 , \48972 , \48973 , \48974 ,
         \48975 , \48976 , \48977 , \48978 , \48979 , \48980 , \48981 , \48982 , \48983 , \48984 ,
         \48985 , \48986 , \48987 , \48988 , \48989 , \48990 , \48991 , \48992 , \48993 , \48994 ,
         \48995 , \48996 , \48997 , \48998 , \48999 , \49000 , \49001 , \49002 , \49003 , \49004 ,
         \49005 , \49006 , \49007 , \49008 , \49009 , \49010 , \49011 , \49012 , \49013 , \49014 ,
         \49015 , \49016 , \49017 , \49018 , \49019 , \49020 , \49021 , \49022 , \49023 , \49024 ,
         \49025 , \49026 , \49027 , \49028 , \49029 , \49030 , \49031 , \49032 , \49033 , \49034 ,
         \49035 , \49036 , \49037 , \49038 , \49039 , \49040 , \49041 , \49042 , \49043 , \49044 ,
         \49045 , \49046 , \49047 , \49048 , \49049 , \49050 , \49051 , \49052 , \49053 , \49054 ,
         \49055 , \49056 , \49057 , \49058 , \49059 , \49060 , \49061 , \49062 , \49063 , \49064 ,
         \49065 , \49066 , \49067 , \49068 , \49069 , \49070 , \49071 , \49072 , \49073 , \49074 ,
         \49075 , \49076 , \49077 , \49078 , \49079 , \49080 , \49081 , \49082 , \49083 , \49084 ,
         \49085 , \49086 , \49087 , \49088 , \49089 , \49090 , \49091 , \49092 , \49093 , \49094 ,
         \49095 , \49096 , \49097 , \49098 , \49099 , \49100 , \49101 , \49102 , \49103 , \49104 ,
         \49105 , \49106 , \49107 , \49108 , \49109 , \49110 , \49111 , \49112 , \49113 , \49114 ,
         \49115 , \49116 , \49117 , \49118 , \49119 , \49120 , \49121 , \49122 , \49123 , \49124 ,
         \49125 , \49126 , \49127 , \49128 , \49129 , \49130 , \49131 , \49132 , \49133 , \49134 ,
         \49135 , \49136 , \49137 , \49138 , \49139 , \49140 , \49141 , \49142 , \49143 , \49144 ,
         \49145 , \49146 , \49147 , \49148 , \49149 , \49150 , \49151 , \49152 , \49153 , \49154 ,
         \49155 , \49156 , \49157 , \49158 , \49159 , \49160 , \49161 , \49162 , \49163 , \49164 ,
         \49165 , \49166 , \49167 , \49168 , \49169 , \49170 , \49171 , \49172 , \49173 , \49174 ,
         \49175 , \49176 , \49177 , \49178 , \49179 , \49180 , \49181 , \49182 , \49183 , \49184 ,
         \49185 , \49186 , \49187 , \49188 , \49189 , \49190 , \49191 , \49192 , \49193 , \49194 ,
         \49195 , \49196 , \49197 , \49198 , \49199 , \49200 , \49201 , \49202 , \49203 , \49204 ,
         \49205 , \49206 , \49207 , \49208 , \49209 , \49210 , \49211 , \49212 , \49213 , \49214 ,
         \49215 , \49216 , \49217 , \49218 , \49219 , \49220 , \49221 , \49222 , \49223 , \49224 ,
         \49225 , \49226 , \49227 , \49228 , \49229 , \49230 , \49231 , \49232 , \49233 , \49234 ,
         \49235 , \49236 , \49237 , \49238 , \49239 , \49240 , \49241 , \49242 , \49243 , \49244 ,
         \49245 , \49246 , \49247 , \49248 , \49249 , \49250 , \49251 , \49252 , \49253 , \49254 ,
         \49255 , \49256 , \49257 , \49258 , \49259 , \49260 , \49261 , \49262 , \49263 , \49264 ,
         \49265 , \49266 , \49267 , \49268 , \49269 , \49270 , \49271 , \49272 , \49273 , \49274 ,
         \49275 , \49276 , \49277 , \49278 , \49279 , \49280 , \49281 , \49282 , \49283 , \49284 ,
         \49285 , \49286 , \49287 , \49288 , \49289 , \49290 , \49291 , \49292 , \49293 , \49294 ,
         \49295 , \49296 , \49297 , \49298 , \49299 , \49300 , \49301 , \49302 , \49303 , \49304 ,
         \49305 , \49306 , \49307 , \49308 , \49309 , \49310 , \49311 , \49312 , \49313 , \49314 ,
         \49315 , \49316 , \49317 , \49318 , \49319 , \49320 , \49321 , \49322 , \49323 , \49324 ,
         \49325 , \49326 , \49327 , \49328 , \49329 , \49330 , \49331 , \49332 , \49333 , \49334 ,
         \49335 , \49336 , \49337 , \49338 , \49339 , \49340 , \49341 , \49342 , \49343 , \49344 ,
         \49345 , \49346 , \49347 , \49348 , \49349 , \49350 , \49351 , \49352 , \49353 , \49354 ,
         \49355 , \49356 , \49357 , \49358 , \49359 , \49360 , \49361 , \49362 , \49363 , \49364 ,
         \49365 , \49366 , \49367 , \49368 , \49369 , \49370 , \49371 , \49372 , \49373 , \49374 ,
         \49375 , \49376 , \49377 , \49378 , \49379 , \49380 , \49381 , \49382 , \49383 , \49384 ,
         \49385 , \49386 , \49387 , \49388 , \49389 , \49390 , \49391 , \49392 , \49393 , \49394 ,
         \49395 , \49396 , \49397 , \49398 , \49399 , \49400 , \49401 , \49402 , \49403 , \49404 ,
         \49405 , \49406 , \49407 , \49408 , \49409 , \49410 , \49411 , \49412 , \49413 , \49414 ,
         \49415 , \49416 , \49417 , \49418 , \49419 , \49420 , \49421 , \49422 , \49423 , \49424 ,
         \49425 , \49426 , \49427 , \49428 , \49429 , \49430 , \49431 , \49432 , \49433 , \49434 ,
         \49435 , \49436 , \49437 , \49438 , \49439 , \49440 , \49441 , \49442 , \49443 , \49444 ,
         \49445 , \49446 , \49447 , \49448 , \49449 , \49450 , \49451 , \49452 , \49453 , \49454 ,
         \49455 , \49456 , \49457 , \49458 , \49459 , \49460 , \49461 , \49462 , \49463 , \49464 ,
         \49465 , \49466 , \49467 , \49468 , \49469 , \49470 , \49471 , \49472 , \49473 , \49474 ,
         \49475 , \49476 , \49477 , \49478 , \49479 , \49480 , \49481 , \49482 , \49483 , \49484 ,
         \49485 , \49486 , \49487 , \49488 , \49489 , \49490 , \49491 , \49492 , \49493 , \49494 ,
         \49495 , \49496 , \49497 , \49498 , \49499 , \49500 , \49501 , \49502 , \49503 , \49504 ,
         \49505 , \49506 , \49507 , \49508 , \49509 , \49510 , \49511 , \49512 , \49513 , \49514 ,
         \49515 , \49516 , \49517 , \49518 , \49519 , \49520 , \49521 , \49522 , \49523 , \49524 ,
         \49525 , \49526 , \49527 , \49528 , \49529 , \49530 , \49531 , \49532 , \49533 , \49534 ,
         \49535 , \49536 , \49537 , \49538 , \49539 , \49540 , \49541 , \49542 , \49543 , \49544 ,
         \49545 , \49546 , \49547 , \49548 , \49549 , \49550 , \49551 , \49552 , \49553 , \49554 ,
         \49555 , \49556 , \49557 , \49558 , \49559 , \49560 , \49561 , \49562 , \49563 , \49564 ,
         \49565 , \49566 , \49567 , \49568 , \49569 , \49570 , \49571 , \49572 , \49573 , \49574 ,
         \49575 , \49576 , \49577 , \49578 , \49579 , \49580 , \49581 , \49582 , \49583 , \49584 ,
         \49585 , \49586 , \49587 , \49588 , \49589 , \49590 , \49591 , \49592 , \49593 , \49594 ,
         \49595 , \49596 , \49597 , \49598 , \49599 , \49600 , \49601 , \49602 , \49603 , \49604 ,
         \49605 , \49606 , \49607 , \49608 , \49609 , \49610 , \49611 , \49612 , \49613 , \49614 ,
         \49615 , \49616 , \49617 , \49618 , \49619 , \49620 , \49621 , \49622 , \49623 , \49624 ,
         \49625 , \49626 , \49627 , \49628 , \49629 , \49630 , \49631 , \49632 , \49633 , \49634 ,
         \49635 , \49636 , \49637 , \49638 , \49639 , \49640 , \49641 , \49642 , \49643 , \49644 ,
         \49645 , \49646 , \49647 , \49648 , \49649 , \49650 , \49651 , \49652 , \49653 , \49654 ,
         \49655 , \49656 , \49657 , \49658 , \49659 , \49660 , \49661 , \49662 , \49663 , \49664 ,
         \49665 , \49666 , \49667 , \49668 , \49669 , \49670 , \49671 , \49672 , \49673 , \49674 ,
         \49675 , \49676 , \49677 , \49678 , \49679 , \49680 , \49681 , \49682 , \49683 , \49684 ,
         \49685 , \49686 , \49687 , \49688 , \49689 , \49690 , \49691 , \49692 , \49693 , \49694 ,
         \49695 , \49696 , \49697 , \49698 , \49699 , \49700 , \49701 , \49702 , \49703 , \49704 ,
         \49705 , \49706 , \49707 , \49708 , \49709 , \49710 , \49711 , \49712 , \49713 , \49714 ,
         \49715 , \49716 , \49717 , \49718 , \49719 , \49720 , \49721 , \49722 , \49723 , \49724 ,
         \49725 , \49726 , \49727 , \49728 , \49729 , \49730 , \49731 , \49732 , \49733 , \49734 ,
         \49735 , \49736 , \49737 , \49738 , \49739 , \49740 , \49741 , \49742 , \49743 , \49744 ,
         \49745 , \49746 , \49747 , \49748 , \49749 , \49750 , \49751 , \49752 , \49753 , \49754 ,
         \49755 , \49756 , \49757 , \49758 , \49759 , \49760 , \49761 , \49762 , \49763 , \49764 ,
         \49765 , \49766 , \49767 , \49768 , \49769 , \49770 , \49771 , \49772 , \49773 , \49774 ,
         \49775 , \49776 , \49777 , \49778 , \49779 , \49780 , \49781 , \49782 , \49783 , \49784 ,
         \49785 , \49786 , \49787 , \49788 , \49789 , \49790 , \49791 , \49792 , \49793 , \49794 ,
         \49795 , \49796 , \49797 , \49798 , \49799 , \49800 , \49801 , \49802 , \49803 , \49804 ,
         \49805 , \49806 , \49807 , \49808 , \49809 , \49810 , \49811 , \49812 , \49813 , \49814 ,
         \49815 , \49816 , \49817 , \49818 , \49819 , \49820 , \49821 , \49822 , \49823 , \49824 ,
         \49825 , \49826 , \49827 , \49828 , \49829 , \49830 , \49831 , \49832 , \49833 , \49834 ,
         \49835 , \49836 , \49837 , \49838 , \49839 , \49840 , \49841 , \49842 , \49843 , \49844 ,
         \49845 , \49846 , \49847 , \49848 , \49849 , \49850 , \49851 , \49852 , \49853 , \49854 ,
         \49855 , \49856 , \49857 , \49858 , \49859 , \49860 , \49861 , \49862 , \49863 , \49864 ,
         \49865 , \49866 , \49867 , \49868 , \49869 , \49870 , \49871 , \49872 , \49873 , \49874 ,
         \49875 , \49876 , \49877 , \49878 , \49879 , \49880 , \49881 , \49882 , \49883 , \49884 ,
         \49885 , \49886 , \49887 , \49888 , \49889 , \49890 , \49891 , \49892 , \49893 , \49894 ,
         \49895 , \49896 , \49897 , \49898 , \49899 , \49900 , \49901 , \49902 , \49903 , \49904 ,
         \49905 , \49906 , \49907 , \49908 , \49909 , \49910 , \49911 , \49912 , \49913 , \49914 ,
         \49915 , \49916 , \49917 , \49918 , \49919 , \49920 , \49921 , \49922 , \49923 , \49924 ,
         \49925 , \49926 , \49927 , \49928 , \49929 , \49930 , \49931 , \49932 , \49933 , \49934 ,
         \49935 , \49936 , \49937 , \49938 , \49939 , \49940 , \49941 , \49942 , \49943 , \49944 ,
         \49945 , \49946 , \49947 , \49948 , \49949 , \49950 , \49951 , \49952 , \49953 , \49954 ,
         \49955 , \49956 , \49957 , \49958 , \49959 , \49960 , \49961 , \49962 , \49963 , \49964 ,
         \49965 , \49966 , \49967 , \49968 , \49969 , \49970 , \49971 , \49972 , \49973 , \49974 ,
         \49975 , \49976 , \49977 , \49978 , \49979 , \49980 , \49981 , \49982 , \49983 , \49984 ,
         \49985 , \49986 , \49987 , \49988 , \49989 , \49990 , \49991 , \49992 , \49993 , \49994 ,
         \49995 , \49996 , \49997 , \49998 , \49999 , \50000 , \50001 , \50002 , \50003 , \50004 ,
         \50005 , \50006 , \50007 , \50008 , \50009 , \50010 , \50011 , \50012 , \50013 , \50014 ,
         \50015 , \50016 , \50017 , \50018 , \50019 , \50020 , \50021 , \50022 , \50023 , \50024 ,
         \50025 , \50026 , \50027 , \50028 , \50029 , \50030 , \50031 , \50032 , \50033 , \50034 ,
         \50035 , \50036 , \50037 , \50038 , \50039 , \50040 , \50041 , \50042 , \50043 , \50044 ,
         \50045 , \50046 , \50047 , \50048 , \50049 , \50050 , \50051 , \50052 , \50053 , \50054 ,
         \50055 , \50056 , \50057 , \50058 , \50059 , \50060 , \50061 , \50062 , \50063 , \50064 ,
         \50065 , \50066 , \50067 , \50068 , \50069 , \50070 , \50071 , \50072 , \50073 , \50074 ,
         \50075 , \50076 , \50077 , \50078 , \50079 , \50080 , \50081 , \50082 , \50083 , \50084 ,
         \50085 , \50086 , \50087 , \50088 , \50089 , \50090 , \50091 , \50092 , \50093 , \50094 ,
         \50095 , \50096 , \50097 , \50098 , \50099 , \50100 , \50101 , \50102 , \50103 , \50104 ,
         \50105 , \50106 , \50107 , \50108 , \50109 , \50110 , \50111 , \50112 , \50113 , \50114 ,
         \50115 , \50116 , \50117 , \50118 , \50119 , \50120 , \50121 , \50122 , \50123 , \50124 ,
         \50125 , \50126 , \50127 , \50128 , \50129 , \50130 , \50131 , \50132 , \50133 , \50134 ,
         \50135 , \50136 , \50137 , \50138 , \50139 , \50140 , \50141 , \50142 , \50143 , \50144 ,
         \50145 , \50146 , \50147 , \50148 , \50149 , \50150 , \50151 , \50152 , \50153 , \50154 ,
         \50155 , \50156 , \50157 , \50158 , \50159 , \50160 , \50161 , \50162 , \50163 , \50164 ,
         \50165 , \50166 , \50167 , \50168 , \50169 , \50170 , \50171 , \50172 , \50173 , \50174 ,
         \50175 , \50176 , \50177 , \50178 , \50179 , \50180 , \50181 , \50182 , \50183 , \50184 ,
         \50185 , \50186 , \50187 , \50188 , \50189 , \50190 , \50191 , \50192 , \50193 , \50194 ,
         \50195 , \50196 , \50197 , \50198 , \50199 , \50200 , \50201 , \50202 , \50203 , \50204 ,
         \50205 , \50206 , \50207 , \50208 , \50209 , \50210 , \50211 , \50212 , \50213 , \50214 ,
         \50215 , \50216 , \50217 , \50218 , \50219 , \50220 , \50221 , \50222 , \50223 , \50224 ,
         \50225 , \50226 , \50227 , \50228 , \50229 , \50230 , \50231 , \50232 , \50233 , \50234 ,
         \50235 , \50236 , \50237 , \50238 , \50239 , \50240 , \50241 , \50242 , \50243 , \50244 ,
         \50245 , \50246 , \50247 , \50248 , \50249 , \50250 , \50251 , \50252 , \50253 , \50254 ,
         \50255 , \50256 , \50257 , \50258 , \50259 , \50260 , \50261 , \50262 , \50263 , \50264 ,
         \50265 , \50266 , \50267 , \50268 , \50269 , \50270 , \50271 , \50272 , \50273 , \50274 ,
         \50275 , \50276 , \50277 , \50278 , \50279 , \50280 , \50281 , \50282 , \50283 , \50284 ,
         \50285 , \50286 , \50287 , \50288 , \50289 , \50290 , \50291 , \50292 , \50293 , \50294 ,
         \50295 , \50296 , \50297 , \50298 , \50299 , \50300 , \50301 , \50302 , \50303 , \50304 ,
         \50305 , \50306 , \50307 , \50308 , \50309 , \50310 , \50311 , \50312 , \50313 , \50314 ,
         \50315 , \50316 , \50317 , \50318 , \50319 , \50320 , \50321 , \50322 , \50323 , \50324 ,
         \50325 , \50326 , \50327 , \50328 , \50329 , \50330 , \50331 , \50332 , \50333 , \50334 ,
         \50335 , \50336 , \50337 , \50338 , \50339 , \50340 , \50341 , \50342 , \50343 , \50344 ,
         \50345 , \50346 , \50347 , \50348 , \50349 , \50350 , \50351 , \50352 , \50353 , \50354 ,
         \50355 , \50356 , \50357 , \50358 , \50359 , \50360 , \50361 , \50362 , \50363 , \50364 ,
         \50365 , \50366 , \50367 , \50368 , \50369 , \50370 , \50371 , \50372 , \50373 , \50374 ,
         \50375 , \50376 , \50377 , \50378 , \50379 , \50380 , \50381 , \50382 , \50383 , \50384 ,
         \50385 , \50386 , \50387 , \50388 , \50389 , \50390 , \50391 , \50392 , \50393 , \50394 ,
         \50395 , \50396 , \50397 , \50398 , \50399 , \50400 , \50401 , \50402 , \50403 , \50404 ,
         \50405 , \50406 , \50407 , \50408 , \50409 , \50410 , \50411 , \50412 , \50413 , \50414 ,
         \50415 , \50416 , \50417 , \50418 , \50419 , \50420 , \50421 , \50422 , \50423 , \50424 ,
         \50425 , \50426 , \50427 , \50428 , \50429 , \50430 , \50431 , \50432 , \50433 , \50434 ,
         \50435 , \50436 , \50437 , \50438 , \50439 , \50440 , \50441 , \50442 , \50443 , \50444 ,
         \50445 , \50446 , \50447 , \50448 , \50449 , \50450 , \50451 , \50452 , \50453 , \50454 ,
         \50455 , \50456 , \50457 , \50458 , \50459 , \50460 , \50461 , \50462 , \50463 , \50464 ,
         \50465 , \50466 , \50467 , \50468 , \50469 , \50470 , \50471 , \50472 , \50473 , \50474 ,
         \50475 , \50476 , \50477 , \50478 , \50479 , \50480 , \50481 , \50482 , \50483 , \50484 ,
         \50485 , \50486 , \50487 , \50488 , \50489 , \50490 , \50491 , \50492 , \50493 , \50494 ,
         \50495 , \50496 , \50497 , \50498 , \50499 , \50500 , \50501 , \50502 , \50503 , \50504 ,
         \50505 , \50506 , \50507 , \50508 , \50509 , \50510 , \50511 , \50512 , \50513 , \50514 ,
         \50515 , \50516 , \50517 , \50518 , \50519 , \50520 , \50521 , \50522 , \50523 , \50524 ,
         \50525 , \50526 , \50527 , \50528 , \50529 , \50530 , \50531 , \50532 , \50533 , \50534 ,
         \50535 , \50536 , \50537 , \50538 , \50539 , \50540 , \50541 , \50542 , \50543 , \50544 ,
         \50545 , \50546 , \50547 , \50548 , \50549 , \50550 , \50551 , \50552 , \50553 , \50554 ,
         \50555 , \50556 , \50557 , \50558 , \50559 , \50560 , \50561 , \50562 , \50563 , \50564 ,
         \50565 , \50566 , \50567 , \50568 , \50569 , \50570 , \50571 , \50572 , \50573 , \50574 ,
         \50575 , \50576 , \50577 , \50578 , \50579 , \50580 , \50581 , \50582 , \50583 , \50584 ,
         \50585 , \50586 , \50587 , \50588 , \50589 , \50590 , \50591 , \50592 , \50593 , \50594 ,
         \50595 , \50596 , \50597 , \50598 , \50599 , \50600 , \50601 , \50602 , \50603 , \50604 ,
         \50605 , \50606 , \50607 , \50608 , \50609 , \50610 , \50611 , \50612 , \50613 , \50614 ,
         \50615 , \50616 , \50617 , \50618 , \50619 , \50620 , \50621 , \50622 , \50623 , \50624 ,
         \50625 , \50626 , \50627 , \50628 , \50629 , \50630 , \50631 , \50632 , \50633 , \50634 ,
         \50635 , \50636 , \50637 , \50638 , \50639 , \50640 , \50641 , \50642 , \50643 , \50644 ,
         \50645 , \50646 , \50647 , \50648 , \50649 , \50650 , \50651 , \50652 , \50653 , \50654 ,
         \50655 , \50656 , \50657 , \50658 , \50659 , \50660 , \50661 , \50662 , \50663 , \50664 ,
         \50665 , \50666 , \50667 , \50668 , \50669 , \50670 , \50671 , \50672 , \50673 , \50674 ,
         \50675 , \50676 , \50677 , \50678 , \50679 , \50680 , \50681 , \50682 , \50683 , \50684 ,
         \50685 , \50686 , \50687 , \50688 , \50689 , \50690 , \50691 , \50692 , \50693 , \50694 ,
         \50695 , \50696 , \50697 , \50698 , \50699 , \50700 , \50701 , \50702 , \50703 , \50704 ,
         \50705 , \50706 , \50707 , \50708 , \50709 , \50710 , \50711 , \50712 , \50713 , \50714 ,
         \50715 , \50716 , \50717 , \50718 , \50719 , \50720 , \50721 , \50722 , \50723 , \50724 ,
         \50725 , \50726 , \50727 , \50728 , \50729 , \50730 , \50731 , \50732 , \50733 , \50734 ,
         \50735 , \50736 , \50737 , \50738 , \50739 , \50740 , \50741 , \50742 , \50743 , \50744 ,
         \50745 , \50746 , \50747 , \50748 , \50749 , \50750 , \50751 , \50752 , \50753 , \50754 ,
         \50755 , \50756 , \50757 , \50758 , \50759 , \50760 , \50761 , \50762 , \50763 , \50764 ,
         \50765 , \50766 , \50767 , \50768 , \50769 , \50770 , \50771 , \50772 , \50773 , \50774 ,
         \50775 , \50776 , \50777 , \50778 , \50779 , \50780 , \50781 , \50782 , \50783 , \50784 ,
         \50785 , \50786 , \50787 , \50788 , \50789 , \50790 , \50791 , \50792 , \50793 , \50794 ,
         \50795 , \50796 , \50797 , \50798 , \50799 , \50800 , \50801 , \50802 , \50803 , \50804 ,
         \50805 , \50806 , \50807 , \50808 , \50809 , \50810 , \50811 , \50812 , \50813 , \50814 ,
         \50815 , \50816 , \50817 , \50818 , \50819 , \50820 , \50821 , \50822 , \50823 , \50824 ,
         \50825 , \50826 , \50827 , \50828 , \50829 , \50830 , \50831 , \50832 , \50833 , \50834 ,
         \50835 , \50836 , \50837 , \50838 , \50839 , \50840 , \50841 , \50842 , \50843 , \50844 ,
         \50845 , \50846 , \50847 , \50848 , \50849 , \50850 , \50851 , \50852 , \50853 , \50854 ,
         \50855 , \50856 , \50857 , \50858 , \50859 , \50860 , \50861 , \50862 , \50863 , \50864 ,
         \50865 , \50866 , \50867 , \50868 , \50869 , \50870 , \50871 , \50872 , \50873 , \50874 ,
         \50875 , \50876 , \50877 , \50878 , \50879 , \50880 , \50881 , \50882 , \50883 , \50884 ,
         \50885 , \50886 , \50887 , \50888 , \50889 , \50890 , \50891 , \50892 , \50893 , \50894 ,
         \50895 , \50896 , \50897 , \50898 , \50899 , \50900 , \50901 , \50902 , \50903 , \50904 ,
         \50905 , \50906 , \50907 , \50908 , \50909 , \50910 , \50911 , \50912 , \50913 , \50914 ,
         \50915 , \50916 , \50917 , \50918 , \50919 , \50920 , \50921 , \50922 , \50923 , \50924 ,
         \50925 , \50926 , \50927 , \50928 , \50929 , \50930 , \50931 , \50932 , \50933 , \50934 ,
         \50935 , \50936 , \50937 , \50938 , \50939 , \50940 , \50941 , \50942 , \50943 , \50944 ,
         \50945 , \50946 , \50947 , \50948 , \50949 , \50950 , \50951 , \50952 , \50953 , \50954 ,
         \50955 , \50956 , \50957 , \50958 , \50959 , \50960 , \50961 , \50962 , \50963 , \50964 ,
         \50965 , \50966 , \50967 , \50968 , \50969 , \50970 , \50971 , \50972 , \50973 , \50974 ,
         \50975 , \50976 , \50977 , \50978 , \50979 , \50980 , \50981 , \50982 , \50983 , \50984 ,
         \50985 , \50986 , \50987 , \50988 , \50989 , \50990 , \50991 , \50992 , \50993 , \50994 ,
         \50995 , \50996 , \50997 , \50998 , \50999 , \51000 , \51001 , \51002 , \51003 , \51004 ,
         \51005 , \51006 , \51007 , \51008 , \51009 , \51010 , \51011 , \51012 , \51013 , \51014 ,
         \51015 , \51016 , \51017 , \51018 , \51019 , \51020 , \51021 , \51022 , \51023 , \51024 ,
         \51025 , \51026 , \51027 , \51028 , \51029 , \51030 , \51031 , \51032 , \51033 , \51034 ,
         \51035 , \51036 , \51037 , \51038 , \51039 , \51040 , \51041 , \51042 , \51043 , \51044 ,
         \51045 , \51046 , \51047 , \51048 , \51049 , \51050 , \51051 , \51052 , \51053 , \51054 ,
         \51055 , \51056 , \51057 , \51058 , \51059 , \51060 , \51061 , \51062 , \51063 , \51064 ,
         \51065 , \51066 , \51067 , \51068 , \51069 , \51070 , \51071 , \51072 , \51073 , \51074 ,
         \51075 , \51076 , \51077 , \51078 , \51079 , \51080 , \51081 , \51082 , \51083 , \51084 ,
         \51085 , \51086 , \51087 , \51088 , \51089 , \51090 , \51091 , \51092 , \51093 , \51094 ,
         \51095 , \51096 , \51097 , \51098 , \51099 , \51100 , \51101 , \51102 , \51103 , \51104 ,
         \51105 , \51106 , \51107 , \51108 , \51109 , \51110 , \51111 , \51112 , \51113 , \51114 ,
         \51115 , \51116 , \51117 , \51118 , \51119 , \51120 , \51121 , \51122 , \51123 , \51124 ,
         \51125 , \51126 , \51127 , \51128 , \51129 , \51130 , \51131 , \51132 , \51133 , \51134 ,
         \51135 , \51136 , \51137 , \51138 , \51139 , \51140 , \51141 , \51142 , \51143 , \51144 ,
         \51145 , \51146 , \51147 , \51148 , \51149 , \51150 , \51151 , \51152 , \51153 , \51154 ,
         \51155 , \51156 , \51157 , \51158 , \51159 , \51160 , \51161 , \51162 , \51163 , \51164 ,
         \51165 , \51166 , \51167 , \51168 , \51169 , \51170 , \51171 , \51172 , \51173 , \51174 ,
         \51175 , \51176 , \51177 , \51178 , \51179 , \51180 , \51181 , \51182 , \51183 , \51184 ,
         \51185 , \51186 , \51187 , \51188 , \51189 , \51190 , \51191 , \51192 , \51193 , \51194 ,
         \51195 , \51196 , \51197 , \51198 , \51199 , \51200 , \51201 , \51202 , \51203 , \51204 ,
         \51205 , \51206 , \51207 , \51208 , \51209 , \51210 , \51211 , \51212 , \51213 , \51214 ,
         \51215 , \51216 , \51217 , \51218 , \51219 , \51220 , \51221 , \51222 , \51223 , \51224 ,
         \51225 , \51226 , \51227 , \51228 , \51229 , \51230 , \51231 , \51232 , \51233 , \51234 ,
         \51235 , \51236 , \51237 , \51238 , \51239 , \51240 , \51241 , \51242 , \51243 , \51244 ,
         \51245 , \51246 , \51247 , \51248 , \51249 , \51250 , \51251 , \51252 , \51253 , \51254 ,
         \51255 , \51256 , \51257 , \51258 , \51259 , \51260 , \51261 , \51262 , \51263 , \51264 ,
         \51265 , \51266 , \51267 , \51268 , \51269 , \51270 , \51271 , \51272 , \51273 , \51274 ,
         \51275 , \51276 , \51277 , \51278 , \51279 , \51280 , \51281 , \51282 , \51283 , \51284 ,
         \51285 , \51286 , \51287 , \51288 , \51289 , \51290 , \51291 , \51292 , \51293 , \51294 ,
         \51295 , \51296 , \51297 , \51298 , \51299 , \51300 , \51301 , \51302 , \51303 , \51304 ,
         \51305 , \51306 , \51307 , \51308 , \51309 , \51310 , \51311 , \51312 , \51313 , \51314 ,
         \51315 , \51316 , \51317 , \51318 , \51319 , \51320 , \51321 , \51322 , \51323 , \51324 ,
         \51325 , \51326 , \51327 , \51328 , \51329 , \51330 , \51331 , \51332 , \51333 , \51334 ,
         \51335 , \51336 , \51337 , \51338 , \51339 , \51340 , \51341 , \51342 , \51343 , \51344 ,
         \51345 , \51346 , \51347 , \51348 , \51349 , \51350 , \51351 , \51352 , \51353 , \51354 ,
         \51355 , \51356 , \51357 , \51358 , \51359 , \51360 , \51361 , \51362 , \51363 , \51364 ,
         \51365 , \51366 , \51367 , \51368 , \51369 , \51370 , \51371 , \51372 , \51373 , \51374 ,
         \51375 , \51376 , \51377 , \51378 , \51379 , \51380 , \51381 , \51382 , \51383 , \51384 ,
         \51385 , \51386 , \51387 , \51388 , \51389 , \51390 , \51391 , \51392 , \51393 , \51394 ,
         \51395 , \51396 , \51397 , \51398 , \51399 , \51400 , \51401 , \51402 , \51403 , \51404 ,
         \51405 , \51406 , \51407 , \51408 , \51409 , \51410 , \51411 , \51412 , \51413 , \51414 ,
         \51415 , \51416 , \51417 , \51418 , \51419 , \51420 , \51421 , \51422 , \51423 , \51424 ,
         \51425 , \51426 , \51427 , \51428 , \51429 , \51430 , \51431 , \51432 , \51433 , \51434 ,
         \51435 , \51436 , \51437 , \51438 , \51439 , \51440 , \51441 , \51442 , \51443 , \51444 ,
         \51445 , \51446 , \51447 , \51448 , \51449 , \51450 , \51451 , \51452 , \51453 , \51454 ,
         \51455 , \51456 , \51457 , \51458 , \51459 , \51460 , \51461 , \51462 , \51463 , \51464 ,
         \51465 , \51466 , \51467 , \51468 , \51469 , \51470 , \51471 , \51472 , \51473 , \51474 ,
         \51475 , \51476 , \51477 , \51478 , \51479 , \51480 , \51481 , \51482 , \51483 , \51484 ,
         \51485 , \51486 , \51487 , \51488 , \51489 , \51490 , \51491 , \51492 , \51493 , \51494 ,
         \51495 , \51496 , \51497 , \51498 , \51499 , \51500 , \51501 , \51502 , \51503 , \51504 ,
         \51505 , \51506 , \51507 , \51508 , \51509 , \51510 , \51511 , \51512 , \51513 , \51514 ,
         \51515 , \51516 , \51517 , \51518 , \51519 , \51520 , \51521 , \51522 , \51523 , \51524 ,
         \51525 , \51526 , \51527 , \51528 , \51529 , \51530 , \51531 , \51532 , \51533 , \51534 ,
         \51535 , \51536 , \51537 , \51538 , \51539 , \51540 , \51541 , \51542 , \51543 , \51544 ,
         \51545 , \51546 , \51547 , \51548 , \51549 , \51550 , \51551 , \51552 , \51553 , \51554 ,
         \51555 , \51556 , \51557 , \51558 , \51559 , \51560 , \51561 , \51562 , \51563 , \51564 ,
         \51565 , \51566 , \51567 , \51568 , \51569 , \51570 , \51571 , \51572 , \51573 , \51574 ,
         \51575 , \51576 , \51577 , \51578 , \51579 , \51580 , \51581 , \51582 , \51583 , \51584 ,
         \51585 , \51586 , \51587 , \51588 , \51589 , \51590 , \51591 , \51592 , \51593 , \51594 ,
         \51595 , \51596 , \51597 , \51598 , \51599 , \51600 , \51601 , \51602 , \51603 , \51604 ,
         \51605 , \51606 , \51607 , \51608 , \51609 , \51610 , \51611 , \51612 , \51613 , \51614 ,
         \51615 , \51616 , \51617 , \51618 , \51619 , \51620 , \51621 , \51622 , \51623 , \51624 ,
         \51625 , \51626 , \51627 , \51628 , \51629 , \51630 , \51631 , \51632 , \51633 , \51634 ,
         \51635 , \51636 , \51637 , \51638 , \51639 , \51640 , \51641 , \51642 , \51643 , \51644 ,
         \51645 , \51646 , \51647 , \51648 , \51649 , \51650 , \51651 , \51652 , \51653 , \51654 ,
         \51655 , \51656 , \51657 , \51658 , \51659 , \51660 , \51661 , \51662 , \51663 , \51664 ,
         \51665 , \51666 , \51667 , \51668 , \51669 , \51670 , \51671 , \51672 , \51673 , \51674 ,
         \51675 , \51676 , \51677 , \51678 , \51679 , \51680 , \51681 , \51682 , \51683 , \51684 ,
         \51685 , \51686 , \51687 , \51688 , \51689 , \51690 , \51691 , \51692 , \51693 , \51694 ,
         \51695 , \51696 , \51697 , \51698 , \51699 , \51700 , \51701 , \51702 , \51703 , \51704 ,
         \51705 , \51706 , \51707 , \51708 , \51709 , \51710 , \51711 , \51712 , \51713 , \51714 ,
         \51715 , \51716 , \51717 , \51718 , \51719 , \51720 , \51721 , \51722 , \51723 , \51724 ,
         \51725 , \51726 , \51727 , \51728 , \51729 , \51730 , \51731 , \51732 , \51733 , \51734 ,
         \51735 , \51736 , \51737 , \51738 , \51739 , \51740 , \51741 , \51742 , \51743 , \51744 ,
         \51745 , \51746 , \51747 , \51748 , \51749 , \51750 , \51751 , \51752 , \51753 , \51754 ,
         \51755 , \51756 , \51757 , \51758 , \51759 , \51760 , \51761 , \51762 , \51763 , \51764 ,
         \51765 , \51766 , \51767 , \51768 , \51769 , \51770 , \51771 , \51772 , \51773 , \51774 ,
         \51775 , \51776 , \51777 , \51778 , \51779 , \51780 , \51781 , \51782 , \51783 , \51784 ,
         \51785 , \51786 , \51787 , \51788 , \51789 , \51790 , \51791 , \51792 , \51793 , \51794 ,
         \51795 , \51796 , \51797 , \51798 , \51799 , \51800 , \51801 , \51802 , \51803 , \51804 ,
         \51805 , \51806 , \51807 , \51808 , \51809 , \51810 , \51811 , \51812 , \51813 , \51814 ,
         \51815 , \51816 , \51817 , \51818 , \51819 , \51820 , \51821 , \51822 , \51823 , \51824 ,
         \51825 , \51826 , \51827 , \51828 , \51829 , \51830 , \51831 , \51832 , \51833 , \51834 ,
         \51835 , \51836 , \51837 , \51838 , \51839 , \51840 , \51841 , \51842 , \51843 , \51844 ,
         \51845 , \51846 , \51847 , \51848 , \51849 , \51850 , \51851 , \51852 , \51853 , \51854 ,
         \51855 , \51856 , \51857 , \51858 , \51859 , \51860 , \51861 , \51862 , \51863 , \51864 ,
         \51865 , \51866 , \51867 , \51868 , \51869 , \51870 , \51871 , \51872 , \51873 , \51874 ,
         \51875 , \51876 , \51877 , \51878 , \51879 , \51880 , \51881 , \51882 , \51883 , \51884 ,
         \51885 , \51886 , \51887 , \51888 , \51889 , \51890 , \51891 , \51892 , \51893 , \51894 ,
         \51895 , \51896 , \51897 , \51898 , \51899 , \51900 , \51901 , \51902 , \51903 , \51904 ,
         \51905 , \51906 , \51907 , \51908 , \51909 , \51910 , \51911 , \51912 , \51913 , \51914 ,
         \51915 , \51916 , \51917 , \51918 , \51919 , \51920 , \51921 , \51922 , \51923 , \51924 ,
         \51925 , \51926 , \51927 , \51928 , \51929 , \51930 , \51931 , \51932 , \51933 , \51934 ,
         \51935 , \51936 , \51937 , \51938 , \51939 , \51940 , \51941 , \51942 , \51943 , \51944 ,
         \51945 , \51946 , \51947 , \51948 , \51949 , \51950 , \51951 , \51952 , \51953 , \51954 ,
         \51955 , \51956 , \51957 , \51958 , \51959 , \51960 , \51961 , \51962 , \51963 , \51964 ,
         \51965 , \51966 , \51967 , \51968 , \51969 , \51970 , \51971 , \51972 , \51973 , \51974 ,
         \51975 , \51976 , \51977 , \51978 , \51979 , \51980 , \51981 , \51982 , \51983 , \51984 ,
         \51985 , \51986 , \51987 , \51988 , \51989 , \51990 , \51991 , \51992 , \51993 , \51994 ,
         \51995 , \51996 , \51997 , \51998 , \51999 , \52000 , \52001 , \52002 , \52003 , \52004 ,
         \52005 , \52006 , \52007 , \52008 , \52009 , \52010 , \52011 , \52012 , \52013 , \52014 ,
         \52015 , \52016 , \52017 , \52018 , \52019 , \52020 , \52021 , \52022 , \52023 , \52024 ,
         \52025 , \52026 , \52027 , \52028 , \52029 , \52030 , \52031 , \52032 , \52033 , \52034 ,
         \52035 , \52036 , \52037 , \52038 , \52039 , \52040 , \52041 , \52042 , \52043 , \52044 ,
         \52045 , \52046 , \52047 , \52048 , \52049 , \52050 , \52051 , \52052 , \52053 , \52054 ,
         \52055 , \52056 , \52057 , \52058 , \52059 , \52060 , \52061 , \52062 , \52063 , \52064 ,
         \52065 , \52066 , \52067 , \52068 , \52069 , \52070 , \52071 , \52072 , \52073 , \52074 ,
         \52075 , \52076 , \52077 , \52078 , \52079 , \52080 , \52081 , \52082 , \52083 , \52084 ,
         \52085 , \52086 , \52087 , \52088 , \52089 , \52090 , \52091 , \52092 , \52093 , \52094 ,
         \52095 , \52096 , \52097 , \52098 , \52099 , \52100 , \52101 , \52102 , \52103 , \52104 ,
         \52105 , \52106 , \52107 , \52108 , \52109 , \52110 , \52111 , \52112 , \52113 , \52114 ,
         \52115 , \52116 , \52117 , \52118 , \52119 , \52120 , \52121 , \52122 , \52123 , \52124 ,
         \52125 , \52126 , \52127 , \52128 , \52129 , \52130 , \52131 , \52132 , \52133 , \52134 ,
         \52135 , \52136 , \52137 , \52138 , \52139 , \52140 , \52141 , \52142 , \52143 , \52144 ,
         \52145 , \52146 , \52147 , \52148 , \52149 , \52150 , \52151 , \52152 , \52153 , \52154 ,
         \52155 , \52156 , \52157 , \52158 , \52159 , \52160 , \52161 , \52162 , \52163 , \52164 ,
         \52165 , \52166 , \52167 , \52168 , \52169 , \52170 , \52171 , \52172 , \52173 , \52174 ,
         \52175 , \52176 , \52177 , \52178 , \52179 , \52180 , \52181 , \52182 , \52183 , \52184 ,
         \52185 , \52186 , \52187 , \52188 , \52189 , \52190 , \52191 , \52192 , \52193 , \52194 ,
         \52195 , \52196 , \52197 , \52198 , \52199 , \52200 , \52201 , \52202 , \52203 , \52204 ,
         \52205 , \52206 , \52207 , \52208 , \52209 , \52210 , \52211 , \52212 , \52213 , \52214 ,
         \52215 , \52216 , \52217 , \52218 , \52219 , \52220 , \52221 , \52222 , \52223 , \52224 ,
         \52225 , \52226 , \52227 , \52228 , \52229 , \52230 , \52231 , \52232 , \52233 , \52234 ,
         \52235 , \52236 , \52237 , \52238 , \52239 , \52240 , \52241 , \52242 , \52243 , \52244 ,
         \52245 , \52246 , \52247 , \52248 , \52249 , \52250 , \52251 , \52252 , \52253 , \52254 ,
         \52255 , \52256 , \52257 , \52258 , \52259 , \52260 , \52261 , \52262 , \52263 , \52264 ,
         \52265 , \52266 , \52267 , \52268 , \52269 , \52270 , \52271 , \52272 , \52273 , \52274 ,
         \52275 , \52276 , \52277 , \52278 , \52279 , \52280 , \52281 , \52282 , \52283 , \52284 ,
         \52285 , \52286 , \52287 , \52288 , \52289 , \52290 , \52291 , \52292 , \52293 , \52294 ,
         \52295 , \52296 , \52297 , \52298 , \52299 , \52300 , \52301 , \52302 , \52303 , \52304 ,
         \52305 , \52306 , \52307 , \52308 , \52309 , \52310 , \52311 , \52312 , \52313 , \52314 ,
         \52315 , \52316 , \52317 , \52318 , \52319 , \52320 , \52321 , \52322 , \52323 , \52324 ,
         \52325 , \52326 , \52327 , \52328 , \52329 , \52330 , \52331 , \52332 , \52333 , \52334 ,
         \52335 , \52336 , \52337 , \52338 , \52339 , \52340 , \52341 , \52342 , \52343 , \52344 ,
         \52345 , \52346 , \52347 , \52348 , \52349 , \52350 , \52351 , \52352 , \52353 , \52354 ,
         \52355 , \52356 , \52357 , \52358 , \52359 , \52360 , \52361 , \52362 , \52363 , \52364 ,
         \52365 , \52366 , \52367 , \52368 , \52369 , \52370 , \52371 , \52372 , \52373 , \52374 ,
         \52375 , \52376 , \52377 , \52378 , \52379 , \52380 , \52381 , \52382 , \52383 , \52384 ,
         \52385 , \52386 , \52387 , \52388 , \52389 , \52390 , \52391 , \52392 , \52393 , \52394 ,
         \52395 , \52396 , \52397 , \52398 , \52399 , \52400 , \52401 , \52402 , \52403 , \52404 ,
         \52405 , \52406 , \52407 , \52408 , \52409 , \52410 , \52411 , \52412 , \52413 , \52414 ,
         \52415 , \52416 , \52417 , \52418 , \52419 , \52420 , \52421 , \52422 , \52423 , \52424 ,
         \52425 , \52426 , \52427 , \52428 , \52429 , \52430 , \52431 , \52432 , \52433 , \52434 ,
         \52435 , \52436 , \52437 , \52438 , \52439 , \52440 , \52441 , \52442 , \52443 , \52444 ,
         \52445 , \52446 , \52447 , \52448 , \52449 , \52450 , \52451 , \52452 , \52453 , \52454 ,
         \52455 , \52456 , \52457 , \52458 , \52459 , \52460 , \52461 , \52462 , \52463 , \52464 ,
         \52465 , \52466 , \52467 , \52468 , \52469 , \52470 , \52471 , \52472 , \52473 , \52474 ,
         \52475 , \52476 , \52477 , \52478 , \52479 , \52480 , \52481 , \52482 , \52483 , \52484 ,
         \52485 , \52486 , \52487 , \52488 , \52489 , \52490 , \52491 , \52492 , \52493 , \52494 ,
         \52495 , \52496 , \52497 , \52498 , \52499 , \52500 , \52501 , \52502 , \52503 , \52504 ,
         \52505 , \52506 , \52507 , \52508 , \52509 , \52510 , \52511 , \52512 , \52513 , \52514 ,
         \52515 , \52516 , \52517 , \52518 , \52519 , \52520 , \52521 , \52522 , \52523 , \52524 ,
         \52525 , \52526 , \52527 , \52528 , \52529 , \52530 , \52531 , \52532 , \52533 , \52534 ,
         \52535 , \52536 , \52537 , \52538 , \52539 , \52540 , \52541 , \52542 , \52543 , \52544 ,
         \52545 , \52546 , \52547 , \52548 , \52549 , \52550 , \52551 , \52552 , \52553 , \52554 ,
         \52555 , \52556 , \52557 , \52558 , \52559 , \52560 , \52561 , \52562 , \52563 , \52564 ,
         \52565 , \52566 , \52567 , \52568 , \52569 , \52570 , \52571 , \52572 , \52573 , \52574 ,
         \52575 , \52576 , \52577 , \52578 , \52579 , \52580 , \52581 , \52582 , \52583 , \52584 ,
         \52585 , \52586 , \52587 , \52588 , \52589 , \52590 , \52591 , \52592 , \52593 , \52594 ,
         \52595 , \52596 , \52597 , \52598 , \52599 , \52600 , \52601 , \52602 , \52603 , \52604 ,
         \52605 , \52606 , \52607 , \52608 , \52609 , \52610 , \52611 , \52612 , \52613 , \52614 ,
         \52615 , \52616 , \52617 , \52618 , \52619 , \52620 , \52621 , \52622 , \52623 , \52624 ,
         \52625 , \52626 , \52627 , \52628 , \52629 , \52630 , \52631 , \52632 , \52633 , \52634 ,
         \52635 , \52636 , \52637 , \52638 , \52639 , \52640 , \52641 , \52642 , \52643 , \52644 ,
         \52645 , \52646 , \52647 , \52648 , \52649 , \52650 , \52651 , \52652 , \52653 , \52654 ,
         \52655 , \52656 , \52657 , \52658 , \52659 , \52660 , \52661 , \52662 , \52663 , \52664 ,
         \52665 , \52666 , \52667 , \52668 , \52669 , \52670 , \52671 , \52672 , \52673 , \52674 ,
         \52675 , \52676 , \52677 , \52678 , \52679 , \52680 , \52681 , \52682 , \52683 , \52684 ,
         \52685 , \52686 , \52687 , \52688 , \52689 , \52690 , \52691 , \52692 , \52693 , \52694 ,
         \52695 , \52696 , \52697 , \52698 , \52699 , \52700 , \52701 , \52702 , \52703 , \52704 ,
         \52705 , \52706 , \52707 , \52708 , \52709 , \52710 , \52711 , \52712 , \52713 , \52714 ,
         \52715 , \52716 , \52717 , \52718 , \52719 , \52720 , \52721 , \52722 , \52723 , \52724 ,
         \52725 , \52726 , \52727 , \52728 , \52729 , \52730 , \52731 , \52732 , \52733 , \52734 ,
         \52735 , \52736 , \52737 , \52738 , \52739 , \52740 , \52741 , \52742 , \52743 , \52744 ,
         \52745 , \52746 , \52747 , \52748 , \52749 , \52750 , \52751 , \52752 , \52753 , \52754 ,
         \52755 , \52756 , \52757 , \52758 , \52759 , \52760 , \52761 , \52762 , \52763 , \52764 ,
         \52765 , \52766 , \52767 , \52768 , \52769 , \52770 , \52771 , \52772 , \52773 , \52774 ,
         \52775 , \52776 , \52777 , \52778 , \52779 , \52780 , \52781 , \52782 , \52783 , \52784 ,
         \52785 , \52786 , \52787 , \52788 , \52789 , \52790 , \52791 , \52792 , \52793 , \52794 ,
         \52795 , \52796 , \52797 , \52798 , \52799 , \52800 , \52801 , \52802 , \52803 , \52804 ,
         \52805 , \52806 , \52807 , \52808 , \52809 , \52810 , \52811 , \52812 , \52813 , \52814 ,
         \52815 , \52816 , \52817 , \52818 , \52819 , \52820 , \52821 , \52822 , \52823 , \52824 ,
         \52825 , \52826 , \52827 , \52828 , \52829 , \52830 , \52831 , \52832 , \52833 , \52834 ,
         \52835 , \52836 , \52837 , \52838 , \52839 , \52840 , \52841 , \52842 , \52843 , \52844 ,
         \52845 , \52846 , \52847 , \52848 , \52849 , \52850 , \52851 , \52852 , \52853 , \52854 ,
         \52855 , \52856 , \52857 , \52858 , \52859 , \52860 , \52861 , \52862 , \52863 , \52864 ,
         \52865 , \52866 , \52867 , \52868 , \52869 , \52870 , \52871 , \52872 , \52873 , \52874 ,
         \52875 , \52876 , \52877 , \52878 , \52879 , \52880 , \52881 , \52882 , \52883 , \52884 ,
         \52885 , \52886 , \52887 , \52888 , \52889 , \52890 , \52891 , \52892 , \52893 , \52894 ,
         \52895 , \52896 , \52897 , \52898 , \52899 , \52900 , \52901 , \52902 , \52903 , \52904 ,
         \52905 , \52906 , \52907 , \52908 , \52909 , \52910 , \52911 , \52912 , \52913 , \52914 ,
         \52915 , \52916 , \52917 , \52918 , \52919 , \52920 , \52921 , \52922 , \52923 , \52924 ,
         \52925 , \52926 , \52927 , \52928 , \52929 , \52930 , \52931 , \52932 , \52933 , \52934 ,
         \52935 , \52936 , \52937 , \52938 , \52939 , \52940 , \52941 , \52942 , \52943 , \52944 ,
         \52945 , \52946 , \52947 , \52948 , \52949 , \52950 , \52951 , \52952 , \52953 , \52954 ,
         \52955 , \52956 , \52957 , \52958 , \52959 , \52960 , \52961 , \52962 , \52963 , \52964 ,
         \52965 , \52966 , \52967 , \52968 , \52969 , \52970 , \52971 , \52972 , \52973 , \52974 ,
         \52975 , \52976 , \52977 , \52978 , \52979 , \52980 , \52981 , \52982 , \52983 , \52984 ,
         \52985 , \52986 , \52987 , \52988 , \52989 , \52990 , \52991 , \52992 , \52993 , \52994 ,
         \52995 , \52996 , \52997 , \52998 , \52999 , \53000 , \53001 , \53002 , \53003 , \53004 ,
         \53005 , \53006 , \53007 , \53008 , \53009 , \53010 , \53011 , \53012 , \53013 , \53014 ,
         \53015 , \53016 , \53017 , \53018 , \53019 , \53020 , \53021 , \53022 , \53023 , \53024 ,
         \53025 , \53026 , \53027 , \53028 , \53029 , \53030 , \53031 , \53032 , \53033 , \53034 ,
         \53035 , \53036 , \53037 , \53038 , \53039 , \53040 , \53041 , \53042 , \53043 , \53044 ,
         \53045 , \53046 , \53047 , \53048 , \53049 , \53050 , \53051 , \53052 , \53053 , \53054 ,
         \53055 , \53056 , \53057 , \53058 , \53059 , \53060 , \53061 , \53062 , \53063 , \53064 ,
         \53065 , \53066 , \53067 , \53068 , \53069 , \53070 , \53071 , \53072 , \53073 , \53074 ,
         \53075 , \53076 , \53077 , \53078 , \53079 , \53080 , \53081 , \53082 , \53083 , \53084 ,
         \53085 , \53086 , \53087 , \53088 , \53089 , \53090 , \53091 , \53092 , \53093 , \53094 ,
         \53095 , \53096 , \53097 , \53098 , \53099 , \53100 , \53101 , \53102 , \53103 , \53104 ,
         \53105 , \53106 , \53107 , \53108 , \53109 , \53110 , \53111 , \53112 , \53113 , \53114 ,
         \53115 , \53116 , \53117 , \53118 , \53119 , \53120 , \53121 , \53122 , \53123 , \53124 ,
         \53125 , \53126 , \53127 , \53128 , \53129 , \53130 , \53131 , \53132 , \53133 , \53134 ,
         \53135 , \53136 , \53137 , \53138 , \53139 , \53140 , \53141 , \53142 , \53143 , \53144 ,
         \53145 , \53146 , \53147 , \53148 , \53149 , \53150 , \53151 , \53152 , \53153 , \53154 ,
         \53155 , \53156 , \53157 , \53158 , \53159 , \53160 , \53161 , \53162 , \53163 , \53164 ,
         \53165 , \53166 , \53167 , \53168 , \53169 , \53170 , \53171 , \53172 , \53173 , \53174 ,
         \53175 , \53176 , \53177 , \53178 , \53179 , \53180 , \53181 , \53182 , \53183 , \53184 ,
         \53185 , \53186 , \53187 , \53188 , \53189 , \53190 , \53191 , \53192 , \53193 , \53194 ,
         \53195 , \53196 , \53197 , \53198 , \53199 , \53200 , \53201 , \53202 , \53203 , \53204 ,
         \53205 , \53206 , \53207 , \53208 , \53209 , \53210 , \53211 , \53212 , \53213 , \53214 ,
         \53215 , \53216 , \53217 , \53218 , \53219 , \53220 , \53221 , \53222 , \53223 , \53224 ,
         \53225 , \53226 , \53227 , \53228 , \53229 , \53230 , \53231 , \53232 , \53233 , \53234 ,
         \53235 , \53236 , \53237 , \53238 , \53239 , \53240 , \53241 , \53242 , \53243 , \53244 ,
         \53245 , \53246 , \53247 , \53248 , \53249 , \53250 , \53251 , \53252 , \53253 , \53254 ,
         \53255 , \53256 , \53257 , \53258 , \53259 , \53260 , \53261 , \53262 , \53263 , \53264 ,
         \53265 , \53266 , \53267 , \53268 , \53269 , \53270 , \53271 , \53272 , \53273 , \53274 ,
         \53275 , \53276 , \53277 , \53278 , \53279 , \53280 , \53281 , \53282 , \53283 , \53284 ,
         \53285 , \53286 , \53287 , \53288 , \53289 , \53290 , \53291 , \53292 , \53293 , \53294 ,
         \53295 , \53296 , \53297 , \53298 , \53299 , \53300 , \53301 , \53302 , \53303 , \53304 ,
         \53305 , \53306 , \53307 , \53308 , \53309 , \53310 , \53311 , \53312 , \53313 , \53314 ,
         \53315 , \53316 , \53317 , \53318 , \53319 , \53320 , \53321 , \53322 , \53323 , \53324 ,
         \53325 , \53326 , \53327 , \53328 , \53329 , \53330 , \53331 , \53332 , \53333 , \53334 ,
         \53335 , \53336 , \53337 , \53338 , \53339 , \53340 , \53341 , \53342 , \53343 , \53344 ,
         \53345 , \53346 , \53347 , \53348 , \53349 , \53350 , \53351 , \53352 , \53353 , \53354 ,
         \53355 , \53356 , \53357 , \53358 , \53359 , \53360 , \53361 , \53362 , \53363 , \53364 ,
         \53365 , \53366 , \53367 , \53368 , \53369 , \53370 , \53371 , \53372 , \53373 , \53374 ,
         \53375 , \53376 , \53377 , \53378 , \53379 , \53380 , \53381 , \53382 , \53383 , \53384 ,
         \53385 , \53386 , \53387 , \53388 , \53389 , \53390 , \53391 , \53392 , \53393 , \53394 ,
         \53395 , \53396 , \53397 , \53398 , \53399 , \53400 , \53401 , \53402 , \53403 , \53404 ,
         \53405 , \53406 , \53407 , \53408 , \53409 , \53410 , \53411 , \53412 , \53413 , \53414 ,
         \53415 , \53416 , \53417 , \53418 , \53419 , \53420 , \53421 , \53422 , \53423 , \53424 ,
         \53425 , \53426 , \53427 , \53428 , \53429 , \53430 , \53431 , \53432 , \53433 , \53434 ,
         \53435 , \53436 , \53437 , \53438 , \53439 , \53440 , \53441 , \53442 , \53443 , \53444 ,
         \53445 , \53446 , \53447 , \53448 , \53449 , \53450 , \53451 , \53452 , \53453 , \53454 ,
         \53455 , \53456 , \53457 , \53458 , \53459 , \53460 , \53461 , \53462 , \53463 , \53464 ,
         \53465 , \53466 , \53467 , \53468 , \53469 , \53470 , \53471 , \53472 , \53473 , \53474 ,
         \53475 , \53476 , \53477 , \53478 , \53479 , \53480 , \53481 , \53482 , \53483 , \53484 ,
         \53485 , \53486 , \53487 , \53488 , \53489 , \53490 , \53491 , \53492 , \53493 , \53494 ,
         \53495 , \53496 , \53497 , \53498 , \53499 , \53500 , \53501 , \53502 , \53503 , \53504 ,
         \53505 , \53506 , \53507 , \53508 , \53509 , \53510 , \53511 , \53512 , \53513 , \53514 ,
         \53515 , \53516 , \53517 , \53518 , \53519 , \53520 , \53521 , \53522 , \53523 , \53524 ,
         \53525 , \53526 , \53527 , \53528 , \53529 , \53530 , \53531 , \53532 , \53533 , \53534 ,
         \53535 , \53536 , \53537 , \53538 , \53539 , \53540 , \53541 , \53542 , \53543 , \53544 ,
         \53545 , \53546 , \53547 , \53548 , \53549 , \53550 , \53551 , \53552 , \53553 , \53554 ,
         \53555 , \53556 , \53557 , \53558 , \53559 , \53560 , \53561 , \53562 , \53563 , \53564 ,
         \53565 , \53566 , \53567 , \53568 , \53569 , \53570 , \53571 , \53572 , \53573 , \53574 ,
         \53575 , \53576 , \53577 , \53578 , \53579 , \53580 , \53581 , \53582 , \53583 , \53584 ,
         \53585 , \53586 , \53587 , \53588 , \53589 , \53590 , \53591 , \53592 , \53593 , \53594 ,
         \53595 , \53596 , \53597 , \53598 , \53599 , \53600 , \53601 , \53602 , \53603 , \53604 ,
         \53605 , \53606 , \53607 , \53608 , \53609 , \53610 , \53611 , \53612 , \53613 , \53614 ,
         \53615 , \53616 , \53617 , \53618 , \53619 , \53620 , \53621 , \53622 , \53623 , \53624 ,
         \53625 , \53626 , \53627 , \53628 , \53629 , \53630 , \53631 , \53632 , \53633 , \53634 ,
         \53635 , \53636 , \53637 , \53638 , \53639 , \53640 , \53641 , \53642 , \53643 , \53644 ,
         \53645 , \53646 , \53647 , \53648 , \53649 , \53650 , \53651 , \53652 , \53653 , \53654 ,
         \53655 , \53656 , \53657 , \53658 , \53659 , \53660 , \53661 , \53662 , \53663 , \53664 ,
         \53665 , \53666 , \53667 , \53668 , \53669 , \53670 , \53671 , \53672 , \53673 , \53674 ,
         \53675 , \53676 , \53677 , \53678 , \53679 , \53680 , \53681 , \53682 , \53683 , \53684 ,
         \53685 , \53686 , \53687 , \53688 , \53689 , \53690 , \53691 , \53692 , \53693 , \53694 ,
         \53695 , \53696 , \53697 , \53698 , \53699 , \53700 , \53701 , \53702 , \53703 , \53704 ,
         \53705 , \53706 , \53707 , \53708 , \53709 , \53710 , \53711 , \53712 , \53713 , \53714 ,
         \53715 , \53716 , \53717 , \53718 , \53719 , \53720 , \53721 , \53722 , \53723 , \53724 ,
         \53725 , \53726 , \53727 , \53728 , \53729 , \53730 , \53731 , \53732 , \53733 , \53734 ,
         \53735 , \53736 , \53737 , \53738 , \53739 , \53740 , \53741 , \53742 , \53743 , \53744 ,
         \53745 , \53746 , \53747 , \53748 , \53749 , \53750 , \53751 , \53752 , \53753 , \53754 ,
         \53755 , \53756 , \53757 , \53758 , \53759 , \53760 , \53761 , \53762 , \53763 , \53764 ,
         \53765 , \53766 , \53767 , \53768 , \53769 , \53770 , \53771 , \53772 , \53773 , \53774 ,
         \53775 , \53776 , \53777 , \53778 , \53779 , \53780 , \53781 , \53782 , \53783 , \53784 ,
         \53785 , \53786 , \53787 , \53788 , \53789 , \53790 , \53791 , \53792 , \53793 , \53794 ,
         \53795 , \53796 , \53797 , \53798 , \53799 , \53800 , \53801 , \53802 , \53803 , \53804 ,
         \53805 , \53806 , \53807 , \53808 , \53809 , \53810 , \53811 , \53812 , \53813 , \53814 ,
         \53815 , \53816 , \53817 , \53818 , \53819 , \53820 , \53821 , \53822 , \53823 , \53824 ,
         \53825 , \53826 , \53827 , \53828 , \53829 , \53830 , \53831 , \53832 , \53833 , \53834 ,
         \53835 , \53836 , \53837 , \53838 , \53839 , \53840 , \53841 , \53842 , \53843 , \53844 ,
         \53845 , \53846 , \53847 , \53848 , \53849 , \53850 , \53851 , \53852 , \53853 , \53854 ,
         \53855 , \53856 , \53857 , \53858 , \53859 , \53860 , \53861 , \53862 , \53863 , \53864 ,
         \53865 , \53866 , \53867 , \53868 , \53869 , \53870 , \53871 , \53872 , \53873 , \53874 ,
         \53875 , \53876 , \53877 , \53878 , \53879 , \53880 , \53881 , \53882 , \53883 , \53884 ,
         \53885 , \53886 , \53887 , \53888 , \53889 , \53890 , \53891 , \53892 , \53893 , \53894 ,
         \53895 , \53896 , \53897 , \53898 , \53899 , \53900 , \53901 , \53902 , \53903 , \53904 ,
         \53905 , \53906 , \53907 , \53908 , \53909 , \53910 , \53911 , \53912 , \53913 , \53914 ,
         \53915 , \53916 , \53917 , \53918 , \53919 , \53920 , \53921 , \53922 , \53923 , \53924 ,
         \53925 , \53926 , \53927 , \53928 , \53929 , \53930 , \53931 , \53932 , \53933 , \53934 ,
         \53935 , \53936 , \53937 , \53938 , \53939 , \53940 , \53941 , \53942 , \53943 , \53944 ,
         \53945 , \53946 , \53947 , \53948 , \53949 , \53950 , \53951 , \53952 , \53953 , \53954 ,
         \53955 , \53956 , \53957 , \53958 , \53959 , \53960 , \53961 , \53962 , \53963 , \53964 ,
         \53965 , \53966 , \53967 , \53968 , \53969 , \53970 , \53971 , \53972 , \53973 , \53974 ,
         \53975 , \53976 , \53977 , \53978 , \53979 , \53980 , \53981 , \53982 , \53983 , \53984 ,
         \53985 , \53986 , \53987 , \53988 , \53989 , \53990 , \53991 , \53992 , \53993 , \53994 ,
         \53995 , \53996 , \53997 , \53998 , \53999 , \54000 , \54001 , \54002 , \54003 , \54004 ,
         \54005 , \54006 , \54007 , \54008 , \54009 , \54010 , \54011 , \54012 , \54013 , \54014 ,
         \54015 , \54016 , \54017 , \54018 , \54019 , \54020 , \54021 , \54022 , \54023 , \54024 ,
         \54025 , \54026 , \54027 , \54028 , \54029 , \54030 , \54031 , \54032 , \54033 , \54034 ,
         \54035 , \54036 , \54037 , \54038 , \54039 , \54040 , \54041 , \54042 , \54043 , \54044 ,
         \54045 , \54046 , \54047 , \54048 , \54049 , \54050 , \54051 , \54052 , \54053 , \54054 ,
         \54055 , \54056 , \54057 , \54058 , \54059 , \54060 , \54061 , \54062 , \54063 , \54064 ,
         \54065 , \54066 , \54067 , \54068 , \54069 , \54070 , \54071 , \54072 , \54073 , \54074 ,
         \54075 , \54076 , \54077 , \54078 , \54079 , \54080 , \54081 , \54082 , \54083 , \54084 ,
         \54085 , \54086 , \54087 , \54088 , \54089 , \54090 , \54091 , \54092 , \54093 , \54094 ,
         \54095 , \54096 , \54097 , \54098 , \54099 , \54100 , \54101 , \54102 , \54103 , \54104 ,
         \54105 , \54106 , \54107 , \54108 , \54109 , \54110 , \54111 , \54112 , \54113 , \54114 ,
         \54115 , \54116 , \54117 , \54118 , \54119 , \54120 , \54121 , \54122 , \54123 , \54124 ,
         \54125 , \54126 , \54127 , \54128 , \54129 , \54130 , \54131 , \54132 , \54133 , \54134 ,
         \54135 , \54136 , \54137 , \54138 , \54139 , \54140 , \54141 , \54142 , \54143 , \54144 ,
         \54145 , \54146 , \54147 , \54148 , \54149 , \54150 , \54151 , \54152 , \54153 , \54154 ,
         \54155 , \54156 , \54157 , \54158 , \54159 , \54160 , \54161 , \54162 , \54163 , \54164 ,
         \54165 , \54166 , \54167 , \54168 , \54169 , \54170 , \54171 , \54172 , \54173 , \54174 ,
         \54175 , \54176 , \54177 , \54178 , \54179 , \54180 , \54181 , \54182 , \54183 , \54184 ,
         \54185 , \54186 , \54187 , \54188 , \54189 , \54190 , \54191 , \54192 , \54193 , \54194 ,
         \54195 , \54196 , \54197 , \54198 , \54199 , \54200 , \54201 , \54202 , \54203 , \54204 ,
         \54205 , \54206 , \54207 , \54208 , \54209 , \54210 , \54211 , \54212 , \54213 , \54214 ,
         \54215 , \54216 , \54217 , \54218 , \54219 , \54220 , \54221 , \54222 , \54223 , \54224 ,
         \54225 , \54226 , \54227 , \54228 , \54229 , \54230 , \54231 , \54232 , \54233 , \54234 ,
         \54235 , \54236 , \54237 , \54238 , \54239 , \54240 , \54241 , \54242 , \54243 , \54244 ,
         \54245 , \54246 , \54247 , \54248 , \54249 , \54250 , \54251 , \54252 , \54253 , \54254 ,
         \54255 , \54256 , \54257 , \54258 , \54259 , \54260 , \54261 , \54262 , \54263 , \54264 ,
         \54265 , \54266 , \54267 , \54268 , \54269 , \54270 , \54271 , \54272 , \54273 , \54274 ,
         \54275 , \54276 , \54277 , \54278 , \54279 , \54280 , \54281 , \54282 , \54283 , \54284 ,
         \54285 , \54286 , \54287 , \54288 , \54289 , \54290 , \54291 , \54292 , \54293 , \54294 ,
         \54295 , \54296 , \54297 , \54298 , \54299 , \54300 , \54301 , \54302 , \54303 , \54304 ,
         \54305 , \54306 , \54307 , \54308 , \54309 , \54310 , \54311 , \54312 , \54313 , \54314 ,
         \54315 , \54316 , \54317 , \54318 , \54319 , \54320 , \54321 , \54322 , \54323 , \54324 ,
         \54325 , \54326 , \54327 , \54328 , \54329 , \54330 , \54331 , \54332 , \54333 , \54334 ,
         \54335 , \54336 , \54337 , \54338 , \54339 , \54340 , \54341 , \54342 , \54343 , \54344 ,
         \54345 , \54346 , \54347 , \54348 , \54349 , \54350 , \54351 , \54352 , \54353 , \54354 ,
         \54355 , \54356 , \54357 , \54358 , \54359 , \54360 , \54361 , \54362 , \54363 , \54364 ,
         \54365 , \54366 , \54367 , \54368 , \54369 , \54370 , \54371 , \54372 , \54373 , \54374 ,
         \54375 , \54376 , \54377 , \54378 , \54379 , \54380 , \54381 , \54382 , \54383 , \54384 ,
         \54385 , \54386 , \54387 , \54388 , \54389 , \54390 , \54391 , \54392 , \54393 , \54394 ,
         \54395 , \54396 , \54397 , \54398 , \54399 , \54400 , \54401 , \54402 , \54403 , \54404 ,
         \54405 , \54406 , \54407 , \54408 , \54409 , \54410 , \54411 , \54412 , \54413 , \54414 ,
         \54415 , \54416 , \54417 , \54418 , \54419 , \54420 , \54421 , \54422 , \54423 , \54424 ,
         \54425 , \54426 , \54427 , \54428 , \54429 , \54430 , \54431 , \54432 , \54433 , \54434 ,
         \54435 , \54436 , \54437 , \54438 , \54439 , \54440 , \54441 , \54442 , \54443 , \54444 ,
         \54445 , \54446 , \54447 , \54448 , \54449 , \54450 , \54451 , \54452 , \54453 , \54454 ,
         \54455 , \54456 , \54457 , \54458 , \54459 , \54460 , \54461 , \54462 , \54463 , \54464 ,
         \54465 , \54466 , \54467 , \54468 , \54469 , \54470 , \54471 , \54472 , \54473 , \54474 ,
         \54475 , \54476 , \54477 , \54478 , \54479 , \54480 , \54481 , \54482 , \54483 , \54484 ,
         \54485 , \54486 , \54487 , \54488 , \54489 , \54490 , \54491 , \54492 , \54493 , \54494 ,
         \54495 , \54496 , \54497 , \54498 , \54499 , \54500 , \54501 , \54502 , \54503 , \54504 ,
         \54505 , \54506 , \54507 , \54508 , \54509 , \54510 , \54511 , \54512 , \54513 , \54514 ,
         \54515 , \54516 , \54517 , \54518 , \54519 , \54520 , \54521 , \54522 , \54523 , \54524 ,
         \54525 , \54526 , \54527 , \54528 , \54529 , \54530 , \54531 , \54532 , \54533 , \54534 ,
         \54535 , \54536 , \54537 , \54538 , \54539 , \54540 , \54541 , \54542 , \54543 , \54544 ,
         \54545 , \54546 , \54547 , \54548 , \54549 , \54550 , \54551 , \54552 , \54553 , \54554 ,
         \54555 , \54556 , \54557 , \54558 , \54559 , \54560 , \54561 , \54562 , \54563 , \54564 ,
         \54565 , \54566 , \54567 , \54568 , \54569 , \54570 , \54571 , \54572 , \54573 , \54574 ,
         \54575 , \54576 , \54577 , \54578 , \54579 , \54580 , \54581 , \54582 , \54583 , \54584 ,
         \54585 , \54586 , \54587 , \54588 , \54589 , \54590 , \54591 , \54592 , \54593 , \54594 ,
         \54595 , \54596 , \54597 , \54598 , \54599 , \54600 , \54601 , \54602 , \54603 , \54604 ,
         \54605 , \54606 , \54607 , \54608 , \54609 , \54610 , \54611 , \54612 , \54613 , \54614 ,
         \54615 , \54616 , \54617 , \54618 , \54619 , \54620 , \54621 , \54622 , \54623 , \54624 ,
         \54625 , \54626 , \54627 , \54628 , \54629 , \54630 , \54631 , \54632 , \54633 , \54634 ,
         \54635 , \54636 , \54637 , \54638 , \54639 , \54640 , \54641 , \54642 , \54643 , \54644 ,
         \54645 , \54646 , \54647 , \54648 , \54649 , \54650 , \54651 , \54652 , \54653 , \54654 ,
         \54655 , \54656 , \54657 , \54658 , \54659 , \54660 , \54661 , \54662 , \54663 , \54664 ,
         \54665 , \54666 , \54667 , \54668 , \54669 , \54670 , \54671 , \54672 , \54673 , \54674 ,
         \54675 , \54676 , \54677 , \54678 , \54679 , \54680 , \54681 , \54682 , \54683 , \54684 ,
         \54685 , \54686 , \54687 , \54688 , \54689 , \54690 , \54691 , \54692 , \54693 , \54694 ,
         \54695 , \54696 , \54697 , \54698 , \54699 , \54700 , \54701 , \54702 , \54703 , \54704 ,
         \54705 , \54706 , \54707 , \54708 , \54709 , \54710 , \54711 , \54712 , \54713 , \54714 ,
         \54715 , \54716 , \54717 , \54718 , \54719 , \54720 , \54721 , \54722 , \54723 , \54724 ,
         \54725 , \54726 , \54727 , \54728 , \54729 , \54730 , \54731 , \54732 , \54733 , \54734 ,
         \54735 , \54736 , \54737 , \54738 , \54739 , \54740 , \54741 , \54742 , \54743 , \54744 ,
         \54745 , \54746 , \54747 , \54748 , \54749 , \54750 , \54751 , \54752 , \54753 , \54754 ,
         \54755 , \54756 , \54757 , \54758 , \54759 , \54760 , \54761 , \54762 , \54763 , \54764 ,
         \54765 , \54766 , \54767 , \54768 , \54769 , \54770 , \54771 , \54772 , \54773 , \54774 ,
         \54775 , \54776 , \54777 , \54778 , \54779 , \54780 , \54781 , \54782 , \54783 , \54784 ,
         \54785 , \54786 , \54787 , \54788 , \54789 , \54790 , \54791 , \54792 , \54793 , \54794 ,
         \54795 , \54796 , \54797 , \54798 , \54799 , \54800 , \54801 , \54802 , \54803 , \54804 ,
         \54805 , \54806 , \54807 , \54808 , \54809 , \54810 , \54811 , \54812 , \54813 , \54814 ,
         \54815 , \54816 , \54817 , \54818 , \54819 , \54820 , \54821 , \54822 , \54823 , \54824 ,
         \54825 , \54826 , \54827 , \54828 , \54829 , \54830 , \54831 , \54832 , \54833 , \54834 ,
         \54835 , \54836 , \54837 , \54838 , \54839 , \54840 , \54841 , \54842 , \54843 , \54844 ,
         \54845 , \54846 , \54847 , \54848 , \54849 , \54850 , \54851 , \54852 , \54853 , \54854 ,
         \54855 , \54856 , \54857 , \54858 , \54859 , \54860 , \54861 , \54862 , \54863 , \54864 ,
         \54865 , \54866 , \54867 , \54868 , \54869 , \54870 , \54871 , \54872 , \54873 , \54874 ,
         \54875 , \54876 , \54877 , \54878 , \54879 , \54880 , \54881 , \54882 , \54883 , \54884 ,
         \54885 , \54886 , \54887 , \54888 , \54889 , \54890 , \54891 , \54892 , \54893 , \54894 ,
         \54895 , \54896 , \54897 , \54898 , \54899 , \54900 , \54901 , \54902 , \54903 , \54904 ,
         \54905 , \54906 , \54907 , \54908 , \54909 , \54910 , \54911 , \54912 , \54913 , \54914 ,
         \54915 , \54916 , \54917 , \54918 , \54919 , \54920 , \54921 , \54922 , \54923 , \54924 ,
         \54925 , \54926 , \54927 , \54928 , \54929 , \54930 , \54931 , \54932 , \54933 , \54934 ,
         \54935 , \54936 , \54937 , \54938 , \54939 , \54940 , \54941 , \54942 , \54943 , \54944 ,
         \54945 , \54946 , \54947 , \54948 , \54949 , \54950 , \54951 , \54952 , \54953 , \54954 ,
         \54955 , \54956 , \54957 , \54958 , \54959 , \54960 , \54961 , \54962 , \54963 , \54964 ,
         \54965 , \54966 , \54967 , \54968 , \54969 , \54970 , \54971 , \54972 , \54973 , \54974 ,
         \54975 , \54976 , \54977 , \54978 , \54979 , \54980 , \54981 , \54982 , \54983 , \54984 ,
         \54985 , \54986 , \54987 , \54988 , \54989 , \54990 , \54991 , \54992 , \54993 , \54994 ,
         \54995 , \54996 , \54997 , \54998 , \54999 , \55000 , \55001 , \55002 , \55003 , \55004 ,
         \55005 , \55006 , \55007 , \55008 , \55009 , \55010 , \55011 , \55012 , \55013 , \55014 ,
         \55015 , \55016 , \55017 , \55018 , \55019 , \55020 , \55021 , \55022 , \55023 , \55024 ,
         \55025 , \55026 , \55027 , \55028 , \55029 , \55030 , \55031 , \55032 , \55033 , \55034 ,
         \55035 , \55036 , \55037 , \55038 , \55039 , \55040 , \55041 , \55042 , \55043 , \55044 ,
         \55045 , \55046 , \55047 , \55048 , \55049 , \55050 , \55051 , \55052 , \55053 , \55054 ,
         \55055 , \55056 , \55057 , \55058 , \55059 , \55060 , \55061 , \55062 , \55063 , \55064 ,
         \55065 , \55066 , \55067 , \55068 , \55069 , \55070 , \55071 , \55072 , \55073 , \55074 ,
         \55075 , \55076 , \55077 , \55078 , \55079 , \55080 , \55081 , \55082 , \55083 , \55084 ,
         \55085 , \55086 , \55087 , \55088 , \55089 , \55090 , \55091 , \55092 , \55093 , \55094 ,
         \55095 , \55096 , \55097 , \55098 , \55099 , \55100 , \55101 , \55102 , \55103 , \55104 ,
         \55105 , \55106 , \55107 , \55108 , \55109 , \55110 , \55111 , \55112 , \55113 , \55114 ,
         \55115 , \55116 , \55117 , \55118 , \55119 , \55120 , \55121 , \55122 , \55123 , \55124 ,
         \55125 , \55126 , \55127 , \55128 , \55129 , \55130 , \55131 , \55132 , \55133 , \55134 ,
         \55135 , \55136 , \55137 , \55138 , \55139 , \55140 , \55141 , \55142 , \55143 , \55144 ,
         \55145 , \55146 , \55147 , \55148 , \55149 , \55150 , \55151 , \55152 , \55153 , \55154 ,
         \55155 , \55156 , \55157 , \55158 , \55159 , \55160 , \55161 , \55162 , \55163 , \55164 ,
         \55165 , \55166 , \55167 , \55168 , \55169 , \55170 , \55171 , \55172 , \55173 , \55174 ,
         \55175 , \55176 , \55177 , \55178 , \55179 , \55180 , \55181 , \55182 , \55183 , \55184 ,
         \55185 , \55186 , \55187 , \55188 , \55189 , \55190 , \55191 , \55192 , \55193 , \55194 ,
         \55195 , \55196 , \55197 , \55198 , \55199 , \55200 , \55201 , \55202 , \55203 , \55204 ,
         \55205 , \55206 , \55207 , \55208 , \55209 , \55210 , \55211 , \55212 , \55213 , \55214 ,
         \55215 , \55216 , \55217 , \55218 , \55219 , \55220 , \55221 , \55222 , \55223 , \55224 ,
         \55225 , \55226 , \55227 , \55228 , \55229 , \55230 , \55231 , \55232 , \55233 , \55234 ,
         \55235 , \55236 , \55237 , \55238 , \55239 , \55240 , \55241 , \55242 , \55243 , \55244 ,
         \55245 , \55246 , \55247 , \55248 , \55249 , \55250 , \55251 , \55252 , \55253 , \55254 ,
         \55255 , \55256 , \55257 , \55258 , \55259 , \55260 , \55261 , \55262 , \55263 , \55264 ,
         \55265 , \55266 , \55267 , \55268 , \55269 , \55270 , \55271 , \55272 , \55273 , \55274 ,
         \55275 , \55276 , \55277 , \55278 , \55279 , \55280 , \55281 , \55282 , \55283 , \55284 ,
         \55285 , \55286 , \55287 , \55288 , \55289 , \55290 , \55291 , \55292 , \55293 , \55294 ,
         \55295 , \55296 , \55297 , \55298 , \55299 , \55300 , \55301 , \55302 , \55303 , \55304 ,
         \55305 , \55306 , \55307 , \55308 , \55309 , \55310 , \55311 , \55312 , \55313 , \55314 ,
         \55315 , \55316 , \55317 , \55318 , \55319 , \55320 , \55321 , \55322 , \55323 , \55324 ,
         \55325 , \55326 , \55327 , \55328 , \55329 , \55330 , \55331 , \55332 , \55333 , \55334 ,
         \55335 , \55336 , \55337 , \55338 , \55339 , \55340 , \55341 , \55342 , \55343 , \55344 ,
         \55345 , \55346 , \55347 , \55348 , \55349 , \55350 , \55351 , \55352 , \55353 , \55354 ,
         \55355 , \55356 , \55357 , \55358 , \55359 , \55360 , \55361 , \55362 , \55363 , \55364 ,
         \55365 , \55366 , \55367 , \55368 , \55369 , \55370 , \55371 , \55372 , \55373 , \55374 ,
         \55375 , \55376 , \55377 , \55378 , \55379 , \55380 , \55381 , \55382 , \55383 , \55384 ,
         \55385 , \55386 , \55387 , \55388 , \55389 , \55390 , \55391 , \55392 , \55393 , \55394 ,
         \55395 , \55396 , \55397 , \55398 , \55399 , \55400 , \55401 , \55402 , \55403 , \55404 ,
         \55405 , \55406 , \55407 , \55408 , \55409 , \55410 , \55411 , \55412 , \55413 , \55414 ,
         \55415 , \55416 , \55417 , \55418 , \55419 , \55420 , \55421 , \55422 , \55423 , \55424 ,
         \55425 , \55426 , \55427 , \55428 , \55429 , \55430 , \55431 , \55432 , \55433 , \55434 ,
         \55435 , \55436 , \55437 , \55438 , \55439 , \55440 , \55441 , \55442 , \55443 , \55444 ,
         \55445 , \55446 , \55447 , \55448 , \55449 , \55450 , \55451 , \55452 , \55453 , \55454 ,
         \55455 , \55456 , \55457 , \55458 , \55459 , \55460 , \55461 , \55462 , \55463 , \55464 ,
         \55465 , \55466 , \55467 , \55468 , \55469 , \55470 , \55471 , \55472 , \55473 , \55474 ,
         \55475 , \55476 , \55477 , \55478 , \55479 , \55480 , \55481 , \55482 , \55483 , \55484 ,
         \55485 , \55486 , \55487 , \55488 , \55489 , \55490 , \55491 , \55492 , \55493 , \55494 ,
         \55495 , \55496 , \55497 , \55498 , \55499 , \55500 , \55501 , \55502 , \55503 , \55504 ,
         \55505 , \55506 , \55507 , \55508 , \55509 , \55510 , \55511 , \55512 , \55513 , \55514 ,
         \55515 , \55516 , \55517 , \55518 , \55519 , \55520 , \55521 , \55522 , \55523 , \55524 ,
         \55525 , \55526 , \55527 , \55528 , \55529 , \55530 , \55531 , \55532 , \55533 , \55534 ,
         \55535 , \55536 , \55537 , \55538 , \55539 , \55540 , \55541 , \55542 , \55543 , \55544 ,
         \55545 , \55546 , \55547 , \55548 , \55549 , \55550 , \55551 , \55552 , \55553 , \55554 ,
         \55555 , \55556 , \55557 , \55558 , \55559 , \55560 , \55561 , \55562 , \55563 , \55564 ,
         \55565 , \55566 , \55567 , \55568 , \55569 , \55570 , \55571 , \55572 , \55573 , \55574 ,
         \55575 , \55576 , \55577 , \55578 , \55579 , \55580 , \55581 , \55582 , \55583 , \55584 ,
         \55585 , \55586 , \55587 , \55588 , \55589 , \55590 , \55591 , \55592 , \55593 , \55594 ,
         \55595 , \55596 , \55597 , \55598 , \55599 , \55600 , \55601 , \55602 , \55603 , \55604 ,
         \55605 , \55606 , \55607 , \55608 , \55609 , \55610 , \55611 , \55612 , \55613 , \55614 ,
         \55615 , \55616 , \55617 , \55618 , \55619 , \55620 , \55621 , \55622 , \55623 , \55624 ,
         \55625 , \55626 , \55627 , \55628 , \55629 , \55630 , \55631 , \55632 , \55633 , \55634 ,
         \55635 , \55636 , \55637 , \55638 , \55639 , \55640 , \55641 , \55642 , \55643 , \55644 ,
         \55645 , \55646 , \55647 , \55648 , \55649 , \55650 , \55651 , \55652 , \55653 , \55654 ,
         \55655 , \55656 , \55657 , \55658 , \55659 , \55660 , \55661 , \55662 , \55663 , \55664 ,
         \55665 , \55666 , \55667 , \55668 , \55669 , \55670 , \55671 , \55672 , \55673 , \55674 ,
         \55675 , \55676 , \55677 , \55678 , \55679 , \55680 , \55681 , \55682 , \55683 , \55684 ,
         \55685 , \55686 , \55687 , \55688 , \55689 , \55690 , \55691 , \55692 , \55693 , \55694 ,
         \55695 , \55696 , \55697 , \55698 , \55699 , \55700 , \55701 , \55702 , \55703 , \55704 ,
         \55705 , \55706 , \55707 , \55708 , \55709 , \55710 , \55711 , \55712 , \55713 , \55714 ,
         \55715 , \55716 , \55717 , \55718 , \55719 , \55720 , \55721 , \55722 , \55723 , \55724 ,
         \55725 , \55726 , \55727 , \55728 , \55729 , \55730 , \55731 , \55732 , \55733 , \55734 ,
         \55735 , \55736 , \55737 , \55738 , \55739 , \55740 , \55741 , \55742 , \55743 , \55744 ,
         \55745 , \55746 , \55747 , \55748 , \55749 , \55750 , \55751 , \55752 , \55753 , \55754 ,
         \55755 , \55756 , \55757 , \55758 , \55759 , \55760 , \55761 , \55762 , \55763 , \55764 ,
         \55765 , \55766 , \55767 , \55768 , \55769 , \55770 , \55771 , \55772 , \55773 , \55774 ,
         \55775 , \55776 , \55777 , \55778 , \55779 , \55780 , \55781 , \55782 , \55783 , \55784 ,
         \55785 , \55786 , \55787 , \55788 , \55789 , \55790 , \55791 , \55792 , \55793 , \55794 ,
         \55795 , \55796 , \55797 , \55798 , \55799 , \55800 , \55801 , \55802 , \55803 , \55804 ,
         \55805 , \55806 , \55807 , \55808 , \55809 , \55810 , \55811 , \55812 , \55813 , \55814 ,
         \55815 , \55816 , \55817 , \55818 , \55819 , \55820 , \55821 , \55822 , \55823 , \55824 ,
         \55825 , \55826 , \55827 , \55828 , \55829 , \55830 , \55831 , \55832 , \55833 , \55834 ,
         \55835 , \55836 , \55837 , \55838 , \55839 , \55840 , \55841 , \55842 , \55843 , \55844 ,
         \55845 , \55846 , \55847 , \55848 , \55849 , \55850 , \55851 , \55852 , \55853 , \55854 ,
         \55855 , \55856 , \55857 , \55858 , \55859 , \55860 , \55861 , \55862 , \55863 , \55864 ,
         \55865 , \55866 , \55867 , \55868 , \55869 , \55870 , \55871 , \55872 , \55873 , \55874 ,
         \55875 , \55876 , \55877 , \55878 , \55879 , \55880 , \55881 , \55882 , \55883 , \55884 ,
         \55885 , \55886 , \55887 , \55888 , \55889 , \55890 , \55891 , \55892 , \55893 , \55894 ,
         \55895 , \55896 , \55897 , \55898 , \55899 , \55900 , \55901 , \55902 , \55903 , \55904 ,
         \55905 , \55906 , \55907 , \55908 , \55909 , \55910 , \55911 , \55912 , \55913 , \55914 ,
         \55915 , \55916 , \55917 , \55918 , \55919 , \55920 , \55921 , \55922 , \55923 , \55924 ,
         \55925 , \55926 , \55927 , \55928 , \55929 , \55930 , \55931 , \55932 , \55933 , \55934 ,
         \55935 , \55936 , \55937 , \55938 , \55939 , \55940 , \55941 , \55942 , \55943 , \55944 ,
         \55945 , \55946 , \55947 , \55948 , \55949 , \55950 , \55951 , \55952 , \55953 , \55954 ,
         \55955 , \55956 , \55957 , \55958 , \55959 , \55960 , \55961 , \55962 , \55963 , \55964 ,
         \55965 , \55966 , \55967 , \55968 , \55969 , \55970 , \55971 , \55972 , \55973 , \55974 ,
         \55975 , \55976 , \55977 , \55978 , \55979 , \55980 , \55981 , \55982 , \55983 , \55984 ,
         \55985 , \55986 , \55987 , \55988 , \55989 , \55990 , \55991 , \55992 , \55993 , \55994 ,
         \55995 , \55996 , \55997 , \55998 , \55999 , \56000 , \56001 , \56002 , \56003 , \56004 ,
         \56005 , \56006 , \56007 , \56008 , \56009 , \56010 , \56011 , \56012 , \56013 , \56014 ,
         \56015 , \56016 , \56017 , \56018 , \56019 , \56020 , \56021 , \56022 , \56023 , \56024 ,
         \56025 , \56026 , \56027 , \56028 , \56029 , \56030 , \56031 , \56032 , \56033 , \56034 ,
         \56035 , \56036 , \56037 , \56038 , \56039 , \56040 , \56041 , \56042 , \56043 , \56044 ,
         \56045 , \56046 , \56047 , \56048 , \56049 , \56050 , \56051 , \56052 , \56053 , \56054 ,
         \56055 , \56056 , \56057 , \56058 , \56059 , \56060 , \56061 , \56062 , \56063 , \56064 ,
         \56065 , \56066 , \56067 , \56068 , \56069 , \56070 , \56071 , \56072 , \56073 , \56074 ,
         \56075 , \56076 , \56077 , \56078 , \56079 , \56080 , \56081 , \56082 , \56083 , \56084 ,
         \56085 , \56086 , \56087 , \56088 , \56089 , \56090 , \56091 , \56092 , \56093 , \56094 ,
         \56095 , \56096 , \56097 , \56098 , \56099 , \56100 , \56101 , \56102 , \56103 , \56104 ,
         \56105 , \56106 , \56107 , \56108 , \56109 , \56110 , \56111 , \56112 , \56113 , \56114 ,
         \56115 , \56116 , \56117 , \56118 , \56119 , \56120 , \56121 , \56122 , \56123 , \56124 ,
         \56125 , \56126 , \56127 , \56128 , \56129 , \56130 , \56131 , \56132 , \56133 , \56134 ,
         \56135 , \56136 , \56137 , \56138 , \56139 , \56140 , \56141 , \56142 , \56143 , \56144 ,
         \56145 , \56146 , \56147 , \56148 , \56149 , \56150 , \56151 , \56152 , \56153 , \56154 ,
         \56155 , \56156 , \56157 , \56158 , \56159 , \56160 , \56161 , \56162 , \56163 , \56164 ,
         \56165 , \56166 , \56167 , \56168 , \56169 , \56170 , \56171 , \56172 , \56173 , \56174 ,
         \56175 , \56176 , \56177 , \56178 , \56179 , \56180 , \56181 , \56182 , \56183 , \56184 ,
         \56185 , \56186 , \56187 , \56188 , \56189 , \56190 , \56191 , \56192 , \56193 , \56194 ,
         \56195 , \56196 , \56197 , \56198 , \56199 , \56200 , \56201 , \56202 , \56203 , \56204 ,
         \56205 , \56206 , \56207 , \56208 , \56209 , \56210 , \56211 , \56212 , \56213 , \56214 ,
         \56215 , \56216 , \56217 , \56218 , \56219 , \56220 , \56221 , \56222 , \56223 , \56224 ,
         \56225 , \56226 , \56227 , \56228 , \56229 , \56230 , \56231 , \56232 , \56233 , \56234 ,
         \56235 , \56236 , \56237 , \56238 , \56239 , \56240 , \56241 , \56242 , \56243 , \56244 ,
         \56245 , \56246 , \56247 , \56248 , \56249 , \56250 , \56251 , \56252 , \56253 , \56254 ,
         \56255 , \56256 , \56257 , \56258 , \56259 , \56260 , \56261 , \56262 , \56263 , \56264 ,
         \56265 , \56266 , \56267 , \56268 , \56269 , \56270 , \56271 , \56272 , \56273 , \56274 ,
         \56275 , \56276 , \56277 , \56278 , \56279 , \56280 , \56281 , \56282 , \56283 , \56284 ,
         \56285 , \56286 , \56287 , \56288 , \56289 , \56290 , \56291 , \56292 , \56293 , \56294 ,
         \56295 , \56296 , \56297 , \56298 , \56299 , \56300 , \56301 , \56302 , \56303 , \56304 ,
         \56305 , \56306 , \56307 , \56308 , \56309 , \56310 , \56311 , \56312 , \56313 , \56314 ,
         \56315 , \56316 , \56317 , \56318 , \56319 , \56320 , \56321 , \56322 , \56323 , \56324 ,
         \56325 , \56326 , \56327 , \56328 , \56329 , \56330 , \56331 , \56332 , \56333 , \56334 ,
         \56335 , \56336 , \56337 , \56338 , \56339 , \56340 , \56341 , \56342 , \56343 , \56344 ,
         \56345 , \56346 , \56347 , \56348 , \56349 , \56350 , \56351 , \56352 , \56353 , \56354 ,
         \56355 , \56356 , \56357 , \56358 , \56359 , \56360 , \56361 , \56362 , \56363 , \56364 ,
         \56365 , \56366 , \56367 , \56368 , \56369 , \56370 , \56371 , \56372 , \56373 , \56374 ,
         \56375 , \56376 , \56377 , \56378 , \56379 , \56380 , \56381 , \56382 , \56383 , \56384 ,
         \56385 , \56386 , \56387 , \56388 , \56389 , \56390 , \56391 , \56392 , \56393 , \56394 ,
         \56395 , \56396 , \56397 , \56398 , \56399 , \56400 , \56401 , \56402 , \56403 , \56404 ,
         \56405 , \56406 , \56407 , \56408 , \56409 , \56410 , \56411 , \56412 , \56413 , \56414 ,
         \56415 , \56416 , \56417 , \56418 , \56419 , \56420 , \56421 , \56422 , \56423 , \56424 ,
         \56425 , \56426 , \56427 , \56428 , \56429 , \56430 , \56431 , \56432 , \56433 , \56434 ,
         \56435 , \56436 , \56437 , \56438 , \56439 , \56440 , \56441 , \56442 , \56443 , \56444 ,
         \56445 , \56446 , \56447 , \56448 , \56449 , \56450 , \56451 , \56452 , \56453 , \56454 ,
         \56455 , \56456 , \56457 , \56458 , \56459 , \56460 , \56461 , \56462 , \56463 , \56464 ,
         \56465 , \56466 , \56467 , \56468 , \56469 , \56470 , \56471 , \56472 , \56473 , \56474 ,
         \56475 , \56476 , \56477 , \56478 , \56479 , \56480 , \56481 , \56482 , \56483 , \56484 ,
         \56485 , \56486 , \56487 , \56488 , \56489 , \56490 , \56491 , \56492 , \56493 , \56494 ,
         \56495 , \56496 , \56497 , \56498 , \56499 , \56500 , \56501 , \56502 , \56503 , \56504 ,
         \56505 , \56506 , \56507 , \56508 , \56509 , \56510 , \56511 , \56512 , \56513 , \56514 ,
         \56515 , \56516 , \56517 , \56518 , \56519 , \56520 , \56521 , \56522 , \56523 , \56524 ,
         \56525 , \56526 , \56527 , \56528 , \56529 , \56530 , \56531 , \56532 , \56533 , \56534 ,
         \56535 , \56536 , \56537 , \56538 , \56539 , \56540 , \56541 , \56542 , \56543 , \56544 ,
         \56545 , \56546 , \56547 , \56548 , \56549 , \56550 , \56551 , \56552 , \56553 , \56554 ,
         \56555 , \56556 , \56557 , \56558 , \56559 , \56560 , \56561 , \56562 , \56563 , \56564 ,
         \56565 , \56566 , \56567 , \56568 , \56569 , \56570 , \56571 , \56572 , \56573 , \56574 ,
         \56575 , \56576 , \56577 , \56578 , \56579 , \56580 , \56581 , \56582 , \56583 , \56584 ,
         \56585 , \56586 , \56587 , \56588 , \56589 , \56590 , \56591 , \56592 , \56593 , \56594 ,
         \56595 , \56596 , \56597 , \56598 , \56599 , \56600 , \56601 , \56602 , \56603 , \56604 ,
         \56605 , \56606 , \56607 , \56608 , \56609 , \56610 , \56611 , \56612 , \56613 , \56614 ,
         \56615 , \56616 , \56617 , \56618 , \56619 , \56620 , \56621 , \56622 , \56623 , \56624 ,
         \56625 , \56626 , \56627 , \56628 , \56629 , \56630 , \56631 , \56632 , \56633 , \56634 ,
         \56635 , \56636 , \56637 , \56638 , \56639 , \56640 , \56641 , \56642 , \56643 , \56644 ,
         \56645 , \56646 , \56647 , \56648 , \56649 , \56650 , \56651 , \56652 , \56653 , \56654 ,
         \56655 , \56656 , \56657 , \56658 , \56659 , \56660 , \56661 , \56662 , \56663 , \56664 ,
         \56665 , \56666 , \56667 , \56668 , \56669 , \56670 , \56671 , \56672 , \56673 , \56674 ,
         \56675 , \56676 , \56677 , \56678 , \56679 , \56680 , \56681 , \56682 , \56683 , \56684 ,
         \56685 , \56686 , \56687 , \56688 , \56689 , \56690 , \56691 , \56692 , \56693 , \56694 ,
         \56695 , \56696 , \56697 , \56698 , \56699 , \56700 , \56701 , \56702 , \56703 , \56704 ,
         \56705 , \56706 , \56707 , \56708 , \56709 , \56710 , \56711 , \56712 , \56713 , \56714 ,
         \56715 , \56716 , \56717 , \56718 , \56719 , \56720 , \56721 , \56722 , \56723 , \56724 ,
         \56725 , \56726 , \56727 , \56728 , \56729 , \56730 , \56731 , \56732 , \56733 , \56734 ,
         \56735 , \56736 , \56737 , \56738 , \56739 , \56740 , \56741 , \56742 , \56743 , \56744 ,
         \56745 , \56746 , \56747 , \56748 , \56749 , \56750 , \56751 , \56752 , \56753 , \56754 ,
         \56755 , \56756 , \56757 , \56758 , \56759 , \56760 , \56761 , \56762 , \56763 , \56764 ,
         \56765 , \56766 , \56767 , \56768 , \56769 , \56770 , \56771 , \56772 , \56773 , \56774 ,
         \56775 , \56776 , \56777 , \56778 , \56779 , \56780 , \56781 , \56782 , \56783 , \56784 ,
         \56785 , \56786 , \56787 , \56788 , \56789 , \56790 , \56791 , \56792 , \56793 , \56794 ,
         \56795 , \56796 , \56797 , \56798 , \56799 , \56800 , \56801 , \56802 , \56803 , \56804 ,
         \56805 , \56806 , \56807 , \56808 , \56809 , \56810 , \56811 , \56812 , \56813 , \56814 ,
         \56815 , \56816 , \56817 , \56818 , \56819 , \56820 , \56821 , \56822 , \56823 , \56824 ,
         \56825 , \56826 , \56827 , \56828 , \56829 , \56830 , \56831 , \56832 , \56833 , \56834 ,
         \56835 , \56836 , \56837 , \56838 , \56839 , \56840 , \56841 , \56842 , \56843 , \56844 ,
         \56845 , \56846 , \56847 , \56848 , \56849 , \56850 , \56851 , \56852 , \56853 , \56854 ,
         \56855 , \56856 , \56857 , \56858 , \56859 , \56860 , \56861 , \56862 , \56863 , \56864 ,
         \56865 , \56866 , \56867 , \56868 , \56869 , \56870 , \56871 , \56872 , \56873 , \56874 ,
         \56875 , \56876 , \56877 , \56878 , \56879 , \56880 , \56881 , \56882 , \56883 , \56884 ,
         \56885 , \56886 , \56887 , \56888 , \56889 , \56890 , \56891 , \56892 , \56893 , \56894 ,
         \56895 , \56896 , \56897 , \56898 , \56899 , \56900 , \56901 , \56902 , \56903 , \56904 ,
         \56905 , \56906 , \56907 , \56908 , \56909 , \56910 , \56911 , \56912 , \56913 , \56914 ,
         \56915 , \56916 , \56917 , \56918 , \56919 , \56920 , \56921 , \56922 , \56923 , \56924 ,
         \56925 , \56926 , \56927 , \56928 , \56929 , \56930 , \56931 , \56932 , \56933 , \56934 ,
         \56935 , \56936 , \56937 , \56938 , \56939 , \56940 , \56941 , \56942 , \56943 , \56944 ,
         \56945 , \56946 , \56947 , \56948 , \56949 , \56950 , \56951 , \56952 , \56953 , \56954 ,
         \56955 , \56956 , \56957 , \56958 , \56959 , \56960 , \56961 , \56962 , \56963 , \56964 ,
         \56965 , \56966 , \56967 , \56968 , \56969 , \56970 , \56971 , \56972 , \56973 , \56974 ,
         \56975 , \56976 , \56977 , \56978 , \56979 , \56980 , \56981 , \56982 , \56983 , \56984 ,
         \56985 , \56986 , \56987 , \56988 , \56989 , \56990 , \56991 , \56992 , \56993 , \56994 ,
         \56995 , \56996 , \56997 , \56998 , \56999 , \57000 , \57001 , \57002 , \57003 , \57004 ,
         \57005 , \57006 , \57007 , \57008 , \57009 , \57010 , \57011 , \57012 , \57013 , \57014 ,
         \57015 , \57016 , \57017 , \57018 , \57019 , \57020 , \57021 , \57022 , \57023 , \57024 ,
         \57025 , \57026 , \57027 , \57028 , \57029 , \57030 , \57031 , \57032 , \57033 , \57034 ,
         \57035 , \57036 , \57037 , \57038 , \57039 , \57040 , \57041 , \57042 , \57043 , \57044 ,
         \57045 , \57046 , \57047 , \57048 , \57049 , \57050 , \57051 , \57052 , \57053 , \57054 ,
         \57055 , \57056 , \57057 , \57058 , \57059 , \57060 , \57061 , \57062 , \57063 , \57064 ,
         \57065 , \57066 , \57067 , \57068 , \57069 , \57070 , \57071 , \57072 , \57073 , \57074 ,
         \57075 , \57076 , \57077 , \57078 , \57079 , \57080 , \57081 , \57082 , \57083 , \57084 ,
         \57085 , \57086 , \57087 , \57088 , \57089 , \57090 , \57091 , \57092 , \57093 , \57094 ,
         \57095 , \57096 , \57097 , \57098 , \57099 , \57100 , \57101 , \57102 , \57103 , \57104 ,
         \57105 , \57106 , \57107 , \57108 , \57109 , \57110 , \57111 , \57112 , \57113 , \57114 ,
         \57115 , \57116 , \57117 , \57118 , \57119 , \57120 , \57121 , \57122 , \57123 , \57124 ,
         \57125 , \57126 , \57127 , \57128 , \57129 , \57130 , \57131 , \57132 , \57133 , \57134 ,
         \57135 , \57136 , \57137 , \57138 , \57139 , \57140 , \57141 , \57142 , \57143 , \57144 ,
         \57145 , \57146 , \57147 , \57148 , \57149 , \57150 , \57151 , \57152 , \57153 , \57154 ,
         \57155 , \57156 , \57157 , \57158 , \57159 , \57160 , \57161 , \57162 , \57163 , \57164 ,
         \57165 , \57166 , \57167 , \57168 , \57169 , \57170 , \57171 , \57172 , \57173 , \57174 ,
         \57175 , \57176 , \57177 , \57178 , \57179 , \57180 , \57181 , \57182 , \57183 , \57184 ,
         \57185 , \57186 , \57187 , \57188 , \57189 , \57190 , \57191 , \57192 , \57193 , \57194 ,
         \57195 , \57196 , \57197 , \57198 , \57199 , \57200 , \57201 , \57202 , \57203 , \57204 ,
         \57205 , \57206 , \57207 , \57208 , \57209 , \57210 , \57211 , \57212 , \57213 , \57214 ,
         \57215 , \57216 , \57217 , \57218 , \57219 , \57220 , \57221 , \57222 , \57223 , \57224 ,
         \57225 , \57226 , \57227 , \57228 , \57229 , \57230 , \57231 , \57232 , \57233 , \57234 ,
         \57235 , \57236 , \57237 , \57238 , \57239 , \57240 , \57241 , \57242 , \57243 , \57244 ,
         \57245 , \57246 , \57247 , \57248 , \57249 , \57250 , \57251 , \57252 , \57253 , \57254 ,
         \57255 , \57256 , \57257 , \57258 , \57259 , \57260 , \57261 , \57262 , \57263 , \57264 ,
         \57265 , \57266 , \57267 , \57268 , \57269 , \57270 , \57271 , \57272 , \57273 , \57274 ,
         \57275 , \57276 , \57277 , \57278 , \57279 , \57280 , \57281 , \57282 , \57283 , \57284 ,
         \57285 , \57286 , \57287 , \57288 , \57289 , \57290 , \57291 , \57292 , \57293 , \57294 ,
         \57295 , \57296 , \57297 , \57298 , \57299 , \57300 , \57301 , \57302 , \57303 , \57304 ,
         \57305 , \57306 , \57307 , \57308 , \57309 , \57310 , \57311 , \57312 , \57313 , \57314 ,
         \57315 , \57316 , \57317 , \57318 , \57319 , \57320 , \57321 , \57322 , \57323 , \57324 ,
         \57325 , \57326 , \57327 , \57328 , \57329 , \57330 , \57331 , \57332 , \57333 , \57334 ,
         \57335 , \57336 , \57337 , \57338 , \57339 , \57340 , \57341 , \57342 , \57343 , \57344 ,
         \57345 , \57346 , \57347 , \57348 , \57349 , \57350 , \57351 , \57352 , \57353 , \57354 ,
         \57355 , \57356 , \57357 , \57358 , \57359 , \57360 , \57361 , \57362 , \57363 , \57364 ,
         \57365 , \57366 , \57367 , \57368 , \57369 , \57370 , \57371 , \57372 , \57373 , \57374 ,
         \57375 , \57376 , \57377 , \57378 , \57379 , \57380 , \57381 , \57382 , \57383 , \57384 ,
         \57385 , \57386 , \57387 , \57388 , \57389 , \57390 , \57391 , \57392 , \57393 , \57394 ,
         \57395 , \57396 , \57397 , \57398 , \57399 , \57400 , \57401 , \57402 , \57403 , \57404 ,
         \57405 , \57406 , \57407 , \57408 , \57409 , \57410 , \57411 , \57412 , \57413 , \57414 ,
         \57415 , \57416 , \57417 , \57418 , \57419 , \57420 , \57421 , \57422 , \57423 , \57424 ,
         \57425 , \57426 , \57427 , \57428 , \57429 , \57430 , \57431 , \57432 , \57433 , \57434 ,
         \57435 , \57436 , \57437 , \57438 , \57439 , \57440 , \57441 , \57442 , \57443 , \57444 ,
         \57445 , \57446 , \57447 , \57448 , \57449 , \57450 , \57451 , \57452 , \57453 , \57454 ,
         \57455 , \57456 , \57457 , \57458 , \57459 , \57460 , \57461 , \57462 , \57463 , \57464 ,
         \57465 , \57466 , \57467 , \57468 , \57469 , \57470 , \57471 , \57472 , \57473 , \57474 ,
         \57475 , \57476 , \57477 , \57478 , \57479 , \57480 , \57481 , \57482 , \57483 , \57484 ,
         \57485 , \57486 , \57487 , \57488 , \57489 , \57490 , \57491 , \57492 , \57493 , \57494 ,
         \57495 , \57496 , \57497 , \57498 , \57499 , \57500 , \57501 , \57502 , \57503 , \57504 ,
         \57505 , \57506 , \57507 , \57508 , \57509 , \57510 , \57511 , \57512 , \57513 , \57514 ,
         \57515 , \57516 , \57517 , \57518 , \57519 , \57520 , \57521 , \57522 , \57523 , \57524 ,
         \57525 , \57526 , \57527 , \57528 , \57529 , \57530 , \57531 , \57532 , \57533 , \57534 ,
         \57535 , \57536 , \57537 , \57538 , \57539 , \57540 , \57541 , \57542 , \57543 , \57544 ,
         \57545 , \57546 , \57547 , \57548 , \57549 , \57550 , \57551 , \57552 , \57553 , \57554 ,
         \57555 , \57556 , \57557 , \57558 , \57559 , \57560 , \57561 , \57562 , \57563 , \57564 ,
         \57565 , \57566 , \57567 , \57568 , \57569 , \57570 , \57571 , \57572 , \57573 , \57574 ,
         \57575 , \57576 , \57577 , \57578 , \57579 , \57580 , \57581 , \57582 , \57583 , \57584 ,
         \57585 , \57586 , \57587 , \57588 , \57589 , \57590 , \57591 , \57592 , \57593 , \57594 ,
         \57595 , \57596 , \57597 , \57598 , \57599 , \57600 , \57601 , \57602 , \57603 , \57604 ,
         \57605 , \57606 , \57607 , \57608 , \57609 , \57610 , \57611 , \57612 , \57613 , \57614 ,
         \57615 , \57616 , \57617 , \57618 , \57619 , \57620 , \57621 , \57622 , \57623 , \57624 ,
         \57625 , \57626 , \57627 , \57628 , \57629 , \57630 , \57631 , \57632 , \57633 , \57634 ,
         \57635 , \57636 , \57637 , \57638 , \57639 , \57640 , \57641 , \57642 , \57643 , \57644 ,
         \57645 , \57646 , \57647 , \57648 , \57649 , \57650 , \57651 , \57652 , \57653 , \57654 ,
         \57655 , \57656 , \57657 , \57658 , \57659 , \57660 , \57661 , \57662 , \57663 , \57664 ,
         \57665 , \57666 , \57667 , \57668 , \57669 , \57670 , \57671 , \57672 , \57673 , \57674 ,
         \57675 , \57676 , \57677 , \57678 , \57679 , \57680 , \57681 , \57682 , \57683 , \57684 ,
         \57685 , \57686 , \57687 , \57688 , \57689 , \57690 , \57691 , \57692 , \57693 , \57694 ,
         \57695 , \57696 , \57697 , \57698 , \57699 , \57700 , \57701 , \57702 , \57703 , \57704 ,
         \57705 , \57706 , \57707 , \57708 , \57709 , \57710 , \57711 , \57712 , \57713 , \57714 ,
         \57715 , \57716 , \57717 , \57718 , \57719 , \57720 , \57721 , \57722 , \57723 , \57724 ,
         \57725 , \57726 , \57727 , \57728 , \57729 , \57730 , \57731 , \57732 , \57733 , \57734 ,
         \57735 , \57736 , \57737 , \57738 , \57739 , \57740 , \57741 , \57742 , \57743 , \57744 ,
         \57745 , \57746 , \57747 , \57748 , \57749 , \57750 , \57751 , \57752 , \57753 , \57754 ,
         \57755 , \57756 , \57757 , \57758 , \57759 , \57760 , \57761 , \57762 , \57763 , \57764 ,
         \57765 , \57766 , \57767 , \57768 , \57769 , \57770 , \57771 , \57772 , \57773 , \57774 ,
         \57775 , \57776 , \57777 , \57778 , \57779 , \57780 , \57781 , \57782 , \57783 , \57784 ,
         \57785 , \57786 , \57787 , \57788 , \57789 , \57790 , \57791 , \57792 , \57793 , \57794 ,
         \57795 , \57796 , \57797 , \57798 , \57799 , \57800 , \57801 , \57802 , \57803 , \57804 ,
         \57805 , \57806 , \57807 , \57808 , \57809 , \57810 , \57811 , \57812 , \57813 , \57814 ,
         \57815 , \57816 , \57817 , \57818 , \57819 , \57820 , \57821 , \57822 , \57823 , \57824 ,
         \57825 , \57826 , \57827 , \57828 , \57829 , \57830 , \57831 , \57832 , \57833 , \57834 ,
         \57835 , \57836 , \57837 , \57838 , \57839 , \57840 , \57841 , \57842 , \57843 , \57844 ,
         \57845 , \57846 , \57847 , \57848 , \57849 , \57850 , \57851 , \57852 , \57853 , \57854 ,
         \57855 , \57856 , \57857 , \57858 , \57859 , \57860 , \57861 , \57862 , \57863 , \57864 ,
         \57865 , \57866 , \57867 , \57868 , \57869 , \57870 , \57871 , \57872 , \57873 , \57874 ,
         \57875 , \57876 , \57877 , \57878 , \57879 , \57880 , \57881 , \57882 , \57883 , \57884 ,
         \57885 , \57886 , \57887 , \57888 , \57889 , \57890 , \57891 , \57892 , \57893 , \57894 ,
         \57895 , \57896 , \57897 , \57898 , \57899 , \57900 , \57901 , \57902 , \57903 , \57904 ,
         \57905 , \57906 , \57907 , \57908 , \57909 , \57910 , \57911 , \57912 , \57913 , \57914 ,
         \57915 , \57916 , \57917 , \57918 , \57919 , \57920 , \57921 , \57922 , \57923 , \57924 ,
         \57925 , \57926 , \57927 , \57928 , \57929 , \57930 , \57931 , \57932 , \57933 , \57934 ,
         \57935 , \57936 , \57937 , \57938 , \57939 , \57940 , \57941 , \57942 , \57943 , \57944 ,
         \57945 , \57946 , \57947 , \57948 , \57949 , \57950 , \57951 , \57952 , \57953 , \57954 ,
         \57955 , \57956 , \57957 , \57958 , \57959 , \57960 , \57961 , \57962 , \57963 , \57964 ,
         \57965 , \57966 , \57967 , \57968 , \57969 , \57970 , \57971 , \57972 , \57973 , \57974 ,
         \57975 , \57976 , \57977 , \57978 , \57979 , \57980 , \57981 , \57982 , \57983 , \57984 ,
         \57985 , \57986 , \57987 , \57988 , \57989 , \57990 , \57991 , \57992 , \57993 , \57994 ,
         \57995 , \57996 , \57997 , \57998 , \57999 , \58000 , \58001 , \58002 , \58003 , \58004 ,
         \58005 , \58006 , \58007 , \58008 , \58009 , \58010 , \58011 , \58012 , \58013 , \58014 ,
         \58015 , \58016 , \58017 , \58018 , \58019 , \58020 , \58021 , \58022 , \58023 , \58024 ,
         \58025 , \58026 , \58027 , \58028 , \58029 , \58030 , \58031 , \58032 , \58033 , \58034 ,
         \58035 , \58036 , \58037 , \58038 , \58039 , \58040 , \58041 , \58042 , \58043 , \58044 ,
         \58045 , \58046 , \58047 , \58048 , \58049 , \58050 , \58051 , \58052 , \58053 , \58054 ,
         \58055 , \58056 , \58057 , \58058 , \58059 , \58060 , \58061 , \58062 , \58063 , \58064 ,
         \58065 , \58066 , \58067 , \58068 , \58069 , \58070 , \58071 , \58072 , \58073 , \58074 ,
         \58075 , \58076 , \58077 , \58078 , \58079 , \58080 , \58081 , \58082 , \58083 , \58084 ,
         \58085 , \58086 , \58087 , \58088 , \58089 , \58090 , \58091 , \58092 , \58093 , \58094 ,
         \58095 , \58096 , \58097 , \58098 , \58099 , \58100 , \58101 , \58102 , \58103 , \58104 ,
         \58105 , \58106 , \58107 , \58108 , \58109 , \58110 , \58111 , \58112 , \58113 , \58114 ,
         \58115 , \58116 , \58117 , \58118 , \58119 , \58120 , \58121 , \58122 , \58123 , \58124 ,
         \58125 , \58126 , \58127 , \58128 , \58129 , \58130 , \58131 , \58132 , \58133 , \58134 ,
         \58135 , \58136 , \58137 , \58138 , \58139 , \58140 , \58141 , \58142 , \58143 , \58144 ,
         \58145 , \58146 , \58147 , \58148 , \58149 , \58150 , \58151 , \58152 , \58153 , \58154 ,
         \58155 , \58156 , \58157 , \58158 , \58159 , \58160 , \58161 , \58162 , \58163 , \58164 ,
         \58165 , \58166 , \58167 , \58168 , \58169 , \58170 , \58171 , \58172 , \58173 , \58174 ,
         \58175 , \58176 , \58177 , \58178 , \58179 , \58180 , \58181 , \58182 , \58183 , \58184 ,
         \58185 , \58186 , \58187 , \58188 , \58189 , \58190 , \58191 , \58192 , \58193 , \58194 ,
         \58195 , \58196 , \58197 , \58198 , \58199 , \58200 , \58201 , \58202 , \58203 , \58204 ,
         \58205 , \58206 , \58207 , \58208 , \58209 , \58210 , \58211 , \58212 , \58213 , \58214 ,
         \58215 , \58216 , \58217 , \58218 , \58219 , \58220 , \58221 , \58222 , \58223 , \58224 ,
         \58225 , \58226 , \58227 , \58228 , \58229 , \58230 , \58231 , \58232 , \58233 , \58234 ,
         \58235 , \58236 , \58237 , \58238 , \58239 , \58240 , \58241 , \58242 , \58243 , \58244 ,
         \58245 , \58246 , \58247 , \58248 , \58249 , \58250 , \58251 , \58252 , \58253 , \58254 ,
         \58255 , \58256 , \58257 , \58258 , \58259 , \58260 , \58261 , \58262 , \58263 , \58264 ,
         \58265 , \58266 , \58267 , \58268 , \58269 , \58270 , \58271 , \58272 , \58273 , \58274 ,
         \58275 , \58276 , \58277 , \58278 , \58279 , \58280 , \58281 , \58282 , \58283 , \58284 ,
         \58285 , \58286 , \58287 , \58288 , \58289 , \58290 , \58291 , \58292 , \58293 , \58294 ,
         \58295 , \58296 , \58297 , \58298 , \58299 , \58300 , \58301 , \58302 , \58303 , \58304 ,
         \58305 , \58306 , \58307 , \58308 , \58309 , \58310 , \58311 , \58312 , \58313 , \58314 ,
         \58315 , \58316 , \58317 , \58318 , \58319 , \58320 , \58321 , \58322 , \58323 , \58324 ,
         \58325 , \58326 , \58327 , \58328 , \58329 , \58330 , \58331 , \58332 , \58333 , \58334 ,
         \58335 , \58336 , \58337 , \58338 , \58339 , \58340 , \58341 , \58342 , \58343 , \58344 ,
         \58345 , \58346 , \58347 , \58348 , \58349 , \58350 , \58351 , \58352 , \58353 , \58354 ,
         \58355 , \58356 , \58357 , \58358 , \58359 , \58360 , \58361 , \58362 , \58363 , \58364 ,
         \58365 , \58366 , \58367 , \58368 , \58369 , \58370 , \58371 , \58372 , \58373 , \58374 ,
         \58375 , \58376 , \58377 , \58378 , \58379 , \58380 , \58381 , \58382 , \58383 , \58384 ,
         \58385 , \58386 , \58387 , \58388 , \58389 , \58390 , \58391 , \58392 , \58393 , \58394 ,
         \58395 , \58396 , \58397 , \58398 , \58399 , \58400 , \58401 , \58402 , \58403 , \58404 ,
         \58405 , \58406 , \58407 , \58408 , \58409 , \58410 , \58411 , \58412 , \58413 , \58414 ,
         \58415 , \58416 , \58417 , \58418 , \58419 , \58420 , \58421 , \58422 , \58423 , \58424 ,
         \58425 , \58426 , \58427 , \58428 , \58429 , \58430 , \58431 , \58432 , \58433 , \58434 ,
         \58435 , \58436 , \58437 , \58438 , \58439 , \58440 , \58441 , \58442 , \58443 , \58444 ,
         \58445 , \58446 , \58447 , \58448 , \58449 , \58450 , \58451 , \58452 , \58453 , \58454 ,
         \58455 , \58456 , \58457 , \58458 , \58459 , \58460 , \58461 , \58462 , \58463 , \58464 ,
         \58465 , \58466 , \58467 , \58468 , \58469 , \58470 , \58471 , \58472 , \58473 , \58474 ,
         \58475 , \58476 , \58477 , \58478 , \58479 , \58480 , \58481 , \58482 , \58483 , \58484 ,
         \58485 , \58486 , \58487 , \58488 , \58489 , \58490 , \58491 , \58492 , \58493 , \58494 ,
         \58495 , \58496 , \58497 , \58498 , \58499 , \58500 , \58501 , \58502 , \58503 , \58504 ,
         \58505 , \58506 , \58507 , \58508 , \58509 , \58510 , \58511 , \58512 , \58513 , \58514 ,
         \58515 , \58516 , \58517 , \58518 , \58519 , \58520 , \58521 , \58522 , \58523 , \58524 ,
         \58525 , \58526 , \58527 , \58528 , \58529 , \58530 , \58531 , \58532 , \58533 , \58534 ,
         \58535 , \58536 , \58537 , \58538 , \58539 , \58540 , \58541 , \58542 , \58543 , \58544 ,
         \58545 , \58546 , \58547 , \58548 , \58549 , \58550 , \58551 , \58552 , \58553 , \58554 ,
         \58555 , \58556 , \58557 , \58558 , \58559 , \58560 , \58561 , \58562 , \58563 , \58564 ,
         \58565 , \58566 , \58567 , \58568 , \58569 , \58570 , \58571 , \58572 , \58573 , \58574 ,
         \58575 , \58576 , \58577 , \58578 , \58579 , \58580 , \58581 , \58582 , \58583 , \58584 ,
         \58585 , \58586 , \58587 , \58588 , \58589 , \58590 , \58591 , \58592 , \58593 , \58594 ,
         \58595 , \58596 , \58597 , \58598 , \58599 , \58600 , \58601 , \58602 , \58603 , \58604 ,
         \58605 , \58606 , \58607 , \58608 , \58609 , \58610 , \58611 , \58612 , \58613 , \58614 ,
         \58615 , \58616 , \58617 , \58618 , \58619 , \58620 , \58621 , \58622 , \58623 , \58624 ,
         \58625 , \58626 , \58627 , \58628 , \58629 , \58630 , \58631 , \58632 , \58633 , \58634 ,
         \58635 , \58636 , \58637 , \58638 , \58639 , \58640 , \58641 , \58642 , \58643 , \58644 ,
         \58645 , \58646 , \58647 , \58648 , \58649 , \58650 , \58651 , \58652 , \58653 , \58654 ,
         \58655 , \58656 , \58657 , \58658 , \58659 , \58660 , \58661 , \58662 , \58663 , \58664 ,
         \58665 , \58666 , \58667 , \58668 , \58669 , \58670 , \58671 , \58672 , \58673 , \58674 ,
         \58675 , \58676 , \58677 , \58678 , \58679 , \58680 , \58681 , \58682 , \58683 , \58684 ,
         \58685 , \58686 , \58687 , \58688 , \58689 , \58690 , \58691 , \58692 , \58693 , \58694 ,
         \58695 , \58696 , \58697 , \58698 , \58699 , \58700 , \58701 , \58702 , \58703 , \58704 ,
         \58705 , \58706 , \58707 , \58708 , \58709 , \58710 , \58711 , \58712 , \58713 , \58714 ,
         \58715 , \58716 , \58717 , \58718 , \58719 , \58720 , \58721 , \58722 , \58723 , \58724 ,
         \58725 , \58726 , \58727 , \58728 , \58729 , \58730 , \58731 , \58732 , \58733 , \58734 ,
         \58735 , \58736 , \58737 , \58738 , \58739 , \58740 , \58741 , \58742 , \58743 , \58744 ,
         \58745 , \58746 , \58747 , \58748 , \58749 , \58750 , \58751 , \58752 , \58753 , \58754 ,
         \58755 , \58756 , \58757 , \58758 , \58759 , \58760 , \58761 , \58762 , \58763 , \58764 ,
         \58765 , \58766 , \58767 , \58768 , \58769 , \58770 , \58771 , \58772 , \58773 , \58774 ,
         \58775 , \58776 , \58777 , \58778 , \58779 , \58780 , \58781 , \58782 , \58783 , \58784 ,
         \58785 , \58786 , \58787 , \58788 , \58789 , \58790 , \58791 , \58792 , \58793 , \58794 ,
         \58795 , \58796 , \58797 , \58798 , \58799 , \58800 , \58801 , \58802 , \58803 , \58804 ,
         \58805 , \58806 , \58807 , \58808 , \58809 , \58810 , \58811 , \58812 , \58813 , \58814 ,
         \58815 , \58816 , \58817 , \58818 , \58819 , \58820 , \58821 , \58822 , \58823 , \58824 ,
         \58825 , \58826 , \58827 , \58828 , \58829 , \58830 , \58831 , \58832 , \58833 , \58834 ,
         \58835 , \58836 , \58837 , \58838 , \58839 , \58840 , \58841 , \58842 , \58843 , \58844 ,
         \58845 , \58846 , \58847 , \58848 , \58849 , \58850 , \58851 , \58852 , \58853 , \58854 ,
         \58855 , \58856 , \58857 , \58858 , \58859 , \58860 , \58861 , \58862 , \58863 , \58864 ,
         \58865 , \58866 , \58867 , \58868 , \58869 , \58870 , \58871 , \58872 , \58873 , \58874 ,
         \58875 , \58876 , \58877 , \58878 , \58879 , \58880 , \58881 , \58882 , \58883 , \58884 ,
         \58885 , \58886 , \58887 , \58888 , \58889 , \58890 , \58891 , \58892 , \58893 , \58894 ,
         \58895 , \58896 , \58897 , \58898 , \58899 , \58900 , \58901 , \58902 , \58903 , \58904 ,
         \58905 , \58906 , \58907 , \58908 , \58909 , \58910 , \58911 , \58912 , \58913 , \58914 ,
         \58915 , \58916 , \58917 , \58918 , \58919 , \58920 , \58921 , \58922 , \58923 , \58924 ,
         \58925 , \58926 , \58927 , \58928 , \58929 , \58930 , \58931 , \58932 , \58933 , \58934 ,
         \58935 , \58936 , \58937 , \58938 , \58939 , \58940 , \58941 , \58942 , \58943 , \58944 ,
         \58945 , \58946 , \58947 , \58948 , \58949 , \58950 , \58951 , \58952 , \58953 , \58954 ,
         \58955 , \58956 , \58957 , \58958 , \58959 , \58960 , \58961 , \58962 , \58963 , \58964 ,
         \58965 , \58966 , \58967 , \58968 , \58969 , \58970 , \58971 , \58972 , \58973 , \58974 ,
         \58975 , \58976 , \58977 , \58978 , \58979 , \58980 , \58981 , \58982 , \58983 , \58984 ,
         \58985 , \58986 , \58987 , \58988 , \58989 , \58990 , \58991 , \58992 , \58993 , \58994 ,
         \58995 , \58996 , \58997 , \58998 , \58999 , \59000 , \59001 , \59002 , \59003 , \59004 ,
         \59005 , \59006 , \59007 , \59008 , \59009 , \59010 , \59011 , \59012 , \59013 , \59014 ,
         \59015 , \59016 , \59017 , \59018 , \59019 , \59020 , \59021 , \59022 , \59023 , \59024 ,
         \59025 , \59026 , \59027 , \59028 , \59029 , \59030 , \59031 , \59032 , \59033 , \59034 ,
         \59035 , \59036 , \59037 , \59038 , \59039 , \59040 , \59041 , \59042 , \59043 , \59044 ,
         \59045 , \59046 , \59047 , \59048 , \59049 , \59050 , \59051 , \59052 , \59053 , \59054 ,
         \59055 , \59056 , \59057 , \59058 , \59059 , \59060 , \59061 , \59062 , \59063 , \59064 ,
         \59065 , \59066 , \59067 , \59068 , \59069 , \59070 , \59071 , \59072 , \59073 , \59074 ,
         \59075 , \59076 , \59077 , \59078 , \59079 , \59080 , \59081 , \59082 , \59083 , \59084 ,
         \59085 , \59086 , \59087 , \59088 , \59089 , \59090 , \59091 , \59092 , \59093 , \59094 ,
         \59095 , \59096 , \59097 , \59098 , \59099 , \59100 , \59101 , \59102 , \59103 , \59104 ,
         \59105 , \59106 , \59107 , \59108 , \59109 , \59110 , \59111 , \59112 , \59113 , \59114 ,
         \59115 , \59116 , \59117 , \59118 , \59119 , \59120 , \59121 , \59122 , \59123 , \59124 ,
         \59125 , \59126 , \59127 , \59128 , \59129 , \59130 , \59131 , \59132 , \59133 , \59134 ,
         \59135 , \59136 , \59137 , \59138 , \59139 , \59140 , \59141 , \59142 , \59143 , \59144 ,
         \59145 , \59146 , \59147 , \59148 , \59149 , \59150 , \59151 , \59152 , \59153 , \59154 ,
         \59155 , \59156 , \59157 , \59158 , \59159 , \59160 , \59161 , \59162 , \59163 , \59164 ,
         \59165 , \59166 , \59167 , \59168 , \59169 , \59170 , \59171 , \59172 , \59173 , \59174 ,
         \59175 , \59176 , \59177 , \59178 , \59179 , \59180 , \59181 , \59182 , \59183 , \59184 ,
         \59185 , \59186 , \59187 , \59188 , \59189 , \59190 , \59191 , \59192 , \59193 , \59194 ,
         \59195 , \59196 , \59197 , \59198 , \59199 , \59200 , \59201 , \59202 , \59203 , \59204 ,
         \59205 , \59206 , \59207 , \59208 , \59209 , \59210 , \59211 , \59212 , \59213 , \59214 ,
         \59215 , \59216 , \59217 , \59218 , \59219 , \59220 , \59221 , \59222 , \59223 , \59224 ,
         \59225 , \59226 , \59227 , \59228 , \59229 , \59230 , \59231 , \59232 , \59233 , \59234 ,
         \59235 , \59236 , \59237 , \59238 , \59239 , \59240 , \59241 , \59242 , \59243 , \59244 ,
         \59245 , \59246 , \59247 , \59248 , \59249 , \59250 , \59251 , \59252 , \59253 , \59254 ,
         \59255 , \59256 , \59257 , \59258 , \59259 , \59260 , \59261 , \59262 , \59263 , \59264 ,
         \59265 , \59266 , \59267 , \59268 , \59269 , \59270 , \59271 , \59272 , \59273 , \59274 ,
         \59275 , \59276 , \59277 , \59278 , \59279 , \59280 , \59281 , \59282 , \59283 , \59284 ,
         \59285 , \59286 , \59287 , \59288 , \59289 , \59290 , \59291 , \59292 , \59293 , \59294 ,
         \59295 , \59296 , \59297 , \59298 , \59299 , \59300 , \59301 , \59302 , \59303 , \59304 ,
         \59305 , \59306 , \59307 , \59308 , \59309 , \59310 , \59311 , \59312 , \59313 , \59314 ,
         \59315 , \59316 , \59317 , \59318 , \59319 , \59320 , \59321 , \59322 , \59323 , \59324 ,
         \59325 , \59326 , \59327 , \59328 , \59329 , \59330 , \59331 , \59332 , \59333 , \59334 ,
         \59335 , \59336 , \59337 , \59338 , \59339 , \59340 , \59341 , \59342 , \59343 , \59344 ,
         \59345 , \59346 , \59347 , \59348 , \59349 , \59350 , \59351 , \59352 , \59353 , \59354 ,
         \59355 , \59356 , \59357 , \59358 , \59359 , \59360 , \59361 , \59362 , \59363 , \59364 ,
         \59365 , \59366 , \59367 , \59368 , \59369 , \59370 , \59371 , \59372 , \59373 , \59374 ,
         \59375 , \59376 , \59377 , \59378 , \59379 , \59380 , \59381 , \59382 , \59383 , \59384 ,
         \59385 , \59386 , \59387 , \59388 , \59389 , \59390 , \59391 , \59392 , \59393 , \59394 ,
         \59395 , \59396 , \59397 , \59398 , \59399 , \59400 , \59401 , \59402 , \59403 , \59404 ,
         \59405 , \59406 , \59407 , \59408 , \59409 , \59410 , \59411 , \59412 , \59413 , \59414 ,
         \59415 , \59416 , \59417 , \59418 , \59419 , \59420 , \59421 , \59422 , \59423 , \59424 ,
         \59425 , \59426 , \59427 , \59428 , \59429 , \59430 , \59431 , \59432 , \59433 , \59434 ,
         \59435 , \59436 , \59437 , \59438 , \59439 , \59440 , \59441 , \59442 , \59443 , \59444 ,
         \59445 , \59446 , \59447 , \59448 , \59449 , \59450 , \59451 , \59452 , \59453 , \59454 ,
         \59455 , \59456 , \59457 , \59458 , \59459 , \59460 , \59461 , \59462 , \59463 , \59464 ,
         \59465 , \59466 , \59467 , \59468 , \59469 , \59470 , \59471 , \59472 , \59473 , \59474 ,
         \59475 , \59476 , \59477 , \59478 , \59479 , \59480 , \59481 , \59482 , \59483 , \59484 ,
         \59485 , \59486 , \59487 , \59488 , \59489 , \59490 , \59491 , \59492 , \59493 , \59494 ,
         \59495 , \59496 , \59497 , \59498 , \59499 , \59500 , \59501 , \59502 , \59503 , \59504 ,
         \59505 , \59506 , \59507 , \59508 , \59509 , \59510 , \59511 , \59512 , \59513 , \59514 ,
         \59515 , \59516 , \59517 , \59518 , \59519 , \59520 , \59521 , \59522 , \59523 , \59524 ,
         \59525 , \59526 , \59527 , \59528 , \59529 , \59530 , \59531 , \59532 , \59533 , \59534 ,
         \59535 , \59536 , \59537 , \59538 , \59539 , \59540 , \59541 , \59542 , \59543 , \59544 ,
         \59545 , \59546 , \59547 , \59548 , \59549 , \59550 , \59551 , \59552 , \59553 , \59554 ,
         \59555 , \59556 , \59557 , \59558 , \59559 , \59560 , \59561 , \59562 , \59563 , \59564 ,
         \59565 , \59566 , \59567 , \59568 , \59569 , \59570 , \59571 , \59572 , \59573 , \59574 ,
         \59575 , \59576 , \59577 , \59578 , \59579 , \59580 , \59581 , \59582 , \59583 , \59584 ,
         \59585 , \59586 , \59587 , \59588 , \59589 , \59590 , \59591 , \59592 , \59593 , \59594 ,
         \59595 , \59596 , \59597 , \59598 , \59599 , \59600 , \59601 , \59602 , \59603 , \59604 ,
         \59605 , \59606 , \59607 , \59608 , \59609 , \59610 , \59611 , \59612 , \59613 , \59614 ,
         \59615 , \59616 , \59617 , \59618 , \59619 , \59620 , \59621 , \59622 , \59623 , \59624 ,
         \59625 , \59626 , \59627 , \59628 , \59629 , \59630 , \59631 , \59632 , \59633 , \59634 ,
         \59635 , \59636 , \59637 , \59638 , \59639 , \59640 , \59641 , \59642 , \59643 , \59644 ,
         \59645 , \59646 , \59647 , \59648 , \59649 , \59650 , \59651 , \59652 , \59653 , \59654 ,
         \59655 , \59656 , \59657 , \59658 , \59659 , \59660 , \59661 , \59662 , \59663 , \59664 ,
         \59665 , \59666 , \59667 , \59668 , \59669 , \59670 , \59671 , \59672 , \59673 , \59674 ,
         \59675 , \59676 , \59677 , \59678 , \59679 , \59680 , \59681 , \59682 , \59683 , \59684 ,
         \59685 , \59686 , \59687 , \59688 , \59689 , \59690 , \59691 , \59692 , \59693 , \59694 ,
         \59695 , \59696 , \59697 , \59698 , \59699 , \59700 , \59701 , \59702 , \59703 , \59704 ,
         \59705 , \59706 , \59707 , \59708 , \59709 , \59710 , \59711 , \59712 , \59713 , \59714 ,
         \59715 , \59716 , \59717 , \59718 , \59719 , \59720 , \59721 , \59722 , \59723 , \59724 ,
         \59725 , \59726 , \59727 , \59728 , \59729 , \59730 , \59731 , \59732 , \59733 , \59734 ,
         \59735 , \59736 , \59737 , \59738 , \59739 , \59740 , \59741 , \59742 , \59743 , \59744 ,
         \59745 , \59746 , \59747 , \59748 , \59749 , \59750 , \59751 , \59752 , \59753 , \59754 ,
         \59755 , \59756 , \59757 , \59758 , \59759 , \59760 , \59761 , \59762 , \59763 , \59764 ,
         \59765 , \59766 , \59767 , \59768 , \59769 , \59770 , \59771 , \59772 , \59773 , \59774 ,
         \59775 , \59776 , \59777 , \59778 , \59779 , \59780 , \59781 , \59782 , \59783 , \59784 ,
         \59785 , \59786 , \59787 , \59788 , \59789 , \59790 , \59791 , \59792 , \59793 , \59794 ,
         \59795 , \59796 , \59797 , \59798 , \59799 , \59800 , \59801 , \59802 , \59803 , \59804 ,
         \59805 , \59806 , \59807 , \59808 , \59809 , \59810 , \59811 , \59812 , \59813 , \59814 ,
         \59815 , \59816 , \59817 , \59818 , \59819 , \59820 , \59821 , \59822 , \59823 , \59824 ,
         \59825 , \59826 , \59827 , \59828 , \59829 , \59830 , \59831 , \59832 , \59833 , \59834 ,
         \59835 , \59836 , \59837 , \59838 , \59839 , \59840 , \59841 , \59842 , \59843 , \59844 ,
         \59845 , \59846 , \59847 , \59848 , \59849 , \59850 , \59851 , \59852 , \59853 , \59854 ,
         \59855 , \59856 , \59857 , \59858 , \59859 , \59860 , \59861 , \59862 , \59863 , \59864 ,
         \59865 , \59866 , \59867 , \59868 , \59869 , \59870 , \59871 , \59872 , \59873 , \59874 ,
         \59875 , \59876 , \59877 , \59878 , \59879 , \59880 , \59881 , \59882 , \59883 , \59884 ,
         \59885 , \59886 , \59887 , \59888 , \59889 , \59890 , \59891 , \59892 , \59893 , \59894 ,
         \59895 , \59896 , \59897 , \59898 , \59899 , \59900 , \59901 , \59902 , \59903 , \59904 ,
         \59905 , \59906 , \59907 , \59908 , \59909 , \59910 , \59911 , \59912 , \59913 , \59914 ,
         \59915 , \59916 , \59917 , \59918 , \59919 , \59920 , \59921 , \59922 , \59923 , \59924 ,
         \59925 , \59926 , \59927 , \59928 , \59929 , \59930 , \59931 , \59932 , \59933 , \59934 ,
         \59935 , \59936 , \59937 , \59938 , \59939 , \59940 , \59941 , \59942 , \59943 , \59944 ,
         \59945 , \59946 , \59947 , \59948 , \59949 , \59950 , \59951 , \59952 , \59953 , \59954 ,
         \59955 , \59956 , \59957 , \59958 , \59959 , \59960 , \59961 , \59962 , \59963 , \59964 ,
         \59965 , \59966 , \59967 , \59968 , \59969 , \59970 , \59971 , \59972 , \59973 , \59974 ,
         \59975 , \59976 , \59977 , \59978 , \59979 , \59980 , \59981 , \59982 , \59983 , \59984 ,
         \59985 , \59986 , \59987 , \59988 , \59989 , \59990 , \59991 , \59992 , \59993 , \59994 ,
         \59995 , \59996 , \59997 , \59998 , \59999 , \60000 , \60001 , \60002 , \60003 , \60004 ,
         \60005 , \60006 , \60007 , \60008 , \60009 , \60010 , \60011 , \60012 , \60013 , \60014 ,
         \60015 , \60016 , \60017 , \60018 , \60019 , \60020 , \60021 , \60022 , \60023 , \60024 ,
         \60025 , \60026 , \60027 , \60028 , \60029 , \60030 , \60031 , \60032 , \60033 , \60034 ,
         \60035 , \60036 , \60037 , \60038 , \60039 , \60040 , \60041 , \60042 , \60043 , \60044 ,
         \60045 , \60046 , \60047 , \60048 , \60049 , \60050 , \60051 , \60052 , \60053 , \60054 ,
         \60055 , \60056 , \60057 , \60058 , \60059 , \60060 , \60061 , \60062 , \60063 , \60064 ,
         \60065 , \60066 , \60067 , \60068 , \60069 , \60070 , \60071 , \60072 , \60073 , \60074 ,
         \60075 , \60076 , \60077 , \60078 , \60079 , \60080 , \60081 , \60082 , \60083 , \60084 ,
         \60085 , \60086 , \60087 , \60088 , \60089 , \60090 , \60091 , \60092 , \60093 , \60094 ,
         \60095 , \60096 , \60097 , \60098 , \60099 , \60100 , \60101 , \60102 , \60103 , \60104 ,
         \60105 , \60106 , \60107 , \60108 , \60109 , \60110 , \60111 , \60112 , \60113 , \60114 ,
         \60115 , \60116 , \60117 , \60118 , \60119 , \60120 , \60121 , \60122 , \60123 , \60124 ,
         \60125 , \60126 , \60127 , \60128 , \60129 , \60130 , \60131 , \60132 , \60133 , \60134 ,
         \60135 , \60136 , \60137 , \60138 , \60139 , \60140 , \60141 , \60142 , \60143 , \60144 ,
         \60145 , \60146 , \60147 , \60148 , \60149 , \60150 , \60151 , \60152 , \60153 , \60154 ,
         \60155 , \60156 , \60157 , \60158 , \60159 , \60160 , \60161 , \60162 , \60163 , \60164 ,
         \60165 , \60166 , \60167 , \60168 , \60169 , \60170 , \60171 , \60172 , \60173 , \60174 ,
         \60175 , \60176 , \60177 , \60178 , \60179 , \60180 , \60181 , \60182 , \60183 , \60184 ,
         \60185 , \60186 , \60187 , \60188 , \60189 , \60190 , \60191 , \60192 , \60193 , \60194 ,
         \60195 , \60196 , \60197 , \60198 , \60199 , \60200 , \60201 , \60202 , \60203 , \60204 ,
         \60205 , \60206 , \60207 , \60208 , \60209 , \60210 , \60211 , \60212 , \60213 , \60214 ,
         \60215 , \60216 , \60217 , \60218 , \60219 , \60220 , \60221 , \60222 , \60223 , \60224 ,
         \60225 , \60226 , \60227 , \60228 , \60229 , \60230 , \60231 , \60232 , \60233 , \60234 ,
         \60235 , \60236 , \60237 , \60238 , \60239 , \60240 , \60241 , \60242 , \60243 , \60244 ,
         \60245 , \60246 , \60247 , \60248 , \60249 , \60250 , \60251 , \60252 , \60253 , \60254 ,
         \60255 , \60256 , \60257 , \60258 , \60259 , \60260 , \60261 , \60262 , \60263 , \60264 ,
         \60265 , \60266 , \60267 , \60268 , \60269 , \60270 , \60271 , \60272 , \60273 , \60274 ,
         \60275 , \60276 , \60277 , \60278 , \60279 , \60280 , \60281 , \60282 , \60283 , \60284 ,
         \60285 , \60286 , \60287 , \60288 , \60289 , \60290 , \60291 , \60292 , \60293 , \60294 ,
         \60295 , \60296 , \60297 , \60298 , \60299 , \60300 , \60301 , \60302 , \60303 , \60304 ,
         \60305 , \60306 , \60307 , \60308 , \60309 , \60310 , \60311 , \60312 , \60313 , \60314 ,
         \60315 , \60316 , \60317 , \60318 , \60319 , \60320 , \60321 , \60322 , \60323 , \60324 ,
         \60325 , \60326 , \60327 , \60328 , \60329 , \60330 , \60331 , \60332 , \60333 , \60334 ,
         \60335 , \60336 , \60337 , \60338 , \60339 , \60340 , \60341 , \60342 , \60343 , \60344 ,
         \60345 , \60346 , \60347 , \60348 , \60349 , \60350 , \60351 , \60352 , \60353 , \60354 ,
         \60355 , \60356 , \60357 , \60358 , \60359 , \60360 , \60361 , \60362 , \60363 , \60364 ,
         \60365 , \60366 , \60367 , \60368 , \60369 , \60370 , \60371 , \60372 , \60373 , \60374 ,
         \60375 , \60376 , \60377 , \60378 , \60379 , \60380 , \60381 , \60382 , \60383 , \60384 ,
         \60385 , \60386 , \60387 , \60388 , \60389 , \60390 , \60391 , \60392 , \60393 , \60394 ,
         \60395 , \60396 , \60397 , \60398 , \60399 , \60400 , \60401 , \60402 , \60403 , \60404 ,
         \60405 , \60406 , \60407 , \60408 , \60409 , \60410 , \60411 , \60412 , \60413 , \60414 ,
         \60415 , \60416 , \60417 , \60418 , \60419 , \60420 , \60421 , \60422 , \60423 , \60424 ,
         \60425 , \60426 , \60427 , \60428 , \60429 , \60430 , \60431 , \60432 , \60433 , \60434 ,
         \60435 , \60436 , \60437 , \60438 , \60439 , \60440 , \60441 , \60442 , \60443 , \60444 ,
         \60445 , \60446 , \60447 , \60448 , \60449 , \60450 , \60451 , \60452 , \60453 , \60454 ,
         \60455 , \60456 , \60457 , \60458 , \60459 , \60460 , \60461 , \60462 , \60463 , \60464 ,
         \60465 , \60466 , \60467 , \60468 , \60469 , \60470 , \60471 , \60472 , \60473 , \60474 ,
         \60475 , \60476 , \60477 , \60478 , \60479 , \60480 , \60481 , \60482 , \60483 , \60484 ,
         \60485 , \60486 , \60487 , \60488 , \60489 , \60490 , \60491 , \60492 , \60493 , \60494 ,
         \60495 , \60496 , \60497 , \60498 , \60499 , \60500 , \60501 , \60502 , \60503 , \60504 ,
         \60505 , \60506 , \60507 , \60508 , \60509 , \60510 , \60511 , \60512 , \60513 , \60514 ,
         \60515 , \60516 , \60517 , \60518 , \60519 , \60520 , \60521 , \60522 , \60523 , \60524 ,
         \60525 , \60526 , \60527 , \60528 , \60529 , \60530 , \60531 , \60532 , \60533 , \60534 ,
         \60535 , \60536 , \60537 , \60538 , \60539 , \60540 , \60541 , \60542 , \60543 , \60544 ,
         \60545 , \60546 , \60547 , \60548 , \60549 , \60550 , \60551 , \60552 , \60553 , \60554 ,
         \60555 , \60556 , \60557 , \60558 , \60559 , \60560 , \60561 , \60562 , \60563 , \60564 ,
         \60565 , \60566 , \60567 , \60568 , \60569 , \60570 , \60571 , \60572 , \60573 , \60574 ,
         \60575 , \60576 , \60577 , \60578 , \60579 , \60580 , \60581 , \60582 , \60583 , \60584 ,
         \60585 , \60586 , \60587 , \60588 , \60589 , \60590 , \60591 , \60592 , \60593 , \60594 ,
         \60595 , \60596 , \60597 , \60598 , \60599 , \60600 , \60601 , \60602 , \60603 , \60604 ,
         \60605 , \60606 , \60607 , \60608 , \60609 , \60610 , \60611 , \60612 , \60613 , \60614 ,
         \60615 , \60616 , \60617 , \60618 , \60619 , \60620 , \60621 , \60622 , \60623 , \60624 ,
         \60625 , \60626 , \60627 , \60628 , \60629 , \60630 , \60631 , \60632 , \60633 , \60634 ,
         \60635 , \60636 , \60637 , \60638 , \60639 , \60640 , \60641 , \60642 , \60643 , \60644 ,
         \60645 , \60646 , \60647 , \60648 , \60649 , \60650 , \60651 , \60652 , \60653 , \60654 ,
         \60655 , \60656 , \60657 , \60658 , \60659 , \60660 , \60661 , \60662 , \60663 , \60664 ,
         \60665 , \60666 , \60667 , \60668 , \60669 , \60670 , \60671 , \60672 , \60673 , \60674 ,
         \60675 , \60676 , \60677 , \60678 , \60679 , \60680 , \60681 , \60682 , \60683 , \60684 ,
         \60685 , \60686 , \60687 , \60688 , \60689 , \60690 , \60691 , \60692 , \60693 , \60694 ,
         \60695 , \60696 , \60697 , \60698 , \60699 , \60700 , \60701 , \60702 , \60703 , \60704 ,
         \60705 , \60706 , \60707 , \60708 , \60709 , \60710 , \60711 , \60712 , \60713 , \60714 ,
         \60715 , \60716 , \60717 , \60718 , \60719 , \60720 , \60721 , \60722 , \60723 , \60724 ,
         \60725 , \60726 , \60727 , \60728 , \60729 , \60730 , \60731 , \60732 , \60733 , \60734 ,
         \60735 , \60736 , \60737 , \60738 , \60739 , \60740 , \60741 , \60742 , \60743 , \60744 ,
         \60745 , \60746 , \60747 , \60748 , \60749 , \60750 , \60751 , \60752 , \60753 , \60754 ,
         \60755 , \60756 , \60757 , \60758 , \60759 , \60760 , \60761 , \60762 , \60763 , \60764 ,
         \60765 , \60766 , \60767 , \60768 , \60769 , \60770 , \60771 , \60772 , \60773 , \60774 ,
         \60775 , \60776 , \60777 , \60778 , \60779 , \60780 , \60781 , \60782 , \60783 , \60784 ,
         \60785 , \60786 , \60787 , \60788 , \60789 , \60790 , \60791 , \60792 , \60793 , \60794 ,
         \60795 , \60796 , \60797 , \60798 , \60799 , \60800 , \60801 , \60802 , \60803 , \60804 ,
         \60805 , \60806 , \60807 , \60808 , \60809 , \60810 , \60811 , \60812 , \60813 , \60814 ,
         \60815 , \60816 , \60817 , \60818 , \60819 , \60820 , \60821 , \60822 , \60823 , \60824 ,
         \60825 , \60826 , \60827 , \60828 , \60829 , \60830 , \60831 , \60832 , \60833 , \60834 ,
         \60835 , \60836 , \60837 , \60838 , \60839 , \60840 , \60841 , \60842 , \60843 , \60844 ,
         \60845 , \60846 , \60847 , \60848 , \60849 , \60850 , \60851 , \60852 , \60853 , \60854 ,
         \60855 , \60856 , \60857 , \60858 , \60859 , \60860 , \60861 , \60862 , \60863 , \60864 ,
         \60865 , \60866 , \60867 , \60868 , \60869 , \60870 , \60871 , \60872 , \60873 , \60874 ,
         \60875 , \60876 , \60877 , \60878 , \60879 , \60880 , \60881 , \60882 , \60883 , \60884 ,
         \60885 , \60886 , \60887 , \60888 , \60889 , \60890 , \60891 , \60892 , \60893 , \60894 ,
         \60895 , \60896 , \60897 , \60898 , \60899 , \60900 , \60901 , \60902 , \60903 , \60904 ,
         \60905 , \60906 , \60907 , \60908 , \60909 , \60910 , \60911 , \60912 , \60913 , \60914 ,
         \60915 , \60916 , \60917 , \60918 , \60919 , \60920 , \60921 , \60922 , \60923 , \60924 ,
         \60925 , \60926 , \60927 , \60928 , \60929 , \60930 , \60931 , \60932 , \60933 , \60934 ,
         \60935 , \60936 , \60937 , \60938 , \60939 , \60940 , \60941 , \60942 , \60943 , \60944 ,
         \60945 , \60946 , \60947 , \60948 , \60949 , \60950 , \60951 , \60952 , \60953 , \60954 ,
         \60955 , \60956 , \60957 , \60958 , \60959 , \60960 , \60961 , \60962 , \60963 , \60964 ,
         \60965 , \60966 , \60967 , \60968 , \60969 , \60970 , \60971 , \60972 , \60973 , \60974 ,
         \60975 , \60976 , \60977 , \60978 , \60979 , \60980 , \60981 , \60982 , \60983 , \60984 ,
         \60985 , \60986 , \60987 , \60988 , \60989 , \60990 , \60991 , \60992 , \60993 , \60994 ,
         \60995 , \60996 , \60997 , \60998 , \60999 , \61000 , \61001 , \61002 , \61003 , \61004 ,
         \61005 , \61006 , \61007 , \61008 , \61009 , \61010 , \61011 , \61012 , \61013 , \61014 ,
         \61015 , \61016 , \61017 , \61018 , \61019 , \61020 , \61021 , \61022 , \61023 , \61024 ,
         \61025 , \61026 , \61027 , \61028 , \61029 , \61030 , \61031 , \61032 , \61033 , \61034 ,
         \61035 , \61036 , \61037 , \61038 , \61039 , \61040 , \61041 , \61042 , \61043 , \61044 ,
         \61045 , \61046 , \61047 , \61048 , \61049 , \61050 , \61051 , \61052 , \61053 , \61054 ,
         \61055 , \61056 , \61057 , \61058 , \61059 , \61060 , \61061 , \61062 , \61063 , \61064 ,
         \61065 , \61066 , \61067 , \61068 , \61069 , \61070 , \61071 , \61072 , \61073 , \61074 ,
         \61075 , \61076 , \61077 , \61078 , \61079 , \61080 , \61081 , \61082 , \61083 , \61084 ,
         \61085 , \61086 , \61087 , \61088 , \61089 , \61090 , \61091 , \61092 , \61093 , \61094 ,
         \61095 , \61096 , \61097 , \61098 , \61099 , \61100 , \61101 , \61102 , \61103 , \61104 ,
         \61105 , \61106 , \61107 , \61108 , \61109 , \61110 , \61111 , \61112 , \61113 , \61114 ,
         \61115 , \61116 , \61117 , \61118 , \61119 , \61120 , \61121 , \61122 , \61123 , \61124 ,
         \61125 , \61126 , \61127 , \61128 , \61129 , \61130 , \61131 , \61132 , \61133 , \61134 ,
         \61135 , \61136 , \61137 , \61138 , \61139 , \61140 , \61141 , \61142 , \61143 , \61144 ,
         \61145 , \61146 , \61147 , \61148 , \61149 , \61150 , \61151 , \61152 , \61153 , \61154 ,
         \61155 , \61156 , \61157 , \61158 , \61159 , \61160 , \61161 , \61162 , \61163 , \61164 ,
         \61165 , \61166 , \61167 , \61168 , \61169 , \61170 , \61171 , \61172 , \61173 , \61174 ,
         \61175 , \61176 , \61177 , \61178 , \61179 , \61180 , \61181 , \61182 , \61183 , \61184 ,
         \61185 , \61186 , \61187 , \61188 , \61189 , \61190 , \61191 , \61192 , \61193 , \61194 ,
         \61195 , \61196 , \61197 , \61198 , \61199 , \61200 , \61201 , \61202 , \61203 , \61204 ,
         \61205 , \61206 , \61207 , \61208 , \61209 , \61210 , \61211 , \61212 , \61213 , \61214 ,
         \61215 , \61216 , \61217 , \61218 , \61219 , \61220 , \61221 , \61222 , \61223 , \61224 ,
         \61225 , \61226 , \61227 , \61228 , \61229 , \61230 , \61231 , \61232 , \61233 , \61234 ,
         \61235 , \61236 , \61237 , \61238 , \61239 , \61240 , \61241 , \61242 , \61243 , \61244 ,
         \61245 , \61246 , \61247 , \61248 , \61249 , \61250 , \61251 , \61252 , \61253 , \61254 ,
         \61255 , \61256 , \61257 , \61258 , \61259 , \61260 , \61261 , \61262 , \61263 , \61264 ,
         \61265 , \61266 , \61267 , \61268 , \61269 , \61270 , \61271 , \61272 , \61273 , \61274 ,
         \61275 , \61276 , \61277 , \61278 , \61279 , \61280 , \61281 , \61282 , \61283 , \61284 ,
         \61285 , \61286 , \61287 , \61288 , \61289 , \61290 , \61291 , \61292 , \61293 , \61294 ,
         \61295 , \61296 , \61297 , \61298 , \61299 , \61300 , \61301 , \61302 , \61303 , \61304 ,
         \61305 , \61306 , \61307 , \61308 , \61309 , \61310 , \61311 , \61312 , \61313 , \61314 ,
         \61315 , \61316 , \61317 , \61318 , \61319 , \61320 , \61321 , \61322 , \61323 , \61324 ,
         \61325 , \61326 , \61327 , \61328 , \61329 , \61330 , \61331 , \61332 , \61333 , \61334 ,
         \61335 , \61336 , \61337 , \61338 , \61339 , \61340 , \61341 , \61342 , \61343 , \61344 ,
         \61345 , \61346 , \61347 , \61348 , \61349 , \61350 , \61351 , \61352 , \61353 , \61354 ,
         \61355 , \61356 , \61357 , \61358 , \61359 , \61360 , \61361 , \61362 , \61363 , \61364 ,
         \61365 , \61366 , \61367 , \61368 , \61369 , \61370 , \61371 , \61372 , \61373 , \61374 ,
         \61375 , \61376 , \61377 , \61378 , \61379 , \61380 , \61381 , \61382 , \61383 , \61384 ,
         \61385 , \61386 , \61387 , \61388 , \61389 , \61390 , \61391 , \61392 , \61393 , \61394 ,
         \61395 , \61396 , \61397 , \61398 , \61399 , \61400 , \61401 , \61402 , \61403 , \61404 ,
         \61405 , \61406 , \61407 , \61408 , \61409 , \61410 , \61411 , \61412 , \61413 , \61414 ,
         \61415 , \61416 , \61417 , \61418 , \61419 , \61420 , \61421 , \61422 , \61423 , \61424 ,
         \61425 , \61426 , \61427 , \61428 , \61429 , \61430 , \61431 , \61432 , \61433 , \61434 ,
         \61435 , \61436 , \61437 , \61438 , \61439 , \61440 , \61441 , \61442 , \61443 , \61444 ,
         \61445 , \61446 , \61447 , \61448 , \61449 , \61450 , \61451 , \61452 , \61453 , \61454 ,
         \61455 , \61456 , \61457 , \61458 , \61459 , \61460 , \61461 , \61462 , \61463 , \61464 ,
         \61465 , \61466 , \61467 , \61468 , \61469 , \61470 , \61471 , \61472 , \61473 , \61474 ,
         \61475 , \61476 , \61477 , \61478 , \61479 , \61480 , \61481 , \61482 , \61483 , \61484 ,
         \61485 , \61486 , \61487 , \61488 , \61489 , \61490 , \61491 , \61492 , \61493 , \61494 ,
         \61495 , \61496 , \61497 , \61498 , \61499 , \61500 , \61501 , \61502 , \61503 , \61504 ,
         \61505 , \61506 , \61507 , \61508 , \61509 , \61510 , \61511 , \61512 , \61513 , \61514 ,
         \61515 , \61516 , \61517 , \61518 , \61519 , \61520 , \61521 , \61522 , \61523 , \61524 ,
         \61525 , \61526 , \61527 , \61528 , \61529 , \61530 , \61531 , \61532 , \61533 , \61534 ,
         \61535 , \61536 , \61537 , \61538 , \61539 , \61540 , \61541 , \61542 , \61543 , \61544 ,
         \61545 , \61546 , \61547 , \61548 , \61549 , \61550 , \61551 , \61552 , \61553 , \61554 ,
         \61555 , \61556 , \61557 , \61558 , \61559 , \61560 , \61561 , \61562 , \61563 , \61564 ,
         \61565 , \61566 , \61567 , \61568 , \61569 , \61570 , \61571 , \61572 , \61573 , \61574 ,
         \61575 , \61576 , \61577 , \61578 , \61579 , \61580 , \61581 , \61582 , \61583 , \61584 ,
         \61585 , \61586 , \61587 , \61588 , \61589 , \61590 , \61591 , \61592 , \61593 , \61594 ,
         \61595 , \61596 , \61597 , \61598 , \61599 , \61600 , \61601 , \61602 , \61603 , \61604 ,
         \61605 , \61606 , \61607 , \61608 , \61609 , \61610 , \61611 , \61612 , \61613 , \61614 ,
         \61615 , \61616 , \61617 , \61618 , \61619 , \61620 , \61621 , \61622 , \61623 , \61624 ,
         \61625 , \61626 , \61627 , \61628 , \61629 , \61630 , \61631 , \61632 , \61633 , \61634 ,
         \61635 , \61636 , \61637 , \61638 , \61639 , \61640 , \61641 , \61642 , \61643 , \61644 ,
         \61645 , \61646 , \61647 , \61648 , \61649 , \61650 , \61651 , \61652 , \61653 , \61654 ,
         \61655 , \61656 , \61657 , \61658 , \61659 , \61660 , \61661 , \61662 , \61663 , \61664 ,
         \61665 , \61666 , \61667 , \61668 , \61669 , \61670 , \61671 , \61672 , \61673 , \61674 ,
         \61675 , \61676 , \61677 , \61678 , \61679 , \61680 , \61681 , \61682 , \61683 , \61684 ,
         \61685 , \61686 , \61687 , \61688 , \61689 , \61690 , \61691 , \61692 , \61693 , \61694 ,
         \61695 , \61696 , \61697 , \61698 , \61699 , \61700 , \61701 , \61702 , \61703 , \61704 ,
         \61705 , \61706 , \61707 , \61708 , \61709 , \61710 , \61711 , \61712 , \61713 , \61714 ,
         \61715 , \61716 , \61717 , \61718 , \61719 , \61720 , \61721 , \61722 , \61723 , \61724 ,
         \61725 , \61726 , \61727 , \61728 , \61729 , \61730 , \61731 , \61732 , \61733 , \61734 ,
         \61735 , \61736 , \61737 , \61738 , \61739 , \61740 , \61741 , \61742 , \61743 , \61744 ,
         \61745 , \61746 , \61747 , \61748 , \61749 , \61750 , \61751 , \61752 , \61753 , \61754 ,
         \61755 , \61756 , \61757 , \61758 , \61759 , \61760 , \61761 , \61762 , \61763 , \61764 ,
         \61765 , \61766 , \61767 , \61768 , \61769 , \61770 , \61771 , \61772 , \61773 , \61774 ,
         \61775 , \61776 , \61777 , \61778 , \61779 , \61780 , \61781 , \61782 , \61783 , \61784 ,
         \61785 , \61786 , \61787 , \61788 , \61789 , \61790 , \61791 , \61792 , \61793 , \61794 ,
         \61795 , \61796 , \61797 , \61798 , \61799 , \61800 , \61801 , \61802 , \61803 , \61804 ,
         \61805 , \61806 , \61807 , \61808 , \61809 , \61810 , \61811 , \61812 , \61813 , \61814 ,
         \61815 , \61816 , \61817 , \61818 , \61819 , \61820 , \61821 , \61822 , \61823 , \61824 ,
         \61825 , \61826 , \61827 , \61828 , \61829 , \61830 , \61831 , \61832 , \61833 , \61834 ,
         \61835 , \61836 , \61837 , \61838 , \61839 , \61840 , \61841 , \61842 , \61843 , \61844 ,
         \61845 , \61846 , \61847 , \61848 , \61849 , \61850 , \61851 , \61852 , \61853 , \61854 ,
         \61855 , \61856 , \61857 , \61858 , \61859 , \61860 , \61861 , \61862 , \61863 , \61864 ,
         \61865 , \61866 , \61867 , \61868 , \61869 , \61870 , \61871 , \61872 , \61873 , \61874 ,
         \61875 , \61876 , \61877 , \61878 , \61879 , \61880 , \61881 , \61882 , \61883 , \61884 ,
         \61885 , \61886 , \61887 , \61888 , \61889 , \61890 , \61891 , \61892 , \61893 , \61894 ,
         \61895 , \61896 , \61897 , \61898 , \61899 , \61900 , \61901 , \61902 , \61903 , \61904 ,
         \61905 , \61906 , \61907 , \61908 , \61909 , \61910 , \61911 , \61912 , \61913 , \61914 ,
         \61915 , \61916 , \61917 , \61918 , \61919 , \61920 , \61921 , \61922 , \61923 , \61924 ,
         \61925 , \61926 , \61927 , \61928 , \61929 , \61930 , \61931 , \61932 , \61933 , \61934 ,
         \61935 , \61936 , \61937 , \61938 , \61939 , \61940 , \61941 , \61942 , \61943 , \61944 ,
         \61945 , \61946 , \61947 , \61948 , \61949 , \61950 , \61951 , \61952 , \61953 , \61954 ,
         \61955 , \61956 , \61957 , \61958 , \61959 , \61960 , \61961 , \61962 , \61963 , \61964 ,
         \61965 , \61966 , \61967 , \61968 , \61969 , \61970 , \61971 , \61972 , \61973 , \61974 ,
         \61975 , \61976 , \61977 , \61978 , \61979 , \61980 , \61981 , \61982 , \61983 , \61984 ,
         \61985 , \61986 , \61987 , \61988 , \61989 , \61990 , \61991 , \61992 , \61993 , \61994 ,
         \61995 , \61996 , \61997 , \61998 , \61999 , \62000 , \62001 , \62002 , \62003 , \62004 ,
         \62005 , \62006 , \62007 , \62008 , \62009 , \62010 , \62011 , \62012 , \62013 , \62014 ,
         \62015 , \62016 , \62017 , \62018 , \62019 , \62020 , \62021 , \62022 , \62023 , \62024 ,
         \62025 , \62026 , \62027 , \62028 , \62029 , \62030 , \62031 , \62032 , \62033 , \62034 ,
         \62035 , \62036 , \62037 , \62038 , \62039 , \62040 , \62041 , \62042 , \62043 , \62044 ,
         \62045 , \62046 , \62047 , \62048 , \62049 , \62050 , \62051 , \62052 , \62053 , \62054 ,
         \62055 , \62056 , \62057 , \62058 , \62059 , \62060 , \62061 , \62062 , \62063 , \62064 ,
         \62065 , \62066 , \62067 , \62068 , \62069 , \62070 , \62071 , \62072 , \62073 , \62074 ,
         \62075 , \62076 , \62077 , \62078 , \62079 , \62080 , \62081 , \62082 , \62083 , \62084 ,
         \62085 , \62086 , \62087 , \62088 , \62089 , \62090 , \62091 , \62092 , \62093 , \62094 ,
         \62095 , \62096 , \62097 , \62098 , \62099 , \62100 , \62101 , \62102 , \62103 , \62104 ,
         \62105 , \62106 , \62107 , \62108 , \62109 , \62110 , \62111 , \62112 , \62113 , \62114 ,
         \62115 , \62116 , \62117 , \62118 , \62119 , \62120 , \62121 , \62122 , \62123 , \62124 ,
         \62125 , \62126 , \62127 , \62128 , \62129 , \62130 , \62131 , \62132 , \62133 , \62134 ,
         \62135 , \62136 , \62137 , \62138 , \62139 , \62140 , \62141 , \62142 , \62143 , \62144 ,
         \62145 , \62146 , \62147 , \62148 , \62149 , \62150 , \62151 , \62152 , \62153 , \62154 ,
         \62155 , \62156 , \62157 , \62158 , \62159 , \62160 , \62161 , \62162 , \62163 , \62164 ,
         \62165 , \62166 , \62167 , \62168 , \62169 , \62170 , \62171 , \62172 , \62173 , \62174 ,
         \62175 , \62176 , \62177 , \62178 , \62179 , \62180 , \62181 , \62182 , \62183 , \62184 ,
         \62185 , \62186 , \62187 , \62188 , \62189 , \62190 , \62191 , \62192 , \62193 , \62194 ,
         \62195 , \62196 , \62197 , \62198 , \62199 , \62200 , \62201 , \62202 , \62203 , \62204 ,
         \62205 , \62206 , \62207 , \62208 , \62209 , \62210 , \62211 , \62212 , \62213 , \62214 ,
         \62215 , \62216 , \62217 , \62218 , \62219 , \62220 , \62221 , \62222 , \62223 , \62224 ,
         \62225 , \62226 , \62227 , \62228 , \62229 , \62230 , \62231 , \62232 , \62233 , \62234 ,
         \62235 , \62236 , \62237 , \62238 , \62239 , \62240 , \62241 , \62242 , \62243 , \62244 ,
         \62245 , \62246 , \62247 , \62248 , \62249 , \62250 , \62251 , \62252 , \62253 , \62254 ,
         \62255 , \62256 , \62257 , \62258 , \62259 , \62260 , \62261 , \62262 , \62263 , \62264 ,
         \62265 , \62266 , \62267 , \62268 , \62269 , \62270 , \62271 , \62272 , \62273 , \62274 ,
         \62275 , \62276 , \62277 , \62278 , \62279 , \62280 , \62281 , \62282 , \62283 , \62284 ,
         \62285 , \62286 , \62287 , \62288 , \62289 , \62290 , \62291 , \62292 , \62293 , \62294 ,
         \62295 , \62296 , \62297 , \62298 , \62299 , \62300 , \62301 , \62302 , \62303 , \62304 ,
         \62305 , \62306 , \62307 , \62308 , \62309 , \62310 , \62311 , \62312 , \62313 , \62314 ,
         \62315 , \62316 , \62317 , \62318 , \62319 , \62320 , \62321 , \62322 , \62323 , \62324 ,
         \62325 , \62326 , \62327 , \62328 , \62329 , \62330 , \62331 , \62332 , \62333 , \62334 ,
         \62335 , \62336 , \62337 , \62338 , \62339 , \62340 , \62341 , \62342 , \62343 , \62344 ,
         \62345 , \62346 , \62347 , \62348 , \62349 , \62350 , \62351 , \62352 , \62353 , \62354 ,
         \62355 , \62356 , \62357 , \62358 , \62359 , \62360 , \62361 , \62362 , \62363 , \62364 ,
         \62365 , \62366 , \62367 , \62368 , \62369 , \62370 , \62371 , \62372 , \62373 , \62374 ,
         \62375 , \62376 , \62377 , \62378 , \62379 , \62380 , \62381 , \62382 , \62383 , \62384 ,
         \62385 , \62386 , \62387 , \62388 , \62389 , \62390 , \62391 , \62392 , \62393 , \62394 ,
         \62395 , \62396 , \62397 , \62398 , \62399 , \62400 , \62401 , \62402 , \62403 , \62404 ,
         \62405 , \62406 , \62407 , \62408 , \62409 , \62410 , \62411 , \62412 , \62413 , \62414 ,
         \62415 , \62416 , \62417 , \62418 , \62419 , \62420 , \62421 , \62422 , \62423 , \62424 ,
         \62425 , \62426 , \62427 , \62428 , \62429 , \62430 , \62431 , \62432 , \62433 , \62434 ,
         \62435 , \62436 , \62437 , \62438 , \62439 , \62440 , \62441 , \62442 , \62443 , \62444 ,
         \62445 , \62446 , \62447 , \62448 , \62449 , \62450 , \62451 , \62452 , \62453 , \62454 ,
         \62455 , \62456 , \62457 , \62458 , \62459 , \62460 , \62461 , \62462 , \62463 , \62464 ,
         \62465 , \62466 , \62467 , \62468 , \62469 , \62470 , \62471 , \62472 , \62473 , \62474 ,
         \62475 , \62476 , \62477 , \62478 , \62479 , \62480 , \62481 , \62482 , \62483 , \62484 ,
         \62485 , \62486 , \62487 , \62488 , \62489 , \62490 , \62491 , \62492 , \62493 , \62494 ,
         \62495 , \62496 , \62497 , \62498 , \62499 , \62500 , \62501 , \62502 , \62503 , \62504 ,
         \62505 , \62506 , \62507 , \62508 , \62509 , \62510 , \62511 , \62512 , \62513 , \62514 ,
         \62515 , \62516 , \62517 , \62518 , \62519 , \62520 , \62521 , \62522 , \62523 , \62524 ,
         \62525 , \62526 , \62527 , \62528 , \62529 , \62530 , \62531 , \62532 , \62533 , \62534 ,
         \62535 , \62536 , \62537 , \62538 , \62539 , \62540 , \62541 , \62542 , \62543 , \62544 ,
         \62545 , \62546 , \62547 , \62548 , \62549 , \62550 , \62551 , \62552 , \62553 , \62554 ,
         \62555 , \62556 , \62557 , \62558 , \62559 , \62560 , \62561 , \62562 , \62563 , \62564 ,
         \62565 , \62566 , \62567 , \62568 , \62569 , \62570 , \62571 , \62572 , \62573 , \62574 ,
         \62575 , \62576 , \62577 , \62578 , \62579 , \62580 , \62581 , \62582 , \62583 , \62584 ,
         \62585 , \62586 , \62587 , \62588 , \62589 , \62590 , \62591 , \62592 , \62593 , \62594 ,
         \62595 , \62596 , \62597 , \62598 , \62599 , \62600 , \62601 , \62602 , \62603 , \62604 ,
         \62605 , \62606 , \62607 , \62608 , \62609 , \62610 , \62611 , \62612 , \62613 , \62614 ,
         \62615 , \62616 , \62617 , \62618 , \62619 , \62620 , \62621 , \62622 , \62623 , \62624 ,
         \62625 , \62626 , \62627 , \62628 , \62629 , \62630 , \62631 , \62632 , \62633 , \62634 ,
         \62635 , \62636 , \62637 , \62638 , \62639 , \62640 , \62641 , \62642 , \62643 , \62644 ,
         \62645 , \62646 , \62647 , \62648 , \62649 , \62650 , \62651 , \62652 , \62653 , \62654 ,
         \62655 , \62656 , \62657 , \62658 , \62659 , \62660 , \62661 , \62662 , \62663 , \62664 ,
         \62665 , \62666 , \62667 , \62668 , \62669 , \62670 , \62671 , \62672 , \62673 , \62674 ,
         \62675 , \62676 , \62677 , \62678 , \62679 , \62680 , \62681 , \62682 , \62683 , \62684 ,
         \62685 , \62686 , \62687 , \62688 , \62689 , \62690 , \62691 , \62692 , \62693 , \62694 ,
         \62695 , \62696 , \62697 , \62698 , \62699 , \62700 , \62701 , \62702 , \62703 , \62704 ,
         \62705 , \62706 , \62707 , \62708 , \62709 , \62710 , \62711 , \62712 , \62713 , \62714 ,
         \62715 , \62716 , \62717 , \62718 , \62719 , \62720 , \62721 , \62722 , \62723 , \62724 ,
         \62725 , \62726 , \62727 , \62728 , \62729 , \62730 , \62731 , \62732 , \62733 , \62734 ,
         \62735 , \62736 , \62737 , \62738 , \62739 , \62740 , \62741 , \62742 , \62743 , \62744 ,
         \62745 , \62746 , \62747 , \62748 , \62749 , \62750 , \62751 , \62752 , \62753 , \62754 ,
         \62755 , \62756 , \62757 , \62758 , \62759 , \62760 , \62761 , \62762 , \62763 , \62764 ,
         \62765 , \62766 , \62767 , \62768 , \62769 , \62770 , \62771 , \62772 , \62773 , \62774 ,
         \62775 , \62776 , \62777 , \62778 , \62779 , \62780 , \62781 , \62782 , \62783 , \62784 ,
         \62785 , \62786 , \62787 , \62788 , \62789 , \62790 , \62791 , \62792 , \62793 , \62794 ,
         \62795 , \62796 , \62797 , \62798 , \62799 , \62800 , \62801 , \62802 , \62803 , \62804 ,
         \62805 , \62806 , \62807 , \62808 , \62809 , \62810 , \62811 , \62812 , \62813 , \62814 ,
         \62815 , \62816 , \62817 , \62818 , \62819 , \62820 , \62821 , \62822 , \62823 , \62824 ,
         \62825 , \62826 , \62827 , \62828 , \62829 , \62830 , \62831 , \62832 , \62833 , \62834 ,
         \62835 , \62836 , \62837 , \62838 , \62839 , \62840 , \62841 , \62842 , \62843 , \62844 ,
         \62845 , \62846 , \62847 , \62848 , \62849 , \62850 , \62851 , \62852 , \62853 , \62854 ,
         \62855 , \62856 , \62857 , \62858 , \62859 , \62860 , \62861 , \62862 , \62863 , \62864 ,
         \62865 , \62866 , \62867 , \62868 , \62869 , \62870 , \62871 , \62872 , \62873 , \62874 ,
         \62875 , \62876 , \62877 , \62878 , \62879 , \62880 , \62881 , \62882 , \62883 , \62884 ,
         \62885 , \62886 , \62887 , \62888 , \62889 , \62890 , \62891 , \62892 , \62893 , \62894 ,
         \62895 , \62896 , \62897 , \62898 , \62899 , \62900 , \62901 , \62902 , \62903 , \62904 ,
         \62905 , \62906 , \62907 , \62908 , \62909 , \62910 , \62911 , \62912 , \62913 , \62914 ,
         \62915 , \62916 , \62917 , \62918 , \62919 , \62920 , \62921 , \62922 , \62923 , \62924 ,
         \62925 , \62926 , \62927 , \62928 , \62929 , \62930 , \62931 , \62932 , \62933 , \62934 ,
         \62935 , \62936 , \62937 , \62938 , \62939 , \62940 , \62941 , \62942 , \62943 , \62944 ,
         \62945 , \62946 , \62947 , \62948 , \62949 , \62950 , \62951 , \62952 , \62953 , \62954 ,
         \62955 , \62956 , \62957 , \62958 , \62959 , \62960 , \62961 , \62962 , \62963 , \62964 ,
         \62965 , \62966 , \62967 , \62968 , \62969 , \62970 , \62971 , \62972 , \62973 , \62974 ,
         \62975 , \62976 , \62977 , \62978 , \62979 , \62980 , \62981 , \62982 , \62983 , \62984 ,
         \62985 , \62986 , \62987 , \62988 , \62989 , \62990 , \62991 , \62992 , \62993 , \62994 ,
         \62995 , \62996 , \62997 , \62998 , \62999 , \63000 , \63001 , \63002 , \63003 , \63004 ,
         \63005 , \63006 , \63007 , \63008 , \63009 , \63010 , \63011 , \63012 , \63013 , \63014 ,
         \63015 , \63016 , \63017 , \63018 , \63019 , \63020 , \63021 , \63022 , \63023 , \63024 ,
         \63025 , \63026 , \63027 , \63028 , \63029 , \63030 , \63031 , \63032 , \63033 , \63034 ,
         \63035 , \63036 , \63037 , \63038 , \63039 , \63040 , \63041 , \63042 , \63043 , \63044 ,
         \63045 , \63046 , \63047 , \63048 , \63049 , \63050 , \63051 , \63052 , \63053 , \63054 ,
         \63055 , \63056 , \63057 , \63058 , \63059 , \63060 , \63061 , \63062 , \63063 , \63064 ,
         \63065 , \63066 , \63067 , \63068 , \63069 , \63070 , \63071 , \63072 , \63073 , \63074 ,
         \63075 , \63076 , \63077 , \63078 , \63079 , \63080 , \63081 , \63082 , \63083 , \63084 ,
         \63085 , \63086 , \63087 , \63088 , \63089 , \63090 , \63091 , \63092 , \63093 , \63094 ,
         \63095 , \63096 , \63097 , \63098 , \63099 , \63100 , \63101 , \63102 , \63103 , \63104 ,
         \63105 , \63106 , \63107 , \63108 , \63109 , \63110 , \63111 , \63112 , \63113 , \63114 ,
         \63115 , \63116 , \63117 , \63118 , \63119 , \63120 , \63121 , \63122 , \63123 , \63124 ,
         \63125 , \63126 , \63127 , \63128 , \63129 , \63130 , \63131 , \63132 , \63133 , \63134 ,
         \63135 , \63136 , \63137 , \63138 , \63139 , \63140 , \63141 , \63142 , \63143 , \63144 ,
         \63145 , \63146 , \63147 , \63148 , \63149 , \63150 , \63151 , \63152 , \63153 , \63154 ,
         \63155 , \63156 , \63157 , \63158 , \63159 , \63160 , \63161 , \63162 , \63163 , \63164 ,
         \63165 , \63166 , \63167 , \63168 , \63169 , \63170 , \63171 , \63172 , \63173 , \63174 ,
         \63175 , \63176 , \63177 , \63178 , \63179 , \63180 , \63181 , \63182 , \63183 , \63184 ,
         \63185 , \63186 , \63187 , \63188 , \63189 , \63190 , \63191 , \63192 , \63193 , \63194 ,
         \63195 , \63196 , \63197 , \63198 , \63199 , \63200 , \63201 , \63202 , \63203 , \63204 ,
         \63205 , \63206 , \63207 , \63208 , \63209 , \63210 , \63211 , \63212 , \63213 , \63214 ,
         \63215 , \63216 , \63217 , \63218 , \63219 , \63220 , \63221 , \63222 , \63223 , \63224 ,
         \63225 , \63226 , \63227 , \63228 , \63229 , \63230 , \63231 , \63232 , \63233 , \63234 ,
         \63235 , \63236 , \63237 , \63238 , \63239 , \63240 , \63241 , \63242 , \63243 , \63244 ,
         \63245 , \63246 , \63247 , \63248 , \63249 , \63250 , \63251 , \63252 , \63253 , \63254 ,
         \63255 , \63256 , \63257 , \63258 , \63259 , \63260 , \63261 , \63262 , \63263 , \63264 ,
         \63265 , \63266 , \63267 , \63268 , \63269 , \63270 , \63271 , \63272 , \63273 , \63274 ,
         \63275 , \63276 , \63277 , \63278 , \63279 , \63280 , \63281 , \63282 , \63283 , \63284 ,
         \63285 , \63286 , \63287 , \63288 , \63289 , \63290 , \63291 , \63292 , \63293 , \63294 ,
         \63295 , \63296 , \63297 , \63298 , \63299 , \63300 , \63301 , \63302 , \63303 , \63304 ,
         \63305 , \63306 , \63307 , \63308 , \63309 , \63310 , \63311 , \63312 , \63313 , \63314 ,
         \63315 , \63316 , \63317 , \63318 , \63319 , \63320 , \63321 , \63322 , \63323 , \63324 ,
         \63325 , \63326 , \63327 , \63328 , \63329 , \63330 , \63331 , \63332 , \63333 , \63334 ,
         \63335 , \63336 , \63337 , \63338 , \63339 , \63340 , \63341 , \63342 , \63343 , \63344 ,
         \63345 , \63346 , \63347 , \63348 , \63349 , \63350 , \63351 , \63352 , \63353 , \63354 ,
         \63355 , \63356 , \63357 , \63358 , \63359 , \63360 , \63361 , \63362 , \63363 , \63364 ,
         \63365 , \63366 , \63367 , \63368 , \63369 , \63370 , \63371 , \63372 , \63373 , \63374 ,
         \63375 , \63376 , \63377 , \63378 , \63379 , \63380 , \63381 , \63382 , \63383 , \63384 ,
         \63385 , \63386 , \63387 , \63388 , \63389 , \63390 , \63391 , \63392 , \63393 , \63394 ,
         \63395 , \63396 , \63397 , \63398 , \63399 , \63400 , \63401 , \63402 , \63403 , \63404 ,
         \63405 , \63406 , \63407 , \63408 , \63409 , \63410 , \63411 , \63412 , \63413 , \63414 ,
         \63415 , \63416 , \63417 , \63418 , \63419 , \63420 , \63421 , \63422 , \63423 , \63424 ,
         \63425 , \63426 , \63427 , \63428 , \63429 , \63430 , \63431 , \63432 , \63433 , \63434 ,
         \63435 , \63436 , \63437 , \63438 , \63439 , \63440 , \63441 , \63442 , \63443 , \63444 ,
         \63445 , \63446 , \63447 , \63448 , \63449 , \63450 , \63451 , \63452 , \63453 , \63454 ,
         \63455 , \63456 , \63457 , \63458 , \63459 , \63460 , \63461 , \63462 , \63463 , \63464 ,
         \63465 , \63466 , \63467 , \63468 , \63469 , \63470 , \63471 , \63472 , \63473 , \63474 ,
         \63475 , \63476 , \63477 , \63478 , \63479 , \63480 , \63481 , \63482 , \63483 , \63484 ,
         \63485 , \63486 , \63487 , \63488 , \63489 , \63490 , \63491 , \63492 , \63493 , \63494 ,
         \63495 , \63496 , \63497 , \63498 , \63499 , \63500 , \63501 , \63502 , \63503 , \63504 ,
         \63505 , \63506 , \63507 , \63508 , \63509 , \63510 , \63511 , \63512 , \63513 , \63514 ,
         \63515 , \63516 , \63517 , \63518 , \63519 , \63520 , \63521 , \63522 , \63523 , \63524 ,
         \63525 , \63526 , \63527 , \63528 , \63529 , \63530 , \63531 , \63532 , \63533 , \63534 ,
         \63535 , \63536 , \63537 , \63538 , \63539 , \63540 , \63541 , \63542 , \63543 , \63544 ,
         \63545 , \63546 , \63547 , \63548 , \63549 , \63550 , \63551 , \63552 , \63553 , \63554 ,
         \63555 , \63556 , \63557 , \63558 , \63559 , \63560 , \63561 , \63562 , \63563 , \63564 ,
         \63565 , \63566 , \63567 , \63568 , \63569 , \63570 , \63571 , \63572 , \63573 , \63574 ,
         \63575 , \63576 , \63577 , \63578 , \63579 , \63580 , \63581 , \63582 , \63583 , \63584 ,
         \63585 , \63586 , \63587 , \63588 , \63589 , \63590 , \63591 , \63592 , \63593 , \63594 ,
         \63595 , \63596 , \63597 , \63598 , \63599 , \63600 , \63601 , \63602 , \63603 , \63604 ,
         \63605 , \63606 , \63607 , \63608 , \63609 , \63610 , \63611 , \63612 , \63613 , \63614 ,
         \63615 , \63616 , \63617 , \63618 , \63619 , \63620 , \63621 , \63622 , \63623 , \63624 ,
         \63625 , \63626 , \63627 , \63628 , \63629 , \63630 , \63631 , \63632 , \63633 , \63634 ,
         \63635 , \63636 , \63637 , \63638 , \63639 , \63640 , \63641 , \63642 , \63643 , \63644 ,
         \63645 , \63646 , \63647 , \63648 , \63649 , \63650 , \63651 , \63652 , \63653 , \63654 ,
         \63655 , \63656 , \63657 , \63658 , \63659 , \63660 , \63661 , \63662 , \63663 , \63664 ,
         \63665 , \63666 , \63667 , \63668 , \63669 , \63670 , \63671 , \63672 , \63673 , \63674 ,
         \63675 , \63676 , \63677 , \63678 , \63679 , \63680 , \63681 , \63682 , \63683 , \63684 ,
         \63685 , \63686 , \63687 , \63688 , \63689 , \63690 , \63691 , \63692 , \63693 , \63694 ,
         \63695 , \63696 , \63697 , \63698 , \63699 , \63700 , \63701 , \63702 , \63703 , \63704 ,
         \63705 , \63706 , \63707 , \63708 , \63709 , \63710 , \63711 , \63712 , \63713 , \63714 ,
         \63715 , \63716 , \63717 , \63718 , \63719 , \63720 , \63721 , \63722 , \63723 , \63724 ,
         \63725 , \63726 , \63727 , \63728 , \63729 , \63730 , \63731 , \63732 , \63733 , \63734 ,
         \63735 , \63736 , \63737 , \63738 , \63739 , \63740 , \63741 , \63742 , \63743 , \63744 ,
         \63745 , \63746 , \63747 , \63748 , \63749 , \63750 , \63751 , \63752 , \63753 , \63754 ,
         \63755 , \63756 , \63757 , \63758 , \63759 , \63760 , \63761 , \63762 , \63763 , \63764 ,
         \63765 , \63766 , \63767 , \63768 , \63769 , \63770 , \63771 , \63772 , \63773 , \63774 ,
         \63775 , \63776 , \63777 , \63778 , \63779 , \63780 , \63781 , \63782 , \63783 , \63784 ,
         \63785 , \63786 , \63787 , \63788 , \63789 , \63790 , \63791 , \63792 , \63793 , \63794 ,
         \63795 , \63796 , \63797 , \63798 , \63799 , \63800 , \63801 , \63802 , \63803 , \63804 ,
         \63805 , \63806 , \63807 , \63808 , \63809 , \63810 , \63811 , \63812 , \63813 , \63814 ,
         \63815 , \63816 , \63817 , \63818 , \63819 , \63820 , \63821 , \63822 , \63823 , \63824 ,
         \63825 , \63826 , \63827 , \63828 , \63829 , \63830 , \63831 , \63832 , \63833 , \63834 ,
         \63835 , \63836 , \63837 , \63838 , \63839 , \63840 , \63841 , \63842 , \63843 , \63844 ,
         \63845 , \63846 , \63847 , \63848 , \63849 , \63850 , \63851 , \63852 , \63853 , \63854 ,
         \63855 , \63856 , \63857 , \63858 , \63859 , \63860 , \63861 , \63862 , \63863 , \63864 ,
         \63865 , \63866 , \63867 , \63868 , \63869 , \63870 , \63871 , \63872 , \63873 , \63874 ,
         \63875 , \63876 , \63877 , \63878 , \63879 , \63880 , \63881 , \63882 , \63883 , \63884 ,
         \63885 , \63886 , \63887 , \63888 , \63889 , \63890 , \63891 , \63892 , \63893 , \63894 ,
         \63895 , \63896 , \63897 , \63898 , \63899 , \63900 , \63901 , \63902 , \63903 , \63904 ,
         \63905 , \63906 , \63907 , \63908 , \63909 , \63910 , \63911 , \63912 , \63913 , \63914 ,
         \63915 , \63916 , \63917 , \63918 , \63919 , \63920 , \63921 , \63922 , \63923 , \63924 ,
         \63925 , \63926 , \63927 , \63928 , \63929 , \63930 , \63931 , \63932 , \63933 , \63934 ,
         \63935 , \63936 , \63937 , \63938 , \63939 , \63940 , \63941 , \63942 , \63943 , \63944 ,
         \63945 , \63946 , \63947 , \63948 , \63949 , \63950 , \63951 , \63952 , \63953 , \63954 ,
         \63955 , \63956 , \63957 , \63958 , \63959 , \63960 , \63961 , \63962 , \63963 , \63964 ,
         \63965 , \63966 , \63967 , \63968 , \63969 , \63970 , \63971 , \63972 , \63973 , \63974 ,
         \63975 , \63976 , \63977 , \63978 , \63979 , \63980 , \63981 , \63982 , \63983 , \63984 ,
         \63985 , \63986 , \63987 , \63988 , \63989 , \63990 , \63991 , \63992 , \63993 , \63994 ,
         \63995 , \63996 , \63997 , \63998 , \63999 , \64000 , \64001 , \64002 , \64003 , \64004 ,
         \64005 , \64006 , \64007 , \64008 , \64009 , \64010 , \64011 , \64012 , \64013 , \64014 ,
         \64015 , \64016 , \64017 , \64018 , \64019 , \64020 , \64021 , \64022 , \64023 , \64024 ,
         \64025 , \64026 , \64027 , \64028 , \64029 , \64030 , \64031 , \64032 , \64033 , \64034 ,
         \64035 , \64036 , \64037 , \64038 , \64039 , \64040 , \64041 , \64042 , \64043 , \64044 ,
         \64045 , \64046 , \64047 , \64048 , \64049 , \64050 , \64051 , \64052 , \64053 , \64054 ,
         \64055 , \64056 , \64057 , \64058 , \64059 , \64060 , \64061 , \64062 , \64063 , \64064 ,
         \64065 , \64066 , \64067 , \64068 , \64069 , \64070 , \64071 , \64072 , \64073 , \64074 ,
         \64075 , \64076 , \64077 , \64078 , \64079 , \64080 , \64081 , \64082 , \64083 , \64084 ,
         \64085 , \64086 , \64087 , \64088 , \64089 , \64090 , \64091 , \64092 , \64093 , \64094 ,
         \64095 , \64096 , \64097 , \64098 , \64099 , \64100 , \64101 , \64102 , \64103 , \64104 ,
         \64105 , \64106 , \64107 , \64108 , \64109 , \64110 , \64111 , \64112 , \64113 , \64114 ,
         \64115 , \64116 , \64117 , \64118 , \64119 , \64120 , \64121 , \64122 , \64123 , \64124 ,
         \64125 , \64126 , \64127 , \64128 , \64129 , \64130 , \64131 , \64132 , \64133 , \64134 ,
         \64135 , \64136 , \64137 , \64138 , \64139 , \64140 , \64141 , \64142 , \64143 , \64144 ,
         \64145 , \64146 , \64147 , \64148 , \64149 , \64150 , \64151 , \64152 , \64153 , \64154 ,
         \64155 , \64156 , \64157 , \64158 , \64159 , \64160 , \64161 , \64162 , \64163 , \64164 ,
         \64165 , \64166 , \64167 , \64168 , \64169 , \64170 , \64171 , \64172 , \64173 , \64174 ,
         \64175 , \64176 , \64177 , \64178 , \64179 , \64180 , \64181 , \64182 , \64183 , \64184 ,
         \64185 , \64186 , \64187 , \64188 , \64189 , \64190 , \64191 , \64192 , \64193 , \64194 ,
         \64195 , \64196 , \64197 , \64198 , \64199 , \64200 , \64201 , \64202 , \64203 , \64204 ,
         \64205 , \64206 , \64207 , \64208 , \64209 , \64210 , \64211 , \64212 , \64213 , \64214 ,
         \64215 , \64216 , \64217 , \64218 , \64219 , \64220 , \64221 , \64222 , \64223 , \64224 ,
         \64225 , \64226 , \64227 , \64228 , \64229 , \64230 , \64231 , \64232 , \64233 , \64234 ,
         \64235 , \64236 , \64237 , \64238 , \64239 , \64240 , \64241 , \64242 , \64243 , \64244 ,
         \64245 , \64246 , \64247 , \64248 , \64249 , \64250 , \64251 , \64252 , \64253 , \64254 ,
         \64255 , \64256 , \64257 , \64258 , \64259 , \64260 , \64261 , \64262 , \64263 , \64264 ,
         \64265 , \64266 , \64267 , \64268 , \64269 , \64270 , \64271 , \64272 , \64273 , \64274 ,
         \64275 , \64276 , \64277 , \64278 , \64279 , \64280 , \64281 , \64282 , \64283 , \64284 ,
         \64285 , \64286 , \64287 , \64288 , \64289 , \64290 , \64291 , \64292 , \64293 , \64294 ,
         \64295 , \64296 , \64297 , \64298 , \64299 , \64300 , \64301 , \64302 , \64303 , \64304 ,
         \64305 , \64306 , \64307 , \64308 , \64309 , \64310 , \64311 , \64312 , \64313 , \64314 ,
         \64315 , \64316 , \64317 , \64318 , \64319 , \64320 , \64321 , \64322 , \64323 , \64324 ,
         \64325 , \64326 , \64327 , \64328 , \64329 , \64330 , \64331 , \64332 , \64333 , \64334 ,
         \64335 , \64336 , \64337 , \64338 , \64339 , \64340 , \64341 , \64342 , \64343 , \64344 ,
         \64345 , \64346 , \64347 , \64348 , \64349 , \64350 , \64351 , \64352 , \64353 , \64354 ,
         \64355 , \64356 , \64357 , \64358 , \64359 , \64360 , \64361 , \64362 , \64363 , \64364 ,
         \64365 , \64366 , \64367 , \64368 , \64369 , \64370 , \64371 , \64372 , \64373 , \64374 ,
         \64375 , \64376 , \64377 , \64378 , \64379 , \64380 , \64381 , \64382 , \64383 , \64384 ,
         \64385 , \64386 , \64387 , \64388 , \64389 , \64390 , \64391 , \64392 , \64393 , \64394 ,
         \64395 , \64396 , \64397 , \64398 , \64399 , \64400 , \64401 , \64402 , \64403 , \64404 ,
         \64405 , \64406 , \64407 , \64408 , \64409 , \64410 , \64411 , \64412 , \64413 , \64414 ,
         \64415 , \64416 , \64417 , \64418 , \64419 , \64420 , \64421 , \64422 , \64423 , \64424 ,
         \64425 , \64426 , \64427 , \64428 , \64429 , \64430 , \64431 , \64432 , \64433 , \64434 ,
         \64435 , \64436 , \64437 , \64438 , \64439 , \64440 , \64441 , \64442 , \64443 , \64444 ,
         \64445 , \64446 , \64447 , \64448 , \64449 , \64450 , \64451 , \64452 , \64453 , \64454 ,
         \64455 , \64456 , \64457 , \64458 , \64459 , \64460 , \64461 , \64462 , \64463 , \64464 ,
         \64465 , \64466 , \64467 , \64468 , \64469 , \64470 , \64471 , \64472 , \64473 , \64474 ,
         \64475 , \64476 , \64477 , \64478 , \64479 , \64480 , \64481 , \64482 , \64483 , \64484 ,
         \64485 , \64486 , \64487 , \64488 , \64489 , \64490 , \64491 , \64492 , \64493 , \64494 ,
         \64495 , \64496 , \64497 , \64498 , \64499 , \64500 , \64501 , \64502 , \64503 , \64504 ,
         \64505 , \64506 , \64507 , \64508 , \64509 , \64510 , \64511 , \64512 , \64513 , \64514 ,
         \64515 , \64516 , \64517 , \64518 , \64519 , \64520 , \64521 , \64522 , \64523 , \64524 ,
         \64525 , \64526 , \64527 , \64528 , \64529 , \64530 , \64531 , \64532 , \64533 , \64534 ,
         \64535 , \64536 , \64537 , \64538 , \64539 , \64540 , \64541 , \64542 , \64543 , \64544 ,
         \64545 , \64546 , \64547 , \64548 , \64549 , \64550 , \64551 , \64552 , \64553 , \64554 ,
         \64555 , \64556 , \64557 , \64558 , \64559 , \64560 , \64561 , \64562 , \64563 , \64564 ,
         \64565 , \64566 , \64567 , \64568 , \64569 , \64570 , \64571 , \64572 , \64573 , \64574 ,
         \64575 , \64576 , \64577 , \64578 , \64579 , \64580 , \64581 , \64582 , \64583 , \64584 ,
         \64585 , \64586 , \64587 , \64588 , \64589 , \64590 , \64591 , \64592 , \64593 , \64594 ,
         \64595 , \64596 , \64597 , \64598 , \64599 , \64600 , \64601 , \64602 , \64603 , \64604 ,
         \64605 , \64606 , \64607 , \64608 , \64609 , \64610 , \64611 , \64612 , \64613 , \64614 ,
         \64615 , \64616 , \64617 , \64618 , \64619 , \64620 , \64621 , \64622 , \64623 , \64624 ,
         \64625 , \64626 , \64627 , \64628 , \64629 , \64630 , \64631 , \64632 , \64633 , \64634 ,
         \64635 , \64636 , \64637 , \64638 , \64639 , \64640 , \64641 , \64642 , \64643 , \64644 ,
         \64645 , \64646 , \64647 , \64648 , \64649 , \64650 , \64651 , \64652 , \64653 , \64654 ,
         \64655 , \64656 , \64657 , \64658 , \64659 , \64660 , \64661 , \64662 , \64663 , \64664 ,
         \64665 , \64666 , \64667 , \64668 , \64669 , \64670 , \64671 , \64672 , \64673 , \64674 ,
         \64675 , \64676 , \64677 , \64678 , \64679 , \64680 , \64681 , \64682 , \64683 , \64684 ,
         \64685 , \64686 , \64687 , \64688 , \64689 , \64690 , \64691 , \64692 , \64693 , \64694 ,
         \64695 , \64696 , \64697 , \64698 , \64699 , \64700 , \64701 , \64702 , \64703 , \64704 ,
         \64705 , \64706 , \64707 , \64708 , \64709 , \64710 , \64711 , \64712 , \64713 , \64714 ,
         \64715 , \64716 , \64717 , \64718 , \64719 , \64720 , \64721 , \64722 , \64723 , \64724 ,
         \64725 , \64726 , \64727 , \64728 , \64729 , \64730 , \64731 , \64732 , \64733 , \64734 ,
         \64735 , \64736 , \64737 , \64738 , \64739 , \64740 , \64741 , \64742 , \64743 , \64744 ,
         \64745 , \64746 , \64747 , \64748 , \64749 , \64750 , \64751 , \64752 , \64753 , \64754 ,
         \64755 , \64756 , \64757 , \64758 , \64759 , \64760 , \64761 , \64762 , \64763 , \64764 ,
         \64765 , \64766 , \64767 , \64768 , \64769 , \64770 , \64771 , \64772 , \64773 , \64774 ,
         \64775 , \64776 , \64777 , \64778 , \64779 , \64780 , \64781 , \64782 , \64783 , \64784 ,
         \64785 , \64786 , \64787 , \64788 , \64789 , \64790 , \64791 , \64792 , \64793 , \64794 ,
         \64795 , \64796 , \64797 , \64798 , \64799 , \64800 , \64801 , \64802 , \64803 , \64804 ,
         \64805 , \64806 , \64807 , \64808 , \64809 , \64810 , \64811 , \64812 , \64813 , \64814 ,
         \64815 , \64816 , \64817 , \64818 , \64819 , \64820 , \64821 , \64822 , \64823 , \64824 ,
         \64825 , \64826 , \64827 , \64828 , \64829 , \64830 , \64831 , \64832 , \64833 , \64834 ,
         \64835 , \64836 , \64837 , \64838 , \64839 , \64840 , \64841 , \64842 , \64843 , \64844 ,
         \64845 , \64846 , \64847 , \64848 , \64849 , \64850 , \64851 , \64852 , \64853 , \64854 ,
         \64855 , \64856 , \64857 , \64858 , \64859 , \64860 , \64861 , \64862 , \64863 , \64864 ,
         \64865 , \64866 , \64867 , \64868 , \64869 , \64870 , \64871 , \64872 , \64873 , \64874 ,
         \64875 , \64876 , \64877 , \64878 , \64879 , \64880 , \64881 , \64882 , \64883 , \64884 ,
         \64885 , \64886 , \64887 , \64888 , \64889 , \64890 , \64891 , \64892 , \64893 , \64894 ,
         \64895 , \64896 , \64897 , \64898 , \64899 , \64900 , \64901 , \64902 , \64903 , \64904 ,
         \64905 , \64906 , \64907 , \64908 , \64909 , \64910 , \64911 , \64912 , \64913 , \64914 ,
         \64915 , \64916 , \64917 , \64918 , \64919 , \64920 , \64921 , \64922 , \64923 , \64924 ,
         \64925 , \64926 , \64927 , \64928 , \64929 , \64930 , \64931 , \64932 , \64933 , \64934 ,
         \64935 , \64936 , \64937 , \64938 , \64939 , \64940 , \64941 , \64942 , \64943 , \64944 ,
         \64945 , \64946 , \64947 , \64948 , \64949 , \64950 , \64951 , \64952 , \64953 , \64954 ,
         \64955 , \64956 , \64957 , \64958 , \64959 , \64960 , \64961 , \64962 , \64963 , \64964 ,
         \64965 , \64966 , \64967 , \64968 , \64969 , \64970 , \64971 , \64972 , \64973 , \64974 ,
         \64975 , \64976 , \64977 , \64978 , \64979 , \64980 , \64981 , \64982 , \64983 , \64984 ,
         \64985 , \64986 , \64987 , \64988 , \64989 , \64990 , \64991 , \64992 , \64993 , \64994 ,
         \64995 , \64996 , \64997 , \64998 , \64999 , \65000 , \65001 , \65002 , \65003 , \65004 ,
         \65005 , \65006 , \65007 , \65008 , \65009 , \65010 , \65011 , \65012 , \65013 , \65014 ,
         \65015 , \65016 , \65017 , \65018 , \65019 , \65020 , \65021 , \65022 , \65023 , \65024 ,
         \65025 , \65026 , \65027 , \65028 , \65029 , \65030 , \65031 , \65032 , \65033 , \65034 ,
         \65035 , \65036 , \65037 , \65038 , \65039 , \65040 , \65041 , \65042 , \65043 , \65044 ,
         \65045 , \65046 , \65047 , \65048 , \65049 , \65050 , \65051 , \65052 , \65053 , \65054 ,
         \65055 , \65056 , \65057 , \65058 , \65059 , \65060 , \65061 , \65062 , \65063 , \65064 ,
         \65065 , \65066 , \65067 , \65068 , \65069 , \65070 , \65071 , \65072 , \65073 , \65074 ,
         \65075 , \65076 , \65077 , \65078 , \65079 , \65080 , \65081 , \65082 , \65083 , \65084 ,
         \65085 , \65086 , \65087 , \65088 , \65089 , \65090 , \65091 , \65092 , \65093 , \65094 ,
         \65095 , \65096 , \65097 , \65098 , \65099 , \65100 , \65101 , \65102 , \65103 , \65104 ,
         \65105 , \65106 , \65107 , \65108 , \65109 , \65110 , \65111 , \65112 , \65113 , \65114 ,
         \65115 , \65116 , \65117 , \65118 , \65119 , \65120 , \65121 , \65122 , \65123 , \65124 ,
         \65125 , \65126 , \65127 , \65128 , \65129 , \65130 , \65131 , \65132 , \65133 , \65134 ,
         \65135 , \65136 , \65137 , \65138 , \65139 , \65140 , \65141 , \65142 , \65143 , \65144 ,
         \65145 , \65146 , \65147 , \65148 , \65149 , \65150 , \65151 , \65152 , \65153 , \65154 ,
         \65155 , \65156 , \65157 , \65158 , \65159 , \65160 , \65161 , \65162 , \65163 , \65164 ,
         \65165 , \65166 , \65167 , \65168 , \65169 , \65170 , \65171 , \65172 , \65173 , \65174 ,
         \65175 , \65176 , \65177 , \65178 , \65179 , \65180 , \65181 , \65182 , \65183 , \65184 ,
         \65185 , \65186 , \65187 , \65188 , \65189 , \65190 , \65191 , \65192 , \65193 , \65194 ,
         \65195 , \65196 , \65197 , \65198 , \65199 , \65200 , \65201 , \65202 , \65203 , \65204 ,
         \65205 , \65206 , \65207 , \65208 , \65209 , \65210 , \65211 , \65212 , \65213 , \65214 ,
         \65215 , \65216 , \65217 , \65218 , \65219 , \65220 , \65221 , \65222 , \65223 , \65224 ,
         \65225 , \65226 , \65227 , \65228 , \65229 , \65230 , \65231 , \65232 , \65233 , \65234 ,
         \65235 , \65236 , \65237 , \65238 , \65239 , \65240 , \65241 , \65242 , \65243 , \65244 ,
         \65245 , \65246 , \65247 , \65248 , \65249 , \65250 , \65251 , \65252 , \65253 , \65254 ,
         \65255 , \65256 , \65257 , \65258 , \65259 , \65260 , \65261 , \65262 , \65263 , \65264 ,
         \65265 , \65266 , \65267 , \65268 , \65269 , \65270 , \65271 , \65272 , \65273 , \65274 ,
         \65275 , \65276 , \65277 , \65278 , \65279 , \65280 , \65281 , \65282 , \65283 , \65284 ,
         \65285 , \65286 , \65287 , \65288 , \65289 , \65290 , \65291 , \65292 , \65293 , \65294 ,
         \65295 , \65296 , \65297 , \65298 , \65299 , \65300 , \65301 , \65302 , \65303 , \65304 ,
         \65305 , \65306 , \65307 , \65308 , \65309 , \65310 , \65311 , \65312 , \65313 , \65314 ,
         \65315 , \65316 , \65317 , \65318 , \65319 , \65320 , \65321 , \65322 , \65323 , \65324 ,
         \65325 , \65326 , \65327 , \65328 , \65329 , \65330 , \65331 , \65332 , \65333 , \65334 ,
         \65335 , \65336 , \65337 , \65338 , \65339 , \65340 , \65341 , \65342 , \65343 , \65344 ,
         \65345 , \65346 , \65347 , \65348 , \65349 , \65350 , \65351 , \65352 , \65353 , \65354 ,
         \65355 , \65356 , \65357 , \65358 , \65359 , \65360 , \65361 , \65362 , \65363 , \65364 ,
         \65365 , \65366 , \65367 , \65368 , \65369 , \65370 , \65371 , \65372 , \65373 , \65374 ,
         \65375 , \65376 , \65377 , \65378 , \65379 , \65380 , \65381 , \65382 , \65383 , \65384 ,
         \65385 , \65386 , \65387 , \65388 , \65389 , \65390 , \65391 , \65392 , \65393 , \65394 ,
         \65395 , \65396 , \65397 , \65398 , \65399 , \65400 , \65401 , \65402 , \65403 , \65404 ,
         \65405 , \65406 , \65407 , \65408 , \65409 , \65410 , \65411 , \65412 , \65413 , \65414 ,
         \65415 , \65416 , \65417 , \65418 , \65419 , \65420 , \65421 , \65422 , \65423 , \65424 ,
         \65425 , \65426 , \65427 , \65428 , \65429 , \65430 , \65431 , \65432 , \65433 , \65434 ,
         \65435 , \65436 , \65437 , \65438 , \65439 , \65440 , \65441 , \65442 , \65443 , \65444 ,
         \65445 , \65446 , \65447 , \65448 , \65449 , \65450 , \65451 , \65452 , \65453 , \65454 ,
         \65455 , \65456 , \65457 , \65458 , \65459 , \65460 , \65461 , \65462 , \65463 , \65464 ,
         \65465 , \65466 , \65467 , \65468 , \65469 , \65470 , \65471 , \65472 , \65473 , \65474 ,
         \65475 , \65476 , \65477 , \65478 , \65479 , \65480 , \65481 , \65482 , \65483 , \65484 ,
         \65485 , \65486 , \65487 , \65488 , \65489 , \65490 , \65491 , \65492 , \65493 , \65494 ,
         \65495 , \65496 , \65497 , \65498 , \65499 , \65500 , \65501 , \65502 , \65503 , \65504 ,
         \65505 , \65506 , \65507 , \65508 , \65509 , \65510 , \65511 , \65512 , \65513 , \65514 ,
         \65515 , \65516 , \65517 , \65518 , \65519 , \65520 , \65521 , \65522 , \65523 , \65524 ,
         \65525 , \65526 , \65527 , \65528 , \65529 , \65530 , \65531 , \65532 , \65533 , \65534 ,
         \65535 , \65536 , \65537 , \65538 , \65539 , \65540 , \65541 , \65542 , \65543 , \65544 ,
         \65545 , \65546 , \65547 , \65548 , \65549 , \65550 , \65551 , \65552 , \65553 , \65554 ,
         \65555 , \65556 , \65557 , \65558 , \65559 , \65560 , \65561 , \65562 , \65563 , \65564 ,
         \65565 , \65566 , \65567 , \65568 , \65569 , \65570 , \65571 , \65572 , \65573 , \65574 ,
         \65575 , \65576 , \65577 , \65578 , \65579 , \65580 , \65581_nG10344 , \65582 , \65583 , \65584 ,
         \65585 , \65586 , \65587 , \65588 , \65589_nG10315 , \65590 , \65591 , \65592 , \65593 , \65594 ,
         \65595 , \65596 , \65597_nG102d0 , \65598 , \65599 , \65600 , \65601 , \65602 , \65603 , \65604 ,
         \65605_nG1026f , \65606 , \65607 , \65608 , \65609 , \65610 , \65611 , \65612 , \65613_nG10201 , \65614 ,
         \65615 , \65616 , \65617 , \65618 , \65619 , \65620 , \65621_nG10176 , \65622 , \65623 , \65624 ,
         \65625 , \65626 , \65627 , \65628 , \65629_nG100f9 , \65630 , \65631 , \65632 , \65633 , \65634 ,
         \65635 , \65636 , \65637_nG1005e , \65638 , \65639 , \65640 , \65641 , \65642 , \65643 , \65644 ,
         \65645_nGff9a , \65646 , \65647 , \65648 , \65649 , \65650 , \65651 , \65652 , \65653_nGfed3 , \65654 ,
         \65655 , \65656 , \65657 , \65658 , \65659 , \65660 , \65661_nGfded , \65662 , \65663 , \65664 ,
         \65665 , \65666 , \65667 , \65668 , \65669_nGfd15 , \65670 , \65671 , \65672 , \65673 , \65674 ,
         \65675 , \65676 , \65677_nGfc38 , \65678 , \65679 , \65680 , \65681 , \65682 , \65683 , \65684 ,
         \65685_nGfb46 , \65686 , \65687 , \65688 , \65689 , \65690 , \65691 , \65692 , \65693_nGfa24 , \65694 ,
         \65695 , \65696 , \65697 , \65698 , \65699 , \65700 , \65701_nGf914 , \65702 , \65703 , \65704 ,
         \65705 , \65706 , \65707 , \65708 , \65709_nGf7e6 , \65710 , \65711 , \65712 , \65713 , \65714 ,
         \65715 , \65716 , \65717_nGf6c6 , \65718 , \65719 , \65720 , \65721 , \65722 , \65723 , \65724 ,
         \65725_nGf581 , \65726 , \65727 , \65728 , \65729 , \65730 , \65731 , \65732 , \65733_nGf429 , \65734 ,
         \65735 , \65736 , \65737 , \65738 , \65739 , \65740 , \65741_nGf2c7 , \65742 , \65743 , \65744 ,
         \65745 , \65746 , \65747 , \65748 , \65749_nGf156 , \65750 , \65751 , \65752 , \65753 , \65754 ,
         \65755 , \65756 , \65757_nGefd8 , \65758 , \65759 , \65760 , \65761 , \65762 , \65763 , \65764 ,
         \65765_nGee3c , \65766 , \65767 , \65768 , \65769 , \65770 , \65771 , \65772 , \65773_nGec7d , \65774 ,
         \65775 , \65776 , \65777 , \65778 , \65779 , \65780 , \65781_nGea87 , \65782 , \65783 , \65784 ,
         \65785 , \65786 , \65787 , \65788 , \65789_nGe8b1 , \65790 , \65791 , \65792 , \65793 , \65794 ,
         \65795 , \65796 , \65797_nGe6d4 , \65798 , \65799 , \65800 , \65801 , \65802 , \65803 , \65804 ,
         \65805_nGe4e7 , \65806 , \65807 , \65808 , \65809 , \65810 , \65811 , \65812 , \65813_nGe2e5 , \65814 ,
         \65815 , \65816 , \65817 , \65818 , \65819 , \65820 , \65821_nGe0da , \65822 , \65823 , \65824 ,
         \65825 , \65826 , \65827 , \65828 , \65829_nGdec8 , \65830 , \65831 , \65832 , \65833 , \65834 ,
         \65835 , \65836 , \65837_nGdcc3 , \65838 , \65839 , \65840 , \65841 , \65842 , \65843 , \65844 ,
         \65845_nGda9d , \65846 , \65847 , \65848 , \65849 , \65850 , \65851 , \65852 , \65853_nGd85e , \65854 ,
         \65855 , \65856 , \65857 , \65858 , \65859 , \65860 , \65861_nGd657 , \65862 , \65863 , \65864 ,
         \65865 , \65866 , \65867 , \65868 , \65869_nGd41d , \65870 , \65871 , \65872 , \65873 , \65874 ,
         \65875 , \65876 , \65877_nGd1fd , \65878 , \65879 , \65880 , \65881 , \65882 , \65883 , \65884 ,
         \65885_nGcfa1 , \65886 , \65887 , \65888 , \65889 , \65890 , \65891 , \65892 , \65893_nGcd2c , \65894 ,
         \65895 , \65896 , \65897 , \65898 , \65899 , \65900 , \65901_nGca99 , \65902 , \65903 , \65904 ,
         \65905 , \65906 , \65907 , \65908 , \65909_nGc812 , \65910 , \65911 , \65912 , \65913 , \65914 ,
         \65915 , \65916 , \65917_nGc589 , \65918 , \65919 , \65920 , \65921 , \65922 , \65923 , \65924 ,
         \65925_nGc2e5 , \65926 , \65927 , \65928 , \65929 , \65930 , \65931 , \65932 , \65933_nGbff1 , \65934 ,
         \65935 , \65936 , \65937 , \65938 , \65939 , \65940 , \65941_nGbcf3 , \65942 , \65943 , \65944 ,
         \65945 , \65946 , \65947 , \65948 , \65949_nGba17 , \65950 , \65951 , \65952 , \65953 , \65954 ,
         \65955 , \65956 , \65957_nGb727 , \65958 , \65959 , \65960 , \65961 , \65962 , \65963 , \65964 ,
         \65965_nGb43a , \65966 , \65967 , \65968 , \65969 , \65970 , \65971 , \65972 , \65973_nGb150 , \65974 ,
         \65975 , \65976 , \65977 , \65978 , \65979 , \65980 , \65981_nGae24 , \65982 , \65983 , \65984 ,
         \65985 , \65986 , \65987 , \65988 , \65989_nGaae2 , \65990 , \65991 , \65992 , \65993 , \65994 ,
         \65995 , \65996 , \65997_nGa7c6 , \65998 , \65999 , \66000 , \66001 , \66002 , \66003 , \66004 ,
         \66005_nGa4a9 , \66006 , \66007 , \66008 , \66009 , \66010 , \66011 , \66012 , \66013_nGa14c , \66014 ,
         \66015 , \66016 , \66017 , \66018 , \66019 , \66020 , \66021_nG9ddd , \66022 , \66023 , \66024 ,
         \66025 , \66026 , \66027 , \66028 , \66029_nG9a6c , \66030 , \66031 , \66032 , \66033 , \66034 ,
         \66035 , \66036 , \66037_nG9704 , \66038 , \66039 , \66040 , \66041 , \66042 , \66043 , \66044 ,
         \66045_nG9381 , \66046 , \66047 , \66048 , \66049 , \66050 , \66051 , \66052 , \66053_nG8ff4 , \66054 ,
         \66055 , \66056 , \66057 , \66058 , \66059 , \66060 , \66061_nG8c7b , \66062 , \66063 , \66064 ,
         \66065 , \66066 , \66067 , \66068 , \66069_nG88e4 , \66070 , \66071 , \66072 , \66073 , \66074 ,
         \66075 , \66076 , \66077_nG850c , \66078 , \66079 , \66080 , \66081 , \66082 , \66083 , \66084 ,
         \66085_nG80dd , \66086 , \66087 , \66088 , \66089 , \66090 , \66091 , \66092 , \66093_nG7cf2 , \66094 ,
         \66095 , \66096 , \66097 , \66098 , \66099 , \66100 , \66101_nG7913 , \66102 , \66103 , \66104 ,
         \66105 , \66106 , \66107 , \66108 , \66109_nG7586 , \66110 , \66111 , \66112 , \66113 , \66114 ,
         \66115 , \66116 , \66117_nG7216 , \66118 , \66119 , \66120 , \66121 , \66122 , \66123 , \66124 ,
         \66125_nG6ea7 , \66126 , \66127 , \66128 , \66129 , \66130 , \66131 , \66132 , \66133_nG6b15 , \66134 ,
         \66135 , \66136 , \66137 , \66138 , \66139 , \66140 , \66141_nG6785 , \66142 , \66143 , \66144 ,
         \66145 , \66146 , \66147 , \66148 , \66149_nG642a , \66150 , \66151 , \66152 , \66153 , \66154 ,
         \66155 , \66156 , \66157_nG60ac , \66158 , \66159 , \66160 , \66161 , \66162 , \66163 , \66164 ,
         \66165_nG5d39 , \66166 , \66167 , \66168 , \66169 , \66170 , \66171 , \66172 , \66173_nG5a0d , \66174 ,
         \66175 , \66176 , \66177 , \66178 , \66179 , \66180 , \66181_nG5705 , \66182 , \66183 , \66184 ,
         \66185 , \66186 , \66187 , \66188 , \66189_nG5400 , \66190 , \66191 , \66192 , \66193 , \66194 ,
         \66195 , \66196 , \66197_nG50b7 , \66198 , \66199 , \66200 , \66201 , \66202 , \66203 , \66204 ,
         \66205_nG4d9f , \66206 , \66207 , \66208 , \66209 , \66210 , \66211 , \66212 , \66213_nG4aba , \66214 ,
         \66215 , \66216 , \66217 , \66218 , \66219 , \66220 , \66221_nG47cd , \66222 , \66223 , \66224 ,
         \66225 , \66226 , \66227 , \66228 , \66229_nG44fd , \66230 , \66231 , \66232 , \66233 , \66234 ,
         \66235 , \66236 , \66237_nG4250 , \66238 , \66239 , \66240 , \66241 , \66242 , \66243 , \66244 ,
         \66245_nG3f85 , \66246 , \66247 , \66248 , \66249 , \66250 , \66251 , \66252 , \66253_nG3cff , \66254 ,
         \66255 , \66256 , \66257 , \66258 , \66259 , \66260 , \66261_nG3a58 , \66262 , \66263 , \66264 ,
         \66265 , \66266 , \66267 , \66268 , \66269_nG37d2 , \66270 , \66271 , \66272 , \66273 , \66274 ,
         \66275 , \66276 , \66277_nG3580 , \66278 , \66279 , \66280 , \66281 , \66282 , \66283 , \66284 ,
         \66285_nG3327 , \66286 , \66287 , \66288 , \66289 , \66290 , \66291 , \66292 , \66293_nG30eb , \66294 ,
         \66295 , \66296 , \66297 , \66298 , \66299 , \66300 , \66301_nG2eb3 , \66302 , \66303 , \66304 ,
         \66305 , \66306 , \66307 , \66308 , \66309_nG2c54 , \66310 , \66311 , \66312 , \66313 , \66314 ,
         \66315 , \66316 , \66317_nG2a16 , \66318 , \66319 , \66320 , \66321 , \66322 , \66323 , \66324 ,
         \66325_nG27e2 , \66326 , \66327 , \66328 , \66329 , \66330 , \66331 , \66332 , \66333_nG25af , \66334 ,
         \66335 , \66336 , \66337 , \66338 , \66339 , \66340 , \66341_nG23ac , \66342 , \66343 , \66344 ,
         \66345 , \66346 , \66347 , \66348 , \66349_nG21c1 , \66350 , \66351 , \66352 , \66353 , \66354 ,
         \66355 , \66356 , \66357_nG1ff9 , \66358 , \66359 , \66360 , \66361 , \66362 , \66363 , \66364 ,
         \66365_nG1e19 , \66366 , \66367 , \66368 , \66369 , \66370 , \66371 , \66372 , \66373_nG1c46 , \66374 ,
         \66375 , \66376 , \66377 , \66378 , \66379 , \66380 , \66381_nG1aa2 , \66382 , \66383 , \66384 ,
         \66385 , \66386 , \66387 , \66388 , \66389_nG190e , \66390 , \66391 , \66392 , \66393 , \66394 ,
         \66395 , \66396 , \66397_nG176a , \66398 , \66399 , \66400 , \66401 , \66402 , \66403 , \66404 ,
         \66405_nG10367 , \66406 , \66407 , \66408 , \66409 , \66410 , \66411 , \66412 , \66413_nG10360 , \66414 ,
         \66415 , \66416 , \66417 , \66418 , \66419 , \66420 , \66421_nG10359 , \66422 , \66423 , \66424 ,
         \66425 , \66426 , \66427 , \66428 , \66429_nG10352 , \66430 , \66431 , \66432 , \66433 , \66434 ,
         \66435 , \66436 , \66437_nG1034b , \66438 , \66439 , \66440 , \66441 , \66442 , \66443 , \66444 ,
         \66445_nG10208 , \66446 , \66447 , \66448 , \66449 , \66450 , \66451 , \66452 , \66453_nGec84 , \66454 ,
         \66455 , \66456 , \66457 , \66458 , \66459 , \66460 , \66461_nGd865 , \66462 , \66463 , \66464 ,
         \66465 , \66466 , \66467 , \66468 , \66469_nGc819 , \66470 , \66471 , \66472 , \66473 , \66474 ,
         \66475 , \66476 , \66477_nGb441 , \66478 , \66479 , \66480 , \66481 , \66482 , \66483 , \66484 ,
         \66485_nGa4b0 , \66486 , \66487 , \66488 , \66489 , \66490 , \66491 , \66492 , \66493_nG970b , \66494 ,
         \66495 , \66496 , \66497 , \66498 , \66499 , \66500 , \66501_nG88eb , \66502 , \66503 , \66504 ,
         \66505 , \66506 , \66507 , \66508 , \66509_nG791a , \66510 , \66511 , \66512 , \66513 , \66514 ,
         \66515 , \66516 , \66517_nG6eae , \66518 , \66519 , \66520 , \66521 , \66522 , \66523 , \66524 ,
         \66525_nG6431 , \66526 ;
buf \U$labajz6697 ( R_101_77c8620, \65582 );
buf \U$labajz6698 ( R_102_af8fd30, \65590 );
buf \U$labajz6699 ( R_103_af901c8, \65598 );
buf \U$labajz6700 ( R_104_af9a140, \65606 );
buf \U$labajz6701 ( R_105_af99768, \65614 );
buf \U$labajz6702 ( R_106_af8be30, \65622 );
buf \U$labajz6703 ( R_107_77c1150, \65630 );
buf \U$labajz6704 ( R_108_af8ddb0, \65638 );
buf \U$labajz6705 ( R_109_af8f010, \65646 );
buf \U$labajz6706 ( R_10a_af996c0, \65654 );
buf \U$labajz6707 ( R_10b_77c34c0, \65662 );
buf \U$labajz6708 ( R_10c_77c28f0, \65670 );
buf \U$labajz6709 ( R_10d_af8d090, \65678 );
buf \U$labajz6710 ( R_10e_77ca5a0, \65686 );
buf \U$labajz6711 ( R_10f_77ce4a0, \65694 );
buf \U$labajz6712 ( R_110_77cd780, \65702 );
buf \U$labajz6713 ( R_111_af8f2b0, \65710 );
buf \U$labajz6714 ( R_112_77c6550, \65718 );
buf \U$labajz6715 ( R_113_af98ee0, \65726 );
buf \U$labajz6716 ( R_114_77c2068, \65734 );
buf \U$labajz6717 ( R_115_af99ea0, \65742 );
buf \U$labajz6718 ( R_116_77c0eb0, \65750 );
buf \U$labajz6719 ( R_117_77cc280, \65758 );
buf \U$labajz6720 ( R_118_77bf860, \65766 );
buf \U$labajz6721 ( R_119_77c9f10, \65774 );
buf \U$labajz6722 ( R_11a_af8bf80, \65782 );
buf \U$labajz6723 ( R_11b_77bf320, \65790 );
buf \U$labajz6724 ( R_11c_77c4fa8, \65798 );
buf \U$labajz6725 ( R_11d_af99ab0, \65806 );
buf \U$labajz6726 ( R_11e_77ca258, \65814 );
buf \U$labajz6727 ( R_11f_af92880, \65822 );
buf \U$labajz6728 ( R_120_af91c08, \65830 );
buf \U$labajz6729 ( R_121_af92298, \65838 );
buf \U$labajz6730 ( R_122_af99ca8, \65846 );
buf \U$labajz6731 ( R_123_af990d8, \65854 );
buf \U$labajz6732 ( R_124_77c5638, \65862 );
buf \U$labajz6733 ( R_125_af8e6e0, \65870 );
buf \U$labajz6734 ( R_126_77c3aa8, \65878 );
buf \U$labajz6735 ( R_127_77c8d58, \65886 );
buf \U$labajz6736 ( R_128_77c1fc0, \65894 );
buf \U$labajz6737 ( R_129_77c6748, \65902 );
buf \U$labajz6738 ( R_12a_77c3370, \65910 );
buf \U$labajz6739 ( R_12b_af99d50, \65918 );
buf \U$labajz6740 ( R_12c_77c5248, \65926 );
buf \U$labajz6741 ( R_12d_77ca840, \65934 );
buf \U$labajz6742 ( R_12e_af8eec0, \65942 );
buf \U$labajz6743 ( R_12f_77c1498, \65950 );
buf \U$labajz6744 ( R_130_77c5398, \65958 );
buf \U$labajz6745 ( R_131_77c0820, \65966 );
buf \U$labajz6746 ( R_132_af8d480, \65974 );
buf \U$labajz6747 ( R_133_77ce890, \65982 );
buf \U$labajz6748 ( R_134_af97c80, \65990 );
buf \U$labajz6749 ( R_135_77c65f8, \65998 );
buf \U$labajz6750 ( R_136_af8d678, \66006 );
buf \U$labajz6751 ( R_137_77c3e98, \66014 );
buf \U$labajz6752 ( R_138_af8e0f8, \66022 );
buf \U$labajz6753 ( R_139_af99378, \66030 );
buf \U$labajz6754 ( R_13a_77c7078, \66038 );
buf \U$labajz6755 ( R_13b_77ce740, \66046 );
buf \U$labajz6756 ( R_13c_af97fc8, \66054 );
buf \U$labajz6757 ( R_13d_77c62b0, \66062 );
buf \U$labajz6758 ( R_13e_77c27a0, \66070 );
buf \U$labajz6759 ( R_13f_af979e0, \66078 );
buf \U$labajz6760 ( R_140_77c25a8, \66086 );
buf \U$labajz6761 ( R_141_af921f0, \66094 );
buf \U$labajz6762 ( R_142_af8b7a0, \66102 );
buf \U$labajz6763 ( R_143_77bfcf8, \66110 );
buf \U$labajz6764 ( R_144_af92148, \66118 );
buf \U$labajz6765 ( R_145_77c1c78, \66126 );
buf \U$labajz6766 ( R_146_77cb560, \66134 );
buf \U$labajz6767 ( R_147_af99960, \66142 );
buf \U$labajz6768 ( R_148_af92490, \66150 );
buf \U$labajz6769 ( R_149_77c9298, \66158 );
buf \U$labajz6770 ( R_14a_77cb170, \66166 );
buf \U$labajz6771 ( R_14b_af98268, \66174 );
buf \U$labajz6772 ( R_14c_77bf9b0, \66182 );
buf \U$labajz6773 ( R_14d_af91b60, \66190 );
buf \U$labajz6774 ( R_14e_af8f208, \66198 );
buf \U$labajz6775 ( R_14f_77c7a50, \66206 );
buf \U$labajz6776 ( R_150_af99030, \66214 );
buf \U$labajz6777 ( R_151_77c67f0, \66222 );
buf \U$labajz6778 ( R_152_af8c370, \66230 );
buf \U$labajz6779 ( R_153_77c8818, \66238 );
buf \U$labajz6780 ( R_154_77c6d30, \66246 );
buf \U$labajz6781 ( R_155_af98c40, \66254 );
buf \U$labajz6782 ( R_156_77c9538, \66262 );
buf \U$labajz6783 ( R_157_af96f60, \66270 );
buf \U$labajz6784 ( R_158_af96d68, \66278 );
buf \U$labajz6785 ( R_159_af8d870, \66286 );
buf \U$labajz6786 ( R_15a_af8e830, \66294 );
buf \U$labajz6787 ( R_15b_77ccbb0, \66302 );
buf \U$labajz6788 ( R_15c_af8c610, \66310 );
buf \U$labajz6789 ( R_15d_77c6898, \66318 );
buf \U$labajz6790 ( R_15e_af8cb50, \66326 );
buf \U$labajz6791 ( R_15f_af92538, \66334 );
buf \U$labajz6792 ( R_160_af975f0, \66342 );
buf \U$labajz6793 ( R_161_77c71c8, \66350 );
buf \U$labajz6794 ( R_162_af8d720, \66358 );
buf \U$labajz6795 ( R_163_77cb608, \66366 );
buf \U$labajz6796 ( R_164_af8b650, \66374 );
buf \U$labajz6797 ( R_165_af988f8, \66382 );
buf \U$labajz6798 ( R_166_77c41e0, \66390 );
buf \U$labajz6799 ( R_167_af8e398, \66398 );
buf \U$labajz6800 ( R_168_af974a0, \66406 );
buf \U$labajz6801 ( R_169_af8d330, \66414 );
buf \U$labajz6802 ( R_16a_af8c0d0, \66422 );
buf \U$labajz6803 ( R_16b_77cc520, \66430 );
buf \U$labajz6804 ( R_16c_77cb8a8, \66438 );
buf \U$labajz6805 ( R_16d_77ccda8, \66446 );
buf \U$labajz6806 ( R_16e_af973f8, \66454 );
buf \U$labajz6807 ( R_16f_77cd6d8, \66462 );
buf \U$labajz6808 ( R_170_af99ff0, \66470 );
buf \U$labajz6809 ( R_171_77c54e8, \66478 );
buf \U$labajz6810 ( R_172_77c3808, \66486 );
buf \U$labajz6811 ( R_173_77c0580, \66494 );
buf \U$labajz6812 ( R_174_af99618, \66502 );
buf \U$labajz6813 ( R_175_77cd198, \66510 );
buf \U$labajz6814 ( R_176_77c0628, \66518 );
buf \U$labajz6815 ( R_177_af97698, \66526 );
and \U$1 ( \378 , RIae78b48_125, RIae78c38_127);
not \U$2 ( \379 , RIae78bc0_126);
and \U$3 ( \380 , \379 , RIae78c38_127);
nor \U$4 ( \381 , \379 , RIae78c38_127);
or \U$5 ( \382 , \380 , \381 );
nor \U$6 ( \383 , RIae78b48_125, RIae78c38_127);
nor \U$7 ( \384 , \378 , \382 , \383 );
nand \U$8 ( \385 , RIae78da0_130, \384 );
not \U$9 ( \386 , \385 );
nand \U$10 ( \387 , RIae78bc0_126, RIae78c38_127);
and \U$11 ( \388 , \387 , RIae78b48_125);
not \U$12 ( \389 , \388 );
and \U$13 ( \390 , \386 , \389 );
not \U$14 ( \391 , \388 );
not \U$15 ( \392 , \391 );
and \U$16 ( \393 , \385 , \392 );
nor \U$17 ( \394 , \390 , \393 );
nand \U$18 ( \395 , RIae78cb0_128, RIae78b48_125);
or \U$19 ( \396 , \394 , \395 );
nand \U$20 ( \397 , \395 , \394 );
nand \U$21 ( \398 , \396 , \397 );
nand \U$22 ( \399 , RIae78e90_132, RIae78ff8_135);
and \U$23 ( \400 , \399 , RIae78bc0_126);
not \U$24 ( \401 , \400 );
not \U$25 ( \402 , \401 );
nand \U$26 ( \403 , RIae78a58_123, RIae78b48_125);
or \U$27 ( \404 , \402 , \403 );
not \U$28 ( \405 , \403 );
not \U$29 ( \406 , \400 );
or \U$30 ( \407 , \405 , \406 );
not \U$31 ( \408 , \392 );
and \U$32 ( \409 , \384 , RIae78cb0_128);
and \U$33 ( \410 , RIae78da0_130, \382 );
nor \U$34 ( \411 , \409 , \410 );
not \U$35 ( \412 , \411 );
or \U$36 ( \413 , \408 , \412 );
or \U$37 ( \414 , \411 , \392 );
nand \U$38 ( \415 , \413 , \414 );
nand \U$39 ( \416 , \407 , \415 );
nand \U$40 ( \417 , \404 , \416 );
xor \U$41 ( \418 , \398 , \417 );
not \U$42 ( \419 , \400 );
not \U$43 ( \420 , \415 );
or \U$44 ( \421 , \419 , \420 );
or \U$45 ( \422 , \415 , \400 );
nand \U$46 ( \423 , \421 , \422 );
not \U$47 ( \424 , \423 );
not \U$48 ( \425 , \403 );
and \U$49 ( \426 , \424 , \425 );
and \U$50 ( \427 , \423 , \403 );
nor \U$51 ( \428 , \426 , \427 );
and \U$52 ( \429 , RIae78bc0_126, RIae78ff8_135);
not \U$53 ( \430 , RIae78ff8_135);
nor \U$54 ( \431 , \430 , RIae78e90_132);
not \U$55 ( \432 , RIae78e90_132);
nor \U$56 ( \433 , \432 , RIae78ff8_135);
or \U$57 ( \434 , \431 , \433 );
nor \U$58 ( \435 , RIae78bc0_126, RIae78ff8_135);
nor \U$59 ( \436 , \429 , \434 , \435 );
nand \U$60 ( \437 , RIae78da0_130, \436 );
not \U$61 ( \438 , \437 );
not \U$62 ( \439 , \402 );
and \U$63 ( \440 , \438 , \439 );
and \U$64 ( \441 , \437 , \400 );
nor \U$65 ( \442 , \440 , \441 );
nand \U$66 ( \443 , RIae76b68_57, RIae78b48_125);
xor \U$67 ( \444 , \442 , \443 );
and \U$68 ( \445 , \384 , RIae78a58_123);
and \U$69 ( \446 , RIae78cb0_128, \382 );
nor \U$70 ( \447 , \445 , \446 );
not \U$71 ( \448 , \447 );
not \U$72 ( \449 , \392 );
and \U$73 ( \450 , \448 , \449 );
and \U$74 ( \451 , \447 , \388 );
nor \U$75 ( \452 , \450 , \451 );
and \U$76 ( \453 , \444 , \452 );
and \U$77 ( \454 , \442 , \443 );
or \U$78 ( \455 , \453 , \454 );
or \U$79 ( \456 , \428 , \455 );
not \U$80 ( \457 , \455 );
not \U$81 ( \458 , \428 );
or \U$82 ( \459 , \457 , \458 );
and \U$83 ( \460 , \436 , RIae78cb0_128);
and \U$84 ( \461 , RIae78da0_130, \434 );
nor \U$85 ( \462 , \460 , \461 );
not \U$86 ( \463 , \462 );
not \U$87 ( \464 , \400 );
and \U$88 ( \465 , \463 , \464 );
and \U$89 ( \466 , \462 , \400 );
nor \U$90 ( \467 , \465 , \466 );
nand \U$91 ( \468 , RIae78f80_134, RIae78f08_133);
and \U$92 ( \469 , \468 , RIae78e90_132);
not \U$93 ( \470 , \469 );
not \U$94 ( \471 , \470 );
xor \U$95 ( \472 , \467 , \471 );
and \U$96 ( \473 , \384 , RIae76b68_57);
and \U$97 ( \474 , RIae78a58_123, \382 );
nor \U$98 ( \475 , \473 , \474 );
not \U$99 ( \476 , \475 );
not \U$100 ( \477 , \388 );
and \U$101 ( \478 , \476 , \477 );
and \U$102 ( \479 , \475 , \392 );
nor \U$103 ( \480 , \478 , \479 );
and \U$104 ( \481 , \472 , \480 );
and \U$105 ( \482 , \467 , \471 );
or \U$106 ( \483 , \481 , \482 );
xor \U$107 ( \484 , \442 , \443 );
xor \U$108 ( \485 , \484 , \452 );
nand \U$109 ( \486 , \483 , \485 );
nand \U$110 ( \487 , \459 , \486 );
nand \U$111 ( \488 , \456 , \487 );
xor \U$112 ( \489 , \418 , \488 );
not \U$113 ( \490 , RIae76988_53);
not \U$114 ( \491 , RIae78b48_125);
nor \U$115 ( \492 , \490 , \491 );
not \U$116 ( \493 , \402 );
and \U$117 ( \494 , \436 , RIae76b68_57);
and \U$118 ( \495 , RIae78a58_123, \434 );
nor \U$119 ( \496 , \494 , \495 );
not \U$120 ( \497 , \496 );
or \U$121 ( \498 , \493 , \497 );
or \U$122 ( \499 , \496 , \402 );
nand \U$123 ( \500 , \498 , \499 );
not \U$124 ( \501 , RIae79070_136);
not \U$125 ( \502 , RIae790e8_137);
or \U$126 ( \503 , \501 , \502 );
nand \U$127 ( \504 , \503 , RIae78f80_134);
xor \U$128 ( \505 , \500 , \504 );
not \U$129 ( \506 , \469 );
and \U$130 ( \507 , RIae78e90_132, RIae78f08_133);
not \U$131 ( \508 , RIae78f08_133);
nor \U$132 ( \509 , \508 , RIae78f80_134);
not \U$133 ( \510 , RIae78f80_134);
nor \U$134 ( \511 , \510 , RIae78f08_133);
or \U$135 ( \512 , \509 , \511 );
nor \U$136 ( \513 , RIae78e90_132, RIae78f08_133);
nor \U$137 ( \514 , \507 , \512 , \513 );
and \U$138 ( \515 , \514 , RIae78cb0_128);
and \U$139 ( \516 , RIae78da0_130, \512 );
nor \U$140 ( \517 , \515 , \516 );
not \U$141 ( \518 , \517 );
or \U$142 ( \519 , \506 , \518 );
or \U$143 ( \520 , \517 , \471 );
nand \U$144 ( \521 , \519 , \520 );
xor \U$145 ( \522 , \505 , \521 );
xor \U$146 ( \523 , \492 , \522 );
not \U$147 ( \524 , \523 );
nand \U$148 ( \525 , RIae76a78_55, RIae78b48_125);
and \U$149 ( \526 , \384 , RIae76988_53);
and \U$150 ( \527 , RIae767a8_49, \382 );
nor \U$151 ( \528 , \526 , \527 );
not \U$152 ( \529 , \528 );
not \U$153 ( \530 , \388 );
and \U$154 ( \531 , \529 , \530 );
and \U$155 ( \532 , \528 , \392 );
nor \U$156 ( \533 , \531 , \532 );
nand \U$157 ( \534 , \525 , \533 );
not \U$158 ( \535 , \388 );
and \U$159 ( \536 , \384 , RIae767a8_49);
and \U$160 ( \537 , RIae76898_51, \382 );
nor \U$161 ( \538 , \536 , \537 );
not \U$162 ( \539 , \538 );
or \U$163 ( \540 , \535 , \539 );
or \U$164 ( \541 , \538 , \392 );
nand \U$165 ( \542 , \540 , \541 );
xor \U$166 ( \543 , \534 , \542 );
not \U$167 ( \544 , \400 );
and \U$168 ( \545 , \436 , RIae76898_51);
and \U$169 ( \546 , RIae76b68_57, \434 );
nor \U$170 ( \547 , \545 , \546 );
not \U$171 ( \548 , \547 );
or \U$172 ( \549 , \544 , \548 );
or \U$173 ( \550 , \547 , \402 );
nand \U$174 ( \551 , \549 , \550 );
and \U$175 ( \552 , RIae78f80_134, RIae790e8_137);
not \U$176 ( \553 , RIae79070_136);
and \U$177 ( \554 , \553 , RIae790e8_137);
nor \U$178 ( \555 , \553 , RIae790e8_137);
or \U$179 ( \556 , \554 , \555 );
nor \U$180 ( \557 , RIae78f80_134, RIae790e8_137);
nor \U$181 ( \558 , \552 , \556 , \557 );
nand \U$182 ( \559 , RIae78da0_130, \558 );
and \U$183 ( \560 , \559 , \504 );
not \U$184 ( \561 , \559 );
not \U$185 ( \562 , \504 );
and \U$186 ( \563 , \561 , \562 );
nor \U$187 ( \564 , \560 , \563 );
xor \U$188 ( \565 , \551 , \564 );
not \U$189 ( \566 , \471 );
and \U$190 ( \567 , \514 , RIae78a58_123);
and \U$191 ( \568 , RIae78cb0_128, \512 );
nor \U$192 ( \569 , \567 , \568 );
not \U$193 ( \570 , \569 );
or \U$194 ( \571 , \566 , \570 );
or \U$195 ( \572 , \569 , \471 );
nand \U$196 ( \573 , \571 , \572 );
and \U$197 ( \574 , \565 , \573 );
and \U$198 ( \575 , \551 , \564 );
or \U$199 ( \576 , \574 , \575 );
xor \U$200 ( \577 , \543 , \576 );
not \U$201 ( \578 , \577 );
and \U$202 ( \579 , \558 , RIae78cb0_128);
and \U$203 ( \580 , RIae78da0_130, \556 );
nor \U$204 ( \581 , \579 , \580 );
and \U$205 ( \582 , \581 , \504 );
not \U$206 ( \583 , \581 );
and \U$207 ( \584 , \583 , \562 );
nor \U$208 ( \585 , \582 , \584 );
nand \U$209 ( \586 , RIae79160_138, RIae792c8_141);
and \U$210 ( \587 , \586 , RIae79070_136);
not \U$211 ( \588 , \587 );
xor \U$212 ( \589 , \585 , \588 );
not \U$213 ( \590 , \469 );
and \U$214 ( \591 , \514 , RIae76b68_57);
and \U$215 ( \592 , RIae78a58_123, \512 );
nor \U$216 ( \593 , \591 , \592 );
not \U$217 ( \594 , \593 );
or \U$218 ( \595 , \590 , \594 );
or \U$219 ( \596 , \593 , \471 );
nand \U$220 ( \597 , \595 , \596 );
and \U$221 ( \598 , \589 , \597 );
and \U$222 ( \599 , \585 , \588 );
or \U$223 ( \600 , \598 , \599 );
and \U$224 ( \601 , \436 , RIae767a8_49);
and \U$225 ( \602 , RIae76898_51, \434 );
nor \U$226 ( \603 , \601 , \602 );
not \U$227 ( \604 , \603 );
not \U$228 ( \605 , \400 );
and \U$229 ( \606 , \604 , \605 );
and \U$230 ( \607 , \603 , \402 );
nor \U$231 ( \608 , \606 , \607 );
nand \U$232 ( \609 , RIae76208_37, RIae78b48_125);
or \U$233 ( \610 , \608 , \609 );
not \U$234 ( \611 , \609 );
not \U$235 ( \612 , \608 );
or \U$236 ( \613 , \611 , \612 );
not \U$237 ( \614 , \388 );
and \U$238 ( \615 , \384 , RIae76a78_55);
and \U$239 ( \616 , RIae76988_53, \382 );
nor \U$240 ( \617 , \615 , \616 );
not \U$241 ( \618 , \617 );
or \U$242 ( \619 , \614 , \618 );
or \U$243 ( \620 , \617 , \388 );
nand \U$244 ( \621 , \619 , \620 );
nand \U$245 ( \622 , \613 , \621 );
nand \U$246 ( \623 , \610 , \622 );
xor \U$247 ( \624 , \600 , \623 );
or \U$248 ( \625 , \533 , \525 );
nand \U$249 ( \626 , \625 , \534 );
and \U$250 ( \627 , \624 , \626 );
and \U$251 ( \628 , \600 , \623 );
nor \U$252 ( \629 , \627 , \628 );
not \U$253 ( \630 , \629 );
and \U$254 ( \631 , \578 , \630 );
and \U$255 ( \632 , \577 , \629 );
nor \U$256 ( \633 , \631 , \632 );
not \U$257 ( \634 , \633 );
or \U$258 ( \635 , \524 , \634 );
or \U$259 ( \636 , \633 , \523 );
nand \U$260 ( \637 , \635 , \636 );
not \U$261 ( \638 , \637 );
xor \U$262 ( \639 , \600 , \623 );
xor \U$263 ( \640 , \639 , \626 );
xor \U$264 ( \641 , \551 , \564 );
xor \U$265 ( \642 , \641 , \573 );
and \U$266 ( \643 , \640 , \642 );
not \U$267 ( \644 , \640 );
not \U$268 ( \645 , \642 );
and \U$269 ( \646 , \644 , \645 );
not \U$270 ( \647 , \608 );
not \U$271 ( \648 , \621 );
or \U$272 ( \649 , \647 , \648 );
or \U$273 ( \650 , \608 , \621 );
nand \U$274 ( \651 , \649 , \650 );
not \U$275 ( \652 , \651 );
not \U$276 ( \653 , \609 );
and \U$277 ( \654 , \652 , \653 );
and \U$278 ( \655 , \651 , \609 );
nor \U$279 ( \656 , \654 , \655 );
not \U$280 ( \657 , \656 );
and \U$281 ( \658 , \514 , RIae76898_51);
and \U$282 ( \659 , RIae76b68_57, \512 );
nor \U$283 ( \660 , \658 , \659 );
not \U$284 ( \661 , \660 );
not \U$285 ( \662 , \469 );
and \U$286 ( \663 , \661 , \662 );
and \U$287 ( \664 , \660 , \471 );
nor \U$288 ( \665 , \663 , \664 );
and \U$289 ( \666 , RIae79070_136, RIae792c8_141);
not \U$290 ( \667 , RIae79160_138);
and \U$291 ( \668 , \667 , RIae792c8_141);
nor \U$292 ( \669 , \667 , RIae792c8_141);
or \U$293 ( \670 , \668 , \669 );
nor \U$294 ( \671 , RIae79070_136, RIae792c8_141);
nor \U$295 ( \672 , \666 , \670 , \671 );
nand \U$296 ( \673 , RIae78da0_130, \672 );
and \U$297 ( \674 , \673 , \587 );
not \U$298 ( \675 , \673 );
and \U$299 ( \676 , \675 , \588 );
nor \U$300 ( \677 , \674 , \676 );
xor \U$301 ( \678 , \665 , \677 );
and \U$302 ( \679 , \558 , RIae78a58_123);
and \U$303 ( \680 , RIae78cb0_128, \556 );
nor \U$304 ( \681 , \679 , \680 );
and \U$305 ( \682 , \681 , \562 );
not \U$306 ( \683 , \681 );
and \U$307 ( \684 , \683 , \504 );
nor \U$308 ( \685 , \682 , \684 );
and \U$309 ( \686 , \678 , \685 );
and \U$310 ( \687 , \665 , \677 );
or \U$311 ( \688 , \686 , \687 );
not \U$312 ( \689 , \688 );
and \U$313 ( \690 , \657 , \689 );
and \U$314 ( \691 , \656 , \688 );
and \U$315 ( \692 , \384 , RIae76208_37);
and \U$316 ( \693 , RIae76a78_55, \382 );
nor \U$317 ( \694 , \692 , \693 );
not \U$318 ( \695 , \694 );
not \U$319 ( \696 , \388 );
and \U$320 ( \697 , \695 , \696 );
and \U$321 ( \698 , \694 , \392 );
nor \U$322 ( \699 , \697 , \698 );
nand \U$323 ( \700 , RIae762f8_39, RIae78b48_125);
xor \U$324 ( \701 , \699 , \700 );
and \U$325 ( \702 , \436 , RIae76988_53);
and \U$326 ( \703 , RIae767a8_49, \434 );
nor \U$327 ( \704 , \702 , \703 );
not \U$328 ( \705 , \704 );
not \U$329 ( \706 , \402 );
and \U$330 ( \707 , \705 , \706 );
and \U$331 ( \708 , \704 , \402 );
nor \U$332 ( \709 , \707 , \708 );
and \U$333 ( \710 , \701 , \709 );
and \U$334 ( \711 , \699 , \700 );
or \U$335 ( \712 , \710 , \711 );
nor \U$336 ( \713 , \691 , \712 );
nor \U$337 ( \714 , \690 , \713 );
nor \U$338 ( \715 , \646 , \714 );
nor \U$339 ( \716 , \643 , \715 );
nor \U$340 ( \717 , \638 , \716 );
and \U$341 ( \718 , \492 , \522 );
xor \U$342 ( \719 , \534 , \542 );
and \U$343 ( \720 , \719 , \576 );
and \U$344 ( \721 , \534 , \542 );
or \U$345 ( \722 , \720 , \721 );
xor \U$346 ( \723 , \718 , \722 );
xor \U$347 ( \724 , \500 , \504 );
and \U$348 ( \725 , \724 , \521 );
and \U$349 ( \726 , \500 , \504 );
or \U$350 ( \727 , \725 , \726 );
nand \U$351 ( \728 , RIae767a8_49, RIae78b48_125);
xor \U$352 ( \729 , \727 , \728 );
not \U$353 ( \730 , \392 );
and \U$354 ( \731 , \384 , RIae76898_51);
and \U$355 ( \732 , RIae76b68_57, \382 );
nor \U$356 ( \733 , \731 , \732 );
not \U$357 ( \734 , \733 );
or \U$358 ( \735 , \730 , \734 );
or \U$359 ( \736 , \733 , \388 );
nand \U$360 ( \737 , \735 , \736 );
not \U$361 ( \738 , \469 );
nand \U$362 ( \739 , RIae78da0_130, \514 );
not \U$363 ( \740 , \739 );
or \U$364 ( \741 , \738 , \740 );
or \U$365 ( \742 , \739 , \471 );
nand \U$366 ( \743 , \741 , \742 );
xor \U$367 ( \744 , \737 , \743 );
not \U$368 ( \745 , \400 );
and \U$369 ( \746 , \436 , RIae78a58_123);
and \U$370 ( \747 , RIae78cb0_128, \434 );
nor \U$371 ( \748 , \746 , \747 );
not \U$372 ( \749 , \748 );
or \U$373 ( \750 , \745 , \749 );
or \U$374 ( \751 , \748 , \402 );
nand \U$375 ( \752 , \750 , \751 );
xor \U$376 ( \753 , \744 , \752 );
xor \U$377 ( \754 , \729 , \753 );
xor \U$378 ( \755 , \723 , \754 );
not \U$379 ( \756 , \755 );
and \U$380 ( \757 , \577 , \523 );
not \U$381 ( \758 , \577 );
not \U$382 ( \759 , \523 );
and \U$383 ( \760 , \758 , \759 );
nor \U$384 ( \761 , \760 , \629 );
nor \U$385 ( \762 , \757 , \761 );
not \U$386 ( \763 , \762 );
or \U$387 ( \764 , \756 , \763 );
or \U$388 ( \765 , \762 , \755 );
nand \U$389 ( \766 , \764 , \765 );
and \U$390 ( \767 , \717 , \766 );
xor \U$391 ( \768 , \717 , \766 );
not \U$392 ( \769 , \640 );
not \U$393 ( \770 , \714 );
not \U$394 ( \771 , \642 );
and \U$395 ( \772 , \770 , \771 );
and \U$396 ( \773 , \714 , \642 );
nor \U$397 ( \774 , \772 , \773 );
not \U$398 ( \775 , \774 );
or \U$399 ( \776 , \769 , \775 );
or \U$400 ( \777 , \774 , \640 );
nand \U$401 ( \778 , \776 , \777 );
and \U$402 ( \779 , \672 , RIae78cb0_128);
and \U$403 ( \780 , RIae78da0_130, \670 );
nor \U$404 ( \781 , \779 , \780 );
and \U$405 ( \782 , \781 , \587 );
not \U$406 ( \783 , \781 );
and \U$407 ( \784 , \783 , \588 );
nor \U$408 ( \785 , \782 , \784 );
nand \U$409 ( \786 , RIae79250_140, RIae791d8_139);
and \U$410 ( \787 , \786 , RIae79160_138);
not \U$411 ( \788 , \787 );
not \U$412 ( \789 , \788 );
xor \U$413 ( \790 , \785 , \789 );
and \U$414 ( \791 , \558 , RIae76b68_57);
and \U$415 ( \792 , RIae78a58_123, \556 );
nor \U$416 ( \793 , \791 , \792 );
and \U$417 ( \794 , \793 , \562 );
not \U$418 ( \795 , \793 );
and \U$419 ( \796 , \795 , \504 );
nor \U$420 ( \797 , \794 , \796 );
and \U$421 ( \798 , \790 , \797 );
and \U$422 ( \799 , \785 , \789 );
or \U$423 ( \800 , \798 , \799 );
and \U$424 ( \801 , \384 , RIae762f8_39);
and \U$425 ( \802 , RIae76208_37, \382 );
nor \U$426 ( \803 , \801 , \802 );
not \U$427 ( \804 , \803 );
not \U$428 ( \805 , \392 );
and \U$429 ( \806 , \804 , \805 );
and \U$430 ( \807 , \803 , \392 );
nor \U$431 ( \808 , \806 , \807 );
and \U$432 ( \809 , \436 , RIae76a78_55);
and \U$433 ( \810 , RIae76988_53, \434 );
nor \U$434 ( \811 , \809 , \810 );
not \U$435 ( \812 , \811 );
not \U$436 ( \813 , \402 );
and \U$437 ( \814 , \812 , \813 );
and \U$438 ( \815 , \811 , \402 );
nor \U$439 ( \816 , \814 , \815 );
xor \U$440 ( \817 , \808 , \816 );
and \U$441 ( \818 , \514 , RIae767a8_49);
and \U$442 ( \819 , RIae76898_51, \512 );
nor \U$443 ( \820 , \818 , \819 );
not \U$444 ( \821 , \820 );
not \U$445 ( \822 , \469 );
and \U$446 ( \823 , \821 , \822 );
and \U$447 ( \824 , \820 , \469 );
nor \U$448 ( \825 , \823 , \824 );
and \U$449 ( \826 , \817 , \825 );
and \U$450 ( \827 , \808 , \816 );
or \U$451 ( \828 , \826 , \827 );
nand \U$452 ( \829 , \800 , \828 );
xor \U$453 ( \830 , \585 , \588 );
xor \U$454 ( \831 , \830 , \597 );
xor \U$455 ( \832 , \829 , \831 );
not \U$456 ( \833 , \656 );
xor \U$457 ( \834 , \712 , \688 );
not \U$458 ( \835 , \834 );
or \U$459 ( \836 , \833 , \835 );
or \U$460 ( \837 , \834 , \656 );
nand \U$461 ( \838 , \836 , \837 );
and \U$462 ( \839 , \832 , \838 );
and \U$463 ( \840 , \829 , \831 );
or \U$464 ( \841 , \839 , \840 );
and \U$465 ( \842 , \778 , \841 );
not \U$466 ( \843 , \778 );
not \U$467 ( \844 , \841 );
and \U$468 ( \845 , \843 , \844 );
xor \U$469 ( \846 , \829 , \831 );
xor \U$470 ( \847 , \846 , \838 );
or \U$471 ( \848 , \828 , \800 );
nand \U$472 ( \849 , \848 , \829 );
not \U$473 ( \850 , \849 );
xor \U$474 ( \851 , \665 , \677 );
xor \U$475 ( \852 , \851 , \685 );
nor \U$476 ( \853 , \850 , \852 );
and \U$477 ( \854 , \847 , \853 );
not \U$478 ( \855 , \847 );
not \U$479 ( \856 , \853 );
and \U$480 ( \857 , \855 , \856 );
and \U$481 ( \858 , \558 , RIae76898_51);
and \U$482 ( \859 , RIae76b68_57, \556 );
nor \U$483 ( \860 , \858 , \859 );
and \U$484 ( \861 , \860 , \562 );
not \U$485 ( \862 , \860 );
and \U$486 ( \863 , \862 , \504 );
nor \U$487 ( \864 , \861 , \863 );
not \U$488 ( \865 , \864 );
and \U$489 ( \866 , \672 , RIae78a58_123);
and \U$490 ( \867 , RIae78cb0_128, \670 );
nor \U$491 ( \868 , \866 , \867 );
and \U$492 ( \869 , \868 , \587 );
not \U$493 ( \870 , \868 );
and \U$494 ( \871 , \870 , \588 );
nor \U$495 ( \872 , \869 , \871 );
not \U$496 ( \873 , \872 );
and \U$497 ( \874 , \865 , \873 );
and \U$498 ( \875 , \872 , \864 );
and \U$499 ( \876 , RIae79160_138, RIae791d8_139);
not \U$500 ( \877 , RIae791d8_139);
nor \U$501 ( \878 , \877 , RIae79250_140);
not \U$502 ( \879 , RIae79250_140);
nor \U$503 ( \880 , \879 , RIae791d8_139);
or \U$504 ( \881 , \878 , \880 );
nor \U$505 ( \882 , RIae79160_138, RIae791d8_139);
nor \U$506 ( \883 , \876 , \881 , \882 );
nand \U$507 ( \884 , RIae78da0_130, \883 );
not \U$508 ( \885 , \884 );
not \U$509 ( \886 , \787 );
and \U$510 ( \887 , \885 , \886 );
and \U$511 ( \888 , \884 , \789 );
nor \U$512 ( \889 , \887 , \888 );
nor \U$513 ( \890 , \875 , \889 );
nor \U$514 ( \891 , \874 , \890 );
nand \U$515 ( \892 , RIae76118_35, RIae78b48_125);
xor \U$516 ( \893 , \891 , \892 );
and \U$517 ( \894 , \384 , RIae76028_33);
and \U$518 ( \895 , RIae762f8_39, \382 );
nor \U$519 ( \896 , \894 , \895 );
not \U$520 ( \897 , \896 );
not \U$521 ( \898 , \388 );
and \U$522 ( \899 , \897 , \898 );
and \U$523 ( \900 , \896 , \392 );
nor \U$524 ( \901 , \899 , \900 );
not \U$525 ( \902 , \901 );
and \U$526 ( \903 , \514 , RIae76988_53);
and \U$527 ( \904 , RIae767a8_49, \512 );
nor \U$528 ( \905 , \903 , \904 );
not \U$529 ( \906 , \905 );
not \U$530 ( \907 , \469 );
and \U$531 ( \908 , \906 , \907 );
and \U$532 ( \909 , \905 , \471 );
nor \U$533 ( \910 , \908 , \909 );
not \U$534 ( \911 , \910 );
and \U$535 ( \912 , \902 , \911 );
and \U$536 ( \913 , \910 , \901 );
and \U$537 ( \914 , \436 , RIae76208_37);
and \U$538 ( \915 , RIae76a78_55, \434 );
nor \U$539 ( \916 , \914 , \915 );
not \U$540 ( \917 , \916 );
not \U$541 ( \918 , \400 );
and \U$542 ( \919 , \917 , \918 );
and \U$543 ( \920 , \916 , \402 );
nor \U$544 ( \921 , \919 , \920 );
nor \U$545 ( \922 , \913 , \921 );
nor \U$546 ( \923 , \912 , \922 );
and \U$547 ( \924 , \893 , \923 );
and \U$548 ( \925 , \891 , \892 );
or \U$549 ( \926 , \924 , \925 );
xor \U$550 ( \927 , \699 , \700 );
xor \U$551 ( \928 , \927 , \709 );
xor \U$552 ( \929 , \926 , \928 );
xor \U$553 ( \930 , \785 , \789 );
xor \U$554 ( \931 , \930 , \797 );
not \U$555 ( \932 , \931 );
nand \U$556 ( \933 , RIae76028_33, RIae78b48_125);
not \U$557 ( \934 , \933 );
and \U$558 ( \935 , \932 , \934 );
and \U$559 ( \936 , \931 , \933 );
xor \U$560 ( \937 , \808 , \816 );
xor \U$561 ( \938 , \937 , \825 );
nor \U$562 ( \939 , \936 , \938 );
nor \U$563 ( \940 , \935 , \939 );
and \U$564 ( \941 , \929 , \940 );
and \U$565 ( \942 , \926 , \928 );
or \U$566 ( \943 , \941 , \942 );
nor \U$567 ( \944 , \857 , \943 );
nor \U$568 ( \945 , \854 , \944 );
nor \U$569 ( \946 , \845 , \945 );
nor \U$570 ( \947 , \842 , \946 );
not \U$571 ( \948 , \637 );
not \U$572 ( \949 , \716 );
and \U$573 ( \950 , \948 , \949 );
and \U$574 ( \951 , \637 , \716 );
nor \U$575 ( \952 , \950 , \951 );
or \U$576 ( \953 , \947 , \952 );
xnor \U$577 ( \954 , \952 , \947 );
not \U$578 ( \955 , \778 );
not \U$579 ( \956 , \945 );
not \U$580 ( \957 , \841 );
and \U$581 ( \958 , \956 , \957 );
and \U$582 ( \959 , \945 , \841 );
nor \U$583 ( \960 , \958 , \959 );
not \U$584 ( \961 , \960 );
or \U$585 ( \962 , \955 , \961 );
or \U$586 ( \963 , \960 , \778 );
nand \U$587 ( \964 , \962 , \963 );
not \U$588 ( \965 , \847 );
not \U$589 ( \966 , \943 );
not \U$590 ( \967 , \853 );
and \U$591 ( \968 , \966 , \967 );
and \U$592 ( \969 , \943 , \853 );
nor \U$593 ( \970 , \968 , \969 );
not \U$594 ( \971 , \970 );
or \U$595 ( \972 , \965 , \971 );
or \U$596 ( \973 , \970 , \847 );
nand \U$597 ( \974 , \972 , \973 );
xor \U$598 ( \975 , \926 , \928 );
xor \U$599 ( \976 , \975 , \940 );
not \U$600 ( \977 , \849 );
not \U$601 ( \978 , \852 );
and \U$602 ( \979 , \977 , \978 );
and \U$603 ( \980 , \849 , \852 );
nor \U$604 ( \981 , \979 , \980 );
or \U$605 ( \982 , \976 , \981 );
not \U$606 ( \983 , \981 );
not \U$607 ( \984 , \976 );
or \U$608 ( \985 , \983 , \984 );
not \U$609 ( \986 , \901 );
xor \U$610 ( \987 , \921 , \910 );
not \U$611 ( \988 , \987 );
or \U$612 ( \989 , \986 , \988 );
or \U$613 ( \990 , \987 , \901 );
nand \U$614 ( \991 , \989 , \990 );
xor \U$615 ( \992 , \991 , \892 );
not \U$616 ( \993 , \864 );
xor \U$617 ( \994 , \889 , \872 );
not \U$618 ( \995 , \994 );
or \U$619 ( \996 , \993 , \995 );
or \U$620 ( \997 , \994 , \864 );
nand \U$621 ( \998 , \996 , \997 );
and \U$622 ( \999 , \992 , \998 );
and \U$623 ( \1000 , \991 , \892 );
or \U$624 ( \1001 , \999 , \1000 );
and \U$625 ( \1002 , \672 , RIae76b68_57);
and \U$626 ( \1003 , RIae78a58_123, \670 );
nor \U$627 ( \1004 , \1002 , \1003 );
and \U$628 ( \1005 , \1004 , \588 );
not \U$629 ( \1006 , \1004 );
and \U$630 ( \1007 , \1006 , \587 );
nor \U$631 ( \1008 , \1005 , \1007 );
not \U$632 ( \1009 , RIae793b8_143);
not \U$633 ( \1010 , RIae79340_142);
or \U$634 ( \1011 , \1009 , \1010 );
nand \U$635 ( \1012 , \1011 , RIae79250_140);
xor \U$636 ( \1013 , \1008 , \1012 );
not \U$637 ( \1014 , \787 );
and \U$638 ( \1015 , \883 , RIae78cb0_128);
and \U$639 ( \1016 , RIae78da0_130, \881 );
nor \U$640 ( \1017 , \1015 , \1016 );
not \U$641 ( \1018 , \1017 );
or \U$642 ( \1019 , \1014 , \1018 );
or \U$643 ( \1020 , \1017 , \787 );
nand \U$644 ( \1021 , \1019 , \1020 );
and \U$645 ( \1022 , \1013 , \1021 );
and \U$646 ( \1023 , \1008 , \1012 );
or \U$647 ( \1024 , \1022 , \1023 );
not \U$648 ( \1025 , RIae765c8_45);
nor \U$649 ( \1026 , \1025 , \491 );
not \U$650 ( \1027 , \388 );
and \U$651 ( \1028 , \384 , RIae76118_35);
and \U$652 ( \1029 , RIae76028_33, \382 );
nor \U$653 ( \1030 , \1028 , \1029 );
not \U$654 ( \1031 , \1030 );
or \U$655 ( \1032 , \1027 , \1031 );
or \U$656 ( \1033 , \1030 , \388 );
nand \U$657 ( \1034 , \1032 , \1033 );
and \U$658 ( \1035 , \1026 , \1034 );
xor \U$659 ( \1036 , \1024 , \1035 );
not \U$660 ( \1037 , \471 );
and \U$661 ( \1038 , \514 , RIae76a78_55);
and \U$662 ( \1039 , RIae76988_53, \512 );
nor \U$663 ( \1040 , \1038 , \1039 );
not \U$664 ( \1041 , \1040 );
or \U$665 ( \1042 , \1037 , \1041 );
or \U$666 ( \1043 , \1040 , \469 );
nand \U$667 ( \1044 , \1042 , \1043 );
not \U$668 ( \1045 , \400 );
and \U$669 ( \1046 , \436 , RIae762f8_39);
and \U$670 ( \1047 , RIae76208_37, \434 );
nor \U$671 ( \1048 , \1046 , \1047 );
not \U$672 ( \1049 , \1048 );
or \U$673 ( \1050 , \1045 , \1049 );
or \U$674 ( \1051 , \1048 , \402 );
nand \U$675 ( \1052 , \1050 , \1051 );
xor \U$676 ( \1053 , \1044 , \1052 );
and \U$677 ( \1054 , \558 , RIae767a8_49);
and \U$678 ( \1055 , RIae76898_51, \556 );
nor \U$679 ( \1056 , \1054 , \1055 );
and \U$680 ( \1057 , \1056 , \504 );
not \U$681 ( \1058 , \1056 );
and \U$682 ( \1059 , \1058 , \562 );
nor \U$683 ( \1060 , \1057 , \1059 );
and \U$684 ( \1061 , \1053 , \1060 );
and \U$685 ( \1062 , \1044 , \1052 );
or \U$686 ( \1063 , \1061 , \1062 );
and \U$687 ( \1064 , \1036 , \1063 );
and \U$688 ( \1065 , \1024 , \1035 );
or \U$689 ( \1066 , \1064 , \1065 );
xor \U$690 ( \1067 , \1001 , \1066 );
not \U$691 ( \1068 , \931 );
xor \U$692 ( \1069 , \933 , \938 );
not \U$693 ( \1070 , \1069 );
or \U$694 ( \1071 , \1068 , \1070 );
or \U$695 ( \1072 , \1069 , \931 );
nand \U$696 ( \1073 , \1071 , \1072 );
and \U$697 ( \1074 , \1067 , \1073 );
and \U$698 ( \1075 , \1001 , \1066 );
or \U$699 ( \1076 , \1074 , \1075 );
nand \U$700 ( \1077 , \985 , \1076 );
nand \U$701 ( \1078 , \982 , \1077 );
and \U$702 ( \1079 , \974 , \1078 );
and \U$703 ( \1080 , \964 , \1079 );
xor \U$704 ( \1081 , \1079 , \964 );
not \U$705 ( \1082 , \1076 );
not \U$706 ( \1083 , \976 );
or \U$707 ( \1084 , \1082 , \1083 );
or \U$708 ( \1085 , \976 , \1076 );
nand \U$709 ( \1086 , \1084 , \1085 );
not \U$710 ( \1087 , \1086 );
not \U$711 ( \1088 , \981 );
and \U$712 ( \1089 , \1087 , \1088 );
and \U$713 ( \1090 , \1086 , \981 );
nor \U$714 ( \1091 , \1089 , \1090 );
not \U$715 ( \1092 , \1091 );
xor \U$716 ( \1093 , \1001 , \1066 );
xor \U$717 ( \1094 , \1093 , \1073 );
not \U$718 ( \1095 , \1094 );
xor \U$719 ( \1096 , \891 , \892 );
xor \U$720 ( \1097 , \1096 , \923 );
or \U$721 ( \1098 , \1095 , \1097 );
not \U$722 ( \1099 , \1097 );
not \U$723 ( \1100 , \1095 );
or \U$724 ( \1101 , \1099 , \1100 );
xor \U$725 ( \1102 , \1026 , \1034 );
xor \U$726 ( \1103 , \1008 , \1012 );
xor \U$727 ( \1104 , \1103 , \1021 );
and \U$728 ( \1105 , \1102 , \1104 );
xor \U$729 ( \1106 , \1044 , \1052 );
xor \U$730 ( \1107 , \1106 , \1060 );
xor \U$731 ( \1108 , \1008 , \1012 );
xor \U$732 ( \1109 , \1108 , \1021 );
and \U$733 ( \1110 , \1107 , \1109 );
and \U$734 ( \1111 , \1102 , \1107 );
or \U$735 ( \1112 , \1105 , \1110 , \1111 );
and \U$736 ( \1113 , \672 , RIae76898_51);
and \U$737 ( \1114 , RIae76b68_57, \670 );
nor \U$738 ( \1115 , \1113 , \1114 );
and \U$739 ( \1116 , \1115 , \587 );
not \U$740 ( \1117 , \1115 );
and \U$741 ( \1118 , \1117 , \588 );
nor \U$742 ( \1119 , \1116 , \1118 );
and \U$743 ( \1120 , \883 , RIae78a58_123);
and \U$744 ( \1121 , RIae78cb0_128, \881 );
nor \U$745 ( \1122 , \1120 , \1121 );
not \U$746 ( \1123 , \1122 );
not \U$747 ( \1124 , \789 );
and \U$748 ( \1125 , \1123 , \1124 );
and \U$749 ( \1126 , \1122 , \787 );
nor \U$750 ( \1127 , \1125 , \1126 );
or \U$751 ( \1128 , \1119 , \1127 );
not \U$752 ( \1129 , \1127 );
not \U$753 ( \1130 , \1119 );
or \U$754 ( \1131 , \1129 , \1130 );
and \U$755 ( \1132 , RIae79250_140, RIae79340_142);
not \U$756 ( \1133 , RIae793b8_143);
and \U$757 ( \1134 , \1133 , RIae79340_142);
nor \U$758 ( \1135 , \1133 , RIae79340_142);
or \U$759 ( \1136 , \1134 , \1135 );
nor \U$760 ( \1137 , RIae79250_140, RIae79340_142);
nor \U$761 ( \1138 , \1132 , \1136 , \1137 );
nand \U$762 ( \1139 , RIae78da0_130, \1138 );
and \U$763 ( \1140 , \1139 , \1012 );
not \U$764 ( \1141 , \1139 );
not \U$765 ( \1142 , \1012 );
and \U$766 ( \1143 , \1141 , \1142 );
nor \U$767 ( \1144 , \1140 , \1143 );
nand \U$768 ( \1145 , \1131 , \1144 );
nand \U$769 ( \1146 , \1128 , \1145 );
nand \U$770 ( \1147 , RIae766b8_47, RIae78b48_125);
and \U$771 ( \1148 , \384 , RIae765c8_45);
and \U$772 ( \1149 , RIae76118_35, \382 );
nor \U$773 ( \1150 , \1148 , \1149 );
not \U$774 ( \1151 , \1150 );
not \U$775 ( \1152 , \392 );
and \U$776 ( \1153 , \1151 , \1152 );
and \U$777 ( \1154 , \1150 , \388 );
nor \U$778 ( \1155 , \1153 , \1154 );
nand \U$779 ( \1156 , \1147 , \1155 );
xor \U$780 ( \1157 , \1146 , \1156 );
and \U$781 ( \1158 , \514 , RIae76208_37);
and \U$782 ( \1159 , RIae76a78_55, \512 );
nor \U$783 ( \1160 , \1158 , \1159 );
not \U$784 ( \1161 , \1160 );
not \U$785 ( \1162 , \469 );
and \U$786 ( \1163 , \1161 , \1162 );
and \U$787 ( \1164 , \1160 , \471 );
nor \U$788 ( \1165 , \1163 , \1164 );
and \U$789 ( \1166 , \558 , RIae76988_53);
and \U$790 ( \1167 , RIae767a8_49, \556 );
nor \U$791 ( \1168 , \1166 , \1167 );
and \U$792 ( \1169 , \1168 , \562 );
not \U$793 ( \1170 , \1168 );
and \U$794 ( \1171 , \1170 , \504 );
nor \U$795 ( \1172 , \1169 , \1171 );
xor \U$796 ( \1173 , \1165 , \1172 );
and \U$797 ( \1174 , \436 , RIae76028_33);
and \U$798 ( \1175 , RIae762f8_39, \434 );
nor \U$799 ( \1176 , \1174 , \1175 );
not \U$800 ( \1177 , \1176 );
not \U$801 ( \1178 , \402 );
and \U$802 ( \1179 , \1177 , \1178 );
and \U$803 ( \1180 , \1176 , \402 );
nor \U$804 ( \1181 , \1179 , \1180 );
and \U$805 ( \1182 , \1173 , \1181 );
and \U$806 ( \1183 , \1165 , \1172 );
nor \U$807 ( \1184 , \1182 , \1183 );
and \U$808 ( \1185 , \1157 , \1184 );
and \U$809 ( \1186 , \1146 , \1156 );
or \U$810 ( \1187 , \1185 , \1186 );
xor \U$811 ( \1188 , \1112 , \1187 );
xor \U$812 ( \1189 , \991 , \892 );
xor \U$813 ( \1190 , \1189 , \998 );
and \U$814 ( \1191 , \1188 , \1190 );
and \U$815 ( \1192 , \1112 , \1187 );
or \U$816 ( \1193 , \1191 , \1192 );
nand \U$817 ( \1194 , \1101 , \1193 );
nand \U$818 ( \1195 , \1098 , \1194 );
not \U$819 ( \1196 , \1195 );
and \U$820 ( \1197 , \1092 , \1196 );
and \U$821 ( \1198 , \1091 , \1195 );
nor \U$822 ( \1199 , \1197 , \1198 );
not \U$823 ( \1200 , \1193 );
not \U$824 ( \1201 , \1097 );
and \U$825 ( \1202 , \1200 , \1201 );
and \U$826 ( \1203 , \1193 , \1097 );
nor \U$827 ( \1204 , \1202 , \1203 );
not \U$828 ( \1205 , \1204 );
not \U$829 ( \1206 , \1094 );
and \U$830 ( \1207 , \1205 , \1206 );
and \U$831 ( \1208 , \1204 , \1094 );
nor \U$832 ( \1209 , \1207 , \1208 );
not \U$833 ( \1210 , \1209 );
not \U$834 ( \1211 , \1144 );
not \U$835 ( \1212 , \1127 );
or \U$836 ( \1213 , \1211 , \1212 );
or \U$837 ( \1214 , \1127 , \1144 );
nand \U$838 ( \1215 , \1213 , \1214 );
not \U$839 ( \1216 , \1215 );
not \U$840 ( \1217 , \1119 );
and \U$841 ( \1218 , \1216 , \1217 );
and \U$842 ( \1219 , \1215 , \1119 );
nor \U$843 ( \1220 , \1218 , \1219 );
xor \U$844 ( \1221 , \1165 , \1172 );
xor \U$845 ( \1222 , \1221 , \1181 );
or \U$846 ( \1223 , \1220 , \1222 );
not \U$847 ( \1224 , \1222 );
not \U$848 ( \1225 , \1220 );
or \U$849 ( \1226 , \1224 , \1225 );
or \U$850 ( \1227 , \1155 , \1147 );
nand \U$851 ( \1228 , \1227 , \1156 );
nand \U$852 ( \1229 , \1226 , \1228 );
nand \U$853 ( \1230 , \1223 , \1229 );
and \U$854 ( \1231 , \436 , RIae76118_35);
and \U$855 ( \1232 , RIae76028_33, \434 );
nor \U$856 ( \1233 , \1231 , \1232 );
not \U$857 ( \1234 , \1233 );
not \U$858 ( \1235 , \400 );
and \U$859 ( \1236 , \1234 , \1235 );
and \U$860 ( \1237 , \1233 , \402 );
nor \U$861 ( \1238 , \1236 , \1237 );
nand \U$862 ( \1239 , RIae764d8_43, RIae78b48_125);
xor \U$863 ( \1240 , \1238 , \1239 );
and \U$864 ( \1241 , \384 , RIae766b8_47);
and \U$865 ( \1242 , RIae765c8_45, \382 );
nor \U$866 ( \1243 , \1241 , \1242 );
not \U$867 ( \1244 , \1243 );
not \U$868 ( \1245 , \388 );
and \U$869 ( \1246 , \1244 , \1245 );
and \U$870 ( \1247 , \1243 , \388 );
nor \U$871 ( \1248 , \1246 , \1247 );
and \U$872 ( \1249 , \1240 , \1248 );
and \U$873 ( \1250 , \1238 , \1239 );
or \U$874 ( \1251 , \1249 , \1250 );
and \U$875 ( \1252 , \883 , RIae76b68_57);
and \U$876 ( \1253 , RIae78a58_123, \881 );
nor \U$877 ( \1254 , \1252 , \1253 );
not \U$878 ( \1255 , \1254 );
not \U$879 ( \1256 , \789 );
and \U$880 ( \1257 , \1255 , \1256 );
and \U$881 ( \1258 , \1254 , \787 );
nor \U$882 ( \1259 , \1257 , \1258 );
nand \U$883 ( \1260 , RIae79610_148, RIae799d0_156);
and \U$884 ( \1261 , \1260 , RIae793b8_143);
xor \U$885 ( \1262 , \1259 , \1261 );
and \U$886 ( \1263 , \1138 , RIae78cb0_128);
and \U$887 ( \1264 , RIae78da0_130, \1136 );
nor \U$888 ( \1265 , \1263 , \1264 );
and \U$889 ( \1266 , \1265 , \1142 );
not \U$890 ( \1267 , \1265 );
and \U$891 ( \1268 , \1267 , \1012 );
nor \U$892 ( \1269 , \1266 , \1268 );
and \U$893 ( \1270 , \1262 , \1269 );
and \U$894 ( \1271 , \1259 , \1261 );
or \U$895 ( \1272 , \1270 , \1271 );
xor \U$896 ( \1273 , \1251 , \1272 );
and \U$897 ( \1274 , \558 , RIae76a78_55);
and \U$898 ( \1275 , RIae76988_53, \556 );
nor \U$899 ( \1276 , \1274 , \1275 );
and \U$900 ( \1277 , \1276 , \562 );
not \U$901 ( \1278 , \1276 );
and \U$902 ( \1279 , \1278 , \504 );
nor \U$903 ( \1280 , \1277 , \1279 );
and \U$904 ( \1281 , \514 , RIae762f8_39);
and \U$905 ( \1282 , RIae76208_37, \512 );
nor \U$906 ( \1283 , \1281 , \1282 );
not \U$907 ( \1284 , \1283 );
not \U$908 ( \1285 , \471 );
and \U$909 ( \1286 , \1284 , \1285 );
and \U$910 ( \1287 , \1283 , \471 );
nor \U$911 ( \1288 , \1286 , \1287 );
xor \U$912 ( \1289 , \1280 , \1288 );
and \U$913 ( \1290 , \672 , RIae767a8_49);
and \U$914 ( \1291 , RIae76898_51, \670 );
nor \U$915 ( \1292 , \1290 , \1291 );
and \U$916 ( \1293 , \1292 , \587 );
not \U$917 ( \1294 , \1292 );
and \U$918 ( \1295 , \1294 , \588 );
nor \U$919 ( \1296 , \1293 , \1295 );
and \U$920 ( \1297 , \1289 , \1296 );
and \U$921 ( \1298 , \1280 , \1288 );
or \U$922 ( \1299 , \1297 , \1298 );
and \U$923 ( \1300 , \1273 , \1299 );
and \U$924 ( \1301 , \1251 , \1272 );
nor \U$925 ( \1302 , \1300 , \1301 );
xor \U$926 ( \1303 , \1230 , \1302 );
xor \U$927 ( \1304 , \1008 , \1012 );
xor \U$928 ( \1305 , \1304 , \1021 );
xor \U$929 ( \1306 , \1102 , \1107 );
xor \U$930 ( \1307 , \1305 , \1306 );
and \U$931 ( \1308 , \1303 , \1307 );
and \U$932 ( \1309 , \1230 , \1302 );
or \U$933 ( \1310 , \1308 , \1309 );
xor \U$934 ( \1311 , \1024 , \1035 );
xor \U$935 ( \1312 , \1311 , \1063 );
xor \U$936 ( \1313 , \1310 , \1312 );
xor \U$937 ( \1314 , \1112 , \1187 );
xor \U$938 ( \1315 , \1314 , \1190 );
and \U$939 ( \1316 , \1313 , \1315 );
and \U$940 ( \1317 , \1310 , \1312 );
or \U$941 ( \1318 , \1316 , \1317 );
nand \U$942 ( \1319 , \1210 , \1318 );
or \U$943 ( \1320 , \1199 , \1319 );
xnor \U$944 ( \1321 , \1319 , \1199 );
not \U$945 ( \1322 , \1318 );
not \U$946 ( \1323 , \1209 );
or \U$947 ( \1324 , \1322 , \1323 );
or \U$948 ( \1325 , \1209 , \1318 );
nand \U$949 ( \1326 , \1324 , \1325 );
xor \U$950 ( \1327 , \1310 , \1312 );
xor \U$951 ( \1328 , \1327 , \1315 );
not \U$952 ( \1329 , \1328 );
xor \U$953 ( \1330 , \1230 , \1302 );
xor \U$954 ( \1331 , \1330 , \1307 );
xor \U$955 ( \1332 , \1146 , \1156 );
xor \U$956 ( \1333 , \1332 , \1184 );
and \U$957 ( \1334 , \1331 , \1333 );
not \U$958 ( \1335 , \1331 );
not \U$959 ( \1336 , \1333 );
and \U$960 ( \1337 , \1335 , \1336 );
xor \U$961 ( \1338 , \1259 , \1261 );
xor \U$962 ( \1339 , \1338 , \1269 );
xor \U$963 ( \1340 , \1238 , \1239 );
xor \U$964 ( \1341 , \1340 , \1248 );
and \U$965 ( \1342 , \1339 , \1341 );
xor \U$966 ( \1343 , \1280 , \1288 );
xor \U$967 ( \1344 , \1343 , \1296 );
xor \U$968 ( \1345 , \1238 , \1239 );
xor \U$969 ( \1346 , \1345 , \1248 );
and \U$970 ( \1347 , \1344 , \1346 );
and \U$971 ( \1348 , \1339 , \1344 );
or \U$972 ( \1349 , \1342 , \1347 , \1348 );
and \U$973 ( \1350 , \883 , RIae76898_51);
and \U$974 ( \1351 , RIae76b68_57, \881 );
nor \U$975 ( \1352 , \1350 , \1351 );
not \U$976 ( \1353 , \1352 );
not \U$977 ( \1354 , \789 );
and \U$978 ( \1355 , \1353 , \1354 );
and \U$979 ( \1356 , \1352 , \789 );
nor \U$980 ( \1357 , \1355 , \1356 );
not \U$981 ( \1358 , \1357 );
and \U$982 ( \1359 , \1138 , RIae78a58_123);
and \U$983 ( \1360 , RIae78cb0_128, \1136 );
nor \U$984 ( \1361 , \1359 , \1360 );
and \U$985 ( \1362 , \1361 , \1142 );
not \U$986 ( \1363 , \1361 );
and \U$987 ( \1364 , \1363 , \1012 );
nor \U$988 ( \1365 , \1362 , \1364 );
not \U$989 ( \1366 , \1365 );
and \U$990 ( \1367 , \1358 , \1366 );
and \U$991 ( \1368 , \1365 , \1357 );
and \U$992 ( \1369 , RIae793b8_143, RIae799d0_156);
not \U$993 ( \1370 , RIae799d0_156);
nor \U$994 ( \1371 , \1370 , RIae79610_148);
not \U$995 ( \1372 , RIae79610_148);
nor \U$996 ( \1373 , \1372 , RIae799d0_156);
or \U$997 ( \1374 , \1371 , \1373 );
nor \U$998 ( \1375 , RIae793b8_143, RIae799d0_156);
nor \U$999 ( \1376 , \1369 , \1374 , \1375 );
nand \U$1000 ( \1377 , RIae78da0_130, \1376 );
and \U$1001 ( \1378 , \1377 , \1261 );
not \U$1002 ( \1379 , \1377 );
not \U$1003 ( \1380 , \1261 );
and \U$1004 ( \1381 , \1379 , \1380 );
nor \U$1005 ( \1382 , \1378 , \1381 );
nor \U$1006 ( \1383 , \1368 , \1382 );
nor \U$1007 ( \1384 , \1367 , \1383 );
and \U$1008 ( \1385 , \436 , RIae765c8_45);
and \U$1009 ( \1386 , RIae76118_35, \434 );
nor \U$1010 ( \1387 , \1385 , \1386 );
not \U$1011 ( \1388 , \1387 );
not \U$1012 ( \1389 , \400 );
and \U$1013 ( \1390 , \1388 , \1389 );
and \U$1014 ( \1391 , \1387 , \400 );
nor \U$1015 ( \1392 , \1390 , \1391 );
nand \U$1016 ( \1393 , RIae763e8_41, RIae78b48_125);
xor \U$1017 ( \1394 , \1392 , \1393 );
and \U$1018 ( \1395 , \384 , RIae764d8_43);
and \U$1019 ( \1396 , RIae766b8_47, \382 );
nor \U$1020 ( \1397 , \1395 , \1396 );
not \U$1021 ( \1398 , \1397 );
not \U$1022 ( \1399 , \392 );
and \U$1023 ( \1400 , \1398 , \1399 );
and \U$1024 ( \1401 , \1397 , \388 );
nor \U$1025 ( \1402 , \1400 , \1401 );
and \U$1026 ( \1403 , \1394 , \1402 );
and \U$1027 ( \1404 , \1392 , \1393 );
or \U$1028 ( \1405 , \1403 , \1404 );
xor \U$1029 ( \1406 , \1384 , \1405 );
and \U$1030 ( \1407 , \514 , RIae76028_33);
and \U$1031 ( \1408 , RIae762f8_39, \512 );
nor \U$1032 ( \1409 , \1407 , \1408 );
not \U$1033 ( \1410 , \1409 );
not \U$1034 ( \1411 , \471 );
and \U$1035 ( \1412 , \1410 , \1411 );
and \U$1036 ( \1413 , \1409 , \469 );
nor \U$1037 ( \1414 , \1412 , \1413 );
and \U$1038 ( \1415 , \558 , RIae76208_37);
and \U$1039 ( \1416 , RIae76a78_55, \556 );
nor \U$1040 ( \1417 , \1415 , \1416 );
and \U$1041 ( \1418 , \1417 , \562 );
not \U$1042 ( \1419 , \1417 );
and \U$1043 ( \1420 , \1419 , \504 );
nor \U$1044 ( \1421 , \1418 , \1420 );
xor \U$1045 ( \1422 , \1414 , \1421 );
and \U$1046 ( \1423 , \672 , RIae76988_53);
and \U$1047 ( \1424 , RIae767a8_49, \670 );
nor \U$1048 ( \1425 , \1423 , \1424 );
and \U$1049 ( \1426 , \1425 , \587 );
not \U$1050 ( \1427 , \1425 );
and \U$1051 ( \1428 , \1427 , \588 );
nor \U$1052 ( \1429 , \1426 , \1428 );
and \U$1053 ( \1430 , \1422 , \1429 );
and \U$1054 ( \1431 , \1414 , \1421 );
or \U$1055 ( \1432 , \1430 , \1431 );
and \U$1056 ( \1433 , \1406 , \1432 );
and \U$1057 ( \1434 , \1384 , \1405 );
or \U$1058 ( \1435 , \1433 , \1434 );
xor \U$1059 ( \1436 , \1349 , \1435 );
xnor \U$1060 ( \1437 , \1220 , \1222 );
not \U$1061 ( \1438 , \1437 );
not \U$1062 ( \1439 , \1228 );
and \U$1063 ( \1440 , \1438 , \1439 );
and \U$1064 ( \1441 , \1437 , \1228 );
nor \U$1065 ( \1442 , \1440 , \1441 );
and \U$1066 ( \1443 , \1436 , \1442 );
and \U$1067 ( \1444 , \1349 , \1435 );
or \U$1068 ( \1445 , \1443 , \1444 );
nor \U$1069 ( \1446 , \1337 , \1445 );
nor \U$1070 ( \1447 , \1334 , \1446 );
nor \U$1071 ( \1448 , \1329 , \1447 );
and \U$1072 ( \1449 , \1326 , \1448 );
xor \U$1073 ( \1450 , \1448 , \1326 );
not \U$1074 ( \1451 , \400 );
and \U$1075 ( \1452 , \436 , RIae766b8_47);
and \U$1076 ( \1453 , RIae765c8_45, \434 );
nor \U$1077 ( \1454 , \1452 , \1453 );
not \U$1078 ( \1455 , \1454 );
or \U$1079 ( \1456 , \1451 , \1455 );
or \U$1080 ( \1457 , \1454 , \400 );
nand \U$1081 ( \1458 , \1456 , \1457 );
not \U$1082 ( \1459 , \469 );
and \U$1083 ( \1460 , \514 , RIae76118_35);
and \U$1084 ( \1461 , RIae76028_33, \512 );
nor \U$1085 ( \1462 , \1460 , \1461 );
not \U$1086 ( \1463 , \1462 );
or \U$1087 ( \1464 , \1459 , \1463 );
or \U$1088 ( \1465 , \1462 , \469 );
nand \U$1089 ( \1466 , \1464 , \1465 );
xor \U$1090 ( \1467 , \1458 , \1466 );
not \U$1091 ( \1468 , \392 );
and \U$1092 ( \1469 , \384 , RIae763e8_41);
and \U$1093 ( \1470 , RIae764d8_43, \382 );
nor \U$1094 ( \1471 , \1469 , \1470 );
not \U$1095 ( \1472 , \1471 );
or \U$1096 ( \1473 , \1468 , \1472 );
or \U$1097 ( \1474 , \1471 , \388 );
nand \U$1098 ( \1475 , \1473 , \1474 );
and \U$1099 ( \1476 , \1467 , \1475 );
and \U$1100 ( \1477 , \1458 , \1466 );
nor \U$1101 ( \1478 , \1476 , \1477 );
and \U$1102 ( \1479 , \1376 , RIae78cb0_128);
and \U$1103 ( \1480 , RIae78da0_130, \1374 );
nor \U$1104 ( \1481 , \1479 , \1480 );
and \U$1105 ( \1482 , \1481 , \1380 );
not \U$1106 ( \1483 , \1481 );
and \U$1107 ( \1484 , \1483 , \1261 );
nor \U$1108 ( \1485 , \1482 , \1484 );
not \U$1109 ( \1486 , \1485 );
nand \U$1110 ( \1487 , RIae79688_149, RIae79598_147);
and \U$1111 ( \1488 , \1487 , RIae79610_148);
nand \U$1112 ( \1489 , \1486 , \1488 );
and \U$1113 ( \1490 , \1138 , RIae76b68_57);
and \U$1114 ( \1491 , RIae78a58_123, \1136 );
nor \U$1115 ( \1492 , \1490 , \1491 );
and \U$1116 ( \1493 , \1492 , \1012 );
not \U$1117 ( \1494 , \1492 );
and \U$1118 ( \1495 , \1494 , \1142 );
nor \U$1119 ( \1496 , \1493 , \1495 );
and \U$1120 ( \1497 , \1489 , \1496 );
not \U$1121 ( \1498 , \1488 );
and \U$1122 ( \1499 , \1498 , \1485 );
nor \U$1123 ( \1500 , \1497 , \1499 );
xor \U$1124 ( \1501 , \1478 , \1500 );
and \U$1125 ( \1502 , \672 , RIae76a78_55);
and \U$1126 ( \1503 , RIae76988_53, \670 );
nor \U$1127 ( \1504 , \1502 , \1503 );
and \U$1128 ( \1505 , \1504 , \588 );
not \U$1129 ( \1506 , \1504 );
and \U$1130 ( \1507 , \1506 , \587 );
nor \U$1131 ( \1508 , \1505 , \1507 );
not \U$1132 ( \1509 , \787 );
and \U$1133 ( \1510 , \883 , RIae767a8_49);
and \U$1134 ( \1511 , RIae76898_51, \881 );
nor \U$1135 ( \1512 , \1510 , \1511 );
not \U$1136 ( \1513 , \1512 );
or \U$1137 ( \1514 , \1509 , \1513 );
or \U$1138 ( \1515 , \1512 , \789 );
nand \U$1139 ( \1516 , \1514 , \1515 );
xor \U$1140 ( \1517 , \1508 , \1516 );
and \U$1141 ( \1518 , \558 , RIae762f8_39);
and \U$1142 ( \1519 , RIae76208_37, \556 );
nor \U$1143 ( \1520 , \1518 , \1519 );
and \U$1144 ( \1521 , \1520 , \504 );
not \U$1145 ( \1522 , \1520 );
and \U$1146 ( \1523 , \1522 , \562 );
nor \U$1147 ( \1524 , \1521 , \1523 );
and \U$1148 ( \1525 , \1517 , \1524 );
and \U$1149 ( \1526 , \1508 , \1516 );
nor \U$1150 ( \1527 , \1525 , \1526 );
and \U$1151 ( \1528 , \1501 , \1527 );
and \U$1152 ( \1529 , \1478 , \1500 );
or \U$1153 ( \1530 , \1528 , \1529 );
xor \U$1154 ( \1531 , \1392 , \1393 );
xor \U$1155 ( \1532 , \1531 , \1402 );
xor \U$1156 ( \1533 , \1414 , \1421 );
xor \U$1157 ( \1534 , \1533 , \1429 );
nand \U$1158 ( \1535 , \1532 , \1534 );
not \U$1159 ( \1536 , \1535 );
xor \U$1160 ( \1537 , \1530 , \1536 );
xor \U$1161 ( \1538 , \1238 , \1239 );
xor \U$1162 ( \1539 , \1538 , \1248 );
xor \U$1163 ( \1540 , \1339 , \1344 );
xor \U$1164 ( \1541 , \1539 , \1540 );
and \U$1165 ( \1542 , \1537 , \1541 );
and \U$1166 ( \1543 , \1530 , \1536 );
or \U$1167 ( \1544 , \1542 , \1543 );
xor \U$1168 ( \1545 , \1251 , \1272 );
xor \U$1169 ( \1546 , \1545 , \1299 );
xor \U$1170 ( \1547 , \1544 , \1546 );
xor \U$1171 ( \1548 , \1349 , \1435 );
xor \U$1172 ( \1549 , \1548 , \1442 );
xor \U$1173 ( \1550 , \1547 , \1549 );
and \U$1174 ( \1551 , \436 , RIae764d8_43);
and \U$1175 ( \1552 , RIae766b8_47, \434 );
nor \U$1176 ( \1553 , \1551 , \1552 );
not \U$1177 ( \1554 , \1553 );
not \U$1178 ( \1555 , \400 );
and \U$1179 ( \1556 , \1554 , \1555 );
and \U$1180 ( \1557 , \1553 , \400 );
nor \U$1181 ( \1558 , \1556 , \1557 );
and \U$1182 ( \1559 , \514 , RIae765c8_45);
and \U$1183 ( \1560 , RIae76118_35, \512 );
nor \U$1184 ( \1561 , \1559 , \1560 );
not \U$1185 ( \1562 , \1561 );
not \U$1186 ( \1563 , \469 );
and \U$1187 ( \1564 , \1562 , \1563 );
and \U$1188 ( \1565 , \1561 , \471 );
nor \U$1189 ( \1566 , \1564 , \1565 );
xor \U$1190 ( \1567 , \1558 , \1566 );
and \U$1191 ( \1568 , \384 , RIae753f8_7);
and \U$1192 ( \1569 , RIae763e8_41, \382 );
nor \U$1193 ( \1570 , \1568 , \1569 );
not \U$1194 ( \1571 , \1570 );
not \U$1195 ( \1572 , \388 );
and \U$1196 ( \1573 , \1571 , \1572 );
and \U$1197 ( \1574 , \1570 , \392 );
nor \U$1198 ( \1575 , \1573 , \1574 );
and \U$1199 ( \1576 , \1567 , \1575 );
and \U$1200 ( \1577 , \1558 , \1566 );
nor \U$1201 ( \1578 , \1576 , \1577 );
and \U$1202 ( \1579 , \1138 , RIae76898_51);
and \U$1203 ( \1580 , RIae76b68_57, \1136 );
nor \U$1204 ( \1581 , \1579 , \1580 );
and \U$1205 ( \1582 , \1581 , \1012 );
not \U$1206 ( \1583 , \1581 );
and \U$1207 ( \1584 , \1583 , \1142 );
nor \U$1208 ( \1585 , \1582 , \1584 );
and \U$1209 ( \1586 , RIae79610_148, RIae79598_147);
not \U$1210 ( \1587 , RIae79598_147);
nor \U$1211 ( \1588 , \1587 , RIae79688_149);
not \U$1212 ( \1589 , RIae79688_149);
nor \U$1213 ( \1590 , \1589 , RIae79598_147);
or \U$1214 ( \1591 , \1588 , \1590 );
nor \U$1215 ( \1592 , RIae79610_148, RIae79598_147);
nor \U$1216 ( \1593 , \1586 , \1591 , \1592 );
nand \U$1217 ( \1594 , RIae78da0_130, \1593 );
and \U$1218 ( \1595 , \1594 , \1498 );
not \U$1219 ( \1596 , \1594 );
and \U$1220 ( \1597 , \1596 , \1488 );
nor \U$1221 ( \1598 , \1595 , \1597 );
xor \U$1222 ( \1599 , \1585 , \1598 );
and \U$1223 ( \1600 , \1376 , RIae78a58_123);
and \U$1224 ( \1601 , RIae78cb0_128, \1374 );
nor \U$1225 ( \1602 , \1600 , \1601 );
and \U$1226 ( \1603 , \1602 , \1380 );
not \U$1227 ( \1604 , \1602 );
and \U$1228 ( \1605 , \1604 , \1261 );
nor \U$1229 ( \1606 , \1603 , \1605 );
and \U$1230 ( \1607 , \1599 , \1606 );
and \U$1231 ( \1608 , \1585 , \1598 );
or \U$1232 ( \1609 , \1607 , \1608 );
xor \U$1233 ( \1610 , \1578 , \1609 );
and \U$1234 ( \1611 , \558 , RIae76028_33);
and \U$1235 ( \1612 , RIae762f8_39, \556 );
nor \U$1236 ( \1613 , \1611 , \1612 );
and \U$1237 ( \1614 , \1613 , \504 );
not \U$1238 ( \1615 , \1613 );
and \U$1239 ( \1616 , \1615 , \562 );
nor \U$1240 ( \1617 , \1614 , \1616 );
and \U$1241 ( \1618 , \672 , RIae76208_37);
and \U$1242 ( \1619 , RIae76a78_55, \670 );
nor \U$1243 ( \1620 , \1618 , \1619 );
and \U$1244 ( \1621 , \1620 , \588 );
not \U$1245 ( \1622 , \1620 );
and \U$1246 ( \1623 , \1622 , \587 );
nor \U$1247 ( \1624 , \1621 , \1623 );
xor \U$1248 ( \1625 , \1617 , \1624 );
not \U$1249 ( \1626 , \789 );
and \U$1250 ( \1627 , \883 , RIae76988_53);
and \U$1251 ( \1628 , RIae767a8_49, \881 );
nor \U$1252 ( \1629 , \1627 , \1628 );
not \U$1253 ( \1630 , \1629 );
or \U$1254 ( \1631 , \1626 , \1630 );
or \U$1255 ( \1632 , \1629 , \787 );
nand \U$1256 ( \1633 , \1631 , \1632 );
and \U$1257 ( \1634 , \1625 , \1633 );
and \U$1258 ( \1635 , \1617 , \1624 );
or \U$1259 ( \1636 , \1634 , \1635 );
and \U$1260 ( \1637 , \1610 , \1636 );
and \U$1261 ( \1638 , \1578 , \1609 );
or \U$1262 ( \1639 , \1637 , \1638 );
not \U$1263 ( \1640 , \1357 );
xor \U$1264 ( \1641 , \1382 , \1365 );
not \U$1265 ( \1642 , \1641 );
or \U$1266 ( \1643 , \1640 , \1642 );
or \U$1267 ( \1644 , \1641 , \1357 );
nand \U$1268 ( \1645 , \1643 , \1644 );
and \U$1269 ( \1646 , \1639 , \1645 );
not \U$1270 ( \1647 , \1639 );
not \U$1271 ( \1648 , \1645 );
and \U$1272 ( \1649 , \1647 , \1648 );
xor \U$1273 ( \1650 , \1508 , \1516 );
xor \U$1274 ( \1651 , \1650 , \1524 );
not \U$1275 ( \1652 , RIae753f8_7);
nor \U$1276 ( \1653 , \1652 , \491 );
xor \U$1277 ( \1654 , \1651 , \1653 );
xor \U$1278 ( \1655 , \1458 , \1466 );
xor \U$1279 ( \1656 , \1655 , \1475 );
and \U$1280 ( \1657 , \1654 , \1656 );
and \U$1281 ( \1658 , \1651 , \1653 );
nor \U$1282 ( \1659 , \1657 , \1658 );
nor \U$1283 ( \1660 , \1649 , \1659 );
nor \U$1284 ( \1661 , \1646 , \1660 );
xor \U$1285 ( \1662 , \1384 , \1405 );
xor \U$1286 ( \1663 , \1662 , \1432 );
xor \U$1287 ( \1664 , \1661 , \1663 );
xor \U$1288 ( \1665 , \1530 , \1536 );
xor \U$1289 ( \1666 , \1665 , \1541 );
and \U$1290 ( \1667 , \1664 , \1666 );
and \U$1291 ( \1668 , \1661 , \1663 );
or \U$1292 ( \1669 , \1667 , \1668 );
or \U$1293 ( \1670 , \1550 , \1669 );
not \U$1294 ( \1671 , \1669 );
not \U$1295 ( \1672 , \1550 );
or \U$1296 ( \1673 , \1671 , \1672 );
xor \U$1297 ( \1674 , \1661 , \1663 );
xor \U$1298 ( \1675 , \1674 , \1666 );
xor \U$1299 ( \1676 , \1478 , \1500 );
xor \U$1300 ( \1677 , \1676 , \1527 );
not \U$1301 ( \1678 , \1677 );
not \U$1302 ( \1679 , \1639 );
not \U$1303 ( \1680 , \1659 );
or \U$1304 ( \1681 , \1679 , \1680 );
or \U$1305 ( \1682 , \1659 , \1639 );
nand \U$1306 ( \1683 , \1681 , \1682 );
xor \U$1307 ( \1684 , \1645 , \1683 );
nand \U$1308 ( \1685 , \1678 , \1684 );
or \U$1309 ( \1686 , \1675 , \1685 );
not \U$1310 ( \1687 , \1685 );
not \U$1311 ( \1688 , \1675 );
or \U$1312 ( \1689 , \1687 , \1688 );
xor \U$1313 ( \1690 , \1617 , \1624 );
xor \U$1314 ( \1691 , \1690 , \1633 );
xor \U$1315 ( \1692 , \1585 , \1598 );
xor \U$1316 ( \1693 , \1692 , \1606 );
and \U$1317 ( \1694 , \1691 , \1693 );
nand \U$1318 ( \1695 , RIae75308_5, RIae78b48_125);
xor \U$1319 ( \1696 , \1558 , \1566 );
xor \U$1320 ( \1697 , \1696 , \1575 );
nand \U$1321 ( \1698 , \1695 , \1697 );
xor \U$1322 ( \1699 , \1694 , \1698 );
and \U$1323 ( \1700 , \672 , RIae762f8_39);
and \U$1324 ( \1701 , RIae76208_37, \670 );
nor \U$1325 ( \1702 , \1700 , \1701 );
and \U$1326 ( \1703 , \1702 , \588 );
not \U$1327 ( \1704 , \1702 );
and \U$1328 ( \1705 , \1704 , \587 );
nor \U$1329 ( \1706 , \1703 , \1705 );
not \U$1330 ( \1707 , \787 );
and \U$1331 ( \1708 , \883 , RIae76a78_55);
and \U$1332 ( \1709 , RIae76988_53, \881 );
nor \U$1333 ( \1710 , \1708 , \1709 );
not \U$1334 ( \1711 , \1710 );
or \U$1335 ( \1712 , \1707 , \1711 );
or \U$1336 ( \1713 , \1710 , \787 );
nand \U$1337 ( \1714 , \1712 , \1713 );
xor \U$1338 ( \1715 , \1706 , \1714 );
and \U$1339 ( \1716 , \1138 , RIae767a8_49);
and \U$1340 ( \1717 , RIae76898_51, \1136 );
nor \U$1341 ( \1718 , \1716 , \1717 );
and \U$1342 ( \1719 , \1718 , \1012 );
not \U$1343 ( \1720 , \1718 );
and \U$1344 ( \1721 , \1720 , \1142 );
nor \U$1345 ( \1722 , \1719 , \1721 );
and \U$1346 ( \1723 , \1715 , \1722 );
and \U$1347 ( \1724 , \1706 , \1714 );
or \U$1348 ( \1725 , \1723 , \1724 );
and \U$1349 ( \1726 , \1593 , RIae78cb0_128);
and \U$1350 ( \1727 , RIae78da0_130, \1591 );
nor \U$1351 ( \1728 , \1726 , \1727 );
and \U$1352 ( \1729 , \1728 , \1498 );
not \U$1353 ( \1730 , \1728 );
and \U$1354 ( \1731 , \1730 , \1488 );
nor \U$1355 ( \1732 , \1729 , \1731 );
nand \U$1356 ( \1733 , RIae79ac0_158, RIae79b38_159);
and \U$1357 ( \1734 , \1733 , RIae79688_149);
not \U$1358 ( \1735 , \1734 );
xor \U$1359 ( \1736 , \1732 , \1735 );
and \U$1360 ( \1737 , \1376 , RIae76b68_57);
and \U$1361 ( \1738 , RIae78a58_123, \1374 );
nor \U$1362 ( \1739 , \1737 , \1738 );
and \U$1363 ( \1740 , \1739 , \1380 );
not \U$1364 ( \1741 , \1739 );
and \U$1365 ( \1742 , \1741 , \1261 );
nor \U$1366 ( \1743 , \1740 , \1742 );
and \U$1367 ( \1744 , \1736 , \1743 );
and \U$1368 ( \1745 , \1732 , \1735 );
or \U$1369 ( \1746 , \1744 , \1745 );
xor \U$1370 ( \1747 , \1725 , \1746 );
not \U$1371 ( \1748 , \402 );
and \U$1372 ( \1749 , \436 , RIae763e8_41);
and \U$1373 ( \1750 , RIae764d8_43, \434 );
nor \U$1374 ( \1751 , \1749 , \1750 );
not \U$1375 ( \1752 , \1751 );
or \U$1376 ( \1753 , \1748 , \1752 );
or \U$1377 ( \1754 , \1751 , \400 );
nand \U$1378 ( \1755 , \1753 , \1754 );
not \U$1379 ( \1756 , \471 );
and \U$1380 ( \1757 , \514 , RIae766b8_47);
and \U$1381 ( \1758 , RIae765c8_45, \512 );
nor \U$1382 ( \1759 , \1757 , \1758 );
not \U$1383 ( \1760 , \1759 );
or \U$1384 ( \1761 , \1756 , \1760 );
or \U$1385 ( \1762 , \1759 , \469 );
nand \U$1386 ( \1763 , \1761 , \1762 );
xor \U$1387 ( \1764 , \1755 , \1763 );
and \U$1388 ( \1765 , \558 , RIae76118_35);
and \U$1389 ( \1766 , RIae76028_33, \556 );
nor \U$1390 ( \1767 , \1765 , \1766 );
and \U$1391 ( \1768 , \1767 , \504 );
not \U$1392 ( \1769 , \1767 );
and \U$1393 ( \1770 , \1769 , \562 );
nor \U$1394 ( \1771 , \1768 , \1770 );
and \U$1395 ( \1772 , \1764 , \1771 );
and \U$1396 ( \1773 , \1755 , \1763 );
or \U$1397 ( \1774 , \1772 , \1773 );
and \U$1398 ( \1775 , \1747 , \1774 );
and \U$1399 ( \1776 , \1725 , \1746 );
or \U$1400 ( \1777 , \1775 , \1776 );
and \U$1401 ( \1778 , \1699 , \1777 );
and \U$1402 ( \1779 , \1694 , \1698 );
or \U$1403 ( \1780 , \1778 , \1779 );
or \U$1404 ( \1781 , \1532 , \1534 );
nand \U$1405 ( \1782 , \1781 , \1535 );
xor \U$1406 ( \1783 , \1780 , \1782 );
not \U$1407 ( \1784 , \1496 );
and \U$1408 ( \1785 , \1485 , \1488 );
not \U$1409 ( \1786 , \1485 );
and \U$1410 ( \1787 , \1786 , \1498 );
nor \U$1411 ( \1788 , \1785 , \1787 );
not \U$1412 ( \1789 , \1788 );
or \U$1413 ( \1790 , \1784 , \1789 );
or \U$1414 ( \1791 , \1788 , \1496 );
nand \U$1415 ( \1792 , \1790 , \1791 );
xor \U$1416 ( \1793 , \1578 , \1609 );
xor \U$1417 ( \1794 , \1793 , \1636 );
and \U$1418 ( \1795 , \1792 , \1794 );
xor \U$1419 ( \1796 , \1651 , \1653 );
xor \U$1420 ( \1797 , \1796 , \1656 );
xor \U$1421 ( \1798 , \1578 , \1609 );
xor \U$1422 ( \1799 , \1798 , \1636 );
and \U$1423 ( \1800 , \1797 , \1799 );
and \U$1424 ( \1801 , \1792 , \1797 );
or \U$1425 ( \1802 , \1795 , \1800 , \1801 );
and \U$1426 ( \1803 , \1783 , \1802 );
and \U$1427 ( \1804 , \1780 , \1782 );
or \U$1428 ( \1805 , \1803 , \1804 );
nand \U$1429 ( \1806 , \1689 , \1805 );
nand \U$1430 ( \1807 , \1686 , \1806 );
nand \U$1431 ( \1808 , \1673 , \1807 );
nand \U$1432 ( \1809 , \1670 , \1808 );
not \U$1433 ( \1810 , \1331 );
not \U$1434 ( \1811 , \1445 );
not \U$1435 ( \1812 , \1333 );
and \U$1436 ( \1813 , \1811 , \1812 );
and \U$1437 ( \1814 , \1445 , \1333 );
nor \U$1438 ( \1815 , \1813 , \1814 );
not \U$1439 ( \1816 , \1815 );
or \U$1440 ( \1817 , \1810 , \1816 );
or \U$1441 ( \1818 , \1815 , \1331 );
nand \U$1442 ( \1819 , \1817 , \1818 );
not \U$1443 ( \1820 , \1819 );
xor \U$1444 ( \1821 , \1544 , \1546 );
and \U$1445 ( \1822 , \1821 , \1549 );
and \U$1446 ( \1823 , \1544 , \1546 );
or \U$1447 ( \1824 , \1822 , \1823 );
not \U$1448 ( \1825 , \1824 );
or \U$1449 ( \1826 , \1820 , \1825 );
or \U$1450 ( \1827 , \1824 , \1819 );
nand \U$1451 ( \1828 , \1826 , \1827 );
and \U$1452 ( \1829 , \1809 , \1828 );
xor \U$1453 ( \1830 , \1828 , \1809 );
not \U$1454 ( \1831 , \1669 );
not \U$1455 ( \1832 , \1807 );
or \U$1456 ( \1833 , \1831 , \1832 );
or \U$1457 ( \1834 , \1807 , \1669 );
nand \U$1458 ( \1835 , \1833 , \1834 );
not \U$1459 ( \1836 , \1835 );
not \U$1460 ( \1837 , \1550 );
and \U$1461 ( \1838 , \1836 , \1837 );
and \U$1462 ( \1839 , \1835 , \1550 );
nor \U$1463 ( \1840 , \1838 , \1839 );
not \U$1464 ( \1841 , \1685 );
not \U$1465 ( \1842 , \1805 );
or \U$1466 ( \1843 , \1841 , \1842 );
or \U$1467 ( \1844 , \1805 , \1685 );
nand \U$1468 ( \1845 , \1843 , \1844 );
not \U$1469 ( \1846 , \1845 );
not \U$1470 ( \1847 , \1675 );
and \U$1471 ( \1848 , \1846 , \1847 );
and \U$1472 ( \1849 , \1845 , \1675 );
nor \U$1473 ( \1850 , \1848 , \1849 );
not \U$1474 ( \1851 , \1850 );
not \U$1475 ( \1852 , \1677 );
not \U$1476 ( \1853 , \1684 );
or \U$1477 ( \1854 , \1852 , \1853 );
or \U$1478 ( \1855 , \1684 , \1677 );
nand \U$1479 ( \1856 , \1854 , \1855 );
not \U$1480 ( \1857 , \1856 );
xor \U$1481 ( \1858 , \1780 , \1782 );
xor \U$1482 ( \1859 , \1858 , \1802 );
not \U$1483 ( \1860 , \1859 );
or \U$1484 ( \1861 , \1857 , \1860 );
or \U$1485 ( \1862 , \1859 , \1856 );
or \U$1486 ( \1863 , \1697 , \1695 );
nand \U$1487 ( \1864 , \1863 , \1698 );
xor \U$1488 ( \1865 , \1691 , \1693 );
xor \U$1489 ( \1866 , \1864 , \1865 );
xor \U$1490 ( \1867 , \1725 , \1746 );
xor \U$1491 ( \1868 , \1867 , \1774 );
and \U$1492 ( \1869 , \1866 , \1868 );
and \U$1493 ( \1870 , \1864 , \1865 );
or \U$1494 ( \1871 , \1869 , \1870 );
and \U$1495 ( \1872 , \672 , RIae76028_33);
and \U$1496 ( \1873 , RIae762f8_39, \670 );
nor \U$1497 ( \1874 , \1872 , \1873 );
and \U$1498 ( \1875 , \1874 , \588 );
not \U$1499 ( \1876 , \1874 );
and \U$1500 ( \1877 , \1876 , \587 );
nor \U$1501 ( \1878 , \1875 , \1877 );
not \U$1502 ( \1879 , \789 );
and \U$1503 ( \1880 , \883 , RIae76208_37);
and \U$1504 ( \1881 , RIae76a78_55, \881 );
nor \U$1505 ( \1882 , \1880 , \1881 );
not \U$1506 ( \1883 , \1882 );
or \U$1507 ( \1884 , \1879 , \1883 );
or \U$1508 ( \1885 , \1882 , \789 );
nand \U$1509 ( \1886 , \1884 , \1885 );
xor \U$1510 ( \1887 , \1878 , \1886 );
and \U$1511 ( \1888 , \1138 , RIae76988_53);
and \U$1512 ( \1889 , RIae767a8_49, \1136 );
nor \U$1513 ( \1890 , \1888 , \1889 );
and \U$1514 ( \1891 , \1890 , \1012 );
not \U$1515 ( \1892 , \1890 );
and \U$1516 ( \1893 , \1892 , \1142 );
nor \U$1517 ( \1894 , \1891 , \1893 );
and \U$1518 ( \1895 , \1887 , \1894 );
and \U$1519 ( \1896 , \1878 , \1886 );
or \U$1520 ( \1897 , \1895 , \1896 );
not \U$1521 ( \1898 , \471 );
and \U$1522 ( \1899 , \514 , RIae764d8_43);
and \U$1523 ( \1900 , RIae766b8_47, \512 );
nor \U$1524 ( \1901 , \1899 , \1900 );
not \U$1525 ( \1902 , \1901 );
or \U$1526 ( \1903 , \1898 , \1902 );
or \U$1527 ( \1904 , \1901 , \469 );
nand \U$1528 ( \1905 , \1903 , \1904 );
not \U$1529 ( \1906 , \402 );
and \U$1530 ( \1907 , \436 , RIae753f8_7);
and \U$1531 ( \1908 , RIae763e8_41, \434 );
nor \U$1532 ( \1909 , \1907 , \1908 );
not \U$1533 ( \1910 , \1909 );
or \U$1534 ( \1911 , \1906 , \1910 );
or \U$1535 ( \1912 , \1909 , \402 );
nand \U$1536 ( \1913 , \1911 , \1912 );
xor \U$1537 ( \1914 , \1905 , \1913 );
and \U$1538 ( \1915 , \558 , RIae765c8_45);
and \U$1539 ( \1916 , RIae76118_35, \556 );
nor \U$1540 ( \1917 , \1915 , \1916 );
and \U$1541 ( \1918 , \1917 , \504 );
not \U$1542 ( \1919 , \1917 );
and \U$1543 ( \1920 , \1919 , \562 );
nor \U$1544 ( \1921 , \1918 , \1920 );
and \U$1545 ( \1922 , \1914 , \1921 );
and \U$1546 ( \1923 , \1905 , \1913 );
or \U$1547 ( \1924 , \1922 , \1923 );
xor \U$1548 ( \1925 , \1897 , \1924 );
and \U$1549 ( \1926 , \1376 , RIae76898_51);
and \U$1550 ( \1927 , RIae76b68_57, \1374 );
nor \U$1551 ( \1928 , \1926 , \1927 );
and \U$1552 ( \1929 , \1928 , \1380 );
not \U$1553 ( \1930 , \1928 );
and \U$1554 ( \1931 , \1930 , \1261 );
nor \U$1555 ( \1932 , \1929 , \1931 );
and \U$1556 ( \1933 , RIae79688_149, RIae79b38_159);
not \U$1557 ( \1934 , RIae79ac0_158);
and \U$1558 ( \1935 , \1934 , RIae79b38_159);
nor \U$1559 ( \1936 , \1934 , RIae79b38_159);
or \U$1560 ( \1937 , \1935 , \1936 );
nor \U$1561 ( \1938 , RIae79688_149, RIae79b38_159);
nor \U$1562 ( \1939 , \1933 , \1937 , \1938 );
nand \U$1563 ( \1940 , RIae78da0_130, \1939 );
and \U$1564 ( \1941 , \1940 , \1735 );
not \U$1565 ( \1942 , \1940 );
and \U$1566 ( \1943 , \1942 , \1734 );
nor \U$1567 ( \1944 , \1941 , \1943 );
xor \U$1568 ( \1945 , \1932 , \1944 );
and \U$1569 ( \1946 , \1593 , RIae78a58_123);
and \U$1570 ( \1947 , RIae78cb0_128, \1591 );
nor \U$1571 ( \1948 , \1946 , \1947 );
and \U$1572 ( \1949 , \1948 , \1498 );
not \U$1573 ( \1950 , \1948 );
and \U$1574 ( \1951 , \1950 , \1488 );
nor \U$1575 ( \1952 , \1949 , \1951 );
and \U$1576 ( \1953 , \1945 , \1952 );
and \U$1577 ( \1954 , \1932 , \1944 );
or \U$1578 ( \1955 , \1953 , \1954 );
and \U$1579 ( \1956 , \1925 , \1955 );
and \U$1580 ( \1957 , \1897 , \1924 );
or \U$1581 ( \1958 , \1956 , \1957 );
not \U$1582 ( \1959 , \388 );
and \U$1583 ( \1960 , \384 , RIae75308_5);
and \U$1584 ( \1961 , RIae753f8_7, \382 );
nor \U$1585 ( \1962 , \1960 , \1961 );
not \U$1586 ( \1963 , \1962 );
or \U$1587 ( \1964 , \1959 , \1963 );
or \U$1588 ( \1965 , \1962 , \392 );
nand \U$1589 ( \1966 , \1964 , \1965 );
not \U$1590 ( \1967 , RIae75128_1);
nor \U$1591 ( \1968 , \1967 , \491 );
xor \U$1592 ( \1969 , \1966 , \1968 );
nand \U$1593 ( \1970 , RIae75218_3, RIae78b48_125);
and \U$1594 ( \1971 , \384 , RIae75128_1);
and \U$1595 ( \1972 , RIae75308_5, \382 );
nor \U$1596 ( \1973 , \1971 , \1972 );
not \U$1597 ( \1974 , \1973 );
not \U$1598 ( \1975 , \392 );
and \U$1599 ( \1976 , \1974 , \1975 );
and \U$1600 ( \1977 , \1973 , \392 );
nor \U$1601 ( \1978 , \1976 , \1977 );
nand \U$1602 ( \1979 , \1970 , \1978 );
and \U$1603 ( \1980 , \1969 , \1979 );
and \U$1604 ( \1981 , \1966 , \1968 );
or \U$1605 ( \1982 , \1980 , \1981 );
xor \U$1606 ( \1983 , \1958 , \1982 );
xor \U$1607 ( \1984 , \1732 , \1735 );
xor \U$1608 ( \1985 , \1984 , \1743 );
xor \U$1609 ( \1986 , \1755 , \1763 );
xor \U$1610 ( \1987 , \1986 , \1771 );
and \U$1611 ( \1988 , \1985 , \1987 );
xor \U$1612 ( \1989 , \1706 , \1714 );
xor \U$1613 ( \1990 , \1989 , \1722 );
xor \U$1614 ( \1991 , \1755 , \1763 );
xor \U$1615 ( \1992 , \1991 , \1771 );
and \U$1616 ( \1993 , \1990 , \1992 );
and \U$1617 ( \1994 , \1985 , \1990 );
or \U$1618 ( \1995 , \1988 , \1993 , \1994 );
and \U$1619 ( \1996 , \1983 , \1995 );
and \U$1620 ( \1997 , \1958 , \1982 );
or \U$1621 ( \1998 , \1996 , \1997 );
xor \U$1622 ( \1999 , \1871 , \1998 );
xor \U$1623 ( \2000 , \1578 , \1609 );
xor \U$1624 ( \2001 , \2000 , \1636 );
xor \U$1625 ( \2002 , \1792 , \1797 );
xor \U$1626 ( \2003 , \2001 , \2002 );
and \U$1627 ( \2004 , \1999 , \2003 );
and \U$1628 ( \2005 , \1871 , \1998 );
or \U$1629 ( \2006 , \2004 , \2005 );
nand \U$1630 ( \2007 , \1862 , \2006 );
nand \U$1631 ( \2008 , \1861 , \2007 );
nand \U$1632 ( \2009 , \1851 , \2008 );
or \U$1633 ( \2010 , \1840 , \2009 );
xnor \U$1634 ( \2011 , \2009 , \1840 );
xor \U$1635 ( \2012 , \1966 , \1968 );
xor \U$1636 ( \2013 , \2012 , \1979 );
xor \U$1637 ( \2014 , \1897 , \1924 );
xor \U$1638 ( \2015 , \2014 , \1955 );
and \U$1639 ( \2016 , \2013 , \2015 );
xor \U$1640 ( \2017 , \1755 , \1763 );
xor \U$1641 ( \2018 , \2017 , \1771 );
xor \U$1642 ( \2019 , \1985 , \1990 );
xor \U$1643 ( \2020 , \2018 , \2019 );
xor \U$1644 ( \2021 , \1897 , \1924 );
xor \U$1645 ( \2022 , \2021 , \1955 );
and \U$1646 ( \2023 , \2020 , \2022 );
and \U$1647 ( \2024 , \2013 , \2020 );
or \U$1648 ( \2025 , \2016 , \2023 , \2024 );
not \U$1649 ( \2026 , \789 );
and \U$1650 ( \2027 , \883 , RIae762f8_39);
and \U$1651 ( \2028 , RIae76208_37, \881 );
nor \U$1652 ( \2029 , \2027 , \2028 );
not \U$1653 ( \2030 , \2029 );
or \U$1654 ( \2031 , \2026 , \2030 );
or \U$1655 ( \2032 , \2029 , \787 );
nand \U$1656 ( \2033 , \2031 , \2032 );
and \U$1657 ( \2034 , \1138 , RIae76a78_55);
and \U$1658 ( \2035 , RIae76988_53, \1136 );
nor \U$1659 ( \2036 , \2034 , \2035 );
and \U$1660 ( \2037 , \2036 , \1012 );
not \U$1661 ( \2038 , \2036 );
and \U$1662 ( \2039 , \2038 , \1142 );
nor \U$1663 ( \2040 , \2037 , \2039 );
xor \U$1664 ( \2041 , \2033 , \2040 );
and \U$1665 ( \2042 , \1376 , RIae767a8_49);
and \U$1666 ( \2043 , RIae76898_51, \1374 );
nor \U$1667 ( \2044 , \2042 , \2043 );
and \U$1668 ( \2045 , \2044 , \1380 );
not \U$1669 ( \2046 , \2044 );
and \U$1670 ( \2047 , \2046 , \1261 );
nor \U$1671 ( \2048 , \2045 , \2047 );
and \U$1672 ( \2049 , \2041 , \2048 );
and \U$1673 ( \2050 , \2033 , \2040 );
or \U$1674 ( \2051 , \2049 , \2050 );
and \U$1675 ( \2052 , \1593 , RIae76b68_57);
and \U$1676 ( \2053 , RIae78a58_123, \1591 );
nor \U$1677 ( \2054 , \2052 , \2053 );
and \U$1678 ( \2055 , \2054 , \1498 );
not \U$1679 ( \2056 , \2054 );
and \U$1680 ( \2057 , \2056 , \1488 );
nor \U$1681 ( \2058 , \2055 , \2057 );
nand \U$1682 ( \2059 , RIae79520_146, RIae79a48_157);
and \U$1683 ( \2060 , \2059 , RIae79ac0_158);
not \U$1684 ( \2061 , \2060 );
xor \U$1685 ( \2062 , \2058 , \2061 );
and \U$1686 ( \2063 , \1939 , RIae78cb0_128);
and \U$1687 ( \2064 , RIae78da0_130, \1937 );
nor \U$1688 ( \2065 , \2063 , \2064 );
and \U$1689 ( \2066 , \2065 , \1735 );
not \U$1690 ( \2067 , \2065 );
and \U$1691 ( \2068 , \2067 , \1734 );
nor \U$1692 ( \2069 , \2066 , \2068 );
and \U$1693 ( \2070 , \2062 , \2069 );
and \U$1694 ( \2071 , \2058 , \2061 );
or \U$1695 ( \2072 , \2070 , \2071 );
xor \U$1696 ( \2073 , \2051 , \2072 );
and \U$1697 ( \2074 , \672 , RIae76118_35);
and \U$1698 ( \2075 , RIae76028_33, \670 );
nor \U$1699 ( \2076 , \2074 , \2075 );
and \U$1700 ( \2077 , \2076 , \588 );
not \U$1701 ( \2078 , \2076 );
and \U$1702 ( \2079 , \2078 , \587 );
nor \U$1703 ( \2080 , \2077 , \2079 );
not \U$1704 ( \2081 , \471 );
and \U$1705 ( \2082 , \514 , RIae763e8_41);
and \U$1706 ( \2083 , RIae764d8_43, \512 );
nor \U$1707 ( \2084 , \2082 , \2083 );
not \U$1708 ( \2085 , \2084 );
or \U$1709 ( \2086 , \2081 , \2085 );
or \U$1710 ( \2087 , \2084 , \471 );
nand \U$1711 ( \2088 , \2086 , \2087 );
xor \U$1712 ( \2089 , \2080 , \2088 );
and \U$1713 ( \2090 , \558 , RIae766b8_47);
and \U$1714 ( \2091 , RIae765c8_45, \556 );
nor \U$1715 ( \2092 , \2090 , \2091 );
and \U$1716 ( \2093 , \2092 , \504 );
not \U$1717 ( \2094 , \2092 );
and \U$1718 ( \2095 , \2094 , \562 );
nor \U$1719 ( \2096 , \2093 , \2095 );
and \U$1720 ( \2097 , \2089 , \2096 );
and \U$1721 ( \2098 , \2080 , \2088 );
or \U$1722 ( \2099 , \2097 , \2098 );
and \U$1723 ( \2100 , \2073 , \2099 );
and \U$1724 ( \2101 , \2051 , \2072 );
or \U$1725 ( \2102 , \2100 , \2101 );
xor \U$1726 ( \2103 , \1878 , \1886 );
xor \U$1727 ( \2104 , \2103 , \1894 );
xor \U$1728 ( \2105 , \1932 , \1944 );
xor \U$1729 ( \2106 , \2105 , \1952 );
and \U$1730 ( \2107 , \2104 , \2106 );
xor \U$1731 ( \2108 , \2102 , \2107 );
not \U$1732 ( \2109 , \388 );
and \U$1733 ( \2110 , \384 , RIae75218_3);
and \U$1734 ( \2111 , RIae75128_1, \382 );
nor \U$1735 ( \2112 , \2110 , \2111 );
not \U$1736 ( \2113 , \2112 );
or \U$1737 ( \2114 , \2109 , \2113 );
or \U$1738 ( \2115 , \2112 , \392 );
nand \U$1739 ( \2116 , \2114 , \2115 );
not \U$1740 ( \2117 , RIae756c8_13);
nor \U$1741 ( \2118 , \2117 , \491 );
xor \U$1742 ( \2119 , \2116 , \2118 );
not \U$1743 ( \2120 , \402 );
and \U$1744 ( \2121 , \436 , RIae75308_5);
and \U$1745 ( \2122 , RIae753f8_7, \434 );
nor \U$1746 ( \2123 , \2121 , \2122 );
not \U$1747 ( \2124 , \2123 );
or \U$1748 ( \2125 , \2120 , \2124 );
or \U$1749 ( \2126 , \2123 , \400 );
nand \U$1750 ( \2127 , \2125 , \2126 );
and \U$1751 ( \2128 , \2119 , \2127 );
and \U$1752 ( \2129 , \2116 , \2118 );
or \U$1753 ( \2130 , \2128 , \2129 );
or \U$1754 ( \2131 , \1978 , \1970 );
nand \U$1755 ( \2132 , \2131 , \1979 );
xor \U$1756 ( \2133 , \2130 , \2132 );
xor \U$1757 ( \2134 , \1905 , \1913 );
xor \U$1758 ( \2135 , \2134 , \1921 );
and \U$1759 ( \2136 , \2133 , \2135 );
and \U$1760 ( \2137 , \2130 , \2132 );
or \U$1761 ( \2138 , \2136 , \2137 );
and \U$1762 ( \2139 , \2108 , \2138 );
and \U$1763 ( \2140 , \2102 , \2107 );
or \U$1764 ( \2141 , \2139 , \2140 );
xor \U$1765 ( \2142 , \2025 , \2141 );
xor \U$1766 ( \2143 , \1864 , \1865 );
xor \U$1767 ( \2144 , \2143 , \1868 );
and \U$1768 ( \2145 , \2142 , \2144 );
and \U$1769 ( \2146 , \2025 , \2141 );
or \U$1770 ( \2147 , \2145 , \2146 );
xor \U$1771 ( \2148 , \1694 , \1698 );
xor \U$1772 ( \2149 , \2148 , \1777 );
xor \U$1773 ( \2150 , \2147 , \2149 );
xor \U$1774 ( \2151 , \1871 , \1998 );
xor \U$1775 ( \2152 , \2151 , \2003 );
and \U$1776 ( \2153 , \2150 , \2152 );
and \U$1777 ( \2154 , \2147 , \2149 );
or \U$1778 ( \2155 , \2153 , \2154 );
not \U$1779 ( \2156 , \2155 );
xnor \U$1780 ( \2157 , \2006 , \1859 );
not \U$1781 ( \2158 , \2157 );
not \U$1782 ( \2159 , \1856 );
and \U$1783 ( \2160 , \2158 , \2159 );
and \U$1784 ( \2161 , \2157 , \1856 );
nor \U$1785 ( \2162 , \2160 , \2161 );
nor \U$1786 ( \2163 , \2156 , \2162 );
not \U$1787 ( \2164 , \1850 );
not \U$1788 ( \2165 , \2008 );
or \U$1789 ( \2166 , \2164 , \2165 );
or \U$1790 ( \2167 , \2008 , \1850 );
nand \U$1791 ( \2168 , \2166 , \2167 );
and \U$1792 ( \2169 , \2163 , \2168 );
xor \U$1793 ( \2170 , \2168 , \2163 );
xor \U$1794 ( \2171 , \2025 , \2141 );
xor \U$1795 ( \2172 , \2171 , \2144 );
not \U$1796 ( \2173 , \2172 );
xor \U$1797 ( \2174 , \1897 , \1924 );
xor \U$1798 ( \2175 , \2174 , \1955 );
xor \U$1799 ( \2176 , \2013 , \2020 );
xor \U$1800 ( \2177 , \2175 , \2176 );
xor \U$1801 ( \2178 , \2033 , \2040 );
xor \U$1802 ( \2179 , \2178 , \2048 );
xor \U$1803 ( \2180 , \2058 , \2061 );
xor \U$1804 ( \2181 , \2180 , \2069 );
and \U$1805 ( \2182 , \2179 , \2181 );
not \U$1806 ( \2183 , \2182 );
and \U$1807 ( \2184 , \1376 , RIae76988_53);
and \U$1808 ( \2185 , RIae767a8_49, \1374 );
nor \U$1809 ( \2186 , \2184 , \2185 );
and \U$1810 ( \2187 , \2186 , \1380 );
not \U$1811 ( \2188 , \2186 );
and \U$1812 ( \2189 , \2188 , \1261 );
nor \U$1813 ( \2190 , \2187 , \2189 );
not \U$1814 ( \2191 , \787 );
and \U$1815 ( \2192 , \883 , RIae76028_33);
and \U$1816 ( \2193 , RIae762f8_39, \881 );
nor \U$1817 ( \2194 , \2192 , \2193 );
not \U$1818 ( \2195 , \2194 );
or \U$1819 ( \2196 , \2191 , \2195 );
or \U$1820 ( \2197 , \2194 , \787 );
nand \U$1821 ( \2198 , \2196 , \2197 );
xor \U$1822 ( \2199 , \2190 , \2198 );
and \U$1823 ( \2200 , \1138 , RIae76208_37);
and \U$1824 ( \2201 , RIae76a78_55, \1136 );
nor \U$1825 ( \2202 , \2200 , \2201 );
and \U$1826 ( \2203 , \2202 , \1012 );
not \U$1827 ( \2204 , \2202 );
and \U$1828 ( \2205 , \2204 , \1142 );
nor \U$1829 ( \2206 , \2203 , \2205 );
and \U$1830 ( \2207 , \2199 , \2206 );
and \U$1831 ( \2208 , \2190 , \2198 );
or \U$1832 ( \2209 , \2207 , \2208 );
and \U$1833 ( \2210 , \1593 , RIae76898_51);
and \U$1834 ( \2211 , RIae76b68_57, \1591 );
nor \U$1835 ( \2212 , \2210 , \2211 );
and \U$1836 ( \2213 , \2212 , \1498 );
not \U$1837 ( \2214 , \2212 );
and \U$1838 ( \2215 , \2214 , \1488 );
nor \U$1839 ( \2216 , \2213 , \2215 );
and \U$1840 ( \2217 , RIae79ac0_158, RIae79a48_157);
not \U$1841 ( \2218 , RIae79520_146);
and \U$1842 ( \2219 , RIae79a48_157, \2218 );
not \U$1843 ( \2220 , RIae79a48_157);
and \U$1844 ( \2221 , \2220 , RIae79520_146);
or \U$1845 ( \2222 , \2219 , \2221 );
nor \U$1846 ( \2223 , RIae79ac0_158, RIae79a48_157);
nor \U$1847 ( \2224 , \2217 , \2222 , \2223 );
nand \U$1848 ( \2225 , RIae78da0_130, \2224 );
and \U$1849 ( \2226 , \2225 , \2061 );
not \U$1850 ( \2227 , \2225 );
and \U$1851 ( \2228 , \2227 , \2060 );
nor \U$1852 ( \2229 , \2226 , \2228 );
xor \U$1853 ( \2230 , \2216 , \2229 );
and \U$1854 ( \2231 , \1939 , RIae78a58_123);
and \U$1855 ( \2232 , RIae78cb0_128, \1937 );
nor \U$1856 ( \2233 , \2231 , \2232 );
and \U$1857 ( \2234 , \2233 , \1735 );
not \U$1858 ( \2235 , \2233 );
and \U$1859 ( \2236 , \2235 , \1734 );
nor \U$1860 ( \2237 , \2234 , \2236 );
and \U$1861 ( \2238 , \2230 , \2237 );
and \U$1862 ( \2239 , \2216 , \2229 );
or \U$1863 ( \2240 , \2238 , \2239 );
xor \U$1864 ( \2241 , \2209 , \2240 );
not \U$1865 ( \2242 , \469 );
and \U$1866 ( \2243 , \514 , RIae753f8_7);
and \U$1867 ( \2244 , RIae763e8_41, \512 );
nor \U$1868 ( \2245 , \2243 , \2244 );
not \U$1869 ( \2246 , \2245 );
or \U$1870 ( \2247 , \2242 , \2246 );
or \U$1871 ( \2248 , \2245 , \471 );
nand \U$1872 ( \2249 , \2247 , \2248 );
and \U$1873 ( \2250 , \558 , RIae764d8_43);
and \U$1874 ( \2251 , RIae766b8_47, \556 );
nor \U$1875 ( \2252 , \2250 , \2251 );
and \U$1876 ( \2253 , \2252 , \504 );
not \U$1877 ( \2254 , \2252 );
and \U$1878 ( \2255 , \2254 , \562 );
nor \U$1879 ( \2256 , \2253 , \2255 );
xor \U$1880 ( \2257 , \2249 , \2256 );
and \U$1881 ( \2258 , \672 , RIae765c8_45);
and \U$1882 ( \2259 , RIae76118_35, \670 );
nor \U$1883 ( \2260 , \2258 , \2259 );
and \U$1884 ( \2261 , \2260 , \588 );
not \U$1885 ( \2262 , \2260 );
and \U$1886 ( \2263 , \2262 , \587 );
nor \U$1887 ( \2264 , \2261 , \2263 );
and \U$1888 ( \2265 , \2257 , \2264 );
and \U$1889 ( \2266 , \2249 , \2256 );
or \U$1890 ( \2267 , \2265 , \2266 );
and \U$1891 ( \2268 , \2241 , \2267 );
and \U$1892 ( \2269 , \2209 , \2240 );
or \U$1893 ( \2270 , \2268 , \2269 );
not \U$1894 ( \2271 , \2270 );
or \U$1895 ( \2272 , \2183 , \2271 );
or \U$1896 ( \2273 , \2270 , \2182 );
and \U$1897 ( \2274 , \384 , RIae756c8_13);
and \U$1898 ( \2275 , RIae75218_3, \382 );
nor \U$1899 ( \2276 , \2274 , \2275 );
not \U$1900 ( \2277 , \2276 );
not \U$1901 ( \2278 , \392 );
and \U$1902 ( \2279 , \2277 , \2278 );
and \U$1903 ( \2280 , \2276 , \392 );
nor \U$1904 ( \2281 , \2279 , \2280 );
nand \U$1905 ( \2282 , RIae757b8_15, RIae78b48_125);
or \U$1906 ( \2283 , \2281 , \2282 );
not \U$1907 ( \2284 , \2282 );
not \U$1908 ( \2285 , \2281 );
or \U$1909 ( \2286 , \2284 , \2285 );
not \U$1910 ( \2287 , \402 );
and \U$1911 ( \2288 , \436 , RIae75128_1);
and \U$1912 ( \2289 , RIae75308_5, \434 );
nor \U$1913 ( \2290 , \2288 , \2289 );
not \U$1914 ( \2291 , \2290 );
or \U$1915 ( \2292 , \2287 , \2291 );
or \U$1916 ( \2293 , \2290 , \400 );
nand \U$1917 ( \2294 , \2292 , \2293 );
nand \U$1918 ( \2295 , \2286 , \2294 );
nand \U$1919 ( \2296 , \2283 , \2295 );
xor \U$1920 ( \2297 , \2116 , \2118 );
xor \U$1921 ( \2298 , \2297 , \2127 );
and \U$1922 ( \2299 , \2296 , \2298 );
xor \U$1923 ( \2300 , \2080 , \2088 );
xor \U$1924 ( \2301 , \2300 , \2096 );
xor \U$1925 ( \2302 , \2116 , \2118 );
xor \U$1926 ( \2303 , \2302 , \2127 );
and \U$1927 ( \2304 , \2301 , \2303 );
and \U$1928 ( \2305 , \2296 , \2301 );
or \U$1929 ( \2306 , \2299 , \2304 , \2305 );
nand \U$1930 ( \2307 , \2273 , \2306 );
nand \U$1931 ( \2308 , \2272 , \2307 );
xor \U$1932 ( \2309 , \2177 , \2308 );
xor \U$1933 ( \2310 , \2104 , \2106 );
xor \U$1934 ( \2311 , \2051 , \2072 );
xor \U$1935 ( \2312 , \2311 , \2099 );
and \U$1936 ( \2313 , \2310 , \2312 );
xor \U$1937 ( \2314 , \2130 , \2132 );
xor \U$1938 ( \2315 , \2314 , \2135 );
xor \U$1939 ( \2316 , \2051 , \2072 );
xor \U$1940 ( \2317 , \2316 , \2099 );
and \U$1941 ( \2318 , \2315 , \2317 );
and \U$1942 ( \2319 , \2310 , \2315 );
or \U$1943 ( \2320 , \2313 , \2318 , \2319 );
and \U$1944 ( \2321 , \2309 , \2320 );
and \U$1945 ( \2322 , \2177 , \2308 );
nor \U$1946 ( \2323 , \2321 , \2322 );
not \U$1947 ( \2324 , \2323 );
xor \U$1948 ( \2325 , \1958 , \1982 );
xor \U$1949 ( \2326 , \2325 , \1995 );
not \U$1950 ( \2327 , \2326 );
and \U$1951 ( \2328 , \2324 , \2327 );
and \U$1952 ( \2329 , \2323 , \2326 );
nor \U$1953 ( \2330 , \2328 , \2329 );
not \U$1954 ( \2331 , \2330 );
or \U$1955 ( \2332 , \2173 , \2331 );
or \U$1956 ( \2333 , \2330 , \2172 );
nand \U$1957 ( \2334 , \2332 , \2333 );
not \U$1958 ( \2335 , \2334 );
xor \U$1959 ( \2336 , \2177 , \2308 );
xor \U$1960 ( \2337 , \2336 , \2320 );
xor \U$1961 ( \2338 , \2102 , \2107 );
xor \U$1962 ( \2339 , \2338 , \2138 );
xor \U$1963 ( \2340 , \2337 , \2339 );
xor \U$1964 ( \2341 , \2179 , \2181 );
xor \U$1965 ( \2342 , \2209 , \2240 );
xor \U$1966 ( \2343 , \2342 , \2267 );
and \U$1967 ( \2344 , \2341 , \2343 );
xor \U$1968 ( \2345 , \2116 , \2118 );
xor \U$1969 ( \2346 , \2345 , \2127 );
xor \U$1970 ( \2347 , \2296 , \2301 );
xor \U$1971 ( \2348 , \2346 , \2347 );
xor \U$1972 ( \2349 , \2209 , \2240 );
xor \U$1973 ( \2350 , \2349 , \2267 );
and \U$1974 ( \2351 , \2348 , \2350 );
and \U$1975 ( \2352 , \2341 , \2348 );
or \U$1976 ( \2353 , \2344 , \2351 , \2352 );
not \U$1977 ( \2354 , \2353 );
xor \U$1978 ( \2355 , \2051 , \2072 );
xor \U$1979 ( \2356 , \2355 , \2099 );
xor \U$1980 ( \2357 , \2310 , \2315 );
xor \U$1981 ( \2358 , \2356 , \2357 );
not \U$1982 ( \2359 , \2358 );
or \U$1983 ( \2360 , \2354 , \2359 );
or \U$1984 ( \2361 , \2358 , \2353 );
and \U$1985 ( \2362 , \672 , RIae766b8_47);
and \U$1986 ( \2363 , RIae765c8_45, \670 );
nor \U$1987 ( \2364 , \2362 , \2363 );
and \U$1988 ( \2365 , \2364 , \587 );
not \U$1989 ( \2366 , \2364 );
and \U$1990 ( \2367 , \2366 , \588 );
nor \U$1991 ( \2368 , \2365 , \2367 );
and \U$1992 ( \2369 , \883 , RIae76118_35);
and \U$1993 ( \2370 , RIae76028_33, \881 );
nor \U$1994 ( \2371 , \2369 , \2370 );
not \U$1995 ( \2372 , \2371 );
not \U$1996 ( \2373 , \789 );
and \U$1997 ( \2374 , \2372 , \2373 );
and \U$1998 ( \2375 , \2371 , \789 );
nor \U$1999 ( \2376 , \2374 , \2375 );
xor \U$2000 ( \2377 , \2368 , \2376 );
and \U$2001 ( \2378 , \558 , RIae763e8_41);
and \U$2002 ( \2379 , RIae764d8_43, \556 );
nor \U$2003 ( \2380 , \2378 , \2379 );
and \U$2004 ( \2381 , \2380 , \562 );
not \U$2005 ( \2382 , \2380 );
and \U$2006 ( \2383 , \2382 , \504 );
nor \U$2007 ( \2384 , \2381 , \2383 );
and \U$2008 ( \2385 , \2377 , \2384 );
and \U$2009 ( \2386 , \2368 , \2376 );
nor \U$2010 ( \2387 , \2385 , \2386 );
and \U$2011 ( \2388 , \1939 , RIae76b68_57);
and \U$2012 ( \2389 , RIae78a58_123, \1937 );
nor \U$2013 ( \2390 , \2388 , \2389 );
and \U$2014 ( \2391 , \2390 , \1734 );
not \U$2015 ( \2392 , \2390 );
and \U$2016 ( \2393 , \2392 , \1735 );
nor \U$2017 ( \2394 , \2391 , \2393 );
and \U$2018 ( \2395 , RIae79430_144, RIae794a8_145);
nor \U$2019 ( \2396 , \2395 , \2218 );
buf \U$2020 ( \2397 , \2396 );
or \U$2021 ( \2398 , \2394 , \2397 );
not \U$2022 ( \2399 , \2397 );
not \U$2023 ( \2400 , \2394 );
or \U$2024 ( \2401 , \2399 , \2400 );
and \U$2025 ( \2402 , \2224 , RIae78cb0_128);
and \U$2026 ( \2403 , RIae78da0_130, \2222 );
nor \U$2027 ( \2404 , \2402 , \2403 );
and \U$2028 ( \2405 , \2404 , \2061 );
not \U$2029 ( \2406 , \2404 );
and \U$2030 ( \2407 , \2406 , \2060 );
nor \U$2031 ( \2408 , \2405 , \2407 );
nand \U$2032 ( \2409 , \2401 , \2408 );
nand \U$2033 ( \2410 , \2398 , \2409 );
xor \U$2034 ( \2411 , \2387 , \2410 );
and \U$2035 ( \2412 , \1138 , RIae762f8_39);
and \U$2036 ( \2413 , RIae76208_37, \1136 );
nor \U$2037 ( \2414 , \2412 , \2413 );
and \U$2038 ( \2415 , \2414 , \1142 );
not \U$2039 ( \2416 , \2414 );
and \U$2040 ( \2417 , \2416 , \1012 );
nor \U$2041 ( \2418 , \2415 , \2417 );
and \U$2042 ( \2419 , \1376 , RIae76a78_55);
and \U$2043 ( \2420 , RIae76988_53, \1374 );
nor \U$2044 ( \2421 , \2419 , \2420 );
and \U$2045 ( \2422 , \2421 , \1261 );
not \U$2046 ( \2423 , \2421 );
and \U$2047 ( \2424 , \2423 , \1380 );
nor \U$2048 ( \2425 , \2422 , \2424 );
or \U$2049 ( \2426 , \2418 , \2425 );
not \U$2050 ( \2427 , \2425 );
not \U$2051 ( \2428 , \2418 );
or \U$2052 ( \2429 , \2427 , \2428 );
and \U$2053 ( \2430 , \1593 , RIae767a8_49);
and \U$2054 ( \2431 , RIae76898_51, \1591 );
nor \U$2055 ( \2432 , \2430 , \2431 );
and \U$2056 ( \2433 , \2432 , \1498 );
not \U$2057 ( \2434 , \2432 );
and \U$2058 ( \2435 , \2434 , \1488 );
nor \U$2059 ( \2436 , \2433 , \2435 );
nand \U$2060 ( \2437 , \2429 , \2436 );
nand \U$2061 ( \2438 , \2426 , \2437 );
and \U$2062 ( \2439 , \2411 , \2438 );
and \U$2063 ( \2440 , \2387 , \2410 );
or \U$2064 ( \2441 , \2439 , \2440 );
and \U$2065 ( \2442 , \514 , RIae75308_5);
and \U$2066 ( \2443 , RIae753f8_7, \512 );
nor \U$2067 ( \2444 , \2442 , \2443 );
not \U$2068 ( \2445 , \2444 );
not \U$2069 ( \2446 , \471 );
and \U$2070 ( \2447 , \2445 , \2446 );
and \U$2071 ( \2448 , \2444 , \469 );
nor \U$2072 ( \2449 , \2447 , \2448 );
and \U$2073 ( \2450 , \384 , RIae757b8_15);
and \U$2074 ( \2451 , RIae756c8_13, \382 );
nor \U$2075 ( \2452 , \2450 , \2451 );
not \U$2076 ( \2453 , \2452 );
not \U$2077 ( \2454 , \392 );
and \U$2078 ( \2455 , \2453 , \2454 );
and \U$2079 ( \2456 , \2452 , \392 );
nor \U$2080 ( \2457 , \2455 , \2456 );
xor \U$2081 ( \2458 , \2449 , \2457 );
and \U$2082 ( \2459 , \436 , RIae75218_3);
and \U$2083 ( \2460 , RIae75128_1, \434 );
nor \U$2084 ( \2461 , \2459 , \2460 );
not \U$2085 ( \2462 , \2461 );
not \U$2086 ( \2463 , \402 );
and \U$2087 ( \2464 , \2462 , \2463 );
and \U$2088 ( \2465 , \2461 , \400 );
nor \U$2089 ( \2466 , \2464 , \2465 );
and \U$2090 ( \2467 , \2458 , \2466 );
and \U$2091 ( \2468 , \2449 , \2457 );
or \U$2092 ( \2469 , \2467 , \2468 );
not \U$2093 ( \2470 , \2281 );
not \U$2094 ( \2471 , \2294 );
or \U$2095 ( \2472 , \2470 , \2471 );
or \U$2096 ( \2473 , \2281 , \2294 );
nand \U$2097 ( \2474 , \2472 , \2473 );
not \U$2098 ( \2475 , \2474 );
not \U$2099 ( \2476 , \2282 );
and \U$2100 ( \2477 , \2475 , \2476 );
and \U$2101 ( \2478 , \2474 , \2282 );
nor \U$2102 ( \2479 , \2477 , \2478 );
nand \U$2103 ( \2480 , \2469 , \2479 );
xor \U$2104 ( \2481 , \2441 , \2480 );
xor \U$2105 ( \2482 , \2216 , \2229 );
xor \U$2106 ( \2483 , \2482 , \2237 );
xor \U$2107 ( \2484 , \2249 , \2256 );
xor \U$2108 ( \2485 , \2484 , \2264 );
and \U$2109 ( \2486 , \2483 , \2485 );
xor \U$2110 ( \2487 , \2190 , \2198 );
xor \U$2111 ( \2488 , \2487 , \2206 );
xor \U$2112 ( \2489 , \2249 , \2256 );
xor \U$2113 ( \2490 , \2489 , \2264 );
and \U$2114 ( \2491 , \2488 , \2490 );
and \U$2115 ( \2492 , \2483 , \2488 );
or \U$2116 ( \2493 , \2486 , \2491 , \2492 );
and \U$2117 ( \2494 , \2481 , \2493 );
and \U$2118 ( \2495 , \2441 , \2480 );
or \U$2119 ( \2496 , \2494 , \2495 );
nand \U$2120 ( \2497 , \2361 , \2496 );
nand \U$2121 ( \2498 , \2360 , \2497 );
and \U$2122 ( \2499 , \2340 , \2498 );
and \U$2123 ( \2500 , \2337 , \2339 );
nor \U$2124 ( \2501 , \2499 , \2500 );
not \U$2125 ( \2502 , \2501 );
and \U$2126 ( \2503 , \2335 , \2502 );
and \U$2127 ( \2504 , \2334 , \2501 );
nor \U$2128 ( \2505 , \2503 , \2504 );
or \U$2129 ( \2506 , \2479 , \2469 );
nand \U$2130 ( \2507 , \2506 , \2480 );
xor \U$2131 ( \2508 , \2387 , \2410 );
xor \U$2132 ( \2509 , \2508 , \2438 );
and \U$2133 ( \2510 , \2507 , \2509 );
xor \U$2134 ( \2511 , \2249 , \2256 );
xor \U$2135 ( \2512 , \2511 , \2264 );
xor \U$2136 ( \2513 , \2483 , \2488 );
xor \U$2137 ( \2514 , \2512 , \2513 );
xor \U$2138 ( \2515 , \2387 , \2410 );
xor \U$2139 ( \2516 , \2515 , \2438 );
and \U$2140 ( \2517 , \2514 , \2516 );
and \U$2141 ( \2518 , \2507 , \2514 );
or \U$2142 ( \2519 , \2510 , \2517 , \2518 );
nand \U$2143 ( \2520 , RIae755d8_11, RIae78b48_125);
nand \U$2144 ( \2521 , RIae754e8_9, RIae78b48_125);
xor \U$2145 ( \2522 , \2520 , \2521 );
and \U$2146 ( \2523 , \384 , RIae754e8_9);
and \U$2147 ( \2524 , RIae757b8_15, \382 );
nor \U$2148 ( \2525 , \2523 , \2524 );
not \U$2149 ( \2526 , \2525 );
not \U$2150 ( \2527 , \388 );
and \U$2151 ( \2528 , \2526 , \2527 );
and \U$2152 ( \2529 , \2525 , \392 );
nor \U$2153 ( \2530 , \2528 , \2529 );
not \U$2154 ( \2531 , \2530 );
and \U$2155 ( \2532 , \436 , RIae756c8_13);
and \U$2156 ( \2533 , RIae75218_3, \434 );
nor \U$2157 ( \2534 , \2532 , \2533 );
not \U$2158 ( \2535 , \2534 );
not \U$2159 ( \2536 , \402 );
and \U$2160 ( \2537 , \2535 , \2536 );
and \U$2161 ( \2538 , \2534 , \400 );
nor \U$2162 ( \2539 , \2537 , \2538 );
not \U$2163 ( \2540 , \2539 );
and \U$2164 ( \2541 , \2531 , \2540 );
and \U$2165 ( \2542 , \2539 , \2530 );
and \U$2166 ( \2543 , \514 , RIae75128_1);
and \U$2167 ( \2544 , RIae75308_5, \512 );
nor \U$2168 ( \2545 , \2543 , \2544 );
not \U$2169 ( \2546 , \2545 );
not \U$2170 ( \2547 , \469 );
and \U$2171 ( \2548 , \2546 , \2547 );
and \U$2172 ( \2549 , \2545 , \469 );
nor \U$2173 ( \2550 , \2548 , \2549 );
nor \U$2174 ( \2551 , \2542 , \2550 );
nor \U$2175 ( \2552 , \2541 , \2551 );
and \U$2176 ( \2553 , \2522 , \2552 );
and \U$2177 ( \2554 , \2520 , \2521 );
or \U$2178 ( \2555 , \2553 , \2554 );
and \U$2179 ( \2556 , \672 , RIae764d8_43);
and \U$2180 ( \2557 , RIae766b8_47, \670 );
nor \U$2181 ( \2558 , \2556 , \2557 );
and \U$2182 ( \2559 , \2558 , \588 );
not \U$2183 ( \2560 , \2558 );
and \U$2184 ( \2561 , \2560 , \587 );
nor \U$2185 ( \2562 , \2559 , \2561 );
not \U$2186 ( \2563 , \789 );
and \U$2187 ( \2564 , \883 , RIae765c8_45);
and \U$2188 ( \2565 , RIae76118_35, \881 );
nor \U$2189 ( \2566 , \2564 , \2565 );
not \U$2190 ( \2567 , \2566 );
or \U$2191 ( \2568 , \2563 , \2567 );
or \U$2192 ( \2569 , \2566 , \789 );
nand \U$2193 ( \2570 , \2568 , \2569 );
xor \U$2194 ( \2571 , \2562 , \2570 );
and \U$2195 ( \2572 , \558 , RIae753f8_7);
and \U$2196 ( \2573 , RIae763e8_41, \556 );
nor \U$2197 ( \2574 , \2572 , \2573 );
and \U$2198 ( \2575 , \2574 , \504 );
not \U$2199 ( \2576 , \2574 );
and \U$2200 ( \2577 , \2576 , \562 );
nor \U$2201 ( \2578 , \2575 , \2577 );
and \U$2202 ( \2579 , \2571 , \2578 );
and \U$2203 ( \2580 , \2562 , \2570 );
nor \U$2204 ( \2581 , \2579 , \2580 );
and \U$2205 ( \2582 , \1939 , RIae76898_51);
and \U$2206 ( \2583 , RIae76b68_57, \1937 );
nor \U$2207 ( \2584 , \2582 , \2583 );
and \U$2208 ( \2585 , \2584 , \1734 );
not \U$2209 ( \2586 , \2584 );
and \U$2210 ( \2587 , \2586 , \1735 );
nor \U$2211 ( \2588 , \2585 , \2587 );
not \U$2212 ( \2589 , \2588 );
and \U$2213 ( \2590 , \2224 , RIae78a58_123);
and \U$2214 ( \2591 , RIae78cb0_128, \2222 );
nor \U$2215 ( \2592 , \2590 , \2591 );
and \U$2216 ( \2593 , \2592 , \2060 );
not \U$2217 ( \2594 , \2592 );
and \U$2218 ( \2595 , \2594 , \2061 );
nor \U$2219 ( \2596 , \2593 , \2595 );
not \U$2220 ( \2597 , \2596 );
and \U$2221 ( \2598 , \2589 , \2597 );
and \U$2222 ( \2599 , \2596 , \2588 );
and \U$2223 ( \2600 , RIae79520_146, RIae79430_144);
not \U$2224 ( \2601 , RIae79430_144);
nor \U$2225 ( \2602 , \2601 , RIae794a8_145);
not \U$2226 ( \2603 , RIae794a8_145);
nor \U$2227 ( \2604 , \2603 , RIae79430_144);
or \U$2228 ( \2605 , \2602 , \2604 );
nor \U$2229 ( \2606 , RIae79520_146, RIae79430_144);
nor \U$2230 ( \2607 , \2600 , \2605 , \2606 );
nand \U$2231 ( \2608 , RIae78da0_130, \2607 );
and \U$2232 ( \2609 , \2608 , \2397 );
not \U$2233 ( \2610 , \2608 );
not \U$2234 ( \2611 , \2396 );
and \U$2235 ( \2612 , \2610 , \2611 );
nor \U$2236 ( \2613 , \2609 , \2612 );
nor \U$2237 ( \2614 , \2599 , \2613 );
nor \U$2238 ( \2615 , \2598 , \2614 );
xor \U$2239 ( \2616 , \2581 , \2615 );
and \U$2240 ( \2617 , \1138 , RIae76028_33);
and \U$2241 ( \2618 , RIae762f8_39, \1136 );
nor \U$2242 ( \2619 , \2617 , \2618 );
and \U$2243 ( \2620 , \2619 , \1142 );
not \U$2244 ( \2621 , \2619 );
and \U$2245 ( \2622 , \2621 , \1012 );
nor \U$2246 ( \2623 , \2620 , \2622 );
not \U$2247 ( \2624 , \2623 );
and \U$2248 ( \2625 , \1376 , RIae76208_37);
and \U$2249 ( \2626 , RIae76a78_55, \1374 );
nor \U$2250 ( \2627 , \2625 , \2626 );
and \U$2251 ( \2628 , \2627 , \1261 );
not \U$2252 ( \2629 , \2627 );
and \U$2253 ( \2630 , \2629 , \1380 );
nor \U$2254 ( \2631 , \2628 , \2630 );
not \U$2255 ( \2632 , \2631 );
and \U$2256 ( \2633 , \2624 , \2632 );
and \U$2257 ( \2634 , \2631 , \2623 );
and \U$2258 ( \2635 , \1593 , RIae76988_53);
and \U$2259 ( \2636 , RIae767a8_49, \1591 );
nor \U$2260 ( \2637 , \2635 , \2636 );
and \U$2261 ( \2638 , \2637 , \1488 );
not \U$2262 ( \2639 , \2637 );
and \U$2263 ( \2640 , \2639 , \1498 );
nor \U$2264 ( \2641 , \2638 , \2640 );
nor \U$2265 ( \2642 , \2634 , \2641 );
nor \U$2266 ( \2643 , \2633 , \2642 );
and \U$2267 ( \2644 , \2616 , \2643 );
and \U$2268 ( \2645 , \2581 , \2615 );
or \U$2269 ( \2646 , \2644 , \2645 );
xor \U$2270 ( \2647 , \2555 , \2646 );
xor \U$2271 ( \2648 , \2368 , \2376 );
xor \U$2272 ( \2649 , \2648 , \2384 );
xor \U$2273 ( \2650 , \2449 , \2457 );
xor \U$2274 ( \2651 , \2650 , \2466 );
xor \U$2275 ( \2652 , \2649 , \2651 );
not \U$2276 ( \2653 , \2425 );
not \U$2277 ( \2654 , \2436 );
or \U$2278 ( \2655 , \2653 , \2654 );
or \U$2279 ( \2656 , \2425 , \2436 );
nand \U$2280 ( \2657 , \2655 , \2656 );
not \U$2281 ( \2658 , \2657 );
not \U$2282 ( \2659 , \2418 );
and \U$2283 ( \2660 , \2658 , \2659 );
and \U$2284 ( \2661 , \2657 , \2418 );
nor \U$2285 ( \2662 , \2660 , \2661 );
and \U$2286 ( \2663 , \2652 , \2662 );
and \U$2287 ( \2664 , \2649 , \2651 );
or \U$2288 ( \2665 , \2663 , \2664 );
and \U$2289 ( \2666 , \2647 , \2665 );
and \U$2290 ( \2667 , \2555 , \2646 );
nor \U$2291 ( \2668 , \2666 , \2667 );
xor \U$2292 ( \2669 , \2519 , \2668 );
xor \U$2293 ( \2670 , \2209 , \2240 );
xor \U$2294 ( \2671 , \2670 , \2267 );
xor \U$2295 ( \2672 , \2341 , \2348 );
xor \U$2296 ( \2673 , \2671 , \2672 );
and \U$2297 ( \2674 , \2669 , \2673 );
and \U$2298 ( \2675 , \2519 , \2668 );
nor \U$2299 ( \2676 , \2674 , \2675 );
xnor \U$2300 ( \2677 , \2270 , \2306 );
not \U$2301 ( \2678 , \2677 );
not \U$2302 ( \2679 , \2182 );
and \U$2303 ( \2680 , \2678 , \2679 );
and \U$2304 ( \2681 , \2677 , \2182 );
nor \U$2305 ( \2682 , \2680 , \2681 );
xor \U$2306 ( \2683 , \2676 , \2682 );
xnor \U$2307 ( \2684 , \2496 , \2353 );
not \U$2308 ( \2685 , \2684 );
not \U$2309 ( \2686 , \2358 );
and \U$2310 ( \2687 , \2685 , \2686 );
and \U$2311 ( \2688 , \2684 , \2358 );
nor \U$2312 ( \2689 , \2687 , \2688 );
and \U$2313 ( \2690 , \2683 , \2689 );
and \U$2314 ( \2691 , \2676 , \2682 );
or \U$2315 ( \2692 , \2690 , \2691 );
not \U$2316 ( \2693 , \2692 );
xor \U$2317 ( \2694 , \2337 , \2339 );
xor \U$2318 ( \2695 , \2694 , \2498 );
nand \U$2319 ( \2696 , \2693 , \2695 );
or \U$2320 ( \2697 , \2505 , \2696 );
xnor \U$2321 ( \2698 , \2696 , \2505 );
and \U$2322 ( \2699 , \436 , RIae755d8_11);
and \U$2323 ( \2700 , RIae754e8_9, \434 );
nor \U$2324 ( \2701 , \2699 , \2700 );
not \U$2325 ( \2702 , \2701 );
not \U$2326 ( \2703 , \402 );
and \U$2327 ( \2704 , \2702 , \2703 );
and \U$2328 ( \2705 , \2701 , \402 );
nor \U$2329 ( \2706 , \2704 , \2705 );
nand \U$2330 ( \2707 , RIae75e48_29, RIae78b48_125);
or \U$2331 ( \2708 , \2706 , \2707 );
not \U$2332 ( \2709 , \2707 );
not \U$2333 ( \2710 , \2706 );
or \U$2334 ( \2711 , \2709 , \2710 );
not \U$2335 ( \2712 , \392 );
and \U$2336 ( \2713 , \384 , RIae75c68_25);
and \U$2337 ( \2714 , RIae75d58_27, \382 );
nor \U$2338 ( \2715 , \2713 , \2714 );
not \U$2339 ( \2716 , \2715 );
or \U$2340 ( \2717 , \2712 , \2716 );
or \U$2341 ( \2718 , \2715 , \392 );
nand \U$2342 ( \2719 , \2717 , \2718 );
nand \U$2343 ( \2720 , \2711 , \2719 );
nand \U$2344 ( \2721 , \2708 , \2720 );
and \U$2345 ( \2722 , \384 , RIae75d58_27);
and \U$2346 ( \2723 , RIae755d8_11, \382 );
nor \U$2347 ( \2724 , \2722 , \2723 );
not \U$2348 ( \2725 , \2724 );
not \U$2349 ( \2726 , \392 );
and \U$2350 ( \2727 , \2725 , \2726 );
and \U$2351 ( \2728 , \2724 , \388 );
nor \U$2352 ( \2729 , \2727 , \2728 );
nand \U$2353 ( \2730 , RIae75c68_25, RIae78b48_125);
or \U$2354 ( \2731 , \2729 , \2730 );
nand \U$2355 ( \2732 , \2730 , \2729 );
nand \U$2356 ( \2733 , \2731 , \2732 );
xor \U$2357 ( \2734 , \2721 , \2733 );
and \U$2358 ( \2735 , \514 , RIae757b8_15);
and \U$2359 ( \2736 , RIae756c8_13, \512 );
nor \U$2360 ( \2737 , \2735 , \2736 );
not \U$2361 ( \2738 , \2737 );
not \U$2362 ( \2739 , \469 );
and \U$2363 ( \2740 , \2738 , \2739 );
and \U$2364 ( \2741 , \2737 , \471 );
nor \U$2365 ( \2742 , \2740 , \2741 );
and \U$2366 ( \2743 , \558 , RIae75218_3);
and \U$2367 ( \2744 , RIae75128_1, \556 );
nor \U$2368 ( \2745 , \2743 , \2744 );
and \U$2369 ( \2746 , \2745 , \562 );
not \U$2370 ( \2747 , \2745 );
and \U$2371 ( \2748 , \2747 , \504 );
nor \U$2372 ( \2749 , \2746 , \2748 );
or \U$2373 ( \2750 , \2742 , \2749 );
not \U$2374 ( \2751 , \2749 );
not \U$2375 ( \2752 , \2742 );
or \U$2376 ( \2753 , \2751 , \2752 );
and \U$2377 ( \2754 , \672 , RIae75308_5);
and \U$2378 ( \2755 , RIae753f8_7, \670 );
nor \U$2379 ( \2756 , \2754 , \2755 );
and \U$2380 ( \2757 , \2756 , \588 );
not \U$2381 ( \2758 , \2756 );
and \U$2382 ( \2759 , \2758 , \587 );
nor \U$2383 ( \2760 , \2757 , \2759 );
nand \U$2384 ( \2761 , \2753 , \2760 );
nand \U$2385 ( \2762 , \2750 , \2761 );
and \U$2386 ( \2763 , \2734 , \2762 );
and \U$2387 ( \2764 , \2721 , \2733 );
or \U$2388 ( \2765 , \2763 , \2764 );
and \U$2389 ( \2766 , \2607 , RIae76b68_57);
and \U$2390 ( \2767 , RIae78a58_123, \2605 );
nor \U$2391 ( \2768 , \2766 , \2767 );
and \U$2392 ( \2769 , \2768 , \2397 );
not \U$2393 ( \2770 , \2768 );
and \U$2394 ( \2771 , \2770 , \2611 );
nor \U$2395 ( \2772 , \2769 , \2771 );
nand \U$2396 ( \2773 , RIae797f0_152, RIae79868_153);
and \U$2397 ( \2774 , \2773 , RIae798e0_154);
xor \U$2398 ( \2775 , \2772 , \2774 );
and \U$2399 ( \2776 , RIae794a8_145, RIae79958_155);
not \U$2400 ( \2777 , RIae79958_155);
nor \U$2401 ( \2778 , \2777 , RIae798e0_154);
not \U$2402 ( \2779 , RIae798e0_154);
nor \U$2403 ( \2780 , \2779 , RIae79958_155);
or \U$2404 ( \2781 , \2778 , \2780 );
nor \U$2405 ( \2782 , RIae794a8_145, RIae79958_155);
nor \U$2406 ( \2783 , \2776 , \2781 , \2782 );
and \U$2407 ( \2784 , \2783 , RIae78cb0_128);
and \U$2408 ( \2785 , RIae78da0_130, \2781 );
nor \U$2409 ( \2786 , \2784 , \2785 );
not \U$2410 ( \2787 , \2786 );
nand \U$2411 ( \2788 , RIae798e0_154, RIae79958_155);
and \U$2412 ( \2789 , \2788 , RIae794a8_145);
not \U$2413 ( \2790 , \2789 );
and \U$2414 ( \2791 , \2787 , \2790 );
and \U$2415 ( \2792 , \2786 , \2789 );
nor \U$2416 ( \2793 , \2791 , \2792 );
and \U$2417 ( \2794 , \2775 , \2793 );
and \U$2418 ( \2795 , \2772 , \2774 );
or \U$2419 ( \2796 , \2794 , \2795 );
and \U$2420 ( \2797 , \2224 , RIae767a8_49);
and \U$2421 ( \2798 , RIae76898_51, \2222 );
nor \U$2422 ( \2799 , \2797 , \2798 );
and \U$2423 ( \2800 , \2799 , \2060 );
not \U$2424 ( \2801 , \2799 );
and \U$2425 ( \2802 , \2801 , \2061 );
nor \U$2426 ( \2803 , \2800 , \2802 );
and \U$2427 ( \2804 , \1593 , RIae762f8_39);
and \U$2428 ( \2805 , RIae76208_37, \1591 );
nor \U$2429 ( \2806 , \2804 , \2805 );
and \U$2430 ( \2807 , \2806 , \1488 );
not \U$2431 ( \2808 , \2806 );
and \U$2432 ( \2809 , \2808 , \1498 );
nor \U$2433 ( \2810 , \2807 , \2809 );
xor \U$2434 ( \2811 , \2803 , \2810 );
and \U$2435 ( \2812 , \1939 , RIae76a78_55);
and \U$2436 ( \2813 , RIae76988_53, \1937 );
nor \U$2437 ( \2814 , \2812 , \2813 );
and \U$2438 ( \2815 , \2814 , \1734 );
not \U$2439 ( \2816 , \2814 );
and \U$2440 ( \2817 , \2816 , \1735 );
nor \U$2441 ( \2818 , \2815 , \2817 );
and \U$2442 ( \2819 , \2811 , \2818 );
and \U$2443 ( \2820 , \2803 , \2810 );
or \U$2444 ( \2821 , \2819 , \2820 );
xor \U$2445 ( \2822 , \2796 , \2821 );
and \U$2446 ( \2823 , \1138 , RIae766b8_47);
and \U$2447 ( \2824 , RIae765c8_45, \1136 );
nor \U$2448 ( \2825 , \2823 , \2824 );
and \U$2449 ( \2826 , \2825 , \1142 );
not \U$2450 ( \2827 , \2825 );
and \U$2451 ( \2828 , \2827 , \1012 );
nor \U$2452 ( \2829 , \2826 , \2828 );
and \U$2453 ( \2830 , \883 , RIae763e8_41);
and \U$2454 ( \2831 , RIae764d8_43, \881 );
nor \U$2455 ( \2832 , \2830 , \2831 );
not \U$2456 ( \2833 , \2832 );
not \U$2457 ( \2834 , \787 );
and \U$2458 ( \2835 , \2833 , \2834 );
and \U$2459 ( \2836 , \2832 , \787 );
nor \U$2460 ( \2837 , \2835 , \2836 );
xor \U$2461 ( \2838 , \2829 , \2837 );
and \U$2462 ( \2839 , \1376 , RIae76118_35);
and \U$2463 ( \2840 , RIae76028_33, \1374 );
nor \U$2464 ( \2841 , \2839 , \2840 );
and \U$2465 ( \2842 , \2841 , \1261 );
not \U$2466 ( \2843 , \2841 );
and \U$2467 ( \2844 , \2843 , \1380 );
nor \U$2468 ( \2845 , \2842 , \2844 );
and \U$2469 ( \2846 , \2838 , \2845 );
and \U$2470 ( \2847 , \2829 , \2837 );
or \U$2471 ( \2848 , \2846 , \2847 );
and \U$2472 ( \2849 , \2822 , \2848 );
and \U$2473 ( \2850 , \2796 , \2821 );
nor \U$2474 ( \2851 , \2849 , \2850 );
xor \U$2475 ( \2852 , \2765 , \2851 );
and \U$2476 ( \2853 , \1138 , RIae765c8_45);
and \U$2477 ( \2854 , RIae76118_35, \1136 );
nor \U$2478 ( \2855 , \2853 , \2854 );
and \U$2479 ( \2856 , \2855 , \1012 );
not \U$2480 ( \2857 , \2855 );
and \U$2481 ( \2858 , \2857 , \1142 );
nor \U$2482 ( \2859 , \2856 , \2858 );
and \U$2483 ( \2860 , \672 , RIae753f8_7);
and \U$2484 ( \2861 , RIae763e8_41, \670 );
nor \U$2485 ( \2862 , \2860 , \2861 );
and \U$2486 ( \2863 , \2862 , \588 );
not \U$2487 ( \2864 , \2862 );
and \U$2488 ( \2865 , \2864 , \587 );
nor \U$2489 ( \2866 , \2863 , \2865 );
xor \U$2490 ( \2867 , \2859 , \2866 );
not \U$2491 ( \2868 , \789 );
and \U$2492 ( \2869 , \883 , RIae764d8_43);
and \U$2493 ( \2870 , RIae766b8_47, \881 );
nor \U$2494 ( \2871 , \2869 , \2870 );
not \U$2495 ( \2872 , \2871 );
or \U$2496 ( \2873 , \2868 , \2872 );
or \U$2497 ( \2874 , \2871 , \789 );
nand \U$2498 ( \2875 , \2873 , \2874 );
xor \U$2499 ( \2876 , \2867 , \2875 );
and \U$2500 ( \2877 , \558 , RIae75128_1);
and \U$2501 ( \2878 , RIae75308_5, \556 );
nor \U$2502 ( \2879 , \2877 , \2878 );
and \U$2503 ( \2880 , \2879 , \504 );
not \U$2504 ( \2881 , \2879 );
and \U$2505 ( \2882 , \2881 , \562 );
nor \U$2506 ( \2883 , \2880 , \2882 );
not \U$2507 ( \2884 , \402 );
and \U$2508 ( \2885 , \436 , RIae754e8_9);
and \U$2509 ( \2886 , RIae757b8_15, \434 );
nor \U$2510 ( \2887 , \2885 , \2886 );
not \U$2511 ( \2888 , \2887 );
or \U$2512 ( \2889 , \2884 , \2888 );
or \U$2513 ( \2890 , \2887 , \402 );
nand \U$2514 ( \2891 , \2889 , \2890 );
xor \U$2515 ( \2892 , \2883 , \2891 );
not \U$2516 ( \2893 , \469 );
and \U$2517 ( \2894 , \514 , RIae756c8_13);
and \U$2518 ( \2895 , RIae75218_3, \512 );
nor \U$2519 ( \2896 , \2894 , \2895 );
not \U$2520 ( \2897 , \2896 );
or \U$2521 ( \2898 , \2893 , \2897 );
or \U$2522 ( \2899 , \2896 , \471 );
nand \U$2523 ( \2900 , \2898 , \2899 );
xor \U$2524 ( \2901 , \2892 , \2900 );
and \U$2525 ( \2902 , \2876 , \2901 );
and \U$2526 ( \2903 , \1376 , RIae76028_33);
and \U$2527 ( \2904 , RIae762f8_39, \1374 );
nor \U$2528 ( \2905 , \2903 , \2904 );
and \U$2529 ( \2906 , \2905 , \1261 );
not \U$2530 ( \2907 , \2905 );
and \U$2531 ( \2908 , \2907 , \1380 );
nor \U$2532 ( \2909 , \2906 , \2908 );
not \U$2533 ( \2910 , \2909 );
and \U$2534 ( \2911 , \1593 , RIae76208_37);
and \U$2535 ( \2912 , RIae76a78_55, \1591 );
nor \U$2536 ( \2913 , \2911 , \2912 );
and \U$2537 ( \2914 , \2913 , \1488 );
not \U$2538 ( \2915 , \2913 );
and \U$2539 ( \2916 , \2915 , \1498 );
nor \U$2540 ( \2917 , \2914 , \2916 );
and \U$2541 ( \2918 , \1939 , RIae76988_53);
and \U$2542 ( \2919 , RIae767a8_49, \1937 );
nor \U$2543 ( \2920 , \2918 , \2919 );
and \U$2544 ( \2921 , \2920 , \1734 );
not \U$2545 ( \2922 , \2920 );
and \U$2546 ( \2923 , \2922 , \1735 );
nor \U$2547 ( \2924 , \2921 , \2923 );
xor \U$2548 ( \2925 , \2917 , \2924 );
not \U$2549 ( \2926 , \2925 );
or \U$2550 ( \2927 , \2910 , \2926 );
or \U$2551 ( \2928 , \2925 , \2909 );
nand \U$2552 ( \2929 , \2927 , \2928 );
xor \U$2553 ( \2930 , \2883 , \2891 );
xor \U$2554 ( \2931 , \2930 , \2900 );
and \U$2555 ( \2932 , \2929 , \2931 );
and \U$2556 ( \2933 , \2876 , \2929 );
or \U$2557 ( \2934 , \2902 , \2932 , \2933 );
and \U$2558 ( \2935 , \2852 , \2934 );
and \U$2559 ( \2936 , \2765 , \2851 );
or \U$2560 ( \2937 , \2935 , \2936 );
not \U$2561 ( \2938 , \2789 );
and \U$2562 ( \2939 , \2607 , RIae78cb0_128);
and \U$2563 ( \2940 , RIae78da0_130, \2605 );
nor \U$2564 ( \2941 , \2939 , \2940 );
and \U$2565 ( \2942 , \2941 , \2611 );
not \U$2566 ( \2943 , \2941 );
and \U$2567 ( \2944 , \2943 , \2397 );
nor \U$2568 ( \2945 , \2942 , \2944 );
not \U$2569 ( \2946 , \2945 );
or \U$2570 ( \2947 , \2938 , \2946 );
or \U$2571 ( \2948 , \2945 , \2789 );
nand \U$2572 ( \2949 , \2947 , \2948 );
not \U$2573 ( \2950 , \2949 );
and \U$2574 ( \2951 , \2224 , RIae76b68_57);
and \U$2575 ( \2952 , RIae78a58_123, \2222 );
nor \U$2576 ( \2953 , \2951 , \2952 );
and \U$2577 ( \2954 , \2953 , \2060 );
not \U$2578 ( \2955 , \2953 );
and \U$2579 ( \2956 , \2955 , \2061 );
nor \U$2580 ( \2957 , \2954 , \2956 );
not \U$2581 ( \2958 , \2957 );
and \U$2582 ( \2959 , \2950 , \2958 );
and \U$2583 ( \2960 , \2949 , \2957 );
nor \U$2584 ( \2961 , \2959 , \2960 );
and \U$2585 ( \2962 , \1593 , RIae76a78_55);
and \U$2586 ( \2963 , RIae76988_53, \1591 );
nor \U$2587 ( \2964 , \2962 , \2963 );
and \U$2588 ( \2965 , \2964 , \1488 );
not \U$2589 ( \2966 , \2964 );
and \U$2590 ( \2967 , \2966 , \1498 );
nor \U$2591 ( \2968 , \2965 , \2967 );
not \U$2592 ( \2969 , \2968 );
and \U$2593 ( \2970 , \1939 , RIae767a8_49);
and \U$2594 ( \2971 , RIae76898_51, \1937 );
nor \U$2595 ( \2972 , \2970 , \2971 );
and \U$2596 ( \2973 , \2972 , \1735 );
not \U$2597 ( \2974 , \2972 );
and \U$2598 ( \2975 , \2974 , \1734 );
nor \U$2599 ( \2976 , \2973 , \2975 );
not \U$2600 ( \2977 , \2976 );
or \U$2601 ( \2978 , \2969 , \2977 );
or \U$2602 ( \2979 , \2968 , \2976 );
nand \U$2603 ( \2980 , \2978 , \2979 );
not \U$2604 ( \2981 , \2980 );
and \U$2605 ( \2982 , \1376 , RIae762f8_39);
and \U$2606 ( \2983 , RIae76208_37, \1374 );
nor \U$2607 ( \2984 , \2982 , \2983 );
and \U$2608 ( \2985 , \2984 , \1261 );
not \U$2609 ( \2986 , \2984 );
and \U$2610 ( \2987 , \2986 , \1380 );
nor \U$2611 ( \2988 , \2985 , \2987 );
not \U$2612 ( \2989 , \2988 );
and \U$2613 ( \2990 , \2981 , \2989 );
and \U$2614 ( \2991 , \2980 , \2988 );
nor \U$2615 ( \2992 , \2990 , \2991 );
or \U$2616 ( \2993 , \2961 , \2992 );
and \U$2617 ( \2994 , \2961 , \2992 );
and \U$2618 ( \2995 , \514 , RIae75218_3);
and \U$2619 ( \2996 , RIae75128_1, \512 );
nor \U$2620 ( \2997 , \2995 , \2996 );
not \U$2621 ( \2998 , \2997 );
not \U$2622 ( \2999 , \469 );
and \U$2623 ( \3000 , \2998 , \2999 );
and \U$2624 ( \3001 , \2997 , \471 );
nor \U$2625 ( \3002 , \3000 , \3001 );
not \U$2626 ( \3003 , \3002 );
and \U$2627 ( \3004 , \558 , RIae75308_5);
and \U$2628 ( \3005 , RIae753f8_7, \556 );
nor \U$2629 ( \3006 , \3004 , \3005 );
and \U$2630 ( \3007 , \3006 , \504 );
not \U$2631 ( \3008 , \3006 );
and \U$2632 ( \3009 , \3008 , \562 );
nor \U$2633 ( \3010 , \3007 , \3009 );
not \U$2634 ( \3011 , \3010 );
or \U$2635 ( \3012 , \3003 , \3011 );
or \U$2636 ( \3013 , \3002 , \3010 );
nand \U$2637 ( \3014 , \3012 , \3013 );
not \U$2638 ( \3015 , \3014 );
and \U$2639 ( \3016 , \436 , RIae757b8_15);
and \U$2640 ( \3017 , RIae756c8_13, \434 );
nor \U$2641 ( \3018 , \3016 , \3017 );
not \U$2642 ( \3019 , \3018 );
not \U$2643 ( \3020 , \400 );
and \U$2644 ( \3021 , \3019 , \3020 );
and \U$2645 ( \3022 , \3018 , \402 );
nor \U$2646 ( \3023 , \3021 , \3022 );
not \U$2647 ( \3024 , \3023 );
and \U$2648 ( \3025 , \3015 , \3024 );
and \U$2649 ( \3026 , \3014 , \3023 );
nor \U$2650 ( \3027 , \3025 , \3026 );
nand \U$2651 ( \3028 , RIae75d58_27, RIae78b48_125);
xor \U$2652 ( \3029 , \3027 , \3028 );
and \U$2653 ( \3030 , \883 , RIae766b8_47);
and \U$2654 ( \3031 , RIae765c8_45, \881 );
nor \U$2655 ( \3032 , \3030 , \3031 );
not \U$2656 ( \3033 , \3032 );
not \U$2657 ( \3034 , \789 );
and \U$2658 ( \3035 , \3033 , \3034 );
and \U$2659 ( \3036 , \3032 , \787 );
nor \U$2660 ( \3037 , \3035 , \3036 );
not \U$2661 ( \3038 , \3037 );
and \U$2662 ( \3039 , \1138 , RIae76118_35);
and \U$2663 ( \3040 , RIae76028_33, \1136 );
nor \U$2664 ( \3041 , \3039 , \3040 );
and \U$2665 ( \3042 , \3041 , \1012 );
not \U$2666 ( \3043 , \3041 );
and \U$2667 ( \3044 , \3043 , \1142 );
nor \U$2668 ( \3045 , \3042 , \3044 );
not \U$2669 ( \3046 , \3045 );
or \U$2670 ( \3047 , \3038 , \3046 );
or \U$2671 ( \3048 , \3037 , \3045 );
nand \U$2672 ( \3049 , \3047 , \3048 );
not \U$2673 ( \3050 , \3049 );
and \U$2674 ( \3051 , \672 , RIae763e8_41);
and \U$2675 ( \3052 , RIae764d8_43, \670 );
nor \U$2676 ( \3053 , \3051 , \3052 );
and \U$2677 ( \3054 , \3053 , \587 );
not \U$2678 ( \3055 , \3053 );
and \U$2679 ( \3056 , \3055 , \588 );
nor \U$2680 ( \3057 , \3054 , \3056 );
not \U$2681 ( \3058 , \3057 );
and \U$2682 ( \3059 , \3050 , \3058 );
and \U$2683 ( \3060 , \3049 , \3057 );
nor \U$2684 ( \3061 , \3059 , \3060 );
xor \U$2685 ( \3062 , \3029 , \3061 );
nor \U$2686 ( \3063 , \2994 , \3062 );
not \U$2687 ( \3064 , \3063 );
nand \U$2688 ( \3065 , \2993 , \3064 );
xor \U$2689 ( \3066 , \2937 , \3065 );
or \U$2690 ( \3067 , \3023 , \3002 );
not \U$2691 ( \3068 , \3002 );
not \U$2692 ( \3069 , \3023 );
or \U$2693 ( \3070 , \3068 , \3069 );
nand \U$2694 ( \3071 , \3070 , \3010 );
nand \U$2695 ( \3072 , \3067 , \3071 );
xor \U$2696 ( \3073 , \3072 , \2520 );
not \U$2697 ( \3074 , \2530 );
xor \U$2698 ( \3075 , \2539 , \2550 );
not \U$2699 ( \3076 , \3075 );
or \U$2700 ( \3077 , \3074 , \3076 );
or \U$2701 ( \3078 , \3075 , \2530 );
nand \U$2702 ( \3079 , \3077 , \3078 );
xor \U$2703 ( \3080 , \3073 , \3079 );
or \U$2704 ( \3081 , \3057 , \3037 );
not \U$2705 ( \3082 , \3037 );
not \U$2706 ( \3083 , \3057 );
or \U$2707 ( \3084 , \3082 , \3083 );
nand \U$2708 ( \3085 , \3084 , \3045 );
nand \U$2709 ( \3086 , \3081 , \3085 );
or \U$2710 ( \3087 , \2957 , \2789 );
not \U$2711 ( \3088 , \2789 );
not \U$2712 ( \3089 , \3088 );
not \U$2713 ( \3090 , \3089 );
not \U$2714 ( \3091 , \2957 );
or \U$2715 ( \3092 , \3090 , \3091 );
nand \U$2716 ( \3093 , \3092 , \2945 );
nand \U$2717 ( \3094 , \3087 , \3093 );
xor \U$2718 ( \3095 , \3086 , \3094 );
or \U$2719 ( \3096 , \2988 , \2968 );
not \U$2720 ( \3097 , \2968 );
not \U$2721 ( \3098 , \2988 );
or \U$2722 ( \3099 , \3097 , \3098 );
nand \U$2723 ( \3100 , \3099 , \2976 );
nand \U$2724 ( \3101 , \3096 , \3100 );
xor \U$2725 ( \3102 , \3095 , \3101 );
xor \U$2726 ( \3103 , \3080 , \3102 );
not \U$2727 ( \3104 , \2623 );
xor \U$2728 ( \3105 , \2631 , \2641 );
not \U$2729 ( \3106 , \3105 );
or \U$2730 ( \3107 , \3104 , \3106 );
or \U$2731 ( \3108 , \3105 , \2623 );
nand \U$2732 ( \3109 , \3107 , \3108 );
not \U$2733 ( \3110 , \2588 );
xor \U$2734 ( \3111 , \2613 , \2596 );
not \U$2735 ( \3112 , \3111 );
or \U$2736 ( \3113 , \3110 , \3112 );
or \U$2737 ( \3114 , \3111 , \2588 );
nand \U$2738 ( \3115 , \3113 , \3114 );
xor \U$2739 ( \3116 , \3109 , \3115 );
xor \U$2740 ( \3117 , \2562 , \2570 );
xor \U$2741 ( \3118 , \3117 , \2578 );
xor \U$2742 ( \3119 , \3116 , \3118 );
xor \U$2743 ( \3120 , \3103 , \3119 );
xor \U$2744 ( \3121 , \3066 , \3120 );
not \U$2745 ( \3122 , \3121 );
not \U$2746 ( \3123 , \2706 );
not \U$2747 ( \3124 , \2719 );
or \U$2748 ( \3125 , \3123 , \3124 );
or \U$2749 ( \3126 , \2706 , \2719 );
nand \U$2750 ( \3127 , \3125 , \3126 );
not \U$2751 ( \3128 , \3127 );
not \U$2752 ( \3129 , \2707 );
and \U$2753 ( \3130 , \3128 , \3129 );
and \U$2754 ( \3131 , \3127 , \2707 );
nor \U$2755 ( \3132 , \3130 , \3131 );
and \U$2756 ( \3133 , \672 , RIae75128_1);
and \U$2757 ( \3134 , RIae75308_5, \670 );
nor \U$2758 ( \3135 , \3133 , \3134 );
and \U$2759 ( \3136 , \3135 , \587 );
not \U$2760 ( \3137 , \3135 );
and \U$2761 ( \3138 , \3137 , \588 );
nor \U$2762 ( \3139 , \3136 , \3138 );
and \U$2763 ( \3140 , \514 , RIae754e8_9);
and \U$2764 ( \3141 , RIae757b8_15, \512 );
nor \U$2765 ( \3142 , \3140 , \3141 );
not \U$2766 ( \3143 , \3142 );
not \U$2767 ( \3144 , \469 );
and \U$2768 ( \3145 , \3143 , \3144 );
and \U$2769 ( \3146 , \3142 , \471 );
nor \U$2770 ( \3147 , \3145 , \3146 );
xor \U$2771 ( \3148 , \3139 , \3147 );
and \U$2772 ( \3149 , \558 , RIae756c8_13);
and \U$2773 ( \3150 , RIae75218_3, \556 );
nor \U$2774 ( \3151 , \3149 , \3150 );
and \U$2775 ( \3152 , \3151 , \562 );
not \U$2776 ( \3153 , \3151 );
and \U$2777 ( \3154 , \3153 , \504 );
nor \U$2778 ( \3155 , \3152 , \3154 );
and \U$2779 ( \3156 , \3148 , \3155 );
and \U$2780 ( \3157 , \3139 , \3147 );
or \U$2781 ( \3158 , \3156 , \3157 );
or \U$2782 ( \3159 , \3132 , \3158 );
not \U$2783 ( \3160 , \3158 );
not \U$2784 ( \3161 , \3132 );
or \U$2785 ( \3162 , \3160 , \3161 );
and \U$2786 ( \3163 , \384 , RIae75e48_29);
and \U$2787 ( \3164 , RIae75c68_25, \382 );
nor \U$2788 ( \3165 , \3163 , \3164 );
not \U$2789 ( \3166 , \3165 );
not \U$2790 ( \3167 , \392 );
and \U$2791 ( \3168 , \3166 , \3167 );
and \U$2792 ( \3169 , \3165 , \392 );
nor \U$2793 ( \3170 , \3168 , \3169 );
nand \U$2794 ( \3171 , RIae75f38_31, RIae78b48_125);
or \U$2795 ( \3172 , \3170 , \3171 );
not \U$2796 ( \3173 , \3171 );
not \U$2797 ( \3174 , \3170 );
or \U$2798 ( \3175 , \3173 , \3174 );
not \U$2799 ( \3176 , \400 );
and \U$2800 ( \3177 , \436 , RIae75d58_27);
and \U$2801 ( \3178 , RIae755d8_11, \434 );
nor \U$2802 ( \3179 , \3177 , \3178 );
not \U$2803 ( \3180 , \3179 );
or \U$2804 ( \3181 , \3176 , \3180 );
or \U$2805 ( \3182 , \3179 , \402 );
nand \U$2806 ( \3183 , \3181 , \3182 );
nand \U$2807 ( \3184 , \3175 , \3183 );
nand \U$2808 ( \3185 , \3172 , \3184 );
nand \U$2809 ( \3186 , \3162 , \3185 );
nand \U$2810 ( \3187 , \3159 , \3186 );
and \U$2811 ( \3188 , \2607 , RIae76898_51);
and \U$2812 ( \3189 , RIae76b68_57, \2605 );
nor \U$2813 ( \3190 , \3188 , \3189 );
and \U$2814 ( \3191 , \3190 , \2397 );
not \U$2815 ( \3192 , \3190 );
and \U$2816 ( \3193 , \3192 , \2611 );
nor \U$2817 ( \3194 , \3191 , \3193 );
not \U$2818 ( \3195 , \3194 );
and \U$2819 ( \3196 , \2783 , RIae78a58_123);
and \U$2820 ( \3197 , RIae78cb0_128, \2781 );
nor \U$2821 ( \3198 , \3196 , \3197 );
not \U$2822 ( \3199 , \3198 );
not \U$2823 ( \3200 , \2789 );
and \U$2824 ( \3201 , \3199 , \3200 );
and \U$2825 ( \3202 , \3198 , \2789 );
nor \U$2826 ( \3203 , \3201 , \3202 );
not \U$2827 ( \3204 , \3203 );
and \U$2828 ( \3205 , \3195 , \3204 );
and \U$2829 ( \3206 , \3203 , \3194 );
and \U$2830 ( \3207 , RIae798e0_154, RIae79868_153);
not \U$2831 ( \3208 , RIae797f0_152);
and \U$2832 ( \3209 , RIae79868_153, \3208 );
not \U$2833 ( \3210 , RIae79868_153);
and \U$2834 ( \3211 , \3210 , RIae797f0_152);
or \U$2835 ( \3212 , \3209 , \3211 );
nor \U$2836 ( \3213 , RIae798e0_154, RIae79868_153);
nor \U$2837 ( \3214 , \3207 , \3212 , \3213 );
nand \U$2838 ( \3215 , RIae78da0_130, \3214 );
not \U$2839 ( \3216 , \3215 );
not \U$2840 ( \3217 , \2774 );
not \U$2841 ( \3218 , \3217 );
not \U$2842 ( \3219 , \3218 );
and \U$2843 ( \3220 , \3216 , \3219 );
and \U$2844 ( \3221 , \3215 , \2774 );
nor \U$2845 ( \3222 , \3220 , \3221 );
nor \U$2846 ( \3223 , \3206 , \3222 );
nor \U$2847 ( \3224 , \3205 , \3223 );
and \U$2848 ( \3225 , \1593 , RIae76028_33);
and \U$2849 ( \3226 , RIae762f8_39, \1591 );
nor \U$2850 ( \3227 , \3225 , \3226 );
and \U$2851 ( \3228 , \3227 , \1488 );
not \U$2852 ( \3229 , \3227 );
and \U$2853 ( \3230 , \3229 , \1498 );
nor \U$2854 ( \3231 , \3228 , \3230 );
not \U$2855 ( \3232 , \3231 );
and \U$2856 ( \3233 , \1939 , RIae76208_37);
and \U$2857 ( \3234 , RIae76a78_55, \1937 );
nor \U$2858 ( \3235 , \3233 , \3234 );
and \U$2859 ( \3236 , \3235 , \1734 );
not \U$2860 ( \3237 , \3235 );
and \U$2861 ( \3238 , \3237 , \1735 );
nor \U$2862 ( \3239 , \3236 , \3238 );
not \U$2863 ( \3240 , \3239 );
and \U$2864 ( \3241 , \3232 , \3240 );
and \U$2865 ( \3242 , \3239 , \3231 );
and \U$2866 ( \3243 , \2224 , RIae76988_53);
and \U$2867 ( \3244 , RIae767a8_49, \2222 );
nor \U$2868 ( \3245 , \3243 , \3244 );
and \U$2869 ( \3246 , \3245 , \2060 );
not \U$2870 ( \3247 , \3245 );
and \U$2871 ( \3248 , \3247 , \2061 );
nor \U$2872 ( \3249 , \3246 , \3248 );
nor \U$2873 ( \3250 , \3242 , \3249 );
nor \U$2874 ( \3251 , \3241 , \3250 );
xor \U$2875 ( \3252 , \3224 , \3251 );
and \U$2876 ( \3253 , \1376 , RIae765c8_45);
and \U$2877 ( \3254 , RIae76118_35, \1374 );
nor \U$2878 ( \3255 , \3253 , \3254 );
and \U$2879 ( \3256 , \3255 , \1261 );
not \U$2880 ( \3257 , \3255 );
and \U$2881 ( \3258 , \3257 , \1380 );
nor \U$2882 ( \3259 , \3256 , \3258 );
and \U$2883 ( \3260 , \883 , RIae753f8_7);
and \U$2884 ( \3261 , RIae763e8_41, \881 );
nor \U$2885 ( \3262 , \3260 , \3261 );
not \U$2886 ( \3263 , \3262 );
not \U$2887 ( \3264 , \789 );
and \U$2888 ( \3265 , \3263 , \3264 );
and \U$2889 ( \3266 , \3262 , \789 );
nor \U$2890 ( \3267 , \3265 , \3266 );
xor \U$2891 ( \3268 , \3259 , \3267 );
and \U$2892 ( \3269 , \1138 , RIae764d8_43);
and \U$2893 ( \3270 , RIae766b8_47, \1136 );
nor \U$2894 ( \3271 , \3269 , \3270 );
and \U$2895 ( \3272 , \3271 , \1142 );
not \U$2896 ( \3273 , \3271 );
and \U$2897 ( \3274 , \3273 , \1012 );
nor \U$2898 ( \3275 , \3272 , \3274 );
and \U$2899 ( \3276 , \3268 , \3275 );
and \U$2900 ( \3277 , \3259 , \3267 );
or \U$2901 ( \3278 , \3276 , \3277 );
and \U$2902 ( \3279 , \3252 , \3278 );
and \U$2903 ( \3280 , \3224 , \3251 );
nor \U$2904 ( \3281 , \3279 , \3280 );
xor \U$2905 ( \3282 , \3187 , \3281 );
not \U$2906 ( \3283 , \2749 );
not \U$2907 ( \3284 , \2760 );
or \U$2908 ( \3285 , \3283 , \3284 );
or \U$2909 ( \3286 , \2749 , \2760 );
nand \U$2910 ( \3287 , \3285 , \3286 );
not \U$2911 ( \3288 , \3287 );
not \U$2912 ( \3289 , \2742 );
and \U$2913 ( \3290 , \3288 , \3289 );
and \U$2914 ( \3291 , \3287 , \2742 );
nor \U$2915 ( \3292 , \3290 , \3291 );
xor \U$2916 ( \3293 , \2803 , \2810 );
xor \U$2917 ( \3294 , \3293 , \2818 );
xor \U$2918 ( \3295 , \3292 , \3294 );
xor \U$2919 ( \3296 , \2829 , \2837 );
xor \U$2920 ( \3297 , \3296 , \2845 );
and \U$2921 ( \3298 , \3295 , \3297 );
and \U$2922 ( \3299 , \3292 , \3294 );
nor \U$2923 ( \3300 , \3298 , \3299 );
and \U$2924 ( \3301 , \3282 , \3300 );
and \U$2925 ( \3302 , \3187 , \3281 );
or \U$2926 ( \3303 , \3301 , \3302 );
and \U$2927 ( \3304 , \2224 , RIae76898_51);
and \U$2928 ( \3305 , RIae76b68_57, \2222 );
nor \U$2929 ( \3306 , \3304 , \3305 );
and \U$2930 ( \3307 , \3306 , \2060 );
not \U$2931 ( \3308 , \3306 );
and \U$2932 ( \3309 , \3308 , \2061 );
nor \U$2933 ( \3310 , \3307 , \3309 );
not \U$2934 ( \3311 , \3310 );
nand \U$2935 ( \3312 , RIae78da0_130, \2783 );
not \U$2936 ( \3313 , \3312 );
not \U$2937 ( \3314 , \2789 );
and \U$2938 ( \3315 , \3313 , \3314 );
and \U$2939 ( \3316 , \3312 , \3089 );
nor \U$2940 ( \3317 , \3315 , \3316 );
and \U$2941 ( \3318 , \2607 , RIae78a58_123);
and \U$2942 ( \3319 , RIae78cb0_128, \2605 );
nor \U$2943 ( \3320 , \3318 , \3319 );
and \U$2944 ( \3321 , \3320 , \2397 );
not \U$2945 ( \3322 , \3320 );
and \U$2946 ( \3323 , \3322 , \2611 );
nor \U$2947 ( \3324 , \3321 , \3323 );
xor \U$2948 ( \3325 , \3317 , \3324 );
not \U$2949 ( \3326 , \3325 );
or \U$2950 ( \3327 , \3311 , \3326 );
or \U$2951 ( \3328 , \3325 , \3310 );
nand \U$2952 ( \3329 , \3327 , \3328 );
xor \U$2953 ( \3330 , \2721 , \2733 );
xor \U$2954 ( \3331 , \3330 , \2762 );
and \U$2955 ( \3332 , \3329 , \3331 );
xor \U$2956 ( \3333 , \2883 , \2891 );
xor \U$2957 ( \3334 , \3333 , \2900 );
xor \U$2958 ( \3335 , \2876 , \2929 );
xor \U$2959 ( \3336 , \3334 , \3335 );
xor \U$2960 ( \3337 , \2721 , \2733 );
xor \U$2961 ( \3338 , \3337 , \2762 );
and \U$2962 ( \3339 , \3336 , \3338 );
and \U$2963 ( \3340 , \3329 , \3336 );
or \U$2964 ( \3341 , \3332 , \3339 , \3340 );
xnor \U$2965 ( \3342 , \3303 , \3341 );
not \U$2966 ( \3343 , \3342 );
not \U$2967 ( \3344 , \388 );
and \U$2968 ( \3345 , \384 , RIae755d8_11);
and \U$2969 ( \3346 , RIae754e8_9, \382 );
nor \U$2970 ( \3347 , \3345 , \3346 );
not \U$2971 ( \3348 , \3347 );
or \U$2972 ( \3349 , \3344 , \3348 );
or \U$2973 ( \3350 , \3347 , \388 );
nand \U$2974 ( \3351 , \3349 , \3350 );
xor \U$2975 ( \3352 , \2732 , \3351 );
xor \U$2976 ( \3353 , \2883 , \2891 );
and \U$2977 ( \3354 , \3353 , \2900 );
and \U$2978 ( \3355 , \2883 , \2891 );
or \U$2979 ( \3356 , \3354 , \3355 );
xor \U$2980 ( \3357 , \3352 , \3356 );
not \U$2981 ( \3358 , \3357 );
and \U$2982 ( \3359 , \3343 , \3358 );
and \U$2983 ( \3360 , \3342 , \3357 );
nor \U$2984 ( \3361 , \3359 , \3360 );
xor \U$2985 ( \3362 , \2772 , \2774 );
xor \U$2986 ( \3363 , \3362 , \2793 );
not \U$2987 ( \3364 , \3185 );
not \U$2988 ( \3365 , \3158 );
or \U$2989 ( \3366 , \3364 , \3365 );
or \U$2990 ( \3367 , \3158 , \3185 );
nand \U$2991 ( \3368 , \3366 , \3367 );
not \U$2992 ( \3369 , \3368 );
not \U$2993 ( \3370 , \3132 );
and \U$2994 ( \3371 , \3369 , \3370 );
and \U$2995 ( \3372 , \3368 , \3132 );
nor \U$2996 ( \3373 , \3371 , \3372 );
xor \U$2997 ( \3374 , \3363 , \3373 );
xor \U$2998 ( \3375 , \3292 , \3294 );
xor \U$2999 ( \3376 , \3375 , \3297 );
and \U$3000 ( \3377 , \3374 , \3376 );
and \U$3001 ( \3378 , \3363 , \3373 );
nor \U$3002 ( \3379 , \3377 , \3378 );
xor \U$3003 ( \3380 , \2796 , \2821 );
xor \U$3004 ( \3381 , \3380 , \2848 );
not \U$3005 ( \3382 , \3381 );
and \U$3006 ( \3383 , \3379 , \3382 );
not \U$3007 ( \3384 , \3379 );
not \U$3008 ( \3385 , \3382 );
and \U$3009 ( \3386 , \3384 , \3385 );
and \U$3010 ( \3387 , \2607 , RIae767a8_49);
and \U$3011 ( \3388 , RIae76898_51, \2605 );
nor \U$3012 ( \3389 , \3387 , \3388 );
and \U$3013 ( \3390 , \3389 , \2397 );
not \U$3014 ( \3391 , \3389 );
and \U$3015 ( \3392 , \3391 , \2611 );
nor \U$3016 ( \3393 , \3390 , \3392 );
and \U$3017 ( \3394 , \1939 , RIae762f8_39);
and \U$3018 ( \3395 , RIae76208_37, \1937 );
nor \U$3019 ( \3396 , \3394 , \3395 );
and \U$3020 ( \3397 , \3396 , \1734 );
not \U$3021 ( \3398 , \3396 );
and \U$3022 ( \3399 , \3398 , \1735 );
nor \U$3023 ( \3400 , \3397 , \3399 );
xor \U$3024 ( \3401 , \3393 , \3400 );
and \U$3025 ( \3402 , \2224 , RIae76a78_55);
and \U$3026 ( \3403 , RIae76988_53, \2222 );
nor \U$3027 ( \3404 , \3402 , \3403 );
and \U$3028 ( \3405 , \3404 , \2060 );
not \U$3029 ( \3406 , \3404 );
and \U$3030 ( \3407 , \3406 , \2061 );
nor \U$3031 ( \3408 , \3405 , \3407 );
and \U$3032 ( \3409 , \3401 , \3408 );
and \U$3033 ( \3410 , \3393 , \3400 );
or \U$3034 ( \3411 , \3409 , \3410 );
and \U$3035 ( \3412 , \2783 , RIae76b68_57);
and \U$3036 ( \3413 , RIae78a58_123, \2781 );
nor \U$3037 ( \3414 , \3412 , \3413 );
not \U$3038 ( \3415 , \3414 );
not \U$3039 ( \3416 , \2789 );
and \U$3040 ( \3417 , \3415 , \3416 );
and \U$3041 ( \3418 , \3414 , \2789 );
nor \U$3042 ( \3419 , \3417 , \3418 );
and \U$3043 ( \3420 , RIae79700_150, RIae79778_151);
nor \U$3044 ( \3421 , \3420 , \3208 );
buf \U$3045 ( \3422 , \3421 );
xor \U$3046 ( \3423 , \3419 , \3422 );
and \U$3047 ( \3424 , \3214 , RIae78cb0_128);
and \U$3048 ( \3425 , RIae78da0_130, \3212 );
nor \U$3049 ( \3426 , \3424 , \3425 );
not \U$3050 ( \3427 , \3426 );
not \U$3051 ( \3428 , \2774 );
and \U$3052 ( \3429 , \3427 , \3428 );
and \U$3053 ( \3430 , \3426 , \3218 );
nor \U$3054 ( \3431 , \3429 , \3430 );
and \U$3055 ( \3432 , \3423 , \3431 );
and \U$3056 ( \3433 , \3419 , \3422 );
or \U$3057 ( \3434 , \3432 , \3433 );
xor \U$3058 ( \3435 , \3411 , \3434 );
and \U$3059 ( \3436 , \1593 , RIae76118_35);
and \U$3060 ( \3437 , RIae76028_33, \1591 );
nor \U$3061 ( \3438 , \3436 , \3437 );
and \U$3062 ( \3439 , \3438 , \1488 );
not \U$3063 ( \3440 , \3438 );
and \U$3064 ( \3441 , \3440 , \1498 );
nor \U$3065 ( \3442 , \3439 , \3441 );
and \U$3066 ( \3443 , \1138 , RIae763e8_41);
and \U$3067 ( \3444 , RIae764d8_43, \1136 );
nor \U$3068 ( \3445 , \3443 , \3444 );
and \U$3069 ( \3446 , \3445 , \1142 );
not \U$3070 ( \3447 , \3445 );
and \U$3071 ( \3448 , \3447 , \1012 );
nor \U$3072 ( \3449 , \3446 , \3448 );
xor \U$3073 ( \3450 , \3442 , \3449 );
and \U$3074 ( \3451 , \1376 , RIae766b8_47);
and \U$3075 ( \3452 , RIae765c8_45, \1374 );
nor \U$3076 ( \3453 , \3451 , \3452 );
and \U$3077 ( \3454 , \3453 , \1261 );
not \U$3078 ( \3455 , \3453 );
and \U$3079 ( \3456 , \3455 , \1380 );
nor \U$3080 ( \3457 , \3454 , \3456 );
and \U$3081 ( \3458 , \3450 , \3457 );
and \U$3082 ( \3459 , \3442 , \3449 );
or \U$3083 ( \3460 , \3458 , \3459 );
and \U$3084 ( \3461 , \3435 , \3460 );
and \U$3085 ( \3462 , \3411 , \3434 );
or \U$3086 ( \3463 , \3461 , \3462 );
and \U$3087 ( \3464 , \384 , RIae75f38_31);
and \U$3088 ( \3465 , RIae75e48_29, \382 );
nor \U$3089 ( \3466 , \3464 , \3465 );
not \U$3090 ( \3467 , \3466 );
not \U$3091 ( \3468 , \388 );
and \U$3092 ( \3469 , \3467 , \3468 );
and \U$3093 ( \3470 , \3466 , \388 );
nor \U$3094 ( \3471 , \3469 , \3470 );
and \U$3095 ( \3472 , \436 , RIae75c68_25);
and \U$3096 ( \3473 , RIae75d58_27, \434 );
nor \U$3097 ( \3474 , \3472 , \3473 );
not \U$3098 ( \3475 , \3474 );
not \U$3099 ( \3476 , \400 );
and \U$3100 ( \3477 , \3475 , \3476 );
and \U$3101 ( \3478 , \3474 , \402 );
nor \U$3102 ( \3479 , \3477 , \3478 );
or \U$3103 ( \3480 , \3471 , \3479 );
not \U$3104 ( \3481 , \3479 );
not \U$3105 ( \3482 , \3471 );
or \U$3106 ( \3483 , \3481 , \3482 );
not \U$3107 ( \3484 , \471 );
and \U$3108 ( \3485 , \514 , RIae755d8_11);
and \U$3109 ( \3486 , RIae754e8_9, \512 );
nor \U$3110 ( \3487 , \3485 , \3486 );
not \U$3111 ( \3488 , \3487 );
or \U$3112 ( \3489 , \3484 , \3488 );
or \U$3113 ( \3490 , \3487 , \471 );
nand \U$3114 ( \3491 , \3489 , \3490 );
nand \U$3115 ( \3492 , \3483 , \3491 );
nand \U$3116 ( \3493 , \3480 , \3492 );
and \U$3117 ( \3494 , \558 , RIae757b8_15);
and \U$3118 ( \3495 , RIae756c8_13, \556 );
nor \U$3119 ( \3496 , \3494 , \3495 );
and \U$3120 ( \3497 , \3496 , \562 );
not \U$3121 ( \3498 , \3496 );
and \U$3122 ( \3499 , \3498 , \504 );
nor \U$3123 ( \3500 , \3497 , \3499 );
and \U$3124 ( \3501 , \672 , RIae75218_3);
and \U$3125 ( \3502 , RIae75128_1, \670 );
nor \U$3126 ( \3503 , \3501 , \3502 );
and \U$3127 ( \3504 , \3503 , \587 );
not \U$3128 ( \3505 , \3503 );
and \U$3129 ( \3506 , \3505 , \588 );
nor \U$3130 ( \3507 , \3504 , \3506 );
or \U$3131 ( \3508 , \3500 , \3507 );
not \U$3132 ( \3509 , \3507 );
not \U$3133 ( \3510 , \3500 );
or \U$3134 ( \3511 , \3509 , \3510 );
not \U$3135 ( \3512 , \789 );
and \U$3136 ( \3513 , \883 , RIae75308_5);
and \U$3137 ( \3514 , RIae753f8_7, \881 );
nor \U$3138 ( \3515 , \3513 , \3514 );
not \U$3139 ( \3516 , \3515 );
or \U$3140 ( \3517 , \3512 , \3516 );
or \U$3141 ( \3518 , \3515 , \789 );
nand \U$3142 ( \3519 , \3517 , \3518 );
nand \U$3143 ( \3520 , \3511 , \3519 );
nand \U$3144 ( \3521 , \3508 , \3520 );
nor \U$3145 ( \3522 , \3493 , \3521 );
xor \U$3146 ( \3523 , \3463 , \3522 );
xor \U$3147 ( \3524 , \3139 , \3147 );
xor \U$3148 ( \3525 , \3524 , \3155 );
xor \U$3149 ( \3526 , \3259 , \3267 );
xor \U$3150 ( \3527 , \3526 , \3275 );
and \U$3151 ( \3528 , \3525 , \3527 );
not \U$3152 ( \3529 , \3170 );
not \U$3153 ( \3530 , \3183 );
or \U$3154 ( \3531 , \3529 , \3530 );
or \U$3155 ( \3532 , \3170 , \3183 );
nand \U$3156 ( \3533 , \3531 , \3532 );
not \U$3157 ( \3534 , \3533 );
not \U$3158 ( \3535 , \3171 );
and \U$3159 ( \3536 , \3534 , \3535 );
and \U$3160 ( \3537 , \3533 , \3171 );
nor \U$3161 ( \3538 , \3536 , \3537 );
xor \U$3162 ( \3539 , \3259 , \3267 );
xor \U$3163 ( \3540 , \3539 , \3275 );
and \U$3164 ( \3541 , \3538 , \3540 );
and \U$3165 ( \3542 , \3525 , \3538 );
or \U$3166 ( \3543 , \3528 , \3541 , \3542 );
and \U$3167 ( \3544 , \3523 , \3543 );
and \U$3168 ( \3545 , \3463 , \3522 );
or \U$3169 ( \3546 , \3544 , \3545 );
nor \U$3170 ( \3547 , \3386 , \3546 );
nor \U$3171 ( \3548 , \3383 , \3547 );
xor \U$3172 ( \3549 , \3361 , \3548 );
xor \U$3173 ( \3550 , \2859 , \2866 );
and \U$3174 ( \3551 , \3550 , \2875 );
and \U$3175 ( \3552 , \2859 , \2866 );
or \U$3176 ( \3553 , \3551 , \3552 );
not \U$3177 ( \3554 , \3553 );
not \U$3178 ( \3555 , \2909 );
not \U$3179 ( \3556 , \2924 );
and \U$3180 ( \3557 , \3555 , \3556 );
and \U$3181 ( \3558 , \2924 , \2909 );
nor \U$3182 ( \3559 , \3558 , \2917 );
nor \U$3183 ( \3560 , \3557 , \3559 );
not \U$3184 ( \3561 , \3560 );
or \U$3185 ( \3562 , \3554 , \3561 );
or \U$3186 ( \3563 , \3560 , \3553 );
nand \U$3187 ( \3564 , \3562 , \3563 );
not \U$3188 ( \3565 , \3564 );
not \U$3189 ( \3566 , \3310 );
not \U$3190 ( \3567 , \3324 );
and \U$3191 ( \3568 , \3566 , \3567 );
and \U$3192 ( \3569 , \3324 , \3310 );
nor \U$3193 ( \3570 , \3569 , \3317 );
nor \U$3194 ( \3571 , \3568 , \3570 );
not \U$3195 ( \3572 , \3571 );
and \U$3196 ( \3573 , \3565 , \3572 );
and \U$3197 ( \3574 , \3564 , \3571 );
nor \U$3198 ( \3575 , \3573 , \3574 );
not \U$3199 ( \3576 , \3575 );
xor \U$3200 ( \3577 , \2765 , \2851 );
xor \U$3201 ( \3578 , \3577 , \2934 );
not \U$3202 ( \3579 , \3578 );
or \U$3203 ( \3580 , \3576 , \3579 );
or \U$3204 ( \3581 , \3578 , \3575 );
nand \U$3205 ( \3582 , \3580 , \3581 );
not \U$3206 ( \3583 , \3582 );
not \U$3207 ( \3584 , \3062 );
xor \U$3208 ( \3585 , \2961 , \2992 );
not \U$3209 ( \3586 , \3585 );
and \U$3210 ( \3587 , \3584 , \3586 );
and \U$3211 ( \3588 , \3062 , \3585 );
nor \U$3212 ( \3589 , \3587 , \3588 );
not \U$3213 ( \3590 , \3589 );
and \U$3214 ( \3591 , \3583 , \3590 );
and \U$3215 ( \3592 , \3582 , \3589 );
nor \U$3216 ( \3593 , \3591 , \3592 );
and \U$3217 ( \3594 , \3549 , \3593 );
and \U$3218 ( \3595 , \3361 , \3548 );
or \U$3219 ( \3596 , \3594 , \3595 );
not \U$3220 ( \3597 , \3596 );
not \U$3221 ( \3598 , \3357 );
not \U$3222 ( \3599 , \3303 );
or \U$3223 ( \3600 , \3598 , \3599 );
or \U$3224 ( \3601 , \3303 , \3357 );
nand \U$3225 ( \3602 , \3601 , \3341 );
nand \U$3226 ( \3603 , \3600 , \3602 );
xor \U$3227 ( \3604 , \3027 , \3028 );
and \U$3228 ( \3605 , \3604 , \3061 );
and \U$3229 ( \3606 , \3027 , \3028 );
or \U$3230 ( \3607 , \3605 , \3606 );
not \U$3231 ( \3608 , \3607 );
xor \U$3232 ( \3609 , \2732 , \3351 );
and \U$3233 ( \3610 , \3609 , \3356 );
and \U$3234 ( \3611 , \2732 , \3351 );
or \U$3235 ( \3612 , \3610 , \3611 );
or \U$3236 ( \3613 , \3571 , \3560 );
not \U$3237 ( \3614 , \3571 );
not \U$3238 ( \3615 , \3560 );
or \U$3239 ( \3616 , \3614 , \3615 );
nand \U$3240 ( \3617 , \3616 , \3553 );
nand \U$3241 ( \3618 , \3613 , \3617 );
xor \U$3242 ( \3619 , \3612 , \3618 );
not \U$3243 ( \3620 , \3619 );
or \U$3244 ( \3621 , \3608 , \3620 );
or \U$3245 ( \3622 , \3619 , \3607 );
nand \U$3246 ( \3623 , \3621 , \3622 );
xor \U$3247 ( \3624 , \3603 , \3623 );
or \U$3248 ( \3625 , \3589 , \3575 );
not \U$3249 ( \3626 , \3575 );
not \U$3250 ( \3627 , \3589 );
or \U$3251 ( \3628 , \3626 , \3627 );
nand \U$3252 ( \3629 , \3628 , \3578 );
nand \U$3253 ( \3630 , \3625 , \3629 );
xor \U$3254 ( \3631 , \3624 , \3630 );
not \U$3255 ( \3632 , \3631 );
and \U$3256 ( \3633 , \3597 , \3632 );
and \U$3257 ( \3634 , \3596 , \3631 );
nor \U$3258 ( \3635 , \3633 , \3634 );
not \U$3259 ( \3636 , \3635 );
or \U$3260 ( \3637 , \3122 , \3636 );
or \U$3261 ( \3638 , \3635 , \3121 );
nand \U$3262 ( \3639 , \3637 , \3638 );
not \U$3263 ( \3640 , \3639 );
xor \U$3264 ( \3641 , \3361 , \3548 );
xor \U$3265 ( \3642 , \3641 , \3593 );
not \U$3266 ( \3643 , \3642 );
xor \U$3267 ( \3644 , \3187 , \3281 );
xor \U$3268 ( \3645 , \3644 , \3300 );
not \U$3269 ( \3646 , \3381 );
not \U$3270 ( \3647 , \3546 );
not \U$3271 ( \3648 , \3379 );
or \U$3272 ( \3649 , \3647 , \3648 );
or \U$3273 ( \3650 , \3379 , \3546 );
nand \U$3274 ( \3651 , \3649 , \3650 );
not \U$3275 ( \3652 , \3651 );
or \U$3276 ( \3653 , \3646 , \3652 );
or \U$3277 ( \3654 , \3651 , \3381 );
nand \U$3278 ( \3655 , \3653 , \3654 );
and \U$3279 ( \3656 , \3645 , \3655 );
and \U$3280 ( \3657 , \3643 , \3656 );
not \U$3281 ( \3658 , \3643 );
not \U$3282 ( \3659 , \3656 );
and \U$3283 ( \3660 , \3658 , \3659 );
xor \U$3284 ( \3661 , \3224 , \3251 );
xor \U$3285 ( \3662 , \3661 , \3278 );
xor \U$3286 ( \3663 , \3463 , \3522 );
xor \U$3287 ( \3664 , \3663 , \3543 );
xor \U$3288 ( \3665 , \3662 , \3664 );
xor \U$3289 ( \3666 , \3363 , \3373 );
xor \U$3290 ( \3667 , \3666 , \3376 );
and \U$3291 ( \3668 , \3665 , \3667 );
and \U$3292 ( \3669 , \3662 , \3664 );
nor \U$3293 ( \3670 , \3668 , \3669 );
xor \U$3294 ( \3671 , \2721 , \2733 );
xor \U$3295 ( \3672 , \3671 , \2762 );
xor \U$3296 ( \3673 , \3329 , \3336 );
xor \U$3297 ( \3674 , \3672 , \3673 );
and \U$3298 ( \3675 , \3670 , \3674 );
not \U$3299 ( \3676 , \3670 );
not \U$3300 ( \3677 , \3674 );
and \U$3301 ( \3678 , \3676 , \3677 );
and \U$3302 ( \3679 , \2224 , RIae76208_37);
and \U$3303 ( \3680 , RIae76a78_55, \2222 );
nor \U$3304 ( \3681 , \3679 , \3680 );
and \U$3305 ( \3682 , \3681 , \2060 );
not \U$3306 ( \3683 , \3681 );
and \U$3307 ( \3684 , \3683 , \2061 );
nor \U$3308 ( \3685 , \3682 , \3684 );
and \U$3309 ( \3686 , \2607 , RIae76988_53);
and \U$3310 ( \3687 , RIae767a8_49, \2605 );
nor \U$3311 ( \3688 , \3686 , \3687 );
and \U$3312 ( \3689 , \3688 , \2397 );
not \U$3313 ( \3690 , \3688 );
and \U$3314 ( \3691 , \3690 , \2611 );
nor \U$3315 ( \3692 , \3689 , \3691 );
xor \U$3316 ( \3693 , \3685 , \3692 );
and \U$3317 ( \3694 , \1939 , RIae76028_33);
and \U$3318 ( \3695 , RIae762f8_39, \1937 );
nor \U$3319 ( \3696 , \3694 , \3695 );
and \U$3320 ( \3697 , \3696 , \1734 );
not \U$3321 ( \3698 , \3696 );
and \U$3322 ( \3699 , \3698 , \1735 );
nor \U$3323 ( \3700 , \3697 , \3699 );
and \U$3324 ( \3701 , \3693 , \3700 );
and \U$3325 ( \3702 , \3685 , \3692 );
nor \U$3326 ( \3703 , \3701 , \3702 );
and \U$3327 ( \3704 , \2783 , RIae76898_51);
and \U$3328 ( \3705 , RIae76b68_57, \2781 );
nor \U$3329 ( \3706 , \3704 , \3705 );
not \U$3330 ( \3707 , \3706 );
not \U$3331 ( \3708 , \3089 );
and \U$3332 ( \3709 , \3707 , \3708 );
and \U$3333 ( \3710 , \3706 , \3089 );
nor \U$3334 ( \3711 , \3709 , \3710 );
and \U$3335 ( \3712 , \3214 , RIae78a58_123);
and \U$3336 ( \3713 , RIae78cb0_128, \3212 );
nor \U$3337 ( \3714 , \3712 , \3713 );
not \U$3338 ( \3715 , \3714 );
not \U$3339 ( \3716 , \3218 );
and \U$3340 ( \3717 , \3715 , \3716 );
and \U$3341 ( \3718 , \3714 , \3218 );
nor \U$3342 ( \3719 , \3717 , \3718 );
or \U$3343 ( \3720 , \3711 , \3719 );
not \U$3344 ( \3721 , \3719 );
not \U$3345 ( \3722 , \3711 );
or \U$3346 ( \3723 , \3721 , \3722 );
and \U$3347 ( \3724 , RIae797f0_152, RIae79700_150);
not \U$3348 ( \3725 , RIae79778_151);
and \U$3349 ( \3726 , \3725 , RIae79700_150);
nor \U$3350 ( \3727 , \3725 , RIae79700_150);
or \U$3351 ( \3728 , \3726 , \3727 );
nor \U$3352 ( \3729 , RIae797f0_152, RIae79700_150);
nor \U$3353 ( \3730 , \3724 , \3728 , \3729 );
nand \U$3354 ( \3731 , RIae78da0_130, \3730 );
not \U$3355 ( \3732 , \3421 );
and \U$3356 ( \3733 , \3731 , \3732 );
not \U$3357 ( \3734 , \3731 );
and \U$3358 ( \3735 , \3734 , \3422 );
nor \U$3359 ( \3736 , \3733 , \3735 );
nand \U$3360 ( \3737 , \3723 , \3736 );
nand \U$3361 ( \3738 , \3720 , \3737 );
xor \U$3362 ( \3739 , \3703 , \3738 );
and \U$3363 ( \3740 , \1138 , RIae753f8_7);
and \U$3364 ( \3741 , RIae763e8_41, \1136 );
nor \U$3365 ( \3742 , \3740 , \3741 );
and \U$3366 ( \3743 , \3742 , \1142 );
not \U$3367 ( \3744 , \3742 );
and \U$3368 ( \3745 , \3744 , \1012 );
nor \U$3369 ( \3746 , \3743 , \3745 );
and \U$3370 ( \3747 , \1376 , RIae764d8_43);
and \U$3371 ( \3748 , RIae766b8_47, \1374 );
nor \U$3372 ( \3749 , \3747 , \3748 );
and \U$3373 ( \3750 , \3749 , \1261 );
not \U$3374 ( \3751 , \3749 );
and \U$3375 ( \3752 , \3751 , \1380 );
nor \U$3376 ( \3753 , \3750 , \3752 );
or \U$3377 ( \3754 , \3746 , \3753 );
not \U$3378 ( \3755 , \3753 );
not \U$3379 ( \3756 , \3746 );
or \U$3380 ( \3757 , \3755 , \3756 );
and \U$3381 ( \3758 , \1593 , RIae765c8_45);
and \U$3382 ( \3759 , RIae76118_35, \1591 );
nor \U$3383 ( \3760 , \3758 , \3759 );
and \U$3384 ( \3761 , \3760 , \1498 );
not \U$3385 ( \3762 , \3760 );
and \U$3386 ( \3763 , \3762 , \1488 );
nor \U$3387 ( \3764 , \3761 , \3763 );
nand \U$3388 ( \3765 , \3757 , \3764 );
nand \U$3389 ( \3766 , \3754 , \3765 );
and \U$3390 ( \3767 , \3739 , \3766 );
and \U$3391 ( \3768 , \3703 , \3738 );
or \U$3392 ( \3769 , \3767 , \3768 );
and \U$3393 ( \3770 , \672 , RIae756c8_13);
and \U$3394 ( \3771 , RIae75218_3, \670 );
nor \U$3395 ( \3772 , \3770 , \3771 );
and \U$3396 ( \3773 , \3772 , \588 );
not \U$3397 ( \3774 , \3772 );
and \U$3398 ( \3775 , \3774 , \587 );
nor \U$3399 ( \3776 , \3773 , \3775 );
and \U$3400 ( \3777 , \558 , RIae754e8_9);
and \U$3401 ( \3778 , RIae757b8_15, \556 );
nor \U$3402 ( \3779 , \3777 , \3778 );
and \U$3403 ( \3780 , \3779 , \504 );
not \U$3404 ( \3781 , \3779 );
and \U$3405 ( \3782 , \3781 , \562 );
nor \U$3406 ( \3783 , \3780 , \3782 );
xor \U$3407 ( \3784 , \3776 , \3783 );
not \U$3408 ( \3785 , \787 );
and \U$3409 ( \3786 , \883 , RIae75128_1);
and \U$3410 ( \3787 , RIae75308_5, \881 );
nor \U$3411 ( \3788 , \3786 , \3787 );
not \U$3412 ( \3789 , \3788 );
or \U$3413 ( \3790 , \3785 , \3789 );
or \U$3414 ( \3791 , \3788 , \787 );
nand \U$3415 ( \3792 , \3790 , \3791 );
and \U$3416 ( \3793 , \3784 , \3792 );
and \U$3417 ( \3794 , \3776 , \3783 );
or \U$3418 ( \3795 , \3793 , \3794 );
nand \U$3419 ( \3796 , RIae75998_19, RIae78b48_125);
not \U$3420 ( \3797 , \3796 );
xor \U$3421 ( \3798 , \3795 , \3797 );
not \U$3422 ( \3799 , \392 );
and \U$3423 ( \3800 , \384 , RIae758a8_17);
and \U$3424 ( \3801 , RIae75f38_31, \382 );
nor \U$3425 ( \3802 , \3800 , \3801 );
not \U$3426 ( \3803 , \3802 );
or \U$3427 ( \3804 , \3799 , \3803 );
or \U$3428 ( \3805 , \3802 , \388 );
nand \U$3429 ( \3806 , \3804 , \3805 );
not \U$3430 ( \3807 , \402 );
and \U$3431 ( \3808 , \436 , RIae75e48_29);
and \U$3432 ( \3809 , RIae75c68_25, \434 );
nor \U$3433 ( \3810 , \3808 , \3809 );
not \U$3434 ( \3811 , \3810 );
or \U$3435 ( \3812 , \3807 , \3811 );
or \U$3436 ( \3813 , \3810 , \402 );
nand \U$3437 ( \3814 , \3812 , \3813 );
xor \U$3438 ( \3815 , \3806 , \3814 );
not \U$3439 ( \3816 , \471 );
and \U$3440 ( \3817 , \514 , RIae75d58_27);
and \U$3441 ( \3818 , RIae755d8_11, \512 );
nor \U$3442 ( \3819 , \3817 , \3818 );
not \U$3443 ( \3820 , \3819 );
or \U$3444 ( \3821 , \3816 , \3820 );
or \U$3445 ( \3822 , \3819 , \469 );
nand \U$3446 ( \3823 , \3821 , \3822 );
and \U$3447 ( \3824 , \3815 , \3823 );
and \U$3448 ( \3825 , \3806 , \3814 );
or \U$3449 ( \3826 , \3824 , \3825 );
and \U$3450 ( \3827 , \3798 , \3826 );
and \U$3451 ( \3828 , \3795 , \3797 );
or \U$3452 ( \3829 , \3827 , \3828 );
and \U$3453 ( \3830 , \3769 , \3829 );
not \U$3454 ( \3831 , \3769 );
not \U$3455 ( \3832 , \3829 );
and \U$3456 ( \3833 , \3831 , \3832 );
not \U$3457 ( \3834 , \3479 );
not \U$3458 ( \3835 , \3491 );
or \U$3459 ( \3836 , \3834 , \3835 );
or \U$3460 ( \3837 , \3479 , \3491 );
nand \U$3461 ( \3838 , \3836 , \3837 );
not \U$3462 ( \3839 , \3838 );
not \U$3463 ( \3840 , \3471 );
and \U$3464 ( \3841 , \3839 , \3840 );
and \U$3465 ( \3842 , \3838 , \3471 );
nor \U$3466 ( \3843 , \3841 , \3842 );
nand \U$3467 ( \3844 , RIae758a8_17, RIae78b48_125);
xor \U$3468 ( \3845 , \3843 , \3844 );
not \U$3469 ( \3846 , \3507 );
not \U$3470 ( \3847 , \3519 );
or \U$3471 ( \3848 , \3846 , \3847 );
or \U$3472 ( \3849 , \3507 , \3519 );
nand \U$3473 ( \3850 , \3848 , \3849 );
not \U$3474 ( \3851 , \3850 );
not \U$3475 ( \3852 , \3500 );
and \U$3476 ( \3853 , \3851 , \3852 );
and \U$3477 ( \3854 , \3850 , \3500 );
nor \U$3478 ( \3855 , \3853 , \3854 );
and \U$3479 ( \3856 , \3845 , \3855 );
and \U$3480 ( \3857 , \3843 , \3844 );
or \U$3481 ( \3858 , \3856 , \3857 );
nor \U$3482 ( \3859 , \3833 , \3858 );
nor \U$3483 ( \3860 , \3830 , \3859 );
not \U$3484 ( \3861 , \3194 );
xor \U$3485 ( \3862 , \3222 , \3203 );
not \U$3486 ( \3863 , \3862 );
or \U$3487 ( \3864 , \3861 , \3863 );
or \U$3488 ( \3865 , \3862 , \3194 );
nand \U$3489 ( \3866 , \3864 , \3865 );
not \U$3490 ( \3867 , \3231 );
xor \U$3491 ( \3868 , \3239 , \3249 );
not \U$3492 ( \3869 , \3868 );
or \U$3493 ( \3870 , \3867 , \3869 );
or \U$3494 ( \3871 , \3868 , \3231 );
nand \U$3495 ( \3872 , \3870 , \3871 );
and \U$3496 ( \3873 , \3866 , \3872 );
not \U$3497 ( \3874 , \3866 );
not \U$3498 ( \3875 , \3872 );
and \U$3499 ( \3876 , \3874 , \3875 );
xor \U$3500 ( \3877 , \3419 , \3422 );
xor \U$3501 ( \3878 , \3877 , \3431 );
xor \U$3502 ( \3879 , \3393 , \3400 );
xor \U$3503 ( \3880 , \3879 , \3408 );
and \U$3504 ( \3881 , \3878 , \3880 );
xor \U$3505 ( \3882 , \3442 , \3449 );
xor \U$3506 ( \3883 , \3882 , \3457 );
xor \U$3507 ( \3884 , \3393 , \3400 );
xor \U$3508 ( \3885 , \3884 , \3408 );
and \U$3509 ( \3886 , \3883 , \3885 );
and \U$3510 ( \3887 , \3878 , \3883 );
or \U$3511 ( \3888 , \3881 , \3886 , \3887 );
nor \U$3512 ( \3889 , \3876 , \3888 );
nor \U$3513 ( \3890 , \3873 , \3889 );
xor \U$3514 ( \3891 , \3860 , \3890 );
and \U$3515 ( \3892 , \3493 , \3521 );
nor \U$3516 ( \3893 , \3892 , \3522 );
xor \U$3517 ( \3894 , \3411 , \3434 );
xor \U$3518 ( \3895 , \3894 , \3460 );
and \U$3519 ( \3896 , \3893 , \3895 );
xor \U$3520 ( \3897 , \3259 , \3267 );
xor \U$3521 ( \3898 , \3897 , \3275 );
xor \U$3522 ( \3899 , \3525 , \3538 );
xor \U$3523 ( \3900 , \3898 , \3899 );
xor \U$3524 ( \3901 , \3411 , \3434 );
xor \U$3525 ( \3902 , \3901 , \3460 );
and \U$3526 ( \3903 , \3900 , \3902 );
and \U$3527 ( \3904 , \3893 , \3900 );
or \U$3528 ( \3905 , \3896 , \3903 , \3904 );
and \U$3529 ( \3906 , \3891 , \3905 );
and \U$3530 ( \3907 , \3860 , \3890 );
or \U$3531 ( \3908 , \3906 , \3907 );
nor \U$3532 ( \3909 , \3678 , \3908 );
nor \U$3533 ( \3910 , \3675 , \3909 );
nor \U$3534 ( \3911 , \3660 , \3910 );
nor \U$3535 ( \3912 , \3657 , \3911 );
not \U$3536 ( \3913 , \3912 );
and \U$3537 ( \3914 , \3640 , \3913 );
and \U$3538 ( \3915 , \3639 , \3912 );
nor \U$3539 ( \3916 , \3914 , \3915 );
not \U$3540 ( \3917 , \3674 );
not \U$3541 ( \3918 , \3670 );
not \U$3542 ( \3919 , \3908 );
and \U$3543 ( \3920 , \3918 , \3919 );
and \U$3544 ( \3921 , \3670 , \3908 );
nor \U$3545 ( \3922 , \3920 , \3921 );
not \U$3546 ( \3923 , \3922 );
or \U$3547 ( \3924 , \3917 , \3923 );
or \U$3548 ( \3925 , \3922 , \3674 );
nand \U$3549 ( \3926 , \3924 , \3925 );
xor \U$3550 ( \3927 , \3645 , \3655 );
and \U$3551 ( \3928 , \3926 , \3927 );
not \U$3552 ( \3929 , \3926 );
not \U$3553 ( \3930 , \3927 );
and \U$3554 ( \3931 , \3929 , \3930 );
not \U$3555 ( \3932 , \3866 );
not \U$3556 ( \3933 , \3888 );
or \U$3557 ( \3934 , \3932 , \3933 );
or \U$3558 ( \3935 , \3888 , \3866 );
nand \U$3559 ( \3936 , \3934 , \3935 );
xor \U$3560 ( \3937 , \3872 , \3936 );
not \U$3561 ( \3938 , \3858 );
xor \U$3562 ( \3939 , \3769 , \3829 );
not \U$3563 ( \3940 , \3939 );
or \U$3564 ( \3941 , \3938 , \3940 );
or \U$3565 ( \3942 , \3939 , \3858 );
nand \U$3566 ( \3943 , \3941 , \3942 );
and \U$3567 ( \3944 , \3937 , \3943 );
not \U$3568 ( \3945 , \3937 );
not \U$3569 ( \3946 , \3943 );
and \U$3570 ( \3947 , \3945 , \3946 );
xor \U$3571 ( \3948 , \3411 , \3434 );
xor \U$3572 ( \3949 , \3948 , \3460 );
xor \U$3573 ( \3950 , \3893 , \3900 );
xor \U$3574 ( \3951 , \3949 , \3950 );
nor \U$3575 ( \3952 , \3947 , \3951 );
nor \U$3576 ( \3953 , \3944 , \3952 );
and \U$3577 ( \3954 , \1376 , RIae763e8_41);
and \U$3578 ( \3955 , RIae764d8_43, \1374 );
nor \U$3579 ( \3956 , \3954 , \3955 );
and \U$3580 ( \3957 , \3956 , \1380 );
not \U$3581 ( \3958 , \3956 );
and \U$3582 ( \3959 , \3958 , \1261 );
nor \U$3583 ( \3960 , \3957 , \3959 );
and \U$3584 ( \3961 , \1593 , RIae766b8_47);
and \U$3585 ( \3962 , RIae765c8_45, \1591 );
nor \U$3586 ( \3963 , \3961 , \3962 );
and \U$3587 ( \3964 , \3963 , \1498 );
not \U$3588 ( \3965 , \3963 );
and \U$3589 ( \3966 , \3965 , \1488 );
nor \U$3590 ( \3967 , \3964 , \3966 );
xor \U$3591 ( \3968 , \3960 , \3967 );
and \U$3592 ( \3969 , \1939 , RIae76118_35);
and \U$3593 ( \3970 , RIae76028_33, \1937 );
nor \U$3594 ( \3971 , \3969 , \3970 );
and \U$3595 ( \3972 , \3971 , \1735 );
not \U$3596 ( \3973 , \3971 );
and \U$3597 ( \3974 , \3973 , \1734 );
nor \U$3598 ( \3975 , \3972 , \3974 );
and \U$3599 ( \3976 , \3968 , \3975 );
and \U$3600 ( \3977 , \3960 , \3967 );
or \U$3601 ( \3978 , \3976 , \3977 );
and \U$3602 ( \3979 , \3730 , RIae78cb0_128);
and \U$3603 ( \3980 , RIae78da0_130, \3728 );
nor \U$3604 ( \3981 , \3979 , \3980 );
and \U$3605 ( \3982 , \3981 , \3732 );
not \U$3606 ( \3983 , \3981 );
and \U$3607 ( \3984 , \3983 , \3422 );
nor \U$3608 ( \3985 , \3982 , \3984 );
not \U$3609 ( \3986 , RIae79c28_161);
not \U$3610 ( \3987 , RIae79bb0_160);
or \U$3611 ( \3988 , \3986 , \3987 );
nand \U$3612 ( \3989 , \3988 , RIae79778_151);
xor \U$3613 ( \3990 , \3985 , \3989 );
not \U$3614 ( \3991 , \3218 );
and \U$3615 ( \3992 , \3214 , RIae76b68_57);
and \U$3616 ( \3993 , RIae78a58_123, \3212 );
nor \U$3617 ( \3994 , \3992 , \3993 );
not \U$3618 ( \3995 , \3994 );
or \U$3619 ( \3996 , \3991 , \3995 );
or \U$3620 ( \3997 , \3994 , \2774 );
nand \U$3621 ( \3998 , \3996 , \3997 );
and \U$3622 ( \3999 , \3990 , \3998 );
and \U$3623 ( \4000 , \3985 , \3989 );
or \U$3624 ( \4001 , \3999 , \4000 );
xor \U$3625 ( \4002 , \3978 , \4001 );
not \U$3626 ( \4003 , \3089 );
and \U$3627 ( \4004 , \2783 , RIae767a8_49);
and \U$3628 ( \4005 , RIae76898_51, \2781 );
nor \U$3629 ( \4006 , \4004 , \4005 );
not \U$3630 ( \4007 , \4006 );
or \U$3631 ( \4008 , \4003 , \4007 );
or \U$3632 ( \4009 , \4006 , \3089 );
nand \U$3633 ( \4010 , \4008 , \4009 );
and \U$3634 ( \4011 , \2224 , RIae762f8_39);
and \U$3635 ( \4012 , RIae76208_37, \2222 );
nor \U$3636 ( \4013 , \4011 , \4012 );
and \U$3637 ( \4014 , \4013 , \2061 );
not \U$3638 ( \4015 , \4013 );
and \U$3639 ( \4016 , \4015 , \2060 );
nor \U$3640 ( \4017 , \4014 , \4016 );
xor \U$3641 ( \4018 , \4010 , \4017 );
and \U$3642 ( \4019 , \2607 , RIae76a78_55);
and \U$3643 ( \4020 , RIae76988_53, \2605 );
nor \U$3644 ( \4021 , \4019 , \4020 );
and \U$3645 ( \4022 , \4021 , \2611 );
not \U$3646 ( \4023 , \4021 );
and \U$3647 ( \4024 , \4023 , \2397 );
nor \U$3648 ( \4025 , \4022 , \4024 );
and \U$3649 ( \4026 , \4018 , \4025 );
and \U$3650 ( \4027 , \4010 , \4017 );
or \U$3651 ( \4028 , \4026 , \4027 );
and \U$3652 ( \4029 , \4002 , \4028 );
and \U$3653 ( \4030 , \3978 , \4001 );
or \U$3654 ( \4031 , \4029 , \4030 );
not \U$3655 ( \4032 , \402 );
and \U$3656 ( \4033 , \436 , RIae75f38_31);
and \U$3657 ( \4034 , RIae75e48_29, \434 );
nor \U$3658 ( \4035 , \4033 , \4034 );
not \U$3659 ( \4036 , \4035 );
or \U$3660 ( \4037 , \4032 , \4036 );
or \U$3661 ( \4038 , \4035 , \402 );
nand \U$3662 ( \4039 , \4037 , \4038 );
not \U$3663 ( \4040 , \471 );
and \U$3664 ( \4041 , \514 , RIae75c68_25);
and \U$3665 ( \4042 , RIae75d58_27, \512 );
nor \U$3666 ( \4043 , \4041 , \4042 );
not \U$3667 ( \4044 , \4043 );
or \U$3668 ( \4045 , \4040 , \4044 );
or \U$3669 ( \4046 , \4043 , \471 );
nand \U$3670 ( \4047 , \4045 , \4046 );
xor \U$3671 ( \4048 , \4039 , \4047 );
and \U$3672 ( \4049 , \558 , RIae755d8_11);
and \U$3673 ( \4050 , RIae754e8_9, \556 );
nor \U$3674 ( \4051 , \4049 , \4050 );
and \U$3675 ( \4052 , \4051 , \504 );
not \U$3676 ( \4053 , \4051 );
and \U$3677 ( \4054 , \4053 , \562 );
nor \U$3678 ( \4055 , \4052 , \4054 );
and \U$3679 ( \4056 , \4048 , \4055 );
and \U$3680 ( \4057 , \4039 , \4047 );
or \U$3681 ( \4058 , \4056 , \4057 );
not \U$3682 ( \4059 , RIae75a88_21);
nor \U$3683 ( \4060 , \4059 , \491 );
not \U$3684 ( \4061 , \388 );
and \U$3685 ( \4062 , \384 , RIae75998_19);
and \U$3686 ( \4063 , RIae758a8_17, \382 );
nor \U$3687 ( \4064 , \4062 , \4063 );
not \U$3688 ( \4065 , \4064 );
or \U$3689 ( \4066 , \4061 , \4065 );
or \U$3690 ( \4067 , \4064 , \392 );
nand \U$3691 ( \4068 , \4066 , \4067 );
and \U$3692 ( \4069 , \4060 , \4068 );
xor \U$3693 ( \4070 , \4058 , \4069 );
and \U$3694 ( \4071 , \1138 , RIae75308_5);
and \U$3695 ( \4072 , RIae753f8_7, \1136 );
nor \U$3696 ( \4073 , \4071 , \4072 );
and \U$3697 ( \4074 , \4073 , \1012 );
not \U$3698 ( \4075 , \4073 );
and \U$3699 ( \4076 , \4075 , \1142 );
nor \U$3700 ( \4077 , \4074 , \4076 );
and \U$3701 ( \4078 , \672 , RIae757b8_15);
and \U$3702 ( \4079 , RIae756c8_13, \670 );
nor \U$3703 ( \4080 , \4078 , \4079 );
and \U$3704 ( \4081 , \4080 , \588 );
not \U$3705 ( \4082 , \4080 );
and \U$3706 ( \4083 , \4082 , \587 );
nor \U$3707 ( \4084 , \4081 , \4083 );
xor \U$3708 ( \4085 , \4077 , \4084 );
not \U$3709 ( \4086 , \787 );
and \U$3710 ( \4087 , \883 , RIae75218_3);
and \U$3711 ( \4088 , RIae75128_1, \881 );
nor \U$3712 ( \4089 , \4087 , \4088 );
not \U$3713 ( \4090 , \4089 );
or \U$3714 ( \4091 , \4086 , \4090 );
or \U$3715 ( \4092 , \4089 , \787 );
nand \U$3716 ( \4093 , \4091 , \4092 );
and \U$3717 ( \4094 , \4085 , \4093 );
and \U$3718 ( \4095 , \4077 , \4084 );
or \U$3719 ( \4096 , \4094 , \4095 );
and \U$3720 ( \4097 , \4070 , \4096 );
and \U$3721 ( \4098 , \4058 , \4069 );
or \U$3722 ( \4099 , \4097 , \4098 );
xor \U$3723 ( \4100 , \4031 , \4099 );
xor \U$3724 ( \4101 , \3776 , \3783 );
xor \U$3725 ( \4102 , \4101 , \3792 );
xor \U$3726 ( \4103 , \4102 , \3796 );
xor \U$3727 ( \4104 , \3806 , \3814 );
xor \U$3728 ( \4105 , \4104 , \3823 );
and \U$3729 ( \4106 , \4103 , \4105 );
and \U$3730 ( \4107 , \4102 , \3796 );
or \U$3731 ( \4108 , \4106 , \4107 );
and \U$3732 ( \4109 , \4100 , \4108 );
and \U$3733 ( \4110 , \4031 , \4099 );
or \U$3734 ( \4111 , \4109 , \4110 );
xor \U$3735 ( \4112 , \3703 , \3738 );
xor \U$3736 ( \4113 , \4112 , \3766 );
xor \U$3737 ( \4114 , \3795 , \3797 );
xor \U$3738 ( \4115 , \4114 , \3826 );
and \U$3739 ( \4116 , \4113 , \4115 );
and \U$3740 ( \4117 , \4111 , \4116 );
not \U$3741 ( \4118 , \4111 );
not \U$3742 ( \4119 , \4116 );
and \U$3743 ( \4120 , \4118 , \4119 );
xor \U$3744 ( \4121 , \3843 , \3844 );
xor \U$3745 ( \4122 , \4121 , \3855 );
not \U$3746 ( \4123 , \4122 );
xor \U$3747 ( \4124 , \3393 , \3400 );
xor \U$3748 ( \4125 , \4124 , \3408 );
xor \U$3749 ( \4126 , \3878 , \3883 );
xor \U$3750 ( \4127 , \4125 , \4126 );
not \U$3751 ( \4128 , \4127 );
and \U$3752 ( \4129 , \4123 , \4128 );
and \U$3753 ( \4130 , \4127 , \4122 );
not \U$3754 ( \4131 , \3736 );
not \U$3755 ( \4132 , \3719 );
or \U$3756 ( \4133 , \4131 , \4132 );
or \U$3757 ( \4134 , \3719 , \3736 );
nand \U$3758 ( \4135 , \4133 , \4134 );
not \U$3759 ( \4136 , \4135 );
not \U$3760 ( \4137 , \3711 );
and \U$3761 ( \4138 , \4136 , \4137 );
and \U$3762 ( \4139 , \4135 , \3711 );
nor \U$3763 ( \4140 , \4138 , \4139 );
not \U$3764 ( \4141 , \4140 );
not \U$3765 ( \4142 , \3753 );
not \U$3766 ( \4143 , \3764 );
or \U$3767 ( \4144 , \4142 , \4143 );
or \U$3768 ( \4145 , \3753 , \3764 );
nand \U$3769 ( \4146 , \4144 , \4145 );
not \U$3770 ( \4147 , \4146 );
not \U$3771 ( \4148 , \3746 );
and \U$3772 ( \4149 , \4147 , \4148 );
and \U$3773 ( \4150 , \4146 , \3746 );
nor \U$3774 ( \4151 , \4149 , \4150 );
not \U$3775 ( \4152 , \4151 );
and \U$3776 ( \4153 , \4141 , \4152 );
and \U$3777 ( \4154 , \4140 , \4151 );
xor \U$3778 ( \4155 , \3685 , \3692 );
xor \U$3779 ( \4156 , \4155 , \3700 );
nor \U$3780 ( \4157 , \4154 , \4156 );
nor \U$3781 ( \4158 , \4153 , \4157 );
nor \U$3782 ( \4159 , \4130 , \4158 );
nor \U$3783 ( \4160 , \4129 , \4159 );
nor \U$3784 ( \4161 , \4120 , \4160 );
nor \U$3785 ( \4162 , \4117 , \4161 );
xor \U$3786 ( \4163 , \3953 , \4162 );
xor \U$3787 ( \4164 , \3662 , \3664 );
xor \U$3788 ( \4165 , \4164 , \3667 );
and \U$3789 ( \4166 , \4163 , \4165 );
and \U$3790 ( \4167 , \3953 , \4162 );
or \U$3791 ( \4168 , \4166 , \4167 );
nor \U$3792 ( \4169 , \3931 , \4168 );
nor \U$3793 ( \4170 , \3928 , \4169 );
not \U$3794 ( \4171 , \4170 );
not \U$3795 ( \4172 , \3642 );
not \U$3796 ( \4173 , \3656 );
not \U$3797 ( \4174 , \3910 );
or \U$3798 ( \4175 , \4173 , \4174 );
or \U$3799 ( \4176 , \3910 , \3656 );
nand \U$3800 ( \4177 , \4175 , \4176 );
not \U$3801 ( \4178 , \4177 );
or \U$3802 ( \4179 , \4172 , \4178 );
or \U$3803 ( \4180 , \4177 , \3642 );
nand \U$3804 ( \4181 , \4179 , \4180 );
nand \U$3805 ( \4182 , \4171 , \4181 );
or \U$3806 ( \4183 , \3916 , \4182 );
xnor \U$3807 ( \4184 , \4182 , \3916 );
not \U$3808 ( \4185 , \4170 );
not \U$3809 ( \4186 , \4181 );
or \U$3810 ( \4187 , \4185 , \4186 );
or \U$3811 ( \4188 , \4181 , \4170 );
nand \U$3812 ( \4189 , \4187 , \4188 );
not \U$3813 ( \4190 , \3927 );
not \U$3814 ( \4191 , \3926 );
not \U$3815 ( \4192 , \4168 );
and \U$3816 ( \4193 , \4191 , \4192 );
and \U$3817 ( \4194 , \4168 , \3926 );
nor \U$3818 ( \4195 , \4193 , \4194 );
not \U$3819 ( \4196 , \4195 );
or \U$3820 ( \4197 , \4190 , \4196 );
or \U$3821 ( \4198 , \4195 , \3927 );
nand \U$3822 ( \4199 , \4197 , \4198 );
not \U$3823 ( \4200 , \4199 );
not \U$3824 ( \4201 , \3951 );
xor \U$3825 ( \4202 , \3943 , \3937 );
not \U$3826 ( \4203 , \4202 );
or \U$3827 ( \4204 , \4201 , \4203 );
or \U$3828 ( \4205 , \4202 , \3951 );
nand \U$3829 ( \4206 , \4204 , \4205 );
and \U$3830 ( \4207 , \1376 , RIae753f8_7);
and \U$3831 ( \4208 , RIae763e8_41, \1374 );
nor \U$3832 ( \4209 , \4207 , \4208 );
and \U$3833 ( \4210 , \4209 , \1380 );
not \U$3834 ( \4211 , \4209 );
and \U$3835 ( \4212 , \4211 , \1261 );
nor \U$3836 ( \4213 , \4210 , \4212 );
and \U$3837 ( \4214 , \1593 , RIae764d8_43);
and \U$3838 ( \4215 , RIae766b8_47, \1591 );
nor \U$3839 ( \4216 , \4214 , \4215 );
and \U$3840 ( \4217 , \4216 , \1498 );
not \U$3841 ( \4218 , \4216 );
and \U$3842 ( \4219 , \4218 , \1488 );
nor \U$3843 ( \4220 , \4217 , \4219 );
xor \U$3844 ( \4221 , \4213 , \4220 );
and \U$3845 ( \4222 , \1939 , RIae765c8_45);
and \U$3846 ( \4223 , RIae76118_35, \1937 );
nor \U$3847 ( \4224 , \4222 , \4223 );
and \U$3848 ( \4225 , \4224 , \1735 );
not \U$3849 ( \4226 , \4224 );
and \U$3850 ( \4227 , \4226 , \1734 );
nor \U$3851 ( \4228 , \4225 , \4227 );
and \U$3852 ( \4229 , \4221 , \4228 );
and \U$3853 ( \4230 , \4213 , \4220 );
or \U$3854 ( \4231 , \4229 , \4230 );
not \U$3855 ( \4232 , \3218 );
and \U$3856 ( \4233 , \3214 , RIae76898_51);
and \U$3857 ( \4234 , RIae76b68_57, \3212 );
nor \U$3858 ( \4235 , \4233 , \4234 );
not \U$3859 ( \4236 , \4235 );
or \U$3860 ( \4237 , \4232 , \4236 );
or \U$3861 ( \4238 , \4235 , \3218 );
nand \U$3862 ( \4239 , \4237 , \4238 );
and \U$3863 ( \4240 , RIae79778_151, RIae79bb0_160);
not \U$3864 ( \4241 , RIae79bb0_160);
nor \U$3865 ( \4242 , \4241 , RIae79c28_161);
not \U$3866 ( \4243 , RIae79c28_161);
nor \U$3867 ( \4244 , \4243 , RIae79bb0_160);
or \U$3868 ( \4245 , \4242 , \4244 );
nor \U$3869 ( \4246 , RIae79778_151, RIae79bb0_160);
nor \U$3870 ( \4247 , \4240 , \4245 , \4246 );
nand \U$3871 ( \4248 , RIae78da0_130, \4247 );
and \U$3872 ( \4249 , \4248 , \3989 );
not \U$3873 ( \4250 , \4248 );
not \U$3874 ( \4251 , \3989 );
and \U$3875 ( \4252 , \4250 , \4251 );
nor \U$3876 ( \4253 , \4249 , \4252 );
xor \U$3877 ( \4254 , \4239 , \4253 );
and \U$3878 ( \4255 , \3730 , RIae78a58_123);
and \U$3879 ( \4256 , RIae78cb0_128, \3728 );
nor \U$3880 ( \4257 , \4255 , \4256 );
and \U$3881 ( \4258 , \4257 , \3732 );
not \U$3882 ( \4259 , \4257 );
and \U$3883 ( \4260 , \4259 , \3422 );
nor \U$3884 ( \4261 , \4258 , \4260 );
and \U$3885 ( \4262 , \4254 , \4261 );
and \U$3886 ( \4263 , \4239 , \4253 );
or \U$3887 ( \4264 , \4262 , \4263 );
xor \U$3888 ( \4265 , \4231 , \4264 );
and \U$3889 ( \4266 , \2224 , RIae76028_33);
and \U$3890 ( \4267 , RIae762f8_39, \2222 );
nor \U$3891 ( \4268 , \4266 , \4267 );
and \U$3892 ( \4269 , \4268 , \2061 );
not \U$3893 ( \4270 , \4268 );
and \U$3894 ( \4271 , \4270 , \2060 );
nor \U$3895 ( \4272 , \4269 , \4271 );
and \U$3896 ( \4273 , \2607 , RIae76208_37);
and \U$3897 ( \4274 , RIae76a78_55, \2605 );
nor \U$3898 ( \4275 , \4273 , \4274 );
and \U$3899 ( \4276 , \4275 , \2611 );
not \U$3900 ( \4277 , \4275 );
and \U$3901 ( \4278 , \4277 , \2397 );
nor \U$3902 ( \4279 , \4276 , \4278 );
xor \U$3903 ( \4280 , \4272 , \4279 );
not \U$3904 ( \4281 , \3089 );
and \U$3905 ( \4282 , \2783 , RIae76988_53);
and \U$3906 ( \4283 , RIae767a8_49, \2781 );
nor \U$3907 ( \4284 , \4282 , \4283 );
not \U$3908 ( \4285 , \4284 );
or \U$3909 ( \4286 , \4281 , \4285 );
or \U$3910 ( \4287 , \4284 , \2789 );
nand \U$3911 ( \4288 , \4286 , \4287 );
and \U$3912 ( \4289 , \4280 , \4288 );
and \U$3913 ( \4290 , \4272 , \4279 );
or \U$3914 ( \4291 , \4289 , \4290 );
and \U$3915 ( \4292 , \4265 , \4291 );
and \U$3916 ( \4293 , \4231 , \4264 );
or \U$3917 ( \4294 , \4292 , \4293 );
not \U$3918 ( \4295 , \787 );
and \U$3919 ( \4296 , \883 , RIae756c8_13);
and \U$3920 ( \4297 , RIae75218_3, \881 );
nor \U$3921 ( \4298 , \4296 , \4297 );
not \U$3922 ( \4299 , \4298 );
or \U$3923 ( \4300 , \4295 , \4299 );
or \U$3924 ( \4301 , \4298 , \787 );
nand \U$3925 ( \4302 , \4300 , \4301 );
and \U$3926 ( \4303 , \672 , RIae754e8_9);
and \U$3927 ( \4304 , RIae757b8_15, \670 );
nor \U$3928 ( \4305 , \4303 , \4304 );
and \U$3929 ( \4306 , \4305 , \588 );
not \U$3930 ( \4307 , \4305 );
and \U$3931 ( \4308 , \4307 , \587 );
nor \U$3932 ( \4309 , \4306 , \4308 );
xor \U$3933 ( \4310 , \4302 , \4309 );
and \U$3934 ( \4311 , \1138 , RIae75128_1);
and \U$3935 ( \4312 , RIae75308_5, \1136 );
nor \U$3936 ( \4313 , \4311 , \4312 );
and \U$3937 ( \4314 , \4313 , \1012 );
not \U$3938 ( \4315 , \4313 );
and \U$3939 ( \4316 , \4315 , \1142 );
nor \U$3940 ( \4317 , \4314 , \4316 );
and \U$3941 ( \4318 , \4310 , \4317 );
and \U$3942 ( \4319 , \4302 , \4309 );
or \U$3943 ( \4320 , \4318 , \4319 );
nand \U$3944 ( \4321 , RIae75b78_23, RIae78b48_125);
and \U$3945 ( \4322 , \384 , RIae75a88_21);
and \U$3946 ( \4323 , RIae75998_19, \382 );
nor \U$3947 ( \4324 , \4322 , \4323 );
not \U$3948 ( \4325 , \4324 );
not \U$3949 ( \4326 , \388 );
and \U$3950 ( \4327 , \4325 , \4326 );
and \U$3951 ( \4328 , \4324 , \392 );
nor \U$3952 ( \4329 , \4327 , \4328 );
nand \U$3953 ( \4330 , \4321 , \4329 );
xor \U$3954 ( \4331 , \4320 , \4330 );
not \U$3955 ( \4332 , \400 );
and \U$3956 ( \4333 , \436 , RIae758a8_17);
and \U$3957 ( \4334 , RIae75f38_31, \434 );
nor \U$3958 ( \4335 , \4333 , \4334 );
not \U$3959 ( \4336 , \4335 );
or \U$3960 ( \4337 , \4332 , \4336 );
or \U$3961 ( \4338 , \4335 , \402 );
nand \U$3962 ( \4339 , \4337 , \4338 );
not \U$3963 ( \4340 , \471 );
and \U$3964 ( \4341 , \514 , RIae75e48_29);
and \U$3965 ( \4342 , RIae75c68_25, \512 );
nor \U$3966 ( \4343 , \4341 , \4342 );
not \U$3967 ( \4344 , \4343 );
or \U$3968 ( \4345 , \4340 , \4344 );
or \U$3969 ( \4346 , \4343 , \471 );
nand \U$3970 ( \4347 , \4345 , \4346 );
xor \U$3971 ( \4348 , \4339 , \4347 );
and \U$3972 ( \4349 , \558 , RIae75d58_27);
and \U$3973 ( \4350 , RIae755d8_11, \556 );
nor \U$3974 ( \4351 , \4349 , \4350 );
and \U$3975 ( \4352 , \4351 , \504 );
not \U$3976 ( \4353 , \4351 );
and \U$3977 ( \4354 , \4353 , \562 );
nor \U$3978 ( \4355 , \4352 , \4354 );
and \U$3979 ( \4356 , \4348 , \4355 );
and \U$3980 ( \4357 , \4339 , \4347 );
or \U$3981 ( \4358 , \4356 , \4357 );
and \U$3982 ( \4359 , \4331 , \4358 );
and \U$3983 ( \4360 , \4320 , \4330 );
or \U$3984 ( \4361 , \4359 , \4360 );
xor \U$3985 ( \4362 , \4294 , \4361 );
xor \U$3986 ( \4363 , \4077 , \4084 );
xor \U$3987 ( \4364 , \4363 , \4093 );
xor \U$3988 ( \4365 , \4060 , \4068 );
xor \U$3989 ( \4366 , \4364 , \4365 );
xor \U$3990 ( \4367 , \4039 , \4047 );
xor \U$3991 ( \4368 , \4367 , \4055 );
and \U$3992 ( \4369 , \4366 , \4368 );
and \U$3993 ( \4370 , \4364 , \4365 );
or \U$3994 ( \4371 , \4369 , \4370 );
and \U$3995 ( \4372 , \4362 , \4371 );
and \U$3996 ( \4373 , \4294 , \4361 );
or \U$3997 ( \4374 , \4372 , \4373 );
xor \U$3998 ( \4375 , \4058 , \4069 );
xor \U$3999 ( \4376 , \4375 , \4096 );
xor \U$4000 ( \4377 , \3978 , \4001 );
xor \U$4001 ( \4378 , \4377 , \4028 );
and \U$4002 ( \4379 , \4376 , \4378 );
xor \U$4003 ( \4380 , \4374 , \4379 );
xor \U$4004 ( \4381 , \3985 , \3989 );
xor \U$4005 ( \4382 , \4381 , \3998 );
xor \U$4006 ( \4383 , \3960 , \3967 );
xor \U$4007 ( \4384 , \4383 , \3975 );
and \U$4008 ( \4385 , \4382 , \4384 );
xor \U$4009 ( \4386 , \4010 , \4017 );
xor \U$4010 ( \4387 , \4386 , \4025 );
xor \U$4011 ( \4388 , \3960 , \3967 );
xor \U$4012 ( \4389 , \4388 , \3975 );
and \U$4013 ( \4390 , \4387 , \4389 );
and \U$4014 ( \4391 , \4382 , \4387 );
or \U$4015 ( \4392 , \4385 , \4390 , \4391 );
xor \U$4016 ( \4393 , \4102 , \3796 );
xor \U$4017 ( \4394 , \4393 , \4105 );
and \U$4018 ( \4395 , \4392 , \4394 );
not \U$4019 ( \4396 , \4151 );
xor \U$4020 ( \4397 , \4156 , \4140 );
not \U$4021 ( \4398 , \4397 );
or \U$4022 ( \4399 , \4396 , \4398 );
or \U$4023 ( \4400 , \4397 , \4151 );
nand \U$4024 ( \4401 , \4399 , \4400 );
xor \U$4025 ( \4402 , \4102 , \3796 );
xor \U$4026 ( \4403 , \4402 , \4105 );
and \U$4027 ( \4404 , \4401 , \4403 );
and \U$4028 ( \4405 , \4392 , \4401 );
or \U$4029 ( \4406 , \4395 , \4404 , \4405 );
and \U$4030 ( \4407 , \4380 , \4406 );
and \U$4031 ( \4408 , \4374 , \4379 );
or \U$4032 ( \4409 , \4407 , \4408 );
xor \U$4033 ( \4410 , \4206 , \4409 );
xor \U$4034 ( \4411 , \4113 , \4115 );
xor \U$4035 ( \4412 , \4031 , \4099 );
xor \U$4036 ( \4413 , \4412 , \4108 );
and \U$4037 ( \4414 , \4411 , \4413 );
not \U$4038 ( \4415 , \4122 );
xor \U$4039 ( \4416 , \4158 , \4127 );
not \U$4040 ( \4417 , \4416 );
or \U$4041 ( \4418 , \4415 , \4417 );
or \U$4042 ( \4419 , \4416 , \4122 );
nand \U$4043 ( \4420 , \4418 , \4419 );
xor \U$4044 ( \4421 , \4031 , \4099 );
xor \U$4045 ( \4422 , \4421 , \4108 );
and \U$4046 ( \4423 , \4420 , \4422 );
and \U$4047 ( \4424 , \4411 , \4420 );
or \U$4048 ( \4425 , \4414 , \4423 , \4424 );
and \U$4049 ( \4426 , \4410 , \4425 );
and \U$4050 ( \4427 , \4206 , \4409 );
nor \U$4051 ( \4428 , \4426 , \4427 );
xor \U$4052 ( \4429 , \3860 , \3890 );
xor \U$4053 ( \4430 , \4429 , \3905 );
xor \U$4054 ( \4431 , \4428 , \4430 );
xor \U$4055 ( \4432 , \3953 , \4162 );
xor \U$4056 ( \4433 , \4432 , \4165 );
and \U$4057 ( \4434 , \4431 , \4433 );
and \U$4058 ( \4435 , \4428 , \4430 );
or \U$4059 ( \4436 , \4434 , \4435 );
nor \U$4060 ( \4437 , \4200 , \4436 );
and \U$4061 ( \4438 , \4189 , \4437 );
xor \U$4062 ( \4439 , \4437 , \4189 );
xor \U$4063 ( \4440 , \4231 , \4264 );
xor \U$4064 ( \4441 , \4440 , \4291 );
xor \U$4065 ( \4442 , \4320 , \4330 );
xor \U$4066 ( \4443 , \4442 , \4358 );
xor \U$4067 ( \4444 , \4441 , \4443 );
not \U$4068 ( \4445 , \4444 );
and \U$4069 ( \4446 , \1939 , RIae766b8_47);
and \U$4070 ( \4447 , RIae765c8_45, \1937 );
nor \U$4071 ( \4448 , \4446 , \4447 );
and \U$4072 ( \4449 , \4448 , \1734 );
not \U$4073 ( \4450 , \4448 );
and \U$4074 ( \4451 , \4450 , \1735 );
nor \U$4075 ( \4452 , \4449 , \4451 );
and \U$4076 ( \4453 , \2224 , RIae76118_35);
and \U$4077 ( \4454 , RIae76028_33, \2222 );
nor \U$4078 ( \4455 , \4453 , \4454 );
and \U$4079 ( \4456 , \4455 , \2060 );
not \U$4080 ( \4457 , \4455 );
and \U$4081 ( \4458 , \4457 , \2061 );
nor \U$4082 ( \4459 , \4456 , \4458 );
xor \U$4083 ( \4460 , \4452 , \4459 );
and \U$4084 ( \4461 , \1593 , RIae763e8_41);
and \U$4085 ( \4462 , RIae764d8_43, \1591 );
nor \U$4086 ( \4463 , \4461 , \4462 );
and \U$4087 ( \4464 , \4463 , \1488 );
not \U$4088 ( \4465 , \4463 );
and \U$4089 ( \4466 , \4465 , \1498 );
nor \U$4090 ( \4467 , \4464 , \4466 );
and \U$4091 ( \4468 , \4460 , \4467 );
and \U$4092 ( \4469 , \4452 , \4459 );
nor \U$4093 ( \4470 , \4468 , \4469 );
and \U$4094 ( \4471 , \3730 , RIae76b68_57);
and \U$4095 ( \4472 , RIae78a58_123, \3728 );
nor \U$4096 ( \4473 , \4471 , \4472 );
and \U$4097 ( \4474 , \4473 , \3422 );
not \U$4098 ( \4475 , \4473 );
and \U$4099 ( \4476 , \4475 , \3732 );
nor \U$4100 ( \4477 , \4474 , \4476 );
not \U$4101 ( \4478 , RIae79ca0_162);
not \U$4102 ( \4479 , RIae79d18_163);
or \U$4103 ( \4480 , \4478 , \4479 );
nand \U$4104 ( \4481 , \4480 , RIae79c28_161);
not \U$4105 ( \4482 , \4481 );
or \U$4106 ( \4483 , \4477 , \4482 );
not \U$4107 ( \4484 , \4482 );
not \U$4108 ( \4485 , \4477 );
or \U$4109 ( \4486 , \4484 , \4485 );
and \U$4110 ( \4487 , \4247 , RIae78cb0_128);
and \U$4111 ( \4488 , RIae78da0_130, \4245 );
nor \U$4112 ( \4489 , \4487 , \4488 );
and \U$4113 ( \4490 , \4489 , \3989 );
not \U$4114 ( \4491 , \4489 );
and \U$4115 ( \4492 , \4491 , \4251 );
nor \U$4116 ( \4493 , \4490 , \4492 );
nand \U$4117 ( \4494 , \4486 , \4493 );
nand \U$4118 ( \4495 , \4483 , \4494 );
xor \U$4119 ( \4496 , \4470 , \4495 );
and \U$4120 ( \4497 , \2607 , RIae762f8_39);
and \U$4121 ( \4498 , RIae76208_37, \2605 );
nor \U$4122 ( \4499 , \4497 , \4498 );
and \U$4123 ( \4500 , \4499 , \2611 );
not \U$4124 ( \4501 , \4499 );
and \U$4125 ( \4502 , \4501 , \2397 );
nor \U$4126 ( \4503 , \4500 , \4502 );
not \U$4127 ( \4504 , \3089 );
and \U$4128 ( \4505 , \2783 , RIae76a78_55);
and \U$4129 ( \4506 , RIae76988_53, \2781 );
nor \U$4130 ( \4507 , \4505 , \4506 );
not \U$4131 ( \4508 , \4507 );
or \U$4132 ( \4509 , \4504 , \4508 );
or \U$4133 ( \4510 , \4507 , \2789 );
nand \U$4134 ( \4511 , \4509 , \4510 );
xor \U$4135 ( \4512 , \4503 , \4511 );
not \U$4136 ( \4513 , \3218 );
and \U$4137 ( \4514 , \3214 , RIae767a8_49);
and \U$4138 ( \4515 , RIae76898_51, \3212 );
nor \U$4139 ( \4516 , \4514 , \4515 );
not \U$4140 ( \4517 , \4516 );
or \U$4141 ( \4518 , \4513 , \4517 );
or \U$4142 ( \4519 , \4516 , \3218 );
nand \U$4143 ( \4520 , \4518 , \4519 );
and \U$4144 ( \4521 , \4512 , \4520 );
and \U$4145 ( \4522 , \4503 , \4511 );
or \U$4146 ( \4523 , \4521 , \4522 );
and \U$4147 ( \4524 , \4496 , \4523 );
and \U$4148 ( \4525 , \4470 , \4495 );
or \U$4149 ( \4526 , \4524 , \4525 );
and \U$4150 ( \4527 , \672 , RIae755d8_11);
and \U$4151 ( \4528 , RIae754e8_9, \670 );
nor \U$4152 ( \4529 , \4527 , \4528 );
and \U$4153 ( \4530 , \4529 , \588 );
not \U$4154 ( \4531 , \4529 );
and \U$4155 ( \4532 , \4531 , \587 );
nor \U$4156 ( \4533 , \4530 , \4532 );
not \U$4157 ( \4534 , \469 );
and \U$4158 ( \4535 , \514 , RIae75f38_31);
and \U$4159 ( \4536 , RIae75e48_29, \512 );
nor \U$4160 ( \4537 , \4535 , \4536 );
not \U$4161 ( \4538 , \4537 );
or \U$4162 ( \4539 , \4534 , \4538 );
or \U$4163 ( \4540 , \4537 , \469 );
nand \U$4164 ( \4541 , \4539 , \4540 );
xor \U$4165 ( \4542 , \4533 , \4541 );
and \U$4166 ( \4543 , \558 , RIae75c68_25);
and \U$4167 ( \4544 , RIae75d58_27, \556 );
nor \U$4168 ( \4545 , \4543 , \4544 );
and \U$4169 ( \4546 , \4545 , \504 );
not \U$4170 ( \4547 , \4545 );
and \U$4171 ( \4548 , \4547 , \562 );
nor \U$4172 ( \4549 , \4546 , \4548 );
and \U$4173 ( \4550 , \4542 , \4549 );
and \U$4174 ( \4551 , \4533 , \4541 );
or \U$4175 ( \4552 , \4550 , \4551 );
and \U$4176 ( \4553 , \436 , RIae75998_19);
and \U$4177 ( \4554 , RIae758a8_17, \434 );
nor \U$4178 ( \4555 , \4553 , \4554 );
not \U$4179 ( \4556 , \4555 );
not \U$4180 ( \4557 , \402 );
and \U$4181 ( \4558 , \4556 , \4557 );
and \U$4182 ( \4559 , \4555 , \400 );
nor \U$4183 ( \4560 , \4558 , \4559 );
nand \U$4184 ( \4561 , RIae78698_115, RIae78b48_125);
or \U$4185 ( \4562 , \4560 , \4561 );
not \U$4186 ( \4563 , \4561 );
not \U$4187 ( \4564 , \4560 );
or \U$4188 ( \4565 , \4563 , \4564 );
not \U$4189 ( \4566 , \392 );
and \U$4190 ( \4567 , \384 , RIae75b78_23);
and \U$4191 ( \4568 , RIae75a88_21, \382 );
nor \U$4192 ( \4569 , \4567 , \4568 );
not \U$4193 ( \4570 , \4569 );
or \U$4194 ( \4571 , \4566 , \4570 );
or \U$4195 ( \4572 , \4569 , \388 );
nand \U$4196 ( \4573 , \4571 , \4572 );
nand \U$4197 ( \4574 , \4565 , \4573 );
nand \U$4198 ( \4575 , \4562 , \4574 );
xor \U$4199 ( \4576 , \4552 , \4575 );
and \U$4200 ( \4577 , \1138 , RIae75218_3);
and \U$4201 ( \4578 , RIae75128_1, \1136 );
nor \U$4202 ( \4579 , \4577 , \4578 );
and \U$4203 ( \4580 , \4579 , \1142 );
not \U$4204 ( \4581 , \4579 );
and \U$4205 ( \4582 , \4581 , \1012 );
nor \U$4206 ( \4583 , \4580 , \4582 );
and \U$4207 ( \4584 , \1376 , RIae75308_5);
and \U$4208 ( \4585 , RIae753f8_7, \1374 );
nor \U$4209 ( \4586 , \4584 , \4585 );
and \U$4210 ( \4587 , \4586 , \1261 );
not \U$4211 ( \4588 , \4586 );
and \U$4212 ( \4589 , \4588 , \1380 );
nor \U$4213 ( \4590 , \4587 , \4589 );
xor \U$4214 ( \4591 , \4583 , \4590 );
and \U$4215 ( \4592 , \883 , RIae757b8_15);
and \U$4216 ( \4593 , RIae756c8_13, \881 );
nor \U$4217 ( \4594 , \4592 , \4593 );
not \U$4218 ( \4595 , \4594 );
not \U$4219 ( \4596 , \789 );
and \U$4220 ( \4597 , \4595 , \4596 );
and \U$4221 ( \4598 , \4594 , \789 );
nor \U$4222 ( \4599 , \4597 , \4598 );
and \U$4223 ( \4600 , \4591 , \4599 );
and \U$4224 ( \4601 , \4583 , \4590 );
nor \U$4225 ( \4602 , \4600 , \4601 );
and \U$4226 ( \4603 , \4576 , \4602 );
and \U$4227 ( \4604 , \4552 , \4575 );
or \U$4228 ( \4605 , \4603 , \4604 );
xor \U$4229 ( \4606 , \4526 , \4605 );
xor \U$4230 ( \4607 , \4339 , \4347 );
xor \U$4231 ( \4608 , \4607 , \4355 );
or \U$4232 ( \4609 , \4329 , \4321 );
nand \U$4233 ( \4610 , \4609 , \4330 );
xor \U$4234 ( \4611 , \4608 , \4610 );
xor \U$4235 ( \4612 , \4302 , \4309 );
xor \U$4236 ( \4613 , \4612 , \4317 );
and \U$4237 ( \4614 , \4611 , \4613 );
and \U$4238 ( \4615 , \4608 , \4610 );
or \U$4239 ( \4616 , \4614 , \4615 );
xor \U$4240 ( \4617 , \4606 , \4616 );
not \U$4241 ( \4618 , \4617 );
or \U$4242 ( \4619 , \4445 , \4618 );
or \U$4243 ( \4620 , \4617 , \4444 );
xor \U$4244 ( \4621 , \4364 , \4365 );
xor \U$4245 ( \4622 , \4621 , \4368 );
xor \U$4246 ( \4623 , \4239 , \4253 );
xor \U$4247 ( \4624 , \4623 , \4261 );
xor \U$4248 ( \4625 , \4272 , \4279 );
xor \U$4249 ( \4626 , \4625 , \4288 );
and \U$4250 ( \4627 , \4624 , \4626 );
xor \U$4251 ( \4628 , \4213 , \4220 );
xor \U$4252 ( \4629 , \4628 , \4228 );
xor \U$4253 ( \4630 , \4272 , \4279 );
xor \U$4254 ( \4631 , \4630 , \4288 );
and \U$4255 ( \4632 , \4629 , \4631 );
and \U$4256 ( \4633 , \4624 , \4629 );
or \U$4257 ( \4634 , \4627 , \4632 , \4633 );
xor \U$4258 ( \4635 , \3960 , \3967 );
xor \U$4259 ( \4636 , \4635 , \3975 );
xor \U$4260 ( \4637 , \4382 , \4387 );
xor \U$4261 ( \4638 , \4636 , \4637 );
xor \U$4262 ( \4639 , \4634 , \4638 );
xor \U$4263 ( \4640 , \4622 , \4639 );
nand \U$4264 ( \4641 , \4620 , \4640 );
nand \U$4265 ( \4642 , \4619 , \4641 );
xor \U$4266 ( \4643 , \4470 , \4495 );
xor \U$4267 ( \4644 , \4643 , \4523 );
xor \U$4268 ( \4645 , \4552 , \4575 );
xor \U$4269 ( \4646 , \4645 , \4602 );
and \U$4270 ( \4647 , \4644 , \4646 );
not \U$4271 ( \4648 , \4647 );
and \U$4272 ( \4649 , \1939 , RIae764d8_43);
and \U$4273 ( \4650 , RIae766b8_47, \1937 );
nor \U$4274 ( \4651 , \4649 , \4650 );
and \U$4275 ( \4652 , \4651 , \1735 );
not \U$4276 ( \4653 , \4651 );
and \U$4277 ( \4654 , \4653 , \1734 );
nor \U$4278 ( \4655 , \4652 , \4654 );
and \U$4279 ( \4656 , \1593 , RIae753f8_7);
and \U$4280 ( \4657 , RIae763e8_41, \1591 );
nor \U$4281 ( \4658 , \4656 , \4657 );
and \U$4282 ( \4659 , \4658 , \1498 );
not \U$4283 ( \4660 , \4658 );
and \U$4284 ( \4661 , \4660 , \1488 );
nor \U$4285 ( \4662 , \4659 , \4661 );
xor \U$4286 ( \4663 , \4655 , \4662 );
and \U$4287 ( \4664 , \2224 , RIae765c8_45);
and \U$4288 ( \4665 , RIae76118_35, \2222 );
nor \U$4289 ( \4666 , \4664 , \4665 );
and \U$4290 ( \4667 , \4666 , \2061 );
not \U$4291 ( \4668 , \4666 );
and \U$4292 ( \4669 , \4668 , \2060 );
nor \U$4293 ( \4670 , \4667 , \4669 );
and \U$4294 ( \4671 , \4663 , \4670 );
and \U$4295 ( \4672 , \4655 , \4662 );
or \U$4296 ( \4673 , \4671 , \4672 );
and \U$4297 ( \4674 , \3730 , RIae76898_51);
and \U$4298 ( \4675 , RIae76b68_57, \3728 );
nor \U$4299 ( \4676 , \4674 , \4675 );
and \U$4300 ( \4677 , \4676 , \3732 );
not \U$4301 ( \4678 , \4676 );
and \U$4302 ( \4679 , \4678 , \3422 );
nor \U$4303 ( \4680 , \4677 , \4679 );
and \U$4304 ( \4681 , RIae79c28_161, RIae79d18_163);
not \U$4305 ( \4682 , RIae79d18_163);
nor \U$4306 ( \4683 , \4682 , RIae79ca0_162);
not \U$4307 ( \4684 , RIae79ca0_162);
nor \U$4308 ( \4685 , \4684 , RIae79d18_163);
or \U$4309 ( \4686 , \4683 , \4685 );
nor \U$4310 ( \4687 , RIae79c28_161, RIae79d18_163);
nor \U$4311 ( \4688 , \4681 , \4686 , \4687 );
nand \U$4312 ( \4689 , RIae78da0_130, \4688 );
and \U$4313 ( \4690 , \4689 , \4481 );
not \U$4314 ( \4691 , \4689 );
and \U$4315 ( \4692 , \4691 , \4482 );
nor \U$4316 ( \4693 , \4690 , \4692 );
xor \U$4317 ( \4694 , \4680 , \4693 );
and \U$4318 ( \4695 , \4247 , RIae78a58_123);
and \U$4319 ( \4696 , RIae78cb0_128, \4245 );
nor \U$4320 ( \4697 , \4695 , \4696 );
and \U$4321 ( \4698 , \4697 , \3989 );
not \U$4322 ( \4699 , \4697 );
and \U$4323 ( \4700 , \4699 , \4251 );
nor \U$4324 ( \4701 , \4698 , \4700 );
and \U$4325 ( \4702 , \4694 , \4701 );
and \U$4326 ( \4703 , \4680 , \4693 );
or \U$4327 ( \4704 , \4702 , \4703 );
xor \U$4328 ( \4705 , \4673 , \4704 );
and \U$4329 ( \4706 , \2607 , RIae76028_33);
and \U$4330 ( \4707 , RIae762f8_39, \2605 );
nor \U$4331 ( \4708 , \4706 , \4707 );
and \U$4332 ( \4709 , \4708 , \2611 );
not \U$4333 ( \4710 , \4708 );
and \U$4334 ( \4711 , \4710 , \2397 );
nor \U$4335 ( \4712 , \4709 , \4711 );
not \U$4336 ( \4713 , \2789 );
and \U$4337 ( \4714 , \2783 , RIae76208_37);
and \U$4338 ( \4715 , RIae76a78_55, \2781 );
nor \U$4339 ( \4716 , \4714 , \4715 );
not \U$4340 ( \4717 , \4716 );
or \U$4341 ( \4718 , \4713 , \4717 );
or \U$4342 ( \4719 , \4716 , \3089 );
nand \U$4343 ( \4720 , \4718 , \4719 );
xor \U$4344 ( \4721 , \4712 , \4720 );
not \U$4345 ( \4722 , \3218 );
and \U$4346 ( \4723 , \3214 , RIae76988_53);
and \U$4347 ( \4724 , RIae767a8_49, \3212 );
nor \U$4348 ( \4725 , \4723 , \4724 );
not \U$4349 ( \4726 , \4725 );
or \U$4350 ( \4727 , \4722 , \4726 );
or \U$4351 ( \4728 , \4725 , \2774 );
nand \U$4352 ( \4729 , \4727 , \4728 );
and \U$4353 ( \4730 , \4721 , \4729 );
and \U$4354 ( \4731 , \4712 , \4720 );
or \U$4355 ( \4732 , \4730 , \4731 );
and \U$4356 ( \4733 , \4705 , \4732 );
and \U$4357 ( \4734 , \4673 , \4704 );
or \U$4358 ( \4735 , \4733 , \4734 );
and \U$4359 ( \4736 , \514 , RIae758a8_17);
and \U$4360 ( \4737 , RIae75f38_31, \512 );
nor \U$4361 ( \4738 , \4736 , \4737 );
not \U$4362 ( \4739 , \4738 );
not \U$4363 ( \4740 , \469 );
and \U$4364 ( \4741 , \4739 , \4740 );
and \U$4365 ( \4742 , \4738 , \471 );
nor \U$4366 ( \4743 , \4741 , \4742 );
and \U$4367 ( \4744 , \672 , RIae75d58_27);
and \U$4368 ( \4745 , RIae755d8_11, \670 );
nor \U$4369 ( \4746 , \4744 , \4745 );
and \U$4370 ( \4747 , \4746 , \587 );
not \U$4371 ( \4748 , \4746 );
and \U$4372 ( \4749 , \4748 , \588 );
nor \U$4373 ( \4750 , \4747 , \4749 );
or \U$4374 ( \4751 , \4743 , \4750 );
not \U$4375 ( \4752 , \4750 );
not \U$4376 ( \4753 , \4743 );
or \U$4377 ( \4754 , \4752 , \4753 );
and \U$4378 ( \4755 , \558 , RIae75e48_29);
and \U$4379 ( \4756 , RIae75c68_25, \556 );
nor \U$4380 ( \4757 , \4755 , \4756 );
and \U$4381 ( \4758 , \4757 , \504 );
not \U$4382 ( \4759 , \4757 );
and \U$4383 ( \4760 , \4759 , \562 );
nor \U$4384 ( \4761 , \4758 , \4760 );
nand \U$4385 ( \4762 , \4754 , \4761 );
nand \U$4386 ( \4763 , \4751 , \4762 );
and \U$4387 ( \4764 , \436 , RIae75a88_21);
and \U$4388 ( \4765 , RIae75998_19, \434 );
nor \U$4389 ( \4766 , \4764 , \4765 );
not \U$4390 ( \4767 , \4766 );
not \U$4391 ( \4768 , \402 );
and \U$4392 ( \4769 , \4767 , \4768 );
and \U$4393 ( \4770 , \4766 , \400 );
nor \U$4394 ( \4771 , \4769 , \4770 );
nand \U$4395 ( \4772 , RIae78788_117, RIae78b48_125);
or \U$4396 ( \4773 , \4771 , \4772 );
not \U$4397 ( \4774 , \4772 );
not \U$4398 ( \4775 , \4771 );
or \U$4399 ( \4776 , \4774 , \4775 );
not \U$4400 ( \4777 , \392 );
and \U$4401 ( \4778 , \384 , RIae78698_115);
and \U$4402 ( \4779 , RIae75b78_23, \382 );
nor \U$4403 ( \4780 , \4778 , \4779 );
not \U$4404 ( \4781 , \4780 );
or \U$4405 ( \4782 , \4777 , \4781 );
or \U$4406 ( \4783 , \4780 , \392 );
nand \U$4407 ( \4784 , \4782 , \4783 );
nand \U$4408 ( \4785 , \4776 , \4784 );
nand \U$4409 ( \4786 , \4773 , \4785 );
xor \U$4410 ( \4787 , \4763 , \4786 );
not \U$4411 ( \4788 , \789 );
and \U$4412 ( \4789 , \883 , RIae754e8_9);
and \U$4413 ( \4790 , RIae757b8_15, \881 );
nor \U$4414 ( \4791 , \4789 , \4790 );
not \U$4415 ( \4792 , \4791 );
or \U$4416 ( \4793 , \4788 , \4792 );
or \U$4417 ( \4794 , \4791 , \787 );
nand \U$4418 ( \4795 , \4793 , \4794 );
and \U$4419 ( \4796 , \1138 , RIae756c8_13);
and \U$4420 ( \4797 , RIae75218_3, \1136 );
nor \U$4421 ( \4798 , \4796 , \4797 );
and \U$4422 ( \4799 , \4798 , \1012 );
not \U$4423 ( \4800 , \4798 );
and \U$4424 ( \4801 , \4800 , \1142 );
nor \U$4425 ( \4802 , \4799 , \4801 );
xor \U$4426 ( \4803 , \4795 , \4802 );
and \U$4427 ( \4804 , \1376 , RIae75128_1);
and \U$4428 ( \4805 , RIae75308_5, \1374 );
nor \U$4429 ( \4806 , \4804 , \4805 );
and \U$4430 ( \4807 , \4806 , \1380 );
not \U$4431 ( \4808 , \4806 );
and \U$4432 ( \4809 , \4808 , \1261 );
nor \U$4433 ( \4810 , \4807 , \4809 );
and \U$4434 ( \4811 , \4803 , \4810 );
and \U$4435 ( \4812 , \4795 , \4802 );
or \U$4436 ( \4813 , \4811 , \4812 );
and \U$4437 ( \4814 , \4787 , \4813 );
and \U$4438 ( \4815 , \4763 , \4786 );
or \U$4439 ( \4816 , \4814 , \4815 );
xor \U$4440 ( \4817 , \4735 , \4816 );
not \U$4441 ( \4818 , \4560 );
not \U$4442 ( \4819 , \4573 );
or \U$4443 ( \4820 , \4818 , \4819 );
or \U$4444 ( \4821 , \4560 , \4573 );
nand \U$4445 ( \4822 , \4820 , \4821 );
not \U$4446 ( \4823 , \4822 );
not \U$4447 ( \4824 , \4561 );
and \U$4448 ( \4825 , \4823 , \4824 );
and \U$4449 ( \4826 , \4822 , \4561 );
nor \U$4450 ( \4827 , \4825 , \4826 );
xor \U$4451 ( \4828 , \4583 , \4590 );
xor \U$4452 ( \4829 , \4828 , \4599 );
or \U$4453 ( \4830 , \4827 , \4829 );
not \U$4454 ( \4831 , \4829 );
not \U$4455 ( \4832 , \4827 );
or \U$4456 ( \4833 , \4831 , \4832 );
xor \U$4457 ( \4834 , \4533 , \4541 );
xor \U$4458 ( \4835 , \4834 , \4549 );
nand \U$4459 ( \4836 , \4833 , \4835 );
nand \U$4460 ( \4837 , \4830 , \4836 );
and \U$4461 ( \4838 , \4817 , \4837 );
and \U$4462 ( \4839 , \4735 , \4816 );
or \U$4463 ( \4840 , \4838 , \4839 );
not \U$4464 ( \4841 , \4840 );
or \U$4465 ( \4842 , \4648 , \4841 );
or \U$4466 ( \4843 , \4840 , \4647 );
and \U$4467 ( \4844 , \4493 , \4481 );
not \U$4468 ( \4845 , \4493 );
and \U$4469 ( \4846 , \4845 , \4482 );
nor \U$4470 ( \4847 , \4844 , \4846 );
not \U$4471 ( \4848 , \4847 );
not \U$4472 ( \4849 , \4477 );
and \U$4473 ( \4850 , \4848 , \4849 );
and \U$4474 ( \4851 , \4847 , \4477 );
nor \U$4475 ( \4852 , \4850 , \4851 );
xor \U$4476 ( \4853 , \4452 , \4459 );
xor \U$4477 ( \4854 , \4853 , \4467 );
or \U$4478 ( \4855 , \4852 , \4854 );
not \U$4479 ( \4856 , \4854 );
not \U$4480 ( \4857 , \4852 );
or \U$4481 ( \4858 , \4856 , \4857 );
xor \U$4482 ( \4859 , \4503 , \4511 );
xor \U$4483 ( \4860 , \4859 , \4520 );
nand \U$4484 ( \4861 , \4858 , \4860 );
nand \U$4485 ( \4862 , \4855 , \4861 );
xor \U$4486 ( \4863 , \4608 , \4610 );
xor \U$4487 ( \4864 , \4863 , \4613 );
and \U$4488 ( \4865 , \4862 , \4864 );
xor \U$4489 ( \4866 , \4272 , \4279 );
xor \U$4490 ( \4867 , \4866 , \4288 );
xor \U$4491 ( \4868 , \4624 , \4629 );
xor \U$4492 ( \4869 , \4867 , \4868 );
xor \U$4493 ( \4870 , \4608 , \4610 );
xor \U$4494 ( \4871 , \4870 , \4613 );
and \U$4495 ( \4872 , \4869 , \4871 );
and \U$4496 ( \4873 , \4862 , \4869 );
or \U$4497 ( \4874 , \4865 , \4872 , \4873 );
nand \U$4498 ( \4875 , \4843 , \4874 );
nand \U$4499 ( \4876 , \4842 , \4875 );
xor \U$4500 ( \4877 , \4642 , \4876 );
xor \U$4501 ( \4878 , \4294 , \4361 );
xor \U$4502 ( \4879 , \4878 , \4371 );
xor \U$4503 ( \4880 , \4376 , \4378 );
xor \U$4504 ( \4881 , \4102 , \3796 );
xor \U$4505 ( \4882 , \4881 , \4105 );
xor \U$4506 ( \4883 , \4392 , \4401 );
xor \U$4507 ( \4884 , \4882 , \4883 );
xor \U$4508 ( \4885 , \4880 , \4884 );
xor \U$4509 ( \4886 , \4879 , \4885 );
and \U$4510 ( \4887 , \4877 , \4886 );
and \U$4511 ( \4888 , \4642 , \4876 );
or \U$4512 ( \4889 , \4887 , \4888 );
xor \U$4513 ( \4890 , \4374 , \4379 );
xor \U$4514 ( \4891 , \4890 , \4406 );
xor \U$4515 ( \4892 , \4889 , \4891 );
xor \U$4516 ( \4893 , \4294 , \4361 );
xor \U$4517 ( \4894 , \4893 , \4371 );
and \U$4518 ( \4895 , \4880 , \4894 );
xor \U$4519 ( \4896 , \4294 , \4361 );
xor \U$4520 ( \4897 , \4896 , \4371 );
and \U$4521 ( \4898 , \4884 , \4897 );
and \U$4522 ( \4899 , \4880 , \4884 );
or \U$4523 ( \4900 , \4895 , \4898 , \4899 );
xor \U$4524 ( \4901 , \4526 , \4605 );
and \U$4525 ( \4902 , \4901 , \4616 );
and \U$4526 ( \4903 , \4526 , \4605 );
or \U$4527 ( \4904 , \4902 , \4903 );
and \U$4528 ( \4905 , \4441 , \4443 );
xor \U$4529 ( \4906 , \4904 , \4905 );
xor \U$4530 ( \4907 , \4364 , \4365 );
xor \U$4531 ( \4908 , \4907 , \4368 );
and \U$4532 ( \4909 , \4634 , \4908 );
xor \U$4533 ( \4910 , \4364 , \4365 );
xor \U$4534 ( \4911 , \4910 , \4368 );
and \U$4535 ( \4912 , \4638 , \4911 );
and \U$4536 ( \4913 , \4634 , \4638 );
or \U$4537 ( \4914 , \4909 , \4912 , \4913 );
and \U$4538 ( \4915 , \4906 , \4914 );
and \U$4539 ( \4916 , \4904 , \4905 );
or \U$4540 ( \4917 , \4915 , \4916 );
xor \U$4541 ( \4918 , \4900 , \4917 );
xor \U$4542 ( \4919 , \4031 , \4099 );
xor \U$4543 ( \4920 , \4919 , \4108 );
xor \U$4544 ( \4921 , \4411 , \4420 );
xor \U$4545 ( \4922 , \4920 , \4921 );
xor \U$4546 ( \4923 , \4918 , \4922 );
and \U$4547 ( \4924 , \4892 , \4923 );
and \U$4548 ( \4925 , \4889 , \4891 );
or \U$4549 ( \4926 , \4924 , \4925 );
xor \U$4550 ( \4927 , \4206 , \4409 );
xor \U$4551 ( \4928 , \4927 , \4425 );
not \U$4552 ( \4929 , \4116 );
not \U$4553 ( \4930 , \4160 );
not \U$4554 ( \4931 , \4111 );
and \U$4555 ( \4932 , \4930 , \4931 );
and \U$4556 ( \4933 , \4160 , \4111 );
nor \U$4557 ( \4934 , \4932 , \4933 );
not \U$4558 ( \4935 , \4934 );
or \U$4559 ( \4936 , \4929 , \4935 );
or \U$4560 ( \4937 , \4934 , \4116 );
nand \U$4561 ( \4938 , \4936 , \4937 );
xor \U$4562 ( \4939 , \4928 , \4938 );
xor \U$4563 ( \4940 , \4900 , \4917 );
and \U$4564 ( \4941 , \4940 , \4922 );
and \U$4565 ( \4942 , \4900 , \4917 );
or \U$4566 ( \4943 , \4941 , \4942 );
xor \U$4567 ( \4944 , \4939 , \4943 );
xor \U$4568 ( \4945 , \4926 , \4944 );
xor \U$4569 ( \4946 , \4889 , \4891 );
xor \U$4570 ( \4947 , \4946 , \4923 );
not \U$4571 ( \4948 , \4947 );
xor \U$4572 ( \4949 , \4642 , \4876 );
xor \U$4573 ( \4950 , \4949 , \4886 );
xor \U$4574 ( \4951 , \4904 , \4905 );
xor \U$4575 ( \4952 , \4951 , \4914 );
xor \U$4576 ( \4953 , \4950 , \4952 );
xnor \U$4577 ( \4954 , \4617 , \4640 );
not \U$4578 ( \4955 , \4954 );
not \U$4579 ( \4956 , \4444 );
and \U$4580 ( \4957 , \4955 , \4956 );
and \U$4581 ( \4958 , \4954 , \4444 );
nor \U$4582 ( \4959 , \4957 , \4958 );
xor \U$4583 ( \4960 , \4644 , \4646 );
xor \U$4584 ( \4961 , \4735 , \4816 );
xor \U$4585 ( \4962 , \4961 , \4837 );
xor \U$4586 ( \4963 , \4960 , \4962 );
xor \U$4587 ( \4964 , \4608 , \4610 );
xor \U$4588 ( \4965 , \4964 , \4613 );
xor \U$4589 ( \4966 , \4862 , \4869 );
xor \U$4590 ( \4967 , \4965 , \4966 );
and \U$4591 ( \4968 , \4963 , \4967 );
and \U$4592 ( \4969 , \4960 , \4962 );
nor \U$4593 ( \4970 , \4968 , \4969 );
or \U$4594 ( \4971 , \4959 , \4970 );
not \U$4595 ( \4972 , \4970 );
not \U$4596 ( \4973 , \4959 );
or \U$4597 ( \4974 , \4972 , \4973 );
xor \U$4598 ( \4975 , \4673 , \4704 );
xor \U$4599 ( \4976 , \4975 , \4732 );
xor \U$4600 ( \4977 , \4763 , \4786 );
xor \U$4601 ( \4978 , \4977 , \4813 );
and \U$4602 ( \4979 , \4976 , \4978 );
not \U$4603 ( \4980 , \4979 );
and \U$4604 ( \4981 , \2224 , RIae766b8_47);
and \U$4605 ( \4982 , RIae765c8_45, \2222 );
nor \U$4606 ( \4983 , \4981 , \4982 );
and \U$4607 ( \4984 , \4983 , \2061 );
not \U$4608 ( \4985 , \4983 );
and \U$4609 ( \4986 , \4985 , \2060 );
nor \U$4610 ( \4987 , \4984 , \4986 );
and \U$4611 ( \4988 , \1939 , RIae763e8_41);
and \U$4612 ( \4989 , RIae764d8_43, \1937 );
nor \U$4613 ( \4990 , \4988 , \4989 );
and \U$4614 ( \4991 , \4990 , \1735 );
not \U$4615 ( \4992 , \4990 );
and \U$4616 ( \4993 , \4992 , \1734 );
nor \U$4617 ( \4994 , \4991 , \4993 );
xor \U$4618 ( \4995 , \4987 , \4994 );
and \U$4619 ( \4996 , \2607 , RIae76118_35);
and \U$4620 ( \4997 , RIae76028_33, \2605 );
nor \U$4621 ( \4998 , \4996 , \4997 );
and \U$4622 ( \4999 , \4998 , \2611 );
not \U$4623 ( \5000 , \4998 );
and \U$4624 ( \5001 , \5000 , \2397 );
nor \U$4625 ( \5002 , \4999 , \5001 );
and \U$4626 ( \5003 , \4995 , \5002 );
and \U$4627 ( \5004 , \4987 , \4994 );
or \U$4628 ( \5005 , \5003 , \5004 );
and \U$4629 ( \5006 , \4688 , RIae78cb0_128);
and \U$4630 ( \5007 , RIae78da0_130, \4686 );
nor \U$4631 ( \5008 , \5006 , \5007 );
and \U$4632 ( \5009 , \5008 , \4481 );
not \U$4633 ( \5010 , \5008 );
and \U$4634 ( \5011 , \5010 , \4482 );
nor \U$4635 ( \5012 , \5009 , \5011 );
not \U$4636 ( \5013 , RIae79d90_164);
not \U$4637 ( \5014 , RIae79e08_165);
or \U$4638 ( \5015 , \5013 , \5014 );
nand \U$4639 ( \5016 , \5015 , RIae79ca0_162);
xor \U$4640 ( \5017 , \5012 , \5016 );
and \U$4641 ( \5018 , \4247 , RIae76b68_57);
and \U$4642 ( \5019 , RIae78a58_123, \4245 );
nor \U$4643 ( \5020 , \5018 , \5019 );
and \U$4644 ( \5021 , \5020 , \3989 );
not \U$4645 ( \5022 , \5020 );
and \U$4646 ( \5023 , \5022 , \4251 );
nor \U$4647 ( \5024 , \5021 , \5023 );
and \U$4648 ( \5025 , \5017 , \5024 );
and \U$4649 ( \5026 , \5012 , \5016 );
or \U$4650 ( \5027 , \5025 , \5026 );
xor \U$4651 ( \5028 , \5005 , \5027 );
and \U$4652 ( \5029 , \3730 , RIae767a8_49);
and \U$4653 ( \5030 , RIae76898_51, \3728 );
nor \U$4654 ( \5031 , \5029 , \5030 );
and \U$4655 ( \5032 , \5031 , \3732 );
not \U$4656 ( \5033 , \5031 );
and \U$4657 ( \5034 , \5033 , \3422 );
nor \U$4658 ( \5035 , \5032 , \5034 );
not \U$4659 ( \5036 , \2789 );
and \U$4660 ( \5037 , \2783 , RIae762f8_39);
and \U$4661 ( \5038 , RIae76208_37, \2781 );
nor \U$4662 ( \5039 , \5037 , \5038 );
not \U$4663 ( \5040 , \5039 );
or \U$4664 ( \5041 , \5036 , \5040 );
or \U$4665 ( \5042 , \5039 , \3089 );
nand \U$4666 ( \5043 , \5041 , \5042 );
xor \U$4667 ( \5044 , \5035 , \5043 );
not \U$4668 ( \5045 , \3218 );
and \U$4669 ( \5046 , \3214 , RIae76a78_55);
and \U$4670 ( \5047 , RIae76988_53, \3212 );
nor \U$4671 ( \5048 , \5046 , \5047 );
not \U$4672 ( \5049 , \5048 );
or \U$4673 ( \5050 , \5045 , \5049 );
or \U$4674 ( \5051 , \5048 , \2774 );
nand \U$4675 ( \5052 , \5050 , \5051 );
and \U$4676 ( \5053 , \5044 , \5052 );
and \U$4677 ( \5054 , \5035 , \5043 );
or \U$4678 ( \5055 , \5053 , \5054 );
and \U$4679 ( \5056 , \5028 , \5055 );
and \U$4680 ( \5057 , \5005 , \5027 );
or \U$4681 ( \5058 , \5056 , \5057 );
not \U$4682 ( \5059 , \4771 );
not \U$4683 ( \5060 , \4784 );
or \U$4684 ( \5061 , \5059 , \5060 );
or \U$4685 ( \5062 , \4771 , \4784 );
nand \U$4686 ( \5063 , \5061 , \5062 );
not \U$4687 ( \5064 , \5063 );
not \U$4688 ( \5065 , \4772 );
and \U$4689 ( \5066 , \5064 , \5065 );
and \U$4690 ( \5067 , \5063 , \4772 );
nor \U$4691 ( \5068 , \5066 , \5067 );
not \U$4692 ( \5069 , \4750 );
not \U$4693 ( \5070 , \4761 );
or \U$4694 ( \5071 , \5069 , \5070 );
or \U$4695 ( \5072 , \4750 , \4761 );
nand \U$4696 ( \5073 , \5071 , \5072 );
not \U$4697 ( \5074 , \5073 );
not \U$4698 ( \5075 , \4743 );
and \U$4699 ( \5076 , \5074 , \5075 );
and \U$4700 ( \5077 , \5073 , \4743 );
nor \U$4701 ( \5078 , \5076 , \5077 );
nand \U$4702 ( \5079 , \5068 , \5078 );
xor \U$4703 ( \5080 , \5058 , \5079 );
and \U$4704 ( \5081 , \1138 , RIae757b8_15);
and \U$4705 ( \5082 , RIae756c8_13, \1136 );
nor \U$4706 ( \5083 , \5081 , \5082 );
and \U$4707 ( \5084 , \5083 , \1012 );
not \U$4708 ( \5085 , \5083 );
and \U$4709 ( \5086 , \5085 , \1142 );
nor \U$4710 ( \5087 , \5084 , \5086 );
and \U$4711 ( \5088 , \1376 , RIae75218_3);
and \U$4712 ( \5089 , RIae75128_1, \1374 );
nor \U$4713 ( \5090 , \5088 , \5089 );
and \U$4714 ( \5091 , \5090 , \1380 );
not \U$4715 ( \5092 , \5090 );
and \U$4716 ( \5093 , \5092 , \1261 );
nor \U$4717 ( \5094 , \5091 , \5093 );
xor \U$4718 ( \5095 , \5087 , \5094 );
and \U$4719 ( \5096 , \1593 , RIae75308_5);
and \U$4720 ( \5097 , RIae753f8_7, \1591 );
nor \U$4721 ( \5098 , \5096 , \5097 );
and \U$4722 ( \5099 , \5098 , \1498 );
not \U$4723 ( \5100 , \5098 );
and \U$4724 ( \5101 , \5100 , \1488 );
nor \U$4725 ( \5102 , \5099 , \5101 );
and \U$4726 ( \5103 , \5095 , \5102 );
and \U$4727 ( \5104 , \5087 , \5094 );
or \U$4728 ( \5105 , \5103 , \5104 );
and \U$4729 ( \5106 , \558 , RIae75f38_31);
and \U$4730 ( \5107 , RIae75e48_29, \556 );
nor \U$4731 ( \5108 , \5106 , \5107 );
and \U$4732 ( \5109 , \5108 , \504 );
not \U$4733 ( \5110 , \5108 );
and \U$4734 ( \5111 , \5110 , \562 );
nor \U$4735 ( \5112 , \5109 , \5111 );
and \U$4736 ( \5113 , \672 , RIae75c68_25);
and \U$4737 ( \5114 , RIae75d58_27, \670 );
nor \U$4738 ( \5115 , \5113 , \5114 );
and \U$4739 ( \5116 , \5115 , \588 );
not \U$4740 ( \5117 , \5115 );
and \U$4741 ( \5118 , \5117 , \587 );
nor \U$4742 ( \5119 , \5116 , \5118 );
xor \U$4743 ( \5120 , \5112 , \5119 );
not \U$4744 ( \5121 , \787 );
and \U$4745 ( \5122 , \883 , RIae755d8_11);
and \U$4746 ( \5123 , RIae754e8_9, \881 );
nor \U$4747 ( \5124 , \5122 , \5123 );
not \U$4748 ( \5125 , \5124 );
or \U$4749 ( \5126 , \5121 , \5125 );
or \U$4750 ( \5127 , \5124 , \789 );
nand \U$4751 ( \5128 , \5126 , \5127 );
and \U$4752 ( \5129 , \5120 , \5128 );
and \U$4753 ( \5130 , \5112 , \5119 );
or \U$4754 ( \5131 , \5129 , \5130 );
xor \U$4755 ( \5132 , \5105 , \5131 );
not \U$4756 ( \5133 , \469 );
and \U$4757 ( \5134 , \514 , RIae75998_19);
and \U$4758 ( \5135 , RIae758a8_17, \512 );
nor \U$4759 ( \5136 , \5134 , \5135 );
not \U$4760 ( \5137 , \5136 );
or \U$4761 ( \5138 , \5133 , \5137 );
or \U$4762 ( \5139 , \5136 , \469 );
nand \U$4763 ( \5140 , \5138 , \5139 );
not \U$4764 ( \5141 , \392 );
and \U$4765 ( \5142 , \384 , RIae78788_117);
and \U$4766 ( \5143 , RIae78698_115, \382 );
nor \U$4767 ( \5144 , \5142 , \5143 );
not \U$4768 ( \5145 , \5144 );
or \U$4769 ( \5146 , \5141 , \5145 );
or \U$4770 ( \5147 , \5144 , \388 );
nand \U$4771 ( \5148 , \5146 , \5147 );
xor \U$4772 ( \5149 , \5140 , \5148 );
not \U$4773 ( \5150 , \400 );
and \U$4774 ( \5151 , \436 , RIae75b78_23);
and \U$4775 ( \5152 , RIae75a88_21, \434 );
nor \U$4776 ( \5153 , \5151 , \5152 );
not \U$4777 ( \5154 , \5153 );
or \U$4778 ( \5155 , \5150 , \5154 );
or \U$4779 ( \5156 , \5153 , \400 );
nand \U$4780 ( \5157 , \5155 , \5156 );
and \U$4781 ( \5158 , \5149 , \5157 );
and \U$4782 ( \5159 , \5140 , \5148 );
or \U$4783 ( \5160 , \5158 , \5159 );
and \U$4784 ( \5161 , \5132 , \5160 );
and \U$4785 ( \5162 , \5105 , \5131 );
or \U$4786 ( \5163 , \5161 , \5162 );
and \U$4787 ( \5164 , \5080 , \5163 );
and \U$4788 ( \5165 , \5058 , \5079 );
or \U$4789 ( \5166 , \5164 , \5165 );
not \U$4790 ( \5167 , \5166 );
or \U$4791 ( \5168 , \4980 , \5167 );
or \U$4792 ( \5169 , \5166 , \4979 );
not \U$4793 ( \5170 , \4835 );
not \U$4794 ( \5171 , \4827 );
or \U$4795 ( \5172 , \5170 , \5171 );
or \U$4796 ( \5173 , \4827 , \4835 );
nand \U$4797 ( \5174 , \5172 , \5173 );
not \U$4798 ( \5175 , \5174 );
not \U$4799 ( \5176 , \4829 );
and \U$4800 ( \5177 , \5175 , \5176 );
and \U$4801 ( \5178 , \5174 , \4829 );
nor \U$4802 ( \5179 , \5177 , \5178 );
not \U$4803 ( \5180 , \4854 );
not \U$4804 ( \5181 , \4860 );
or \U$4805 ( \5182 , \5180 , \5181 );
or \U$4806 ( \5183 , \4854 , \4860 );
nand \U$4807 ( \5184 , \5182 , \5183 );
not \U$4808 ( \5185 , \5184 );
not \U$4809 ( \5186 , \4852 );
and \U$4810 ( \5187 , \5185 , \5186 );
and \U$4811 ( \5188 , \5184 , \4852 );
nor \U$4812 ( \5189 , \5187 , \5188 );
or \U$4813 ( \5190 , \5179 , \5189 );
not \U$4814 ( \5191 , \5189 );
not \U$4815 ( \5192 , \5179 );
or \U$4816 ( \5193 , \5191 , \5192 );
xor \U$4817 ( \5194 , \4795 , \4802 );
xor \U$4818 ( \5195 , \5194 , \4810 );
xor \U$4819 ( \5196 , \4655 , \4662 );
xor \U$4820 ( \5197 , \5196 , \4670 );
and \U$4821 ( \5198 , \5195 , \5197 );
xor \U$4822 ( \5199 , \4712 , \4720 );
xor \U$4823 ( \5200 , \5199 , \4729 );
xor \U$4824 ( \5201 , \4655 , \4662 );
xor \U$4825 ( \5202 , \5201 , \4670 );
and \U$4826 ( \5203 , \5200 , \5202 );
and \U$4827 ( \5204 , \5195 , \5200 );
or \U$4828 ( \5205 , \5198 , \5203 , \5204 );
nand \U$4829 ( \5206 , \5193 , \5205 );
nand \U$4830 ( \5207 , \5190 , \5206 );
nand \U$4831 ( \5208 , \5169 , \5207 );
nand \U$4832 ( \5209 , \5168 , \5208 );
nand \U$4833 ( \5210 , \4974 , \5209 );
nand \U$4834 ( \5211 , \4971 , \5210 );
and \U$4835 ( \5212 , \4953 , \5211 );
and \U$4836 ( \5213 , \4950 , \4952 );
nor \U$4837 ( \5214 , \5212 , \5213 );
nor \U$4838 ( \5215 , \4948 , \5214 );
and \U$4839 ( \5216 , \4945 , \5215 );
xor \U$4840 ( \5217 , \5215 , \4945 );
not \U$4841 ( \5218 , \4947 );
not \U$4842 ( \5219 , \5214 );
and \U$4843 ( \5220 , \5218 , \5219 );
and \U$4844 ( \5221 , \4947 , \5214 );
nor \U$4845 ( \5222 , \5220 , \5221 );
not \U$4846 ( \5223 , \5209 );
not \U$4847 ( \5224 , \4970 );
or \U$4848 ( \5225 , \5223 , \5224 );
or \U$4849 ( \5226 , \4970 , \5209 );
nand \U$4850 ( \5227 , \5225 , \5226 );
not \U$4851 ( \5228 , \5227 );
not \U$4852 ( \5229 , \4959 );
and \U$4853 ( \5230 , \5228 , \5229 );
and \U$4854 ( \5231 , \5227 , \4959 );
nor \U$4855 ( \5232 , \5230 , \5231 );
xnor \U$4856 ( \5233 , \4840 , \4874 );
not \U$4857 ( \5234 , \5233 );
not \U$4858 ( \5235 , \4647 );
and \U$4859 ( \5236 , \5234 , \5235 );
and \U$4860 ( \5237 , \5233 , \4647 );
nor \U$4861 ( \5238 , \5236 , \5237 );
xor \U$4862 ( \5239 , \5232 , \5238 );
xor \U$4863 ( \5240 , \4960 , \4962 );
xor \U$4864 ( \5241 , \5240 , \4967 );
not \U$4865 ( \5242 , \5241 );
xor \U$4866 ( \5243 , \5058 , \5079 );
xor \U$4867 ( \5244 , \5243 , \5163 );
xor \U$4868 ( \5245 , \4976 , \4978 );
and \U$4869 ( \5246 , \5244 , \5245 );
not \U$4870 ( \5247 , \5244 );
not \U$4871 ( \5248 , \5245 );
and \U$4872 ( \5249 , \5247 , \5248 );
not \U$4873 ( \5250 , \5205 );
not \U$4874 ( \5251 , \5179 );
or \U$4875 ( \5252 , \5250 , \5251 );
or \U$4876 ( \5253 , \5179 , \5205 );
nand \U$4877 ( \5254 , \5252 , \5253 );
not \U$4878 ( \5255 , \5254 );
not \U$4879 ( \5256 , \5189 );
and \U$4880 ( \5257 , \5255 , \5256 );
and \U$4881 ( \5258 , \5254 , \5189 );
nor \U$4882 ( \5259 , \5257 , \5258 );
nor \U$4883 ( \5260 , \5249 , \5259 );
nor \U$4884 ( \5261 , \5246 , \5260 );
nand \U$4885 ( \5262 , \5242 , \5261 );
or \U$4886 ( \5263 , \5068 , \5078 );
nand \U$4887 ( \5264 , \5263 , \5079 );
xor \U$4888 ( \5265 , \5005 , \5027 );
xor \U$4889 ( \5266 , \5265 , \5055 );
and \U$4890 ( \5267 , \5264 , \5266 );
xor \U$4891 ( \5268 , \5105 , \5131 );
xor \U$4892 ( \5269 , \5268 , \5160 );
xor \U$4893 ( \5270 , \5005 , \5027 );
xor \U$4894 ( \5271 , \5270 , \5055 );
and \U$4895 ( \5272 , \5269 , \5271 );
and \U$4896 ( \5273 , \5264 , \5269 );
or \U$4897 ( \5274 , \5267 , \5272 , \5273 );
and \U$4898 ( \5275 , \1138 , RIae754e8_9);
and \U$4899 ( \5276 , RIae757b8_15, \1136 );
nor \U$4900 ( \5277 , \5275 , \5276 );
and \U$4901 ( \5278 , \5277 , \1012 );
not \U$4902 ( \5279 , \5277 );
and \U$4903 ( \5280 , \5279 , \1142 );
nor \U$4904 ( \5281 , \5278 , \5280 );
and \U$4905 ( \5282 , \1376 , RIae756c8_13);
and \U$4906 ( \5283 , RIae75218_3, \1374 );
nor \U$4907 ( \5284 , \5282 , \5283 );
and \U$4908 ( \5285 , \5284 , \1380 );
not \U$4909 ( \5286 , \5284 );
and \U$4910 ( \5287 , \5286 , \1261 );
nor \U$4911 ( \5288 , \5285 , \5287 );
xor \U$4912 ( \5289 , \5281 , \5288 );
and \U$4913 ( \5290 , \1593 , RIae75128_1);
and \U$4914 ( \5291 , RIae75308_5, \1591 );
nor \U$4915 ( \5292 , \5290 , \5291 );
and \U$4916 ( \5293 , \5292 , \1498 );
not \U$4917 ( \5294 , \5292 );
and \U$4918 ( \5295 , \5294 , \1488 );
nor \U$4919 ( \5296 , \5293 , \5295 );
and \U$4920 ( \5297 , \5289 , \5296 );
and \U$4921 ( \5298 , \5281 , \5288 );
or \U$4922 ( \5299 , \5297 , \5298 );
and \U$4923 ( \5300 , \436 , RIae78698_115);
and \U$4924 ( \5301 , RIae75b78_23, \434 );
nor \U$4925 ( \5302 , \5300 , \5301 );
not \U$4926 ( \5303 , \5302 );
not \U$4927 ( \5304 , \400 );
and \U$4928 ( \5305 , \5303 , \5304 );
and \U$4929 ( \5306 , \5302 , \402 );
nor \U$4930 ( \5307 , \5305 , \5306 );
and \U$4931 ( \5308 , \514 , RIae75a88_21);
and \U$4932 ( \5309 , RIae75998_19, \512 );
nor \U$4933 ( \5310 , \5308 , \5309 );
not \U$4934 ( \5311 , \5310 );
not \U$4935 ( \5312 , \469 );
and \U$4936 ( \5313 , \5311 , \5312 );
and \U$4937 ( \5314 , \5310 , \469 );
nor \U$4938 ( \5315 , \5313 , \5314 );
xor \U$4939 ( \5316 , \5307 , \5315 );
and \U$4940 ( \5317 , \384 , RIae78878_119);
and \U$4941 ( \5318 , RIae78788_117, \382 );
nor \U$4942 ( \5319 , \5317 , \5318 );
not \U$4943 ( \5320 , \5319 );
not \U$4944 ( \5321 , \392 );
and \U$4945 ( \5322 , \5320 , \5321 );
and \U$4946 ( \5323 , \5319 , \392 );
nor \U$4947 ( \5324 , \5322 , \5323 );
and \U$4948 ( \5325 , \5316 , \5324 );
and \U$4949 ( \5326 , \5307 , \5315 );
nor \U$4950 ( \5327 , \5325 , \5326 );
xor \U$4951 ( \5328 , \5299 , \5327 );
and \U$4952 ( \5329 , \558 , RIae758a8_17);
and \U$4953 ( \5330 , RIae75f38_31, \556 );
nor \U$4954 ( \5331 , \5329 , \5330 );
and \U$4955 ( \5332 , \5331 , \504 );
not \U$4956 ( \5333 , \5331 );
and \U$4957 ( \5334 , \5333 , \562 );
nor \U$4958 ( \5335 , \5332 , \5334 );
and \U$4959 ( \5336 , \672 , RIae75e48_29);
and \U$4960 ( \5337 , RIae75c68_25, \670 );
nor \U$4961 ( \5338 , \5336 , \5337 );
and \U$4962 ( \5339 , \5338 , \588 );
not \U$4963 ( \5340 , \5338 );
and \U$4964 ( \5341 , \5340 , \587 );
nor \U$4965 ( \5342 , \5339 , \5341 );
xor \U$4966 ( \5343 , \5335 , \5342 );
not \U$4967 ( \5344 , \787 );
and \U$4968 ( \5345 , \883 , RIae75d58_27);
and \U$4969 ( \5346 , RIae755d8_11, \881 );
nor \U$4970 ( \5347 , \5345 , \5346 );
not \U$4971 ( \5348 , \5347 );
or \U$4972 ( \5349 , \5344 , \5348 );
or \U$4973 ( \5350 , \5347 , \787 );
nand \U$4974 ( \5351 , \5349 , \5350 );
and \U$4975 ( \5352 , \5343 , \5351 );
and \U$4976 ( \5353 , \5335 , \5342 );
or \U$4977 ( \5354 , \5352 , \5353 );
and \U$4978 ( \5355 , \5328 , \5354 );
and \U$4979 ( \5356 , \5299 , \5327 );
or \U$4980 ( \5357 , \5355 , \5356 );
not \U$4981 ( \5358 , \3089 );
and \U$4982 ( \5359 , \2783 , RIae76028_33);
and \U$4983 ( \5360 , RIae762f8_39, \2781 );
nor \U$4984 ( \5361 , \5359 , \5360 );
not \U$4985 ( \5362 , \5361 );
or \U$4986 ( \5363 , \5358 , \5362 );
or \U$4987 ( \5364 , \5361 , \2789 );
nand \U$4988 ( \5365 , \5363 , \5364 );
not \U$4989 ( \5366 , \3218 );
and \U$4990 ( \5367 , \3214 , RIae76208_37);
and \U$4991 ( \5368 , RIae76a78_55, \3212 );
nor \U$4992 ( \5369 , \5367 , \5368 );
not \U$4993 ( \5370 , \5369 );
or \U$4994 ( \5371 , \5366 , \5370 );
or \U$4995 ( \5372 , \5369 , \3218 );
nand \U$4996 ( \5373 , \5371 , \5372 );
xor \U$4997 ( \5374 , \5365 , \5373 );
and \U$4998 ( \5375 , \3730 , RIae76988_53);
and \U$4999 ( \5376 , RIae767a8_49, \3728 );
nor \U$5000 ( \5377 , \5375 , \5376 );
and \U$5001 ( \5378 , \5377 , \3732 );
not \U$5002 ( \5379 , \5377 );
and \U$5003 ( \5380 , \5379 , \3422 );
nor \U$5004 ( \5381 , \5378 , \5380 );
and \U$5005 ( \5382 , \5374 , \5381 );
and \U$5006 ( \5383 , \5365 , \5373 );
or \U$5007 ( \5384 , \5382 , \5383 );
and \U$5008 ( \5385 , \4247 , RIae76898_51);
and \U$5009 ( \5386 , RIae76b68_57, \4245 );
nor \U$5010 ( \5387 , \5385 , \5386 );
and \U$5011 ( \5388 , \5387 , \3989 );
not \U$5012 ( \5389 , \5387 );
and \U$5013 ( \5390 , \5389 , \4251 );
nor \U$5014 ( \5391 , \5388 , \5390 );
and \U$5015 ( \5392 , RIae79ca0_162, RIae79e08_165);
not \U$5016 ( \5393 , RIae79e08_165);
nor \U$5017 ( \5394 , \5393 , RIae79d90_164);
not \U$5018 ( \5395 , RIae79d90_164);
nor \U$5019 ( \5396 , \5395 , RIae79e08_165);
or \U$5020 ( \5397 , \5394 , \5396 );
nor \U$5021 ( \5398 , RIae79ca0_162, RIae79e08_165);
nor \U$5022 ( \5399 , \5392 , \5397 , \5398 );
nand \U$5023 ( \5400 , RIae78da0_130, \5399 );
and \U$5024 ( \5401 , \5400 , \5016 );
not \U$5025 ( \5402 , \5400 );
not \U$5026 ( \5403 , \5016 );
and \U$5027 ( \5404 , \5402 , \5403 );
nor \U$5028 ( \5405 , \5401 , \5404 );
xor \U$5029 ( \5406 , \5391 , \5405 );
and \U$5030 ( \5407 , \4688 , RIae78a58_123);
and \U$5031 ( \5408 , RIae78cb0_128, \4686 );
nor \U$5032 ( \5409 , \5407 , \5408 );
and \U$5033 ( \5410 , \5409 , \4481 );
not \U$5034 ( \5411 , \5409 );
and \U$5035 ( \5412 , \5411 , \4482 );
nor \U$5036 ( \5413 , \5410 , \5412 );
and \U$5037 ( \5414 , \5406 , \5413 );
and \U$5038 ( \5415 , \5391 , \5405 );
or \U$5039 ( \5416 , \5414 , \5415 );
xor \U$5040 ( \5417 , \5384 , \5416 );
and \U$5041 ( \5418 , \2607 , RIae765c8_45);
and \U$5042 ( \5419 , RIae76118_35, \2605 );
nor \U$5043 ( \5420 , \5418 , \5419 );
and \U$5044 ( \5421 , \5420 , \2611 );
not \U$5045 ( \5422 , \5420 );
and \U$5046 ( \5423 , \5422 , \2397 );
nor \U$5047 ( \5424 , \5421 , \5423 );
and \U$5048 ( \5425 , \1939 , RIae753f8_7);
and \U$5049 ( \5426 , RIae763e8_41, \1937 );
nor \U$5050 ( \5427 , \5425 , \5426 );
and \U$5051 ( \5428 , \5427 , \1735 );
not \U$5052 ( \5429 , \5427 );
and \U$5053 ( \5430 , \5429 , \1734 );
nor \U$5054 ( \5431 , \5428 , \5430 );
xor \U$5055 ( \5432 , \5424 , \5431 );
and \U$5056 ( \5433 , \2224 , RIae764d8_43);
and \U$5057 ( \5434 , RIae766b8_47, \2222 );
nor \U$5058 ( \5435 , \5433 , \5434 );
and \U$5059 ( \5436 , \5435 , \2061 );
not \U$5060 ( \5437 , \5435 );
and \U$5061 ( \5438 , \5437 , \2060 );
nor \U$5062 ( \5439 , \5436 , \5438 );
and \U$5063 ( \5440 , \5432 , \5439 );
and \U$5064 ( \5441 , \5424 , \5431 );
or \U$5065 ( \5442 , \5440 , \5441 );
and \U$5066 ( \5443 , \5417 , \5442 );
and \U$5067 ( \5444 , \5384 , \5416 );
or \U$5068 ( \5445 , \5443 , \5444 );
xor \U$5069 ( \5446 , \5357 , \5445 );
not \U$5070 ( \5447 , RIae78878_119);
nor \U$5071 ( \5448 , \5447 , \491 );
xor \U$5072 ( \5449 , \5112 , \5119 );
xor \U$5073 ( \5450 , \5449 , \5128 );
and \U$5074 ( \5451 , \5448 , \5450 );
xor \U$5075 ( \5452 , \5140 , \5148 );
xor \U$5076 ( \5453 , \5452 , \5157 );
xor \U$5077 ( \5454 , \5112 , \5119 );
xor \U$5078 ( \5455 , \5454 , \5128 );
and \U$5079 ( \5456 , \5453 , \5455 );
and \U$5080 ( \5457 , \5448 , \5453 );
or \U$5081 ( \5458 , \5451 , \5456 , \5457 );
and \U$5082 ( \5459 , \5446 , \5458 );
and \U$5083 ( \5460 , \5357 , \5445 );
or \U$5084 ( \5461 , \5459 , \5460 );
xor \U$5085 ( \5462 , \5274 , \5461 );
xor \U$5086 ( \5463 , \5087 , \5094 );
xor \U$5087 ( \5464 , \5463 , \5102 );
xor \U$5088 ( \5465 , \5035 , \5043 );
xor \U$5089 ( \5466 , \5465 , \5052 );
and \U$5090 ( \5467 , \5464 , \5466 );
xor \U$5091 ( \5468 , \4987 , \4994 );
xor \U$5092 ( \5469 , \5468 , \5002 );
xor \U$5093 ( \5470 , \5035 , \5043 );
xor \U$5094 ( \5471 , \5470 , \5052 );
and \U$5095 ( \5472 , \5469 , \5471 );
and \U$5096 ( \5473 , \5464 , \5469 );
or \U$5097 ( \5474 , \5467 , \5472 , \5473 );
xor \U$5098 ( \5475 , \4680 , \4693 );
xor \U$5099 ( \5476 , \5475 , \4701 );
xor \U$5100 ( \5477 , \5474 , \5476 );
xor \U$5101 ( \5478 , \4655 , \4662 );
xor \U$5102 ( \5479 , \5478 , \4670 );
xor \U$5103 ( \5480 , \5195 , \5200 );
xor \U$5104 ( \5481 , \5479 , \5480 );
and \U$5105 ( \5482 , \5477 , \5481 );
and \U$5106 ( \5483 , \5474 , \5476 );
or \U$5107 ( \5484 , \5482 , \5483 );
and \U$5108 ( \5485 , \5462 , \5484 );
and \U$5109 ( \5486 , \5274 , \5461 );
or \U$5110 ( \5487 , \5485 , \5486 );
and \U$5111 ( \5488 , \5262 , \5487 );
not \U$5112 ( \5489 , \5261 );
and \U$5113 ( \5490 , \5489 , \5241 );
nor \U$5114 ( \5491 , \5488 , \5490 );
and \U$5115 ( \5492 , \5239 , \5491 );
and \U$5116 ( \5493 , \5232 , \5238 );
or \U$5117 ( \5494 , \5492 , \5493 );
not \U$5118 ( \5495 , \5494 );
xor \U$5119 ( \5496 , \4950 , \4952 );
xor \U$5120 ( \5497 , \5496 , \5211 );
nand \U$5121 ( \5498 , \5495 , \5497 );
or \U$5122 ( \5499 , \5222 , \5498 );
xnor \U$5123 ( \5500 , \5222 , \5498 );
not \U$5124 ( \5501 , \5494 );
not \U$5125 ( \5502 , \5497 );
or \U$5126 ( \5503 , \5501 , \5502 );
or \U$5127 ( \5504 , \5497 , \5494 );
nand \U$5128 ( \5505 , \5503 , \5504 );
not \U$5129 ( \5506 , \5241 );
not \U$5130 ( \5507 , \5261 );
not \U$5131 ( \5508 , \5487 );
and \U$5132 ( \5509 , \5507 , \5508 );
and \U$5133 ( \5510 , \5261 , \5487 );
nor \U$5134 ( \5511 , \5509 , \5510 );
not \U$5135 ( \5512 , \5511 );
or \U$5136 ( \5513 , \5506 , \5512 );
or \U$5137 ( \5514 , \5511 , \5241 );
nand \U$5138 ( \5515 , \5513 , \5514 );
not \U$5139 ( \5516 , \5515 );
xnor \U$5140 ( \5517 , \5166 , \5207 );
not \U$5141 ( \5518 , \5517 );
not \U$5142 ( \5519 , \4979 );
and \U$5143 ( \5520 , \5518 , \5519 );
and \U$5144 ( \5521 , \5517 , \4979 );
nor \U$5145 ( \5522 , \5520 , \5521 );
or \U$5146 ( \5523 , \5516 , \5522 );
not \U$5147 ( \5524 , \5522 );
not \U$5148 ( \5525 , \5516 );
or \U$5149 ( \5526 , \5524 , \5525 );
xor \U$5150 ( \5527 , \5357 , \5445 );
xor \U$5151 ( \5528 , \5527 , \5458 );
xor \U$5152 ( \5529 , \5474 , \5476 );
xor \U$5153 ( \5530 , \5529 , \5481 );
and \U$5154 ( \5531 , \5528 , \5530 );
xor \U$5155 ( \5532 , \5005 , \5027 );
xor \U$5156 ( \5533 , \5532 , \5055 );
xor \U$5157 ( \5534 , \5264 , \5269 );
xor \U$5158 ( \5535 , \5533 , \5534 );
xor \U$5159 ( \5536 , \5474 , \5476 );
xor \U$5160 ( \5537 , \5536 , \5481 );
and \U$5161 ( \5538 , \5535 , \5537 );
and \U$5162 ( \5539 , \5528 , \5535 );
or \U$5163 ( \5540 , \5531 , \5538 , \5539 );
xor \U$5164 ( \5541 , \5384 , \5416 );
xor \U$5165 ( \5542 , \5541 , \5442 );
xor \U$5166 ( \5543 , \5299 , \5327 );
xor \U$5167 ( \5544 , \5543 , \5354 );
and \U$5168 ( \5545 , \5542 , \5544 );
xor \U$5169 ( \5546 , \5112 , \5119 );
xor \U$5170 ( \5547 , \5546 , \5128 );
xor \U$5171 ( \5548 , \5448 , \5453 );
xor \U$5172 ( \5549 , \5547 , \5548 );
xor \U$5173 ( \5550 , \5299 , \5327 );
xor \U$5174 ( \5551 , \5550 , \5354 );
and \U$5175 ( \5552 , \5549 , \5551 );
and \U$5176 ( \5553 , \5542 , \5549 );
or \U$5177 ( \5554 , \5545 , \5552 , \5553 );
and \U$5178 ( \5555 , \2224 , RIae763e8_41);
and \U$5179 ( \5556 , RIae764d8_43, \2222 );
nor \U$5180 ( \5557 , \5555 , \5556 );
and \U$5181 ( \5558 , \5557 , \2061 );
not \U$5182 ( \5559 , \5557 );
and \U$5183 ( \5560 , \5559 , \2060 );
nor \U$5184 ( \5561 , \5558 , \5560 );
and \U$5185 ( \5562 , \2607 , RIae766b8_47);
and \U$5186 ( \5563 , RIae765c8_45, \2605 );
nor \U$5187 ( \5564 , \5562 , \5563 );
and \U$5188 ( \5565 , \5564 , \2611 );
not \U$5189 ( \5566 , \5564 );
and \U$5190 ( \5567 , \5566 , \2397 );
nor \U$5191 ( \5568 , \5565 , \5567 );
xor \U$5192 ( \5569 , \5561 , \5568 );
not \U$5193 ( \5570 , \2789 );
and \U$5194 ( \5571 , \2783 , RIae76118_35);
and \U$5195 ( \5572 , RIae76028_33, \2781 );
nor \U$5196 ( \5573 , \5571 , \5572 );
not \U$5197 ( \5574 , \5573 );
or \U$5198 ( \5575 , \5570 , \5574 );
or \U$5199 ( \5576 , \5573 , \3089 );
nand \U$5200 ( \5577 , \5575 , \5576 );
and \U$5201 ( \5578 , \5569 , \5577 );
and \U$5202 ( \5579 , \5561 , \5568 );
or \U$5203 ( \5580 , \5578 , \5579 );
and \U$5204 ( \5581 , \4688 , RIae76b68_57);
and \U$5205 ( \5582 , RIae78a58_123, \4686 );
nor \U$5206 ( \5583 , \5581 , \5582 );
and \U$5207 ( \5584 , \5583 , \4481 );
not \U$5208 ( \5585 , \5583 );
and \U$5209 ( \5586 , \5585 , \4482 );
nor \U$5210 ( \5587 , \5584 , \5586 );
nand \U$5211 ( \5588 , RIae79ef8_167, RIae79e80_166);
and \U$5212 ( \5589 , \5588 , RIae79d90_164);
not \U$5213 ( \5590 , \5589 );
xor \U$5214 ( \5591 , \5587 , \5590 );
and \U$5215 ( \5592 , \5399 , RIae78cb0_128);
and \U$5216 ( \5593 , RIae78da0_130, \5397 );
nor \U$5217 ( \5594 , \5592 , \5593 );
and \U$5218 ( \5595 , \5594 , \5016 );
not \U$5219 ( \5596 , \5594 );
and \U$5220 ( \5597 , \5596 , \5403 );
nor \U$5221 ( \5598 , \5595 , \5597 );
and \U$5222 ( \5599 , \5591 , \5598 );
and \U$5223 ( \5600 , \5587 , \5590 );
or \U$5224 ( \5601 , \5599 , \5600 );
xor \U$5225 ( \5602 , \5580 , \5601 );
and \U$5226 ( \5603 , \3730 , RIae76a78_55);
and \U$5227 ( \5604 , RIae76988_53, \3728 );
nor \U$5228 ( \5605 , \5603 , \5604 );
and \U$5229 ( \5606 , \5605 , \3732 );
not \U$5230 ( \5607 , \5605 );
and \U$5231 ( \5608 , \5607 , \3422 );
nor \U$5232 ( \5609 , \5606 , \5608 );
not \U$5233 ( \5610 , \3218 );
and \U$5234 ( \5611 , \3214 , RIae762f8_39);
and \U$5235 ( \5612 , RIae76208_37, \3212 );
nor \U$5236 ( \5613 , \5611 , \5612 );
not \U$5237 ( \5614 , \5613 );
or \U$5238 ( \5615 , \5610 , \5614 );
or \U$5239 ( \5616 , \5613 , \2774 );
nand \U$5240 ( \5617 , \5615 , \5616 );
xor \U$5241 ( \5618 , \5609 , \5617 );
and \U$5242 ( \5619 , \4247 , RIae767a8_49);
and \U$5243 ( \5620 , RIae76898_51, \4245 );
nor \U$5244 ( \5621 , \5619 , \5620 );
and \U$5245 ( \5622 , \5621 , \3989 );
not \U$5246 ( \5623 , \5621 );
and \U$5247 ( \5624 , \5623 , \4251 );
nor \U$5248 ( \5625 , \5622 , \5624 );
and \U$5249 ( \5626 , \5618 , \5625 );
and \U$5250 ( \5627 , \5609 , \5617 );
or \U$5251 ( \5628 , \5626 , \5627 );
and \U$5252 ( \5629 , \5602 , \5628 );
and \U$5253 ( \5630 , \5580 , \5601 );
or \U$5254 ( \5631 , \5629 , \5630 );
nand \U$5255 ( \5632 , RIae78968_121, RIae78b48_125);
xor \U$5256 ( \5633 , \5307 , \5315 );
xor \U$5257 ( \5634 , \5633 , \5324 );
nand \U$5258 ( \5635 , \5632 , \5634 );
xor \U$5259 ( \5636 , \5631 , \5635 );
and \U$5260 ( \5637 , \1138 , RIae755d8_11);
and \U$5261 ( \5638 , RIae754e8_9, \1136 );
nor \U$5262 ( \5639 , \5637 , \5638 );
and \U$5263 ( \5640 , \5639 , \1012 );
not \U$5264 ( \5641 , \5639 );
and \U$5265 ( \5642 , \5641 , \1142 );
nor \U$5266 ( \5643 , \5640 , \5642 );
and \U$5267 ( \5644 , \672 , RIae75f38_31);
and \U$5268 ( \5645 , RIae75e48_29, \670 );
nor \U$5269 ( \5646 , \5644 , \5645 );
and \U$5270 ( \5647 , \5646 , \588 );
not \U$5271 ( \5648 , \5646 );
and \U$5272 ( \5649 , \5648 , \587 );
nor \U$5273 ( \5650 , \5647 , \5649 );
xor \U$5274 ( \5651 , \5643 , \5650 );
not \U$5275 ( \5652 , \787 );
and \U$5276 ( \5653 , \883 , RIae75c68_25);
and \U$5277 ( \5654 , RIae75d58_27, \881 );
nor \U$5278 ( \5655 , \5653 , \5654 );
not \U$5279 ( \5656 , \5655 );
or \U$5280 ( \5657 , \5652 , \5656 );
or \U$5281 ( \5658 , \5655 , \789 );
nand \U$5282 ( \5659 , \5657 , \5658 );
and \U$5283 ( \5660 , \5651 , \5659 );
and \U$5284 ( \5661 , \5643 , \5650 );
or \U$5285 ( \5662 , \5660 , \5661 );
not \U$5286 ( \5663 , \400 );
and \U$5287 ( \5664 , \436 , RIae78788_117);
and \U$5288 ( \5665 , RIae78698_115, \434 );
nor \U$5289 ( \5666 , \5664 , \5665 );
not \U$5290 ( \5667 , \5666 );
or \U$5291 ( \5668 , \5663 , \5667 );
or \U$5292 ( \5669 , \5666 , \400 );
nand \U$5293 ( \5670 , \5668 , \5669 );
not \U$5294 ( \5671 , \471 );
and \U$5295 ( \5672 , \514 , RIae75b78_23);
and \U$5296 ( \5673 , RIae75a88_21, \512 );
nor \U$5297 ( \5674 , \5672 , \5673 );
not \U$5298 ( \5675 , \5674 );
or \U$5299 ( \5676 , \5671 , \5675 );
or \U$5300 ( \5677 , \5674 , \469 );
nand \U$5301 ( \5678 , \5676 , \5677 );
xor \U$5302 ( \5679 , \5670 , \5678 );
and \U$5303 ( \5680 , \558 , RIae75998_19);
and \U$5304 ( \5681 , RIae758a8_17, \556 );
nor \U$5305 ( \5682 , \5680 , \5681 );
and \U$5306 ( \5683 , \5682 , \504 );
not \U$5307 ( \5684 , \5682 );
and \U$5308 ( \5685 , \5684 , \562 );
nor \U$5309 ( \5686 , \5683 , \5685 );
and \U$5310 ( \5687 , \5679 , \5686 );
and \U$5311 ( \5688 , \5670 , \5678 );
or \U$5312 ( \5689 , \5687 , \5688 );
xor \U$5313 ( \5690 , \5662 , \5689 );
and \U$5314 ( \5691 , \1376 , RIae757b8_15);
and \U$5315 ( \5692 , RIae756c8_13, \1374 );
nor \U$5316 ( \5693 , \5691 , \5692 );
and \U$5317 ( \5694 , \5693 , \1380 );
not \U$5318 ( \5695 , \5693 );
and \U$5319 ( \5696 , \5695 , \1261 );
nor \U$5320 ( \5697 , \5694 , \5696 );
and \U$5321 ( \5698 , \1593 , RIae75218_3);
and \U$5322 ( \5699 , RIae75128_1, \1591 );
nor \U$5323 ( \5700 , \5698 , \5699 );
and \U$5324 ( \5701 , \5700 , \1498 );
not \U$5325 ( \5702 , \5700 );
and \U$5326 ( \5703 , \5702 , \1488 );
nor \U$5327 ( \5704 , \5701 , \5703 );
xor \U$5328 ( \5705 , \5697 , \5704 );
and \U$5329 ( \5706 , \1939 , RIae75308_5);
and \U$5330 ( \5707 , RIae753f8_7, \1937 );
nor \U$5331 ( \5708 , \5706 , \5707 );
and \U$5332 ( \5709 , \5708 , \1735 );
not \U$5333 ( \5710 , \5708 );
and \U$5334 ( \5711 , \5710 , \1734 );
nor \U$5335 ( \5712 , \5709 , \5711 );
and \U$5336 ( \5713 , \5705 , \5712 );
and \U$5337 ( \5714 , \5697 , \5704 );
or \U$5338 ( \5715 , \5713 , \5714 );
and \U$5339 ( \5716 , \5690 , \5715 );
and \U$5340 ( \5717 , \5662 , \5689 );
or \U$5341 ( \5718 , \5716 , \5717 );
and \U$5342 ( \5719 , \5636 , \5718 );
and \U$5343 ( \5720 , \5631 , \5635 );
or \U$5344 ( \5721 , \5719 , \5720 );
xor \U$5345 ( \5722 , \5554 , \5721 );
xor \U$5346 ( \5723 , \5281 , \5288 );
xor \U$5347 ( \5724 , \5723 , \5296 );
xor \U$5348 ( \5725 , \5335 , \5342 );
xor \U$5349 ( \5726 , \5725 , \5351 );
and \U$5350 ( \5727 , \5724 , \5726 );
xor \U$5351 ( \5728 , \5424 , \5431 );
xor \U$5352 ( \5729 , \5728 , \5439 );
xor \U$5353 ( \5730 , \5335 , \5342 );
xor \U$5354 ( \5731 , \5730 , \5351 );
and \U$5355 ( \5732 , \5729 , \5731 );
and \U$5356 ( \5733 , \5724 , \5729 );
or \U$5357 ( \5734 , \5727 , \5732 , \5733 );
xor \U$5358 ( \5735 , \5012 , \5016 );
xor \U$5359 ( \5736 , \5735 , \5024 );
xor \U$5360 ( \5737 , \5734 , \5736 );
xor \U$5361 ( \5738 , \5035 , \5043 );
xor \U$5362 ( \5739 , \5738 , \5052 );
xor \U$5363 ( \5740 , \5464 , \5469 );
xor \U$5364 ( \5741 , \5739 , \5740 );
and \U$5365 ( \5742 , \5737 , \5741 );
and \U$5366 ( \5743 , \5734 , \5736 );
or \U$5367 ( \5744 , \5742 , \5743 );
and \U$5368 ( \5745 , \5722 , \5744 );
and \U$5369 ( \5746 , \5554 , \5721 );
or \U$5370 ( \5747 , \5745 , \5746 );
xor \U$5371 ( \5748 , \5540 , \5747 );
not \U$5372 ( \5749 , \5245 );
not \U$5373 ( \5750 , \5259 );
not \U$5374 ( \5751 , \5244 );
and \U$5375 ( \5752 , \5750 , \5751 );
and \U$5376 ( \5753 , \5259 , \5244 );
nor \U$5377 ( \5754 , \5752 , \5753 );
not \U$5378 ( \5755 , \5754 );
or \U$5379 ( \5756 , \5749 , \5755 );
or \U$5380 ( \5757 , \5754 , \5245 );
nand \U$5381 ( \5758 , \5756 , \5757 );
and \U$5382 ( \5759 , \5748 , \5758 );
and \U$5383 ( \5760 , \5540 , \5747 );
or \U$5384 ( \5761 , \5759 , \5760 );
nand \U$5385 ( \5762 , \5526 , \5761 );
nand \U$5386 ( \5763 , \5523 , \5762 );
not \U$5387 ( \5764 , \5763 );
xor \U$5388 ( \5765 , \5232 , \5238 );
xor \U$5389 ( \5766 , \5765 , \5491 );
nor \U$5390 ( \5767 , \5764 , \5766 );
and \U$5391 ( \5768 , \5505 , \5767 );
xor \U$5392 ( \5769 , \5767 , \5505 );
not \U$5393 ( \5770 , \5766 );
not \U$5394 ( \5771 , \5763 );
and \U$5395 ( \5772 , \5770 , \5771 );
and \U$5396 ( \5773 , \5766 , \5763 );
nor \U$5397 ( \5774 , \5772 , \5773 );
not \U$5398 ( \5775 , \5761 );
not \U$5399 ( \5776 , \5522 );
and \U$5400 ( \5777 , \5775 , \5776 );
and \U$5401 ( \5778 , \5761 , \5522 );
nor \U$5402 ( \5779 , \5777 , \5778 );
not \U$5403 ( \5780 , \5779 );
not \U$5404 ( \5781 , \5515 );
and \U$5405 ( \5782 , \5780 , \5781 );
and \U$5406 ( \5783 , \5779 , \5515 );
nor \U$5407 ( \5784 , \5782 , \5783 );
not \U$5408 ( \5785 , \5784 );
xor \U$5409 ( \5786 , \5631 , \5635 );
xor \U$5410 ( \5787 , \5786 , \5718 );
xor \U$5411 ( \5788 , \5734 , \5736 );
xor \U$5412 ( \5789 , \5788 , \5741 );
and \U$5413 ( \5790 , \5787 , \5789 );
xor \U$5414 ( \5791 , \5299 , \5327 );
xor \U$5415 ( \5792 , \5791 , \5354 );
xor \U$5416 ( \5793 , \5542 , \5549 );
xor \U$5417 ( \5794 , \5792 , \5793 );
xor \U$5418 ( \5795 , \5734 , \5736 );
xor \U$5419 ( \5796 , \5795 , \5741 );
and \U$5420 ( \5797 , \5794 , \5796 );
and \U$5421 ( \5798 , \5787 , \5794 );
or \U$5422 ( \5799 , \5790 , \5797 , \5798 );
xor \U$5423 ( \5800 , \5587 , \5590 );
xor \U$5424 ( \5801 , \5800 , \5598 );
xor \U$5425 ( \5802 , \5609 , \5617 );
xor \U$5426 ( \5803 , \5802 , \5625 );
and \U$5427 ( \5804 , \5801 , \5803 );
xor \U$5428 ( \5805 , \5561 , \5568 );
xor \U$5429 ( \5806 , \5805 , \5577 );
xor \U$5430 ( \5807 , \5609 , \5617 );
xor \U$5431 ( \5808 , \5807 , \5625 );
and \U$5432 ( \5809 , \5806 , \5808 );
and \U$5433 ( \5810 , \5801 , \5806 );
or \U$5434 ( \5811 , \5804 , \5809 , \5810 );
xor \U$5435 ( \5812 , \5365 , \5373 );
xor \U$5436 ( \5813 , \5812 , \5381 );
xor \U$5437 ( \5814 , \5811 , \5813 );
xor \U$5438 ( \5815 , \5643 , \5650 );
xor \U$5439 ( \5816 , \5815 , \5659 );
xor \U$5440 ( \5817 , \5670 , \5678 );
xor \U$5441 ( \5818 , \5817 , \5686 );
and \U$5442 ( \5819 , \5816 , \5818 );
xor \U$5443 ( \5820 , \5697 , \5704 );
xor \U$5444 ( \5821 , \5820 , \5712 );
xor \U$5445 ( \5822 , \5670 , \5678 );
xor \U$5446 ( \5823 , \5822 , \5686 );
and \U$5447 ( \5824 , \5821 , \5823 );
and \U$5448 ( \5825 , \5816 , \5821 );
or \U$5449 ( \5826 , \5819 , \5824 , \5825 );
and \U$5450 ( \5827 , \5814 , \5826 );
and \U$5451 ( \5828 , \5811 , \5813 );
or \U$5452 ( \5829 , \5827 , \5828 );
and \U$5453 ( \5830 , \4247 , RIae76988_53);
and \U$5454 ( \5831 , RIae767a8_49, \4245 );
nor \U$5455 ( \5832 , \5830 , \5831 );
and \U$5456 ( \5833 , \5832 , \3989 );
not \U$5457 ( \5834 , \5832 );
and \U$5458 ( \5835 , \5834 , \4251 );
nor \U$5459 ( \5836 , \5833 , \5835 );
not \U$5460 ( \5837 , \3218 );
and \U$5461 ( \5838 , \3214 , RIae76028_33);
and \U$5462 ( \5839 , RIae762f8_39, \3212 );
nor \U$5463 ( \5840 , \5838 , \5839 );
not \U$5464 ( \5841 , \5840 );
or \U$5465 ( \5842 , \5837 , \5841 );
or \U$5466 ( \5843 , \5840 , \2774 );
nand \U$5467 ( \5844 , \5842 , \5843 );
xor \U$5468 ( \5845 , \5836 , \5844 );
and \U$5469 ( \5846 , \3730 , RIae76208_37);
and \U$5470 ( \5847 , RIae76a78_55, \3728 );
nor \U$5471 ( \5848 , \5846 , \5847 );
and \U$5472 ( \5849 , \5848 , \3732 );
not \U$5473 ( \5850 , \5848 );
and \U$5474 ( \5851 , \5850 , \3422 );
nor \U$5475 ( \5852 , \5849 , \5851 );
and \U$5476 ( \5853 , \5845 , \5852 );
and \U$5477 ( \5854 , \5836 , \5844 );
or \U$5478 ( \5855 , \5853 , \5854 );
and \U$5479 ( \5856 , \2224 , RIae753f8_7);
and \U$5480 ( \5857 , RIae763e8_41, \2222 );
nor \U$5481 ( \5858 , \5856 , \5857 );
and \U$5482 ( \5859 , \5858 , \2061 );
not \U$5483 ( \5860 , \5858 );
and \U$5484 ( \5861 , \5860 , \2060 );
nor \U$5485 ( \5862 , \5859 , \5861 );
and \U$5486 ( \5863 , \2607 , RIae764d8_43);
and \U$5487 ( \5864 , RIae766b8_47, \2605 );
nor \U$5488 ( \5865 , \5863 , \5864 );
and \U$5489 ( \5866 , \5865 , \2611 );
not \U$5490 ( \5867 , \5865 );
and \U$5491 ( \5868 , \5867 , \2397 );
nor \U$5492 ( \5869 , \5866 , \5868 );
xor \U$5493 ( \5870 , \5862 , \5869 );
not \U$5494 ( \5871 , \2789 );
and \U$5495 ( \5872 , \2783 , RIae765c8_45);
and \U$5496 ( \5873 , RIae76118_35, \2781 );
nor \U$5497 ( \5874 , \5872 , \5873 );
not \U$5498 ( \5875 , \5874 );
or \U$5499 ( \5876 , \5871 , \5875 );
or \U$5500 ( \5877 , \5874 , \2789 );
nand \U$5501 ( \5878 , \5876 , \5877 );
and \U$5502 ( \5879 , \5870 , \5878 );
and \U$5503 ( \5880 , \5862 , \5869 );
or \U$5504 ( \5881 , \5879 , \5880 );
xor \U$5505 ( \5882 , \5855 , \5881 );
and \U$5506 ( \5883 , \4688 , RIae76898_51);
and \U$5507 ( \5884 , RIae76b68_57, \4686 );
nor \U$5508 ( \5885 , \5883 , \5884 );
and \U$5509 ( \5886 , \5885 , \4481 );
not \U$5510 ( \5887 , \5885 );
and \U$5511 ( \5888 , \5887 , \4482 );
nor \U$5512 ( \5889 , \5886 , \5888 );
and \U$5513 ( \5890 , RIae79d90_164, RIae79e80_166);
not \U$5514 ( \5891 , RIae79ef8_167);
and \U$5515 ( \5892 , \5891 , RIae79e80_166);
nor \U$5516 ( \5893 , \5891 , RIae79e80_166);
or \U$5517 ( \5894 , \5892 , \5893 );
nor \U$5518 ( \5895 , RIae79d90_164, RIae79e80_166);
nor \U$5519 ( \5896 , \5890 , \5894 , \5895 );
nand \U$5520 ( \5897 , RIae78da0_130, \5896 );
and \U$5521 ( \5898 , \5897 , \5590 );
not \U$5522 ( \5899 , \5897 );
and \U$5523 ( \5900 , \5899 , \5589 );
nor \U$5524 ( \5901 , \5898 , \5900 );
xor \U$5525 ( \5902 , \5889 , \5901 );
and \U$5526 ( \5903 , \5399 , RIae78a58_123);
and \U$5527 ( \5904 , RIae78cb0_128, \5397 );
nor \U$5528 ( \5905 , \5903 , \5904 );
and \U$5529 ( \5906 , \5905 , \5016 );
not \U$5530 ( \5907 , \5905 );
and \U$5531 ( \5908 , \5907 , \5403 );
nor \U$5532 ( \5909 , \5906 , \5908 );
and \U$5533 ( \5910 , \5902 , \5909 );
and \U$5534 ( \5911 , \5889 , \5901 );
or \U$5535 ( \5912 , \5910 , \5911 );
and \U$5536 ( \5913 , \5882 , \5912 );
and \U$5537 ( \5914 , \5855 , \5881 );
or \U$5538 ( \5915 , \5913 , \5914 );
not \U$5539 ( \5916 , \388 );
and \U$5540 ( \5917 , \384 , RIae78968_121);
and \U$5541 ( \5918 , RIae78878_119, \382 );
nor \U$5542 ( \5919 , \5917 , \5918 );
not \U$5543 ( \5920 , \5919 );
or \U$5544 ( \5921 , \5916 , \5920 );
or \U$5545 ( \5922 , \5919 , \392 );
nand \U$5546 ( \5923 , \5921 , \5922 );
not \U$5547 ( \5924 , RIae77e28_97);
nor \U$5548 ( \5925 , \5924 , \491 );
xor \U$5549 ( \5926 , \5923 , \5925 );
nand \U$5550 ( \5927 , RIae77d38_95, RIae78b48_125);
and \U$5551 ( \5928 , \384 , RIae77e28_97);
and \U$5552 ( \5929 , RIae78968_121, \382 );
nor \U$5553 ( \5930 , \5928 , \5929 );
not \U$5554 ( \5931 , \5930 );
not \U$5555 ( \5932 , \388 );
and \U$5556 ( \5933 , \5931 , \5932 );
and \U$5557 ( \5934 , \5930 , \388 );
nor \U$5558 ( \5935 , \5933 , \5934 );
nand \U$5559 ( \5936 , \5927 , \5935 );
and \U$5560 ( \5937 , \5926 , \5936 );
and \U$5561 ( \5938 , \5923 , \5925 );
or \U$5562 ( \5939 , \5937 , \5938 );
xor \U$5563 ( \5940 , \5915 , \5939 );
and \U$5564 ( \5941 , \1939 , RIae75128_1);
and \U$5565 ( \5942 , RIae75308_5, \1937 );
nor \U$5566 ( \5943 , \5941 , \5942 );
and \U$5567 ( \5944 , \5943 , \1735 );
not \U$5568 ( \5945 , \5943 );
and \U$5569 ( \5946 , \5945 , \1734 );
nor \U$5570 ( \5947 , \5944 , \5946 );
and \U$5571 ( \5948 , \1376 , RIae754e8_9);
and \U$5572 ( \5949 , RIae757b8_15, \1374 );
nor \U$5573 ( \5950 , \5948 , \5949 );
and \U$5574 ( \5951 , \5950 , \1380 );
not \U$5575 ( \5952 , \5950 );
and \U$5576 ( \5953 , \5952 , \1261 );
nor \U$5577 ( \5954 , \5951 , \5953 );
xor \U$5578 ( \5955 , \5947 , \5954 );
and \U$5579 ( \5956 , \1593 , RIae756c8_13);
and \U$5580 ( \5957 , RIae75218_3, \1591 );
nor \U$5581 ( \5958 , \5956 , \5957 );
and \U$5582 ( \5959 , \5958 , \1498 );
not \U$5583 ( \5960 , \5958 );
and \U$5584 ( \5961 , \5960 , \1488 );
nor \U$5585 ( \5962 , \5959 , \5961 );
and \U$5586 ( \5963 , \5955 , \5962 );
and \U$5587 ( \5964 , \5947 , \5954 );
or \U$5588 ( \5965 , \5963 , \5964 );
and \U$5589 ( \5966 , \672 , RIae758a8_17);
and \U$5590 ( \5967 , RIae75f38_31, \670 );
nor \U$5591 ( \5968 , \5966 , \5967 );
and \U$5592 ( \5969 , \5968 , \588 );
not \U$5593 ( \5970 , \5968 );
and \U$5594 ( \5971 , \5970 , \587 );
nor \U$5595 ( \5972 , \5969 , \5971 );
not \U$5596 ( \5973 , \789 );
and \U$5597 ( \5974 , \883 , RIae75e48_29);
and \U$5598 ( \5975 , RIae75c68_25, \881 );
nor \U$5599 ( \5976 , \5974 , \5975 );
not \U$5600 ( \5977 , \5976 );
or \U$5601 ( \5978 , \5973 , \5977 );
or \U$5602 ( \5979 , \5976 , \787 );
nand \U$5603 ( \5980 , \5978 , \5979 );
xor \U$5604 ( \5981 , \5972 , \5980 );
and \U$5605 ( \5982 , \1138 , RIae75d58_27);
and \U$5606 ( \5983 , RIae755d8_11, \1136 );
nor \U$5607 ( \5984 , \5982 , \5983 );
and \U$5608 ( \5985 , \5984 , \1012 );
not \U$5609 ( \5986 , \5984 );
and \U$5610 ( \5987 , \5986 , \1142 );
nor \U$5611 ( \5988 , \5985 , \5987 );
and \U$5612 ( \5989 , \5981 , \5988 );
and \U$5613 ( \5990 , \5972 , \5980 );
or \U$5614 ( \5991 , \5989 , \5990 );
xor \U$5615 ( \5992 , \5965 , \5991 );
not \U$5616 ( \5993 , \400 );
and \U$5617 ( \5994 , \436 , RIae78878_119);
and \U$5618 ( \5995 , RIae78788_117, \434 );
nor \U$5619 ( \5996 , \5994 , \5995 );
not \U$5620 ( \5997 , \5996 );
or \U$5621 ( \5998 , \5993 , \5997 );
or \U$5622 ( \5999 , \5996 , \400 );
nand \U$5623 ( \6000 , \5998 , \5999 );
not \U$5624 ( \6001 , \469 );
and \U$5625 ( \6002 , \514 , RIae78698_115);
and \U$5626 ( \6003 , RIae75b78_23, \512 );
nor \U$5627 ( \6004 , \6002 , \6003 );
not \U$5628 ( \6005 , \6004 );
or \U$5629 ( \6006 , \6001 , \6005 );
or \U$5630 ( \6007 , \6004 , \471 );
nand \U$5631 ( \6008 , \6006 , \6007 );
xor \U$5632 ( \6009 , \6000 , \6008 );
and \U$5633 ( \6010 , \558 , RIae75a88_21);
and \U$5634 ( \6011 , RIae75998_19, \556 );
nor \U$5635 ( \6012 , \6010 , \6011 );
and \U$5636 ( \6013 , \6012 , \504 );
not \U$5637 ( \6014 , \6012 );
and \U$5638 ( \6015 , \6014 , \562 );
nor \U$5639 ( \6016 , \6013 , \6015 );
and \U$5640 ( \6017 , \6009 , \6016 );
and \U$5641 ( \6018 , \6000 , \6008 );
or \U$5642 ( \6019 , \6017 , \6018 );
and \U$5643 ( \6020 , \5992 , \6019 );
and \U$5644 ( \6021 , \5965 , \5991 );
or \U$5645 ( \6022 , \6020 , \6021 );
and \U$5646 ( \6023 , \5940 , \6022 );
and \U$5647 ( \6024 , \5915 , \5939 );
or \U$5648 ( \6025 , \6023 , \6024 );
xor \U$5649 ( \6026 , \5829 , \6025 );
or \U$5650 ( \6027 , \5634 , \5632 );
nand \U$5651 ( \6028 , \6027 , \5635 );
xor \U$5652 ( \6029 , \5391 , \5405 );
xor \U$5653 ( \6030 , \6029 , \5413 );
xor \U$5654 ( \6031 , \6028 , \6030 );
xor \U$5655 ( \6032 , \5335 , \5342 );
xor \U$5656 ( \6033 , \6032 , \5351 );
xor \U$5657 ( \6034 , \5724 , \5729 );
xor \U$5658 ( \6035 , \6033 , \6034 );
and \U$5659 ( \6036 , \6031 , \6035 );
and \U$5660 ( \6037 , \6028 , \6030 );
or \U$5661 ( \6038 , \6036 , \6037 );
and \U$5662 ( \6039 , \6026 , \6038 );
and \U$5663 ( \6040 , \5829 , \6025 );
or \U$5664 ( \6041 , \6039 , \6040 );
xor \U$5665 ( \6042 , \5799 , \6041 );
xor \U$5666 ( \6043 , \5474 , \5476 );
xor \U$5667 ( \6044 , \6043 , \5481 );
xor \U$5668 ( \6045 , \5528 , \5535 );
xor \U$5669 ( \6046 , \6044 , \6045 );
and \U$5670 ( \6047 , \6042 , \6046 );
and \U$5671 ( \6048 , \5799 , \6041 );
or \U$5672 ( \6049 , \6047 , \6048 );
xor \U$5673 ( \6050 , \5274 , \5461 );
xor \U$5674 ( \6051 , \6050 , \5484 );
xor \U$5675 ( \6052 , \6049 , \6051 );
xor \U$5676 ( \6053 , \5540 , \5747 );
xor \U$5677 ( \6054 , \6053 , \5758 );
and \U$5678 ( \6055 , \6052 , \6054 );
and \U$5679 ( \6056 , \6049 , \6051 );
or \U$5680 ( \6057 , \6055 , \6056 );
nand \U$5681 ( \6058 , \5785 , \6057 );
or \U$5682 ( \6059 , \5774 , \6058 );
xnor \U$5683 ( \6060 , \6058 , \5774 );
and \U$5684 ( \6061 , \1593 , RIae754e8_9);
and \U$5685 ( \6062 , RIae757b8_15, \1591 );
nor \U$5686 ( \6063 , \6061 , \6062 );
and \U$5687 ( \6064 , \6063 , \1498 );
not \U$5688 ( \6065 , \6063 );
and \U$5689 ( \6066 , \6065 , \1488 );
nor \U$5690 ( \6067 , \6064 , \6066 );
and \U$5691 ( \6068 , \1939 , RIae756c8_13);
and \U$5692 ( \6069 , RIae75218_3, \1937 );
nor \U$5693 ( \6070 , \6068 , \6069 );
and \U$5694 ( \6071 , \6070 , \1735 );
not \U$5695 ( \6072 , \6070 );
and \U$5696 ( \6073 , \6072 , \1734 );
nor \U$5697 ( \6074 , \6071 , \6073 );
xor \U$5698 ( \6075 , \6067 , \6074 );
and \U$5699 ( \6076 , \2224 , RIae75128_1);
and \U$5700 ( \6077 , RIae75308_5, \2222 );
nor \U$5701 ( \6078 , \6076 , \6077 );
and \U$5702 ( \6079 , \6078 , \2061 );
not \U$5703 ( \6080 , \6078 );
and \U$5704 ( \6081 , \6080 , \2060 );
nor \U$5705 ( \6082 , \6079 , \6081 );
xor \U$5706 ( \6083 , \6075 , \6082 );
not \U$5707 ( \6084 , \471 );
and \U$5708 ( \6085 , \514 , RIae78878_119);
and \U$5709 ( \6086 , RIae78788_117, \512 );
nor \U$5710 ( \6087 , \6085 , \6086 );
not \U$5711 ( \6088 , \6087 );
or \U$5712 ( \6089 , \6084 , \6088 );
or \U$5713 ( \6090 , \6087 , \471 );
nand \U$5714 ( \6091 , \6089 , \6090 );
and \U$5715 ( \6092 , \558 , RIae78698_115);
and \U$5716 ( \6093 , RIae75b78_23, \556 );
nor \U$5717 ( \6094 , \6092 , \6093 );
and \U$5718 ( \6095 , \6094 , \504 );
not \U$5719 ( \6096 , \6094 );
and \U$5720 ( \6097 , \6096 , \562 );
nor \U$5721 ( \6098 , \6095 , \6097 );
xor \U$5722 ( \6099 , \6091 , \6098 );
and \U$5723 ( \6100 , \672 , RIae75a88_21);
and \U$5724 ( \6101 , RIae75998_19, \670 );
nor \U$5725 ( \6102 , \6100 , \6101 );
and \U$5726 ( \6103 , \6102 , \588 );
not \U$5727 ( \6104 , \6102 );
and \U$5728 ( \6105 , \6104 , \587 );
nor \U$5729 ( \6106 , \6103 , \6105 );
xor \U$5730 ( \6107 , \6099 , \6106 );
and \U$5731 ( \6108 , \6083 , \6107 );
and \U$5732 ( \6109 , \1138 , RIae75e48_29);
and \U$5733 ( \6110 , RIae75c68_25, \1136 );
nor \U$5734 ( \6111 , \6109 , \6110 );
and \U$5735 ( \6112 , \6111 , \1012 );
not \U$5736 ( \6113 , \6111 );
and \U$5737 ( \6114 , \6113 , \1142 );
nor \U$5738 ( \6115 , \6112 , \6114 );
not \U$5739 ( \6116 , \787 );
and \U$5740 ( \6117 , \883 , RIae758a8_17);
and \U$5741 ( \6118 , RIae75f38_31, \881 );
nor \U$5742 ( \6119 , \6117 , \6118 );
not \U$5743 ( \6120 , \6119 );
or \U$5744 ( \6121 , \6116 , \6120 );
or \U$5745 ( \6122 , \6119 , \787 );
nand \U$5746 ( \6123 , \6121 , \6122 );
xor \U$5747 ( \6124 , \6115 , \6123 );
and \U$5748 ( \6125 , \1376 , RIae75d58_27);
and \U$5749 ( \6126 , RIae755d8_11, \1374 );
nor \U$5750 ( \6127 , \6125 , \6126 );
and \U$5751 ( \6128 , \6127 , \1380 );
not \U$5752 ( \6129 , \6127 );
and \U$5753 ( \6130 , \6129 , \1261 );
nor \U$5754 ( \6131 , \6128 , \6130 );
xor \U$5755 ( \6132 , \6124 , \6131 );
xor \U$5756 ( \6133 , \6091 , \6098 );
xor \U$5757 ( \6134 , \6133 , \6106 );
and \U$5758 ( \6135 , \6132 , \6134 );
and \U$5759 ( \6136 , \6083 , \6132 );
or \U$5760 ( \6137 , \6108 , \6135 , \6136 );
not \U$5761 ( \6138 , \6137 );
and \U$5762 ( \6139 , \4247 , RIae76a78_55);
and \U$5763 ( \6140 , RIae76988_53, \4245 );
nor \U$5764 ( \6141 , \6139 , \6140 );
and \U$5765 ( \6142 , \6141 , \4251 );
not \U$5766 ( \6143 , \6141 );
and \U$5767 ( \6144 , \6143 , \3989 );
nor \U$5768 ( \6145 , \6142 , \6144 );
and \U$5769 ( \6146 , \4688 , RIae767a8_49);
and \U$5770 ( \6147 , RIae76898_51, \4686 );
nor \U$5771 ( \6148 , \6146 , \6147 );
and \U$5772 ( \6149 , \6148 , \4482 );
not \U$5773 ( \6150 , \6148 );
and \U$5774 ( \6151 , \6150 , \4481 );
nor \U$5775 ( \6152 , \6149 , \6151 );
xor \U$5776 ( \6153 , \6145 , \6152 );
and \U$5777 ( \6154 , \3730 , RIae762f8_39);
and \U$5778 ( \6155 , RIae76208_37, \3728 );
nor \U$5779 ( \6156 , \6154 , \6155 );
and \U$5780 ( \6157 , \6156 , \3422 );
not \U$5781 ( \6158 , \6156 );
and \U$5782 ( \6159 , \6158 , \3732 );
nor \U$5783 ( \6160 , \6157 , \6159 );
xor \U$5784 ( \6161 , \6153 , \6160 );
or \U$5785 ( \6162 , \6138 , \6161 );
not \U$5786 ( \6163 , \6161 );
not \U$5787 ( \6164 , \6138 );
or \U$5788 ( \6165 , \6163 , \6164 );
and \U$5789 ( \6166 , RIae79ef8_167, RIae79f70_168);
not \U$5790 ( \6167 , RIae79fe8_169);
and \U$5791 ( \6168 , \6167 , RIae79f70_168);
nor \U$5792 ( \6169 , \6167 , RIae79f70_168);
or \U$5793 ( \6170 , \6168 , \6169 );
nor \U$5794 ( \6171 , RIae79ef8_167, RIae79f70_168);
nor \U$5795 ( \6172 , \6166 , \6170 , \6171 );
nand \U$5796 ( \6173 , RIae78da0_130, \6172 );
nand \U$5797 ( \6174 , RIae79fe8_169, RIae79f70_168);
and \U$5798 ( \6175 , \6174 , RIae79ef8_167);
not \U$5799 ( \6176 , \6175 );
and \U$5800 ( \6177 , \6173 , \6176 );
not \U$5801 ( \6178 , \6173 );
and \U$5802 ( \6179 , \6178 , \6175 );
nor \U$5803 ( \6180 , \6177 , \6179 );
not \U$5804 ( \6181 , \6180 );
and \U$5805 ( \6182 , \5896 , RIae78a58_123);
and \U$5806 ( \6183 , RIae78cb0_128, \5894 );
nor \U$5807 ( \6184 , \6182 , \6183 );
and \U$5808 ( \6185 , \6184 , \5589 );
not \U$5809 ( \6186 , \6184 );
and \U$5810 ( \6187 , \6186 , \5590 );
nor \U$5811 ( \6188 , \6185 , \6187 );
not \U$5812 ( \6189 , \6188 );
or \U$5813 ( \6190 , \6181 , \6189 );
or \U$5814 ( \6191 , \6188 , \6180 );
nand \U$5815 ( \6192 , \6190 , \6191 );
not \U$5816 ( \6193 , \6192 );
and \U$5817 ( \6194 , \5399 , RIae76898_51);
and \U$5818 ( \6195 , RIae76b68_57, \5397 );
nor \U$5819 ( \6196 , \6194 , \6195 );
and \U$5820 ( \6197 , \6196 , \5403 );
not \U$5821 ( \6198 , \6196 );
and \U$5822 ( \6199 , \6198 , \5016 );
nor \U$5823 ( \6200 , \6197 , \6199 );
not \U$5824 ( \6201 , \6200 );
and \U$5825 ( \6202 , \6193 , \6201 );
and \U$5826 ( \6203 , \6192 , \6200 );
nor \U$5827 ( \6204 , \6202 , \6203 );
and \U$5828 ( \6205 , \4247 , RIae76208_37);
and \U$5829 ( \6206 , RIae76a78_55, \4245 );
nor \U$5830 ( \6207 , \6205 , \6206 );
and \U$5831 ( \6208 , \6207 , \4251 );
not \U$5832 ( \6209 , \6207 );
and \U$5833 ( \6210 , \6209 , \3989 );
nor \U$5834 ( \6211 , \6208 , \6210 );
not \U$5835 ( \6212 , \6211 );
and \U$5836 ( \6213 , \4688 , RIae76988_53);
and \U$5837 ( \6214 , RIae767a8_49, \4686 );
nor \U$5838 ( \6215 , \6213 , \6214 );
and \U$5839 ( \6216 , \6215 , \4481 );
not \U$5840 ( \6217 , \6215 );
and \U$5841 ( \6218 , \6217 , \4482 );
nor \U$5842 ( \6219 , \6216 , \6218 );
not \U$5843 ( \6220 , \6219 );
or \U$5844 ( \6221 , \6212 , \6220 );
or \U$5845 ( \6222 , \6211 , \6219 );
nand \U$5846 ( \6223 , \6221 , \6222 );
not \U$5847 ( \6224 , \6223 );
and \U$5848 ( \6225 , \3730 , RIae76028_33);
and \U$5849 ( \6226 , RIae762f8_39, \3728 );
nor \U$5850 ( \6227 , \6225 , \6226 );
and \U$5851 ( \6228 , \6227 , \3422 );
not \U$5852 ( \6229 , \6227 );
and \U$5853 ( \6230 , \6229 , \3732 );
nor \U$5854 ( \6231 , \6228 , \6230 );
not \U$5855 ( \6232 , \6231 );
and \U$5856 ( \6233 , \6224 , \6232 );
and \U$5857 ( \6234 , \6223 , \6231 );
nor \U$5858 ( \6235 , \6233 , \6234 );
xor \U$5859 ( \6236 , \6204 , \6235 );
and \U$5860 ( \6237 , \3214 , RIae765c8_45);
and \U$5861 ( \6238 , RIae76118_35, \3212 );
nor \U$5862 ( \6239 , \6237 , \6238 );
not \U$5863 ( \6240 , \6239 );
not \U$5864 ( \6241 , \2774 );
and \U$5865 ( \6242 , \6240 , \6241 );
and \U$5866 ( \6243 , \6239 , \2774 );
nor \U$5867 ( \6244 , \6242 , \6243 );
not \U$5868 ( \6245 , \6244 );
not \U$5869 ( \6246 , \3089 );
and \U$5870 ( \6247 , \2783 , RIae764d8_43);
and \U$5871 ( \6248 , RIae766b8_47, \2781 );
nor \U$5872 ( \6249 , \6247 , \6248 );
not \U$5873 ( \6250 , \6249 );
or \U$5874 ( \6251 , \6246 , \6250 );
or \U$5875 ( \6252 , \6249 , \2789 );
nand \U$5876 ( \6253 , \6251 , \6252 );
not \U$5877 ( \6254 , \6253 );
or \U$5878 ( \6255 , \6245 , \6254 );
or \U$5879 ( \6256 , \6244 , \6253 );
nand \U$5880 ( \6257 , \6255 , \6256 );
not \U$5881 ( \6258 , \6257 );
and \U$5882 ( \6259 , \2607 , RIae753f8_7);
and \U$5883 ( \6260 , RIae763e8_41, \2605 );
nor \U$5884 ( \6261 , \6259 , \6260 );
and \U$5885 ( \6262 , \6261 , \2397 );
not \U$5886 ( \6263 , \6261 );
and \U$5887 ( \6264 , \6263 , \2611 );
nor \U$5888 ( \6265 , \6262 , \6264 );
not \U$5889 ( \6266 , \6265 );
and \U$5890 ( \6267 , \6258 , \6266 );
and \U$5891 ( \6268 , \6257 , \6265 );
nor \U$5892 ( \6269 , \6267 , \6268 );
and \U$5893 ( \6270 , \6236 , \6269 );
and \U$5894 ( \6271 , \6204 , \6235 );
nor \U$5895 ( \6272 , \6270 , \6271 );
nand \U$5896 ( \6273 , \6165 , \6272 );
nand \U$5897 ( \6274 , \6162 , \6273 );
and \U$5898 ( \6275 , \2783 , RIae763e8_41);
and \U$5899 ( \6276 , RIae764d8_43, \2781 );
nor \U$5900 ( \6277 , \6275 , \6276 );
not \U$5901 ( \6278 , \6277 );
not \U$5902 ( \6279 , \3089 );
and \U$5903 ( \6280 , \6278 , \6279 );
and \U$5904 ( \6281 , \6277 , \2789 );
nor \U$5905 ( \6282 , \6280 , \6281 );
and \U$5906 ( \6283 , \3730 , RIae76118_35);
and \U$5907 ( \6284 , RIae76028_33, \3728 );
nor \U$5908 ( \6285 , \6283 , \6284 );
and \U$5909 ( \6286 , \6285 , \3422 );
not \U$5910 ( \6287 , \6285 );
and \U$5911 ( \6288 , \6287 , \3732 );
nor \U$5912 ( \6289 , \6286 , \6288 );
or \U$5913 ( \6290 , \6282 , \6289 );
not \U$5914 ( \6291 , \6289 );
not \U$5915 ( \6292 , \6282 );
or \U$5916 ( \6293 , \6291 , \6292 );
not \U$5917 ( \6294 , \3218 );
and \U$5918 ( \6295 , \3214 , RIae766b8_47);
and \U$5919 ( \6296 , RIae765c8_45, \3212 );
nor \U$5920 ( \6297 , \6295 , \6296 );
not \U$5921 ( \6298 , \6297 );
or \U$5922 ( \6299 , \6294 , \6298 );
or \U$5923 ( \6300 , \6297 , \2774 );
nand \U$5924 ( \6301 , \6299 , \6300 );
nand \U$5925 ( \6302 , \6293 , \6301 );
nand \U$5926 ( \6303 , \6290 , \6302 );
and \U$5927 ( \6304 , \6172 , RIae78cb0_128);
and \U$5928 ( \6305 , RIae78da0_130, \6170 );
nor \U$5929 ( \6306 , \6304 , \6305 );
and \U$5930 ( \6307 , \6306 , \6176 );
not \U$5931 ( \6308 , \6306 );
and \U$5932 ( \6309 , \6308 , \6175 );
nor \U$5933 ( \6310 , \6307 , \6309 );
not \U$5934 ( \6311 , RIae7a2b8_175);
not \U$5935 ( \6312 , RIae7a678_183);
or \U$5936 ( \6313 , \6311 , \6312 );
nand \U$5937 ( \6314 , \6313 , RIae79fe8_169);
xor \U$5938 ( \6315 , \6310 , \6314 );
and \U$5939 ( \6316 , \5896 , RIae76b68_57);
and \U$5940 ( \6317 , RIae78a58_123, \5894 );
nor \U$5941 ( \6318 , \6316 , \6317 );
and \U$5942 ( \6319 , \6318 , \5590 );
not \U$5943 ( \6320 , \6318 );
and \U$5944 ( \6321 , \6320 , \5589 );
nor \U$5945 ( \6322 , \6319 , \6321 );
and \U$5946 ( \6323 , \6315 , \6322 );
and \U$5947 ( \6324 , \6310 , \6314 );
or \U$5948 ( \6325 , \6323 , \6324 );
xor \U$5949 ( \6326 , \6303 , \6325 );
and \U$5950 ( \6327 , \4688 , RIae76a78_55);
and \U$5951 ( \6328 , RIae76988_53, \4686 );
nor \U$5952 ( \6329 , \6327 , \6328 );
and \U$5953 ( \6330 , \6329 , \4482 );
not \U$5954 ( \6331 , \6329 );
and \U$5955 ( \6332 , \6331 , \4481 );
nor \U$5956 ( \6333 , \6330 , \6332 );
and \U$5957 ( \6334 , \5399 , RIae767a8_49);
and \U$5958 ( \6335 , RIae76898_51, \5397 );
nor \U$5959 ( \6336 , \6334 , \6335 );
and \U$5960 ( \6337 , \6336 , \5403 );
not \U$5961 ( \6338 , \6336 );
and \U$5962 ( \6339 , \6338 , \5016 );
nor \U$5963 ( \6340 , \6337 , \6339 );
xor \U$5964 ( \6341 , \6333 , \6340 );
and \U$5965 ( \6342 , \4247 , RIae762f8_39);
and \U$5966 ( \6343 , RIae76208_37, \4245 );
nor \U$5967 ( \6344 , \6342 , \6343 );
and \U$5968 ( \6345 , \6344 , \4251 );
not \U$5969 ( \6346 , \6344 );
and \U$5970 ( \6347 , \6346 , \3989 );
nor \U$5971 ( \6348 , \6345 , \6347 );
and \U$5972 ( \6349 , \6341 , \6348 );
and \U$5973 ( \6350 , \6333 , \6340 );
nor \U$5974 ( \6351 , \6349 , \6350 );
and \U$5975 ( \6352 , \6326 , \6351 );
and \U$5976 ( \6353 , \6303 , \6325 );
or \U$5977 ( \6354 , \6352 , \6353 );
and \U$5978 ( \6355 , \384 , RIae77c48_93);
and \U$5979 ( \6356 , RIae77b58_91, \382 );
nor \U$5980 ( \6357 , \6355 , \6356 );
not \U$5981 ( \6358 , \6357 );
not \U$5982 ( \6359 , \392 );
and \U$5983 ( \6360 , \6358 , \6359 );
and \U$5984 ( \6361 , \6357 , \388 );
nor \U$5985 ( \6362 , \6360 , \6361 );
and \U$5986 ( \6363 , \436 , RIae77d38_95);
and \U$5987 ( \6364 , RIae77e28_97, \434 );
nor \U$5988 ( \6365 , \6363 , \6364 );
not \U$5989 ( \6366 , \6365 );
not \U$5990 ( \6367 , \400 );
and \U$5991 ( \6368 , \6366 , \6367 );
and \U$5992 ( \6369 , \6365 , \402 );
nor \U$5993 ( \6370 , \6368 , \6369 );
xor \U$5994 ( \6371 , \6362 , \6370 );
and \U$5995 ( \6372 , \514 , RIae78968_121);
and \U$5996 ( \6373 , RIae78878_119, \512 );
nor \U$5997 ( \6374 , \6372 , \6373 );
not \U$5998 ( \6375 , \6374 );
not \U$5999 ( \6376 , \471 );
and \U$6000 ( \6377 , \6375 , \6376 );
and \U$6001 ( \6378 , \6374 , \469 );
nor \U$6002 ( \6379 , \6377 , \6378 );
and \U$6003 ( \6380 , \6371 , \6379 );
and \U$6004 ( \6381 , \6362 , \6370 );
or \U$6005 ( \6382 , \6380 , \6381 );
and \U$6006 ( \6383 , \384 , RIae77b58_91);
and \U$6007 ( \6384 , RIae77d38_95, \382 );
nor \U$6008 ( \6385 , \6383 , \6384 );
not \U$6009 ( \6386 , \6385 );
not \U$6010 ( \6387 , \388 );
and \U$6011 ( \6388 , \6386 , \6387 );
and \U$6012 ( \6389 , \6385 , \392 );
nor \U$6013 ( \6390 , \6388 , \6389 );
not \U$6014 ( \6391 , \6390 );
not \U$6015 ( \6392 , \400 );
and \U$6016 ( \6393 , \436 , RIae77e28_97);
and \U$6017 ( \6394 , RIae78968_121, \434 );
nor \U$6018 ( \6395 , \6393 , \6394 );
not \U$6019 ( \6396 , \6395 );
or \U$6020 ( \6397 , \6392 , \6396 );
or \U$6021 ( \6398 , \6395 , \400 );
nand \U$6022 ( \6399 , \6397 , \6398 );
not \U$6023 ( \6400 , \6399 );
or \U$6024 ( \6401 , \6391 , \6400 );
or \U$6025 ( \6402 , \6390 , \6399 );
nand \U$6026 ( \6403 , \6401 , \6402 );
not \U$6027 ( \6404 , \6403 );
nand \U$6028 ( \6405 , RIae77c48_93, RIae78b48_125);
not \U$6029 ( \6406 , \6405 );
and \U$6030 ( \6407 , \6404 , \6406 );
and \U$6031 ( \6408 , \6403 , \6405 );
nor \U$6032 ( \6409 , \6407 , \6408 );
nand \U$6033 ( \6410 , \6382 , \6409 );
xor \U$6034 ( \6411 , \6354 , \6410 );
and \U$6035 ( \6412 , \2224 , RIae75218_3);
and \U$6036 ( \6413 , RIae75128_1, \2222 );
nor \U$6037 ( \6414 , \6412 , \6413 );
and \U$6038 ( \6415 , \6414 , \2060 );
not \U$6039 ( \6416 , \6414 );
and \U$6040 ( \6417 , \6416 , \2061 );
nor \U$6041 ( \6418 , \6415 , \6417 );
and \U$6042 ( \6419 , \2607 , RIae75308_5);
and \U$6043 ( \6420 , RIae753f8_7, \2605 );
nor \U$6044 ( \6421 , \6419 , \6420 );
and \U$6045 ( \6422 , \6421 , \2397 );
not \U$6046 ( \6423 , \6421 );
and \U$6047 ( \6424 , \6423 , \2611 );
nor \U$6048 ( \6425 , \6422 , \6424 );
xor \U$6049 ( \6426 , \6418 , \6425 );
and \U$6050 ( \6427 , \1939 , RIae757b8_15);
and \U$6051 ( \6428 , RIae756c8_13, \1937 );
nor \U$6052 ( \6429 , \6427 , \6428 );
and \U$6053 ( \6430 , \6429 , \1734 );
not \U$6054 ( \6431 , \6429 );
and \U$6055 ( \6432 , \6431 , \1735 );
nor \U$6056 ( \6433 , \6430 , \6432 );
and \U$6057 ( \6434 , \6426 , \6433 );
and \U$6058 ( \6435 , \6418 , \6425 );
nor \U$6059 ( \6436 , \6434 , \6435 );
and \U$6060 ( \6437 , \672 , RIae75b78_23);
and \U$6061 ( \6438 , RIae75a88_21, \670 );
nor \U$6062 ( \6439 , \6437 , \6438 );
and \U$6063 ( \6440 , \6439 , \587 );
not \U$6064 ( \6441 , \6439 );
and \U$6065 ( \6442 , \6441 , \588 );
nor \U$6066 ( \6443 , \6440 , \6442 );
and \U$6067 ( \6444 , \883 , RIae75998_19);
and \U$6068 ( \6445 , RIae758a8_17, \881 );
nor \U$6069 ( \6446 , \6444 , \6445 );
not \U$6070 ( \6447 , \6446 );
not \U$6071 ( \6448 , \787 );
and \U$6072 ( \6449 , \6447 , \6448 );
and \U$6073 ( \6450 , \6446 , \787 );
nor \U$6074 ( \6451 , \6449 , \6450 );
xor \U$6075 ( \6452 , \6443 , \6451 );
and \U$6076 ( \6453 , \558 , RIae78788_117);
and \U$6077 ( \6454 , RIae78698_115, \556 );
nor \U$6078 ( \6455 , \6453 , \6454 );
and \U$6079 ( \6456 , \6455 , \562 );
not \U$6080 ( \6457 , \6455 );
and \U$6081 ( \6458 , \6457 , \504 );
nor \U$6082 ( \6459 , \6456 , \6458 );
and \U$6083 ( \6460 , \6452 , \6459 );
and \U$6084 ( \6461 , \6443 , \6451 );
nor \U$6085 ( \6462 , \6460 , \6461 );
xor \U$6086 ( \6463 , \6436 , \6462 );
and \U$6087 ( \6464 , \1138 , RIae75f38_31);
and \U$6088 ( \6465 , RIae75e48_29, \1136 );
nor \U$6089 ( \6466 , \6464 , \6465 );
and \U$6090 ( \6467 , \6466 , \1142 );
not \U$6091 ( \6468 , \6466 );
and \U$6092 ( \6469 , \6468 , \1012 );
nor \U$6093 ( \6470 , \6467 , \6469 );
and \U$6094 ( \6471 , \1376 , RIae75c68_25);
and \U$6095 ( \6472 , RIae75d58_27, \1374 );
nor \U$6096 ( \6473 , \6471 , \6472 );
and \U$6097 ( \6474 , \6473 , \1261 );
not \U$6098 ( \6475 , \6473 );
and \U$6099 ( \6476 , \6475 , \1380 );
nor \U$6100 ( \6477 , \6474 , \6476 );
or \U$6101 ( \6478 , \6470 , \6477 );
not \U$6102 ( \6479 , \6477 );
not \U$6103 ( \6480 , \6470 );
or \U$6104 ( \6481 , \6479 , \6480 );
and \U$6105 ( \6482 , \1593 , RIae755d8_11);
and \U$6106 ( \6483 , RIae754e8_9, \1591 );
nor \U$6107 ( \6484 , \6482 , \6483 );
and \U$6108 ( \6485 , \6484 , \1498 );
not \U$6109 ( \6486 , \6484 );
and \U$6110 ( \6487 , \6486 , \1488 );
nor \U$6111 ( \6488 , \6485 , \6487 );
nand \U$6112 ( \6489 , \6481 , \6488 );
nand \U$6113 ( \6490 , \6478 , \6489 );
and \U$6114 ( \6491 , \6463 , \6490 );
and \U$6115 ( \6492 , \6436 , \6462 );
or \U$6116 ( \6493 , \6491 , \6492 );
and \U$6117 ( \6494 , \6411 , \6493 );
and \U$6118 ( \6495 , \6354 , \6410 );
or \U$6119 ( \6496 , \6494 , \6495 );
xor \U$6120 ( \6497 , \6274 , \6496 );
and \U$6121 ( \6498 , \5896 , RIae78cb0_128);
and \U$6122 ( \6499 , RIae78da0_130, \5894 );
nor \U$6123 ( \6500 , \6498 , \6499 );
and \U$6124 ( \6501 , \6500 , \5590 );
not \U$6125 ( \6502 , \6500 );
and \U$6126 ( \6503 , \6502 , \5589 );
nor \U$6127 ( \6504 , \6501 , \6503 );
xor \U$6128 ( \6505 , \6504 , \6176 );
and \U$6129 ( \6506 , \5399 , RIae76b68_57);
and \U$6130 ( \6507 , RIae78a58_123, \5397 );
nor \U$6131 ( \6508 , \6506 , \6507 );
and \U$6132 ( \6509 , \6508 , \5016 );
not \U$6133 ( \6510 , \6508 );
and \U$6134 ( \6511 , \6510 , \5403 );
nor \U$6135 ( \6512 , \6509 , \6511 );
xor \U$6136 ( \6513 , \6505 , \6512 );
not \U$6137 ( \6514 , \400 );
and \U$6138 ( \6515 , \436 , RIae78968_121);
and \U$6139 ( \6516 , RIae78878_119, \434 );
nor \U$6140 ( \6517 , \6515 , \6516 );
not \U$6141 ( \6518 , \6517 );
or \U$6142 ( \6519 , \6514 , \6518 );
or \U$6143 ( \6520 , \6517 , \402 );
nand \U$6144 ( \6521 , \6519 , \6520 );
not \U$6145 ( \6522 , RIae77b58_91);
nor \U$6146 ( \6523 , \6522 , \491 );
xor \U$6147 ( \6524 , \6521 , \6523 );
not \U$6148 ( \6525 , \388 );
and \U$6149 ( \6526 , \384 , RIae77d38_95);
and \U$6150 ( \6527 , RIae77e28_97, \382 );
nor \U$6151 ( \6528 , \6526 , \6527 );
not \U$6152 ( \6529 , \6528 );
or \U$6153 ( \6530 , \6525 , \6529 );
or \U$6154 ( \6531 , \6528 , \392 );
nand \U$6155 ( \6532 , \6530 , \6531 );
xor \U$6156 ( \6533 , \6524 , \6532 );
or \U$6157 ( \6534 , \6390 , \6405 );
not \U$6158 ( \6535 , \6405 );
not \U$6159 ( \6536 , \6390 );
or \U$6160 ( \6537 , \6535 , \6536 );
nand \U$6161 ( \6538 , \6537 , \6399 );
nand \U$6162 ( \6539 , \6534 , \6538 );
xor \U$6163 ( \6540 , \6533 , \6539 );
and \U$6164 ( \6541 , \558 , RIae75b78_23);
and \U$6165 ( \6542 , RIae75a88_21, \556 );
nor \U$6166 ( \6543 , \6541 , \6542 );
and \U$6167 ( \6544 , \6543 , \504 );
not \U$6168 ( \6545 , \6543 );
and \U$6169 ( \6546 , \6545 , \562 );
nor \U$6170 ( \6547 , \6544 , \6546 );
not \U$6171 ( \6548 , \469 );
and \U$6172 ( \6549 , \514 , RIae78788_117);
and \U$6173 ( \6550 , RIae78698_115, \512 );
nor \U$6174 ( \6551 , \6549 , \6550 );
not \U$6175 ( \6552 , \6551 );
or \U$6176 ( \6553 , \6548 , \6552 );
or \U$6177 ( \6554 , \6551 , \469 );
nand \U$6178 ( \6555 , \6553 , \6554 );
xor \U$6179 ( \6556 , \6547 , \6555 );
and \U$6180 ( \6557 , \672 , RIae75998_19);
and \U$6181 ( \6558 , RIae758a8_17, \670 );
nor \U$6182 ( \6559 , \6557 , \6558 );
and \U$6183 ( \6560 , \6559 , \588 );
not \U$6184 ( \6561 , \6559 );
and \U$6185 ( \6562 , \6561 , \587 );
nor \U$6186 ( \6563 , \6560 , \6562 );
xor \U$6187 ( \6564 , \6556 , \6563 );
xor \U$6188 ( \6565 , \6540 , \6564 );
and \U$6189 ( \6566 , \6513 , \6565 );
and \U$6190 ( \6567 , \1138 , RIae75c68_25);
and \U$6191 ( \6568 , RIae75d58_27, \1136 );
nor \U$6192 ( \6569 , \6567 , \6568 );
and \U$6193 ( \6570 , \6569 , \1012 );
not \U$6194 ( \6571 , \6569 );
and \U$6195 ( \6572 , \6571 , \1142 );
nor \U$6196 ( \6573 , \6570 , \6572 );
not \U$6197 ( \6574 , \789 );
and \U$6198 ( \6575 , \883 , RIae75f38_31);
and \U$6199 ( \6576 , RIae75e48_29, \881 );
nor \U$6200 ( \6577 , \6575 , \6576 );
not \U$6201 ( \6578 , \6577 );
or \U$6202 ( \6579 , \6574 , \6578 );
or \U$6203 ( \6580 , \6577 , \787 );
nand \U$6204 ( \6581 , \6579 , \6580 );
xor \U$6205 ( \6582 , \6573 , \6581 );
and \U$6206 ( \6583 , \1376 , RIae755d8_11);
and \U$6207 ( \6584 , RIae754e8_9, \1374 );
nor \U$6208 ( \6585 , \6583 , \6584 );
and \U$6209 ( \6586 , \6585 , \1380 );
not \U$6210 ( \6587 , \6585 );
and \U$6211 ( \6588 , \6587 , \1261 );
nor \U$6212 ( \6589 , \6586 , \6588 );
xor \U$6213 ( \6590 , \6582 , \6589 );
and \U$6214 ( \6591 , \2224 , RIae75308_5);
and \U$6215 ( \6592 , RIae753f8_7, \2222 );
nor \U$6216 ( \6593 , \6591 , \6592 );
and \U$6217 ( \6594 , \6593 , \2061 );
not \U$6218 ( \6595 , \6593 );
and \U$6219 ( \6596 , \6595 , \2060 );
nor \U$6220 ( \6597 , \6594 , \6596 );
and \U$6221 ( \6598 , \1593 , RIae757b8_15);
and \U$6222 ( \6599 , RIae756c8_13, \1591 );
nor \U$6223 ( \6600 , \6598 , \6599 );
and \U$6224 ( \6601 , \6600 , \1498 );
not \U$6225 ( \6602 , \6600 );
and \U$6226 ( \6603 , \6602 , \1488 );
nor \U$6227 ( \6604 , \6601 , \6603 );
xor \U$6228 ( \6605 , \6597 , \6604 );
and \U$6229 ( \6606 , \1939 , RIae75218_3);
and \U$6230 ( \6607 , RIae75128_1, \1937 );
nor \U$6231 ( \6608 , \6606 , \6607 );
and \U$6232 ( \6609 , \6608 , \1735 );
not \U$6233 ( \6610 , \6608 );
and \U$6234 ( \6611 , \6610 , \1734 );
nor \U$6235 ( \6612 , \6609 , \6611 );
xor \U$6236 ( \6613 , \6605 , \6612 );
not \U$6237 ( \6614 , \3218 );
and \U$6238 ( \6615 , \3214 , RIae76118_35);
and \U$6239 ( \6616 , RIae76028_33, \3212 );
nor \U$6240 ( \6617 , \6615 , \6616 );
not \U$6241 ( \6618 , \6617 );
or \U$6242 ( \6619 , \6614 , \6618 );
or \U$6243 ( \6620 , \6617 , \2774 );
nand \U$6244 ( \6621 , \6619 , \6620 );
and \U$6245 ( \6622 , \2607 , RIae763e8_41);
and \U$6246 ( \6623 , RIae764d8_43, \2605 );
nor \U$6247 ( \6624 , \6622 , \6623 );
and \U$6248 ( \6625 , \6624 , \2611 );
not \U$6249 ( \6626 , \6624 );
and \U$6250 ( \6627 , \6626 , \2396 );
nor \U$6251 ( \6628 , \6625 , \6627 );
xor \U$6252 ( \6629 , \6621 , \6628 );
not \U$6253 ( \6630 , \3089 );
and \U$6254 ( \6631 , \2783 , RIae766b8_47);
and \U$6255 ( \6632 , RIae765c8_45, \2781 );
nor \U$6256 ( \6633 , \6631 , \6632 );
not \U$6257 ( \6634 , \6633 );
or \U$6258 ( \6635 , \6630 , \6634 );
or \U$6259 ( \6636 , \6633 , \2789 );
nand \U$6260 ( \6637 , \6635 , \6636 );
xor \U$6261 ( \6638 , \6629 , \6637 );
xor \U$6262 ( \6639 , \6613 , \6638 );
xor \U$6263 ( \6640 , \6590 , \6639 );
xor \U$6264 ( \6641 , \6533 , \6539 );
xor \U$6265 ( \6642 , \6641 , \6564 );
and \U$6266 ( \6643 , \6640 , \6642 );
and \U$6267 ( \6644 , \6513 , \6640 );
or \U$6268 ( \6645 , \6566 , \6643 , \6644 );
and \U$6269 ( \6646 , \6497 , \6645 );
and \U$6270 ( \6647 , \6274 , \6496 );
or \U$6271 ( \6648 , \6646 , \6647 );
xor \U$6272 ( \6649 , \6597 , \6604 );
and \U$6273 ( \6650 , \6649 , \6612 );
and \U$6274 ( \6651 , \6597 , \6604 );
or \U$6275 ( \6652 , \6650 , \6651 );
xor \U$6276 ( \6653 , \6573 , \6581 );
and \U$6277 ( \6654 , \6653 , \6589 );
and \U$6278 ( \6655 , \6573 , \6581 );
or \U$6279 ( \6656 , \6654 , \6655 );
xor \U$6280 ( \6657 , \6652 , \6656 );
xor \U$6281 ( \6658 , \6547 , \6555 );
and \U$6282 ( \6659 , \6658 , \6563 );
and \U$6283 ( \6660 , \6547 , \6555 );
or \U$6284 ( \6661 , \6659 , \6660 );
and \U$6285 ( \6662 , \6657 , \6661 );
and \U$6286 ( \6663 , \6652 , \6656 );
or \U$6287 ( \6664 , \6662 , \6663 );
xor \U$6288 ( \6665 , \6145 , \6152 );
and \U$6289 ( \6666 , \6665 , \6160 );
and \U$6290 ( \6667 , \6145 , \6152 );
nor \U$6291 ( \6668 , \6666 , \6667 );
xor \U$6292 ( \6669 , \6504 , \6176 );
and \U$6293 ( \6670 , \6669 , \6512 );
and \U$6294 ( \6671 , \6504 , \6176 );
or \U$6295 ( \6672 , \6670 , \6671 );
xor \U$6296 ( \6673 , \6668 , \6672 );
xor \U$6297 ( \6674 , \6621 , \6628 );
and \U$6298 ( \6675 , \6674 , \6637 );
and \U$6299 ( \6676 , \6621 , \6628 );
or \U$6300 ( \6677 , \6675 , \6676 );
and \U$6301 ( \6678 , \6673 , \6677 );
and \U$6302 ( \6679 , \6668 , \6672 );
or \U$6303 ( \6680 , \6678 , \6679 );
xor \U$6304 ( \6681 , \6664 , \6680 );
xor \U$6305 ( \6682 , \6521 , \6523 );
and \U$6306 ( \6683 , \6682 , \6532 );
and \U$6307 ( \6684 , \6521 , \6523 );
or \U$6308 ( \6685 , \6683 , \6684 );
or \U$6309 ( \6686 , \5935 , \5927 );
nand \U$6310 ( \6687 , \6686 , \5936 );
xor \U$6311 ( \6688 , \6685 , \6687 );
xor \U$6312 ( \6689 , \6000 , \6008 );
xor \U$6313 ( \6690 , \6689 , \6016 );
and \U$6314 ( \6691 , \6688 , \6690 );
and \U$6315 ( \6692 , \6685 , \6687 );
or \U$6316 ( \6693 , \6691 , \6692 );
xor \U$6317 ( \6694 , \6681 , \6693 );
xor \U$6318 ( \6695 , \6648 , \6694 );
xor \U$6319 ( \6696 , \6067 , \6074 );
and \U$6320 ( \6697 , \6696 , \6082 );
and \U$6321 ( \6698 , \6067 , \6074 );
or \U$6322 ( \6699 , \6697 , \6698 );
xor \U$6323 ( \6700 , \6115 , \6123 );
and \U$6324 ( \6701 , \6700 , \6131 );
and \U$6325 ( \6702 , \6115 , \6123 );
or \U$6326 ( \6703 , \6701 , \6702 );
xor \U$6327 ( \6704 , \6699 , \6703 );
xor \U$6328 ( \6705 , \6091 , \6098 );
and \U$6329 ( \6706 , \6705 , \6106 );
and \U$6330 ( \6707 , \6091 , \6098 );
or \U$6331 ( \6708 , \6706 , \6707 );
and \U$6332 ( \6709 , \6704 , \6708 );
and \U$6333 ( \6710 , \6699 , \6703 );
or \U$6334 ( \6711 , \6709 , \6710 );
or \U$6335 ( \6712 , \6265 , \6244 );
not \U$6336 ( \6713 , \6244 );
not \U$6337 ( \6714 , \6265 );
or \U$6338 ( \6715 , \6713 , \6714 );
nand \U$6339 ( \6716 , \6715 , \6253 );
nand \U$6340 ( \6717 , \6712 , \6716 );
or \U$6341 ( \6718 , \6200 , \6188 );
not \U$6342 ( \6719 , \6188 );
not \U$6343 ( \6720 , \6200 );
or \U$6344 ( \6721 , \6719 , \6720 );
nand \U$6345 ( \6722 , \6721 , \6180 );
nand \U$6346 ( \6723 , \6718 , \6722 );
xor \U$6347 ( \6724 , \6717 , \6723 );
or \U$6348 ( \6725 , \6231 , \6211 );
not \U$6349 ( \6726 , \6211 );
not \U$6350 ( \6727 , \6231 );
or \U$6351 ( \6728 , \6726 , \6727 );
nand \U$6352 ( \6729 , \6728 , \6219 );
nand \U$6353 ( \6730 , \6725 , \6729 );
and \U$6354 ( \6731 , \6724 , \6730 );
and \U$6355 ( \6732 , \6717 , \6723 );
or \U$6356 ( \6733 , \6731 , \6732 );
xor \U$6357 ( \6734 , \6711 , \6733 );
xor \U$6358 ( \6735 , \6533 , \6539 );
and \U$6359 ( \6736 , \6735 , \6564 );
and \U$6360 ( \6737 , \6533 , \6539 );
or \U$6361 ( \6738 , \6736 , \6737 );
xor \U$6362 ( \6739 , \6734 , \6738 );
xor \U$6363 ( \6740 , \6668 , \6672 );
xor \U$6364 ( \6741 , \6740 , \6677 );
xor \U$6365 ( \6742 , \6652 , \6656 );
xor \U$6366 ( \6743 , \6742 , \6661 );
xor \U$6367 ( \6744 , \6741 , \6743 );
xor \U$6368 ( \6745 , \6685 , \6687 );
xor \U$6369 ( \6746 , \6745 , \6690 );
xor \U$6370 ( \6747 , \6744 , \6746 );
and \U$6371 ( \6748 , \6739 , \6747 );
xor \U$6372 ( \6749 , \6573 , \6581 );
xor \U$6373 ( \6750 , \6749 , \6589 );
and \U$6374 ( \6751 , \6613 , \6750 );
xor \U$6375 ( \6752 , \6573 , \6581 );
xor \U$6376 ( \6753 , \6752 , \6589 );
and \U$6377 ( \6754 , \6638 , \6753 );
and \U$6378 ( \6755 , \6613 , \6638 );
or \U$6379 ( \6756 , \6751 , \6754 , \6755 );
xor \U$6380 ( \6757 , \5836 , \5844 );
xor \U$6381 ( \6758 , \6757 , \5852 );
xor \U$6382 ( \6759 , \5889 , \5901 );
xor \U$6383 ( \6760 , \6759 , \5909 );
xor \U$6384 ( \6761 , \6758 , \6760 );
xor \U$6385 ( \6762 , \6756 , \6761 );
xor \U$6386 ( \6763 , \5862 , \5869 );
xor \U$6387 ( \6764 , \6763 , \5878 );
xor \U$6388 ( \6765 , \5972 , \5980 );
xor \U$6389 ( \6766 , \6765 , \5988 );
xor \U$6390 ( \6767 , \5947 , \5954 );
xor \U$6391 ( \6768 , \6767 , \5962 );
xor \U$6392 ( \6769 , \6766 , \6768 );
xor \U$6393 ( \6770 , \6764 , \6769 );
xor \U$6394 ( \6771 , \6762 , \6770 );
xor \U$6395 ( \6772 , \6741 , \6743 );
xor \U$6396 ( \6773 , \6772 , \6746 );
and \U$6397 ( \6774 , \6771 , \6773 );
and \U$6398 ( \6775 , \6739 , \6771 );
or \U$6399 ( \6776 , \6748 , \6774 , \6775 );
and \U$6400 ( \6777 , \6695 , \6776 );
and \U$6401 ( \6778 , \6648 , \6694 );
or \U$6402 ( \6779 , \6777 , \6778 );
xor \U$6403 ( \6780 , \6741 , \6743 );
and \U$6404 ( \6781 , \6780 , \6746 );
and \U$6405 ( \6782 , \6741 , \6743 );
or \U$6406 ( \6783 , \6781 , \6782 );
xor \U$6407 ( \6784 , \6711 , \6733 );
and \U$6408 ( \6785 , \6784 , \6738 );
and \U$6409 ( \6786 , \6711 , \6733 );
or \U$6410 ( \6787 , \6785 , \6786 );
xor \U$6411 ( \6788 , \6783 , \6787 );
xor \U$6412 ( \6789 , \6756 , \6761 );
and \U$6413 ( \6790 , \6789 , \6770 );
and \U$6414 ( \6791 , \6756 , \6761 );
or \U$6415 ( \6792 , \6790 , \6791 );
xor \U$6416 ( \6793 , \6788 , \6792 );
xor \U$6417 ( \6794 , \5862 , \5869 );
xor \U$6418 ( \6795 , \6794 , \5878 );
and \U$6419 ( \6796 , \6766 , \6795 );
xor \U$6420 ( \6797 , \5862 , \5869 );
xor \U$6421 ( \6798 , \6797 , \5878 );
and \U$6422 ( \6799 , \6768 , \6798 );
and \U$6423 ( \6800 , \6766 , \6768 );
or \U$6424 ( \6801 , \6796 , \6799 , \6800 );
and \U$6425 ( \6802 , \6758 , \6760 );
xor \U$6426 ( \6803 , \6801 , \6802 );
xor \U$6427 ( \6804 , \5609 , \5617 );
xor \U$6428 ( \6805 , \6804 , \5625 );
xor \U$6429 ( \6806 , \5801 , \5806 );
xor \U$6430 ( \6807 , \6805 , \6806 );
xor \U$6431 ( \6808 , \6803 , \6807 );
xor \U$6432 ( \6809 , \5855 , \5881 );
xor \U$6433 ( \6810 , \6809 , \5912 );
xor \U$6434 ( \6811 , \5965 , \5991 );
xor \U$6435 ( \6812 , \6811 , \6019 );
xor \U$6436 ( \6813 , \5923 , \5925 );
xor \U$6437 ( \6814 , \6813 , \5936 );
xor \U$6438 ( \6815 , \5670 , \5678 );
xor \U$6439 ( \6816 , \6815 , \5686 );
xor \U$6440 ( \6817 , \5816 , \5821 );
xor \U$6441 ( \6818 , \6816 , \6817 );
xor \U$6442 ( \6819 , \6814 , \6818 );
xor \U$6443 ( \6820 , \6812 , \6819 );
xor \U$6444 ( \6821 , \6810 , \6820 );
xor \U$6445 ( \6822 , \6808 , \6821 );
and \U$6446 ( \6823 , \6793 , \6822 );
xor \U$6447 ( \6824 , \6779 , \6823 );
xor \U$6448 ( \6825 , \5580 , \5601 );
xor \U$6449 ( \6826 , \6825 , \5628 );
xor \U$6450 ( \6827 , \5662 , \5689 );
xor \U$6451 ( \6828 , \6827 , \5715 );
xor \U$6452 ( \6829 , \6826 , \6828 );
xor \U$6453 ( \6830 , \6028 , \6030 );
xor \U$6454 ( \6831 , \6830 , \6035 );
xor \U$6455 ( \6832 , \6829 , \6831 );
xor \U$6456 ( \6833 , \5915 , \5939 );
xor \U$6457 ( \6834 , \6833 , \6022 );
xor \U$6458 ( \6835 , \5965 , \5991 );
xor \U$6459 ( \6836 , \6835 , \6019 );
and \U$6460 ( \6837 , \6814 , \6836 );
xor \U$6461 ( \6838 , \5965 , \5991 );
xor \U$6462 ( \6839 , \6838 , \6019 );
and \U$6463 ( \6840 , \6818 , \6839 );
and \U$6464 ( \6841 , \6814 , \6818 );
or \U$6465 ( \6842 , \6837 , \6840 , \6841 );
xor \U$6466 ( \6843 , \6664 , \6680 );
and \U$6467 ( \6844 , \6843 , \6693 );
and \U$6468 ( \6845 , \6664 , \6680 );
or \U$6469 ( \6846 , \6844 , \6845 );
xor \U$6470 ( \6847 , \6842 , \6846 );
xor \U$6471 ( \6848 , \6801 , \6802 );
and \U$6472 ( \6849 , \6848 , \6807 );
and \U$6473 ( \6850 , \6801 , \6802 );
or \U$6474 ( \6851 , \6849 , \6850 );
xor \U$6475 ( \6852 , \6847 , \6851 );
xor \U$6476 ( \6853 , \6834 , \6852 );
xor \U$6477 ( \6854 , \6832 , \6853 );
and \U$6478 ( \6855 , \6824 , \6854 );
and \U$6479 ( \6856 , \6779 , \6823 );
or \U$6480 ( \6857 , \6855 , \6856 );
xor \U$6481 ( \6858 , \6842 , \6846 );
and \U$6482 ( \6859 , \6858 , \6851 );
and \U$6483 ( \6860 , \6842 , \6846 );
or \U$6484 ( \6861 , \6859 , \6860 );
xor \U$6485 ( \6862 , \6826 , \6828 );
and \U$6486 ( \6863 , \6862 , \6831 );
and \U$6487 ( \6864 , \6826 , \6828 );
or \U$6488 ( \6865 , \6863 , \6864 );
xor \U$6489 ( \6866 , \6861 , \6865 );
xor \U$6490 ( \6867 , \5734 , \5736 );
xor \U$6491 ( \6868 , \6867 , \5741 );
xor \U$6492 ( \6869 , \5787 , \5794 );
xor \U$6493 ( \6870 , \6868 , \6869 );
xor \U$6494 ( \6871 , \6866 , \6870 );
xor \U$6495 ( \6872 , \6857 , \6871 );
xor \U$6496 ( \6873 , \5829 , \6025 );
xor \U$6497 ( \6874 , \6873 , \6038 );
xor \U$6498 ( \6875 , \6826 , \6828 );
xor \U$6499 ( \6876 , \6875 , \6831 );
and \U$6500 ( \6877 , \6834 , \6876 );
xor \U$6501 ( \6878 , \6826 , \6828 );
xor \U$6502 ( \6879 , \6878 , \6831 );
and \U$6503 ( \6880 , \6852 , \6879 );
and \U$6504 ( \6881 , \6834 , \6852 );
or \U$6505 ( \6882 , \6877 , \6880 , \6881 );
xor \U$6506 ( \6883 , \6874 , \6882 );
xor \U$6507 ( \6884 , \6783 , \6787 );
and \U$6508 ( \6885 , \6884 , \6792 );
and \U$6509 ( \6886 , \6783 , \6787 );
or \U$6510 ( \6887 , \6885 , \6886 );
xor \U$6511 ( \6888 , \5811 , \5813 );
xor \U$6512 ( \6889 , \6888 , \5826 );
xor \U$6513 ( \6890 , \6887 , \6889 );
xor \U$6514 ( \6891 , \6801 , \6802 );
xor \U$6515 ( \6892 , \6891 , \6807 );
and \U$6516 ( \6893 , \6810 , \6892 );
xor \U$6517 ( \6894 , \6801 , \6802 );
xor \U$6518 ( \6895 , \6894 , \6807 );
and \U$6519 ( \6896 , \6820 , \6895 );
and \U$6520 ( \6897 , \6810 , \6820 );
or \U$6521 ( \6898 , \6893 , \6896 , \6897 );
and \U$6522 ( \6899 , \6890 , \6898 );
and \U$6523 ( \6900 , \6887 , \6889 );
or \U$6524 ( \6901 , \6899 , \6900 );
xor \U$6525 ( \6902 , \6883 , \6901 );
and \U$6526 ( \6903 , \6872 , \6902 );
and \U$6527 ( \6904 , \6857 , \6871 );
or \U$6528 ( \6905 , \6903 , \6904 );
xor \U$6529 ( \6906 , \6874 , \6882 );
and \U$6530 ( \6907 , \6906 , \6901 );
and \U$6531 ( \6908 , \6874 , \6882 );
nor \U$6532 ( \6909 , \6907 , \6908 );
not \U$6533 ( \6910 , \6909 );
xor \U$6534 ( \6911 , \6861 , \6865 );
and \U$6535 ( \6912 , \6911 , \6870 );
and \U$6536 ( \6913 , \6861 , \6865 );
or \U$6537 ( \6914 , \6912 , \6913 );
xor \U$6538 ( \6915 , \5554 , \5721 );
xor \U$6539 ( \6916 , \6915 , \5744 );
xor \U$6540 ( \6917 , \6914 , \6916 );
xor \U$6541 ( \6918 , \5799 , \6041 );
xor \U$6542 ( \6919 , \6918 , \6046 );
xor \U$6543 ( \6920 , \6917 , \6919 );
not \U$6544 ( \6921 , \6920 );
or \U$6545 ( \6922 , \6910 , \6921 );
or \U$6546 ( \6923 , \6920 , \6909 );
nand \U$6547 ( \6924 , \6922 , \6923 );
and \U$6548 ( \6925 , \6905 , \6924 );
xor \U$6549 ( \6926 , \6924 , \6905 );
and \U$6550 ( \6927 , \5896 , RIae76898_51);
and \U$6551 ( \6928 , RIae76b68_57, \5894 );
nor \U$6552 ( \6929 , \6927 , \6928 );
and \U$6553 ( \6930 , \6929 , \5590 );
not \U$6554 ( \6931 , \6929 );
and \U$6555 ( \6932 , \6931 , \5589 );
nor \U$6556 ( \6933 , \6930 , \6932 );
and \U$6557 ( \6934 , RIae79fe8_169, RIae7a678_183);
not \U$6558 ( \6935 , RIae7a678_183);
nor \U$6559 ( \6936 , \6935 , RIae7a2b8_175);
not \U$6560 ( \6937 , RIae7a2b8_175);
nor \U$6561 ( \6938 , \6937 , RIae7a678_183);
or \U$6562 ( \6939 , \6936 , \6938 );
nor \U$6563 ( \6940 , RIae79fe8_169, RIae7a678_183);
nor \U$6564 ( \6941 , \6934 , \6939 , \6940 );
nand \U$6565 ( \6942 , RIae78da0_130, \6941 );
and \U$6566 ( \6943 , \6942 , \6314 );
not \U$6567 ( \6944 , \6942 );
not \U$6568 ( \6945 , \6314 );
and \U$6569 ( \6946 , \6944 , \6945 );
nor \U$6570 ( \6947 , \6943 , \6946 );
xor \U$6571 ( \6948 , \6933 , \6947 );
and \U$6572 ( \6949 , \6172 , RIae78a58_123);
and \U$6573 ( \6950 , RIae78cb0_128, \6170 );
nor \U$6574 ( \6951 , \6949 , \6950 );
and \U$6575 ( \6952 , \6951 , \6176 );
not \U$6576 ( \6953 , \6951 );
and \U$6577 ( \6954 , \6953 , \6175 );
nor \U$6578 ( \6955 , \6952 , \6954 );
xor \U$6579 ( \6956 , \6948 , \6955 );
and \U$6580 ( \6957 , \5399 , RIae76988_53);
and \U$6581 ( \6958 , RIae767a8_49, \5397 );
nor \U$6582 ( \6959 , \6957 , \6958 );
and \U$6583 ( \6960 , \6959 , \5016 );
not \U$6584 ( \6961 , \6959 );
and \U$6585 ( \6962 , \6961 , \5403 );
nor \U$6586 ( \6963 , \6960 , \6962 );
and \U$6587 ( \6964 , \4247 , RIae76028_33);
and \U$6588 ( \6965 , RIae762f8_39, \4245 );
nor \U$6589 ( \6966 , \6964 , \6965 );
and \U$6590 ( \6967 , \6966 , \3989 );
not \U$6591 ( \6968 , \6966 );
and \U$6592 ( \6969 , \6968 , \4251 );
nor \U$6593 ( \6970 , \6967 , \6969 );
xor \U$6594 ( \6971 , \6963 , \6970 );
and \U$6595 ( \6972 , \4688 , RIae76208_37);
and \U$6596 ( \6973 , RIae76a78_55, \4686 );
nor \U$6597 ( \6974 , \6972 , \6973 );
and \U$6598 ( \6975 , \6974 , \4481 );
not \U$6599 ( \6976 , \6974 );
and \U$6600 ( \6977 , \6976 , \4482 );
nor \U$6601 ( \6978 , \6975 , \6977 );
xor \U$6602 ( \6979 , \6971 , \6978 );
and \U$6603 ( \6980 , \6956 , \6979 );
and \U$6604 ( \6981 , \3730 , RIae765c8_45);
and \U$6605 ( \6982 , RIae76118_35, \3728 );
nor \U$6606 ( \6983 , \6981 , \6982 );
and \U$6607 ( \6984 , \6983 , \3732 );
not \U$6608 ( \6985 , \6983 );
and \U$6609 ( \6986 , \6985 , \3422 );
nor \U$6610 ( \6987 , \6984 , \6986 );
not \U$6611 ( \6988 , \2789 );
and \U$6612 ( \6989 , \2783 , RIae753f8_7);
and \U$6613 ( \6990 , RIae763e8_41, \2781 );
nor \U$6614 ( \6991 , \6989 , \6990 );
not \U$6615 ( \6992 , \6991 );
or \U$6616 ( \6993 , \6988 , \6992 );
or \U$6617 ( \6994 , \6991 , \3089 );
nand \U$6618 ( \6995 , \6993 , \6994 );
xor \U$6619 ( \6996 , \6987 , \6995 );
not \U$6620 ( \6997 , \2774 );
and \U$6621 ( \6998 , \3214 , RIae764d8_43);
and \U$6622 ( \6999 , RIae766b8_47, \3212 );
nor \U$6623 ( \7000 , \6998 , \6999 );
not \U$6624 ( \7001 , \7000 );
or \U$6625 ( \7002 , \6997 , \7001 );
or \U$6626 ( \7003 , \7000 , \3218 );
nand \U$6627 ( \7004 , \7002 , \7003 );
xor \U$6628 ( \7005 , \6996 , \7004 );
xor \U$6629 ( \7006 , \6963 , \6970 );
xor \U$6630 ( \7007 , \7006 , \6978 );
and \U$6631 ( \7008 , \7005 , \7007 );
and \U$6632 ( \7009 , \6956 , \7005 );
or \U$6633 ( \7010 , \6980 , \7008 , \7009 );
xor \U$6634 ( \7011 , \6310 , \6314 );
xor \U$6635 ( \7012 , \7011 , \6322 );
xor \U$6636 ( \7013 , \7010 , \7012 );
not \U$6637 ( \7014 , \789 );
and \U$6638 ( \7015 , \883 , RIae75a88_21);
and \U$6639 ( \7016 , RIae75998_19, \881 );
nor \U$6640 ( \7017 , \7015 , \7016 );
not \U$6641 ( \7018 , \7017 );
or \U$6642 ( \7019 , \7014 , \7018 );
or \U$6643 ( \7020 , \7017 , \787 );
nand \U$6644 ( \7021 , \7019 , \7020 );
and \U$6645 ( \7022 , \558 , RIae78878_119);
and \U$6646 ( \7023 , RIae78788_117, \556 );
nor \U$6647 ( \7024 , \7022 , \7023 );
and \U$6648 ( \7025 , \7024 , \504 );
not \U$6649 ( \7026 , \7024 );
and \U$6650 ( \7027 , \7026 , \562 );
nor \U$6651 ( \7028 , \7025 , \7027 );
xor \U$6652 ( \7029 , \7021 , \7028 );
and \U$6653 ( \7030 , \672 , RIae78698_115);
and \U$6654 ( \7031 , RIae75b78_23, \670 );
nor \U$6655 ( \7032 , \7030 , \7031 );
and \U$6656 ( \7033 , \7032 , \588 );
not \U$6657 ( \7034 , \7032 );
and \U$6658 ( \7035 , \7034 , \587 );
nor \U$6659 ( \7036 , \7033 , \7035 );
xor \U$6660 ( \7037 , \7029 , \7036 );
and \U$6661 ( \7038 , \1376 , RIae75e48_29);
and \U$6662 ( \7039 , RIae75c68_25, \1374 );
nor \U$6663 ( \7040 , \7038 , \7039 );
and \U$6664 ( \7041 , \7040 , \1380 );
not \U$6665 ( \7042 , \7040 );
and \U$6666 ( \7043 , \7042 , \1261 );
nor \U$6667 ( \7044 , \7041 , \7043 );
and \U$6668 ( \7045 , \1138 , RIae758a8_17);
and \U$6669 ( \7046 , RIae75f38_31, \1136 );
nor \U$6670 ( \7047 , \7045 , \7046 );
and \U$6671 ( \7048 , \7047 , \1012 );
not \U$6672 ( \7049 , \7047 );
and \U$6673 ( \7050 , \7049 , \1142 );
nor \U$6674 ( \7051 , \7048 , \7050 );
xor \U$6675 ( \7052 , \7044 , \7051 );
and \U$6676 ( \7053 , \1593 , RIae75d58_27);
and \U$6677 ( \7054 , RIae755d8_11, \1591 );
nor \U$6678 ( \7055 , \7053 , \7054 );
and \U$6679 ( \7056 , \7055 , \1498 );
not \U$6680 ( \7057 , \7055 );
and \U$6681 ( \7058 , \7057 , \1488 );
nor \U$6682 ( \7059 , \7056 , \7058 );
xor \U$6683 ( \7060 , \7052 , \7059 );
xor \U$6684 ( \7061 , \7037 , \7060 );
and \U$6685 ( \7062 , \1939 , RIae754e8_9);
and \U$6686 ( \7063 , RIae757b8_15, \1937 );
nor \U$6687 ( \7064 , \7062 , \7063 );
and \U$6688 ( \7065 , \7064 , \1735 );
not \U$6689 ( \7066 , \7064 );
and \U$6690 ( \7067 , \7066 , \1734 );
nor \U$6691 ( \7068 , \7065 , \7067 );
and \U$6692 ( \7069 , \2224 , RIae756c8_13);
and \U$6693 ( \7070 , RIae75218_3, \2222 );
nor \U$6694 ( \7071 , \7069 , \7070 );
and \U$6695 ( \7072 , \7071 , \2061 );
not \U$6696 ( \7073 , \7071 );
and \U$6697 ( \7074 , \7073 , \2060 );
nor \U$6698 ( \7075 , \7072 , \7074 );
xor \U$6699 ( \7076 , \7068 , \7075 );
and \U$6700 ( \7077 , \2607 , RIae75128_1);
and \U$6701 ( \7078 , RIae75308_5, \2605 );
nor \U$6702 ( \7079 , \7077 , \7078 );
and \U$6703 ( \7080 , \7079 , \2611 );
not \U$6704 ( \7081 , \7079 );
and \U$6705 ( \7082 , \7081 , \2397 );
nor \U$6706 ( \7083 , \7080 , \7082 );
xor \U$6707 ( \7084 , \7076 , \7083 );
and \U$6708 ( \7085 , \7061 , \7084 );
and \U$6709 ( \7086 , \7037 , \7060 );
or \U$6710 ( \7087 , \7085 , \7086 );
and \U$6711 ( \7088 , \7013 , \7087 );
and \U$6712 ( \7089 , \7010 , \7012 );
or \U$6713 ( \7090 , \7088 , \7089 );
and \U$6714 ( \7091 , \1939 , RIae755d8_11);
and \U$6715 ( \7092 , RIae754e8_9, \1937 );
nor \U$6716 ( \7093 , \7091 , \7092 );
and \U$6717 ( \7094 , \7093 , \1735 );
not \U$6718 ( \7095 , \7093 );
and \U$6719 ( \7096 , \7095 , \1734 );
nor \U$6720 ( \7097 , \7094 , \7096 );
and \U$6721 ( \7098 , \1376 , RIae75f38_31);
and \U$6722 ( \7099 , RIae75e48_29, \1374 );
nor \U$6723 ( \7100 , \7098 , \7099 );
and \U$6724 ( \7101 , \7100 , \1380 );
not \U$6725 ( \7102 , \7100 );
and \U$6726 ( \7103 , \7102 , \1261 );
nor \U$6727 ( \7104 , \7101 , \7103 );
xor \U$6728 ( \7105 , \7097 , \7104 );
and \U$6729 ( \7106 , \1593 , RIae75c68_25);
and \U$6730 ( \7107 , RIae75d58_27, \1591 );
nor \U$6731 ( \7108 , \7106 , \7107 );
and \U$6732 ( \7109 , \7108 , \1498 );
not \U$6733 ( \7110 , \7108 );
and \U$6734 ( \7111 , \7110 , \1488 );
nor \U$6735 ( \7112 , \7109 , \7111 );
and \U$6736 ( \7113 , \7105 , \7112 );
and \U$6737 ( \7114 , \7097 , \7104 );
or \U$6738 ( \7115 , \7113 , \7114 );
not \U$6739 ( \7116 , \789 );
and \U$6740 ( \7117 , \883 , RIae75b78_23);
and \U$6741 ( \7118 , RIae75a88_21, \881 );
nor \U$6742 ( \7119 , \7117 , \7118 );
not \U$6743 ( \7120 , \7119 );
or \U$6744 ( \7121 , \7116 , \7120 );
or \U$6745 ( \7122 , \7119 , \787 );
nand \U$6746 ( \7123 , \7121 , \7122 );
and \U$6747 ( \7124 , \672 , RIae78788_117);
and \U$6748 ( \7125 , RIae78698_115, \670 );
nor \U$6749 ( \7126 , \7124 , \7125 );
and \U$6750 ( \7127 , \7126 , \588 );
not \U$6751 ( \7128 , \7126 );
and \U$6752 ( \7129 , \7128 , \587 );
nor \U$6753 ( \7130 , \7127 , \7129 );
xor \U$6754 ( \7131 , \7123 , \7130 );
and \U$6755 ( \7132 , \1138 , RIae75998_19);
and \U$6756 ( \7133 , RIae758a8_17, \1136 );
nor \U$6757 ( \7134 , \7132 , \7133 );
and \U$6758 ( \7135 , \7134 , \1012 );
not \U$6759 ( \7136 , \7134 );
and \U$6760 ( \7137 , \7136 , \1142 );
nor \U$6761 ( \7138 , \7135 , \7137 );
and \U$6762 ( \7139 , \7131 , \7138 );
and \U$6763 ( \7140 , \7123 , \7130 );
or \U$6764 ( \7141 , \7139 , \7140 );
xor \U$6765 ( \7142 , \7115 , \7141 );
not \U$6766 ( \7143 , \2789 );
and \U$6767 ( \7144 , \2783 , RIae75308_5);
and \U$6768 ( \7145 , RIae753f8_7, \2781 );
nor \U$6769 ( \7146 , \7144 , \7145 );
not \U$6770 ( \7147 , \7146 );
or \U$6771 ( \7148 , \7143 , \7147 );
or \U$6772 ( \7149 , \7146 , \2789 );
nand \U$6773 ( \7150 , \7148 , \7149 );
and \U$6774 ( \7151 , \2224 , RIae757b8_15);
and \U$6775 ( \7152 , RIae756c8_13, \2222 );
nor \U$6776 ( \7153 , \7151 , \7152 );
and \U$6777 ( \7154 , \7153 , \2061 );
not \U$6778 ( \7155 , \7153 );
and \U$6779 ( \7156 , \7155 , \2060 );
nor \U$6780 ( \7157 , \7154 , \7156 );
xor \U$6781 ( \7158 , \7150 , \7157 );
and \U$6782 ( \7159 , \2607 , RIae75218_3);
and \U$6783 ( \7160 , RIae75128_1, \2605 );
nor \U$6784 ( \7161 , \7159 , \7160 );
and \U$6785 ( \7162 , \7161 , \2611 );
not \U$6786 ( \7163 , \7161 );
and \U$6787 ( \7164 , \7163 , \2397 );
nor \U$6788 ( \7165 , \7162 , \7164 );
and \U$6789 ( \7166 , \7158 , \7165 );
and \U$6790 ( \7167 , \7150 , \7157 );
or \U$6791 ( \7168 , \7166 , \7167 );
and \U$6792 ( \7169 , \7142 , \7168 );
and \U$6793 ( \7170 , \7115 , \7141 );
or \U$6794 ( \7171 , \7169 , \7170 );
and \U$6795 ( \7172 , \5399 , RIae76a78_55);
and \U$6796 ( \7173 , RIae76988_53, \5397 );
nor \U$6797 ( \7174 , \7172 , \7173 );
and \U$6798 ( \7175 , \7174 , \5016 );
not \U$6799 ( \7176 , \7174 );
and \U$6800 ( \7177 , \7176 , \5403 );
nor \U$6801 ( \7178 , \7175 , \7177 );
and \U$6802 ( \7179 , \4688 , RIae762f8_39);
and \U$6803 ( \7180 , RIae76208_37, \4686 );
nor \U$6804 ( \7181 , \7179 , \7180 );
and \U$6805 ( \7182 , \7181 , \4481 );
not \U$6806 ( \7183 , \7181 );
and \U$6807 ( \7184 , \7183 , \4482 );
nor \U$6808 ( \7185 , \7182 , \7184 );
xor \U$6809 ( \7186 , \7178 , \7185 );
and \U$6810 ( \7187 , \5896 , RIae767a8_49);
and \U$6811 ( \7188 , RIae76898_51, \5894 );
nor \U$6812 ( \7189 , \7187 , \7188 );
and \U$6813 ( \7190 , \7189 , \5590 );
not \U$6814 ( \7191 , \7189 );
and \U$6815 ( \7192 , \7191 , \5589 );
nor \U$6816 ( \7193 , \7190 , \7192 );
and \U$6817 ( \7194 , \7186 , \7193 );
and \U$6818 ( \7195 , \7178 , \7185 );
or \U$6819 ( \7196 , \7194 , \7195 );
and \U$6820 ( \7197 , \6172 , RIae76b68_57);
and \U$6821 ( \7198 , RIae78a58_123, \6170 );
nor \U$6822 ( \7199 , \7197 , \7198 );
and \U$6823 ( \7200 , \7199 , \6176 );
not \U$6824 ( \7201 , \7199 );
and \U$6825 ( \7202 , \7201 , \6175 );
nor \U$6826 ( \7203 , \7200 , \7202 );
nand \U$6827 ( \7204 , RIae7a240_174, RIae7a1c8_173);
and \U$6828 ( \7205 , \7204 , RIae7a2b8_175);
not \U$6829 ( \7206 , \7205 );
xor \U$6830 ( \7207 , \7203 , \7206 );
and \U$6831 ( \7208 , \6941 , RIae78cb0_128);
and \U$6832 ( \7209 , RIae78da0_130, \6939 );
nor \U$6833 ( \7210 , \7208 , \7209 );
and \U$6834 ( \7211 , \7210 , \6314 );
not \U$6835 ( \7212 , \7210 );
and \U$6836 ( \7213 , \7212 , \6945 );
nor \U$6837 ( \7214 , \7211 , \7213 );
and \U$6838 ( \7215 , \7207 , \7214 );
and \U$6839 ( \7216 , \7203 , \7206 );
or \U$6840 ( \7217 , \7215 , \7216 );
xor \U$6841 ( \7218 , \7196 , \7217 );
not \U$6842 ( \7219 , \3218 );
and \U$6843 ( \7220 , \3214 , RIae763e8_41);
and \U$6844 ( \7221 , RIae764d8_43, \3212 );
nor \U$6845 ( \7222 , \7220 , \7221 );
not \U$6846 ( \7223 , \7222 );
or \U$6847 ( \7224 , \7219 , \7223 );
or \U$6848 ( \7225 , \7222 , \2774 );
nand \U$6849 ( \7226 , \7224 , \7225 );
and \U$6850 ( \7227 , \3730 , RIae766b8_47);
and \U$6851 ( \7228 , RIae765c8_45, \3728 );
nor \U$6852 ( \7229 , \7227 , \7228 );
and \U$6853 ( \7230 , \7229 , \3732 );
not \U$6854 ( \7231 , \7229 );
and \U$6855 ( \7232 , \7231 , \3422 );
nor \U$6856 ( \7233 , \7230 , \7232 );
xor \U$6857 ( \7234 , \7226 , \7233 );
and \U$6858 ( \7235 , \4247 , RIae76118_35);
and \U$6859 ( \7236 , RIae76028_33, \4245 );
nor \U$6860 ( \7237 , \7235 , \7236 );
and \U$6861 ( \7238 , \7237 , \3989 );
not \U$6862 ( \7239 , \7237 );
and \U$6863 ( \7240 , \7239 , \4251 );
nor \U$6864 ( \7241 , \7238 , \7240 );
and \U$6865 ( \7242 , \7234 , \7241 );
and \U$6866 ( \7243 , \7226 , \7233 );
or \U$6867 ( \7244 , \7242 , \7243 );
and \U$6868 ( \7245 , \7218 , \7244 );
and \U$6869 ( \7246 , \7196 , \7217 );
or \U$6870 ( \7247 , \7245 , \7246 );
xor \U$6871 ( \7248 , \7171 , \7247 );
and \U$6872 ( \7249 , \558 , RIae78968_121);
and \U$6873 ( \7250 , RIae78878_119, \556 );
nor \U$6874 ( \7251 , \7249 , \7250 );
and \U$6875 ( \7252 , \7251 , \504 );
not \U$6876 ( \7253 , \7251 );
and \U$6877 ( \7254 , \7253 , \562 );
nor \U$6878 ( \7255 , \7252 , \7254 );
not \U$6879 ( \7256 , \402 );
and \U$6880 ( \7257 , \436 , RIae77c48_93);
and \U$6881 ( \7258 , RIae77b58_91, \434 );
nor \U$6882 ( \7259 , \7257 , \7258 );
not \U$6883 ( \7260 , \7259 );
or \U$6884 ( \7261 , \7256 , \7260 );
or \U$6885 ( \7262 , \7259 , \400 );
nand \U$6886 ( \7263 , \7261 , \7262 );
xor \U$6887 ( \7264 , \7255 , \7263 );
not \U$6888 ( \7265 , \471 );
and \U$6889 ( \7266 , \514 , RIae77d38_95);
and \U$6890 ( \7267 , RIae77e28_97, \512 );
nor \U$6891 ( \7268 , \7266 , \7267 );
not \U$6892 ( \7269 , \7268 );
or \U$6893 ( \7270 , \7265 , \7269 );
or \U$6894 ( \7271 , \7268 , \469 );
nand \U$6895 ( \7272 , \7270 , \7271 );
and \U$6896 ( \7273 , \7264 , \7272 );
and \U$6897 ( \7274 , \7255 , \7263 );
or \U$6898 ( \7275 , \7273 , \7274 );
nand \U$6899 ( \7276 , RIae783c8_109, RIae78b48_125);
xor \U$6900 ( \7277 , \7275 , \7276 );
and \U$6901 ( \7278 , \384 , RIae78530_112);
and \U$6902 ( \7279 , RIae77c48_93, \382 );
nor \U$6903 ( \7280 , \7278 , \7279 );
not \U$6904 ( \7281 , \7280 );
not \U$6905 ( \7282 , \388 );
and \U$6906 ( \7283 , \7281 , \7282 );
and \U$6907 ( \7284 , \7280 , \392 );
nor \U$6908 ( \7285 , \7283 , \7284 );
not \U$6909 ( \7286 , \7285 );
and \U$6910 ( \7287 , \436 , RIae77b58_91);
and \U$6911 ( \7288 , RIae77d38_95, \434 );
nor \U$6912 ( \7289 , \7287 , \7288 );
not \U$6913 ( \7290 , \7289 );
not \U$6914 ( \7291 , \402 );
and \U$6915 ( \7292 , \7290 , \7291 );
and \U$6916 ( \7293 , \7289 , \402 );
nor \U$6917 ( \7294 , \7292 , \7293 );
and \U$6918 ( \7295 , \514 , RIae77e28_97);
and \U$6919 ( \7296 , RIae78968_121, \512 );
nor \U$6920 ( \7297 , \7295 , \7296 );
not \U$6921 ( \7298 , \7297 );
not \U$6922 ( \7299 , \471 );
and \U$6923 ( \7300 , \7298 , \7299 );
and \U$6924 ( \7301 , \7297 , \469 );
nor \U$6925 ( \7302 , \7300 , \7301 );
xor \U$6926 ( \7303 , \7294 , \7302 );
not \U$6927 ( \7304 , \7303 );
or \U$6928 ( \7305 , \7286 , \7304 );
or \U$6929 ( \7306 , \7303 , \7285 );
nand \U$6930 ( \7307 , \7305 , \7306 );
and \U$6931 ( \7308 , \7277 , \7307 );
and \U$6932 ( \7309 , \7275 , \7276 );
or \U$6933 ( \7310 , \7308 , \7309 );
and \U$6934 ( \7311 , \7248 , \7310 );
and \U$6935 ( \7312 , \7171 , \7247 );
or \U$6936 ( \7313 , \7311 , \7312 );
and \U$6937 ( \7314 , \7090 , \7313 );
not \U$6938 ( \7315 , \7090 );
not \U$6939 ( \7316 , \7313 );
and \U$6940 ( \7317 , \7315 , \7316 );
nand \U$6941 ( \7318 , RIae78530_112, RIae78b48_125);
xor \U$6942 ( \7319 , \7276 , \7318 );
not \U$6943 ( \7320 , \7285 );
not \U$6944 ( \7321 , \7302 );
and \U$6945 ( \7322 , \7320 , \7321 );
and \U$6946 ( \7323 , \7302 , \7285 );
nor \U$6947 ( \7324 , \7323 , \7294 );
nor \U$6948 ( \7325 , \7322 , \7324 );
xor \U$6949 ( \7326 , \7319 , \7325 );
xor \U$6950 ( \7327 , \6362 , \6370 );
xor \U$6951 ( \7328 , \7327 , \6379 );
xor \U$6952 ( \7329 , \6443 , \6451 );
xor \U$6953 ( \7330 , \7329 , \6459 );
xor \U$6954 ( \7331 , \7328 , \7330 );
not \U$6955 ( \7332 , \6477 );
not \U$6956 ( \7333 , \6488 );
or \U$6957 ( \7334 , \7332 , \7333 );
or \U$6958 ( \7335 , \6477 , \6488 );
nand \U$6959 ( \7336 , \7334 , \7335 );
not \U$6960 ( \7337 , \7336 );
not \U$6961 ( \7338 , \6470 );
and \U$6962 ( \7339 , \7337 , \7338 );
and \U$6963 ( \7340 , \7336 , \6470 );
nor \U$6964 ( \7341 , \7339 , \7340 );
xor \U$6965 ( \7342 , \7331 , \7341 );
and \U$6966 ( \7343 , \7326 , \7342 );
xor \U$6967 ( \7344 , \6333 , \6340 );
xor \U$6968 ( \7345 , \7344 , \6348 );
xor \U$6969 ( \7346 , \6418 , \6425 );
xor \U$6970 ( \7347 , \7346 , \6433 );
xor \U$6971 ( \7348 , \7345 , \7347 );
not \U$6972 ( \7349 , \6289 );
not \U$6973 ( \7350 , \6301 );
or \U$6974 ( \7351 , \7349 , \7350 );
or \U$6975 ( \7352 , \6289 , \6301 );
nand \U$6976 ( \7353 , \7351 , \7352 );
not \U$6977 ( \7354 , \7353 );
not \U$6978 ( \7355 , \6282 );
and \U$6979 ( \7356 , \7354 , \7355 );
and \U$6980 ( \7357 , \7353 , \6282 );
nor \U$6981 ( \7358 , \7356 , \7357 );
xor \U$6982 ( \7359 , \7348 , \7358 );
xor \U$6983 ( \7360 , \7328 , \7330 );
xor \U$6984 ( \7361 , \7360 , \7341 );
and \U$6985 ( \7362 , \7359 , \7361 );
and \U$6986 ( \7363 , \7326 , \7359 );
or \U$6987 ( \7364 , \7343 , \7362 , \7363 );
nor \U$6988 ( \7365 , \7317 , \7364 );
nor \U$6989 ( \7366 , \7314 , \7365 );
not \U$6990 ( \7367 , \6272 );
not \U$6991 ( \7368 , \6138 );
or \U$6992 ( \7369 , \7367 , \7368 );
or \U$6993 ( \7370 , \6138 , \6272 );
nand \U$6994 ( \7371 , \7369 , \7370 );
not \U$6995 ( \7372 , \7371 );
not \U$6996 ( \7373 , \6161 );
and \U$6997 ( \7374 , \7372 , \7373 );
and \U$6998 ( \7375 , \7371 , \6161 );
nor \U$6999 ( \7376 , \7374 , \7375 );
or \U$7000 ( \7377 , \7366 , \7376 );
not \U$7001 ( \7378 , \7376 );
not \U$7002 ( \7379 , \7366 );
or \U$7003 ( \7380 , \7378 , \7379 );
xor \U$7004 ( \7381 , \6204 , \6235 );
xor \U$7005 ( \7382 , \7381 , \6269 );
not \U$7006 ( \7383 , \7382 );
xor \U$7007 ( \7384 , \7328 , \7330 );
and \U$7008 ( \7385 , \7384 , \7341 );
and \U$7009 ( \7386 , \7328 , \7330 );
or \U$7010 ( \7387 , \7385 , \7386 );
xor \U$7011 ( \7388 , \7345 , \7347 );
and \U$7012 ( \7389 , \7388 , \7358 );
and \U$7013 ( \7390 , \7345 , \7347 );
or \U$7014 ( \7391 , \7389 , \7390 );
xor \U$7015 ( \7392 , \7387 , \7391 );
not \U$7016 ( \7393 , \7392 );
or \U$7017 ( \7394 , \7383 , \7393 );
or \U$7018 ( \7395 , \7392 , \7382 );
nand \U$7019 ( \7396 , \7394 , \7395 );
xor \U$7020 ( \7397 , \6303 , \6325 );
xor \U$7021 ( \7398 , \7397 , \6351 );
xor \U$7022 ( \7399 , \7396 , \7398 );
xor \U$7023 ( \7400 , \6436 , \6462 );
xor \U$7024 ( \7401 , \7400 , \6490 );
or \U$7025 ( \7402 , \6409 , \6382 );
nand \U$7026 ( \7403 , \7402 , \6410 );
xor \U$7027 ( \7404 , \6091 , \6098 );
xor \U$7028 ( \7405 , \7404 , \6106 );
xor \U$7029 ( \7406 , \6083 , \6132 );
xor \U$7030 ( \7407 , \7405 , \7406 );
xor \U$7031 ( \7408 , \7403 , \7407 );
xor \U$7032 ( \7409 , \7401 , \7408 );
and \U$7033 ( \7410 , \7399 , \7409 );
and \U$7034 ( \7411 , \7396 , \7398 );
or \U$7035 ( \7412 , \7410 , \7411 );
nand \U$7036 ( \7413 , \7380 , \7412 );
nand \U$7037 ( \7414 , \7377 , \7413 );
xor \U$7038 ( \7415 , \6274 , \6496 );
xor \U$7039 ( \7416 , \7415 , \6645 );
xor \U$7040 ( \7417 , \7414 , \7416 );
xor \U$7041 ( \7418 , \6354 , \6410 );
xor \U$7042 ( \7419 , \7418 , \6493 );
not \U$7043 ( \7420 , \7419 );
xor \U$7044 ( \7421 , \6699 , \6703 );
xor \U$7045 ( \7422 , \7421 , \6708 );
xor \U$7046 ( \7423 , \6717 , \6723 );
xor \U$7047 ( \7424 , \7423 , \6730 );
xor \U$7048 ( \7425 , \6533 , \6539 );
xor \U$7049 ( \7426 , \7425 , \6564 );
xor \U$7050 ( \7427 , \6513 , \6640 );
xor \U$7051 ( \7428 , \7426 , \7427 );
xor \U$7052 ( \7429 , \7424 , \7428 );
xor \U$7053 ( \7430 , \7422 , \7429 );
not \U$7054 ( \7431 , \7430 );
or \U$7055 ( \7432 , \7420 , \7431 );
or \U$7056 ( \7433 , \7430 , \7419 );
xor \U$7057 ( \7434 , \6987 , \6995 );
and \U$7058 ( \7435 , \7434 , \7004 );
and \U$7059 ( \7436 , \6987 , \6995 );
or \U$7060 ( \7437 , \7435 , \7436 );
xor \U$7061 ( \7438 , \6933 , \6947 );
and \U$7062 ( \7439 , \7438 , \6955 );
and \U$7063 ( \7440 , \6933 , \6947 );
or \U$7064 ( \7441 , \7439 , \7440 );
xor \U$7065 ( \7442 , \7437 , \7441 );
xor \U$7066 ( \7443 , \6963 , \6970 );
and \U$7067 ( \7444 , \7443 , \6978 );
and \U$7068 ( \7445 , \6963 , \6970 );
or \U$7069 ( \7446 , \7444 , \7445 );
and \U$7070 ( \7447 , \7442 , \7446 );
and \U$7071 ( \7448 , \7437 , \7441 );
nor \U$7072 ( \7449 , \7447 , \7448 );
xor \U$7073 ( \7450 , \7276 , \7318 );
and \U$7074 ( \7451 , \7450 , \7325 );
and \U$7075 ( \7452 , \7276 , \7318 );
or \U$7076 ( \7453 , \7451 , \7452 );
xor \U$7077 ( \7454 , \7449 , \7453 );
xor \U$7078 ( \7455 , \7044 , \7051 );
and \U$7079 ( \7456 , \7455 , \7059 );
and \U$7080 ( \7457 , \7044 , \7051 );
or \U$7081 ( \7458 , \7456 , \7457 );
xor \U$7082 ( \7459 , \7021 , \7028 );
and \U$7083 ( \7460 , \7459 , \7036 );
and \U$7084 ( \7461 , \7021 , \7028 );
or \U$7085 ( \7462 , \7460 , \7461 );
xor \U$7086 ( \7463 , \7458 , \7462 );
xor \U$7087 ( \7464 , \7068 , \7075 );
and \U$7088 ( \7465 , \7464 , \7083 );
and \U$7089 ( \7466 , \7068 , \7075 );
or \U$7090 ( \7467 , \7465 , \7466 );
and \U$7091 ( \7468 , \7463 , \7467 );
and \U$7092 ( \7469 , \7458 , \7462 );
nor \U$7093 ( \7470 , \7468 , \7469 );
and \U$7094 ( \7471 , \7454 , \7470 );
and \U$7095 ( \7472 , \7449 , \7453 );
or \U$7096 ( \7473 , \7471 , \7472 );
not \U$7097 ( \7474 , \7382 );
not \U$7098 ( \7475 , \7391 );
and \U$7099 ( \7476 , \7474 , \7475 );
and \U$7100 ( \7477 , \7382 , \7391 );
nor \U$7101 ( \7478 , \7477 , \7387 );
nor \U$7102 ( \7479 , \7476 , \7478 );
xnor \U$7103 ( \7480 , \7473 , \7479 );
not \U$7104 ( \7481 , \7480 );
xor \U$7105 ( \7482 , \6436 , \6462 );
xor \U$7106 ( \7483 , \7482 , \6490 );
and \U$7107 ( \7484 , \7403 , \7483 );
xor \U$7108 ( \7485 , \6436 , \6462 );
xor \U$7109 ( \7486 , \7485 , \6490 );
and \U$7110 ( \7487 , \7407 , \7486 );
and \U$7111 ( \7488 , \7403 , \7407 );
or \U$7112 ( \7489 , \7484 , \7487 , \7488 );
not \U$7113 ( \7490 , \7489 );
and \U$7114 ( \7491 , \7481 , \7490 );
and \U$7115 ( \7492 , \7480 , \7489 );
nor \U$7116 ( \7493 , \7491 , \7492 );
not \U$7117 ( \7494 , \7493 );
nand \U$7118 ( \7495 , \7433 , \7494 );
nand \U$7119 ( \7496 , \7432 , \7495 );
and \U$7120 ( \7497 , \7417 , \7496 );
and \U$7121 ( \7498 , \7414 , \7416 );
or \U$7122 ( \7499 , \7497 , \7498 );
or \U$7123 ( \7500 , \7479 , \7473 );
not \U$7124 ( \7501 , \7473 );
not \U$7125 ( \7502 , \7479 );
or \U$7126 ( \7503 , \7501 , \7502 );
nand \U$7127 ( \7504 , \7503 , \7489 );
nand \U$7128 ( \7505 , \7500 , \7504 );
xor \U$7129 ( \7506 , \6699 , \6703 );
xor \U$7130 ( \7507 , \7506 , \6708 );
and \U$7131 ( \7508 , \7424 , \7507 );
xor \U$7132 ( \7509 , \6699 , \6703 );
xor \U$7133 ( \7510 , \7509 , \6708 );
and \U$7134 ( \7511 , \7428 , \7510 );
and \U$7135 ( \7512 , \7424 , \7428 );
or \U$7136 ( \7513 , \7508 , \7511 , \7512 );
xor \U$7137 ( \7514 , \7505 , \7513 );
xor \U$7138 ( \7515 , \6741 , \6743 );
xor \U$7139 ( \7516 , \7515 , \6746 );
xor \U$7140 ( \7517 , \6739 , \6771 );
xor \U$7141 ( \7518 , \7516 , \7517 );
and \U$7142 ( \7519 , \7514 , \7518 );
and \U$7143 ( \7520 , \7505 , \7513 );
or \U$7144 ( \7521 , \7519 , \7520 );
xor \U$7145 ( \7522 , \6793 , \6822 );
xor \U$7146 ( \7523 , \7521 , \7522 );
xor \U$7147 ( \7524 , \6648 , \6694 );
xor \U$7148 ( \7525 , \7524 , \6776 );
xor \U$7149 ( \7526 , \7523 , \7525 );
and \U$7150 ( \7527 , \7499 , \7526 );
xor \U$7151 ( \7528 , \7505 , \7513 );
xor \U$7152 ( \7529 , \7528 , \7518 );
not \U$7153 ( \7530 , \7529 );
xor \U$7154 ( \7531 , \7414 , \7416 );
xor \U$7155 ( \7532 , \7531 , \7496 );
not \U$7156 ( \7533 , \7532 );
or \U$7157 ( \7534 , \7530 , \7533 );
or \U$7158 ( \7535 , \7532 , \7529 );
not \U$7159 ( \7536 , \7366 );
not \U$7160 ( \7537 , \7412 );
or \U$7161 ( \7538 , \7536 , \7537 );
or \U$7162 ( \7539 , \7412 , \7366 );
nand \U$7163 ( \7540 , \7538 , \7539 );
not \U$7164 ( \7541 , \7540 );
not \U$7165 ( \7542 , \7376 );
and \U$7166 ( \7543 , \7541 , \7542 );
and \U$7167 ( \7544 , \7540 , \7376 );
nor \U$7168 ( \7545 , \7543 , \7544 );
xor \U$7169 ( \7546 , \7458 , \7462 );
xor \U$7170 ( \7547 , \7546 , \7467 );
xor \U$7171 ( \7548 , \7437 , \7441 );
xor \U$7172 ( \7549 , \7548 , \7446 );
and \U$7173 ( \7550 , \7547 , \7549 );
not \U$7174 ( \7551 , \7549 );
not \U$7175 ( \7552 , \7547 );
and \U$7176 ( \7553 , \7551 , \7552 );
xor \U$7177 ( \7554 , \7328 , \7330 );
xor \U$7178 ( \7555 , \7554 , \7341 );
xor \U$7179 ( \7556 , \7326 , \7359 );
xor \U$7180 ( \7557 , \7555 , \7556 );
nor \U$7181 ( \7558 , \7553 , \7557 );
nor \U$7182 ( \7559 , \7550 , \7558 );
xor \U$7183 ( \7560 , \7449 , \7453 );
xor \U$7184 ( \7561 , \7560 , \7470 );
xor \U$7185 ( \7562 , \7559 , \7561 );
xor \U$7186 ( \7563 , \7150 , \7157 );
xor \U$7187 ( \7564 , \7563 , \7165 );
xor \U$7188 ( \7565 , \7097 , \7104 );
xor \U$7189 ( \7566 , \7565 , \7112 );
and \U$7190 ( \7567 , \7564 , \7566 );
xor \U$7191 ( \7568 , \7226 , \7233 );
xor \U$7192 ( \7569 , \7568 , \7241 );
xor \U$7193 ( \7570 , \7097 , \7104 );
xor \U$7194 ( \7571 , \7570 , \7112 );
and \U$7195 ( \7572 , \7569 , \7571 );
and \U$7196 ( \7573 , \7564 , \7569 );
or \U$7197 ( \7574 , \7567 , \7572 , \7573 );
xor \U$7198 ( \7575 , \7123 , \7130 );
xor \U$7199 ( \7576 , \7575 , \7138 );
not \U$7200 ( \7577 , RIae785a8_113);
nor \U$7201 ( \7578 , \7577 , \491 );
xor \U$7202 ( \7579 , \7576 , \7578 );
xor \U$7203 ( \7580 , \7255 , \7263 );
xor \U$7204 ( \7581 , \7580 , \7272 );
and \U$7205 ( \7582 , \7579 , \7581 );
and \U$7206 ( \7583 , \7576 , \7578 );
or \U$7207 ( \7584 , \7582 , \7583 );
xor \U$7208 ( \7585 , \7574 , \7584 );
xor \U$7209 ( \7586 , \6963 , \6970 );
xor \U$7210 ( \7587 , \7586 , \6978 );
xor \U$7211 ( \7588 , \6956 , \7005 );
xor \U$7212 ( \7589 , \7587 , \7588 );
and \U$7213 ( \7590 , \7585 , \7589 );
and \U$7214 ( \7591 , \7574 , \7584 );
or \U$7215 ( \7592 , \7590 , \7591 );
and \U$7216 ( \7593 , \3730 , RIae764d8_43);
and \U$7217 ( \7594 , RIae766b8_47, \3728 );
nor \U$7218 ( \7595 , \7593 , \7594 );
and \U$7219 ( \7596 , \7595 , \3732 );
not \U$7220 ( \7597 , \7595 );
and \U$7221 ( \7598 , \7597 , \3422 );
nor \U$7222 ( \7599 , \7596 , \7598 );
not \U$7223 ( \7600 , \2774 );
and \U$7224 ( \7601 , \3214 , RIae753f8_7);
and \U$7225 ( \7602 , RIae763e8_41, \3212 );
nor \U$7226 ( \7603 , \7601 , \7602 );
not \U$7227 ( \7604 , \7603 );
or \U$7228 ( \7605 , \7600 , \7604 );
or \U$7229 ( \7606 , \7603 , \2774 );
nand \U$7230 ( \7607 , \7605 , \7606 );
xor \U$7231 ( \7608 , \7599 , \7607 );
and \U$7232 ( \7609 , \4247 , RIae765c8_45);
and \U$7233 ( \7610 , RIae76118_35, \4245 );
nor \U$7234 ( \7611 , \7609 , \7610 );
and \U$7235 ( \7612 , \7611 , \3989 );
not \U$7236 ( \7613 , \7611 );
and \U$7237 ( \7614 , \7613 , \4251 );
nor \U$7238 ( \7615 , \7612 , \7614 );
and \U$7239 ( \7616 , \7608 , \7615 );
and \U$7240 ( \7617 , \7599 , \7607 );
or \U$7241 ( \7618 , \7616 , \7617 );
and \U$7242 ( \7619 , \6172 , RIae76898_51);
and \U$7243 ( \7620 , RIae76b68_57, \6170 );
nor \U$7244 ( \7621 , \7619 , \7620 );
and \U$7245 ( \7622 , \7621 , \6176 );
not \U$7246 ( \7623 , \7621 );
and \U$7247 ( \7624 , \7623 , \6175 );
nor \U$7248 ( \7625 , \7622 , \7624 );
and \U$7249 ( \7626 , RIae7a2b8_175, RIae7a1c8_173);
not \U$7250 ( \7627 , RIae7a1c8_173);
nor \U$7251 ( \7628 , \7627 , RIae7a240_174);
not \U$7252 ( \7629 , RIae7a240_174);
nor \U$7253 ( \7630 , \7629 , RIae7a1c8_173);
or \U$7254 ( \7631 , \7628 , \7630 );
nor \U$7255 ( \7632 , RIae7a2b8_175, RIae7a1c8_173);
nor \U$7256 ( \7633 , \7626 , \7631 , \7632 );
nand \U$7257 ( \7634 , RIae78da0_130, \7633 );
and \U$7258 ( \7635 , \7634 , \7206 );
not \U$7259 ( \7636 , \7634 );
and \U$7260 ( \7637 , \7636 , \7205 );
nor \U$7261 ( \7638 , \7635 , \7637 );
xor \U$7262 ( \7639 , \7625 , \7638 );
and \U$7263 ( \7640 , \6941 , RIae78a58_123);
and \U$7264 ( \7641 , RIae78cb0_128, \6939 );
nor \U$7265 ( \7642 , \7640 , \7641 );
and \U$7266 ( \7643 , \7642 , \6314 );
not \U$7267 ( \7644 , \7642 );
and \U$7268 ( \7645 , \7644 , \6945 );
nor \U$7269 ( \7646 , \7643 , \7645 );
and \U$7270 ( \7647 , \7639 , \7646 );
and \U$7271 ( \7648 , \7625 , \7638 );
or \U$7272 ( \7649 , \7647 , \7648 );
xor \U$7273 ( \7650 , \7618 , \7649 );
and \U$7274 ( \7651 , \5896 , RIae76988_53);
and \U$7275 ( \7652 , RIae767a8_49, \5894 );
nor \U$7276 ( \7653 , \7651 , \7652 );
and \U$7277 ( \7654 , \7653 , \5590 );
not \U$7278 ( \7655 , \7653 );
and \U$7279 ( \7656 , \7655 , \5589 );
nor \U$7280 ( \7657 , \7654 , \7656 );
and \U$7281 ( \7658 , \4688 , RIae76028_33);
and \U$7282 ( \7659 , RIae762f8_39, \4686 );
nor \U$7283 ( \7660 , \7658 , \7659 );
and \U$7284 ( \7661 , \7660 , \4481 );
not \U$7285 ( \7662 , \7660 );
and \U$7286 ( \7663 , \7662 , \4482 );
nor \U$7287 ( \7664 , \7661 , \7663 );
xor \U$7288 ( \7665 , \7657 , \7664 );
and \U$7289 ( \7666 , \5399 , RIae76208_37);
and \U$7290 ( \7667 , RIae76a78_55, \5397 );
nor \U$7291 ( \7668 , \7666 , \7667 );
and \U$7292 ( \7669 , \7668 , \5016 );
not \U$7293 ( \7670 , \7668 );
and \U$7294 ( \7671 , \7670 , \5403 );
nor \U$7295 ( \7672 , \7669 , \7671 );
and \U$7296 ( \7673 , \7665 , \7672 );
and \U$7297 ( \7674 , \7657 , \7664 );
or \U$7298 ( \7675 , \7673 , \7674 );
and \U$7299 ( \7676 , \7650 , \7675 );
and \U$7300 ( \7677 , \7618 , \7649 );
or \U$7301 ( \7678 , \7676 , \7677 );
nand \U$7302 ( \7679 , RIae781e8_105, RIae78b48_125);
and \U$7303 ( \7680 , \384 , RIae785a8_113);
and \U$7304 ( \7681 , RIae783c8_109, \382 );
nor \U$7305 ( \7682 , \7680 , \7681 );
not \U$7306 ( \7683 , \7682 );
not \U$7307 ( \7684 , \392 );
and \U$7308 ( \7685 , \7683 , \7684 );
and \U$7309 ( \7686 , \7682 , \388 );
nor \U$7310 ( \7687 , \7685 , \7686 );
nand \U$7311 ( \7688 , \7679 , \7687 );
not \U$7312 ( \7689 , \392 );
and \U$7313 ( \7690 , \384 , RIae783c8_109);
and \U$7314 ( \7691 , RIae78530_112, \382 );
nor \U$7315 ( \7692 , \7690 , \7691 );
not \U$7316 ( \7693 , \7692 );
or \U$7317 ( \7694 , \7689 , \7693 );
or \U$7318 ( \7695 , \7692 , \392 );
nand \U$7319 ( \7696 , \7694 , \7695 );
xor \U$7320 ( \7697 , \7688 , \7696 );
and \U$7321 ( \7698 , \558 , RIae77e28_97);
and \U$7322 ( \7699 , RIae78968_121, \556 );
nor \U$7323 ( \7700 , \7698 , \7699 );
and \U$7324 ( \7701 , \7700 , \504 );
not \U$7325 ( \7702 , \7700 );
and \U$7326 ( \7703 , \7702 , \562 );
nor \U$7327 ( \7704 , \7701 , \7703 );
not \U$7328 ( \7705 , \402 );
and \U$7329 ( \7706 , \436 , RIae78530_112);
and \U$7330 ( \7707 , RIae77c48_93, \434 );
nor \U$7331 ( \7708 , \7706 , \7707 );
not \U$7332 ( \7709 , \7708 );
or \U$7333 ( \7710 , \7705 , \7709 );
or \U$7334 ( \7711 , \7708 , \400 );
nand \U$7335 ( \7712 , \7710 , \7711 );
xor \U$7336 ( \7713 , \7704 , \7712 );
not \U$7337 ( \7714 , \471 );
and \U$7338 ( \7715 , \514 , RIae77b58_91);
and \U$7339 ( \7716 , RIae77d38_95, \512 );
nor \U$7340 ( \7717 , \7715 , \7716 );
not \U$7341 ( \7718 , \7717 );
or \U$7342 ( \7719 , \7714 , \7718 );
or \U$7343 ( \7720 , \7717 , \471 );
nand \U$7344 ( \7721 , \7719 , \7720 );
and \U$7345 ( \7722 , \7713 , \7721 );
and \U$7346 ( \7723 , \7704 , \7712 );
or \U$7347 ( \7724 , \7722 , \7723 );
and \U$7348 ( \7725 , \7697 , \7724 );
and \U$7349 ( \7726 , \7688 , \7696 );
or \U$7350 ( \7727 , \7725 , \7726 );
xor \U$7351 ( \7728 , \7678 , \7727 );
and \U$7352 ( \7729 , \2607 , RIae756c8_13);
and \U$7353 ( \7730 , RIae75218_3, \2605 );
nor \U$7354 ( \7731 , \7729 , \7730 );
and \U$7355 ( \7732 , \7731 , \2611 );
not \U$7356 ( \7733 , \7731 );
and \U$7357 ( \7734 , \7733 , \2397 );
nor \U$7358 ( \7735 , \7732 , \7734 );
and \U$7359 ( \7736 , \2224 , RIae754e8_9);
and \U$7360 ( \7737 , RIae757b8_15, \2222 );
nor \U$7361 ( \7738 , \7736 , \7737 );
and \U$7362 ( \7739 , \7738 , \2061 );
not \U$7363 ( \7740 , \7738 );
and \U$7364 ( \7741 , \7740 , \2060 );
nor \U$7365 ( \7742 , \7739 , \7741 );
xor \U$7366 ( \7743 , \7735 , \7742 );
not \U$7367 ( \7744 , \2789 );
and \U$7368 ( \7745 , \2783 , RIae75128_1);
and \U$7369 ( \7746 , RIae75308_5, \2781 );
nor \U$7370 ( \7747 , \7745 , \7746 );
not \U$7371 ( \7748 , \7747 );
or \U$7372 ( \7749 , \7744 , \7748 );
or \U$7373 ( \7750 , \7747 , \3089 );
nand \U$7374 ( \7751 , \7749 , \7750 );
and \U$7375 ( \7752 , \7743 , \7751 );
and \U$7376 ( \7753 , \7735 , \7742 );
or \U$7377 ( \7754 , \7752 , \7753 );
and \U$7378 ( \7755 , \1593 , RIae75e48_29);
and \U$7379 ( \7756 , RIae75c68_25, \1591 );
nor \U$7380 ( \7757 , \7755 , \7756 );
and \U$7381 ( \7758 , \7757 , \1498 );
not \U$7382 ( \7759 , \7757 );
and \U$7383 ( \7760 , \7759 , \1488 );
nor \U$7384 ( \7761 , \7758 , \7760 );
and \U$7385 ( \7762 , \1376 , RIae758a8_17);
and \U$7386 ( \7763 , RIae75f38_31, \1374 );
nor \U$7387 ( \7764 , \7762 , \7763 );
and \U$7388 ( \7765 , \7764 , \1380 );
not \U$7389 ( \7766 , \7764 );
and \U$7390 ( \7767 , \7766 , \1261 );
nor \U$7391 ( \7768 , \7765 , \7767 );
xor \U$7392 ( \7769 , \7761 , \7768 );
and \U$7393 ( \7770 , \1939 , RIae75d58_27);
and \U$7394 ( \7771 , RIae755d8_11, \1937 );
nor \U$7395 ( \7772 , \7770 , \7771 );
and \U$7396 ( \7773 , \7772 , \1735 );
not \U$7397 ( \7774 , \7772 );
and \U$7398 ( \7775 , \7774 , \1734 );
nor \U$7399 ( \7776 , \7773 , \7775 );
and \U$7400 ( \7777 , \7769 , \7776 );
and \U$7401 ( \7778 , \7761 , \7768 );
or \U$7402 ( \7779 , \7777 , \7778 );
xor \U$7403 ( \7780 , \7754 , \7779 );
and \U$7404 ( \7781 , \672 , RIae78878_119);
and \U$7405 ( \7782 , RIae78788_117, \670 );
nor \U$7406 ( \7783 , \7781 , \7782 );
and \U$7407 ( \7784 , \7783 , \588 );
not \U$7408 ( \7785 , \7783 );
and \U$7409 ( \7786 , \7785 , \587 );
nor \U$7410 ( \7787 , \7784 , \7786 );
not \U$7411 ( \7788 , \789 );
and \U$7412 ( \7789 , \883 , RIae78698_115);
and \U$7413 ( \7790 , RIae75b78_23, \881 );
nor \U$7414 ( \7791 , \7789 , \7790 );
not \U$7415 ( \7792 , \7791 );
or \U$7416 ( \7793 , \7788 , \7792 );
or \U$7417 ( \7794 , \7791 , \789 );
nand \U$7418 ( \7795 , \7793 , \7794 );
xor \U$7419 ( \7796 , \7787 , \7795 );
and \U$7420 ( \7797 , \1138 , RIae75a88_21);
and \U$7421 ( \7798 , RIae75998_19, \1136 );
nor \U$7422 ( \7799 , \7797 , \7798 );
and \U$7423 ( \7800 , \7799 , \1012 );
not \U$7424 ( \7801 , \7799 );
and \U$7425 ( \7802 , \7801 , \1142 );
nor \U$7426 ( \7803 , \7800 , \7802 );
and \U$7427 ( \7804 , \7796 , \7803 );
and \U$7428 ( \7805 , \7787 , \7795 );
or \U$7429 ( \7806 , \7804 , \7805 );
and \U$7430 ( \7807 , \7780 , \7806 );
and \U$7431 ( \7808 , \7754 , \7779 );
or \U$7432 ( \7809 , \7807 , \7808 );
and \U$7433 ( \7810 , \7728 , \7809 );
and \U$7434 ( \7811 , \7678 , \7727 );
or \U$7435 ( \7812 , \7810 , \7811 );
xor \U$7436 ( \7813 , \7592 , \7812 );
xor \U$7437 ( \7814 , \7115 , \7141 );
xor \U$7438 ( \7815 , \7814 , \7168 );
xor \U$7439 ( \7816 , \7037 , \7060 );
xor \U$7440 ( \7817 , \7816 , \7084 );
and \U$7441 ( \7818 , \7815 , \7817 );
xor \U$7442 ( \7819 , \7275 , \7276 );
xor \U$7443 ( \7820 , \7819 , \7307 );
xor \U$7444 ( \7821 , \7037 , \7060 );
xor \U$7445 ( \7822 , \7821 , \7084 );
and \U$7446 ( \7823 , \7820 , \7822 );
and \U$7447 ( \7824 , \7815 , \7820 );
or \U$7448 ( \7825 , \7818 , \7823 , \7824 );
and \U$7449 ( \7826 , \7813 , \7825 );
and \U$7450 ( \7827 , \7592 , \7812 );
nor \U$7451 ( \7828 , \7826 , \7827 );
and \U$7452 ( \7829 , \7562 , \7828 );
and \U$7453 ( \7830 , \7559 , \7561 );
or \U$7454 ( \7831 , \7829 , \7830 );
xor \U$7455 ( \7832 , \7545 , \7831 );
not \U$7456 ( \7833 , \7493 );
not \U$7457 ( \7834 , \7419 );
and \U$7458 ( \7835 , \7833 , \7834 );
and \U$7459 ( \7836 , \7493 , \7419 );
nor \U$7460 ( \7837 , \7835 , \7836 );
not \U$7461 ( \7838 , \7837 );
not \U$7462 ( \7839 , \7430 );
and \U$7463 ( \7840 , \7838 , \7839 );
and \U$7464 ( \7841 , \7837 , \7430 );
nor \U$7465 ( \7842 , \7840 , \7841 );
and \U$7466 ( \7843 , \7832 , \7842 );
and \U$7467 ( \7844 , \7545 , \7831 );
or \U$7468 ( \7845 , \7843 , \7844 );
not \U$7469 ( \7846 , \7845 );
nand \U$7470 ( \7847 , \7535 , \7846 );
nand \U$7471 ( \7848 , \7534 , \7847 );
xor \U$7472 ( \7849 , \7521 , \7522 );
xor \U$7473 ( \7850 , \7849 , \7525 );
and \U$7474 ( \7851 , \7848 , \7850 );
and \U$7475 ( \7852 , \7499 , \7848 );
or \U$7476 ( \7853 , \7527 , \7851 , \7852 );
xor \U$7477 ( \7854 , \7521 , \7522 );
and \U$7478 ( \7855 , \7854 , \7525 );
and \U$7479 ( \7856 , \7521 , \7522 );
or \U$7480 ( \7857 , \7855 , \7856 );
xor \U$7481 ( \7858 , \6887 , \6889 );
xor \U$7482 ( \7859 , \7858 , \6898 );
xor \U$7483 ( \7860 , \7857 , \7859 );
xor \U$7484 ( \7861 , \6779 , \6823 );
xor \U$7485 ( \7862 , \7861 , \6854 );
xor \U$7486 ( \7863 , \7860 , \7862 );
and \U$7487 ( \7864 , \7853 , \7863 );
xor \U$7488 ( \7865 , \7863 , \7853 );
xor \U$7489 ( \7866 , \7521 , \7522 );
xor \U$7490 ( \7867 , \7866 , \7525 );
xor \U$7491 ( \7868 , \7499 , \7848 );
xor \U$7492 ( \7869 , \7867 , \7868 );
xor \U$7493 ( \7870 , \7545 , \7831 );
xor \U$7494 ( \7871 , \7870 , \7842 );
xor \U$7495 ( \7872 , \7559 , \7561 );
xor \U$7496 ( \7873 , \7872 , \7828 );
not \U$7497 ( \7874 , \7873 );
not \U$7498 ( \7875 , \7364 );
xor \U$7499 ( \7876 , \7313 , \7090 );
not \U$7500 ( \7877 , \7876 );
or \U$7501 ( \7878 , \7875 , \7877 );
or \U$7502 ( \7879 , \7876 , \7364 );
nand \U$7503 ( \7880 , \7878 , \7879 );
nand \U$7504 ( \7881 , \7874 , \7880 );
or \U$7505 ( \7882 , \7871 , \7881 );
not \U$7506 ( \7883 , \7881 );
not \U$7507 ( \7884 , \7871 );
or \U$7508 ( \7885 , \7883 , \7884 );
xor \U$7509 ( \7886 , \7547 , \7549 );
not \U$7510 ( \7887 , \7886 );
not \U$7511 ( \7888 , \7557 );
or \U$7512 ( \7889 , \7887 , \7888 );
or \U$7513 ( \7890 , \7557 , \7886 );
nand \U$7514 ( \7891 , \7889 , \7890 );
xor \U$7515 ( \7892 , \7171 , \7247 );
xor \U$7516 ( \7893 , \7892 , \7310 );
xor \U$7517 ( \7894 , \7891 , \7893 );
xor \U$7518 ( \7895 , \7592 , \7812 );
xor \U$7519 ( \7896 , \7895 , \7825 );
and \U$7520 ( \7897 , \7894 , \7896 );
and \U$7521 ( \7898 , \7891 , \7893 );
or \U$7522 ( \7899 , \7897 , \7898 );
xor \U$7523 ( \7900 , \7396 , \7398 );
xor \U$7524 ( \7901 , \7900 , \7409 );
xor \U$7525 ( \7902 , \7899 , \7901 );
xor \U$7526 ( \7903 , \7735 , \7742 );
xor \U$7527 ( \7904 , \7903 , \7751 );
xor \U$7528 ( \7905 , \7657 , \7664 );
xor \U$7529 ( \7906 , \7905 , \7672 );
and \U$7530 ( \7907 , \7904 , \7906 );
xor \U$7531 ( \7908 , \7599 , \7607 );
xor \U$7532 ( \7909 , \7908 , \7615 );
xor \U$7533 ( \7910 , \7657 , \7664 );
xor \U$7534 ( \7911 , \7910 , \7672 );
and \U$7535 ( \7912 , \7909 , \7911 );
and \U$7536 ( \7913 , \7904 , \7909 );
or \U$7537 ( \7914 , \7907 , \7912 , \7913 );
xor \U$7538 ( \7915 , \7178 , \7185 );
xor \U$7539 ( \7916 , \7915 , \7193 );
xor \U$7540 ( \7917 , \7914 , \7916 );
xor \U$7541 ( \7918 , \7761 , \7768 );
xor \U$7542 ( \7919 , \7918 , \7776 );
xor \U$7543 ( \7920 , \7704 , \7712 );
xor \U$7544 ( \7921 , \7920 , \7721 );
xor \U$7545 ( \7922 , \7919 , \7921 );
xor \U$7546 ( \7923 , \7787 , \7795 );
xor \U$7547 ( \7924 , \7923 , \7803 );
and \U$7548 ( \7925 , \7922 , \7924 );
and \U$7549 ( \7926 , \7919 , \7921 );
or \U$7550 ( \7927 , \7925 , \7926 );
and \U$7551 ( \7928 , \7917 , \7927 );
and \U$7552 ( \7929 , \7914 , \7916 );
or \U$7553 ( \7930 , \7928 , \7929 );
and \U$7554 ( \7931 , \436 , RIae783c8_109);
and \U$7555 ( \7932 , RIae78530_112, \434 );
nor \U$7556 ( \7933 , \7931 , \7932 );
not \U$7557 ( \7934 , \7933 );
not \U$7558 ( \7935 , \400 );
and \U$7559 ( \7936 , \7934 , \7935 );
and \U$7560 ( \7937 , \7933 , \402 );
nor \U$7561 ( \7938 , \7936 , \7937 );
nand \U$7562 ( \7939 , RIae78008_101, RIae78b48_125);
or \U$7563 ( \7940 , \7938 , \7939 );
not \U$7564 ( \7941 , \7939 );
not \U$7565 ( \7942 , \7938 );
or \U$7566 ( \7943 , \7941 , \7942 );
not \U$7567 ( \7944 , \388 );
and \U$7568 ( \7945 , \384 , RIae781e8_105);
and \U$7569 ( \7946 , RIae785a8_113, \382 );
nor \U$7570 ( \7947 , \7945 , \7946 );
not \U$7571 ( \7948 , \7947 );
or \U$7572 ( \7949 , \7944 , \7948 );
or \U$7573 ( \7950 , \7947 , \392 );
nand \U$7574 ( \7951 , \7949 , \7950 );
nand \U$7575 ( \7952 , \7943 , \7951 );
nand \U$7576 ( \7953 , \7940 , \7952 );
or \U$7577 ( \7954 , \7687 , \7679 );
nand \U$7578 ( \7955 , \7954 , \7688 );
xor \U$7579 ( \7956 , \7953 , \7955 );
and \U$7580 ( \7957 , \672 , RIae78968_121);
and \U$7581 ( \7958 , RIae78878_119, \670 );
nor \U$7582 ( \7959 , \7957 , \7958 );
and \U$7583 ( \7960 , \7959 , \588 );
not \U$7584 ( \7961 , \7959 );
and \U$7585 ( \7962 , \7961 , \587 );
nor \U$7586 ( \7963 , \7960 , \7962 );
not \U$7587 ( \7964 , \469 );
and \U$7588 ( \7965 , \514 , RIae77c48_93);
and \U$7589 ( \7966 , RIae77b58_91, \512 );
nor \U$7590 ( \7967 , \7965 , \7966 );
not \U$7591 ( \7968 , \7967 );
or \U$7592 ( \7969 , \7964 , \7968 );
or \U$7593 ( \7970 , \7967 , \471 );
nand \U$7594 ( \7971 , \7969 , \7970 );
xor \U$7595 ( \7972 , \7963 , \7971 );
and \U$7596 ( \7973 , \558 , RIae77d38_95);
and \U$7597 ( \7974 , RIae77e28_97, \556 );
nor \U$7598 ( \7975 , \7973 , \7974 );
and \U$7599 ( \7976 , \7975 , \504 );
not \U$7600 ( \7977 , \7975 );
and \U$7601 ( \7978 , \7977 , \562 );
nor \U$7602 ( \7979 , \7976 , \7978 );
and \U$7603 ( \7980 , \7972 , \7979 );
and \U$7604 ( \7981 , \7963 , \7971 );
or \U$7605 ( \7982 , \7980 , \7981 );
and \U$7606 ( \7983 , \7956 , \7982 );
and \U$7607 ( \7984 , \7953 , \7955 );
or \U$7608 ( \7985 , \7983 , \7984 );
and \U$7609 ( \7986 , \6172 , RIae767a8_49);
and \U$7610 ( \7987 , RIae76898_51, \6170 );
nor \U$7611 ( \7988 , \7986 , \7987 );
and \U$7612 ( \7989 , \7988 , \6176 );
not \U$7613 ( \7990 , \7988 );
and \U$7614 ( \7991 , \7990 , \6175 );
nor \U$7615 ( \7992 , \7989 , \7991 );
and \U$7616 ( \7993 , \5399 , RIae762f8_39);
and \U$7617 ( \7994 , RIae76208_37, \5397 );
nor \U$7618 ( \7995 , \7993 , \7994 );
and \U$7619 ( \7996 , \7995 , \5016 );
not \U$7620 ( \7997 , \7995 );
and \U$7621 ( \7998 , \7997 , \5403 );
nor \U$7622 ( \7999 , \7996 , \7998 );
xor \U$7623 ( \8000 , \7992 , \7999 );
and \U$7624 ( \8001 , \5896 , RIae76a78_55);
and \U$7625 ( \8002 , RIae76988_53, \5894 );
nor \U$7626 ( \8003 , \8001 , \8002 );
and \U$7627 ( \8004 , \8003 , \5590 );
not \U$7628 ( \8005 , \8003 );
and \U$7629 ( \8006 , \8005 , \5589 );
nor \U$7630 ( \8007 , \8004 , \8006 );
and \U$7631 ( \8008 , \8000 , \8007 );
and \U$7632 ( \8009 , \7992 , \7999 );
or \U$7633 ( \8010 , \8008 , \8009 );
and \U$7634 ( \8011 , \7633 , RIae78cb0_128);
and \U$7635 ( \8012 , RIae78da0_130, \7631 );
nor \U$7636 ( \8013 , \8011 , \8012 );
and \U$7637 ( \8014 , \8013 , \7206 );
not \U$7638 ( \8015 , \8013 );
and \U$7639 ( \8016 , \8015 , \7205 );
nor \U$7640 ( \8017 , \8014 , \8016 );
nand \U$7641 ( \8018 , RIae7a3a8_177, RIae7a330_176);
and \U$7642 ( \8019 , \8018 , RIae7a240_174);
not \U$7643 ( \8020 , \8019 );
xor \U$7644 ( \8021 , \8017 , \8020 );
and \U$7645 ( \8022 , \6941 , RIae76b68_57);
and \U$7646 ( \8023 , RIae78a58_123, \6939 );
nor \U$7647 ( \8024 , \8022 , \8023 );
and \U$7648 ( \8025 , \8024 , \6314 );
not \U$7649 ( \8026 , \8024 );
and \U$7650 ( \8027 , \8026 , \6945 );
nor \U$7651 ( \8028 , \8025 , \8027 );
and \U$7652 ( \8029 , \8021 , \8028 );
and \U$7653 ( \8030 , \8017 , \8020 );
or \U$7654 ( \8031 , \8029 , \8030 );
xor \U$7655 ( \8032 , \8010 , \8031 );
and \U$7656 ( \8033 , \4688 , RIae76118_35);
and \U$7657 ( \8034 , RIae76028_33, \4686 );
nor \U$7658 ( \8035 , \8033 , \8034 );
and \U$7659 ( \8036 , \8035 , \4481 );
not \U$7660 ( \8037 , \8035 );
and \U$7661 ( \8038 , \8037 , \4482 );
nor \U$7662 ( \8039 , \8036 , \8038 );
and \U$7663 ( \8040 , \3730 , RIae763e8_41);
and \U$7664 ( \8041 , RIae764d8_43, \3728 );
nor \U$7665 ( \8042 , \8040 , \8041 );
and \U$7666 ( \8043 , \8042 , \3732 );
not \U$7667 ( \8044 , \8042 );
and \U$7668 ( \8045 , \8044 , \3422 );
nor \U$7669 ( \8046 , \8043 , \8045 );
xor \U$7670 ( \8047 , \8039 , \8046 );
and \U$7671 ( \8048 , \4247 , RIae766b8_47);
and \U$7672 ( \8049 , RIae765c8_45, \4245 );
nor \U$7673 ( \8050 , \8048 , \8049 );
and \U$7674 ( \8051 , \8050 , \3989 );
not \U$7675 ( \8052 , \8050 );
and \U$7676 ( \8053 , \8052 , \4251 );
nor \U$7677 ( \8054 , \8051 , \8053 );
and \U$7678 ( \8055 , \8047 , \8054 );
and \U$7679 ( \8056 , \8039 , \8046 );
or \U$7680 ( \8057 , \8055 , \8056 );
and \U$7681 ( \8058 , \8032 , \8057 );
and \U$7682 ( \8059 , \8010 , \8031 );
or \U$7683 ( \8060 , \8058 , \8059 );
xor \U$7684 ( \8061 , \7985 , \8060 );
and \U$7685 ( \8062 , \1593 , RIae75f38_31);
and \U$7686 ( \8063 , RIae75e48_29, \1591 );
nor \U$7687 ( \8064 , \8062 , \8063 );
and \U$7688 ( \8065 , \8064 , \1488 );
not \U$7689 ( \8066 , \8064 );
and \U$7690 ( \8067 , \8066 , \1498 );
nor \U$7691 ( \8068 , \8065 , \8067 );
not \U$7692 ( \8069 , \8068 );
and \U$7693 ( \8070 , \1939 , RIae75c68_25);
and \U$7694 ( \8071 , RIae75d58_27, \1937 );
nor \U$7695 ( \8072 , \8070 , \8071 );
and \U$7696 ( \8073 , \8072 , \1734 );
not \U$7697 ( \8074 , \8072 );
and \U$7698 ( \8075 , \8074 , \1735 );
nor \U$7699 ( \8076 , \8073 , \8075 );
not \U$7700 ( \8077 , \8076 );
and \U$7701 ( \8078 , \8069 , \8077 );
and \U$7702 ( \8079 , \8076 , \8068 );
and \U$7703 ( \8080 , \2224 , RIae755d8_11);
and \U$7704 ( \8081 , RIae754e8_9, \2222 );
nor \U$7705 ( \8082 , \8080 , \8081 );
and \U$7706 ( \8083 , \8082 , \2060 );
not \U$7707 ( \8084 , \8082 );
and \U$7708 ( \8085 , \8084 , \2061 );
nor \U$7709 ( \8086 , \8083 , \8085 );
nor \U$7710 ( \8087 , \8079 , \8086 );
nor \U$7711 ( \8088 , \8078 , \8087 );
and \U$7712 ( \8089 , \2607 , RIae757b8_15);
and \U$7713 ( \8090 , RIae756c8_13, \2605 );
nor \U$7714 ( \8091 , \8089 , \8090 );
and \U$7715 ( \8092 , \8091 , \2397 );
not \U$7716 ( \8093 , \8091 );
and \U$7717 ( \8094 , \8093 , \2611 );
nor \U$7718 ( \8095 , \8092 , \8094 );
not \U$7719 ( \8096 , \8095 );
and \U$7720 ( \8097 , \2783 , RIae75218_3);
and \U$7721 ( \8098 , RIae75128_1, \2781 );
nor \U$7722 ( \8099 , \8097 , \8098 );
not \U$7723 ( \8100 , \8099 );
not \U$7724 ( \8101 , \2789 );
and \U$7725 ( \8102 , \8100 , \8101 );
and \U$7726 ( \8103 , \8099 , \3089 );
nor \U$7727 ( \8104 , \8102 , \8103 );
not \U$7728 ( \8105 , \8104 );
and \U$7729 ( \8106 , \8096 , \8105 );
and \U$7730 ( \8107 , \8104 , \8095 );
and \U$7731 ( \8108 , \3214 , RIae75308_5);
and \U$7732 ( \8109 , RIae753f8_7, \3212 );
nor \U$7733 ( \8110 , \8108 , \8109 );
not \U$7734 ( \8111 , \8110 );
not \U$7735 ( \8112 , \3218 );
and \U$7736 ( \8113 , \8111 , \8112 );
and \U$7737 ( \8114 , \8110 , \3218 );
nor \U$7738 ( \8115 , \8113 , \8114 );
nor \U$7739 ( \8116 , \8107 , \8115 );
nor \U$7740 ( \8117 , \8106 , \8116 );
xor \U$7741 ( \8118 , \8088 , \8117 );
and \U$7742 ( \8119 , \883 , RIae78788_117);
and \U$7743 ( \8120 , RIae78698_115, \881 );
nor \U$7744 ( \8121 , \8119 , \8120 );
not \U$7745 ( \8122 , \8121 );
not \U$7746 ( \8123 , \789 );
and \U$7747 ( \8124 , \8122 , \8123 );
and \U$7748 ( \8125 , \8121 , \787 );
nor \U$7749 ( \8126 , \8124 , \8125 );
not \U$7750 ( \8127 , \8126 );
and \U$7751 ( \8128 , \1138 , RIae75b78_23);
and \U$7752 ( \8129 , RIae75a88_21, \1136 );
nor \U$7753 ( \8130 , \8128 , \8129 );
and \U$7754 ( \8131 , \8130 , \1142 );
not \U$7755 ( \8132 , \8130 );
and \U$7756 ( \8133 , \8132 , \1012 );
nor \U$7757 ( \8134 , \8131 , \8133 );
not \U$7758 ( \8135 , \8134 );
and \U$7759 ( \8136 , \8127 , \8135 );
and \U$7760 ( \8137 , \8134 , \8126 );
and \U$7761 ( \8138 , \1376 , RIae75998_19);
and \U$7762 ( \8139 , RIae758a8_17, \1374 );
nor \U$7763 ( \8140 , \8138 , \8139 );
and \U$7764 ( \8141 , \8140 , \1261 );
not \U$7765 ( \8142 , \8140 );
and \U$7766 ( \8143 , \8142 , \1380 );
nor \U$7767 ( \8144 , \8141 , \8143 );
nor \U$7768 ( \8145 , \8137 , \8144 );
nor \U$7769 ( \8146 , \8136 , \8145 );
and \U$7770 ( \8147 , \8118 , \8146 );
and \U$7771 ( \8148 , \8088 , \8117 );
nor \U$7772 ( \8149 , \8147 , \8148 );
and \U$7773 ( \8150 , \8061 , \8149 );
and \U$7774 ( \8151 , \7985 , \8060 );
or \U$7775 ( \8152 , \8150 , \8151 );
xor \U$7776 ( \8153 , \7930 , \8152 );
xor \U$7777 ( \8154 , \7203 , \7206 );
xor \U$7778 ( \8155 , \8154 , \7214 );
xor \U$7779 ( \8156 , \7576 , \7578 );
xor \U$7780 ( \8157 , \8156 , \7581 );
and \U$7781 ( \8158 , \8155 , \8157 );
xor \U$7782 ( \8159 , \7097 , \7104 );
xor \U$7783 ( \8160 , \8159 , \7112 );
xor \U$7784 ( \8161 , \7564 , \7569 );
xor \U$7785 ( \8162 , \8160 , \8161 );
xor \U$7786 ( \8163 , \7576 , \7578 );
xor \U$7787 ( \8164 , \8163 , \7581 );
and \U$7788 ( \8165 , \8162 , \8164 );
and \U$7789 ( \8166 , \8155 , \8162 );
or \U$7790 ( \8167 , \8158 , \8165 , \8166 );
and \U$7791 ( \8168 , \8153 , \8167 );
and \U$7792 ( \8169 , \7930 , \8152 );
or \U$7793 ( \8170 , \8168 , \8169 );
xor \U$7794 ( \8171 , \7010 , \7012 );
xor \U$7795 ( \8172 , \8171 , \7087 );
xor \U$7796 ( \8173 , \8170 , \8172 );
xor \U$7797 ( \8174 , \7754 , \7779 );
xor \U$7798 ( \8175 , \8174 , \7806 );
xor \U$7799 ( \8176 , \7688 , \7696 );
xor \U$7800 ( \8177 , \8176 , \7724 );
xor \U$7801 ( \8178 , \8175 , \8177 );
xor \U$7802 ( \8179 , \7618 , \7649 );
xor \U$7803 ( \8180 , \8179 , \7675 );
and \U$7804 ( \8181 , \8178 , \8180 );
and \U$7805 ( \8182 , \8175 , \8177 );
or \U$7806 ( \8183 , \8181 , \8182 );
xor \U$7807 ( \8184 , \7196 , \7217 );
xor \U$7808 ( \8185 , \8184 , \7244 );
xor \U$7809 ( \8186 , \8183 , \8185 );
xor \U$7810 ( \8187 , \7037 , \7060 );
xor \U$7811 ( \8188 , \8187 , \7084 );
xor \U$7812 ( \8189 , \7815 , \7820 );
xor \U$7813 ( \8190 , \8188 , \8189 );
and \U$7814 ( \8191 , \8186 , \8190 );
and \U$7815 ( \8192 , \8183 , \8185 );
or \U$7816 ( \8193 , \8191 , \8192 );
and \U$7817 ( \8194 , \8173 , \8193 );
and \U$7818 ( \8195 , \8170 , \8172 );
or \U$7819 ( \8196 , \8194 , \8195 );
and \U$7820 ( \8197 , \7902 , \8196 );
and \U$7821 ( \8198 , \7899 , \7901 );
or \U$7822 ( \8199 , \8197 , \8198 );
nand \U$7823 ( \8200 , \7885 , \8199 );
nand \U$7824 ( \8201 , \7882 , \8200 );
not \U$7825 ( \8202 , \8201 );
not \U$7826 ( \8203 , \7845 );
not \U$7827 ( \8204 , \7532 );
and \U$7828 ( \8205 , \8203 , \8204 );
and \U$7829 ( \8206 , \7845 , \7532 );
nor \U$7830 ( \8207 , \8205 , \8206 );
not \U$7831 ( \8208 , \8207 );
not \U$7832 ( \8209 , \7529 );
and \U$7833 ( \8210 , \8208 , \8209 );
and \U$7834 ( \8211 , \8207 , \7529 );
nor \U$7835 ( \8212 , \8210 , \8211 );
nor \U$7836 ( \8213 , \8202 , \8212 );
and \U$7837 ( \8214 , \7869 , \8213 );
xor \U$7838 ( \8215 , \8213 , \7869 );
not \U$7839 ( \8216 , \8212 );
not \U$7840 ( \8217 , \8201 );
and \U$7841 ( \8218 , \8216 , \8217 );
and \U$7842 ( \8219 , \8212 , \8201 );
nor \U$7843 ( \8220 , \8218 , \8219 );
not \U$7844 ( \8221 , \7881 );
not \U$7845 ( \8222 , \8199 );
or \U$7846 ( \8223 , \8221 , \8222 );
or \U$7847 ( \8224 , \8199 , \7881 );
nand \U$7848 ( \8225 , \8223 , \8224 );
not \U$7849 ( \8226 , \8225 );
not \U$7850 ( \8227 , \7871 );
and \U$7851 ( \8228 , \8226 , \8227 );
and \U$7852 ( \8229 , \8225 , \7871 );
nor \U$7853 ( \8230 , \8228 , \8229 );
not \U$7854 ( \8231 , \8230 );
not \U$7855 ( \8232 , \8095 );
xor \U$7856 ( \8233 , \8104 , \8115 );
not \U$7857 ( \8234 , \8233 );
or \U$7858 ( \8235 , \8232 , \8234 );
or \U$7859 ( \8236 , \8233 , \8095 );
nand \U$7860 ( \8237 , \8235 , \8236 );
xor \U$7861 ( \8238 , \8039 , \8046 );
xor \U$7862 ( \8239 , \8238 , \8054 );
xor \U$7863 ( \8240 , \8237 , \8239 );
xor \U$7864 ( \8241 , \7992 , \7999 );
xor \U$7865 ( \8242 , \8241 , \8007 );
and \U$7866 ( \8243 , \8240 , \8242 );
and \U$7867 ( \8244 , \8237 , \8239 );
or \U$7868 ( \8245 , \8243 , \8244 );
xor \U$7869 ( \8246 , \7625 , \7638 );
xor \U$7870 ( \8247 , \8246 , \7646 );
xor \U$7871 ( \8248 , \8245 , \8247 );
not \U$7872 ( \8249 , \8126 );
xor \U$7873 ( \8250 , \8134 , \8144 );
not \U$7874 ( \8251 , \8250 );
or \U$7875 ( \8252 , \8249 , \8251 );
or \U$7876 ( \8253 , \8250 , \8126 );
nand \U$7877 ( \8254 , \8252 , \8253 );
xor \U$7878 ( \8255 , \7963 , \7971 );
xor \U$7879 ( \8256 , \8255 , \7979 );
and \U$7880 ( \8257 , \8254 , \8256 );
not \U$7881 ( \8258 , \8068 );
xor \U$7882 ( \8259 , \8076 , \8086 );
not \U$7883 ( \8260 , \8259 );
or \U$7884 ( \8261 , \8258 , \8260 );
or \U$7885 ( \8262 , \8259 , \8068 );
nand \U$7886 ( \8263 , \8261 , \8262 );
xor \U$7887 ( \8264 , \7963 , \7971 );
xor \U$7888 ( \8265 , \8264 , \7979 );
and \U$7889 ( \8266 , \8263 , \8265 );
and \U$7890 ( \8267 , \8254 , \8263 );
or \U$7891 ( \8268 , \8257 , \8266 , \8267 );
and \U$7892 ( \8269 , \8248 , \8268 );
and \U$7893 ( \8270 , \8245 , \8247 );
or \U$7894 ( \8271 , \8269 , \8270 );
and \U$7895 ( \8272 , \883 , RIae78878_119);
and \U$7896 ( \8273 , RIae78788_117, \881 );
nor \U$7897 ( \8274 , \8272 , \8273 );
not \U$7898 ( \8275 , \8274 );
not \U$7899 ( \8276 , \787 );
and \U$7900 ( \8277 , \8275 , \8276 );
and \U$7901 ( \8278 , \8274 , \789 );
nor \U$7902 ( \8279 , \8277 , \8278 );
and \U$7903 ( \8280 , \1138 , RIae78698_115);
and \U$7904 ( \8281 , RIae75b78_23, \1136 );
nor \U$7905 ( \8282 , \8280 , \8281 );
and \U$7906 ( \8283 , \8282 , \1142 );
not \U$7907 ( \8284 , \8282 );
and \U$7908 ( \8285 , \8284 , \1012 );
nor \U$7909 ( \8286 , \8283 , \8285 );
xor \U$7910 ( \8287 , \8279 , \8286 );
and \U$7911 ( \8288 , \1376 , RIae75a88_21);
and \U$7912 ( \8289 , RIae75998_19, \1374 );
nor \U$7913 ( \8290 , \8288 , \8289 );
and \U$7914 ( \8291 , \8290 , \1261 );
not \U$7915 ( \8292 , \8290 );
and \U$7916 ( \8293 , \8292 , \1380 );
nor \U$7917 ( \8294 , \8291 , \8293 );
and \U$7918 ( \8295 , \8287 , \8294 );
and \U$7919 ( \8296 , \8279 , \8286 );
or \U$7920 ( \8297 , \8295 , \8296 );
and \U$7921 ( \8298 , \2607 , RIae754e8_9);
and \U$7922 ( \8299 , RIae757b8_15, \2605 );
nor \U$7923 ( \8300 , \8298 , \8299 );
and \U$7924 ( \8301 , \8300 , \2397 );
not \U$7925 ( \8302 , \8300 );
and \U$7926 ( \8303 , \8302 , \2611 );
nor \U$7927 ( \8304 , \8301 , \8303 );
not \U$7928 ( \8305 , \8304 );
and \U$7929 ( \8306 , \2783 , RIae756c8_13);
and \U$7930 ( \8307 , RIae75218_3, \2781 );
nor \U$7931 ( \8308 , \8306 , \8307 );
not \U$7932 ( \8309 , \8308 );
not \U$7933 ( \8310 , \3089 );
and \U$7934 ( \8311 , \8309 , \8310 );
and \U$7935 ( \8312 , \8308 , \3089 );
nor \U$7936 ( \8313 , \8311 , \8312 );
not \U$7937 ( \8314 , \8313 );
and \U$7938 ( \8315 , \8305 , \8314 );
and \U$7939 ( \8316 , \8313 , \8304 );
and \U$7940 ( \8317 , \3214 , RIae75128_1);
and \U$7941 ( \8318 , RIae75308_5, \3212 );
nor \U$7942 ( \8319 , \8317 , \8318 );
not \U$7943 ( \8320 , \8319 );
not \U$7944 ( \8321 , \2774 );
and \U$7945 ( \8322 , \8320 , \8321 );
and \U$7946 ( \8323 , \8319 , \2774 );
nor \U$7947 ( \8324 , \8322 , \8323 );
nor \U$7948 ( \8325 , \8316 , \8324 );
nor \U$7949 ( \8326 , \8315 , \8325 );
or \U$7950 ( \8327 , \8297 , \8326 );
not \U$7951 ( \8328 , \8297 );
not \U$7952 ( \8329 , \8326 );
or \U$7953 ( \8330 , \8328 , \8329 );
and \U$7954 ( \8331 , \2224 , RIae75d58_27);
and \U$7955 ( \8332 , RIae755d8_11, \2222 );
nor \U$7956 ( \8333 , \8331 , \8332 );
and \U$7957 ( \8334 , \8333 , \2061 );
not \U$7958 ( \8335 , \8333 );
and \U$7959 ( \8336 , \8335 , \2060 );
nor \U$7960 ( \8337 , \8334 , \8336 );
and \U$7961 ( \8338 , \1593 , RIae758a8_17);
and \U$7962 ( \8339 , RIae75f38_31, \1591 );
nor \U$7963 ( \8340 , \8338 , \8339 );
and \U$7964 ( \8341 , \8340 , \1498 );
not \U$7965 ( \8342 , \8340 );
and \U$7966 ( \8343 , \8342 , \1488 );
nor \U$7967 ( \8344 , \8341 , \8343 );
xor \U$7968 ( \8345 , \8337 , \8344 );
and \U$7969 ( \8346 , \1939 , RIae75e48_29);
and \U$7970 ( \8347 , RIae75c68_25, \1937 );
nor \U$7971 ( \8348 , \8346 , \8347 );
and \U$7972 ( \8349 , \8348 , \1735 );
not \U$7973 ( \8350 , \8348 );
and \U$7974 ( \8351 , \8350 , \1734 );
nor \U$7975 ( \8352 , \8349 , \8351 );
and \U$7976 ( \8353 , \8345 , \8352 );
and \U$7977 ( \8354 , \8337 , \8344 );
or \U$7978 ( \8355 , \8353 , \8354 );
nand \U$7979 ( \8356 , \8330 , \8355 );
nand \U$7980 ( \8357 , \8327 , \8356 );
and \U$7981 ( \8358 , \6941 , RIae76898_51);
and \U$7982 ( \8359 , RIae76b68_57, \6939 );
nor \U$7983 ( \8360 , \8358 , \8359 );
and \U$7984 ( \8361 , \8360 , \6945 );
not \U$7985 ( \8362 , \8360 );
and \U$7986 ( \8363 , \8362 , \6314 );
nor \U$7987 ( \8364 , \8361 , \8363 );
and \U$7988 ( \8365 , RIae7a240_174, RIae7a330_176);
not \U$7989 ( \8366 , RIae7a3a8_177);
and \U$7990 ( \8367 , \8366 , RIae7a330_176);
nor \U$7991 ( \8368 , \8366 , RIae7a330_176);
or \U$7992 ( \8369 , \8367 , \8368 );
nor \U$7993 ( \8370 , RIae7a240_174, RIae7a330_176);
nor \U$7994 ( \8371 , \8365 , \8369 , \8370 );
nand \U$7995 ( \8372 , RIae78da0_130, \8371 );
and \U$7996 ( \8373 , \8372 , \8019 );
not \U$7997 ( \8374 , \8372 );
and \U$7998 ( \8375 , \8374 , \8020 );
nor \U$7999 ( \8376 , \8373 , \8375 );
xor \U$8000 ( \8377 , \8364 , \8376 );
and \U$8001 ( \8378 , \7633 , RIae78a58_123);
and \U$8002 ( \8379 , RIae78cb0_128, \7631 );
nor \U$8003 ( \8380 , \8378 , \8379 );
and \U$8004 ( \8381 , \8380 , \7205 );
not \U$8005 ( \8382 , \8380 );
and \U$8006 ( \8383 , \8382 , \7206 );
nor \U$8007 ( \8384 , \8381 , \8383 );
and \U$8008 ( \8385 , \8377 , \8384 );
and \U$8009 ( \8386 , \8364 , \8376 );
or \U$8010 ( \8387 , \8385 , \8386 );
and \U$8011 ( \8388 , \4247 , RIae764d8_43);
and \U$8012 ( \8389 , RIae766b8_47, \4245 );
nor \U$8013 ( \8390 , \8388 , \8389 );
and \U$8014 ( \8391 , \8390 , \3989 );
not \U$8015 ( \8392 , \8390 );
and \U$8016 ( \8393 , \8392 , \4251 );
nor \U$8017 ( \8394 , \8391 , \8393 );
and \U$8018 ( \8395 , \4688 , RIae765c8_45);
and \U$8019 ( \8396 , RIae76118_35, \4686 );
nor \U$8020 ( \8397 , \8395 , \8396 );
and \U$8021 ( \8398 , \8397 , \4481 );
not \U$8022 ( \8399 , \8397 );
and \U$8023 ( \8400 , \8399 , \4482 );
nor \U$8024 ( \8401 , \8398 , \8400 );
xor \U$8025 ( \8402 , \8394 , \8401 );
and \U$8026 ( \8403 , \3730 , RIae753f8_7);
and \U$8027 ( \8404 , RIae763e8_41, \3728 );
nor \U$8028 ( \8405 , \8403 , \8404 );
and \U$8029 ( \8406 , \8405 , \3732 );
not \U$8030 ( \8407 , \8405 );
and \U$8031 ( \8408 , \8407 , \3422 );
nor \U$8032 ( \8409 , \8406 , \8408 );
and \U$8033 ( \8410 , \8402 , \8409 );
and \U$8034 ( \8411 , \8394 , \8401 );
nor \U$8035 ( \8412 , \8410 , \8411 );
or \U$8036 ( \8413 , \8387 , \8412 );
not \U$8037 ( \8414 , \8387 );
not \U$8038 ( \8415 , \8412 );
or \U$8039 ( \8416 , \8414 , \8415 );
and \U$8040 ( \8417 , \5399 , RIae76028_33);
and \U$8041 ( \8418 , RIae762f8_39, \5397 );
nor \U$8042 ( \8419 , \8417 , \8418 );
and \U$8043 ( \8420 , \8419 , \5016 );
not \U$8044 ( \8421 , \8419 );
and \U$8045 ( \8422 , \8421 , \5403 );
nor \U$8046 ( \8423 , \8420 , \8422 );
and \U$8047 ( \8424 , \5896 , RIae76208_37);
and \U$8048 ( \8425 , RIae76a78_55, \5894 );
nor \U$8049 ( \8426 , \8424 , \8425 );
and \U$8050 ( \8427 , \8426 , \5590 );
not \U$8051 ( \8428 , \8426 );
and \U$8052 ( \8429 , \8428 , \5589 );
nor \U$8053 ( \8430 , \8427 , \8429 );
xor \U$8054 ( \8431 , \8423 , \8430 );
and \U$8055 ( \8432 , \6172 , RIae76988_53);
and \U$8056 ( \8433 , RIae767a8_49, \6170 );
nor \U$8057 ( \8434 , \8432 , \8433 );
and \U$8058 ( \8435 , \8434 , \6176 );
not \U$8059 ( \8436 , \8434 );
and \U$8060 ( \8437 , \8436 , \6175 );
nor \U$8061 ( \8438 , \8435 , \8437 );
and \U$8062 ( \8439 , \8431 , \8438 );
and \U$8063 ( \8440 , \8423 , \8430 );
or \U$8064 ( \8441 , \8439 , \8440 );
nand \U$8065 ( \8442 , \8416 , \8441 );
nand \U$8066 ( \8443 , \8413 , \8442 );
xor \U$8067 ( \8444 , \8357 , \8443 );
not \U$8068 ( \8445 , \7938 );
not \U$8069 ( \8446 , \7951 );
or \U$8070 ( \8447 , \8445 , \8446 );
or \U$8071 ( \8448 , \7938 , \7951 );
nand \U$8072 ( \8449 , \8447 , \8448 );
not \U$8073 ( \8450 , \8449 );
not \U$8074 ( \8451 , \7939 );
and \U$8075 ( \8452 , \8450 , \8451 );
and \U$8076 ( \8453 , \8449 , \7939 );
nor \U$8077 ( \8454 , \8452 , \8453 );
and \U$8078 ( \8455 , \436 , RIae785a8_113);
and \U$8079 ( \8456 , RIae783c8_109, \434 );
nor \U$8080 ( \8457 , \8455 , \8456 );
not \U$8081 ( \8458 , \8457 );
not \U$8082 ( \8459 , \402 );
and \U$8083 ( \8460 , \8458 , \8459 );
and \U$8084 ( \8461 , \8457 , \402 );
nor \U$8085 ( \8462 , \8460 , \8461 );
nand \U$8086 ( \8463 , RIae77f18_99, RIae78b48_125);
xor \U$8087 ( \8464 , \8462 , \8463 );
and \U$8088 ( \8465 , \384 , RIae78008_101);
and \U$8089 ( \8466 , RIae781e8_105, \382 );
nor \U$8090 ( \8467 , \8465 , \8466 );
not \U$8091 ( \8468 , \8467 );
not \U$8092 ( \8469 , \392 );
and \U$8093 ( \8470 , \8468 , \8469 );
and \U$8094 ( \8471 , \8467 , \388 );
nor \U$8095 ( \8472 , \8470 , \8471 );
and \U$8096 ( \8473 , \8464 , \8472 );
and \U$8097 ( \8474 , \8462 , \8463 );
or \U$8098 ( \8475 , \8473 , \8474 );
or \U$8099 ( \8476 , \8454 , \8475 );
not \U$8100 ( \8477 , \8475 );
not \U$8101 ( \8478 , \8454 );
or \U$8102 ( \8479 , \8477 , \8478 );
and \U$8103 ( \8480 , \558 , RIae77b58_91);
and \U$8104 ( \8481 , RIae77d38_95, \556 );
nor \U$8105 ( \8482 , \8480 , \8481 );
and \U$8106 ( \8483 , \8482 , \562 );
not \U$8107 ( \8484 , \8482 );
and \U$8108 ( \8485 , \8484 , \504 );
nor \U$8109 ( \8486 , \8483 , \8485 );
and \U$8110 ( \8487 , \672 , RIae77e28_97);
and \U$8111 ( \8488 , RIae78968_121, \670 );
nor \U$8112 ( \8489 , \8487 , \8488 );
and \U$8113 ( \8490 , \8489 , \587 );
not \U$8114 ( \8491 , \8489 );
and \U$8115 ( \8492 , \8491 , \588 );
nor \U$8116 ( \8493 , \8490 , \8492 );
xor \U$8117 ( \8494 , \8486 , \8493 );
and \U$8118 ( \8495 , \514 , RIae78530_112);
and \U$8119 ( \8496 , RIae77c48_93, \512 );
nor \U$8120 ( \8497 , \8495 , \8496 );
not \U$8121 ( \8498 , \8497 );
not \U$8122 ( \8499 , \469 );
and \U$8123 ( \8500 , \8498 , \8499 );
and \U$8124 ( \8501 , \8497 , \469 );
nor \U$8125 ( \8502 , \8500 , \8501 );
and \U$8126 ( \8503 , \8494 , \8502 );
and \U$8127 ( \8504 , \8486 , \8493 );
nor \U$8128 ( \8505 , \8503 , \8504 );
nand \U$8129 ( \8506 , \8479 , \8505 );
nand \U$8130 ( \8507 , \8476 , \8506 );
and \U$8131 ( \8508 , \8444 , \8507 );
and \U$8132 ( \8509 , \8357 , \8443 );
or \U$8133 ( \8510 , \8508 , \8509 );
xor \U$8134 ( \8511 , \8271 , \8510 );
xor \U$8135 ( \8512 , \7953 , \7955 );
xor \U$8136 ( \8513 , \8512 , \7982 );
xor \U$8137 ( \8514 , \7919 , \7921 );
xor \U$8138 ( \8515 , \8514 , \7924 );
and \U$8139 ( \8516 , \8513 , \8515 );
xor \U$8140 ( \8517 , \7657 , \7664 );
xor \U$8141 ( \8518 , \8517 , \7672 );
xor \U$8142 ( \8519 , \7904 , \7909 );
xor \U$8143 ( \8520 , \8518 , \8519 );
xor \U$8144 ( \8521 , \7919 , \7921 );
xor \U$8145 ( \8522 , \8521 , \7924 );
and \U$8146 ( \8523 , \8520 , \8522 );
and \U$8147 ( \8524 , \8513 , \8520 );
or \U$8148 ( \8525 , \8516 , \8523 , \8524 );
and \U$8149 ( \8526 , \8511 , \8525 );
and \U$8150 ( \8527 , \8271 , \8510 );
or \U$8151 ( \8528 , \8526 , \8527 );
xor \U$8152 ( \8529 , \7574 , \7584 );
xor \U$8153 ( \8530 , \8529 , \7589 );
xor \U$8154 ( \8531 , \8528 , \8530 );
xor \U$8155 ( \8532 , \7914 , \7916 );
xor \U$8156 ( \8533 , \8532 , \7927 );
xor \U$8157 ( \8534 , \8175 , \8177 );
xor \U$8158 ( \8535 , \8534 , \8180 );
and \U$8159 ( \8536 , \8533 , \8535 );
xor \U$8160 ( \8537 , \7576 , \7578 );
xor \U$8161 ( \8538 , \8537 , \7581 );
xor \U$8162 ( \8539 , \8155 , \8162 );
xor \U$8163 ( \8540 , \8538 , \8539 );
xor \U$8164 ( \8541 , \8175 , \8177 );
xor \U$8165 ( \8542 , \8541 , \8180 );
and \U$8166 ( \8543 , \8540 , \8542 );
and \U$8167 ( \8544 , \8533 , \8540 );
or \U$8168 ( \8545 , \8536 , \8543 , \8544 );
and \U$8169 ( \8546 , \8531 , \8545 );
and \U$8170 ( \8547 , \8528 , \8530 );
or \U$8171 ( \8548 , \8546 , \8547 );
xor \U$8172 ( \8549 , \7678 , \7727 );
xor \U$8173 ( \8550 , \8549 , \7809 );
xor \U$8174 ( \8551 , \8183 , \8185 );
xor \U$8175 ( \8552 , \8551 , \8190 );
and \U$8176 ( \8553 , \8550 , \8552 );
xor \U$8177 ( \8554 , \7930 , \8152 );
xor \U$8178 ( \8555 , \8554 , \8167 );
xor \U$8179 ( \8556 , \8183 , \8185 );
xor \U$8180 ( \8557 , \8556 , \8190 );
and \U$8181 ( \8558 , \8555 , \8557 );
and \U$8182 ( \8559 , \8550 , \8555 );
or \U$8183 ( \8560 , \8553 , \8558 , \8559 );
xor \U$8184 ( \8561 , \8548 , \8560 );
xor \U$8185 ( \8562 , \7891 , \7893 );
xor \U$8186 ( \8563 , \8562 , \7896 );
and \U$8187 ( \8564 , \8561 , \8563 );
and \U$8188 ( \8565 , \8548 , \8560 );
or \U$8189 ( \8566 , \8564 , \8565 );
not \U$8190 ( \8567 , \7880 );
not \U$8191 ( \8568 , \7873 );
or \U$8192 ( \8569 , \8567 , \8568 );
or \U$8193 ( \8570 , \7873 , \7880 );
nand \U$8194 ( \8571 , \8569 , \8570 );
xor \U$8195 ( \8572 , \8566 , \8571 );
xor \U$8196 ( \8573 , \7899 , \7901 );
xor \U$8197 ( \8574 , \8573 , \8196 );
and \U$8198 ( \8575 , \8572 , \8574 );
and \U$8199 ( \8576 , \8566 , \8571 );
or \U$8200 ( \8577 , \8575 , \8576 );
nand \U$8201 ( \8578 , \8231 , \8577 );
or \U$8202 ( \8579 , \8220 , \8578 );
xnor \U$8203 ( \8580 , \8578 , \8220 );
and \U$8204 ( \8581 , \2607 , RIae755d8_11);
and \U$8205 ( \8582 , RIae754e8_9, \2605 );
nor \U$8206 ( \8583 , \8581 , \8582 );
and \U$8207 ( \8584 , \8583 , \2611 );
not \U$8208 ( \8585 , \8583 );
and \U$8209 ( \8586 , \8585 , \2397 );
nor \U$8210 ( \8587 , \8584 , \8586 );
and \U$8211 ( \8588 , \1939 , RIae75f38_31);
and \U$8212 ( \8589 , RIae75e48_29, \1937 );
nor \U$8213 ( \8590 , \8588 , \8589 );
and \U$8214 ( \8591 , \8590 , \1735 );
not \U$8215 ( \8592 , \8590 );
and \U$8216 ( \8593 , \8592 , \1734 );
nor \U$8217 ( \8594 , \8591 , \8593 );
xor \U$8218 ( \8595 , \8587 , \8594 );
and \U$8219 ( \8596 , \2224 , RIae75c68_25);
and \U$8220 ( \8597 , RIae75d58_27, \2222 );
nor \U$8221 ( \8598 , \8596 , \8597 );
and \U$8222 ( \8599 , \8598 , \2061 );
not \U$8223 ( \8600 , \8598 );
and \U$8224 ( \8601 , \8600 , \2060 );
nor \U$8225 ( \8602 , \8599 , \8601 );
and \U$8226 ( \8603 , \8595 , \8602 );
and \U$8227 ( \8604 , \8587 , \8594 );
or \U$8228 ( \8605 , \8603 , \8604 );
and \U$8229 ( \8606 , \1593 , RIae75998_19);
and \U$8230 ( \8607 , RIae758a8_17, \1591 );
nor \U$8231 ( \8608 , \8606 , \8607 );
and \U$8232 ( \8609 , \8608 , \1498 );
not \U$8233 ( \8610 , \8608 );
and \U$8234 ( \8611 , \8610 , \1488 );
nor \U$8235 ( \8612 , \8609 , \8611 );
and \U$8236 ( \8613 , \1138 , RIae78788_117);
and \U$8237 ( \8614 , RIae78698_115, \1136 );
nor \U$8238 ( \8615 , \8613 , \8614 );
and \U$8239 ( \8616 , \8615 , \1012 );
not \U$8240 ( \8617 , \8615 );
and \U$8241 ( \8618 , \8617 , \1142 );
nor \U$8242 ( \8619 , \8616 , \8618 );
xor \U$8243 ( \8620 , \8612 , \8619 );
and \U$8244 ( \8621 , \1376 , RIae75b78_23);
and \U$8245 ( \8622 , RIae75a88_21, \1374 );
nor \U$8246 ( \8623 , \8621 , \8622 );
and \U$8247 ( \8624 , \8623 , \1380 );
not \U$8248 ( \8625 , \8623 );
and \U$8249 ( \8626 , \8625 , \1261 );
nor \U$8250 ( \8627 , \8624 , \8626 );
and \U$8251 ( \8628 , \8620 , \8627 );
and \U$8252 ( \8629 , \8612 , \8619 );
or \U$8253 ( \8630 , \8628 , \8629 );
xor \U$8254 ( \8631 , \8605 , \8630 );
not \U$8255 ( \8632 , \3218 );
and \U$8256 ( \8633 , \3214 , RIae75218_3);
and \U$8257 ( \8634 , RIae75128_1, \3212 );
nor \U$8258 ( \8635 , \8633 , \8634 );
not \U$8259 ( \8636 , \8635 );
or \U$8260 ( \8637 , \8632 , \8636 );
or \U$8261 ( \8638 , \8635 , \2774 );
nand \U$8262 ( \8639 , \8637 , \8638 );
not \U$8263 ( \8640 , \2789 );
and \U$8264 ( \8641 , \2783 , RIae757b8_15);
and \U$8265 ( \8642 , RIae756c8_13, \2781 );
nor \U$8266 ( \8643 , \8641 , \8642 );
not \U$8267 ( \8644 , \8643 );
or \U$8268 ( \8645 , \8640 , \8644 );
or \U$8269 ( \8646 , \8643 , \2789 );
nand \U$8270 ( \8647 , \8645 , \8646 );
xor \U$8271 ( \8648 , \8639 , \8647 );
and \U$8272 ( \8649 , \3730 , RIae75308_5);
and \U$8273 ( \8650 , RIae753f8_7, \3728 );
nor \U$8274 ( \8651 , \8649 , \8650 );
and \U$8275 ( \8652 , \8651 , \3732 );
not \U$8276 ( \8653 , \8651 );
and \U$8277 ( \8654 , \8653 , \3422 );
nor \U$8278 ( \8655 , \8652 , \8654 );
and \U$8279 ( \8656 , \8648 , \8655 );
and \U$8280 ( \8657 , \8639 , \8647 );
or \U$8281 ( \8658 , \8656 , \8657 );
and \U$8282 ( \8659 , \8631 , \8658 );
and \U$8283 ( \8660 , \8605 , \8630 );
nor \U$8284 ( \8661 , \8659 , \8660 );
not \U$8285 ( \8662 , \8661 );
and \U$8286 ( \8663 , \672 , RIae77d38_95);
and \U$8287 ( \8664 , RIae77e28_97, \670 );
nor \U$8288 ( \8665 , \8663 , \8664 );
and \U$8289 ( \8666 , \8665 , \588 );
not \U$8290 ( \8667 , \8665 );
and \U$8291 ( \8668 , \8667 , \587 );
nor \U$8292 ( \8669 , \8666 , \8668 );
not \U$8293 ( \8670 , \787 );
and \U$8294 ( \8671 , \883 , RIae78968_121);
and \U$8295 ( \8672 , RIae78878_119, \881 );
nor \U$8296 ( \8673 , \8671 , \8672 );
not \U$8297 ( \8674 , \8673 );
or \U$8298 ( \8675 , \8670 , \8674 );
or \U$8299 ( \8676 , \8673 , \789 );
nand \U$8300 ( \8677 , \8675 , \8676 );
xor \U$8301 ( \8678 , \8669 , \8677 );
and \U$8302 ( \8679 , \558 , RIae77c48_93);
and \U$8303 ( \8680 , RIae77b58_91, \556 );
nor \U$8304 ( \8681 , \8679 , \8680 );
and \U$8305 ( \8682 , \8681 , \504 );
not \U$8306 ( \8683 , \8681 );
and \U$8307 ( \8684 , \8683 , \562 );
nor \U$8308 ( \8685 , \8682 , \8684 );
and \U$8309 ( \8686 , \8678 , \8685 );
and \U$8310 ( \8687 , \8669 , \8677 );
nor \U$8311 ( \8688 , \8686 , \8687 );
and \U$8312 ( \8689 , \384 , RIae77f18_99);
and \U$8313 ( \8690 , RIae78008_101, \382 );
nor \U$8314 ( \8691 , \8689 , \8690 );
not \U$8315 ( \8692 , \8691 );
not \U$8316 ( \8693 , \392 );
and \U$8317 ( \8694 , \8692 , \8693 );
and \U$8318 ( \8695 , \8691 , \392 );
nor \U$8319 ( \8696 , \8694 , \8695 );
not \U$8320 ( \8697 , \8696 );
and \U$8321 ( \8698 , \436 , RIae781e8_105);
and \U$8322 ( \8699 , RIae785a8_113, \434 );
nor \U$8323 ( \8700 , \8698 , \8699 );
not \U$8324 ( \8701 , \8700 );
not \U$8325 ( \8702 , \400 );
and \U$8326 ( \8703 , \8701 , \8702 );
and \U$8327 ( \8704 , \8700 , \402 );
nor \U$8328 ( \8705 , \8703 , \8704 );
not \U$8329 ( \8706 , \8705 );
and \U$8330 ( \8707 , \8697 , \8706 );
and \U$8331 ( \8708 , \8705 , \8696 );
and \U$8332 ( \8709 , \514 , RIae783c8_109);
and \U$8333 ( \8710 , RIae78530_112, \512 );
nor \U$8334 ( \8711 , \8709 , \8710 );
not \U$8335 ( \8712 , \8711 );
not \U$8336 ( \8713 , \469 );
and \U$8337 ( \8714 , \8712 , \8713 );
and \U$8338 ( \8715 , \8711 , \471 );
nor \U$8339 ( \8716 , \8714 , \8715 );
nor \U$8340 ( \8717 , \8708 , \8716 );
nor \U$8341 ( \8718 , \8707 , \8717 );
nand \U$8342 ( \8719 , \8688 , \8718 );
not \U$8343 ( \8720 , \8719 );
not \U$8344 ( \8721 , \8720 );
and \U$8345 ( \8722 , \8662 , \8721 );
and \U$8346 ( \8723 , \8661 , \8720 );
and \U$8347 ( \8724 , \4688 , RIae766b8_47);
and \U$8348 ( \8725 , RIae765c8_45, \4686 );
nor \U$8349 ( \8726 , \8724 , \8725 );
and \U$8350 ( \8727 , \8726 , \4481 );
not \U$8351 ( \8728 , \8726 );
and \U$8352 ( \8729 , \8728 , \4482 );
nor \U$8353 ( \8730 , \8727 , \8729 );
and \U$8354 ( \8731 , \5399 , RIae76118_35);
and \U$8355 ( \8732 , RIae76028_33, \5397 );
nor \U$8356 ( \8733 , \8731 , \8732 );
and \U$8357 ( \8734 , \8733 , \5016 );
not \U$8358 ( \8735 , \8733 );
and \U$8359 ( \8736 , \8735 , \5403 );
nor \U$8360 ( \8737 , \8734 , \8736 );
xor \U$8361 ( \8738 , \8730 , \8737 );
and \U$8362 ( \8739 , \4247 , RIae763e8_41);
and \U$8363 ( \8740 , RIae764d8_43, \4245 );
nor \U$8364 ( \8741 , \8739 , \8740 );
and \U$8365 ( \8742 , \8741 , \3989 );
not \U$8366 ( \8743 , \8741 );
and \U$8367 ( \8744 , \8743 , \4251 );
nor \U$8368 ( \8745 , \8742 , \8744 );
and \U$8369 ( \8746 , \8738 , \8745 );
and \U$8370 ( \8747 , \8730 , \8737 );
nor \U$8371 ( \8748 , \8746 , \8747 );
not \U$8372 ( \8749 , \8748 );
and \U$8373 ( \8750 , \5896 , RIae762f8_39);
and \U$8374 ( \8751 , RIae76208_37, \5894 );
nor \U$8375 ( \8752 , \8750 , \8751 );
and \U$8376 ( \8753 , \8752 , \5589 );
not \U$8377 ( \8754 , \8752 );
and \U$8378 ( \8755 , \8754 , \5590 );
nor \U$8379 ( \8756 , \8753 , \8755 );
not \U$8380 ( \8757 , \8756 );
and \U$8381 ( \8758 , \6172 , RIae76a78_55);
and \U$8382 ( \8759 , RIae76988_53, \6170 );
nor \U$8383 ( \8760 , \8758 , \8759 );
and \U$8384 ( \8761 , \8760 , \6175 );
not \U$8385 ( \8762 , \8760 );
and \U$8386 ( \8763 , \8762 , \6176 );
nor \U$8387 ( \8764 , \8761 , \8763 );
not \U$8388 ( \8765 , \8764 );
and \U$8389 ( \8766 , \8757 , \8765 );
and \U$8390 ( \8767 , \8764 , \8756 );
and \U$8391 ( \8768 , \6941 , RIae767a8_49);
and \U$8392 ( \8769 , RIae76898_51, \6939 );
nor \U$8393 ( \8770 , \8768 , \8769 );
and \U$8394 ( \8771 , \8770 , \6945 );
not \U$8395 ( \8772 , \8770 );
and \U$8396 ( \8773 , \8772 , \6314 );
nor \U$8397 ( \8774 , \8771 , \8773 );
nor \U$8398 ( \8775 , \8767 , \8774 );
nor \U$8399 ( \8776 , \8766 , \8775 );
not \U$8400 ( \8777 , \8776 );
and \U$8401 ( \8778 , \8749 , \8777 );
and \U$8402 ( \8779 , \8748 , \8776 );
and \U$8403 ( \8780 , \8371 , RIae78cb0_128);
and \U$8404 ( \8781 , RIae78da0_130, \8369 );
nor \U$8405 ( \8782 , \8780 , \8781 );
and \U$8406 ( \8783 , \8782 , \8020 );
not \U$8407 ( \8784 , \8782 );
and \U$8408 ( \8785 , \8784 , \8019 );
nor \U$8409 ( \8786 , \8783 , \8785 );
not \U$8410 ( \8787 , \8786 );
nand \U$8411 ( \8788 , RIae7a510_180, RIae7a600_182);
and \U$8412 ( \8789 , \8788 , RIae7a3a8_177);
nand \U$8413 ( \8790 , \8787 , \8789 );
and \U$8414 ( \8791 , \7633 , RIae76b68_57);
and \U$8415 ( \8792 , RIae78a58_123, \7631 );
nor \U$8416 ( \8793 , \8791 , \8792 );
and \U$8417 ( \8794 , \8793 , \7206 );
not \U$8418 ( \8795 , \8793 );
and \U$8419 ( \8796 , \8795 , \7205 );
nor \U$8420 ( \8797 , \8794 , \8796 );
and \U$8421 ( \8798 , \8790 , \8797 );
not \U$8422 ( \8799 , \8789 );
and \U$8423 ( \8800 , \8799 , \8786 );
nor \U$8424 ( \8801 , \8798 , \8800 );
nor \U$8425 ( \8802 , \8779 , \8801 );
nor \U$8426 ( \8803 , \8778 , \8802 );
nor \U$8427 ( \8804 , \8723 , \8803 );
nor \U$8428 ( \8805 , \8722 , \8804 );
xor \U$8429 ( \8806 , \8462 , \8463 );
xor \U$8430 ( \8807 , \8806 , \8472 );
not \U$8431 ( \8808 , \8807 );
xor \U$8432 ( \8809 , \8486 , \8493 );
xor \U$8433 ( \8810 , \8809 , \8502 );
not \U$8434 ( \8811 , \8810 );
and \U$8435 ( \8812 , \8808 , \8811 );
and \U$8436 ( \8813 , \8810 , \8807 );
xor \U$8437 ( \8814 , \8279 , \8286 );
xor \U$8438 ( \8815 , \8814 , \8294 );
nor \U$8439 ( \8816 , \8813 , \8815 );
nor \U$8440 ( \8817 , \8812 , \8816 );
not \U$8441 ( \8818 , \8817 );
xor \U$8442 ( \8819 , \8364 , \8376 );
xor \U$8443 ( \8820 , \8819 , \8384 );
not \U$8444 ( \8821 , \8820 );
xor \U$8445 ( \8822 , \8423 , \8430 );
xor \U$8446 ( \8823 , \8822 , \8438 );
nand \U$8447 ( \8824 , \8821 , \8823 );
not \U$8448 ( \8825 , \8824 );
and \U$8449 ( \8826 , \8818 , \8825 );
and \U$8450 ( \8827 , \8817 , \8824 );
xor \U$8451 ( \8828 , \8394 , \8401 );
xor \U$8452 ( \8829 , \8828 , \8409 );
xor \U$8453 ( \8830 , \8337 , \8344 );
xor \U$8454 ( \8831 , \8830 , \8352 );
and \U$8455 ( \8832 , \8829 , \8831 );
not \U$8456 ( \8833 , \8304 );
xor \U$8457 ( \8834 , \8313 , \8324 );
not \U$8458 ( \8835 , \8834 );
or \U$8459 ( \8836 , \8833 , \8835 );
or \U$8460 ( \8837 , \8834 , \8304 );
nand \U$8461 ( \8838 , \8836 , \8837 );
xor \U$8462 ( \8839 , \8337 , \8344 );
xor \U$8463 ( \8840 , \8839 , \8352 );
and \U$8464 ( \8841 , \8838 , \8840 );
and \U$8465 ( \8842 , \8829 , \8838 );
or \U$8466 ( \8843 , \8832 , \8841 , \8842 );
not \U$8467 ( \8844 , \8843 );
nor \U$8468 ( \8845 , \8827 , \8844 );
nor \U$8469 ( \8846 , \8826 , \8845 );
xor \U$8470 ( \8847 , \8805 , \8846 );
xor \U$8471 ( \8848 , \8237 , \8239 );
xor \U$8472 ( \8849 , \8848 , \8242 );
xor \U$8473 ( \8850 , \8017 , \8020 );
xor \U$8474 ( \8851 , \8850 , \8028 );
xor \U$8475 ( \8852 , \8849 , \8851 );
xor \U$8476 ( \8853 , \7963 , \7971 );
xor \U$8477 ( \8854 , \8853 , \7979 );
xor \U$8478 ( \8855 , \8254 , \8263 );
xor \U$8479 ( \8856 , \8854 , \8855 );
and \U$8480 ( \8857 , \8852 , \8856 );
and \U$8481 ( \8858 , \8849 , \8851 );
nor \U$8482 ( \8859 , \8857 , \8858 );
xor \U$8483 ( \8860 , \8847 , \8859 );
xor \U$8484 ( \8861 , \8010 , \8031 );
xor \U$8485 ( \8862 , \8861 , \8057 );
not \U$8486 ( \8863 , \8862 );
not \U$8487 ( \8864 , \8505 );
not \U$8488 ( \8865 , \8475 );
or \U$8489 ( \8866 , \8864 , \8865 );
or \U$8490 ( \8867 , \8475 , \8505 );
nand \U$8491 ( \8868 , \8866 , \8867 );
not \U$8492 ( \8869 , \8868 );
not \U$8493 ( \8870 , \8454 );
and \U$8494 ( \8871 , \8869 , \8870 );
and \U$8495 ( \8872 , \8868 , \8454 );
nor \U$8496 ( \8873 , \8871 , \8872 );
not \U$8497 ( \8874 , \8873 );
not \U$8498 ( \8875 , \8355 );
not \U$8499 ( \8876 , \8326 );
or \U$8500 ( \8877 , \8875 , \8876 );
or \U$8501 ( \8878 , \8326 , \8355 );
nand \U$8502 ( \8879 , \8877 , \8878 );
not \U$8503 ( \8880 , \8879 );
not \U$8504 ( \8881 , \8297 );
and \U$8505 ( \8882 , \8880 , \8881 );
and \U$8506 ( \8883 , \8879 , \8297 );
nor \U$8507 ( \8884 , \8882 , \8883 );
not \U$8508 ( \8885 , \8884 );
and \U$8509 ( \8886 , \8874 , \8885 );
and \U$8510 ( \8887 , \8873 , \8884 );
not \U$8511 ( \8888 , \8441 );
not \U$8512 ( \8889 , \8387 );
or \U$8513 ( \8890 , \8888 , \8889 );
or \U$8514 ( \8891 , \8387 , \8441 );
nand \U$8515 ( \8892 , \8890 , \8891 );
not \U$8516 ( \8893 , \8892 );
not \U$8517 ( \8894 , \8412 );
and \U$8518 ( \8895 , \8893 , \8894 );
and \U$8519 ( \8896 , \8892 , \8412 );
nor \U$8520 ( \8897 , \8895 , \8896 );
nor \U$8521 ( \8898 , \8887 , \8897 );
nor \U$8522 ( \8899 , \8886 , \8898 );
not \U$8523 ( \8900 , \8899 );
or \U$8524 ( \8901 , \8863 , \8900 );
or \U$8525 ( \8902 , \8899 , \8862 );
nand \U$8526 ( \8903 , \8901 , \8902 );
not \U$8527 ( \8904 , \8903 );
xor \U$8528 ( \8905 , \8088 , \8117 );
xor \U$8529 ( \8906 , \8905 , \8146 );
not \U$8530 ( \8907 , \8906 );
and \U$8531 ( \8908 , \8904 , \8907 );
and \U$8532 ( \8909 , \8903 , \8906 );
nor \U$8533 ( \8910 , \8908 , \8909 );
xnor \U$8534 ( \8911 , \8860 , \8910 );
not \U$8535 ( \8912 , \8911 );
xor \U$8536 ( \8913 , \8245 , \8247 );
xor \U$8537 ( \8914 , \8913 , \8268 );
xor \U$8538 ( \8915 , \8357 , \8443 );
xor \U$8539 ( \8916 , \8915 , \8507 );
xor \U$8540 ( \8917 , \7919 , \7921 );
xor \U$8541 ( \8918 , \8917 , \7924 );
xor \U$8542 ( \8919 , \8513 , \8520 );
xor \U$8543 ( \8920 , \8918 , \8919 );
xor \U$8544 ( \8921 , \8916 , \8920 );
xor \U$8545 ( \8922 , \8914 , \8921 );
not \U$8546 ( \8923 , \8922 );
and \U$8547 ( \8924 , \8912 , \8923 );
and \U$8548 ( \8925 , \8911 , \8922 );
nor \U$8549 ( \8926 , \8924 , \8925 );
and \U$8550 ( \8927 , \5896 , RIae76028_33);
and \U$8551 ( \8928 , RIae762f8_39, \5894 );
nor \U$8552 ( \8929 , \8927 , \8928 );
and \U$8553 ( \8930 , \8929 , \5590 );
not \U$8554 ( \8931 , \8929 );
and \U$8555 ( \8932 , \8931 , \5589 );
nor \U$8556 ( \8933 , \8930 , \8932 );
and \U$8557 ( \8934 , \6172 , RIae76208_37);
and \U$8558 ( \8935 , RIae76a78_55, \6170 );
nor \U$8559 ( \8936 , \8934 , \8935 );
and \U$8560 ( \8937 , \8936 , \6176 );
not \U$8561 ( \8938 , \8936 );
and \U$8562 ( \8939 , \8938 , \6175 );
nor \U$8563 ( \8940 , \8937 , \8939 );
xor \U$8564 ( \8941 , \8933 , \8940 );
and \U$8565 ( \8942 , \6941 , RIae76988_53);
and \U$8566 ( \8943 , RIae767a8_49, \6939 );
nor \U$8567 ( \8944 , \8942 , \8943 );
and \U$8568 ( \8945 , \8944 , \6314 );
not \U$8569 ( \8946 , \8944 );
and \U$8570 ( \8947 , \8946 , \6945 );
nor \U$8571 ( \8948 , \8945 , \8947 );
and \U$8572 ( \8949 , \8941 , \8948 );
and \U$8573 ( \8950 , \8933 , \8940 );
or \U$8574 ( \8951 , \8949 , \8950 );
and \U$8575 ( \8952 , \7633 , RIae76898_51);
and \U$8576 ( \8953 , RIae76b68_57, \7631 );
nor \U$8577 ( \8954 , \8952 , \8953 );
and \U$8578 ( \8955 , \8954 , \7206 );
not \U$8579 ( \8956 , \8954 );
and \U$8580 ( \8957 , \8956 , \7205 );
nor \U$8581 ( \8958 , \8955 , \8957 );
and \U$8582 ( \8959 , RIae7a3a8_177, RIae7a600_182);
not \U$8583 ( \8960 , RIae7a510_180);
and \U$8584 ( \8961 , RIae7a600_182, \8960 );
not \U$8585 ( \8962 , RIae7a600_182);
and \U$8586 ( \8963 , \8962 , RIae7a510_180);
or \U$8587 ( \8964 , \8961 , \8963 );
nor \U$8588 ( \8965 , RIae7a3a8_177, RIae7a600_182);
nor \U$8589 ( \8966 , \8959 , \8964 , \8965 );
nand \U$8590 ( \8967 , RIae78da0_130, \8966 );
and \U$8591 ( \8968 , \8967 , \8799 );
not \U$8592 ( \8969 , \8967 );
and \U$8593 ( \8970 , \8969 , \8789 );
nor \U$8594 ( \8971 , \8968 , \8970 );
xor \U$8595 ( \8972 , \8958 , \8971 );
and \U$8596 ( \8973 , \8371 , RIae78a58_123);
and \U$8597 ( \8974 , RIae78cb0_128, \8369 );
nor \U$8598 ( \8975 , \8973 , \8974 );
and \U$8599 ( \8976 , \8975 , \8020 );
not \U$8600 ( \8977 , \8975 );
and \U$8601 ( \8978 , \8977 , \8019 );
nor \U$8602 ( \8979 , \8976 , \8978 );
and \U$8603 ( \8980 , \8972 , \8979 );
and \U$8604 ( \8981 , \8958 , \8971 );
or \U$8605 ( \8982 , \8980 , \8981 );
xor \U$8606 ( \8983 , \8951 , \8982 );
and \U$8607 ( \8984 , \4247 , RIae753f8_7);
and \U$8608 ( \8985 , RIae763e8_41, \4245 );
nor \U$8609 ( \8986 , \8984 , \8985 );
and \U$8610 ( \8987 , \8986 , \3989 );
not \U$8611 ( \8988 , \8986 );
and \U$8612 ( \8989 , \8988 , \4251 );
nor \U$8613 ( \8990 , \8987 , \8989 );
and \U$8614 ( \8991 , \4688 , RIae764d8_43);
and \U$8615 ( \8992 , RIae766b8_47, \4686 );
nor \U$8616 ( \8993 , \8991 , \8992 );
and \U$8617 ( \8994 , \8993 , \4481 );
not \U$8618 ( \8995 , \8993 );
and \U$8619 ( \8996 , \8995 , \4482 );
nor \U$8620 ( \8997 , \8994 , \8996 );
xor \U$8621 ( \8998 , \8990 , \8997 );
and \U$8622 ( \8999 , \5399 , RIae765c8_45);
and \U$8623 ( \9000 , RIae76118_35, \5397 );
nor \U$8624 ( \9001 , \8999 , \9000 );
and \U$8625 ( \9002 , \9001 , \5016 );
not \U$8626 ( \9003 , \9001 );
and \U$8627 ( \9004 , \9003 , \5403 );
nor \U$8628 ( \9005 , \9002 , \9004 );
and \U$8629 ( \9006 , \8998 , \9005 );
and \U$8630 ( \9007 , \8990 , \8997 );
or \U$8631 ( \9008 , \9006 , \9007 );
and \U$8632 ( \9009 , \8983 , \9008 );
and \U$8633 ( \9010 , \8951 , \8982 );
or \U$8634 ( \9011 , \9009 , \9010 );
and \U$8635 ( \9012 , \558 , RIae78530_112);
and \U$8636 ( \9013 , RIae77c48_93, \556 );
nor \U$8637 ( \9014 , \9012 , \9013 );
and \U$8638 ( \9015 , \9014 , \504 );
not \U$8639 ( \9016 , \9014 );
and \U$8640 ( \9017 , \9016 , \562 );
nor \U$8641 ( \9018 , \9015 , \9017 );
and \U$8642 ( \9019 , \672 , RIae77b58_91);
and \U$8643 ( \9020 , RIae77d38_95, \670 );
nor \U$8644 ( \9021 , \9019 , \9020 );
and \U$8645 ( \9022 , \9021 , \588 );
not \U$8646 ( \9023 , \9021 );
and \U$8647 ( \9024 , \9023 , \587 );
nor \U$8648 ( \9025 , \9022 , \9024 );
xor \U$8649 ( \9026 , \9018 , \9025 );
not \U$8650 ( \9027 , \789 );
and \U$8651 ( \9028 , \883 , RIae77e28_97);
and \U$8652 ( \9029 , RIae78968_121, \881 );
nor \U$8653 ( \9030 , \9028 , \9029 );
not \U$8654 ( \9031 , \9030 );
or \U$8655 ( \9032 , \9027 , \9031 );
or \U$8656 ( \9033 , \9030 , \789 );
nand \U$8657 ( \9034 , \9032 , \9033 );
and \U$8658 ( \9035 , \9026 , \9034 );
and \U$8659 ( \9036 , \9018 , \9025 );
or \U$8660 ( \9037 , \9035 , \9036 );
nand \U$8661 ( \9038 , RIae782d8_107, RIae78b48_125);
not \U$8662 ( \9039 , \9038 );
xor \U$8663 ( \9040 , \9037 , \9039 );
not \U$8664 ( \9041 , \392 );
and \U$8665 ( \9042 , \384 , RIae780f8_103);
and \U$8666 ( \9043 , RIae77f18_99, \382 );
nor \U$8667 ( \9044 , \9042 , \9043 );
not \U$8668 ( \9045 , \9044 );
or \U$8669 ( \9046 , \9041 , \9045 );
or \U$8670 ( \9047 , \9044 , \388 );
nand \U$8671 ( \9048 , \9046 , \9047 );
not \U$8672 ( \9049 , \400 );
and \U$8673 ( \9050 , \436 , RIae78008_101);
and \U$8674 ( \9051 , RIae781e8_105, \434 );
nor \U$8675 ( \9052 , \9050 , \9051 );
not \U$8676 ( \9053 , \9052 );
or \U$8677 ( \9054 , \9049 , \9053 );
or \U$8678 ( \9055 , \9052 , \400 );
nand \U$8679 ( \9056 , \9054 , \9055 );
xor \U$8680 ( \9057 , \9048 , \9056 );
not \U$8681 ( \9058 , \469 );
and \U$8682 ( \9059 , \514 , RIae785a8_113);
and \U$8683 ( \9060 , RIae783c8_109, \512 );
nor \U$8684 ( \9061 , \9059 , \9060 );
not \U$8685 ( \9062 , \9061 );
or \U$8686 ( \9063 , \9058 , \9062 );
or \U$8687 ( \9064 , \9061 , \469 );
nand \U$8688 ( \9065 , \9063 , \9064 );
and \U$8689 ( \9066 , \9057 , \9065 );
and \U$8690 ( \9067 , \9048 , \9056 );
or \U$8691 ( \9068 , \9066 , \9067 );
and \U$8692 ( \9069 , \9040 , \9068 );
and \U$8693 ( \9070 , \9037 , \9039 );
or \U$8694 ( \9071 , \9069 , \9070 );
xor \U$8695 ( \9072 , \9011 , \9071 );
and \U$8696 ( \9073 , \2607 , RIae75d58_27);
and \U$8697 ( \9074 , RIae755d8_11, \2605 );
nor \U$8698 ( \9075 , \9073 , \9074 );
and \U$8699 ( \9076 , \9075 , \2611 );
not \U$8700 ( \9077 , \9075 );
and \U$8701 ( \9078 , \9077 , \2397 );
nor \U$8702 ( \9079 , \9076 , \9078 );
and \U$8703 ( \9080 , \1939 , RIae758a8_17);
and \U$8704 ( \9081 , RIae75f38_31, \1937 );
nor \U$8705 ( \9082 , \9080 , \9081 );
and \U$8706 ( \9083 , \9082 , \1735 );
not \U$8707 ( \9084 , \9082 );
and \U$8708 ( \9085 , \9084 , \1734 );
nor \U$8709 ( \9086 , \9083 , \9085 );
xor \U$8710 ( \9087 , \9079 , \9086 );
and \U$8711 ( \9088 , \2224 , RIae75e48_29);
and \U$8712 ( \9089 , RIae75c68_25, \2222 );
nor \U$8713 ( \9090 , \9088 , \9089 );
and \U$8714 ( \9091 , \9090 , \2061 );
not \U$8715 ( \9092 , \9090 );
and \U$8716 ( \9093 , \9092 , \2060 );
nor \U$8717 ( \9094 , \9091 , \9093 );
and \U$8718 ( \9095 , \9087 , \9094 );
and \U$8719 ( \9096 , \9079 , \9086 );
or \U$8720 ( \9097 , \9095 , \9096 );
and \U$8721 ( \9098 , \1138 , RIae78878_119);
and \U$8722 ( \9099 , RIae78788_117, \1136 );
nor \U$8723 ( \9100 , \9098 , \9099 );
and \U$8724 ( \9101 , \9100 , \1012 );
not \U$8725 ( \9102 , \9100 );
and \U$8726 ( \9103 , \9102 , \1142 );
nor \U$8727 ( \9104 , \9101 , \9103 );
and \U$8728 ( \9105 , \1376 , RIae78698_115);
and \U$8729 ( \9106 , RIae75b78_23, \1374 );
nor \U$8730 ( \9107 , \9105 , \9106 );
and \U$8731 ( \9108 , \9107 , \1380 );
not \U$8732 ( \9109 , \9107 );
and \U$8733 ( \9110 , \9109 , \1261 );
nor \U$8734 ( \9111 , \9108 , \9110 );
xor \U$8735 ( \9112 , \9104 , \9111 );
and \U$8736 ( \9113 , \1593 , RIae75a88_21);
and \U$8737 ( \9114 , RIae75998_19, \1591 );
nor \U$8738 ( \9115 , \9113 , \9114 );
and \U$8739 ( \9116 , \9115 , \1498 );
not \U$8740 ( \9117 , \9115 );
and \U$8741 ( \9118 , \9117 , \1488 );
nor \U$8742 ( \9119 , \9116 , \9118 );
and \U$8743 ( \9120 , \9112 , \9119 );
and \U$8744 ( \9121 , \9104 , \9111 );
or \U$8745 ( \9122 , \9120 , \9121 );
xor \U$8746 ( \9123 , \9097 , \9122 );
and \U$8747 ( \9124 , \3730 , RIae75128_1);
and \U$8748 ( \9125 , RIae75308_5, \3728 );
nor \U$8749 ( \9126 , \9124 , \9125 );
and \U$8750 ( \9127 , \9126 , \3732 );
not \U$8751 ( \9128 , \9126 );
and \U$8752 ( \9129 , \9128 , \3422 );
nor \U$8753 ( \9130 , \9127 , \9129 );
not \U$8754 ( \9131 , \3089 );
and \U$8755 ( \9132 , \2783 , RIae754e8_9);
and \U$8756 ( \9133 , RIae757b8_15, \2781 );
nor \U$8757 ( \9134 , \9132 , \9133 );
not \U$8758 ( \9135 , \9134 );
or \U$8759 ( \9136 , \9131 , \9135 );
or \U$8760 ( \9137 , \9134 , \2789 );
nand \U$8761 ( \9138 , \9136 , \9137 );
xor \U$8762 ( \9139 , \9130 , \9138 );
not \U$8763 ( \9140 , \2774 );
and \U$8764 ( \9141 , \3214 , RIae756c8_13);
and \U$8765 ( \9142 , RIae75218_3, \3212 );
nor \U$8766 ( \9143 , \9141 , \9142 );
not \U$8767 ( \9144 , \9143 );
or \U$8768 ( \9145 , \9140 , \9144 );
or \U$8769 ( \9146 , \9143 , \3218 );
nand \U$8770 ( \9147 , \9145 , \9146 );
and \U$8771 ( \9148 , \9139 , \9147 );
and \U$8772 ( \9149 , \9130 , \9138 );
or \U$8773 ( \9150 , \9148 , \9149 );
and \U$8774 ( \9151 , \9123 , \9150 );
and \U$8775 ( \9152 , \9097 , \9122 );
or \U$8776 ( \9153 , \9151 , \9152 );
xor \U$8777 ( \9154 , \9072 , \9153 );
xor \U$8778 ( \9155 , \8730 , \8737 );
xor \U$8779 ( \9156 , \9155 , \8745 );
not \U$8780 ( \9157 , \8797 );
and \U$8781 ( \9158 , \8786 , \8789 );
not \U$8782 ( \9159 , \8786 );
and \U$8783 ( \9160 , \9159 , \8799 );
nor \U$8784 ( \9161 , \9158 , \9160 );
not \U$8785 ( \9162 , \9161 );
or \U$8786 ( \9163 , \9157 , \9162 );
or \U$8787 ( \9164 , \9161 , \8797 );
nand \U$8788 ( \9165 , \9163 , \9164 );
xor \U$8789 ( \9166 , \9156 , \9165 );
not \U$8790 ( \9167 , \8756 );
xor \U$8791 ( \9168 , \8764 , \8774 );
not \U$8792 ( \9169 , \9168 );
or \U$8793 ( \9170 , \9167 , \9169 );
or \U$8794 ( \9171 , \9168 , \8756 );
nand \U$8795 ( \9172 , \9170 , \9171 );
and \U$8796 ( \9173 , \9166 , \9172 );
and \U$8797 ( \9174 , \9156 , \9165 );
or \U$8798 ( \9175 , \9173 , \9174 );
not \U$8799 ( \9176 , \8696 );
xor \U$8800 ( \9177 , \8705 , \8716 );
not \U$8801 ( \9178 , \9177 );
or \U$8802 ( \9179 , \9176 , \9178 );
or \U$8803 ( \9180 , \9177 , \8696 );
nand \U$8804 ( \9181 , \9179 , \9180 );
not \U$8805 ( \9182 , RIae780f8_103);
nor \U$8806 ( \9183 , \9182 , \491 );
xor \U$8807 ( \9184 , \9181 , \9183 );
xor \U$8808 ( \9185 , \8669 , \8677 );
xor \U$8809 ( \9186 , \9185 , \8685 );
and \U$8810 ( \9187 , \9184 , \9186 );
and \U$8811 ( \9188 , \9181 , \9183 );
or \U$8812 ( \9189 , \9187 , \9188 );
xor \U$8813 ( \9190 , \9175 , \9189 );
xor \U$8814 ( \9191 , \8612 , \8619 );
xor \U$8815 ( \9192 , \9191 , \8627 );
xor \U$8816 ( \9193 , \8587 , \8594 );
xor \U$8817 ( \9194 , \9193 , \8602 );
xor \U$8818 ( \9195 , \9192 , \9194 );
xor \U$8819 ( \9196 , \8639 , \8647 );
xor \U$8820 ( \9197 , \9196 , \8655 );
and \U$8821 ( \9198 , \9195 , \9197 );
and \U$8822 ( \9199 , \9192 , \9194 );
or \U$8823 ( \9200 , \9198 , \9199 );
xor \U$8824 ( \9201 , \9190 , \9200 );
and \U$8825 ( \9202 , \9154 , \9201 );
xor \U$8826 ( \9203 , \8990 , \8997 );
xor \U$8827 ( \9204 , \9203 , \9005 );
xor \U$8828 ( \9205 , \8958 , \8971 );
xor \U$8829 ( \9206 , \9205 , \8979 );
and \U$8830 ( \9207 , \9204 , \9206 );
xor \U$8831 ( \9208 , \8933 , \8940 );
xor \U$8832 ( \9209 , \9208 , \8948 );
xor \U$8833 ( \9210 , \8958 , \8971 );
xor \U$8834 ( \9211 , \9210 , \8979 );
and \U$8835 ( \9212 , \9209 , \9211 );
and \U$8836 ( \9213 , \9204 , \9209 );
or \U$8837 ( \9214 , \9207 , \9212 , \9213 );
xor \U$8838 ( \9215 , \9018 , \9025 );
xor \U$8839 ( \9216 , \9215 , \9034 );
xor \U$8840 ( \9217 , \9216 , \9038 );
xor \U$8841 ( \9218 , \9048 , \9056 );
xor \U$8842 ( \9219 , \9218 , \9065 );
and \U$8843 ( \9220 , \9217 , \9219 );
and \U$8844 ( \9221 , \9216 , \9038 );
or \U$8845 ( \9222 , \9220 , \9221 );
xor \U$8846 ( \9223 , \9214 , \9222 );
xor \U$8847 ( \9224 , \9079 , \9086 );
xor \U$8848 ( \9225 , \9224 , \9094 );
xor \U$8849 ( \9226 , \9104 , \9111 );
xor \U$8850 ( \9227 , \9226 , \9119 );
and \U$8851 ( \9228 , \9225 , \9227 );
xor \U$8852 ( \9229 , \9130 , \9138 );
xor \U$8853 ( \9230 , \9229 , \9147 );
xor \U$8854 ( \9231 , \9104 , \9111 );
xor \U$8855 ( \9232 , \9231 , \9119 );
and \U$8856 ( \9233 , \9230 , \9232 );
and \U$8857 ( \9234 , \9225 , \9230 );
or \U$8858 ( \9235 , \9228 , \9233 , \9234 );
and \U$8859 ( \9236 , \9223 , \9235 );
and \U$8860 ( \9237 , \9214 , \9222 );
or \U$8861 ( \9238 , \9236 , \9237 );
and \U$8862 ( \9239 , \5896 , RIae76118_35);
and \U$8863 ( \9240 , RIae76028_33, \5894 );
nor \U$8864 ( \9241 , \9239 , \9240 );
and \U$8865 ( \9242 , \9241 , \5590 );
not \U$8866 ( \9243 , \9241 );
and \U$8867 ( \9244 , \9243 , \5589 );
nor \U$8868 ( \9245 , \9242 , \9244 );
and \U$8869 ( \9246 , \4688 , RIae763e8_41);
and \U$8870 ( \9247 , RIae764d8_43, \4686 );
nor \U$8871 ( \9248 , \9246 , \9247 );
and \U$8872 ( \9249 , \9248 , \4481 );
not \U$8873 ( \9250 , \9248 );
and \U$8874 ( \9251 , \9250 , \4482 );
nor \U$8875 ( \9252 , \9249 , \9251 );
xor \U$8876 ( \9253 , \9245 , \9252 );
and \U$8877 ( \9254 , \5399 , RIae766b8_47);
and \U$8878 ( \9255 , RIae765c8_45, \5397 );
nor \U$8879 ( \9256 , \9254 , \9255 );
and \U$8880 ( \9257 , \9256 , \5016 );
not \U$8881 ( \9258 , \9256 );
and \U$8882 ( \9259 , \9258 , \5403 );
nor \U$8883 ( \9260 , \9257 , \9259 );
and \U$8884 ( \9261 , \9253 , \9260 );
and \U$8885 ( \9262 , \9245 , \9252 );
or \U$8886 ( \9263 , \9261 , \9262 );
and \U$8887 ( \9264 , \8966 , RIae78cb0_128);
and \U$8888 ( \9265 , RIae78da0_130, \8964 );
nor \U$8889 ( \9266 , \9264 , \9265 );
and \U$8890 ( \9267 , \9266 , \8799 );
not \U$8891 ( \9268 , \9266 );
and \U$8892 ( \9269 , \9268 , \8789 );
nor \U$8893 ( \9270 , \9267 , \9269 );
and \U$8894 ( \9271 , RIae7a588_181, RIae7a498_179);
nor \U$8895 ( \9272 , \9271 , \8960 );
not \U$8896 ( \9273 , \9272 );
xor \U$8897 ( \9274 , \9270 , \9273 );
and \U$8898 ( \9275 , \8371 , RIae76b68_57);
and \U$8899 ( \9276 , RIae78a58_123, \8369 );
nor \U$8900 ( \9277 , \9275 , \9276 );
and \U$8901 ( \9278 , \9277 , \8020 );
not \U$8902 ( \9279 , \9277 );
and \U$8903 ( \9280 , \9279 , \8019 );
nor \U$8904 ( \9281 , \9278 , \9280 );
and \U$8905 ( \9282 , \9274 , \9281 );
and \U$8906 ( \9283 , \9270 , \9273 );
or \U$8907 ( \9284 , \9282 , \9283 );
xor \U$8908 ( \9285 , \9263 , \9284 );
and \U$8909 ( \9286 , \6941 , RIae76a78_55);
and \U$8910 ( \9287 , RIae76988_53, \6939 );
nor \U$8911 ( \9288 , \9286 , \9287 );
and \U$8912 ( \9289 , \9288 , \6314 );
not \U$8913 ( \9290 , \9288 );
and \U$8914 ( \9291 , \9290 , \6945 );
nor \U$8915 ( \9292 , \9289 , \9291 );
and \U$8916 ( \9293 , \6172 , RIae762f8_39);
and \U$8917 ( \9294 , RIae76208_37, \6170 );
nor \U$8918 ( \9295 , \9293 , \9294 );
and \U$8919 ( \9296 , \9295 , \6176 );
not \U$8920 ( \9297 , \9295 );
and \U$8921 ( \9298 , \9297 , \6175 );
nor \U$8922 ( \9299 , \9296 , \9298 );
xor \U$8923 ( \9300 , \9292 , \9299 );
and \U$8924 ( \9301 , \7633 , RIae767a8_49);
and \U$8925 ( \9302 , RIae76898_51, \7631 );
nor \U$8926 ( \9303 , \9301 , \9302 );
and \U$8927 ( \9304 , \9303 , \7206 );
not \U$8928 ( \9305 , \9303 );
and \U$8929 ( \9306 , \9305 , \7205 );
nor \U$8930 ( \9307 , \9304 , \9306 );
and \U$8931 ( \9308 , \9300 , \9307 );
and \U$8932 ( \9309 , \9292 , \9299 );
or \U$8933 ( \9310 , \9308 , \9309 );
and \U$8934 ( \9311 , \9285 , \9310 );
and \U$8935 ( \9312 , \9263 , \9284 );
or \U$8936 ( \9313 , \9311 , \9312 );
and \U$8937 ( \9314 , \672 , RIae77c48_93);
and \U$8938 ( \9315 , RIae77b58_91, \670 );
nor \U$8939 ( \9316 , \9314 , \9315 );
and \U$8940 ( \9317 , \9316 , \588 );
not \U$8941 ( \9318 , \9316 );
and \U$8942 ( \9319 , \9318 , \587 );
nor \U$8943 ( \9320 , \9317 , \9319 );
not \U$8944 ( \9321 , \787 );
and \U$8945 ( \9322 , \883 , RIae77d38_95);
and \U$8946 ( \9323 , RIae77e28_97, \881 );
nor \U$8947 ( \9324 , \9322 , \9323 );
not \U$8948 ( \9325 , \9324 );
or \U$8949 ( \9326 , \9321 , \9325 );
or \U$8950 ( \9327 , \9324 , \789 );
nand \U$8951 ( \9328 , \9326 , \9327 );
xor \U$8952 ( \9329 , \9320 , \9328 );
and \U$8953 ( \9330 , \1138 , RIae78968_121);
and \U$8954 ( \9331 , RIae78878_119, \1136 );
nor \U$8955 ( \9332 , \9330 , \9331 );
and \U$8956 ( \9333 , \9332 , \1012 );
not \U$8957 ( \9334 , \9332 );
and \U$8958 ( \9335 , \9334 , \1142 );
nor \U$8959 ( \9336 , \9333 , \9335 );
and \U$8960 ( \9337 , \9329 , \9336 );
and \U$8961 ( \9338 , \9320 , \9328 );
or \U$8962 ( \9339 , \9337 , \9338 );
not \U$8963 ( \9340 , RIae772e8_73);
nor \U$8964 ( \9341 , \9340 , \491 );
not \U$8965 ( \9342 , \388 );
and \U$8966 ( \9343 , \384 , RIae782d8_107);
and \U$8967 ( \9344 , RIae780f8_103, \382 );
nor \U$8968 ( \9345 , \9343 , \9344 );
not \U$8969 ( \9346 , \9345 );
or \U$8970 ( \9347 , \9342 , \9346 );
or \U$8971 ( \9348 , \9345 , \388 );
nand \U$8972 ( \9349 , \9347 , \9348 );
and \U$8973 ( \9350 , \9341 , \9349 );
xor \U$8974 ( \9351 , \9339 , \9350 );
not \U$8975 ( \9352 , \469 );
and \U$8976 ( \9353 , \514 , RIae781e8_105);
and \U$8977 ( \9354 , RIae785a8_113, \512 );
nor \U$8978 ( \9355 , \9353 , \9354 );
not \U$8979 ( \9356 , \9355 );
or \U$8980 ( \9357 , \9352 , \9356 );
or \U$8981 ( \9358 , \9355 , \469 );
nand \U$8982 ( \9359 , \9357 , \9358 );
not \U$8983 ( \9360 , \402 );
and \U$8984 ( \9361 , \436 , RIae77f18_99);
and \U$8985 ( \9362 , RIae78008_101, \434 );
nor \U$8986 ( \9363 , \9361 , \9362 );
not \U$8987 ( \9364 , \9363 );
or \U$8988 ( \9365 , \9360 , \9364 );
or \U$8989 ( \9366 , \9363 , \402 );
nand \U$8990 ( \9367 , \9365 , \9366 );
xor \U$8991 ( \9368 , \9359 , \9367 );
and \U$8992 ( \9369 , \558 , RIae783c8_109);
and \U$8993 ( \9370 , RIae78530_112, \556 );
nor \U$8994 ( \9371 , \9369 , \9370 );
and \U$8995 ( \9372 , \9371 , \504 );
not \U$8996 ( \9373 , \9371 );
and \U$8997 ( \9374 , \9373 , \562 );
nor \U$8998 ( \9375 , \9372 , \9374 );
and \U$8999 ( \9376 , \9368 , \9375 );
and \U$9000 ( \9377 , \9359 , \9367 );
or \U$9001 ( \9378 , \9376 , \9377 );
and \U$9002 ( \9379 , \9351 , \9378 );
and \U$9003 ( \9380 , \9339 , \9350 );
or \U$9004 ( \9381 , \9379 , \9380 );
xor \U$9005 ( \9382 , \9313 , \9381 );
and \U$9006 ( \9383 , \2607 , RIae75c68_25);
and \U$9007 ( \9384 , RIae75d58_27, \2605 );
nor \U$9008 ( \9385 , \9383 , \9384 );
and \U$9009 ( \9386 , \9385 , \2611 );
not \U$9010 ( \9387 , \9385 );
and \U$9011 ( \9388 , \9387 , \2397 );
nor \U$9012 ( \9389 , \9386 , \9388 );
and \U$9013 ( \9390 , \2224 , RIae75f38_31);
and \U$9014 ( \9391 , RIae75e48_29, \2222 );
nor \U$9015 ( \9392 , \9390 , \9391 );
and \U$9016 ( \9393 , \9392 , \2061 );
not \U$9017 ( \9394 , \9392 );
and \U$9018 ( \9395 , \9394 , \2060 );
nor \U$9019 ( \9396 , \9393 , \9395 );
xor \U$9020 ( \9397 , \9389 , \9396 );
not \U$9021 ( \9398 , \3089 );
and \U$9022 ( \9399 , \2783 , RIae755d8_11);
and \U$9023 ( \9400 , RIae754e8_9, \2781 );
nor \U$9024 ( \9401 , \9399 , \9400 );
not \U$9025 ( \9402 , \9401 );
or \U$9026 ( \9403 , \9398 , \9402 );
or \U$9027 ( \9404 , \9401 , \2789 );
nand \U$9028 ( \9405 , \9403 , \9404 );
and \U$9029 ( \9406 , \9397 , \9405 );
and \U$9030 ( \9407 , \9389 , \9396 );
or \U$9031 ( \9408 , \9406 , \9407 );
and \U$9032 ( \9409 , \1939 , RIae75998_19);
and \U$9033 ( \9410 , RIae758a8_17, \1937 );
nor \U$9034 ( \9411 , \9409 , \9410 );
and \U$9035 ( \9412 , \9411 , \1735 );
not \U$9036 ( \9413 , \9411 );
and \U$9037 ( \9414 , \9413 , \1734 );
nor \U$9038 ( \9415 , \9412 , \9414 );
and \U$9039 ( \9416 , \1376 , RIae78788_117);
and \U$9040 ( \9417 , RIae78698_115, \1374 );
nor \U$9041 ( \9418 , \9416 , \9417 );
and \U$9042 ( \9419 , \9418 , \1380 );
not \U$9043 ( \9420 , \9418 );
and \U$9044 ( \9421 , \9420 , \1261 );
nor \U$9045 ( \9422 , \9419 , \9421 );
xor \U$9046 ( \9423 , \9415 , \9422 );
and \U$9047 ( \9424 , \1593 , RIae75b78_23);
and \U$9048 ( \9425 , RIae75a88_21, \1591 );
nor \U$9049 ( \9426 , \9424 , \9425 );
and \U$9050 ( \9427 , \9426 , \1498 );
not \U$9051 ( \9428 , \9426 );
and \U$9052 ( \9429 , \9428 , \1488 );
nor \U$9053 ( \9430 , \9427 , \9429 );
and \U$9054 ( \9431 , \9423 , \9430 );
and \U$9055 ( \9432 , \9415 , \9422 );
or \U$9056 ( \9433 , \9431 , \9432 );
xor \U$9057 ( \9434 , \9408 , \9433 );
and \U$9058 ( \9435 , \4247 , RIae75308_5);
and \U$9059 ( \9436 , RIae753f8_7, \4245 );
nor \U$9060 ( \9437 , \9435 , \9436 );
and \U$9061 ( \9438 , \9437 , \3989 );
not \U$9062 ( \9439 , \9437 );
and \U$9063 ( \9440 , \9439 , \4251 );
nor \U$9064 ( \9441 , \9438 , \9440 );
not \U$9065 ( \9442 , \2774 );
and \U$9066 ( \9443 , \3214 , RIae757b8_15);
and \U$9067 ( \9444 , RIae756c8_13, \3212 );
nor \U$9068 ( \9445 , \9443 , \9444 );
not \U$9069 ( \9446 , \9445 );
or \U$9070 ( \9447 , \9442 , \9446 );
or \U$9071 ( \9448 , \9445 , \2774 );
nand \U$9072 ( \9449 , \9447 , \9448 );
xor \U$9073 ( \9450 , \9441 , \9449 );
and \U$9074 ( \9451 , \3730 , RIae75218_3);
and \U$9075 ( \9452 , RIae75128_1, \3728 );
nor \U$9076 ( \9453 , \9451 , \9452 );
and \U$9077 ( \9454 , \9453 , \3732 );
not \U$9078 ( \9455 , \9453 );
and \U$9079 ( \9456 , \9455 , \3421 );
nor \U$9080 ( \9457 , \9454 , \9456 );
and \U$9081 ( \9458 , \9450 , \9457 );
and \U$9082 ( \9459 , \9441 , \9449 );
or \U$9083 ( \9460 , \9458 , \9459 );
and \U$9084 ( \9461 , \9434 , \9460 );
and \U$9085 ( \9462 , \9408 , \9433 );
or \U$9086 ( \9463 , \9461 , \9462 );
and \U$9087 ( \9464 , \9382 , \9463 );
and \U$9088 ( \9465 , \9313 , \9381 );
or \U$9089 ( \9466 , \9464 , \9465 );
xor \U$9090 ( \9467 , \9238 , \9466 );
xor \U$9091 ( \9468 , \9181 , \9183 );
xor \U$9092 ( \9469 , \9468 , \9186 );
xor \U$9093 ( \9470 , \9192 , \9194 );
xor \U$9094 ( \9471 , \9470 , \9197 );
and \U$9095 ( \9472 , \9469 , \9471 );
xor \U$9096 ( \9473 , \9156 , \9165 );
xor \U$9097 ( \9474 , \9473 , \9172 );
xor \U$9098 ( \9475 , \9192 , \9194 );
xor \U$9099 ( \9476 , \9475 , \9197 );
and \U$9100 ( \9477 , \9474 , \9476 );
and \U$9101 ( \9478 , \9469 , \9474 );
or \U$9102 ( \9479 , \9472 , \9477 , \9478 );
and \U$9103 ( \9480 , \9467 , \9479 );
and \U$9104 ( \9481 , \9238 , \9466 );
or \U$9105 ( \9482 , \9480 , \9481 );
xor \U$9106 ( \9483 , \9202 , \9482 );
xor \U$9107 ( \9484 , \9037 , \9039 );
xor \U$9108 ( \9485 , \9484 , \9068 );
xor \U$9109 ( \9486 , \8951 , \8982 );
xor \U$9110 ( \9487 , \9486 , \9008 );
xor \U$9111 ( \9488 , \9485 , \9487 );
xor \U$9112 ( \9489 , \9097 , \9122 );
xor \U$9113 ( \9490 , \9489 , \9150 );
and \U$9114 ( \9491 , \9488 , \9490 );
and \U$9115 ( \9492 , \9485 , \9487 );
or \U$9116 ( \9493 , \9491 , \9492 );
xor \U$9117 ( \9494 , \8605 , \8630 );
xor \U$9118 ( \9495 , \9494 , \8658 );
or \U$9119 ( \9496 , \8688 , \8718 );
nand \U$9120 ( \9497 , \9496 , \8719 );
xor \U$9121 ( \9498 , \9495 , \9497 );
not \U$9122 ( \9499 , \8748 );
xor \U$9123 ( \9500 , \8801 , \8776 );
not \U$9124 ( \9501 , \9500 );
or \U$9125 ( \9502 , \9499 , \9501 );
or \U$9126 ( \9503 , \9500 , \8748 );
nand \U$9127 ( \9504 , \9502 , \9503 );
xor \U$9128 ( \9505 , \9498 , \9504 );
and \U$9129 ( \9506 , \9493 , \9505 );
xor \U$9130 ( \9507 , \8337 , \8344 );
xor \U$9131 ( \9508 , \9507 , \8352 );
xor \U$9132 ( \9509 , \8829 , \8838 );
xor \U$9133 ( \9510 , \9508 , \9509 );
not \U$9134 ( \9511 , \8823 );
not \U$9135 ( \9512 , \8820 );
or \U$9136 ( \9513 , \9511 , \9512 );
or \U$9137 ( \9514 , \8820 , \8823 );
nand \U$9138 ( \9515 , \9513 , \9514 );
xor \U$9139 ( \9516 , \9510 , \9515 );
not \U$9140 ( \9517 , \8807 );
xor \U$9141 ( \9518 , \8810 , \8815 );
not \U$9142 ( \9519 , \9518 );
or \U$9143 ( \9520 , \9517 , \9519 );
or \U$9144 ( \9521 , \9518 , \8807 );
nand \U$9145 ( \9522 , \9520 , \9521 );
xor \U$9146 ( \9523 , \9516 , \9522 );
xor \U$9147 ( \9524 , \9495 , \9497 );
xor \U$9148 ( \9525 , \9524 , \9504 );
and \U$9149 ( \9526 , \9523 , \9525 );
and \U$9150 ( \9527 , \9493 , \9523 );
or \U$9151 ( \9528 , \9506 , \9526 , \9527 );
and \U$9152 ( \9529 , \9483 , \9528 );
and \U$9153 ( \9530 , \9202 , \9482 );
nor \U$9154 ( \9531 , \9529 , \9530 );
or \U$9155 ( \9532 , \8926 , \9531 );
not \U$9156 ( \9533 , \9531 );
not \U$9157 ( \9534 , \8926 );
or \U$9158 ( \9535 , \9533 , \9534 );
not \U$9159 ( \9536 , \8720 );
xor \U$9160 ( \9537 , \8803 , \8661 );
not \U$9161 ( \9538 , \9537 );
or \U$9162 ( \9539 , \9536 , \9538 );
or \U$9163 ( \9540 , \9537 , \8720 );
nand \U$9164 ( \9541 , \9539 , \9540 );
not \U$9165 ( \9542 , \8824 );
xor \U$9166 ( \9543 , \8844 , \8817 );
not \U$9167 ( \9544 , \9543 );
or \U$9168 ( \9545 , \9542 , \9544 );
or \U$9169 ( \9546 , \9543 , \8824 );
nand \U$9170 ( \9547 , \9545 , \9546 );
xor \U$9171 ( \9548 , \9541 , \9547 );
not \U$9172 ( \9549 , \9548 );
xor \U$9173 ( \9550 , \9175 , \9189 );
and \U$9174 ( \9551 , \9550 , \9200 );
and \U$9175 ( \9552 , \9175 , \9189 );
or \U$9176 ( \9553 , \9551 , \9552 );
xor \U$9177 ( \9554 , \9011 , \9071 );
and \U$9178 ( \9555 , \9554 , \9153 );
and \U$9179 ( \9556 , \9011 , \9071 );
or \U$9180 ( \9557 , \9555 , \9556 );
xor \U$9181 ( \9558 , \9553 , \9557 );
xor \U$9182 ( \9559 , \9510 , \9515 );
and \U$9183 ( \9560 , \9559 , \9522 );
and \U$9184 ( \9561 , \9510 , \9515 );
or \U$9185 ( \9562 , \9560 , \9561 );
xor \U$9186 ( \9563 , \9558 , \9562 );
not \U$9187 ( \9564 , \9563 );
or \U$9188 ( \9565 , \9549 , \9564 );
or \U$9189 ( \9566 , \9563 , \9548 );
not \U$9190 ( \9567 , \8873 );
xor \U$9191 ( \9568 , \8897 , \8884 );
not \U$9192 ( \9569 , \9568 );
or \U$9193 ( \9570 , \9567 , \9569 );
or \U$9194 ( \9571 , \9568 , \8873 );
nand \U$9195 ( \9572 , \9570 , \9571 );
xor \U$9196 ( \9573 , \9495 , \9497 );
and \U$9197 ( \9574 , \9573 , \9504 );
and \U$9198 ( \9575 , \9495 , \9497 );
or \U$9199 ( \9576 , \9574 , \9575 );
xor \U$9200 ( \9577 , \9572 , \9576 );
xor \U$9201 ( \9578 , \8849 , \8851 );
xor \U$9202 ( \9579 , \9578 , \8856 );
xor \U$9203 ( \9580 , \9577 , \9579 );
nand \U$9204 ( \9581 , \9566 , \9580 );
nand \U$9205 ( \9582 , \9565 , \9581 );
nand \U$9206 ( \9583 , \9535 , \9582 );
nand \U$9207 ( \9584 , \9532 , \9583 );
xor \U$9208 ( \9585 , \8805 , \8846 );
and \U$9209 ( \9586 , \9585 , \8859 );
and \U$9210 ( \9587 , \8805 , \8846 );
nor \U$9211 ( \9588 , \9586 , \9587 );
not \U$9212 ( \9589 , \8906 );
nor \U$9213 ( \9590 , \9589 , \8862 );
or \U$9214 ( \9591 , \8899 , \9590 );
not \U$9215 ( \9592 , \8906 );
nand \U$9216 ( \9593 , \9592 , \8862 );
nand \U$9217 ( \9594 , \9591 , \9593 );
xor \U$9218 ( \9595 , \9588 , \9594 );
xor \U$9219 ( \9596 , \8245 , \8247 );
xor \U$9220 ( \9597 , \9596 , \8268 );
and \U$9221 ( \9598 , \8916 , \9597 );
xor \U$9222 ( \9599 , \8245 , \8247 );
xor \U$9223 ( \9600 , \9599 , \8268 );
and \U$9224 ( \9601 , \8920 , \9600 );
and \U$9225 ( \9602 , \8916 , \8920 );
or \U$9226 ( \9603 , \9598 , \9601 , \9602 );
xor \U$9227 ( \9604 , \9595 , \9603 );
xor \U$9228 ( \9605 , \9584 , \9604 );
or \U$9229 ( \9606 , \8910 , \8860 );
not \U$9230 ( \9607 , \8860 );
not \U$9231 ( \9608 , \8910 );
or \U$9232 ( \9609 , \9607 , \9608 );
nand \U$9233 ( \9610 , \9609 , \8922 );
nand \U$9234 ( \9611 , \9606 , \9610 );
and \U$9235 ( \9612 , \9541 , \9547 );
not \U$9236 ( \9613 , \9612 );
xor \U$9237 ( \9614 , \9553 , \9557 );
and \U$9238 ( \9615 , \9614 , \9562 );
and \U$9239 ( \9616 , \9553 , \9557 );
or \U$9240 ( \9617 , \9615 , \9616 );
not \U$9241 ( \9618 , \9617 );
or \U$9242 ( \9619 , \9613 , \9618 );
or \U$9243 ( \9620 , \9617 , \9612 );
xor \U$9244 ( \9621 , \9572 , \9576 );
and \U$9245 ( \9622 , \9621 , \9579 );
and \U$9246 ( \9623 , \9572 , \9576 );
or \U$9247 ( \9624 , \9622 , \9623 );
nand \U$9248 ( \9625 , \9620 , \9624 );
nand \U$9249 ( \9626 , \9619 , \9625 );
xor \U$9250 ( \9627 , \9611 , \9626 );
xor \U$9251 ( \9628 , \8271 , \8510 );
xor \U$9252 ( \9629 , \9628 , \8525 );
xor \U$9253 ( \9630 , \7985 , \8060 );
xor \U$9254 ( \9631 , \9630 , \8149 );
xor \U$9255 ( \9632 , \8175 , \8177 );
xor \U$9256 ( \9633 , \9632 , \8180 );
xor \U$9257 ( \9634 , \8533 , \8540 );
xor \U$9258 ( \9635 , \9633 , \9634 );
xor \U$9259 ( \9636 , \9631 , \9635 );
xor \U$9260 ( \9637 , \9629 , \9636 );
xor \U$9261 ( \9638 , \9627 , \9637 );
and \U$9262 ( \9639 , \9605 , \9638 );
and \U$9263 ( \9640 , \9584 , \9604 );
or \U$9264 ( \9641 , \9639 , \9640 );
xor \U$9265 ( \9642 , \9611 , \9626 );
and \U$9266 ( \9643 , \9642 , \9637 );
and \U$9267 ( \9644 , \9611 , \9626 );
or \U$9268 ( \9645 , \9643 , \9644 );
xor \U$9269 ( \9646 , \8528 , \8530 );
xor \U$9270 ( \9647 , \9646 , \8545 );
xor \U$9271 ( \9648 , \9645 , \9647 );
xor \U$9272 ( \9649 , \9588 , \9594 );
and \U$9273 ( \9650 , \9649 , \9603 );
and \U$9274 ( \9651 , \9588 , \9594 );
or \U$9275 ( \9652 , \9650 , \9651 );
xor \U$9276 ( \9653 , \8271 , \8510 );
xor \U$9277 ( \9654 , \9653 , \8525 );
and \U$9278 ( \9655 , \9631 , \9654 );
xor \U$9279 ( \9656 , \8271 , \8510 );
xor \U$9280 ( \9657 , \9656 , \8525 );
and \U$9281 ( \9658 , \9635 , \9657 );
and \U$9282 ( \9659 , \9631 , \9635 );
or \U$9283 ( \9660 , \9655 , \9658 , \9659 );
xor \U$9284 ( \9661 , \9652 , \9660 );
xor \U$9285 ( \9662 , \8183 , \8185 );
xor \U$9286 ( \9663 , \9662 , \8190 );
xor \U$9287 ( \9664 , \8550 , \8555 );
xor \U$9288 ( \9665 , \9663 , \9664 );
xor \U$9289 ( \9666 , \9661 , \9665 );
xor \U$9290 ( \9667 , \9648 , \9666 );
xor \U$9291 ( \9668 , \9641 , \9667 );
xor \U$9292 ( \9669 , \9584 , \9604 );
xor \U$9293 ( \9670 , \9669 , \9638 );
not \U$9294 ( \9671 , \9670 );
xor \U$9295 ( \9672 , \9154 , \9201 );
xor \U$9296 ( \9673 , \9238 , \9466 );
xor \U$9297 ( \9674 , \9673 , \9479 );
and \U$9298 ( \9675 , \9672 , \9674 );
xor \U$9299 ( \9676 , \9495 , \9497 );
xor \U$9300 ( \9677 , \9676 , \9504 );
xor \U$9301 ( \9678 , \9493 , \9523 );
xor \U$9302 ( \9679 , \9677 , \9678 );
xor \U$9303 ( \9680 , \9238 , \9466 );
xor \U$9304 ( \9681 , \9680 , \9479 );
and \U$9305 ( \9682 , \9679 , \9681 );
and \U$9306 ( \9683 , \9672 , \9679 );
or \U$9307 ( \9684 , \9675 , \9682 , \9683 );
xor \U$9308 ( \9685 , \9245 , \9252 );
xor \U$9309 ( \9686 , \9685 , \9260 );
xor \U$9310 ( \9687 , \9270 , \9273 );
xor \U$9311 ( \9688 , \9687 , \9281 );
and \U$9312 ( \9689 , \9686 , \9688 );
xor \U$9313 ( \9690 , \9292 , \9299 );
xor \U$9314 ( \9691 , \9690 , \9307 );
xor \U$9315 ( \9692 , \9270 , \9273 );
xor \U$9316 ( \9693 , \9692 , \9281 );
and \U$9317 ( \9694 , \9691 , \9693 );
and \U$9318 ( \9695 , \9686 , \9691 );
or \U$9319 ( \9696 , \9689 , \9694 , \9695 );
xor \U$9320 ( \9697 , \9359 , \9367 );
xor \U$9321 ( \9698 , \9697 , \9375 );
xor \U$9322 ( \9699 , \9341 , \9349 );
xor \U$9323 ( \9700 , \9698 , \9699 );
xor \U$9324 ( \9701 , \9320 , \9328 );
xor \U$9325 ( \9702 , \9701 , \9336 );
and \U$9326 ( \9703 , \9700 , \9702 );
and \U$9327 ( \9704 , \9698 , \9699 );
or \U$9328 ( \9705 , \9703 , \9704 );
xor \U$9329 ( \9706 , \9696 , \9705 );
xor \U$9330 ( \9707 , \9415 , \9422 );
xor \U$9331 ( \9708 , \9707 , \9430 );
xor \U$9332 ( \9709 , \9389 , \9396 );
xor \U$9333 ( \9710 , \9709 , \9405 );
and \U$9334 ( \9711 , \9708 , \9710 );
xor \U$9335 ( \9712 , \9441 , \9449 );
xor \U$9336 ( \9713 , \9712 , \9457 );
xor \U$9337 ( \9714 , \9389 , \9396 );
xor \U$9338 ( \9715 , \9714 , \9405 );
and \U$9339 ( \9716 , \9713 , \9715 );
and \U$9340 ( \9717 , \9708 , \9713 );
or \U$9341 ( \9718 , \9711 , \9716 , \9717 );
and \U$9342 ( \9719 , \9706 , \9718 );
and \U$9343 ( \9720 , \9696 , \9705 );
or \U$9344 ( \9721 , \9719 , \9720 );
and \U$9345 ( \9722 , \4688 , RIae753f8_7);
and \U$9346 ( \9723 , RIae763e8_41, \4686 );
nor \U$9347 ( \9724 , \9722 , \9723 );
and \U$9348 ( \9725 , \9724 , \4481 );
not \U$9349 ( \9726 , \9724 );
and \U$9350 ( \9727 , \9726 , \4482 );
nor \U$9351 ( \9728 , \9725 , \9727 );
and \U$9352 ( \9729 , \5399 , RIae764d8_43);
and \U$9353 ( \9730 , RIae766b8_47, \5397 );
nor \U$9354 ( \9731 , \9729 , \9730 );
and \U$9355 ( \9732 , \9731 , \5016 );
not \U$9356 ( \9733 , \9731 );
and \U$9357 ( \9734 , \9733 , \5403 );
nor \U$9358 ( \9735 , \9732 , \9734 );
xor \U$9359 ( \9736 , \9728 , \9735 );
and \U$9360 ( \9737 , \5896 , RIae765c8_45);
and \U$9361 ( \9738 , RIae76118_35, \5894 );
nor \U$9362 ( \9739 , \9737 , \9738 );
and \U$9363 ( \9740 , \9739 , \5590 );
not \U$9364 ( \9741 , \9739 );
and \U$9365 ( \9742 , \9741 , \5589 );
nor \U$9366 ( \9743 , \9740 , \9742 );
and \U$9367 ( \9744 , \9736 , \9743 );
and \U$9368 ( \9745 , \9728 , \9735 );
or \U$9369 ( \9746 , \9744 , \9745 );
and \U$9370 ( \9747 , \8371 , RIae76898_51);
and \U$9371 ( \9748 , RIae76b68_57, \8369 );
nor \U$9372 ( \9749 , \9747 , \9748 );
and \U$9373 ( \9750 , \9749 , \8020 );
not \U$9374 ( \9751 , \9749 );
and \U$9375 ( \9752 , \9751 , \8019 );
nor \U$9376 ( \9753 , \9750 , \9752 );
and \U$9377 ( \9754 , RIae7a510_180, RIae7a588_181);
not \U$9378 ( \9755 , RIae7a498_179);
and \U$9379 ( \9756 , \9755 , RIae7a588_181);
nor \U$9380 ( \9757 , \9755 , RIae7a588_181);
or \U$9381 ( \9758 , \9756 , \9757 );
nor \U$9382 ( \9759 , RIae7a510_180, RIae7a588_181);
nor \U$9383 ( \9760 , \9754 , \9758 , \9759 );
nand \U$9384 ( \9761 , RIae78da0_130, \9760 );
and \U$9385 ( \9762 , \9761 , \9273 );
not \U$9386 ( \9763 , \9761 );
buf \U$9387 ( \9764 , \9272 );
and \U$9388 ( \9765 , \9763 , \9764 );
nor \U$9389 ( \9766 , \9762 , \9765 );
xor \U$9390 ( \9767 , \9753 , \9766 );
and \U$9391 ( \9768 , \8966 , RIae78a58_123);
and \U$9392 ( \9769 , RIae78cb0_128, \8964 );
nor \U$9393 ( \9770 , \9768 , \9769 );
and \U$9394 ( \9771 , \9770 , \8799 );
not \U$9395 ( \9772 , \9770 );
and \U$9396 ( \9773 , \9772 , \8789 );
nor \U$9397 ( \9774 , \9771 , \9773 );
and \U$9398 ( \9775 , \9767 , \9774 );
and \U$9399 ( \9776 , \9753 , \9766 );
or \U$9400 ( \9777 , \9775 , \9776 );
xor \U$9401 ( \9778 , \9746 , \9777 );
and \U$9402 ( \9779 , \6941 , RIae76208_37);
and \U$9403 ( \9780 , RIae76a78_55, \6939 );
nor \U$9404 ( \9781 , \9779 , \9780 );
and \U$9405 ( \9782 , \9781 , \6314 );
not \U$9406 ( \9783 , \9781 );
and \U$9407 ( \9784 , \9783 , \6945 );
nor \U$9408 ( \9785 , \9782 , \9784 );
and \U$9409 ( \9786 , \6172 , RIae76028_33);
and \U$9410 ( \9787 , RIae762f8_39, \6170 );
nor \U$9411 ( \9788 , \9786 , \9787 );
and \U$9412 ( \9789 , \9788 , \6176 );
not \U$9413 ( \9790 , \9788 );
and \U$9414 ( \9791 , \9790 , \6175 );
nor \U$9415 ( \9792 , \9789 , \9791 );
xor \U$9416 ( \9793 , \9785 , \9792 );
and \U$9417 ( \9794 , \7633 , RIae76988_53);
and \U$9418 ( \9795 , RIae767a8_49, \7631 );
nor \U$9419 ( \9796 , \9794 , \9795 );
and \U$9420 ( \9797 , \9796 , \7206 );
not \U$9421 ( \9798 , \9796 );
and \U$9422 ( \9799 , \9798 , \7205 );
nor \U$9423 ( \9800 , \9797 , \9799 );
and \U$9424 ( \9801 , \9793 , \9800 );
and \U$9425 ( \9802 , \9785 , \9792 );
or \U$9426 ( \9803 , \9801 , \9802 );
and \U$9427 ( \9804 , \9778 , \9803 );
and \U$9428 ( \9805 , \9746 , \9777 );
or \U$9429 ( \9806 , \9804 , \9805 );
not \U$9430 ( \9807 , \400 );
and \U$9431 ( \9808 , \436 , RIae780f8_103);
and \U$9432 ( \9809 , RIae77f18_99, \434 );
nor \U$9433 ( \9810 , \9808 , \9809 );
not \U$9434 ( \9811 , \9810 );
or \U$9435 ( \9812 , \9807 , \9811 );
or \U$9436 ( \9813 , \9810 , \402 );
nand \U$9437 ( \9814 , \9812 , \9813 );
not \U$9438 ( \9815 , \471 );
and \U$9439 ( \9816 , \514 , RIae78008_101);
and \U$9440 ( \9817 , RIae781e8_105, \512 );
nor \U$9441 ( \9818 , \9816 , \9817 );
not \U$9442 ( \9819 , \9818 );
or \U$9443 ( \9820 , \9815 , \9819 );
or \U$9444 ( \9821 , \9818 , \469 );
nand \U$9445 ( \9822 , \9820 , \9821 );
xor \U$9446 ( \9823 , \9814 , \9822 );
and \U$9447 ( \9824 , \558 , RIae785a8_113);
and \U$9448 ( \9825 , RIae783c8_109, \556 );
nor \U$9449 ( \9826 , \9824 , \9825 );
and \U$9450 ( \9827 , \9826 , \504 );
not \U$9451 ( \9828 , \9826 );
and \U$9452 ( \9829 , \9828 , \562 );
nor \U$9453 ( \9830 , \9827 , \9829 );
and \U$9454 ( \9831 , \9823 , \9830 );
and \U$9455 ( \9832 , \9814 , \9822 );
or \U$9456 ( \9833 , \9831 , \9832 );
nand \U$9457 ( \9834 , RIae771f8_71, RIae78b48_125);
and \U$9458 ( \9835 , \384 , RIae772e8_73);
and \U$9459 ( \9836 , RIae782d8_107, \382 );
nor \U$9460 ( \9837 , \9835 , \9836 );
not \U$9461 ( \9838 , \9837 );
not \U$9462 ( \9839 , \392 );
and \U$9463 ( \9840 , \9838 , \9839 );
and \U$9464 ( \9841 , \9837 , \392 );
nor \U$9465 ( \9842 , \9840 , \9841 );
nand \U$9466 ( \9843 , \9834 , \9842 );
xor \U$9467 ( \9844 , \9833 , \9843 );
and \U$9468 ( \9845 , \1138 , RIae77e28_97);
and \U$9469 ( \9846 , RIae78968_121, \1136 );
nor \U$9470 ( \9847 , \9845 , \9846 );
and \U$9471 ( \9848 , \9847 , \1012 );
not \U$9472 ( \9849 , \9847 );
and \U$9473 ( \9850 , \9849 , \1142 );
nor \U$9474 ( \9851 , \9848 , \9850 );
and \U$9475 ( \9852 , \672 , RIae78530_112);
and \U$9476 ( \9853 , RIae77c48_93, \670 );
nor \U$9477 ( \9854 , \9852 , \9853 );
and \U$9478 ( \9855 , \9854 , \588 );
not \U$9479 ( \9856 , \9854 );
and \U$9480 ( \9857 , \9856 , \587 );
nor \U$9481 ( \9858 , \9855 , \9857 );
xor \U$9482 ( \9859 , \9851 , \9858 );
not \U$9483 ( \9860 , \789 );
and \U$9484 ( \9861 , \883 , RIae77b58_91);
and \U$9485 ( \9862 , RIae77d38_95, \881 );
nor \U$9486 ( \9863 , \9861 , \9862 );
not \U$9487 ( \9864 , \9863 );
or \U$9488 ( \9865 , \9860 , \9864 );
or \U$9489 ( \9866 , \9863 , \787 );
nand \U$9490 ( \9867 , \9865 , \9866 );
and \U$9491 ( \9868 , \9859 , \9867 );
and \U$9492 ( \9869 , \9851 , \9858 );
or \U$9493 ( \9870 , \9868 , \9869 );
and \U$9494 ( \9871 , \9844 , \9870 );
and \U$9495 ( \9872 , \9833 , \9843 );
or \U$9496 ( \9873 , \9871 , \9872 );
xor \U$9497 ( \9874 , \9806 , \9873 );
not \U$9498 ( \9875 , \2774 );
and \U$9499 ( \9876 , \3214 , RIae754e8_9);
and \U$9500 ( \9877 , RIae757b8_15, \3212 );
nor \U$9501 ( \9878 , \9876 , \9877 );
not \U$9502 ( \9879 , \9878 );
or \U$9503 ( \9880 , \9875 , \9879 );
or \U$9504 ( \9881 , \9878 , \3218 );
nand \U$9505 ( \9882 , \9880 , \9881 );
and \U$9506 ( \9883 , \3730 , RIae756c8_13);
and \U$9507 ( \9884 , RIae75218_3, \3728 );
nor \U$9508 ( \9885 , \9883 , \9884 );
and \U$9509 ( \9886 , \9885 , \3732 );
not \U$9510 ( \9887 , \9885 );
and \U$9511 ( \9888 , \9887 , \3421 );
nor \U$9512 ( \9889 , \9886 , \9888 );
xor \U$9513 ( \9890 , \9882 , \9889 );
and \U$9514 ( \9891 , \4247 , RIae75128_1);
and \U$9515 ( \9892 , RIae75308_5, \4245 );
nor \U$9516 ( \9893 , \9891 , \9892 );
and \U$9517 ( \9894 , \9893 , \3989 );
not \U$9518 ( \9895 , \9893 );
and \U$9519 ( \9896 , \9895 , \4251 );
nor \U$9520 ( \9897 , \9894 , \9896 );
and \U$9521 ( \9898 , \9890 , \9897 );
and \U$9522 ( \9899 , \9882 , \9889 );
or \U$9523 ( \9900 , \9898 , \9899 );
and \U$9524 ( \9901 , \1376 , RIae78878_119);
and \U$9525 ( \9902 , RIae78788_117, \1374 );
nor \U$9526 ( \9903 , \9901 , \9902 );
and \U$9527 ( \9904 , \9903 , \1380 );
not \U$9528 ( \9905 , \9903 );
and \U$9529 ( \9906 , \9905 , \1261 );
nor \U$9530 ( \9907 , \9904 , \9906 );
and \U$9531 ( \9908 , \1593 , RIae78698_115);
and \U$9532 ( \9909 , RIae75b78_23, \1591 );
nor \U$9533 ( \9910 , \9908 , \9909 );
and \U$9534 ( \9911 , \9910 , \1498 );
not \U$9535 ( \9912 , \9910 );
and \U$9536 ( \9913 , \9912 , \1488 );
nor \U$9537 ( \9914 , \9911 , \9913 );
xor \U$9538 ( \9915 , \9907 , \9914 );
and \U$9539 ( \9916 , \1939 , RIae75a88_21);
and \U$9540 ( \9917 , RIae75998_19, \1937 );
nor \U$9541 ( \9918 , \9916 , \9917 );
and \U$9542 ( \9919 , \9918 , \1735 );
not \U$9543 ( \9920 , \9918 );
and \U$9544 ( \9921 , \9920 , \1734 );
nor \U$9545 ( \9922 , \9919 , \9921 );
and \U$9546 ( \9923 , \9915 , \9922 );
and \U$9547 ( \9924 , \9907 , \9914 );
or \U$9548 ( \9925 , \9923 , \9924 );
xor \U$9549 ( \9926 , \9900 , \9925 );
not \U$9550 ( \9927 , \2789 );
and \U$9551 ( \9928 , \2783 , RIae75d58_27);
and \U$9552 ( \9929 , RIae755d8_11, \2781 );
nor \U$9553 ( \9930 , \9928 , \9929 );
not \U$9554 ( \9931 , \9930 );
or \U$9555 ( \9932 , \9927 , \9931 );
or \U$9556 ( \9933 , \9930 , \2789 );
nand \U$9557 ( \9934 , \9932 , \9933 );
and \U$9558 ( \9935 , \2224 , RIae758a8_17);
and \U$9559 ( \9936 , RIae75f38_31, \2222 );
nor \U$9560 ( \9937 , \9935 , \9936 );
and \U$9561 ( \9938 , \9937 , \2061 );
not \U$9562 ( \9939 , \9937 );
and \U$9563 ( \9940 , \9939 , \2060 );
nor \U$9564 ( \9941 , \9938 , \9940 );
xor \U$9565 ( \9942 , \9934 , \9941 );
and \U$9566 ( \9943 , \2607 , RIae75e48_29);
and \U$9567 ( \9944 , RIae75c68_25, \2605 );
nor \U$9568 ( \9945 , \9943 , \9944 );
and \U$9569 ( \9946 , \9945 , \2611 );
not \U$9570 ( \9947 , \9945 );
and \U$9571 ( \9948 , \9947 , \2397 );
nor \U$9572 ( \9949 , \9946 , \9948 );
and \U$9573 ( \9950 , \9942 , \9949 );
and \U$9574 ( \9951 , \9934 , \9941 );
or \U$9575 ( \9952 , \9950 , \9951 );
and \U$9576 ( \9953 , \9926 , \9952 );
and \U$9577 ( \9954 , \9900 , \9925 );
or \U$9578 ( \9955 , \9953 , \9954 );
and \U$9579 ( \9956 , \9874 , \9955 );
and \U$9580 ( \9957 , \9806 , \9873 );
or \U$9581 ( \9958 , \9956 , \9957 );
xor \U$9582 ( \9959 , \9721 , \9958 );
xor \U$9583 ( \9960 , \9104 , \9111 );
xor \U$9584 ( \9961 , \9960 , \9119 );
xor \U$9585 ( \9962 , \9225 , \9230 );
xor \U$9586 ( \9963 , \9961 , \9962 );
xor \U$9587 ( \9964 , \9216 , \9038 );
xor \U$9588 ( \9965 , \9964 , \9219 );
and \U$9589 ( \9966 , \9963 , \9965 );
xor \U$9590 ( \9967 , \8958 , \8971 );
xor \U$9591 ( \9968 , \9967 , \8979 );
xor \U$9592 ( \9969 , \9204 , \9209 );
xor \U$9593 ( \9970 , \9968 , \9969 );
xor \U$9594 ( \9971 , \9216 , \9038 );
xor \U$9595 ( \9972 , \9971 , \9219 );
and \U$9596 ( \9973 , \9970 , \9972 );
and \U$9597 ( \9974 , \9963 , \9970 );
or \U$9598 ( \9975 , \9966 , \9973 , \9974 );
and \U$9599 ( \9976 , \9959 , \9975 );
and \U$9600 ( \9977 , \9721 , \9958 );
or \U$9601 ( \9978 , \9976 , \9977 );
xor \U$9602 ( \9979 , \9313 , \9381 );
xor \U$9603 ( \9980 , \9979 , \9463 );
xor \U$9604 ( \9981 , \9214 , \9222 );
xor \U$9605 ( \9982 , \9981 , \9235 );
and \U$9606 ( \9983 , \9980 , \9982 );
xor \U$9607 ( \9984 , \9978 , \9983 );
xor \U$9608 ( \9985 , \9263 , \9284 );
xor \U$9609 ( \9986 , \9985 , \9310 );
xor \U$9610 ( \9987 , \9408 , \9433 );
xor \U$9611 ( \9988 , \9987 , \9460 );
xor \U$9612 ( \9989 , \9986 , \9988 );
xor \U$9613 ( \9990 , \9339 , \9350 );
xor \U$9614 ( \9991 , \9990 , \9378 );
and \U$9615 ( \9992 , \9989 , \9991 );
and \U$9616 ( \9993 , \9986 , \9988 );
or \U$9617 ( \9994 , \9992 , \9993 );
xor \U$9618 ( \9995 , \9485 , \9487 );
xor \U$9619 ( \9996 , \9995 , \9490 );
and \U$9620 ( \9997 , \9994 , \9996 );
xor \U$9621 ( \9998 , \9192 , \9194 );
xor \U$9622 ( \9999 , \9998 , \9197 );
xor \U$9623 ( \10000 , \9469 , \9474 );
xor \U$9624 ( \10001 , \9999 , \10000 );
xor \U$9625 ( \10002 , \9485 , \9487 );
xor \U$9626 ( \10003 , \10002 , \9490 );
and \U$9627 ( \10004 , \10001 , \10003 );
and \U$9628 ( \10005 , \9994 , \10001 );
or \U$9629 ( \10006 , \9997 , \10004 , \10005 );
and \U$9630 ( \10007 , \9984 , \10006 );
and \U$9631 ( \10008 , \9978 , \9983 );
or \U$9632 ( \10009 , \10007 , \10008 );
and \U$9633 ( \10010 , \9684 , \10009 );
not \U$9634 ( \10011 , \9684 );
not \U$9635 ( \10012 , \10009 );
and \U$9636 ( \10013 , \10011 , \10012 );
xnor \U$9637 ( \10014 , \9563 , \9580 );
not \U$9638 ( \10015 , \10014 );
not \U$9639 ( \10016 , \9548 );
and \U$9640 ( \10017 , \10015 , \10016 );
and \U$9641 ( \10018 , \10014 , \9548 );
nor \U$9642 ( \10019 , \10017 , \10018 );
nor \U$9643 ( \10020 , \10013 , \10019 );
nor \U$9644 ( \10021 , \10010 , \10020 );
xnor \U$9645 ( \10022 , \9617 , \9624 );
not \U$9646 ( \10023 , \10022 );
not \U$9647 ( \10024 , \9612 );
and \U$9648 ( \10025 , \10023 , \10024 );
and \U$9649 ( \10026 , \10022 , \9612 );
nor \U$9650 ( \10027 , \10025 , \10026 );
xor \U$9651 ( \10028 , \10021 , \10027 );
not \U$9652 ( \10029 , \9582 );
not \U$9653 ( \10030 , \9531 );
or \U$9654 ( \10031 , \10029 , \10030 );
or \U$9655 ( \10032 , \9531 , \9582 );
nand \U$9656 ( \10033 , \10031 , \10032 );
not \U$9657 ( \10034 , \10033 );
not \U$9658 ( \10035 , \8926 );
and \U$9659 ( \10036 , \10034 , \10035 );
and \U$9660 ( \10037 , \10033 , \8926 );
nor \U$9661 ( \10038 , \10036 , \10037 );
and \U$9662 ( \10039 , \10028 , \10038 );
and \U$9663 ( \10040 , \10021 , \10027 );
or \U$9664 ( \10041 , \10039 , \10040 );
nor \U$9665 ( \10042 , \9671 , \10041 );
and \U$9666 ( \10043 , \9668 , \10042 );
xor \U$9667 ( \10044 , \10042 , \9668 );
or \U$9668 ( \10045 , \9842 , \9834 );
nand \U$9669 ( \10046 , \10045 , \9843 );
xor \U$9670 ( \10047 , \9814 , \9822 );
xor \U$9671 ( \10048 , \10047 , \9830 );
and \U$9672 ( \10049 , \10046 , \10048 );
xor \U$9673 ( \10050 , \9851 , \9858 );
xor \U$9674 ( \10051 , \10050 , \9867 );
xor \U$9675 ( \10052 , \9814 , \9822 );
xor \U$9676 ( \10053 , \10052 , \9830 );
and \U$9677 ( \10054 , \10051 , \10053 );
and \U$9678 ( \10055 , \10046 , \10051 );
or \U$9679 ( \10056 , \10049 , \10054 , \10055 );
xor \U$9680 ( \10057 , \9753 , \9766 );
xor \U$9681 ( \10058 , \10057 , \9774 );
xor \U$9682 ( \10059 , \9785 , \9792 );
xor \U$9683 ( \10060 , \10059 , \9800 );
and \U$9684 ( \10061 , \10058 , \10060 );
xor \U$9685 ( \10062 , \9728 , \9735 );
xor \U$9686 ( \10063 , \10062 , \9743 );
xor \U$9687 ( \10064 , \9785 , \9792 );
xor \U$9688 ( \10065 , \10064 , \9800 );
and \U$9689 ( \10066 , \10063 , \10065 );
and \U$9690 ( \10067 , \10058 , \10063 );
or \U$9691 ( \10068 , \10061 , \10066 , \10067 );
xor \U$9692 ( \10069 , \10056 , \10068 );
xor \U$9693 ( \10070 , \9934 , \9941 );
xor \U$9694 ( \10071 , \10070 , \9949 );
xor \U$9695 ( \10072 , \9907 , \9914 );
xor \U$9696 ( \10073 , \10072 , \9922 );
xor \U$9697 ( \10074 , \10071 , \10073 );
xor \U$9698 ( \10075 , \9882 , \9889 );
xor \U$9699 ( \10076 , \10075 , \9897 );
and \U$9700 ( \10077 , \10074 , \10076 );
and \U$9701 ( \10078 , \10071 , \10073 );
or \U$9702 ( \10079 , \10077 , \10078 );
and \U$9703 ( \10080 , \10069 , \10079 );
and \U$9704 ( \10081 , \10056 , \10068 );
or \U$9705 ( \10082 , \10080 , \10081 );
and \U$9706 ( \10083 , \5399 , RIae763e8_41);
and \U$9707 ( \10084 , RIae764d8_43, \5397 );
nor \U$9708 ( \10085 , \10083 , \10084 );
and \U$9709 ( \10086 , \10085 , \5403 );
not \U$9710 ( \10087 , \10085 );
and \U$9711 ( \10088 , \10087 , \5016 );
nor \U$9712 ( \10089 , \10086 , \10088 );
and \U$9713 ( \10090 , \5896 , RIae766b8_47);
and \U$9714 ( \10091 , RIae765c8_45, \5894 );
nor \U$9715 ( \10092 , \10090 , \10091 );
and \U$9716 ( \10093 , \10092 , \5589 );
not \U$9717 ( \10094 , \10092 );
and \U$9718 ( \10095 , \10094 , \5590 );
nor \U$9719 ( \10096 , \10093 , \10095 );
or \U$9720 ( \10097 , \10089 , \10096 );
not \U$9721 ( \10098 , \10096 );
not \U$9722 ( \10099 , \10089 );
or \U$9723 ( \10100 , \10098 , \10099 );
and \U$9724 ( \10101 , \6172 , RIae76118_35);
and \U$9725 ( \10102 , RIae76028_33, \6170 );
nor \U$9726 ( \10103 , \10101 , \10102 );
and \U$9727 ( \10104 , \10103 , \6176 );
not \U$9728 ( \10105 , \10103 );
and \U$9729 ( \10106 , \10105 , \6175 );
nor \U$9730 ( \10107 , \10104 , \10106 );
nand \U$9731 ( \10108 , \10100 , \10107 );
nand \U$9732 ( \10109 , \10097 , \10108 );
and \U$9733 ( \10110 , \9760 , RIae78cb0_128);
and \U$9734 ( \10111 , RIae78da0_130, \9758 );
nor \U$9735 ( \10112 , \10110 , \10111 );
and \U$9736 ( \10113 , \10112 , \9272 );
not \U$9737 ( \10114 , \10112 );
and \U$9738 ( \10115 , \10114 , \9273 );
nor \U$9739 ( \10116 , \10113 , \10115 );
nand \U$9740 ( \10117 , RIae7a150_172, RIae7a420_178);
and \U$9741 ( \10118 , \10117 , RIae7a498_179);
or \U$9742 ( \10119 , \10116 , \10118 );
and \U$9743 ( \10120 , \10116 , \10118 );
and \U$9744 ( \10121 , \8966 , RIae76b68_57);
and \U$9745 ( \10122 , RIae78a58_123, \8964 );
nor \U$9746 ( \10123 , \10121 , \10122 );
and \U$9747 ( \10124 , \10123 , \8789 );
not \U$9748 ( \10125 , \10123 );
and \U$9749 ( \10126 , \10125 , \8799 );
nor \U$9750 ( \10127 , \10124 , \10126 );
nor \U$9751 ( \10128 , \10120 , \10127 );
not \U$9752 ( \10129 , \10128 );
nand \U$9753 ( \10130 , \10119 , \10129 );
xor \U$9754 ( \10131 , \10109 , \10130 );
and \U$9755 ( \10132 , \7633 , RIae76a78_55);
and \U$9756 ( \10133 , RIae76988_53, \7631 );
nor \U$9757 ( \10134 , \10132 , \10133 );
and \U$9758 ( \10135 , \10134 , \7206 );
not \U$9759 ( \10136 , \10134 );
and \U$9760 ( \10137 , \10136 , \7205 );
nor \U$9761 ( \10138 , \10135 , \10137 );
and \U$9762 ( \10139 , \6941 , RIae762f8_39);
and \U$9763 ( \10140 , RIae76208_37, \6939 );
nor \U$9764 ( \10141 , \10139 , \10140 );
and \U$9765 ( \10142 , \10141 , \6314 );
not \U$9766 ( \10143 , \10141 );
and \U$9767 ( \10144 , \10143 , \6945 );
nor \U$9768 ( \10145 , \10142 , \10144 );
xor \U$9769 ( \10146 , \10138 , \10145 );
and \U$9770 ( \10147 , \8371 , RIae767a8_49);
and \U$9771 ( \10148 , RIae76898_51, \8369 );
nor \U$9772 ( \10149 , \10147 , \10148 );
and \U$9773 ( \10150 , \10149 , \8020 );
not \U$9774 ( \10151 , \10149 );
and \U$9775 ( \10152 , \10151 , \8019 );
nor \U$9776 ( \10153 , \10150 , \10152 );
and \U$9777 ( \10154 , \10146 , \10153 );
and \U$9778 ( \10155 , \10138 , \10145 );
or \U$9779 ( \10156 , \10154 , \10155 );
and \U$9780 ( \10157 , \10131 , \10156 );
and \U$9781 ( \10158 , \10109 , \10130 );
or \U$9782 ( \10159 , \10157 , \10158 );
and \U$9783 ( \10160 , \384 , RIae771f8_71);
and \U$9784 ( \10161 , RIae772e8_73, \382 );
nor \U$9785 ( \10162 , \10160 , \10161 );
not \U$9786 ( \10163 , \10162 );
not \U$9787 ( \10164 , \392 );
and \U$9788 ( \10165 , \10163 , \10164 );
and \U$9789 ( \10166 , \10162 , \388 );
nor \U$9790 ( \10167 , \10165 , \10166 );
nand \U$9791 ( \10168 , RIae77018_67, RIae78b48_125);
xor \U$9792 ( \10169 , \10167 , \10168 );
and \U$9793 ( \10170 , \436 , RIae782d8_107);
and \U$9794 ( \10171 , RIae780f8_103, \434 );
nor \U$9795 ( \10172 , \10170 , \10171 );
not \U$9796 ( \10173 , \10172 );
not \U$9797 ( \10174 , \402 );
and \U$9798 ( \10175 , \10173 , \10174 );
and \U$9799 ( \10176 , \10172 , \402 );
nor \U$9800 ( \10177 , \10175 , \10176 );
and \U$9801 ( \10178 , \10169 , \10177 );
and \U$9802 ( \10179 , \10167 , \10168 );
or \U$9803 ( \10180 , \10178 , \10179 );
and \U$9804 ( \10181 , \1376 , RIae78968_121);
and \U$9805 ( \10182 , RIae78878_119, \1374 );
nor \U$9806 ( \10183 , \10181 , \10182 );
and \U$9807 ( \10184 , \10183 , \1261 );
not \U$9808 ( \10185 , \10183 );
and \U$9809 ( \10186 , \10185 , \1380 );
nor \U$9810 ( \10187 , \10184 , \10186 );
and \U$9811 ( \10188 , \883 , RIae77c48_93);
and \U$9812 ( \10189 , RIae77b58_91, \881 );
nor \U$9813 ( \10190 , \10188 , \10189 );
not \U$9814 ( \10191 , \10190 );
not \U$9815 ( \10192 , \787 );
and \U$9816 ( \10193 , \10191 , \10192 );
and \U$9817 ( \10194 , \10190 , \789 );
nor \U$9818 ( \10195 , \10193 , \10194 );
xor \U$9819 ( \10196 , \10187 , \10195 );
and \U$9820 ( \10197 , \1138 , RIae77d38_95);
and \U$9821 ( \10198 , RIae77e28_97, \1136 );
nor \U$9822 ( \10199 , \10197 , \10198 );
and \U$9823 ( \10200 , \10199 , \1142 );
not \U$9824 ( \10201 , \10199 );
and \U$9825 ( \10202 , \10201 , \1012 );
nor \U$9826 ( \10203 , \10200 , \10202 );
and \U$9827 ( \10204 , \10196 , \10203 );
and \U$9828 ( \10205 , \10187 , \10195 );
or \U$9829 ( \10206 , \10204 , \10205 );
xor \U$9830 ( \10207 , \10180 , \10206 );
and \U$9831 ( \10208 , \514 , RIae77f18_99);
and \U$9832 ( \10209 , RIae78008_101, \512 );
nor \U$9833 ( \10210 , \10208 , \10209 );
not \U$9834 ( \10211 , \10210 );
not \U$9835 ( \10212 , \471 );
and \U$9836 ( \10213 , \10211 , \10212 );
and \U$9837 ( \10214 , \10210 , \471 );
nor \U$9838 ( \10215 , \10213 , \10214 );
and \U$9839 ( \10216 , \558 , RIae781e8_105);
and \U$9840 ( \10217 , RIae785a8_113, \556 );
nor \U$9841 ( \10218 , \10216 , \10217 );
and \U$9842 ( \10219 , \10218 , \562 );
not \U$9843 ( \10220 , \10218 );
and \U$9844 ( \10221 , \10220 , \504 );
nor \U$9845 ( \10222 , \10219 , \10221 );
xor \U$9846 ( \10223 , \10215 , \10222 );
and \U$9847 ( \10224 , \672 , RIae783c8_109);
and \U$9848 ( \10225 , RIae78530_112, \670 );
nor \U$9849 ( \10226 , \10224 , \10225 );
and \U$9850 ( \10227 , \10226 , \587 );
not \U$9851 ( \10228 , \10226 );
and \U$9852 ( \10229 , \10228 , \588 );
nor \U$9853 ( \10230 , \10227 , \10229 );
and \U$9854 ( \10231 , \10223 , \10230 );
and \U$9855 ( \10232 , \10215 , \10222 );
or \U$9856 ( \10233 , \10231 , \10232 );
and \U$9857 ( \10234 , \10207 , \10233 );
and \U$9858 ( \10235 , \10180 , \10206 );
nor \U$9859 ( \10236 , \10234 , \10235 );
xor \U$9860 ( \10237 , \10159 , \10236 );
and \U$9861 ( \10238 , \2607 , RIae75f38_31);
and \U$9862 ( \10239 , RIae75e48_29, \2605 );
nor \U$9863 ( \10240 , \10238 , \10239 );
and \U$9864 ( \10241 , \10240 , \2397 );
not \U$9865 ( \10242 , \10240 );
and \U$9866 ( \10243 , \10242 , \2611 );
nor \U$9867 ( \10244 , \10241 , \10243 );
not \U$9868 ( \10245 , \10244 );
and \U$9869 ( \10246 , \2783 , RIae75c68_25);
and \U$9870 ( \10247 , RIae75d58_27, \2781 );
nor \U$9871 ( \10248 , \10246 , \10247 );
not \U$9872 ( \10249 , \10248 );
not \U$9873 ( \10250 , \3089 );
and \U$9874 ( \10251 , \10249 , \10250 );
and \U$9875 ( \10252 , \10248 , \2789 );
nor \U$9876 ( \10253 , \10251 , \10252 );
not \U$9877 ( \10254 , \10253 );
and \U$9878 ( \10255 , \10245 , \10254 );
and \U$9879 ( \10256 , \10253 , \10244 );
and \U$9880 ( \10257 , \3214 , RIae755d8_11);
and \U$9881 ( \10258 , RIae754e8_9, \3212 );
nor \U$9882 ( \10259 , \10257 , \10258 );
not \U$9883 ( \10260 , \10259 );
not \U$9884 ( \10261 , \3218 );
and \U$9885 ( \10262 , \10260 , \10261 );
and \U$9886 ( \10263 , \10259 , \2774 );
nor \U$9887 ( \10264 , \10262 , \10263 );
nor \U$9888 ( \10265 , \10256 , \10264 );
nor \U$9889 ( \10266 , \10255 , \10265 );
and \U$9890 ( \10267 , \3730 , RIae757b8_15);
and \U$9891 ( \10268 , RIae756c8_13, \3728 );
nor \U$9892 ( \10269 , \10267 , \10268 );
and \U$9893 ( \10270 , \10269 , \3422 );
not \U$9894 ( \10271 , \10269 );
and \U$9895 ( \10272 , \10271 , \3732 );
nor \U$9896 ( \10273 , \10270 , \10272 );
not \U$9897 ( \10274 , \10273 );
and \U$9898 ( \10275 , \4247 , RIae75218_3);
and \U$9899 ( \10276 , RIae75128_1, \4245 );
nor \U$9900 ( \10277 , \10275 , \10276 );
and \U$9901 ( \10278 , \10277 , \4251 );
not \U$9902 ( \10279 , \10277 );
and \U$9903 ( \10280 , \10279 , \3989 );
nor \U$9904 ( \10281 , \10278 , \10280 );
not \U$9905 ( \10282 , \10281 );
and \U$9906 ( \10283 , \10274 , \10282 );
and \U$9907 ( \10284 , \10281 , \10273 );
and \U$9908 ( \10285 , \4688 , RIae75308_5);
and \U$9909 ( \10286 , RIae753f8_7, \4686 );
nor \U$9910 ( \10287 , \10285 , \10286 );
and \U$9911 ( \10288 , \10287 , \4482 );
not \U$9912 ( \10289 , \10287 );
and \U$9913 ( \10290 , \10289 , \4481 );
nor \U$9914 ( \10291 , \10288 , \10290 );
nor \U$9915 ( \10292 , \10284 , \10291 );
nor \U$9916 ( \10293 , \10283 , \10292 );
xor \U$9917 ( \10294 , \10266 , \10293 );
and \U$9918 ( \10295 , \1593 , RIae78788_117);
and \U$9919 ( \10296 , RIae78698_115, \1591 );
nor \U$9920 ( \10297 , \10295 , \10296 );
and \U$9921 ( \10298 , \10297 , \1488 );
not \U$9922 ( \10299 , \10297 );
and \U$9923 ( \10300 , \10299 , \1498 );
nor \U$9924 ( \10301 , \10298 , \10300 );
not \U$9925 ( \10302 , \10301 );
and \U$9926 ( \10303 , \1939 , RIae75b78_23);
and \U$9927 ( \10304 , RIae75a88_21, \1937 );
nor \U$9928 ( \10305 , \10303 , \10304 );
and \U$9929 ( \10306 , \10305 , \1734 );
not \U$9930 ( \10307 , \10305 );
and \U$9931 ( \10308 , \10307 , \1735 );
nor \U$9932 ( \10309 , \10306 , \10308 );
not \U$9933 ( \10310 , \10309 );
and \U$9934 ( \10311 , \10302 , \10310 );
and \U$9935 ( \10312 , \10309 , \10301 );
and \U$9936 ( \10313 , \2224 , RIae75998_19);
and \U$9937 ( \10314 , RIae758a8_17, \2222 );
nor \U$9938 ( \10315 , \10313 , \10314 );
and \U$9939 ( \10316 , \10315 , \2060 );
not \U$9940 ( \10317 , \10315 );
and \U$9941 ( \10318 , \10317 , \2061 );
nor \U$9942 ( \10319 , \10316 , \10318 );
nor \U$9943 ( \10320 , \10312 , \10319 );
nor \U$9944 ( \10321 , \10311 , \10320 );
and \U$9945 ( \10322 , \10294 , \10321 );
and \U$9946 ( \10323 , \10266 , \10293 );
nor \U$9947 ( \10324 , \10322 , \10323 );
and \U$9948 ( \10325 , \10237 , \10324 );
and \U$9949 ( \10326 , \10159 , \10236 );
or \U$9950 ( \10327 , \10325 , \10326 );
xor \U$9951 ( \10328 , \10082 , \10327 );
xor \U$9952 ( \10329 , \9270 , \9273 );
xor \U$9953 ( \10330 , \10329 , \9281 );
xor \U$9954 ( \10331 , \9686 , \9691 );
xor \U$9955 ( \10332 , \10330 , \10331 );
xor \U$9956 ( \10333 , \9698 , \9699 );
xor \U$9957 ( \10334 , \10333 , \9702 );
and \U$9958 ( \10335 , \10332 , \10334 );
xor \U$9959 ( \10336 , \9389 , \9396 );
xor \U$9960 ( \10337 , \10336 , \9405 );
xor \U$9961 ( \10338 , \9708 , \9713 );
xor \U$9962 ( \10339 , \10337 , \10338 );
xor \U$9963 ( \10340 , \9698 , \9699 );
xor \U$9964 ( \10341 , \10340 , \9702 );
and \U$9965 ( \10342 , \10339 , \10341 );
and \U$9966 ( \10343 , \10332 , \10339 );
or \U$9967 ( \10344 , \10335 , \10342 , \10343 );
and \U$9968 ( \10345 , \10328 , \10344 );
and \U$9969 ( \10346 , \10082 , \10327 );
or \U$9970 ( \10347 , \10345 , \10346 );
xor \U$9971 ( \10348 , \9806 , \9873 );
xor \U$9972 ( \10349 , \10348 , \9955 );
xor \U$9973 ( \10350 , \9696 , \9705 );
xor \U$9974 ( \10351 , \10350 , \9718 );
and \U$9975 ( \10352 , \10349 , \10351 );
xor \U$9976 ( \10353 , \10347 , \10352 );
xor \U$9977 ( \10354 , \9746 , \9777 );
xor \U$9978 ( \10355 , \10354 , \9803 );
xor \U$9979 ( \10356 , \9833 , \9843 );
xor \U$9980 ( \10357 , \10356 , \9870 );
xor \U$9981 ( \10358 , \10355 , \10357 );
xor \U$9982 ( \10359 , \9900 , \9925 );
xor \U$9983 ( \10360 , \10359 , \9952 );
and \U$9984 ( \10361 , \10358 , \10360 );
and \U$9985 ( \10362 , \10355 , \10357 );
or \U$9986 ( \10363 , \10361 , \10362 );
xor \U$9987 ( \10364 , \9986 , \9988 );
xor \U$9988 ( \10365 , \10364 , \9991 );
and \U$9989 ( \10366 , \10363 , \10365 );
xor \U$9990 ( \10367 , \9216 , \9038 );
xor \U$9991 ( \10368 , \10367 , \9219 );
xor \U$9992 ( \10369 , \9963 , \9970 );
xor \U$9993 ( \10370 , \10368 , \10369 );
xor \U$9994 ( \10371 , \9986 , \9988 );
xor \U$9995 ( \10372 , \10371 , \9991 );
and \U$9996 ( \10373 , \10370 , \10372 );
and \U$9997 ( \10374 , \10363 , \10370 );
or \U$9998 ( \10375 , \10366 , \10373 , \10374 );
and \U$9999 ( \10376 , \10353 , \10375 );
and \U$10000 ( \10377 , \10347 , \10352 );
or \U$10001 ( \10378 , \10376 , \10377 );
xor \U$10002 ( \10379 , \9980 , \9982 );
xor \U$10003 ( \10380 , \9721 , \9958 );
xor \U$10004 ( \10381 , \10380 , \9975 );
and \U$10005 ( \10382 , \10379 , \10381 );
xor \U$10006 ( \10383 , \9485 , \9487 );
xor \U$10007 ( \10384 , \10383 , \9490 );
xor \U$10008 ( \10385 , \9994 , \10001 );
xor \U$10009 ( \10386 , \10384 , \10385 );
xor \U$10010 ( \10387 , \9721 , \9958 );
xor \U$10011 ( \10388 , \10387 , \9975 );
and \U$10012 ( \10389 , \10386 , \10388 );
and \U$10013 ( \10390 , \10379 , \10386 );
or \U$10014 ( \10391 , \10382 , \10389 , \10390 );
xor \U$10015 ( \10392 , \10378 , \10391 );
xor \U$10016 ( \10393 , \9238 , \9466 );
xor \U$10017 ( \10394 , \10393 , \9479 );
xor \U$10018 ( \10395 , \9672 , \9679 );
xor \U$10019 ( \10396 , \10394 , \10395 );
and \U$10020 ( \10397 , \10392 , \10396 );
and \U$10021 ( \10398 , \10378 , \10391 );
or \U$10022 ( \10399 , \10397 , \10398 );
xor \U$10023 ( \10400 , \9202 , \9482 );
xor \U$10024 ( \10401 , \10400 , \9528 );
xor \U$10025 ( \10402 , \10399 , \10401 );
not \U$10026 ( \10403 , \10019 );
xor \U$10027 ( \10404 , \10009 , \9684 );
not \U$10028 ( \10405 , \10404 );
or \U$10029 ( \10406 , \10403 , \10405 );
or \U$10030 ( \10407 , \10404 , \10019 );
nand \U$10031 ( \10408 , \10406 , \10407 );
and \U$10032 ( \10409 , \10402 , \10408 );
and \U$10033 ( \10410 , \10399 , \10401 );
or \U$10034 ( \10411 , \10409 , \10410 );
not \U$10035 ( \10412 , \10411 );
xor \U$10036 ( \10413 , \10021 , \10027 );
xor \U$10037 ( \10414 , \10413 , \10038 );
not \U$10038 ( \10415 , \10414 );
or \U$10039 ( \10416 , \10412 , \10415 );
or \U$10040 ( \10417 , \10414 , \10411 );
nand \U$10041 ( \10418 , \10416 , \10417 );
and \U$10042 ( \10419 , \10116 , \10118 );
not \U$10043 ( \10420 , \10116 );
not \U$10044 ( \10421 , \10118 );
and \U$10045 ( \10422 , \10420 , \10421 );
nor \U$10046 ( \10423 , \10419 , \10422 );
not \U$10047 ( \10424 , \10423 );
not \U$10048 ( \10425 , \10127 );
and \U$10049 ( \10426 , \10424 , \10425 );
and \U$10050 ( \10427 , \10423 , \10127 );
nor \U$10051 ( \10428 , \10426 , \10427 );
not \U$10052 ( \10429 , \10096 );
not \U$10053 ( \10430 , \10107 );
or \U$10054 ( \10431 , \10429 , \10430 );
or \U$10055 ( \10432 , \10096 , \10107 );
nand \U$10056 ( \10433 , \10431 , \10432 );
not \U$10057 ( \10434 , \10433 );
not \U$10058 ( \10435 , \10089 );
and \U$10059 ( \10436 , \10434 , \10435 );
and \U$10060 ( \10437 , \10433 , \10089 );
nor \U$10061 ( \10438 , \10436 , \10437 );
or \U$10062 ( \10439 , \10428 , \10438 );
not \U$10063 ( \10440 , \10438 );
not \U$10064 ( \10441 , \10428 );
or \U$10065 ( \10442 , \10440 , \10441 );
xor \U$10066 ( \10443 , \10138 , \10145 );
xor \U$10067 ( \10444 , \10443 , \10153 );
nand \U$10068 ( \10445 , \10442 , \10444 );
nand \U$10069 ( \10446 , \10439 , \10445 );
xor \U$10070 ( \10447 , \10187 , \10195 );
xor \U$10071 ( \10448 , \10447 , \10203 );
xor \U$10072 ( \10449 , \10167 , \10168 );
xor \U$10073 ( \10450 , \10449 , \10177 );
xor \U$10074 ( \10451 , \10448 , \10450 );
xor \U$10075 ( \10452 , \10215 , \10222 );
xor \U$10076 ( \10453 , \10452 , \10230 );
and \U$10077 ( \10454 , \10451 , \10453 );
and \U$10078 ( \10455 , \10448 , \10450 );
nor \U$10079 ( \10456 , \10454 , \10455 );
xor \U$10080 ( \10457 , \10446 , \10456 );
not \U$10081 ( \10458 , \10244 );
xor \U$10082 ( \10459 , \10253 , \10264 );
not \U$10083 ( \10460 , \10459 );
or \U$10084 ( \10461 , \10458 , \10460 );
or \U$10085 ( \10462 , \10459 , \10244 );
nand \U$10086 ( \10463 , \10461 , \10462 );
not \U$10087 ( \10464 , \10301 );
xor \U$10088 ( \10465 , \10309 , \10319 );
not \U$10089 ( \10466 , \10465 );
or \U$10090 ( \10467 , \10464 , \10466 );
or \U$10091 ( \10468 , \10465 , \10301 );
nand \U$10092 ( \10469 , \10467 , \10468 );
xor \U$10093 ( \10470 , \10463 , \10469 );
not \U$10094 ( \10471 , \10273 );
xor \U$10095 ( \10472 , \10281 , \10291 );
not \U$10096 ( \10473 , \10472 );
or \U$10097 ( \10474 , \10471 , \10473 );
or \U$10098 ( \10475 , \10472 , \10273 );
nand \U$10099 ( \10476 , \10474 , \10475 );
and \U$10100 ( \10477 , \10470 , \10476 );
and \U$10101 ( \10478 , \10463 , \10469 );
or \U$10102 ( \10479 , \10477 , \10478 );
and \U$10103 ( \10480 , \10457 , \10479 );
and \U$10104 ( \10481 , \10446 , \10456 );
or \U$10105 ( \10482 , \10480 , \10481 );
and \U$10106 ( \10483 , \6941 , RIae76028_33);
and \U$10107 ( \10484 , RIae762f8_39, \6939 );
nor \U$10108 ( \10485 , \10483 , \10484 );
and \U$10109 ( \10486 , \10485 , \6314 );
not \U$10110 ( \10487 , \10485 );
and \U$10111 ( \10488 , \10487 , \6945 );
nor \U$10112 ( \10489 , \10486 , \10488 );
and \U$10113 ( \10490 , \7633 , RIae76208_37);
and \U$10114 ( \10491 , RIae76a78_55, \7631 );
nor \U$10115 ( \10492 , \10490 , \10491 );
and \U$10116 ( \10493 , \10492 , \7206 );
not \U$10117 ( \10494 , \10492 );
and \U$10118 ( \10495 , \10494 , \7205 );
nor \U$10119 ( \10496 , \10493 , \10495 );
xor \U$10120 ( \10497 , \10489 , \10496 );
and \U$10121 ( \10498 , \8371 , RIae76988_53);
and \U$10122 ( \10499 , RIae767a8_49, \8369 );
nor \U$10123 ( \10500 , \10498 , \10499 );
and \U$10124 ( \10501 , \10500 , \8020 );
not \U$10125 ( \10502 , \10500 );
and \U$10126 ( \10503 , \10502 , \8019 );
nor \U$10127 ( \10504 , \10501 , \10503 );
and \U$10128 ( \10505 , \10497 , \10504 );
and \U$10129 ( \10506 , \10489 , \10496 );
or \U$10130 ( \10507 , \10505 , \10506 );
and \U$10131 ( \10508 , \5399 , RIae753f8_7);
and \U$10132 ( \10509 , RIae763e8_41, \5397 );
nor \U$10133 ( \10510 , \10508 , \10509 );
and \U$10134 ( \10511 , \10510 , \5016 );
not \U$10135 ( \10512 , \10510 );
and \U$10136 ( \10513 , \10512 , \5403 );
nor \U$10137 ( \10514 , \10511 , \10513 );
and \U$10138 ( \10515 , \5896 , RIae764d8_43);
and \U$10139 ( \10516 , RIae766b8_47, \5894 );
nor \U$10140 ( \10517 , \10515 , \10516 );
and \U$10141 ( \10518 , \10517 , \5590 );
not \U$10142 ( \10519 , \10517 );
and \U$10143 ( \10520 , \10519 , \5589 );
nor \U$10144 ( \10521 , \10518 , \10520 );
xor \U$10145 ( \10522 , \10514 , \10521 );
and \U$10146 ( \10523 , \6172 , RIae765c8_45);
and \U$10147 ( \10524 , RIae76118_35, \6170 );
nor \U$10148 ( \10525 , \10523 , \10524 );
and \U$10149 ( \10526 , \10525 , \6176 );
not \U$10150 ( \10527 , \10525 );
and \U$10151 ( \10528 , \10527 , \6175 );
nor \U$10152 ( \10529 , \10526 , \10528 );
and \U$10153 ( \10530 , \10522 , \10529 );
and \U$10154 ( \10531 , \10514 , \10521 );
or \U$10155 ( \10532 , \10530 , \10531 );
xor \U$10156 ( \10533 , \10507 , \10532 );
and \U$10157 ( \10534 , \8966 , RIae76898_51);
and \U$10158 ( \10535 , RIae76b68_57, \8964 );
nor \U$10159 ( \10536 , \10534 , \10535 );
and \U$10160 ( \10537 , \10536 , \8799 );
not \U$10161 ( \10538 , \10536 );
and \U$10162 ( \10539 , \10538 , \8789 );
nor \U$10163 ( \10540 , \10537 , \10539 );
and \U$10164 ( \10541 , RIae7a498_179, RIae7a420_178);
not \U$10165 ( \10542 , RIae7a420_178);
nor \U$10166 ( \10543 , \10542 , RIae7a150_172);
not \U$10167 ( \10544 , RIae7a150_172);
nor \U$10168 ( \10545 , \10544 , RIae7a420_178);
or \U$10169 ( \10546 , \10543 , \10545 );
nor \U$10170 ( \10547 , RIae7a498_179, RIae7a420_178);
nor \U$10171 ( \10548 , \10541 , \10546 , \10547 );
nand \U$10172 ( \10549 , RIae78da0_130, \10548 );
and \U$10173 ( \10550 , \10549 , \10421 );
not \U$10174 ( \10551 , \10549 );
and \U$10175 ( \10552 , \10551 , \10118 );
nor \U$10176 ( \10553 , \10550 , \10552 );
xor \U$10177 ( \10554 , \10540 , \10553 );
and \U$10178 ( \10555 , \9760 , RIae78a58_123);
and \U$10179 ( \10556 , RIae78cb0_128, \9758 );
nor \U$10180 ( \10557 , \10555 , \10556 );
and \U$10181 ( \10558 , \10557 , \9273 );
not \U$10182 ( \10559 , \10557 );
and \U$10183 ( \10560 , \10559 , \9764 );
nor \U$10184 ( \10561 , \10558 , \10560 );
and \U$10185 ( \10562 , \10554 , \10561 );
and \U$10186 ( \10563 , \10540 , \10553 );
or \U$10187 ( \10564 , \10562 , \10563 );
and \U$10188 ( \10565 , \10533 , \10564 );
and \U$10189 ( \10566 , \10507 , \10532 );
or \U$10190 ( \10567 , \10565 , \10566 );
and \U$10191 ( \10568 , \1138 , RIae77b58_91);
and \U$10192 ( \10569 , RIae77d38_95, \1136 );
nor \U$10193 ( \10570 , \10568 , \10569 );
and \U$10194 ( \10571 , \10570 , \1012 );
not \U$10195 ( \10572 , \10570 );
and \U$10196 ( \10573 , \10572 , \1142 );
nor \U$10197 ( \10574 , \10571 , \10573 );
not \U$10198 ( \10575 , \789 );
and \U$10199 ( \10576 , \883 , RIae78530_112);
and \U$10200 ( \10577 , RIae77c48_93, \881 );
nor \U$10201 ( \10578 , \10576 , \10577 );
not \U$10202 ( \10579 , \10578 );
or \U$10203 ( \10580 , \10575 , \10579 );
or \U$10204 ( \10581 , \10578 , \787 );
nand \U$10205 ( \10582 , \10580 , \10581 );
xor \U$10206 ( \10583 , \10574 , \10582 );
and \U$10207 ( \10584 , \1376 , RIae77e28_97);
and \U$10208 ( \10585 , RIae78968_121, \1374 );
nor \U$10209 ( \10586 , \10584 , \10585 );
and \U$10210 ( \10587 , \10586 , \1380 );
not \U$10211 ( \10588 , \10586 );
and \U$10212 ( \10589 , \10588 , \1261 );
nor \U$10213 ( \10590 , \10587 , \10589 );
and \U$10214 ( \10591 , \10583 , \10590 );
and \U$10215 ( \10592 , \10574 , \10582 );
or \U$10216 ( \10593 , \10591 , \10592 );
and \U$10217 ( \10594 , \436 , RIae772e8_73);
and \U$10218 ( \10595 , RIae782d8_107, \434 );
nor \U$10219 ( \10596 , \10594 , \10595 );
not \U$10220 ( \10597 , \10596 );
not \U$10221 ( \10598 , \400 );
and \U$10222 ( \10599 , \10597 , \10598 );
and \U$10223 ( \10600 , \10596 , \400 );
nor \U$10224 ( \10601 , \10599 , \10600 );
nand \U$10225 ( \10602 , RIae77180_70, RIae78b48_125);
or \U$10226 ( \10603 , \10601 , \10602 );
not \U$10227 ( \10604 , \10602 );
not \U$10228 ( \10605 , \10601 );
or \U$10229 ( \10606 , \10604 , \10605 );
not \U$10230 ( \10607 , \388 );
and \U$10231 ( \10608 , \384 , RIae77018_67);
and \U$10232 ( \10609 , RIae771f8_71, \382 );
nor \U$10233 ( \10610 , \10608 , \10609 );
not \U$10234 ( \10611 , \10610 );
or \U$10235 ( \10612 , \10607 , \10611 );
or \U$10236 ( \10613 , \10610 , \392 );
nand \U$10237 ( \10614 , \10612 , \10613 );
nand \U$10238 ( \10615 , \10606 , \10614 );
nand \U$10239 ( \10616 , \10603 , \10615 );
xor \U$10240 ( \10617 , \10593 , \10616 );
and \U$10241 ( \10618 , \558 , RIae78008_101);
and \U$10242 ( \10619 , RIae781e8_105, \556 );
nor \U$10243 ( \10620 , \10618 , \10619 );
and \U$10244 ( \10621 , \10620 , \562 );
not \U$10245 ( \10622 , \10620 );
and \U$10246 ( \10623 , \10622 , \504 );
nor \U$10247 ( \10624 , \10621 , \10623 );
and \U$10248 ( \10625 , \672 , RIae785a8_113);
and \U$10249 ( \10626 , RIae783c8_109, \670 );
nor \U$10250 ( \10627 , \10625 , \10626 );
and \U$10251 ( \10628 , \10627 , \587 );
not \U$10252 ( \10629 , \10627 );
and \U$10253 ( \10630 , \10629 , \588 );
nor \U$10254 ( \10631 , \10628 , \10630 );
xor \U$10255 ( \10632 , \10624 , \10631 );
and \U$10256 ( \10633 , \514 , RIae780f8_103);
and \U$10257 ( \10634 , RIae77f18_99, \512 );
nor \U$10258 ( \10635 , \10633 , \10634 );
not \U$10259 ( \10636 , \10635 );
not \U$10260 ( \10637 , \471 );
and \U$10261 ( \10638 , \10636 , \10637 );
and \U$10262 ( \10639 , \10635 , \469 );
nor \U$10263 ( \10640 , \10638 , \10639 );
and \U$10264 ( \10641 , \10632 , \10640 );
and \U$10265 ( \10642 , \10624 , \10631 );
nor \U$10266 ( \10643 , \10641 , \10642 );
and \U$10267 ( \10644 , \10617 , \10643 );
and \U$10268 ( \10645 , \10593 , \10616 );
or \U$10269 ( \10646 , \10644 , \10645 );
xor \U$10270 ( \10647 , \10567 , \10646 );
and \U$10271 ( \10648 , \3730 , RIae754e8_9);
and \U$10272 ( \10649 , RIae757b8_15, \3728 );
nor \U$10273 ( \10650 , \10648 , \10649 );
and \U$10274 ( \10651 , \10650 , \3732 );
not \U$10275 ( \10652 , \10650 );
and \U$10276 ( \10653 , \10652 , \3422 );
nor \U$10277 ( \10654 , \10651 , \10653 );
and \U$10278 ( \10655 , \4247 , RIae756c8_13);
and \U$10279 ( \10656 , RIae75218_3, \4245 );
nor \U$10280 ( \10657 , \10655 , \10656 );
and \U$10281 ( \10658 , \10657 , \3989 );
not \U$10282 ( \10659 , \10657 );
and \U$10283 ( \10660 , \10659 , \4251 );
nor \U$10284 ( \10661 , \10658 , \10660 );
xor \U$10285 ( \10662 , \10654 , \10661 );
and \U$10286 ( \10663 , \4688 , RIae75128_1);
and \U$10287 ( \10664 , RIae75308_5, \4686 );
nor \U$10288 ( \10665 , \10663 , \10664 );
and \U$10289 ( \10666 , \10665 , \4481 );
not \U$10290 ( \10667 , \10665 );
and \U$10291 ( \10668 , \10667 , \4482 );
nor \U$10292 ( \10669 , \10666 , \10668 );
and \U$10293 ( \10670 , \10662 , \10669 );
and \U$10294 ( \10671 , \10654 , \10661 );
or \U$10295 ( \10672 , \10670 , \10671 );
and \U$10296 ( \10673 , \2607 , RIae758a8_17);
and \U$10297 ( \10674 , RIae75f38_31, \2605 );
nor \U$10298 ( \10675 , \10673 , \10674 );
and \U$10299 ( \10676 , \10675 , \2611 );
not \U$10300 ( \10677 , \10675 );
and \U$10301 ( \10678 , \10677 , \2397 );
nor \U$10302 ( \10679 , \10676 , \10678 );
not \U$10303 ( \10680 , \3089 );
and \U$10304 ( \10681 , \2783 , RIae75e48_29);
and \U$10305 ( \10682 , RIae75c68_25, \2781 );
nor \U$10306 ( \10683 , \10681 , \10682 );
not \U$10307 ( \10684 , \10683 );
or \U$10308 ( \10685 , \10680 , \10684 );
or \U$10309 ( \10686 , \10683 , \3089 );
nand \U$10310 ( \10687 , \10685 , \10686 );
xor \U$10311 ( \10688 , \10679 , \10687 );
not \U$10312 ( \10689 , \3218 );
and \U$10313 ( \10690 , \3214 , RIae75d58_27);
and \U$10314 ( \10691 , RIae755d8_11, \3212 );
nor \U$10315 ( \10692 , \10690 , \10691 );
not \U$10316 ( \10693 , \10692 );
or \U$10317 ( \10694 , \10689 , \10693 );
or \U$10318 ( \10695 , \10692 , \3218 );
nand \U$10319 ( \10696 , \10694 , \10695 );
and \U$10320 ( \10697 , \10688 , \10696 );
and \U$10321 ( \10698 , \10679 , \10687 );
or \U$10322 ( \10699 , \10697 , \10698 );
xor \U$10323 ( \10700 , \10672 , \10699 );
and \U$10324 ( \10701 , \1939 , RIae78698_115);
and \U$10325 ( \10702 , RIae75b78_23, \1937 );
nor \U$10326 ( \10703 , \10701 , \10702 );
and \U$10327 ( \10704 , \10703 , \1735 );
not \U$10328 ( \10705 , \10703 );
and \U$10329 ( \10706 , \10705 , \1734 );
nor \U$10330 ( \10707 , \10704 , \10706 );
and \U$10331 ( \10708 , \1593 , RIae78878_119);
and \U$10332 ( \10709 , RIae78788_117, \1591 );
nor \U$10333 ( \10710 , \10708 , \10709 );
and \U$10334 ( \10711 , \10710 , \1498 );
not \U$10335 ( \10712 , \10710 );
and \U$10336 ( \10713 , \10712 , \1488 );
nor \U$10337 ( \10714 , \10711 , \10713 );
xor \U$10338 ( \10715 , \10707 , \10714 );
and \U$10339 ( \10716 , \2224 , RIae75a88_21);
and \U$10340 ( \10717 , RIae75998_19, \2222 );
nor \U$10341 ( \10718 , \10716 , \10717 );
and \U$10342 ( \10719 , \10718 , \2061 );
not \U$10343 ( \10720 , \10718 );
and \U$10344 ( \10721 , \10720 , \2060 );
nor \U$10345 ( \10722 , \10719 , \10721 );
and \U$10346 ( \10723 , \10715 , \10722 );
and \U$10347 ( \10724 , \10707 , \10714 );
or \U$10348 ( \10725 , \10723 , \10724 );
and \U$10349 ( \10726 , \10700 , \10725 );
and \U$10350 ( \10727 , \10672 , \10699 );
or \U$10351 ( \10728 , \10726 , \10727 );
and \U$10352 ( \10729 , \10647 , \10728 );
and \U$10353 ( \10730 , \10567 , \10646 );
or \U$10354 ( \10731 , \10729 , \10730 );
xor \U$10355 ( \10732 , \10482 , \10731 );
xor \U$10356 ( \10733 , \9814 , \9822 );
xor \U$10357 ( \10734 , \10733 , \9830 );
xor \U$10358 ( \10735 , \10046 , \10051 );
xor \U$10359 ( \10736 , \10734 , \10735 );
xor \U$10360 ( \10737 , \10071 , \10073 );
xor \U$10361 ( \10738 , \10737 , \10076 );
and \U$10362 ( \10739 , \10736 , \10738 );
xor \U$10363 ( \10740 , \9785 , \9792 );
xor \U$10364 ( \10741 , \10740 , \9800 );
xor \U$10365 ( \10742 , \10058 , \10063 );
xor \U$10366 ( \10743 , \10741 , \10742 );
xor \U$10367 ( \10744 , \10071 , \10073 );
xor \U$10368 ( \10745 , \10744 , \10076 );
and \U$10369 ( \10746 , \10743 , \10745 );
and \U$10370 ( \10747 , \10736 , \10743 );
or \U$10371 ( \10748 , \10739 , \10746 , \10747 );
and \U$10372 ( \10749 , \10732 , \10748 );
and \U$10373 ( \10750 , \10482 , \10731 );
or \U$10374 ( \10751 , \10749 , \10750 );
xor \U$10375 ( \10752 , \10159 , \10236 );
xor \U$10376 ( \10753 , \10752 , \10324 );
xor \U$10377 ( \10754 , \10056 , \10068 );
xor \U$10378 ( \10755 , \10754 , \10079 );
and \U$10379 ( \10756 , \10753 , \10755 );
xor \U$10380 ( \10757 , \10751 , \10756 );
xor \U$10381 ( \10758 , \10180 , \10206 );
xor \U$10382 ( \10759 , \10758 , \10233 );
xor \U$10383 ( \10760 , \10266 , \10293 );
xor \U$10384 ( \10761 , \10760 , \10321 );
or \U$10385 ( \10762 , \10759 , \10761 );
not \U$10386 ( \10763 , \10761 );
not \U$10387 ( \10764 , \10759 );
or \U$10388 ( \10765 , \10763 , \10764 );
xor \U$10389 ( \10766 , \10109 , \10130 );
xor \U$10390 ( \10767 , \10766 , \10156 );
nand \U$10391 ( \10768 , \10765 , \10767 );
nand \U$10392 ( \10769 , \10762 , \10768 );
xor \U$10393 ( \10770 , \10355 , \10357 );
xor \U$10394 ( \10771 , \10770 , \10360 );
and \U$10395 ( \10772 , \10769 , \10771 );
xor \U$10396 ( \10773 , \9698 , \9699 );
xor \U$10397 ( \10774 , \10773 , \9702 );
xor \U$10398 ( \10775 , \10332 , \10339 );
xor \U$10399 ( \10776 , \10774 , \10775 );
xor \U$10400 ( \10777 , \10355 , \10357 );
xor \U$10401 ( \10778 , \10777 , \10360 );
and \U$10402 ( \10779 , \10776 , \10778 );
and \U$10403 ( \10780 , \10769 , \10776 );
or \U$10404 ( \10781 , \10772 , \10779 , \10780 );
and \U$10405 ( \10782 , \10757 , \10781 );
and \U$10406 ( \10783 , \10751 , \10756 );
or \U$10407 ( \10784 , \10782 , \10783 );
xor \U$10408 ( \10785 , \10349 , \10351 );
xor \U$10409 ( \10786 , \10082 , \10327 );
xor \U$10410 ( \10787 , \10786 , \10344 );
and \U$10411 ( \10788 , \10785 , \10787 );
xor \U$10412 ( \10789 , \9986 , \9988 );
xor \U$10413 ( \10790 , \10789 , \9991 );
xor \U$10414 ( \10791 , \10363 , \10370 );
xor \U$10415 ( \10792 , \10790 , \10791 );
xor \U$10416 ( \10793 , \10082 , \10327 );
xor \U$10417 ( \10794 , \10793 , \10344 );
and \U$10418 ( \10795 , \10792 , \10794 );
and \U$10419 ( \10796 , \10785 , \10792 );
or \U$10420 ( \10797 , \10788 , \10795 , \10796 );
xor \U$10421 ( \10798 , \10784 , \10797 );
xor \U$10422 ( \10799 , \9721 , \9958 );
xor \U$10423 ( \10800 , \10799 , \9975 );
xor \U$10424 ( \10801 , \10379 , \10386 );
xor \U$10425 ( \10802 , \10800 , \10801 );
and \U$10426 ( \10803 , \10798 , \10802 );
and \U$10427 ( \10804 , \10784 , \10797 );
or \U$10428 ( \10805 , \10803 , \10804 );
xor \U$10429 ( \10806 , \9978 , \9983 );
xor \U$10430 ( \10807 , \10806 , \10006 );
xor \U$10431 ( \10808 , \10805 , \10807 );
xor \U$10432 ( \10809 , \10378 , \10391 );
xor \U$10433 ( \10810 , \10809 , \10396 );
and \U$10434 ( \10811 , \10808 , \10810 );
and \U$10435 ( \10812 , \10805 , \10807 );
or \U$10436 ( \10813 , \10811 , \10812 );
xor \U$10437 ( \10814 , \10399 , \10401 );
xor \U$10438 ( \10815 , \10814 , \10408 );
and \U$10439 ( \10816 , \10813 , \10815 );
and \U$10440 ( \10817 , \10418 , \10816 );
xor \U$10441 ( \10818 , \10816 , \10418 );
xor \U$10442 ( \10819 , \10813 , \10815 );
xor \U$10443 ( \10820 , \10567 , \10646 );
xor \U$10444 ( \10821 , \10820 , \10728 );
xor \U$10445 ( \10822 , \10446 , \10456 );
xor \U$10446 ( \10823 , \10822 , \10479 );
and \U$10447 ( \10824 , \10821 , \10823 );
not \U$10448 ( \10825 , \10824 );
not \U$10449 ( \10826 , \10761 );
not \U$10450 ( \10827 , \10767 );
or \U$10451 ( \10828 , \10826 , \10827 );
or \U$10452 ( \10829 , \10767 , \10761 );
nand \U$10453 ( \10830 , \10828 , \10829 );
not \U$10454 ( \10831 , \10830 );
not \U$10455 ( \10832 , \10759 );
and \U$10456 ( \10833 , \10831 , \10832 );
and \U$10457 ( \10834 , \10830 , \10759 );
nor \U$10458 ( \10835 , \10833 , \10834 );
xor \U$10459 ( \10836 , \10507 , \10532 );
xor \U$10460 ( \10837 , \10836 , \10564 );
xor \U$10461 ( \10838 , \10593 , \10616 );
xor \U$10462 ( \10839 , \10838 , \10643 );
and \U$10463 ( \10840 , \10837 , \10839 );
xor \U$10464 ( \10841 , \10672 , \10699 );
xor \U$10465 ( \10842 , \10841 , \10725 );
xor \U$10466 ( \10843 , \10593 , \10616 );
xor \U$10467 ( \10844 , \10843 , \10643 );
and \U$10468 ( \10845 , \10842 , \10844 );
and \U$10469 ( \10846 , \10837 , \10842 );
or \U$10470 ( \10847 , \10840 , \10845 , \10846 );
not \U$10471 ( \10848 , \10847 );
or \U$10472 ( \10849 , \10835 , \10848 );
not \U$10473 ( \10850 , \10848 );
not \U$10474 ( \10851 , \10835 );
or \U$10475 ( \10852 , \10850 , \10851 );
xor \U$10476 ( \10853 , \10071 , \10073 );
xor \U$10477 ( \10854 , \10853 , \10076 );
xor \U$10478 ( \10855 , \10736 , \10743 );
xor \U$10479 ( \10856 , \10854 , \10855 );
nand \U$10480 ( \10857 , \10852 , \10856 );
nand \U$10481 ( \10858 , \10849 , \10857 );
not \U$10482 ( \10859 , \10858 );
or \U$10483 ( \10860 , \10825 , \10859 );
or \U$10484 ( \10861 , \10858 , \10824 );
xor \U$10485 ( \10862 , \10514 , \10521 );
xor \U$10486 ( \10863 , \10862 , \10529 );
xor \U$10487 ( \10864 , \10654 , \10661 );
xor \U$10488 ( \10865 , \10864 , \10669 );
xor \U$10489 ( \10866 , \10863 , \10865 );
xor \U$10490 ( \10867 , \10489 , \10496 );
xor \U$10491 ( \10868 , \10867 , \10504 );
and \U$10492 ( \10869 , \10866 , \10868 );
and \U$10493 ( \10870 , \10863 , \10865 );
or \U$10494 ( \10871 , \10869 , \10870 );
not \U$10495 ( \10872 , \10601 );
not \U$10496 ( \10873 , \10614 );
or \U$10497 ( \10874 , \10872 , \10873 );
or \U$10498 ( \10875 , \10601 , \10614 );
nand \U$10499 ( \10876 , \10874 , \10875 );
not \U$10500 ( \10877 , \10876 );
not \U$10501 ( \10878 , \10602 );
and \U$10502 ( \10879 , \10877 , \10878 );
and \U$10503 ( \10880 , \10876 , \10602 );
nor \U$10504 ( \10881 , \10879 , \10880 );
xor \U$10505 ( \10882 , \10624 , \10631 );
xor \U$10506 ( \10883 , \10882 , \10640 );
nand \U$10507 ( \10884 , \10881 , \10883 );
xor \U$10508 ( \10885 , \10871 , \10884 );
xor \U$10509 ( \10886 , \10574 , \10582 );
xor \U$10510 ( \10887 , \10886 , \10590 );
xor \U$10511 ( \10888 , \10679 , \10687 );
xor \U$10512 ( \10889 , \10888 , \10696 );
and \U$10513 ( \10890 , \10887 , \10889 );
xor \U$10514 ( \10891 , \10707 , \10714 );
xor \U$10515 ( \10892 , \10891 , \10722 );
xor \U$10516 ( \10893 , \10679 , \10687 );
xor \U$10517 ( \10894 , \10893 , \10696 );
and \U$10518 ( \10895 , \10892 , \10894 );
and \U$10519 ( \10896 , \10887 , \10892 );
or \U$10520 ( \10897 , \10890 , \10895 , \10896 );
and \U$10521 ( \10898 , \10885 , \10897 );
and \U$10522 ( \10899 , \10871 , \10884 );
or \U$10523 ( \10900 , \10898 , \10899 );
and \U$10524 ( \10901 , \8371 , RIae76a78_55);
and \U$10525 ( \10902 , RIae76988_53, \8369 );
nor \U$10526 ( \10903 , \10901 , \10902 );
and \U$10527 ( \10904 , \10903 , \8020 );
not \U$10528 ( \10905 , \10903 );
and \U$10529 ( \10906 , \10905 , \8019 );
nor \U$10530 ( \10907 , \10904 , \10906 );
and \U$10531 ( \10908 , \7633 , RIae762f8_39);
and \U$10532 ( \10909 , RIae76208_37, \7631 );
nor \U$10533 ( \10910 , \10908 , \10909 );
and \U$10534 ( \10911 , \10910 , \7206 );
not \U$10535 ( \10912 , \10910 );
and \U$10536 ( \10913 , \10912 , \7205 );
nor \U$10537 ( \10914 , \10911 , \10913 );
xor \U$10538 ( \10915 , \10907 , \10914 );
and \U$10539 ( \10916 , \8966 , RIae767a8_49);
and \U$10540 ( \10917 , RIae76898_51, \8964 );
nor \U$10541 ( \10918 , \10916 , \10917 );
and \U$10542 ( \10919 , \10918 , \8799 );
not \U$10543 ( \10920 , \10918 );
and \U$10544 ( \10921 , \10920 , \8789 );
nor \U$10545 ( \10922 , \10919 , \10921 );
and \U$10546 ( \10923 , \10915 , \10922 );
and \U$10547 ( \10924 , \10907 , \10914 );
or \U$10548 ( \10925 , \10923 , \10924 );
and \U$10549 ( \10926 , \10548 , RIae78cb0_128);
and \U$10550 ( \10927 , RIae78da0_130, \10546 );
nor \U$10551 ( \10928 , \10926 , \10927 );
and \U$10552 ( \10929 , \10928 , \10421 );
not \U$10553 ( \10930 , \10928 );
and \U$10554 ( \10931 , \10930 , \10118 );
nor \U$10555 ( \10932 , \10929 , \10931 );
not \U$10556 ( \10933 , RIae7a060_170);
not \U$10557 ( \10934 , RIae7a0d8_171);
or \U$10558 ( \10935 , \10933 , \10934 );
nand \U$10559 ( \10936 , \10935 , RIae7a150_172);
xor \U$10560 ( \10937 , \10932 , \10936 );
and \U$10561 ( \10938 , \9760 , RIae76b68_57);
and \U$10562 ( \10939 , RIae78a58_123, \9758 );
nor \U$10563 ( \10940 , \10938 , \10939 );
and \U$10564 ( \10941 , \10940 , \9273 );
not \U$10565 ( \10942 , \10940 );
and \U$10566 ( \10943 , \10942 , \9764 );
nor \U$10567 ( \10944 , \10941 , \10943 );
and \U$10568 ( \10945 , \10937 , \10944 );
and \U$10569 ( \10946 , \10932 , \10936 );
or \U$10570 ( \10947 , \10945 , \10946 );
xor \U$10571 ( \10948 , \10925 , \10947 );
and \U$10572 ( \10949 , \6172 , RIae766b8_47);
and \U$10573 ( \10950 , RIae765c8_45, \6170 );
nor \U$10574 ( \10951 , \10949 , \10950 );
and \U$10575 ( \10952 , \10951 , \6176 );
not \U$10576 ( \10953 , \10951 );
and \U$10577 ( \10954 , \10953 , \6175 );
nor \U$10578 ( \10955 , \10952 , \10954 );
and \U$10579 ( \10956 , \5896 , RIae763e8_41);
and \U$10580 ( \10957 , RIae764d8_43, \5894 );
nor \U$10581 ( \10958 , \10956 , \10957 );
and \U$10582 ( \10959 , \10958 , \5590 );
not \U$10583 ( \10960 , \10958 );
and \U$10584 ( \10961 , \10960 , \5589 );
nor \U$10585 ( \10962 , \10959 , \10961 );
xor \U$10586 ( \10963 , \10955 , \10962 );
and \U$10587 ( \10964 , \6941 , RIae76118_35);
and \U$10588 ( \10965 , RIae76028_33, \6939 );
nor \U$10589 ( \10966 , \10964 , \10965 );
and \U$10590 ( \10967 , \10966 , \6314 );
not \U$10591 ( \10968 , \10966 );
and \U$10592 ( \10969 , \10968 , \6945 );
nor \U$10593 ( \10970 , \10967 , \10969 );
and \U$10594 ( \10971 , \10963 , \10970 );
and \U$10595 ( \10972 , \10955 , \10962 );
or \U$10596 ( \10973 , \10971 , \10972 );
and \U$10597 ( \10974 , \10948 , \10973 );
and \U$10598 ( \10975 , \10925 , \10947 );
nor \U$10599 ( \10976 , \10974 , \10975 );
and \U$10600 ( \10977 , \4688 , RIae75218_3);
and \U$10601 ( \10978 , RIae75128_1, \4686 );
nor \U$10602 ( \10979 , \10977 , \10978 );
and \U$10603 ( \10980 , \10979 , \4481 );
not \U$10604 ( \10981 , \10979 );
and \U$10605 ( \10982 , \10981 , \4482 );
nor \U$10606 ( \10983 , \10980 , \10982 );
and \U$10607 ( \10984 , \4247 , RIae757b8_15);
and \U$10608 ( \10985 , RIae756c8_13, \4245 );
nor \U$10609 ( \10986 , \10984 , \10985 );
and \U$10610 ( \10987 , \10986 , \3989 );
not \U$10611 ( \10988 , \10986 );
and \U$10612 ( \10989 , \10988 , \4251 );
nor \U$10613 ( \10990 , \10987 , \10989 );
xor \U$10614 ( \10991 , \10983 , \10990 );
and \U$10615 ( \10992 , \5399 , RIae75308_5);
and \U$10616 ( \10993 , RIae753f8_7, \5397 );
nor \U$10617 ( \10994 , \10992 , \10993 );
and \U$10618 ( \10995 , \10994 , \5016 );
not \U$10619 ( \10996 , \10994 );
and \U$10620 ( \10997 , \10996 , \5403 );
nor \U$10621 ( \10998 , \10995 , \10997 );
and \U$10622 ( \10999 , \10991 , \10998 );
and \U$10623 ( \11000 , \10983 , \10990 );
or \U$10624 ( \11001 , \10999 , \11000 );
and \U$10625 ( \11002 , \1939 , RIae78788_117);
and \U$10626 ( \11003 , RIae78698_115, \1937 );
nor \U$10627 ( \11004 , \11002 , \11003 );
and \U$10628 ( \11005 , \11004 , \1735 );
not \U$10629 ( \11006 , \11004 );
and \U$10630 ( \11007 , \11006 , \1734 );
nor \U$10631 ( \11008 , \11005 , \11007 );
and \U$10632 ( \11009 , \2224 , RIae75b78_23);
and \U$10633 ( \11010 , RIae75a88_21, \2222 );
nor \U$10634 ( \11011 , \11009 , \11010 );
and \U$10635 ( \11012 , \11011 , \2061 );
not \U$10636 ( \11013 , \11011 );
and \U$10637 ( \11014 , \11013 , \2060 );
nor \U$10638 ( \11015 , \11012 , \11014 );
xor \U$10639 ( \11016 , \11008 , \11015 );
and \U$10640 ( \11017 , \2607 , RIae75998_19);
and \U$10641 ( \11018 , RIae758a8_17, \2605 );
nor \U$10642 ( \11019 , \11017 , \11018 );
and \U$10643 ( \11020 , \11019 , \2611 );
not \U$10644 ( \11021 , \11019 );
and \U$10645 ( \11022 , \11021 , \2397 );
nor \U$10646 ( \11023 , \11020 , \11022 );
and \U$10647 ( \11024 , \11016 , \11023 );
and \U$10648 ( \11025 , \11008 , \11015 );
or \U$10649 ( \11026 , \11024 , \11025 );
xor \U$10650 ( \11027 , \11001 , \11026 );
not \U$10651 ( \11028 , \2774 );
and \U$10652 ( \11029 , \3214 , RIae75c68_25);
and \U$10653 ( \11030 , RIae75d58_27, \3212 );
nor \U$10654 ( \11031 , \11029 , \11030 );
not \U$10655 ( \11032 , \11031 );
or \U$10656 ( \11033 , \11028 , \11032 );
or \U$10657 ( \11034 , \11031 , \2774 );
nand \U$10658 ( \11035 , \11033 , \11034 );
not \U$10659 ( \11036 , \2789 );
and \U$10660 ( \11037 , \2783 , RIae75f38_31);
and \U$10661 ( \11038 , RIae75e48_29, \2781 );
nor \U$10662 ( \11039 , \11037 , \11038 );
not \U$10663 ( \11040 , \11039 );
or \U$10664 ( \11041 , \11036 , \11040 );
or \U$10665 ( \11042 , \11039 , \3089 );
nand \U$10666 ( \11043 , \11041 , \11042 );
xor \U$10667 ( \11044 , \11035 , \11043 );
and \U$10668 ( \11045 , \3730 , RIae755d8_11);
and \U$10669 ( \11046 , RIae754e8_9, \3728 );
nor \U$10670 ( \11047 , \11045 , \11046 );
and \U$10671 ( \11048 , \11047 , \3732 );
not \U$10672 ( \11049 , \11047 );
and \U$10673 ( \11050 , \11049 , \3422 );
nor \U$10674 ( \11051 , \11048 , \11050 );
and \U$10675 ( \11052 , \11044 , \11051 );
and \U$10676 ( \11053 , \11035 , \11043 );
or \U$10677 ( \11054 , \11052 , \11053 );
and \U$10678 ( \11055 , \11027 , \11054 );
and \U$10679 ( \11056 , \11001 , \11026 );
nor \U$10680 ( \11057 , \11055 , \11056 );
xor \U$10681 ( \11058 , \10976 , \11057 );
and \U$10682 ( \11059 , \1593 , RIae78968_121);
and \U$10683 ( \11060 , RIae78878_119, \1591 );
nor \U$10684 ( \11061 , \11059 , \11060 );
and \U$10685 ( \11062 , \11061 , \1498 );
not \U$10686 ( \11063 , \11061 );
and \U$10687 ( \11064 , \11063 , \1488 );
nor \U$10688 ( \11065 , \11062 , \11064 );
and \U$10689 ( \11066 , \1138 , RIae77c48_93);
and \U$10690 ( \11067 , RIae77b58_91, \1136 );
nor \U$10691 ( \11068 , \11066 , \11067 );
and \U$10692 ( \11069 , \11068 , \1012 );
not \U$10693 ( \11070 , \11068 );
and \U$10694 ( \11071 , \11070 , \1142 );
nor \U$10695 ( \11072 , \11069 , \11071 );
xor \U$10696 ( \11073 , \11065 , \11072 );
and \U$10697 ( \11074 , \1376 , RIae77d38_95);
and \U$10698 ( \11075 , RIae77e28_97, \1374 );
nor \U$10699 ( \11076 , \11074 , \11075 );
and \U$10700 ( \11077 , \11076 , \1380 );
not \U$10701 ( \11078 , \11076 );
and \U$10702 ( \11079 , \11078 , \1261 );
nor \U$10703 ( \11080 , \11077 , \11079 );
and \U$10704 ( \11081 , \11073 , \11080 );
and \U$10705 ( \11082 , \11065 , \11072 );
or \U$10706 ( \11083 , \11081 , \11082 );
and \U$10707 ( \11084 , \672 , RIae781e8_105);
and \U$10708 ( \11085 , RIae785a8_113, \670 );
nor \U$10709 ( \11086 , \11084 , \11085 );
and \U$10710 ( \11087 , \11086 , \588 );
not \U$10711 ( \11088 , \11086 );
and \U$10712 ( \11089 , \11088 , \587 );
nor \U$10713 ( \11090 , \11087 , \11089 );
and \U$10714 ( \11091 , \558 , RIae77f18_99);
and \U$10715 ( \11092 , RIae78008_101, \556 );
nor \U$10716 ( \11093 , \11091 , \11092 );
and \U$10717 ( \11094 , \11093 , \504 );
not \U$10718 ( \11095 , \11093 );
and \U$10719 ( \11096 , \11095 , \562 );
nor \U$10720 ( \11097 , \11094 , \11096 );
xor \U$10721 ( \11098 , \11090 , \11097 );
not \U$10722 ( \11099 , \787 );
and \U$10723 ( \11100 , \883 , RIae783c8_109);
and \U$10724 ( \11101 , RIae78530_112, \881 );
nor \U$10725 ( \11102 , \11100 , \11101 );
not \U$10726 ( \11103 , \11102 );
or \U$10727 ( \11104 , \11099 , \11103 );
or \U$10728 ( \11105 , \11102 , \789 );
nand \U$10729 ( \11106 , \11104 , \11105 );
and \U$10730 ( \11107 , \11098 , \11106 );
and \U$10731 ( \11108 , \11090 , \11097 );
or \U$10732 ( \11109 , \11107 , \11108 );
xor \U$10733 ( \11110 , \11083 , \11109 );
not \U$10734 ( \11111 , \402 );
and \U$10735 ( \11112 , \436 , RIae771f8_71);
and \U$10736 ( \11113 , RIae772e8_73, \434 );
nor \U$10737 ( \11114 , \11112 , \11113 );
not \U$10738 ( \11115 , \11114 );
or \U$10739 ( \11116 , \11111 , \11115 );
or \U$10740 ( \11117 , \11114 , \402 );
nand \U$10741 ( \11118 , \11116 , \11117 );
not \U$10742 ( \11119 , \388 );
and \U$10743 ( \11120 , \384 , RIae77180_70);
and \U$10744 ( \11121 , RIae77018_67, \382 );
nor \U$10745 ( \11122 , \11120 , \11121 );
not \U$10746 ( \11123 , \11122 );
or \U$10747 ( \11124 , \11119 , \11123 );
or \U$10748 ( \11125 , \11122 , \388 );
nand \U$10749 ( \11126 , \11124 , \11125 );
xor \U$10750 ( \11127 , \11118 , \11126 );
not \U$10751 ( \11128 , \471 );
and \U$10752 ( \11129 , \514 , RIae782d8_107);
and \U$10753 ( \11130 , RIae780f8_103, \512 );
nor \U$10754 ( \11131 , \11129 , \11130 );
not \U$10755 ( \11132 , \11131 );
or \U$10756 ( \11133 , \11128 , \11132 );
or \U$10757 ( \11134 , \11131 , \469 );
nand \U$10758 ( \11135 , \11133 , \11134 );
and \U$10759 ( \11136 , \11127 , \11135 );
and \U$10760 ( \11137 , \11118 , \11126 );
or \U$10761 ( \11138 , \11136 , \11137 );
and \U$10762 ( \11139 , \11110 , \11138 );
and \U$10763 ( \11140 , \11083 , \11109 );
nor \U$10764 ( \11141 , \11139 , \11140 );
and \U$10765 ( \11142 , \11058 , \11141 );
and \U$10766 ( \11143 , \10976 , \11057 );
nor \U$10767 ( \11144 , \11142 , \11143 );
xor \U$10768 ( \11145 , \10900 , \11144 );
xor \U$10769 ( \11146 , \10448 , \10450 );
xor \U$10770 ( \11147 , \11146 , \10453 );
not \U$10771 ( \11148 , \10438 );
not \U$10772 ( \11149 , \10444 );
or \U$10773 ( \11150 , \11148 , \11149 );
or \U$10774 ( \11151 , \10438 , \10444 );
nand \U$10775 ( \11152 , \11150 , \11151 );
not \U$10776 ( \11153 , \11152 );
not \U$10777 ( \11154 , \10428 );
and \U$10778 ( \11155 , \11153 , \11154 );
and \U$10779 ( \11156 , \11152 , \10428 );
nor \U$10780 ( \11157 , \11155 , \11156 );
or \U$10781 ( \11158 , \11147 , \11157 );
not \U$10782 ( \11159 , \11157 );
not \U$10783 ( \11160 , \11147 );
or \U$10784 ( \11161 , \11159 , \11160 );
xor \U$10785 ( \11162 , \10463 , \10469 );
xor \U$10786 ( \11163 , \11162 , \10476 );
nand \U$10787 ( \11164 , \11161 , \11163 );
nand \U$10788 ( \11165 , \11158 , \11164 );
and \U$10789 ( \11166 , \11145 , \11165 );
and \U$10790 ( \11167 , \10900 , \11144 );
or \U$10791 ( \11168 , \11166 , \11167 );
nand \U$10792 ( \11169 , \10861 , \11168 );
nand \U$10793 ( \11170 , \10860 , \11169 );
xor \U$10794 ( \11171 , \10753 , \10755 );
not \U$10795 ( \11172 , \11171 );
xor \U$10796 ( \11173 , \10482 , \10731 );
xor \U$10797 ( \11174 , \11173 , \10748 );
not \U$10798 ( \11175 , \11174 );
or \U$10799 ( \11176 , \11172 , \11175 );
or \U$10800 ( \11177 , \11174 , \11171 );
xor \U$10801 ( \11178 , \10355 , \10357 );
xor \U$10802 ( \11179 , \11178 , \10360 );
xor \U$10803 ( \11180 , \10769 , \10776 );
xor \U$10804 ( \11181 , \11179 , \11180 );
nand \U$10805 ( \11182 , \11177 , \11181 );
nand \U$10806 ( \11183 , \11176 , \11182 );
xor \U$10807 ( \11184 , \11170 , \11183 );
xor \U$10808 ( \11185 , \10082 , \10327 );
xor \U$10809 ( \11186 , \11185 , \10344 );
xor \U$10810 ( \11187 , \10785 , \10792 );
xor \U$10811 ( \11188 , \11186 , \11187 );
and \U$10812 ( \11189 , \11184 , \11188 );
and \U$10813 ( \11190 , \11170 , \11183 );
or \U$10814 ( \11191 , \11189 , \11190 );
xor \U$10815 ( \11192 , \10347 , \10352 );
xor \U$10816 ( \11193 , \11192 , \10375 );
xor \U$10817 ( \11194 , \11191 , \11193 );
xor \U$10818 ( \11195 , \10784 , \10797 );
xor \U$10819 ( \11196 , \11195 , \10802 );
and \U$10820 ( \11197 , \11194 , \11196 );
and \U$10821 ( \11198 , \11191 , \11193 );
or \U$10822 ( \11199 , \11197 , \11198 );
xor \U$10823 ( \11200 , \10805 , \10807 );
xor \U$10824 ( \11201 , \11200 , \10810 );
and \U$10825 ( \11202 , \11199 , \11201 );
and \U$10826 ( \11203 , \10819 , \11202 );
xor \U$10827 ( \11204 , \11202 , \10819 );
xor \U$10828 ( \11205 , \11191 , \11193 );
xor \U$10829 ( \11206 , \11205 , \11196 );
not \U$10830 ( \11207 , \11206 );
xor \U$10831 ( \11208 , \11170 , \11183 );
xor \U$10832 ( \11209 , \11208 , \11188 );
xor \U$10833 ( \11210 , \10751 , \10756 );
xor \U$10834 ( \11211 , \11210 , \10781 );
and \U$10835 ( \11212 , \11209 , \11211 );
not \U$10836 ( \11213 , \11209 );
not \U$10837 ( \11214 , \11211 );
and \U$10838 ( \11215 , \11213 , \11214 );
xor \U$10839 ( \11216 , \10900 , \11144 );
xor \U$10840 ( \11217 , \11216 , \11165 );
xor \U$10841 ( \11218 , \10821 , \10823 );
and \U$10842 ( \11219 , \11217 , \11218 );
not \U$10843 ( \11220 , \11217 );
not \U$10844 ( \11221 , \11218 );
and \U$10845 ( \11222 , \11220 , \11221 );
xnor \U$10846 ( \11223 , \10848 , \10835 );
not \U$10847 ( \11224 , \11223 );
not \U$10848 ( \11225 , \10856 );
and \U$10849 ( \11226 , \11224 , \11225 );
and \U$10850 ( \11227 , \11223 , \10856 );
nor \U$10851 ( \11228 , \11226 , \11227 );
nor \U$10852 ( \11229 , \11222 , \11228 );
nor \U$10853 ( \11230 , \11219 , \11229 );
xor \U$10854 ( \11231 , \10593 , \10616 );
xor \U$10855 ( \11232 , \11231 , \10643 );
xor \U$10856 ( \11233 , \10837 , \10842 );
xor \U$10857 ( \11234 , \11232 , \11233 );
xor \U$10858 ( \11235 , \11083 , \11109 );
xor \U$10859 ( \11236 , \11235 , \11138 );
or \U$10860 ( \11237 , \10881 , \10883 );
nand \U$10861 ( \11238 , \11237 , \10884 );
xor \U$10862 ( \11239 , \11236 , \11238 );
xor \U$10863 ( \11240 , \11001 , \11026 );
xor \U$10864 ( \11241 , \11240 , \11054 );
and \U$10865 ( \11242 , \11239 , \11241 );
and \U$10866 ( \11243 , \11236 , \11238 );
or \U$10867 ( \11244 , \11242 , \11243 );
and \U$10868 ( \11245 , \11234 , \11244 );
not \U$10869 ( \11246 , \11234 );
not \U$10870 ( \11247 , \11244 );
and \U$10871 ( \11248 , \11246 , \11247 );
not \U$10872 ( \11249 , \11163 );
not \U$10873 ( \11250 , \11147 );
or \U$10874 ( \11251 , \11249 , \11250 );
or \U$10875 ( \11252 , \11147 , \11163 );
nand \U$10876 ( \11253 , \11251 , \11252 );
not \U$10877 ( \11254 , \11253 );
not \U$10878 ( \11255 , \11157 );
and \U$10879 ( \11256 , \11254 , \11255 );
and \U$10880 ( \11257 , \11253 , \11157 );
nor \U$10881 ( \11258 , \11256 , \11257 );
nor \U$10882 ( \11259 , \11248 , \11258 );
nor \U$10883 ( \11260 , \11245 , \11259 );
not \U$10884 ( \11261 , \11260 );
xor \U$10885 ( \11262 , \10976 , \11057 );
xor \U$10886 ( \11263 , \11262 , \11141 );
not \U$10887 ( \11264 , \11263 );
xor \U$10888 ( \11265 , \10871 , \10884 );
xor \U$10889 ( \11266 , \11265 , \10897 );
nand \U$10890 ( \11267 , \11264 , \11266 );
not \U$10891 ( \11268 , \11267 );
and \U$10892 ( \11269 , \11261 , \11268 );
and \U$10893 ( \11270 , \11260 , \11267 );
xor \U$10894 ( \11271 , \11065 , \11072 );
xor \U$10895 ( \11272 , \11271 , \11080 );
xor \U$10896 ( \11273 , \11008 , \11015 );
xor \U$10897 ( \11274 , \11273 , \11023 );
and \U$10898 ( \11275 , \11272 , \11274 );
xor \U$10899 ( \11276 , \11035 , \11043 );
xor \U$10900 ( \11277 , \11276 , \11051 );
xor \U$10901 ( \11278 , \11008 , \11015 );
xor \U$10902 ( \11279 , \11278 , \11023 );
and \U$10903 ( \11280 , \11277 , \11279 );
and \U$10904 ( \11281 , \11272 , \11277 );
or \U$10905 ( \11282 , \11275 , \11280 , \11281 );
not \U$10906 ( \11283 , RIae76c58_59);
nor \U$10907 ( \11284 , \11283 , \491 );
xor \U$10908 ( \11285 , \11118 , \11126 );
xor \U$10909 ( \11286 , \11285 , \11135 );
and \U$10910 ( \11287 , \11284 , \11286 );
xor \U$10911 ( \11288 , \11090 , \11097 );
xor \U$10912 ( \11289 , \11288 , \11106 );
xor \U$10913 ( \11290 , \11118 , \11126 );
xor \U$10914 ( \11291 , \11290 , \11135 );
and \U$10915 ( \11292 , \11289 , \11291 );
and \U$10916 ( \11293 , \11284 , \11289 );
or \U$10917 ( \11294 , \11287 , \11292 , \11293 );
xor \U$10918 ( \11295 , \11282 , \11294 );
xor \U$10919 ( \11296 , \10955 , \10962 );
xor \U$10920 ( \11297 , \11296 , \10970 );
xor \U$10921 ( \11298 , \10983 , \10990 );
xor \U$10922 ( \11299 , \11298 , \10998 );
xor \U$10923 ( \11300 , \11297 , \11299 );
xor \U$10924 ( \11301 , \10907 , \10914 );
xor \U$10925 ( \11302 , \11301 , \10922 );
and \U$10926 ( \11303 , \11300 , \11302 );
and \U$10927 ( \11304 , \11297 , \11299 );
or \U$10928 ( \11305 , \11303 , \11304 );
and \U$10929 ( \11306 , \11295 , \11305 );
and \U$10930 ( \11307 , \11282 , \11294 );
or \U$10931 ( \11308 , \11306 , \11307 );
and \U$10932 ( \11309 , \1138 , RIae78530_112);
and \U$10933 ( \11310 , RIae77c48_93, \1136 );
nor \U$10934 ( \11311 , \11309 , \11310 );
and \U$10935 ( \11312 , \11311 , \1012 );
not \U$10936 ( \11313 , \11311 );
and \U$10937 ( \11314 , \11313 , \1142 );
nor \U$10938 ( \11315 , \11312 , \11314 );
and \U$10939 ( \11316 , \1376 , RIae77b58_91);
and \U$10940 ( \11317 , RIae77d38_95, \1374 );
nor \U$10941 ( \11318 , \11316 , \11317 );
and \U$10942 ( \11319 , \11318 , \1380 );
not \U$10943 ( \11320 , \11318 );
and \U$10944 ( \11321 , \11320 , \1261 );
nor \U$10945 ( \11322 , \11319 , \11321 );
xor \U$10946 ( \11323 , \11315 , \11322 );
and \U$10947 ( \11324 , \1593 , RIae77e28_97);
and \U$10948 ( \11325 , RIae78968_121, \1591 );
nor \U$10949 ( \11326 , \11324 , \11325 );
and \U$10950 ( \11327 , \11326 , \1498 );
not \U$10951 ( \11328 , \11326 );
and \U$10952 ( \11329 , \11328 , \1488 );
nor \U$10953 ( \11330 , \11327 , \11329 );
and \U$10954 ( \11331 , \11323 , \11330 );
and \U$10955 ( \11332 , \11315 , \11322 );
or \U$10956 ( \11333 , \11331 , \11332 );
and \U$10957 ( \11334 , \384 , RIae76c58_59);
and \U$10958 ( \11335 , RIae77180_70, \382 );
nor \U$10959 ( \11336 , \11334 , \11335 );
not \U$10960 ( \11337 , \11336 );
not \U$10961 ( \11338 , \392 );
and \U$10962 ( \11339 , \11337 , \11338 );
and \U$10963 ( \11340 , \11336 , \392 );
nor \U$10964 ( \11341 , \11339 , \11340 );
and \U$10965 ( \11342 , \436 , RIae77018_67);
and \U$10966 ( \11343 , RIae771f8_71, \434 );
nor \U$10967 ( \11344 , \11342 , \11343 );
not \U$10968 ( \11345 , \11344 );
not \U$10969 ( \11346 , \400 );
and \U$10970 ( \11347 , \11345 , \11346 );
and \U$10971 ( \11348 , \11344 , \402 );
nor \U$10972 ( \11349 , \11347 , \11348 );
or \U$10973 ( \11350 , \11341 , \11349 );
not \U$10974 ( \11351 , \11349 );
not \U$10975 ( \11352 , \11341 );
or \U$10976 ( \11353 , \11351 , \11352 );
not \U$10977 ( \11354 , \469 );
and \U$10978 ( \11355 , \514 , RIae772e8_73);
and \U$10979 ( \11356 , RIae782d8_107, \512 );
nor \U$10980 ( \11357 , \11355 , \11356 );
not \U$10981 ( \11358 , \11357 );
or \U$10982 ( \11359 , \11354 , \11358 );
or \U$10983 ( \11360 , \11357 , \469 );
nand \U$10984 ( \11361 , \11359 , \11360 );
nand \U$10985 ( \11362 , \11353 , \11361 );
nand \U$10986 ( \11363 , \11350 , \11362 );
xor \U$10987 ( \11364 , \11333 , \11363 );
not \U$10988 ( \11365 , \787 );
and \U$10989 ( \11366 , \883 , RIae785a8_113);
and \U$10990 ( \11367 , RIae783c8_109, \881 );
nor \U$10991 ( \11368 , \11366 , \11367 );
not \U$10992 ( \11369 , \11368 );
or \U$10993 ( \11370 , \11365 , \11369 );
or \U$10994 ( \11371 , \11368 , \789 );
nand \U$10995 ( \11372 , \11370 , \11371 );
and \U$10996 ( \11373 , \558 , RIae780f8_103);
and \U$10997 ( \11374 , RIae77f18_99, \556 );
nor \U$10998 ( \11375 , \11373 , \11374 );
and \U$10999 ( \11376 , \11375 , \504 );
not \U$11000 ( \11377 , \11375 );
and \U$11001 ( \11378 , \11377 , \562 );
nor \U$11002 ( \11379 , \11376 , \11378 );
xor \U$11003 ( \11380 , \11372 , \11379 );
and \U$11004 ( \11381 , \672 , RIae78008_101);
and \U$11005 ( \11382 , RIae781e8_105, \670 );
nor \U$11006 ( \11383 , \11381 , \11382 );
and \U$11007 ( \11384 , \11383 , \588 );
not \U$11008 ( \11385 , \11383 );
and \U$11009 ( \11386 , \11385 , \587 );
nor \U$11010 ( \11387 , \11384 , \11386 );
and \U$11011 ( \11388 , \11380 , \11387 );
and \U$11012 ( \11389 , \11372 , \11379 );
or \U$11013 ( \11390 , \11388 , \11389 );
and \U$11014 ( \11391 , \11364 , \11390 );
and \U$11015 ( \11392 , \11333 , \11363 );
or \U$11016 ( \11393 , \11391 , \11392 );
and \U$11017 ( \11394 , \7633 , RIae76028_33);
and \U$11018 ( \11395 , RIae762f8_39, \7631 );
nor \U$11019 ( \11396 , \11394 , \11395 );
and \U$11020 ( \11397 , \11396 , \7206 );
not \U$11021 ( \11398 , \11396 );
and \U$11022 ( \11399 , \11398 , \7205 );
nor \U$11023 ( \11400 , \11397 , \11399 );
and \U$11024 ( \11401 , \8371 , RIae76208_37);
and \U$11025 ( \11402 , RIae76a78_55, \8369 );
nor \U$11026 ( \11403 , \11401 , \11402 );
and \U$11027 ( \11404 , \11403 , \8020 );
not \U$11028 ( \11405 , \11403 );
and \U$11029 ( \11406 , \11405 , \8019 );
nor \U$11030 ( \11407 , \11404 , \11406 );
xor \U$11031 ( \11408 , \11400 , \11407 );
and \U$11032 ( \11409 , \8966 , RIae76988_53);
and \U$11033 ( \11410 , RIae767a8_49, \8964 );
nor \U$11034 ( \11411 , \11409 , \11410 );
and \U$11035 ( \11412 , \11411 , \8799 );
not \U$11036 ( \11413 , \11411 );
and \U$11037 ( \11414 , \11413 , \8789 );
nor \U$11038 ( \11415 , \11412 , \11414 );
and \U$11039 ( \11416 , \11408 , \11415 );
and \U$11040 ( \11417 , \11400 , \11407 );
or \U$11041 ( \11418 , \11416 , \11417 );
and \U$11042 ( \11419 , \6172 , RIae764d8_43);
and \U$11043 ( \11420 , RIae766b8_47, \6170 );
nor \U$11044 ( \11421 , \11419 , \11420 );
and \U$11045 ( \11422 , \11421 , \6176 );
not \U$11046 ( \11423 , \11421 );
and \U$11047 ( \11424 , \11423 , \6175 );
nor \U$11048 ( \11425 , \11422 , \11424 );
and \U$11049 ( \11426 , \5896 , RIae753f8_7);
and \U$11050 ( \11427 , RIae763e8_41, \5894 );
nor \U$11051 ( \11428 , \11426 , \11427 );
and \U$11052 ( \11429 , \11428 , \5590 );
not \U$11053 ( \11430 , \11428 );
and \U$11054 ( \11431 , \11430 , \5589 );
nor \U$11055 ( \11432 , \11429 , \11431 );
xor \U$11056 ( \11433 , \11425 , \11432 );
and \U$11057 ( \11434 , \6941 , RIae765c8_45);
and \U$11058 ( \11435 , RIae76118_35, \6939 );
nor \U$11059 ( \11436 , \11434 , \11435 );
and \U$11060 ( \11437 , \11436 , \6314 );
not \U$11061 ( \11438 , \11436 );
and \U$11062 ( \11439 , \11438 , \6945 );
nor \U$11063 ( \11440 , \11437 , \11439 );
and \U$11064 ( \11441 , \11433 , \11440 );
and \U$11065 ( \11442 , \11425 , \11432 );
or \U$11066 ( \11443 , \11441 , \11442 );
xor \U$11067 ( \11444 , \11418 , \11443 );
and \U$11068 ( \11445 , \9760 , RIae76898_51);
and \U$11069 ( \11446 , RIae76b68_57, \9758 );
nor \U$11070 ( \11447 , \11445 , \11446 );
and \U$11071 ( \11448 , \11447 , \9272 );
not \U$11072 ( \11449 , \11447 );
and \U$11073 ( \11450 , \11449 , \9273 );
nor \U$11074 ( \11451 , \11448 , \11450 );
and \U$11075 ( \11452 , \10548 , RIae78a58_123);
and \U$11076 ( \11453 , RIae78cb0_128, \10546 );
nor \U$11077 ( \11454 , \11452 , \11453 );
and \U$11078 ( \11455 , \11454 , \10118 );
not \U$11079 ( \11456 , \11454 );
and \U$11080 ( \11457 , \11456 , \10421 );
nor \U$11081 ( \11458 , \11455 , \11457 );
or \U$11082 ( \11459 , \11451 , \11458 );
not \U$11083 ( \11460 , \11458 );
not \U$11084 ( \11461 , \11451 );
or \U$11085 ( \11462 , \11460 , \11461 );
and \U$11086 ( \11463 , RIae7a150_172, RIae7a0d8_171);
not \U$11087 ( \11464 , RIae7a0d8_171);
nor \U$11088 ( \11465 , \11464 , RIae7a060_170);
not \U$11089 ( \11466 , RIae7a060_170);
nor \U$11090 ( \11467 , \11466 , RIae7a0d8_171);
or \U$11091 ( \11468 , \11465 , \11467 );
nor \U$11092 ( \11469 , RIae7a150_172, RIae7a0d8_171);
nor \U$11093 ( \11470 , \11463 , \11468 , \11469 );
nand \U$11094 ( \11471 , RIae78da0_130, \11470 );
and \U$11095 ( \11472 , \11471 , \10936 );
not \U$11096 ( \11473 , \11471 );
not \U$11097 ( \11474 , \10936 );
and \U$11098 ( \11475 , \11473 , \11474 );
nor \U$11099 ( \11476 , \11472 , \11475 );
nand \U$11100 ( \11477 , \11462 , \11476 );
nand \U$11101 ( \11478 , \11459 , \11477 );
and \U$11102 ( \11479 , \11444 , \11478 );
and \U$11103 ( \11480 , \11418 , \11443 );
or \U$11104 ( \11481 , \11479 , \11480 );
xor \U$11105 ( \11482 , \11393 , \11481 );
not \U$11106 ( \11483 , \3089 );
and \U$11107 ( \11484 , \2783 , RIae758a8_17);
and \U$11108 ( \11485 , RIae75f38_31, \2781 );
nor \U$11109 ( \11486 , \11484 , \11485 );
not \U$11110 ( \11487 , \11486 );
or \U$11111 ( \11488 , \11483 , \11487 );
or \U$11112 ( \11489 , \11486 , \2789 );
nand \U$11113 ( \11490 , \11488 , \11489 );
not \U$11114 ( \11491 , \2774 );
and \U$11115 ( \11492 , \3214 , RIae75e48_29);
and \U$11116 ( \11493 , RIae75c68_25, \3212 );
nor \U$11117 ( \11494 , \11492 , \11493 );
not \U$11118 ( \11495 , \11494 );
or \U$11119 ( \11496 , \11491 , \11495 );
or \U$11120 ( \11497 , \11494 , \2774 );
nand \U$11121 ( \11498 , \11496 , \11497 );
xor \U$11122 ( \11499 , \11490 , \11498 );
and \U$11123 ( \11500 , \3730 , RIae75d58_27);
and \U$11124 ( \11501 , RIae755d8_11, \3728 );
nor \U$11125 ( \11502 , \11500 , \11501 );
and \U$11126 ( \11503 , \11502 , \3732 );
not \U$11127 ( \11504 , \11502 );
and \U$11128 ( \11505 , \11504 , \3422 );
nor \U$11129 ( \11506 , \11503 , \11505 );
and \U$11130 ( \11507 , \11499 , \11506 );
and \U$11131 ( \11508 , \11490 , \11498 );
or \U$11132 ( \11509 , \11507 , \11508 );
and \U$11133 ( \11510 , \2607 , RIae75a88_21);
and \U$11134 ( \11511 , RIae75998_19, \2605 );
nor \U$11135 ( \11512 , \11510 , \11511 );
and \U$11136 ( \11513 , \11512 , \2611 );
not \U$11137 ( \11514 , \11512 );
and \U$11138 ( \11515 , \11514 , \2397 );
nor \U$11139 ( \11516 , \11513 , \11515 );
and \U$11140 ( \11517 , \1939 , RIae78878_119);
and \U$11141 ( \11518 , RIae78788_117, \1937 );
nor \U$11142 ( \11519 , \11517 , \11518 );
and \U$11143 ( \11520 , \11519 , \1735 );
not \U$11144 ( \11521 , \11519 );
and \U$11145 ( \11522 , \11521 , \1734 );
nor \U$11146 ( \11523 , \11520 , \11522 );
xor \U$11147 ( \11524 , \11516 , \11523 );
and \U$11148 ( \11525 , \2224 , RIae78698_115);
and \U$11149 ( \11526 , RIae75b78_23, \2222 );
nor \U$11150 ( \11527 , \11525 , \11526 );
and \U$11151 ( \11528 , \11527 , \2061 );
not \U$11152 ( \11529 , \11527 );
and \U$11153 ( \11530 , \11529 , \2060 );
nor \U$11154 ( \11531 , \11528 , \11530 );
and \U$11155 ( \11532 , \11524 , \11531 );
and \U$11156 ( \11533 , \11516 , \11523 );
or \U$11157 ( \11534 , \11532 , \11533 );
xor \U$11158 ( \11535 , \11509 , \11534 );
and \U$11159 ( \11536 , \5399 , RIae75128_1);
and \U$11160 ( \11537 , RIae75308_5, \5397 );
nor \U$11161 ( \11538 , \11536 , \11537 );
and \U$11162 ( \11539 , \11538 , \5016 );
not \U$11163 ( \11540 , \11538 );
and \U$11164 ( \11541 , \11540 , \5403 );
nor \U$11165 ( \11542 , \11539 , \11541 );
and \U$11166 ( \11543 , \4247 , RIae754e8_9);
and \U$11167 ( \11544 , RIae757b8_15, \4245 );
nor \U$11168 ( \11545 , \11543 , \11544 );
and \U$11169 ( \11546 , \11545 , \3989 );
not \U$11170 ( \11547 , \11545 );
and \U$11171 ( \11548 , \11547 , \4251 );
nor \U$11172 ( \11549 , \11546 , \11548 );
xor \U$11173 ( \11550 , \11542 , \11549 );
and \U$11174 ( \11551 , \4688 , RIae756c8_13);
and \U$11175 ( \11552 , RIae75218_3, \4686 );
nor \U$11176 ( \11553 , \11551 , \11552 );
and \U$11177 ( \11554 , \11553 , \4481 );
not \U$11178 ( \11555 , \11553 );
and \U$11179 ( \11556 , \11555 , \4482 );
nor \U$11180 ( \11557 , \11554 , \11556 );
and \U$11181 ( \11558 , \11550 , \11557 );
and \U$11182 ( \11559 , \11542 , \11549 );
or \U$11183 ( \11560 , \11558 , \11559 );
and \U$11184 ( \11561 , \11535 , \11560 );
and \U$11185 ( \11562 , \11509 , \11534 );
or \U$11186 ( \11563 , \11561 , \11562 );
and \U$11187 ( \11564 , \11482 , \11563 );
and \U$11188 ( \11565 , \11393 , \11481 );
or \U$11189 ( \11566 , \11564 , \11565 );
xor \U$11190 ( \11567 , \11308 , \11566 );
xor \U$11191 ( \11568 , \10540 , \10553 );
xor \U$11192 ( \11569 , \11568 , \10561 );
xor \U$11193 ( \11570 , \10863 , \10865 );
xor \U$11194 ( \11571 , \11570 , \10868 );
and \U$11195 ( \11572 , \11569 , \11571 );
xor \U$11196 ( \11573 , \10679 , \10687 );
xor \U$11197 ( \11574 , \11573 , \10696 );
xor \U$11198 ( \11575 , \10887 , \10892 );
xor \U$11199 ( \11576 , \11574 , \11575 );
xor \U$11200 ( \11577 , \10863 , \10865 );
xor \U$11201 ( \11578 , \11577 , \10868 );
and \U$11202 ( \11579 , \11576 , \11578 );
and \U$11203 ( \11580 , \11569 , \11576 );
or \U$11204 ( \11581 , \11572 , \11579 , \11580 );
and \U$11205 ( \11582 , \11567 , \11581 );
and \U$11206 ( \11583 , \11308 , \11566 );
nor \U$11207 ( \11584 , \11582 , \11583 );
nor \U$11208 ( \11585 , \11270 , \11584 );
nor \U$11209 ( \11586 , \11269 , \11585 );
xor \U$11210 ( \11587 , \11230 , \11586 );
xnor \U$11211 ( \11588 , \11174 , \11181 );
not \U$11212 ( \11589 , \11588 );
not \U$11213 ( \11590 , \11171 );
and \U$11214 ( \11591 , \11589 , \11590 );
and \U$11215 ( \11592 , \11588 , \11171 );
nor \U$11216 ( \11593 , \11591 , \11592 );
and \U$11217 ( \11594 , \11587 , \11593 );
and \U$11218 ( \11595 , \11230 , \11586 );
or \U$11219 ( \11596 , \11594 , \11595 );
nor \U$11220 ( \11597 , \11215 , \11596 );
nor \U$11221 ( \11598 , \11212 , \11597 );
not \U$11222 ( \11599 , \11598 );
or \U$11223 ( \11600 , \11207 , \11599 );
or \U$11224 ( \11601 , \11598 , \11206 );
nand \U$11225 ( \11602 , \11600 , \11601 );
not \U$11226 ( \11603 , \11209 );
not \U$11227 ( \11604 , \11596 );
not \U$11228 ( \11605 , \11211 );
and \U$11229 ( \11606 , \11604 , \11605 );
and \U$11230 ( \11607 , \11596 , \11211 );
nor \U$11231 ( \11608 , \11606 , \11607 );
not \U$11232 ( \11609 , \11608 );
or \U$11233 ( \11610 , \11603 , \11609 );
or \U$11234 ( \11611 , \11608 , \11209 );
nand \U$11235 ( \11612 , \11610 , \11611 );
not \U$11236 ( \11613 , \11612 );
xnor \U$11237 ( \11614 , \11168 , \10858 );
not \U$11238 ( \11615 , \11614 );
not \U$11239 ( \11616 , \10824 );
and \U$11240 ( \11617 , \11615 , \11616 );
and \U$11241 ( \11618 , \11614 , \10824 );
nor \U$11242 ( \11619 , \11617 , \11618 );
xor \U$11243 ( \11620 , \11230 , \11586 );
xor \U$11244 ( \11621 , \11620 , \11593 );
and \U$11245 ( \11622 , \11619 , \11621 );
not \U$11246 ( \11623 , \11218 );
not \U$11247 ( \11624 , \11228 );
not \U$11248 ( \11625 , \11217 );
and \U$11249 ( \11626 , \11624 , \11625 );
and \U$11250 ( \11627 , \11228 , \11217 );
nor \U$11251 ( \11628 , \11626 , \11627 );
not \U$11252 ( \11629 , \11628 );
or \U$11253 ( \11630 , \11623 , \11629 );
or \U$11254 ( \11631 , \11628 , \11218 );
nand \U$11255 ( \11632 , \11630 , \11631 );
xor \U$11256 ( \11633 , \11308 , \11566 );
xor \U$11257 ( \11634 , \11633 , \11581 );
not \U$11258 ( \11635 , \11263 );
not \U$11259 ( \11636 , \11266 );
or \U$11260 ( \11637 , \11635 , \11636 );
or \U$11261 ( \11638 , \11266 , \11263 );
nand \U$11262 ( \11639 , \11637 , \11638 );
xor \U$11263 ( \11640 , \11634 , \11639 );
not \U$11264 ( \11641 , \11258 );
xor \U$11265 ( \11642 , \11244 , \11234 );
not \U$11266 ( \11643 , \11642 );
or \U$11267 ( \11644 , \11641 , \11643 );
or \U$11268 ( \11645 , \11642 , \11258 );
nand \U$11269 ( \11646 , \11644 , \11645 );
and \U$11270 ( \11647 , \11640 , \11646 );
and \U$11271 ( \11648 , \11634 , \11639 );
or \U$11272 ( \11649 , \11647 , \11648 );
xor \U$11273 ( \11650 , \11632 , \11649 );
xor \U$11274 ( \11651 , \11333 , \11363 );
xor \U$11275 ( \11652 , \11651 , \11390 );
xor \U$11276 ( \11653 , \11509 , \11534 );
xor \U$11277 ( \11654 , \11653 , \11560 );
and \U$11278 ( \11655 , \11652 , \11654 );
xor \U$11279 ( \11656 , \11118 , \11126 );
xor \U$11280 ( \11657 , \11656 , \11135 );
xor \U$11281 ( \11658 , \11284 , \11289 );
xor \U$11282 ( \11659 , \11657 , \11658 );
xor \U$11283 ( \11660 , \11509 , \11534 );
xor \U$11284 ( \11661 , \11660 , \11560 );
and \U$11285 ( \11662 , \11659 , \11661 );
and \U$11286 ( \11663 , \11652 , \11659 );
or \U$11287 ( \11664 , \11655 , \11662 , \11663 );
xor \U$11288 ( \11665 , \10925 , \10947 );
xor \U$11289 ( \11666 , \11665 , \10973 );
xor \U$11290 ( \11667 , \11664 , \11666 );
xor \U$11291 ( \11668 , \11236 , \11238 );
xor \U$11292 ( \11669 , \11668 , \11241 );
and \U$11293 ( \11670 , \11667 , \11669 );
and \U$11294 ( \11671 , \11664 , \11666 );
or \U$11295 ( \11672 , \11670 , \11671 );
xor \U$11296 ( \11673 , \11490 , \11498 );
xor \U$11297 ( \11674 , \11673 , \11506 );
xor \U$11298 ( \11675 , \11542 , \11549 );
xor \U$11299 ( \11676 , \11675 , \11557 );
and \U$11300 ( \11677 , \11674 , \11676 );
xor \U$11301 ( \11678 , \11425 , \11432 );
xor \U$11302 ( \11679 , \11678 , \11440 );
xor \U$11303 ( \11680 , \11542 , \11549 );
xor \U$11304 ( \11681 , \11680 , \11557 );
and \U$11305 ( \11682 , \11679 , \11681 );
and \U$11306 ( \11683 , \11674 , \11679 );
or \U$11307 ( \11684 , \11677 , \11682 , \11683 );
nand \U$11308 ( \11685 , RIae76d48_61, RIae78b48_125);
not \U$11309 ( \11686 , \11349 );
not \U$11310 ( \11687 , \11361 );
or \U$11311 ( \11688 , \11686 , \11687 );
or \U$11312 ( \11689 , \11349 , \11361 );
nand \U$11313 ( \11690 , \11688 , \11689 );
not \U$11314 ( \11691 , \11690 );
not \U$11315 ( \11692 , \11341 );
and \U$11316 ( \11693 , \11691 , \11692 );
and \U$11317 ( \11694 , \11690 , \11341 );
nor \U$11318 ( \11695 , \11693 , \11694 );
nand \U$11319 ( \11696 , \11685 , \11695 );
xor \U$11320 ( \11697 , \11684 , \11696 );
xor \U$11321 ( \11698 , \11516 , \11523 );
xor \U$11322 ( \11699 , \11698 , \11531 );
xor \U$11323 ( \11700 , \11372 , \11379 );
xor \U$11324 ( \11701 , \11700 , \11387 );
xor \U$11325 ( \11702 , \11699 , \11701 );
xor \U$11326 ( \11703 , \11315 , \11322 );
xor \U$11327 ( \11704 , \11703 , \11330 );
and \U$11328 ( \11705 , \11702 , \11704 );
and \U$11329 ( \11706 , \11699 , \11701 );
or \U$11330 ( \11707 , \11705 , \11706 );
and \U$11331 ( \11708 , \11697 , \11707 );
and \U$11332 ( \11709 , \11684 , \11696 );
or \U$11333 ( \11710 , \11708 , \11709 );
and \U$11334 ( \11711 , \5399 , RIae75218_3);
and \U$11335 ( \11712 , RIae75128_1, \5397 );
nor \U$11336 ( \11713 , \11711 , \11712 );
and \U$11337 ( \11714 , \11713 , \5403 );
not \U$11338 ( \11715 , \11713 );
and \U$11339 ( \11716 , \11715 , \5016 );
nor \U$11340 ( \11717 , \11714 , \11716 );
and \U$11341 ( \11718 , \5896 , RIae75308_5);
and \U$11342 ( \11719 , RIae753f8_7, \5894 );
nor \U$11343 ( \11720 , \11718 , \11719 );
and \U$11344 ( \11721 , \11720 , \5589 );
not \U$11345 ( \11722 , \11720 );
and \U$11346 ( \11723 , \11722 , \5590 );
nor \U$11347 ( \11724 , \11721 , \11723 );
xor \U$11348 ( \11725 , \11717 , \11724 );
and \U$11349 ( \11726 , \4688 , RIae757b8_15);
and \U$11350 ( \11727 , RIae756c8_13, \4686 );
nor \U$11351 ( \11728 , \11726 , \11727 );
and \U$11352 ( \11729 , \11728 , \4482 );
not \U$11353 ( \11730 , \11728 );
and \U$11354 ( \11731 , \11730 , \4481 );
nor \U$11355 ( \11732 , \11729 , \11731 );
and \U$11356 ( \11733 , \11725 , \11732 );
and \U$11357 ( \11734 , \11717 , \11724 );
nor \U$11358 ( \11735 , \11733 , \11734 );
and \U$11359 ( \11736 , \2607 , RIae75b78_23);
and \U$11360 ( \11737 , RIae75a88_21, \2605 );
nor \U$11361 ( \11738 , \11736 , \11737 );
and \U$11362 ( \11739 , \11738 , \2397 );
not \U$11363 ( \11740 , \11738 );
and \U$11364 ( \11741 , \11740 , \2611 );
nor \U$11365 ( \11742 , \11739 , \11741 );
and \U$11366 ( \11743 , \2783 , RIae75998_19);
and \U$11367 ( \11744 , RIae758a8_17, \2781 );
nor \U$11368 ( \11745 , \11743 , \11744 );
not \U$11369 ( \11746 , \11745 );
not \U$11370 ( \11747 , \3089 );
and \U$11371 ( \11748 , \11746 , \11747 );
and \U$11372 ( \11749 , \11745 , \3089 );
nor \U$11373 ( \11750 , \11748 , \11749 );
xor \U$11374 ( \11751 , \11742 , \11750 );
and \U$11375 ( \11752 , \2224 , RIae78788_117);
and \U$11376 ( \11753 , RIae78698_115, \2222 );
nor \U$11377 ( \11754 , \11752 , \11753 );
and \U$11378 ( \11755 , \11754 , \2060 );
not \U$11379 ( \11756 , \11754 );
and \U$11380 ( \11757 , \11756 , \2061 );
nor \U$11381 ( \11758 , \11755 , \11757 );
and \U$11382 ( \11759 , \11751 , \11758 );
and \U$11383 ( \11760 , \11742 , \11750 );
nor \U$11384 ( \11761 , \11759 , \11760 );
xor \U$11385 ( \11762 , \11735 , \11761 );
and \U$11386 ( \11763 , \3214 , RIae75f38_31);
and \U$11387 ( \11764 , RIae75e48_29, \3212 );
nor \U$11388 ( \11765 , \11763 , \11764 );
not \U$11389 ( \11766 , \11765 );
not \U$11390 ( \11767 , \2774 );
and \U$11391 ( \11768 , \11766 , \11767 );
and \U$11392 ( \11769 , \11765 , \2774 );
nor \U$11393 ( \11770 , \11768 , \11769 );
and \U$11394 ( \11771 , \3730 , RIae75c68_25);
and \U$11395 ( \11772 , RIae75d58_27, \3728 );
nor \U$11396 ( \11773 , \11771 , \11772 );
and \U$11397 ( \11774 , \11773 , \3422 );
not \U$11398 ( \11775 , \11773 );
and \U$11399 ( \11776 , \11775 , \3732 );
nor \U$11400 ( \11777 , \11774 , \11776 );
or \U$11401 ( \11778 , \11770 , \11777 );
not \U$11402 ( \11779 , \11777 );
not \U$11403 ( \11780 , \11770 );
or \U$11404 ( \11781 , \11779 , \11780 );
and \U$11405 ( \11782 , \4247 , RIae755d8_11);
and \U$11406 ( \11783 , RIae754e8_9, \4245 );
nor \U$11407 ( \11784 , \11782 , \11783 );
and \U$11408 ( \11785 , \11784 , \3989 );
not \U$11409 ( \11786 , \11784 );
and \U$11410 ( \11787 , \11786 , \4251 );
nor \U$11411 ( \11788 , \11785 , \11787 );
nand \U$11412 ( \11789 , \11781 , \11788 );
nand \U$11413 ( \11790 , \11778 , \11789 );
and \U$11414 ( \11791 , \11762 , \11790 );
and \U$11415 ( \11792 , \11735 , \11761 );
or \U$11416 ( \11793 , \11791 , \11792 );
and \U$11417 ( \11794 , \6941 , RIae766b8_47);
and \U$11418 ( \11795 , RIae765c8_45, \6939 );
nor \U$11419 ( \11796 , \11794 , \11795 );
and \U$11420 ( \11797 , \11796 , \6945 );
not \U$11421 ( \11798 , \11796 );
and \U$11422 ( \11799 , \11798 , \6314 );
nor \U$11423 ( \11800 , \11797 , \11799 );
and \U$11424 ( \11801 , \7633 , RIae76118_35);
and \U$11425 ( \11802 , RIae76028_33, \7631 );
nor \U$11426 ( \11803 , \11801 , \11802 );
and \U$11427 ( \11804 , \11803 , \7205 );
not \U$11428 ( \11805 , \11803 );
and \U$11429 ( \11806 , \11805 , \7206 );
nor \U$11430 ( \11807 , \11804 , \11806 );
xor \U$11431 ( \11808 , \11800 , \11807 );
and \U$11432 ( \11809 , \6172 , RIae763e8_41);
and \U$11433 ( \11810 , RIae764d8_43, \6170 );
nor \U$11434 ( \11811 , \11809 , \11810 );
and \U$11435 ( \11812 , \11811 , \6175 );
not \U$11436 ( \11813 , \11811 );
and \U$11437 ( \11814 , \11813 , \6176 );
nor \U$11438 ( \11815 , \11812 , \11814 );
and \U$11439 ( \11816 , \11808 , \11815 );
and \U$11440 ( \11817 , \11800 , \11807 );
nor \U$11441 ( \11818 , \11816 , \11817 );
and \U$11442 ( \11819 , \10548 , RIae76b68_57);
and \U$11443 ( \11820 , RIae78a58_123, \10546 );
nor \U$11444 ( \11821 , \11819 , \11820 );
and \U$11445 ( \11822 , \11821 , \10118 );
not \U$11446 ( \11823 , \11821 );
and \U$11447 ( \11824 , \11823 , \10421 );
nor \U$11448 ( \11825 , \11822 , \11824 );
nand \U$11449 ( \11826 , RIae7a7e0_186, RIae7a948_189);
and \U$11450 ( \11827 , \11826 , RIae7a060_170);
or \U$11451 ( \11828 , \11825 , \11827 );
not \U$11452 ( \11829 , \11827 );
not \U$11453 ( \11830 , \11825 );
or \U$11454 ( \11831 , \11829 , \11830 );
and \U$11455 ( \11832 , \11470 , RIae78cb0_128);
and \U$11456 ( \11833 , RIae78da0_130, \11468 );
nor \U$11457 ( \11834 , \11832 , \11833 );
and \U$11458 ( \11835 , \11834 , \10936 );
not \U$11459 ( \11836 , \11834 );
and \U$11460 ( \11837 , \11836 , \11474 );
nor \U$11461 ( \11838 , \11835 , \11837 );
nand \U$11462 ( \11839 , \11831 , \11838 );
nand \U$11463 ( \11840 , \11828 , \11839 );
xor \U$11464 ( \11841 , \11818 , \11840 );
and \U$11465 ( \11842 , \8371 , RIae762f8_39);
and \U$11466 ( \11843 , RIae76208_37, \8369 );
nor \U$11467 ( \11844 , \11842 , \11843 );
and \U$11468 ( \11845 , \11844 , \8019 );
not \U$11469 ( \11846 , \11844 );
and \U$11470 ( \11847 , \11846 , \8020 );
nor \U$11471 ( \11848 , \11845 , \11847 );
and \U$11472 ( \11849 , \8966 , RIae76a78_55);
and \U$11473 ( \11850 , RIae76988_53, \8964 );
nor \U$11474 ( \11851 , \11849 , \11850 );
and \U$11475 ( \11852 , \11851 , \8789 );
not \U$11476 ( \11853 , \11851 );
and \U$11477 ( \11854 , \11853 , \8799 );
nor \U$11478 ( \11855 , \11852 , \11854 );
or \U$11479 ( \11856 , \11848 , \11855 );
not \U$11480 ( \11857 , \11855 );
not \U$11481 ( \11858 , \11848 );
or \U$11482 ( \11859 , \11857 , \11858 );
and \U$11483 ( \11860 , \9760 , RIae767a8_49);
and \U$11484 ( \11861 , RIae76898_51, \9758 );
nor \U$11485 ( \11862 , \11860 , \11861 );
and \U$11486 ( \11863 , \11862 , \9273 );
not \U$11487 ( \11864 , \11862 );
and \U$11488 ( \11865 , \11864 , \9764 );
nor \U$11489 ( \11866 , \11863 , \11865 );
nand \U$11490 ( \11867 , \11859 , \11866 );
nand \U$11491 ( \11868 , \11856 , \11867 );
and \U$11492 ( \11869 , \11841 , \11868 );
and \U$11493 ( \11870 , \11818 , \11840 );
or \U$11494 ( \11871 , \11869 , \11870 );
xor \U$11495 ( \11872 , \11793 , \11871 );
and \U$11496 ( \11873 , \1593 , RIae77d38_95);
and \U$11497 ( \11874 , RIae77e28_97, \1591 );
nor \U$11498 ( \11875 , \11873 , \11874 );
and \U$11499 ( \11876 , \11875 , \1498 );
not \U$11500 ( \11877 , \11875 );
and \U$11501 ( \11878 , \11877 , \1488 );
nor \U$11502 ( \11879 , \11876 , \11878 );
and \U$11503 ( \11880 , \1376 , RIae77c48_93);
and \U$11504 ( \11881 , RIae77b58_91, \1374 );
nor \U$11505 ( \11882 , \11880 , \11881 );
and \U$11506 ( \11883 , \11882 , \1380 );
not \U$11507 ( \11884 , \11882 );
and \U$11508 ( \11885 , \11884 , \1261 );
nor \U$11509 ( \11886 , \11883 , \11885 );
xor \U$11510 ( \11887 , \11879 , \11886 );
and \U$11511 ( \11888 , \1939 , RIae78968_121);
and \U$11512 ( \11889 , RIae78878_119, \1937 );
nor \U$11513 ( \11890 , \11888 , \11889 );
and \U$11514 ( \11891 , \11890 , \1735 );
not \U$11515 ( \11892 , \11890 );
and \U$11516 ( \11893 , \11892 , \1734 );
nor \U$11517 ( \11894 , \11891 , \11893 );
and \U$11518 ( \11895 , \11887 , \11894 );
and \U$11519 ( \11896 , \11879 , \11886 );
or \U$11520 ( \11897 , \11895 , \11896 );
not \U$11521 ( \11898 , \789 );
and \U$11522 ( \11899 , \883 , RIae781e8_105);
and \U$11523 ( \11900 , RIae785a8_113, \881 );
nor \U$11524 ( \11901 , \11899 , \11900 );
not \U$11525 ( \11902 , \11901 );
or \U$11526 ( \11903 , \11898 , \11902 );
or \U$11527 ( \11904 , \11901 , \787 );
nand \U$11528 ( \11905 , \11903 , \11904 );
and \U$11529 ( \11906 , \672 , RIae77f18_99);
and \U$11530 ( \11907 , RIae78008_101, \670 );
nor \U$11531 ( \11908 , \11906 , \11907 );
and \U$11532 ( \11909 , \11908 , \588 );
not \U$11533 ( \11910 , \11908 );
and \U$11534 ( \11911 , \11910 , \587 );
nor \U$11535 ( \11912 , \11909 , \11911 );
xor \U$11536 ( \11913 , \11905 , \11912 );
and \U$11537 ( \11914 , \1138 , RIae783c8_109);
and \U$11538 ( \11915 , RIae78530_112, \1136 );
nor \U$11539 ( \11916 , \11914 , \11915 );
and \U$11540 ( \11917 , \11916 , \1012 );
not \U$11541 ( \11918 , \11916 );
and \U$11542 ( \11919 , \11918 , \1142 );
nor \U$11543 ( \11920 , \11917 , \11919 );
and \U$11544 ( \11921 , \11913 , \11920 );
and \U$11545 ( \11922 , \11905 , \11912 );
or \U$11546 ( \11923 , \11921 , \11922 );
xor \U$11547 ( \11924 , \11897 , \11923 );
and \U$11548 ( \11925 , \514 , RIae771f8_71);
and \U$11549 ( \11926 , RIae772e8_73, \512 );
nor \U$11550 ( \11927 , \11925 , \11926 );
not \U$11551 ( \11928 , \11927 );
not \U$11552 ( \11929 , \471 );
and \U$11553 ( \11930 , \11928 , \11929 );
and \U$11554 ( \11931 , \11927 , \471 );
nor \U$11555 ( \11932 , \11930 , \11931 );
and \U$11556 ( \11933 , \558 , RIae782d8_107);
and \U$11557 ( \11934 , RIae780f8_103, \556 );
nor \U$11558 ( \11935 , \11933 , \11934 );
and \U$11559 ( \11936 , \11935 , \562 );
not \U$11560 ( \11937 , \11935 );
and \U$11561 ( \11938 , \11937 , \504 );
nor \U$11562 ( \11939 , \11936 , \11938 );
xor \U$11563 ( \11940 , \11932 , \11939 );
and \U$11564 ( \11941 , \436 , RIae77180_70);
and \U$11565 ( \11942 , RIae77018_67, \434 );
nor \U$11566 ( \11943 , \11941 , \11942 );
not \U$11567 ( \11944 , \11943 );
not \U$11568 ( \11945 , \400 );
and \U$11569 ( \11946 , \11944 , \11945 );
and \U$11570 ( \11947 , \11943 , \400 );
nor \U$11571 ( \11948 , \11946 , \11947 );
and \U$11572 ( \11949 , \11940 , \11948 );
and \U$11573 ( \11950 , \11932 , \11939 );
nor \U$11574 ( \11951 , \11949 , \11950 );
and \U$11575 ( \11952 , \11924 , \11951 );
and \U$11576 ( \11953 , \11897 , \11923 );
or \U$11577 ( \11954 , \11952 , \11953 );
and \U$11578 ( \11955 , \11872 , \11954 );
and \U$11579 ( \11956 , \11793 , \11871 );
or \U$11580 ( \11957 , \11955 , \11956 );
xor \U$11581 ( \11958 , \11710 , \11957 );
xor \U$11582 ( \11959 , \10932 , \10936 );
xor \U$11583 ( \11960 , \11959 , \10944 );
xor \U$11584 ( \11961 , \11297 , \11299 );
xor \U$11585 ( \11962 , \11961 , \11302 );
and \U$11586 ( \11963 , \11960 , \11962 );
xor \U$11587 ( \11964 , \11008 , \11015 );
xor \U$11588 ( \11965 , \11964 , \11023 );
xor \U$11589 ( \11966 , \11272 , \11277 );
xor \U$11590 ( \11967 , \11965 , \11966 );
xor \U$11591 ( \11968 , \11297 , \11299 );
xor \U$11592 ( \11969 , \11968 , \11302 );
and \U$11593 ( \11970 , \11967 , \11969 );
and \U$11594 ( \11971 , \11960 , \11967 );
or \U$11595 ( \11972 , \11963 , \11970 , \11971 );
and \U$11596 ( \11973 , \11958 , \11972 );
and \U$11597 ( \11974 , \11710 , \11957 );
or \U$11598 ( \11975 , \11973 , \11974 );
xor \U$11599 ( \11976 , \11672 , \11975 );
xor \U$11600 ( \11977 , \11393 , \11481 );
xor \U$11601 ( \11978 , \11977 , \11563 );
xor \U$11602 ( \11979 , \11282 , \11294 );
xor \U$11603 ( \11980 , \11979 , \11305 );
and \U$11604 ( \11981 , \11978 , \11980 );
xor \U$11605 ( \11982 , \10863 , \10865 );
xor \U$11606 ( \11983 , \11982 , \10868 );
xor \U$11607 ( \11984 , \11569 , \11576 );
xor \U$11608 ( \11985 , \11983 , \11984 );
xor \U$11609 ( \11986 , \11282 , \11294 );
xor \U$11610 ( \11987 , \11986 , \11305 );
and \U$11611 ( \11988 , \11985 , \11987 );
and \U$11612 ( \11989 , \11978 , \11985 );
or \U$11613 ( \11990 , \11981 , \11988 , \11989 );
and \U$11614 ( \11991 , \11976 , \11990 );
and \U$11615 ( \11992 , \11672 , \11975 );
or \U$11616 ( \11993 , \11991 , \11992 );
and \U$11617 ( \11994 , \11650 , \11993 );
and \U$11618 ( \11995 , \11632 , \11649 );
nor \U$11619 ( \11996 , \11994 , \11995 );
xor \U$11620 ( \11997 , \11230 , \11586 );
xor \U$11621 ( \11998 , \11997 , \11593 );
and \U$11622 ( \11999 , \11996 , \11998 );
and \U$11623 ( \12000 , \11619 , \11996 );
or \U$11624 ( \12001 , \11622 , \11999 , \12000 );
nor \U$11625 ( \12002 , \11613 , \12001 );
and \U$11626 ( \12003 , \11602 , \12002 );
xor \U$11627 ( \12004 , \12002 , \11602 );
not \U$11628 ( \12005 , \11267 );
xor \U$11629 ( \12006 , \11584 , \11260 );
not \U$11630 ( \12007 , \12006 );
or \U$11631 ( \12008 , \12005 , \12007 );
or \U$11632 ( \12009 , \12006 , \11267 );
nand \U$11633 ( \12010 , \12008 , \12009 );
not \U$11634 ( \12011 , \12010 );
xor \U$11635 ( \12012 , \11632 , \11649 );
xor \U$11636 ( \12013 , \12012 , \11993 );
not \U$11637 ( \12014 , \12013 );
or \U$11638 ( \12015 , \12011 , \12014 );
or \U$11639 ( \12016 , \12013 , \12010 );
xor \U$11640 ( \12017 , \11710 , \11957 );
xor \U$11641 ( \12018 , \12017 , \11972 );
xor \U$11642 ( \12019 , \11664 , \11666 );
xor \U$11643 ( \12020 , \12019 , \11669 );
and \U$11644 ( \12021 , \12018 , \12020 );
xor \U$11645 ( \12022 , \11282 , \11294 );
xor \U$11646 ( \12023 , \12022 , \11305 );
xor \U$11647 ( \12024 , \11978 , \11985 );
xor \U$11648 ( \12025 , \12023 , \12024 );
xor \U$11649 ( \12026 , \11664 , \11666 );
xor \U$11650 ( \12027 , \12026 , \11669 );
and \U$11651 ( \12028 , \12025 , \12027 );
and \U$11652 ( \12029 , \12018 , \12025 );
or \U$11653 ( \12030 , \12021 , \12028 , \12029 );
xor \U$11654 ( \12031 , \11897 , \11923 );
xor \U$11655 ( \12032 , \12031 , \11951 );
xor \U$11656 ( \12033 , \11818 , \11840 );
xor \U$11657 ( \12034 , \12033 , \11868 );
xor \U$11658 ( \12035 , \12032 , \12034 );
xor \U$11659 ( \12036 , \11735 , \11761 );
xor \U$11660 ( \12037 , \12036 , \11790 );
and \U$11661 ( \12038 , \12035 , \12037 );
and \U$11662 ( \12039 , \12032 , \12034 );
or \U$11663 ( \12040 , \12038 , \12039 );
xor \U$11664 ( \12041 , \11418 , \11443 );
xor \U$11665 ( \12042 , \12041 , \11478 );
xor \U$11666 ( \12043 , \12040 , \12042 );
or \U$11667 ( \12044 , \11695 , \11685 );
nand \U$11668 ( \12045 , \12044 , \11696 );
xor \U$11669 ( \12046 , \11699 , \11701 );
xor \U$11670 ( \12047 , \12046 , \11704 );
and \U$11671 ( \12048 , \12045 , \12047 );
xor \U$11672 ( \12049 , \11542 , \11549 );
xor \U$11673 ( \12050 , \12049 , \11557 );
xor \U$11674 ( \12051 , \11674 , \11679 );
xor \U$11675 ( \12052 , \12050 , \12051 );
xor \U$11676 ( \12053 , \11699 , \11701 );
xor \U$11677 ( \12054 , \12053 , \11704 );
and \U$11678 ( \12055 , \12052 , \12054 );
and \U$11679 ( \12056 , \12045 , \12052 );
or \U$11680 ( \12057 , \12048 , \12055 , \12056 );
and \U$11681 ( \12058 , \12043 , \12057 );
and \U$11682 ( \12059 , \12040 , \12042 );
or \U$11683 ( \12060 , \12058 , \12059 );
and \U$11684 ( \12061 , \3730 , RIae75e48_29);
and \U$11685 ( \12062 , RIae75c68_25, \3728 );
nor \U$11686 ( \12063 , \12061 , \12062 );
and \U$11687 ( \12064 , \12063 , \3422 );
not \U$11688 ( \12065 , \12063 );
and \U$11689 ( \12066 , \12065 , \3732 );
nor \U$11690 ( \12067 , \12064 , \12066 );
and \U$11691 ( \12068 , \4247 , RIae75d58_27);
and \U$11692 ( \12069 , RIae755d8_11, \4245 );
nor \U$11693 ( \12070 , \12068 , \12069 );
and \U$11694 ( \12071 , \12070 , \4251 );
not \U$11695 ( \12072 , \12070 );
and \U$11696 ( \12073 , \12072 , \3989 );
nor \U$11697 ( \12074 , \12071 , \12073 );
xor \U$11698 ( \12075 , \12067 , \12074 );
and \U$11699 ( \12076 , \3214 , RIae758a8_17);
and \U$11700 ( \12077 , RIae75f38_31, \3212 );
nor \U$11701 ( \12078 , \12076 , \12077 );
not \U$11702 ( \12079 , \12078 );
not \U$11703 ( \12080 , \3218 );
and \U$11704 ( \12081 , \12079 , \12080 );
and \U$11705 ( \12082 , \12078 , \3218 );
nor \U$11706 ( \12083 , \12081 , \12082 );
and \U$11707 ( \12084 , \12075 , \12083 );
and \U$11708 ( \12085 , \12067 , \12074 );
nor \U$11709 ( \12086 , \12084 , \12085 );
not \U$11710 ( \12087 , \3089 );
and \U$11711 ( \12088 , \2783 , RIae75a88_21);
and \U$11712 ( \12089 , RIae75998_19, \2781 );
nor \U$11713 ( \12090 , \12088 , \12089 );
not \U$11714 ( \12091 , \12090 );
or \U$11715 ( \12092 , \12087 , \12091 );
or \U$11716 ( \12093 , \12090 , \2789 );
nand \U$11717 ( \12094 , \12092 , \12093 );
and \U$11718 ( \12095 , \2224 , RIae78878_119);
and \U$11719 ( \12096 , RIae78788_117, \2222 );
nor \U$11720 ( \12097 , \12095 , \12096 );
and \U$11721 ( \12098 , \12097 , \2061 );
not \U$11722 ( \12099 , \12097 );
and \U$11723 ( \12100 , \12099 , \2060 );
nor \U$11724 ( \12101 , \12098 , \12100 );
xor \U$11725 ( \12102 , \12094 , \12101 );
and \U$11726 ( \12103 , \2607 , RIae78698_115);
and \U$11727 ( \12104 , RIae75b78_23, \2605 );
nor \U$11728 ( \12105 , \12103 , \12104 );
and \U$11729 ( \12106 , \12105 , \2611 );
not \U$11730 ( \12107 , \12105 );
and \U$11731 ( \12108 , \12107 , \2397 );
nor \U$11732 ( \12109 , \12106 , \12108 );
and \U$11733 ( \12110 , \12102 , \12109 );
and \U$11734 ( \12111 , \12094 , \12101 );
or \U$11735 ( \12112 , \12110 , \12111 );
xor \U$11736 ( \12113 , \12086 , \12112 );
and \U$11737 ( \12114 , \5399 , RIae756c8_13);
and \U$11738 ( \12115 , RIae75218_3, \5397 );
nor \U$11739 ( \12116 , \12114 , \12115 );
and \U$11740 ( \12117 , \12116 , \5403 );
not \U$11741 ( \12118 , \12116 );
and \U$11742 ( \12119 , \12118 , \5016 );
nor \U$11743 ( \12120 , \12117 , \12119 );
and \U$11744 ( \12121 , \5896 , RIae75128_1);
and \U$11745 ( \12122 , RIae75308_5, \5894 );
nor \U$11746 ( \12123 , \12121 , \12122 );
and \U$11747 ( \12124 , \12123 , \5589 );
not \U$11748 ( \12125 , \12123 );
and \U$11749 ( \12126 , \12125 , \5590 );
nor \U$11750 ( \12127 , \12124 , \12126 );
xor \U$11751 ( \12128 , \12120 , \12127 );
and \U$11752 ( \12129 , \4688 , RIae754e8_9);
and \U$11753 ( \12130 , RIae757b8_15, \4686 );
nor \U$11754 ( \12131 , \12129 , \12130 );
and \U$11755 ( \12132 , \12131 , \4482 );
not \U$11756 ( \12133 , \12131 );
and \U$11757 ( \12134 , \12133 , \4481 );
nor \U$11758 ( \12135 , \12132 , \12134 );
and \U$11759 ( \12136 , \12128 , \12135 );
and \U$11760 ( \12137 , \12120 , \12127 );
nor \U$11761 ( \12138 , \12136 , \12137 );
and \U$11762 ( \12139 , \12113 , \12138 );
and \U$11763 ( \12140 , \12086 , \12112 );
nor \U$11764 ( \12141 , \12139 , \12140 );
and \U$11765 ( \12142 , \6941 , RIae764d8_43);
and \U$11766 ( \12143 , RIae766b8_47, \6939 );
nor \U$11767 ( \12144 , \12142 , \12143 );
and \U$11768 ( \12145 , \12144 , \6314 );
not \U$11769 ( \12146 , \12144 );
and \U$11770 ( \12147 , \12146 , \6945 );
nor \U$11771 ( \12148 , \12145 , \12147 );
and \U$11772 ( \12149 , \7633 , RIae765c8_45);
and \U$11773 ( \12150 , RIae76118_35, \7631 );
nor \U$11774 ( \12151 , \12149 , \12150 );
and \U$11775 ( \12152 , \12151 , \7206 );
not \U$11776 ( \12153 , \12151 );
and \U$11777 ( \12154 , \12153 , \7205 );
nor \U$11778 ( \12155 , \12152 , \12154 );
xor \U$11779 ( \12156 , \12148 , \12155 );
and \U$11780 ( \12157 , \6172 , RIae753f8_7);
and \U$11781 ( \12158 , RIae763e8_41, \6170 );
nor \U$11782 ( \12159 , \12157 , \12158 );
and \U$11783 ( \12160 , \12159 , \6176 );
not \U$11784 ( \12161 , \12159 );
and \U$11785 ( \12162 , \12161 , \6175 );
nor \U$11786 ( \12163 , \12160 , \12162 );
and \U$11787 ( \12164 , \12156 , \12163 );
and \U$11788 ( \12165 , \12148 , \12155 );
nor \U$11789 ( \12166 , \12164 , \12165 );
and \U$11790 ( \12167 , \10548 , RIae76898_51);
and \U$11791 ( \12168 , RIae76b68_57, \10546 );
nor \U$11792 ( \12169 , \12167 , \12168 );
and \U$11793 ( \12170 , \12169 , \10118 );
not \U$11794 ( \12171 , \12169 );
and \U$11795 ( \12172 , \12171 , \10421 );
nor \U$11796 ( \12173 , \12170 , \12172 );
and \U$11797 ( \12174 , RIae7a060_170, RIae7a948_189);
not \U$11798 ( \12175 , RIae7a7e0_186);
and \U$11799 ( \12176 , \12175 , RIae7a948_189);
nor \U$11800 ( \12177 , \12175 , RIae7a948_189);
or \U$11801 ( \12178 , \12176 , \12177 );
nor \U$11802 ( \12179 , RIae7a060_170, RIae7a948_189);
nor \U$11803 ( \12180 , \12174 , \12178 , \12179 );
nand \U$11804 ( \12181 , RIae78da0_130, \12180 );
and \U$11805 ( \12182 , \12181 , \11827 );
not \U$11806 ( \12183 , \12181 );
not \U$11807 ( \12184 , \11827 );
and \U$11808 ( \12185 , \12183 , \12184 );
nor \U$11809 ( \12186 , \12182 , \12185 );
xor \U$11810 ( \12187 , \12173 , \12186 );
and \U$11811 ( \12188 , \11470 , RIae78a58_123);
and \U$11812 ( \12189 , RIae78cb0_128, \11468 );
nor \U$11813 ( \12190 , \12188 , \12189 );
and \U$11814 ( \12191 , \12190 , \11474 );
not \U$11815 ( \12192 , \12190 );
and \U$11816 ( \12193 , \12192 , \10936 );
nor \U$11817 ( \12194 , \12191 , \12193 );
and \U$11818 ( \12195 , \12187 , \12194 );
and \U$11819 ( \12196 , \12173 , \12186 );
or \U$11820 ( \12197 , \12195 , \12196 );
xor \U$11821 ( \12198 , \12166 , \12197 );
and \U$11822 ( \12199 , \8371 , RIae76028_33);
and \U$11823 ( \12200 , RIae762f8_39, \8369 );
nor \U$11824 ( \12201 , \12199 , \12200 );
and \U$11825 ( \12202 , \12201 , \8019 );
not \U$11826 ( \12203 , \12201 );
and \U$11827 ( \12204 , \12203 , \8020 );
nor \U$11828 ( \12205 , \12202 , \12204 );
and \U$11829 ( \12206 , \8966 , RIae76208_37);
and \U$11830 ( \12207 , RIae76a78_55, \8964 );
nor \U$11831 ( \12208 , \12206 , \12207 );
and \U$11832 ( \12209 , \12208 , \8789 );
not \U$11833 ( \12210 , \12208 );
and \U$11834 ( \12211 , \12210 , \8799 );
nor \U$11835 ( \12212 , \12209 , \12211 );
xor \U$11836 ( \12213 , \12205 , \12212 );
and \U$11837 ( \12214 , \9760 , RIae76988_53);
and \U$11838 ( \12215 , RIae767a8_49, \9758 );
nor \U$11839 ( \12216 , \12214 , \12215 );
and \U$11840 ( \12217 , \12216 , \9272 );
not \U$11841 ( \12218 , \12216 );
and \U$11842 ( \12219 , \12218 , \9273 );
nor \U$11843 ( \12220 , \12217 , \12219 );
and \U$11844 ( \12221 , \12213 , \12220 );
and \U$11845 ( \12222 , \12205 , \12212 );
or \U$11846 ( \12223 , \12221 , \12222 );
and \U$11847 ( \12224 , \12198 , \12223 );
and \U$11848 ( \12225 , \12166 , \12197 );
or \U$11849 ( \12226 , \12224 , \12225 );
or \U$11850 ( \12227 , \12141 , \12226 );
not \U$11851 ( \12228 , \12141 );
not \U$11852 ( \12229 , \12226 );
or \U$11853 ( \12230 , \12228 , \12229 );
not \U$11854 ( \12231 , \789 );
and \U$11855 ( \12232 , \883 , RIae78008_101);
and \U$11856 ( \12233 , RIae781e8_105, \881 );
nor \U$11857 ( \12234 , \12232 , \12233 );
not \U$11858 ( \12235 , \12234 );
or \U$11859 ( \12236 , \12231 , \12235 );
or \U$11860 ( \12237 , \12234 , \789 );
nand \U$11861 ( \12238 , \12236 , \12237 );
and \U$11862 ( \12239 , \1138 , RIae785a8_113);
and \U$11863 ( \12240 , RIae783c8_109, \1136 );
nor \U$11864 ( \12241 , \12239 , \12240 );
and \U$11865 ( \12242 , \12241 , \1012 );
not \U$11866 ( \12243 , \12241 );
and \U$11867 ( \12244 , \12243 , \1142 );
nor \U$11868 ( \12245 , \12242 , \12244 );
xor \U$11869 ( \12246 , \12238 , \12245 );
and \U$11870 ( \12247 , \672 , RIae780f8_103);
and \U$11871 ( \12248 , RIae77f18_99, \670 );
nor \U$11872 ( \12249 , \12247 , \12248 );
and \U$11873 ( \12250 , \12249 , \588 );
not \U$11874 ( \12251 , \12249 );
and \U$11875 ( \12252 , \12251 , \587 );
nor \U$11876 ( \12253 , \12250 , \12252 );
and \U$11877 ( \12254 , \12246 , \12253 );
and \U$11878 ( \12255 , \12238 , \12245 );
nor \U$11879 ( \12256 , \12254 , \12255 );
and \U$11880 ( \12257 , \1593 , RIae77b58_91);
and \U$11881 ( \12258 , RIae77d38_95, \1591 );
nor \U$11882 ( \12259 , \12257 , \12258 );
and \U$11883 ( \12260 , \12259 , \1498 );
not \U$11884 ( \12261 , \12259 );
and \U$11885 ( \12262 , \12261 , \1488 );
nor \U$11886 ( \12263 , \12260 , \12262 );
and \U$11887 ( \12264 , \1939 , RIae77e28_97);
and \U$11888 ( \12265 , RIae78968_121, \1937 );
nor \U$11889 ( \12266 , \12264 , \12265 );
and \U$11890 ( \12267 , \12266 , \1735 );
not \U$11891 ( \12268 , \12266 );
and \U$11892 ( \12269 , \12268 , \1734 );
nor \U$11893 ( \12270 , \12267 , \12269 );
xor \U$11894 ( \12271 , \12263 , \12270 );
and \U$11895 ( \12272 , \1376 , RIae78530_112);
and \U$11896 ( \12273 , RIae77c48_93, \1374 );
nor \U$11897 ( \12274 , \12272 , \12273 );
and \U$11898 ( \12275 , \12274 , \1380 );
not \U$11899 ( \12276 , \12274 );
and \U$11900 ( \12277 , \12276 , \1261 );
nor \U$11901 ( \12278 , \12275 , \12277 );
and \U$11902 ( \12279 , \12271 , \12278 );
and \U$11903 ( \12280 , \12263 , \12270 );
nor \U$11904 ( \12281 , \12279 , \12280 );
xor \U$11905 ( \12282 , \12256 , \12281 );
and \U$11906 ( \12283 , \436 , RIae76c58_59);
and \U$11907 ( \12284 , RIae77180_70, \434 );
nor \U$11908 ( \12285 , \12283 , \12284 );
not \U$11909 ( \12286 , \12285 );
not \U$11910 ( \12287 , \402 );
and \U$11911 ( \12288 , \12286 , \12287 );
and \U$11912 ( \12289 , \12285 , \400 );
nor \U$11913 ( \12290 , \12288 , \12289 );
not \U$11914 ( \12291 , \12290 );
and \U$11915 ( \12292 , \558 , RIae772e8_73);
and \U$11916 ( \12293 , RIae782d8_107, \556 );
nor \U$11917 ( \12294 , \12292 , \12293 );
and \U$11918 ( \12295 , \12294 , \562 );
not \U$11919 ( \12296 , \12294 );
and \U$11920 ( \12297 , \12296 , \504 );
nor \U$11921 ( \12298 , \12295 , \12297 );
not \U$11922 ( \12299 , \12298 );
and \U$11923 ( \12300 , \12291 , \12299 );
and \U$11924 ( \12301 , \12298 , \12290 );
and \U$11925 ( \12302 , \514 , RIae77018_67);
and \U$11926 ( \12303 , RIae771f8_71, \512 );
nor \U$11927 ( \12304 , \12302 , \12303 );
not \U$11928 ( \12305 , \12304 );
not \U$11929 ( \12306 , \471 );
and \U$11930 ( \12307 , \12305 , \12306 );
and \U$11931 ( \12308 , \12304 , \471 );
nor \U$11932 ( \12309 , \12307 , \12308 );
nor \U$11933 ( \12310 , \12301 , \12309 );
nor \U$11934 ( \12311 , \12300 , \12310 );
and \U$11935 ( \12312 , \12282 , \12311 );
and \U$11936 ( \12313 , \12256 , \12281 );
nor \U$11937 ( \12314 , \12312 , \12313 );
nand \U$11938 ( \12315 , \12230 , \12314 );
nand \U$11939 ( \12316 , \12227 , \12315 );
xor \U$11940 ( \12317 , \11800 , \11807 );
xor \U$11941 ( \12318 , \12317 , \11815 );
not \U$11942 ( \12319 , \12318 );
not \U$11943 ( \12320 , \11855 );
not \U$11944 ( \12321 , \11866 );
or \U$11945 ( \12322 , \12320 , \12321 );
or \U$11946 ( \12323 , \11855 , \11866 );
nand \U$11947 ( \12324 , \12322 , \12323 );
not \U$11948 ( \12325 , \12324 );
not \U$11949 ( \12326 , \11848 );
and \U$11950 ( \12327 , \12325 , \12326 );
and \U$11951 ( \12328 , \12324 , \11848 );
nor \U$11952 ( \12329 , \12327 , \12328 );
not \U$11953 ( \12330 , \12329 );
and \U$11954 ( \12331 , \12319 , \12330 );
and \U$11955 ( \12332 , \12329 , \12318 );
and \U$11956 ( \12333 , \11838 , \12184 );
not \U$11957 ( \12334 , \11838 );
and \U$11958 ( \12335 , \12334 , \11827 );
nor \U$11959 ( \12336 , \12333 , \12335 );
not \U$11960 ( \12337 , \12336 );
not \U$11961 ( \12338 , \11825 );
and \U$11962 ( \12339 , \12337 , \12338 );
and \U$11963 ( \12340 , \12336 , \11825 );
nor \U$11964 ( \12341 , \12339 , \12340 );
nor \U$11965 ( \12342 , \12332 , \12341 );
nor \U$11966 ( \12343 , \12331 , \12342 );
not \U$11967 ( \12344 , \11476 );
not \U$11968 ( \12345 , \11458 );
or \U$11969 ( \12346 , \12344 , \12345 );
or \U$11970 ( \12347 , \11458 , \11476 );
nand \U$11971 ( \12348 , \12346 , \12347 );
not \U$11972 ( \12349 , \12348 );
not \U$11973 ( \12350 , \11451 );
and \U$11974 ( \12351 , \12349 , \12350 );
and \U$11975 ( \12352 , \12348 , \11451 );
nor \U$11976 ( \12353 , \12351 , \12352 );
not \U$11977 ( \12354 , \12353 );
xor \U$11978 ( \12355 , \11400 , \11407 );
xor \U$11979 ( \12356 , \12355 , \11415 );
nor \U$11980 ( \12357 , \12354 , \12356 );
or \U$11981 ( \12358 , \12343 , \12357 );
not \U$11982 ( \12359 , \12353 );
nand \U$11983 ( \12360 , \12359 , \12356 );
nand \U$11984 ( \12361 , \12358 , \12360 );
xor \U$11985 ( \12362 , \12316 , \12361 );
and \U$11986 ( \12363 , \384 , RIae76d48_61);
and \U$11987 ( \12364 , RIae76c58_59, \382 );
nor \U$11988 ( \12365 , \12363 , \12364 );
not \U$11989 ( \12366 , \12365 );
not \U$11990 ( \12367 , \392 );
and \U$11991 ( \12368 , \12366 , \12367 );
and \U$11992 ( \12369 , \12365 , \388 );
nor \U$11993 ( \12370 , \12368 , \12369 );
nand \U$11994 ( \12371 , RIae76e38_63, RIae78b48_125);
xor \U$11995 ( \12372 , \12370 , \12371 );
nand \U$11996 ( \12373 , RIae76f28_65, RIae78b48_125);
and \U$11997 ( \12374 , \384 , RIae76e38_63);
and \U$11998 ( \12375 , RIae76d48_61, \382 );
nor \U$11999 ( \12376 , \12374 , \12375 );
not \U$12000 ( \12377 , \12376 );
not \U$12001 ( \12378 , \388 );
and \U$12002 ( \12379 , \12377 , \12378 );
and \U$12003 ( \12380 , \12376 , \388 );
nor \U$12004 ( \12381 , \12379 , \12380 );
nand \U$12005 ( \12382 , \12373 , \12381 );
not \U$12006 ( \12383 , \12382 );
and \U$12007 ( \12384 , \12372 , \12383 );
and \U$12008 ( \12385 , \12370 , \12371 );
or \U$12009 ( \12386 , \12384 , \12385 );
xor \U$12010 ( \12387 , \11879 , \11886 );
xor \U$12011 ( \12388 , \12387 , \11894 );
xor \U$12012 ( \12389 , \11905 , \11912 );
xor \U$12013 ( \12390 , \12389 , \11920 );
and \U$12014 ( \12391 , \12388 , \12390 );
not \U$12015 ( \12392 , \12390 );
not \U$12016 ( \12393 , \12388 );
and \U$12017 ( \12394 , \12392 , \12393 );
xor \U$12018 ( \12395 , \11932 , \11939 );
xor \U$12019 ( \12396 , \12395 , \11948 );
nor \U$12020 ( \12397 , \12394 , \12396 );
nor \U$12021 ( \12398 , \12391 , \12397 );
xor \U$12022 ( \12399 , \12386 , \12398 );
xor \U$12023 ( \12400 , \11742 , \11750 );
xor \U$12024 ( \12401 , \12400 , \11758 );
not \U$12025 ( \12402 , \12401 );
not \U$12026 ( \12403 , \11777 );
not \U$12027 ( \12404 , \11788 );
or \U$12028 ( \12405 , \12403 , \12404 );
or \U$12029 ( \12406 , \11777 , \11788 );
nand \U$12030 ( \12407 , \12405 , \12406 );
not \U$12031 ( \12408 , \12407 );
not \U$12032 ( \12409 , \11770 );
and \U$12033 ( \12410 , \12408 , \12409 );
and \U$12034 ( \12411 , \12407 , \11770 );
nor \U$12035 ( \12412 , \12410 , \12411 );
not \U$12036 ( \12413 , \12412 );
and \U$12037 ( \12414 , \12402 , \12413 );
and \U$12038 ( \12415 , \12412 , \12401 );
xor \U$12039 ( \12416 , \11717 , \11724 );
xor \U$12040 ( \12417 , \12416 , \11732 );
nor \U$12041 ( \12418 , \12415 , \12417 );
nor \U$12042 ( \12419 , \12414 , \12418 );
and \U$12043 ( \12420 , \12399 , \12419 );
and \U$12044 ( \12421 , \12386 , \12398 );
nor \U$12045 ( \12422 , \12420 , \12421 );
and \U$12046 ( \12423 , \12362 , \12422 );
and \U$12047 ( \12424 , \12316 , \12361 );
or \U$12048 ( \12425 , \12423 , \12424 );
xor \U$12049 ( \12426 , \12060 , \12425 );
xor \U$12050 ( \12427 , \11509 , \11534 );
xor \U$12051 ( \12428 , \12427 , \11560 );
xor \U$12052 ( \12429 , \11652 , \11659 );
xor \U$12053 ( \12430 , \12428 , \12429 );
xor \U$12054 ( \12431 , \11684 , \11696 );
xor \U$12055 ( \12432 , \12431 , \11707 );
and \U$12056 ( \12433 , \12430 , \12432 );
xor \U$12057 ( \12434 , \11297 , \11299 );
xor \U$12058 ( \12435 , \12434 , \11302 );
xor \U$12059 ( \12436 , \11960 , \11967 );
xor \U$12060 ( \12437 , \12435 , \12436 );
xor \U$12061 ( \12438 , \11684 , \11696 );
xor \U$12062 ( \12439 , \12438 , \11707 );
and \U$12063 ( \12440 , \12437 , \12439 );
and \U$12064 ( \12441 , \12430 , \12437 );
or \U$12065 ( \12442 , \12433 , \12440 , \12441 );
and \U$12066 ( \12443 , \12426 , \12442 );
and \U$12067 ( \12444 , \12060 , \12425 );
or \U$12068 ( \12445 , \12443 , \12444 );
xor \U$12069 ( \12446 , \12030 , \12445 );
xor \U$12070 ( \12447 , \11634 , \11639 );
xor \U$12071 ( \12448 , \12447 , \11646 );
and \U$12072 ( \12449 , \12446 , \12448 );
and \U$12073 ( \12450 , \12030 , \12445 );
or \U$12074 ( \12451 , \12449 , \12450 );
nand \U$12075 ( \12452 , \12016 , \12451 );
nand \U$12076 ( \12453 , \12015 , \12452 );
not \U$12077 ( \12454 , \12453 );
xor \U$12078 ( \12455 , \11230 , \11586 );
xor \U$12079 ( \12456 , \12455 , \11593 );
xor \U$12080 ( \12457 , \11619 , \11996 );
xor \U$12081 ( \12458 , \12456 , \12457 );
not \U$12082 ( \12459 , \12458 );
or \U$12083 ( \12460 , \12454 , \12459 );
or \U$12084 ( \12461 , \12458 , \12453 );
nand \U$12085 ( \12462 , \12460 , \12461 );
xor \U$12086 ( \12463 , \11672 , \11975 );
xor \U$12087 ( \12464 , \12463 , \11990 );
xor \U$12088 ( \12465 , \12030 , \12445 );
xor \U$12089 ( \12466 , \12465 , \12448 );
and \U$12090 ( \12467 , \12464 , \12466 );
xor \U$12091 ( \12468 , \11793 , \11871 );
xor \U$12092 ( \12469 , \12468 , \11954 );
xor \U$12093 ( \12470 , \12040 , \12042 );
xor \U$12094 ( \12471 , \12470 , \12057 );
and \U$12095 ( \12472 , \12469 , \12471 );
xor \U$12096 ( \12473 , \11684 , \11696 );
xor \U$12097 ( \12474 , \12473 , \11707 );
xor \U$12098 ( \12475 , \12430 , \12437 );
xor \U$12099 ( \12476 , \12474 , \12475 );
xor \U$12100 ( \12477 , \12040 , \12042 );
xor \U$12101 ( \12478 , \12477 , \12057 );
and \U$12102 ( \12479 , \12476 , \12478 );
and \U$12103 ( \12480 , \12469 , \12476 );
or \U$12104 ( \12481 , \12472 , \12479 , \12480 );
xor \U$12105 ( \12482 , \12256 , \12281 );
xor \U$12106 ( \12483 , \12482 , \12311 );
xor \U$12107 ( \12484 , \12370 , \12371 );
xor \U$12108 ( \12485 , \12484 , \12383 );
or \U$12109 ( \12486 , \12483 , \12485 );
not \U$12110 ( \12487 , \12485 );
not \U$12111 ( \12488 , \12483 );
or \U$12112 ( \12489 , \12487 , \12488 );
xor \U$12113 ( \12490 , \12086 , \12112 );
xor \U$12114 ( \12491 , \12490 , \12138 );
nand \U$12115 ( \12492 , \12489 , \12491 );
nand \U$12116 ( \12493 , \12486 , \12492 );
xor \U$12117 ( \12494 , \12032 , \12034 );
xor \U$12118 ( \12495 , \12494 , \12037 );
and \U$12119 ( \12496 , \12493 , \12495 );
xor \U$12120 ( \12497 , \11699 , \11701 );
xor \U$12121 ( \12498 , \12497 , \11704 );
xor \U$12122 ( \12499 , \12045 , \12052 );
xor \U$12123 ( \12500 , \12498 , \12499 );
xor \U$12124 ( \12501 , \12032 , \12034 );
xor \U$12125 ( \12502 , \12501 , \12037 );
and \U$12126 ( \12503 , \12500 , \12502 );
and \U$12127 ( \12504 , \12493 , \12500 );
or \U$12128 ( \12505 , \12496 , \12503 , \12504 );
not \U$12129 ( \12506 , \12505 );
not \U$12130 ( \12507 , \12356 );
not \U$12131 ( \12508 , \12343 );
or \U$12132 ( \12509 , \12507 , \12508 );
or \U$12133 ( \12510 , \12343 , \12356 );
nand \U$12134 ( \12511 , \12509 , \12510 );
not \U$12135 ( \12512 , \12511 );
not \U$12136 ( \12513 , \12353 );
and \U$12137 ( \12514 , \12512 , \12513 );
and \U$12138 ( \12515 , \12511 , \12353 );
nor \U$12139 ( \12516 , \12514 , \12515 );
not \U$12140 ( \12517 , \12516 );
not \U$12141 ( \12518 , \12141 );
not \U$12142 ( \12519 , \12314 );
or \U$12143 ( \12520 , \12518 , \12519 );
or \U$12144 ( \12521 , \12314 , \12141 );
nand \U$12145 ( \12522 , \12520 , \12521 );
not \U$12146 ( \12523 , \12522 );
not \U$12147 ( \12524 , \12226 );
and \U$12148 ( \12525 , \12523 , \12524 );
and \U$12149 ( \12526 , \12522 , \12226 );
nor \U$12150 ( \12527 , \12525 , \12526 );
not \U$12151 ( \12528 , \12527 );
and \U$12152 ( \12529 , \12517 , \12528 );
and \U$12153 ( \12530 , \12516 , \12527 );
xor \U$12154 ( \12531 , \12386 , \12398 );
xor \U$12155 ( \12532 , \12531 , \12419 );
nor \U$12156 ( \12533 , \12530 , \12532 );
nor \U$12157 ( \12534 , \12529 , \12533 );
or \U$12158 ( \12535 , \12506 , \12534 );
not \U$12159 ( \12536 , \12534 );
not \U$12160 ( \12537 , \12506 );
or \U$12161 ( \12538 , \12536 , \12537 );
xor \U$12162 ( \12539 , \12238 , \12245 );
xor \U$12163 ( \12540 , \12539 , \12253 );
xor \U$12164 ( \12541 , \12094 , \12101 );
xor \U$12165 ( \12542 , \12541 , \12109 );
and \U$12166 ( \12543 , \12540 , \12542 );
xor \U$12167 ( \12544 , \12263 , \12270 );
xor \U$12168 ( \12545 , \12544 , \12278 );
xor \U$12169 ( \12546 , \12094 , \12101 );
xor \U$12170 ( \12547 , \12546 , \12109 );
and \U$12171 ( \12548 , \12545 , \12547 );
and \U$12172 ( \12549 , \12540 , \12545 );
or \U$12173 ( \12550 , \12543 , \12548 , \12549 );
and \U$12174 ( \12551 , \384 , RIae76f28_65);
and \U$12175 ( \12552 , RIae76e38_63, \382 );
nor \U$12176 ( \12553 , \12551 , \12552 );
not \U$12177 ( \12554 , \12553 );
not \U$12178 ( \12555 , \388 );
and \U$12179 ( \12556 , \12554 , \12555 );
and \U$12180 ( \12557 , \12553 , \388 );
nor \U$12181 ( \12558 , \12556 , \12557 );
nand \U$12182 ( \12559 , RIae77888_85, RIae78b48_125);
or \U$12183 ( \12560 , \12558 , \12559 );
not \U$12184 ( \12561 , \12559 );
not \U$12185 ( \12562 , \12558 );
or \U$12186 ( \12563 , \12561 , \12562 );
not \U$12187 ( \12564 , \400 );
and \U$12188 ( \12565 , \436 , RIae76d48_61);
and \U$12189 ( \12566 , RIae76c58_59, \434 );
nor \U$12190 ( \12567 , \12565 , \12566 );
not \U$12191 ( \12568 , \12567 );
or \U$12192 ( \12569 , \12564 , \12568 );
or \U$12193 ( \12570 , \12567 , \400 );
nand \U$12194 ( \12571 , \12569 , \12570 );
nand \U$12195 ( \12572 , \12563 , \12571 );
nand \U$12196 ( \12573 , \12560 , \12572 );
or \U$12197 ( \12574 , \12381 , \12373 );
nand \U$12198 ( \12575 , \12574 , \12382 );
xor \U$12199 ( \12576 , \12573 , \12575 );
not \U$12200 ( \12577 , \12290 );
xor \U$12201 ( \12578 , \12309 , \12298 );
not \U$12202 ( \12579 , \12578 );
or \U$12203 ( \12580 , \12577 , \12579 );
or \U$12204 ( \12581 , \12578 , \12290 );
nand \U$12205 ( \12582 , \12580 , \12581 );
and \U$12206 ( \12583 , \12576 , \12582 );
and \U$12207 ( \12584 , \12573 , \12575 );
or \U$12208 ( \12585 , \12583 , \12584 );
xor \U$12209 ( \12586 , \12550 , \12585 );
xor \U$12210 ( \12587 , \12067 , \12074 );
xor \U$12211 ( \12588 , \12587 , \12083 );
xor \U$12212 ( \12589 , \12120 , \12127 );
xor \U$12213 ( \12590 , \12589 , \12135 );
or \U$12214 ( \12591 , \12588 , \12590 );
not \U$12215 ( \12592 , \12590 );
not \U$12216 ( \12593 , \12588 );
or \U$12217 ( \12594 , \12592 , \12593 );
xor \U$12218 ( \12595 , \12148 , \12155 );
xor \U$12219 ( \12596 , \12595 , \12163 );
nand \U$12220 ( \12597 , \12594 , \12596 );
nand \U$12221 ( \12598 , \12591 , \12597 );
and \U$12222 ( \12599 , \12586 , \12598 );
and \U$12223 ( \12600 , \12550 , \12585 );
or \U$12224 ( \12601 , \12599 , \12600 );
and \U$12225 ( \12602 , \1593 , RIae77c48_93);
and \U$12226 ( \12603 , RIae77b58_91, \1591 );
nor \U$12227 ( \12604 , \12602 , \12603 );
and \U$12228 ( \12605 , \12604 , \1488 );
not \U$12229 ( \12606 , \12604 );
and \U$12230 ( \12607 , \12606 , \1498 );
nor \U$12231 ( \12608 , \12605 , \12607 );
and \U$12232 ( \12609 , \2224 , RIae78968_121);
and \U$12233 ( \12610 , RIae78878_119, \2222 );
nor \U$12234 ( \12611 , \12609 , \12610 );
and \U$12235 ( \12612 , \12611 , \2060 );
not \U$12236 ( \12613 , \12611 );
and \U$12237 ( \12614 , \12613 , \2061 );
nor \U$12238 ( \12615 , \12612 , \12614 );
or \U$12239 ( \12616 , \12608 , \12615 );
not \U$12240 ( \12617 , \12615 );
not \U$12241 ( \12618 , \12608 );
or \U$12242 ( \12619 , \12617 , \12618 );
and \U$12243 ( \12620 , \1939 , RIae77d38_95);
and \U$12244 ( \12621 , RIae77e28_97, \1937 );
nor \U$12245 ( \12622 , \12620 , \12621 );
and \U$12246 ( \12623 , \12622 , \1735 );
not \U$12247 ( \12624 , \12622 );
and \U$12248 ( \12625 , \12624 , \1734 );
nor \U$12249 ( \12626 , \12623 , \12625 );
nand \U$12250 ( \12627 , \12619 , \12626 );
nand \U$12251 ( \12628 , \12616 , \12627 );
and \U$12252 ( \12629 , \1138 , RIae781e8_105);
and \U$12253 ( \12630 , RIae785a8_113, \1136 );
nor \U$12254 ( \12631 , \12629 , \12630 );
and \U$12255 ( \12632 , \12631 , \1142 );
not \U$12256 ( \12633 , \12631 );
and \U$12257 ( \12634 , \12633 , \1012 );
nor \U$12258 ( \12635 , \12632 , \12634 );
and \U$12259 ( \12636 , \1376 , RIae783c8_109);
and \U$12260 ( \12637 , RIae78530_112, \1374 );
nor \U$12261 ( \12638 , \12636 , \12637 );
and \U$12262 ( \12639 , \12638 , \1261 );
not \U$12263 ( \12640 , \12638 );
and \U$12264 ( \12641 , \12640 , \1380 );
nor \U$12265 ( \12642 , \12639 , \12641 );
xor \U$12266 ( \12643 , \12635 , \12642 );
and \U$12267 ( \12644 , \883 , RIae77f18_99);
and \U$12268 ( \12645 , RIae78008_101, \881 );
nor \U$12269 ( \12646 , \12644 , \12645 );
not \U$12270 ( \12647 , \12646 );
not \U$12271 ( \12648 , \789 );
and \U$12272 ( \12649 , \12647 , \12648 );
and \U$12273 ( \12650 , \12646 , \789 );
nor \U$12274 ( \12651 , \12649 , \12650 );
and \U$12275 ( \12652 , \12643 , \12651 );
and \U$12276 ( \12653 , \12635 , \12642 );
nor \U$12277 ( \12654 , \12652 , \12653 );
xor \U$12278 ( \12655 , \12628 , \12654 );
and \U$12279 ( \12656 , \558 , RIae771f8_71);
and \U$12280 ( \12657 , RIae772e8_73, \556 );
nor \U$12281 ( \12658 , \12656 , \12657 );
and \U$12282 ( \12659 , \12658 , \562 );
not \U$12283 ( \12660 , \12658 );
and \U$12284 ( \12661 , \12660 , \504 );
nor \U$12285 ( \12662 , \12659 , \12661 );
and \U$12286 ( \12663 , \672 , RIae782d8_107);
and \U$12287 ( \12664 , RIae780f8_103, \670 );
nor \U$12288 ( \12665 , \12663 , \12664 );
and \U$12289 ( \12666 , \12665 , \587 );
not \U$12290 ( \12667 , \12665 );
and \U$12291 ( \12668 , \12667 , \588 );
nor \U$12292 ( \12669 , \12666 , \12668 );
xor \U$12293 ( \12670 , \12662 , \12669 );
and \U$12294 ( \12671 , \514 , RIae77180_70);
and \U$12295 ( \12672 , RIae77018_67, \512 );
nor \U$12296 ( \12673 , \12671 , \12672 );
not \U$12297 ( \12674 , \12673 );
not \U$12298 ( \12675 , \471 );
and \U$12299 ( \12676 , \12674 , \12675 );
and \U$12300 ( \12677 , \12673 , \469 );
nor \U$12301 ( \12678 , \12676 , \12677 );
and \U$12302 ( \12679 , \12670 , \12678 );
and \U$12303 ( \12680 , \12662 , \12669 );
nor \U$12304 ( \12681 , \12679 , \12680 );
and \U$12305 ( \12682 , \12655 , \12681 );
and \U$12306 ( \12683 , \12628 , \12654 );
or \U$12307 ( \12684 , \12682 , \12683 );
and \U$12308 ( \12685 , \6941 , RIae763e8_41);
and \U$12309 ( \12686 , RIae764d8_43, \6939 );
nor \U$12310 ( \12687 , \12685 , \12686 );
and \U$12311 ( \12688 , \12687 , \6945 );
not \U$12312 ( \12689 , \12687 );
and \U$12313 ( \12690 , \12689 , \6314 );
nor \U$12314 ( \12691 , \12688 , \12690 );
and \U$12315 ( \12692 , \7633 , RIae766b8_47);
and \U$12316 ( \12693 , RIae765c8_45, \7631 );
nor \U$12317 ( \12694 , \12692 , \12693 );
and \U$12318 ( \12695 , \12694 , \7205 );
not \U$12319 ( \12696 , \12694 );
and \U$12320 ( \12697 , \12696 , \7206 );
nor \U$12321 ( \12698 , \12695 , \12697 );
xor \U$12322 ( \12699 , \12691 , \12698 );
and \U$12323 ( \12700 , \8371 , RIae76118_35);
and \U$12324 ( \12701 , RIae76028_33, \8369 );
nor \U$12325 ( \12702 , \12700 , \12701 );
and \U$12326 ( \12703 , \12702 , \8019 );
not \U$12327 ( \12704 , \12702 );
and \U$12328 ( \12705 , \12704 , \8020 );
nor \U$12329 ( \12706 , \12703 , \12705 );
and \U$12330 ( \12707 , \12699 , \12706 );
and \U$12331 ( \12708 , \12691 , \12698 );
or \U$12332 ( \12709 , \12707 , \12708 );
and \U$12333 ( \12710 , \11470 , RIae76b68_57);
and \U$12334 ( \12711 , RIae78a58_123, \11468 );
nor \U$12335 ( \12712 , \12710 , \12711 );
and \U$12336 ( \12713 , \12712 , \11474 );
not \U$12337 ( \12714 , \12712 );
and \U$12338 ( \12715 , \12714 , \10936 );
nor \U$12339 ( \12716 , \12713 , \12715 );
nand \U$12340 ( \12717 , RIae7a6f0_184, RIae7a768_185);
and \U$12341 ( \12718 , \12717 , RIae7a7e0_186);
xor \U$12342 ( \12719 , \12716 , \12718 );
and \U$12343 ( \12720 , \12180 , RIae78cb0_128);
and \U$12344 ( \12721 , RIae78da0_130, \12178 );
nor \U$12345 ( \12722 , \12720 , \12721 );
and \U$12346 ( \12723 , \12722 , \11827 );
not \U$12347 ( \12724 , \12722 );
and \U$12348 ( \12725 , \12724 , \12184 );
nor \U$12349 ( \12726 , \12723 , \12725 );
and \U$12350 ( \12727 , \12719 , \12726 );
and \U$12351 ( \12728 , \12716 , \12718 );
or \U$12352 ( \12729 , \12727 , \12728 );
or \U$12353 ( \12730 , \12709 , \12729 );
not \U$12354 ( \12731 , \12729 );
not \U$12355 ( \12732 , \12709 );
or \U$12356 ( \12733 , \12731 , \12732 );
and \U$12357 ( \12734 , \9760 , RIae76a78_55);
and \U$12358 ( \12735 , RIae76988_53, \9758 );
nor \U$12359 ( \12736 , \12734 , \12735 );
and \U$12360 ( \12737 , \12736 , \9764 );
not \U$12361 ( \12738 , \12736 );
and \U$12362 ( \12739 , \12738 , \9273 );
nor \U$12363 ( \12740 , \12737 , \12739 );
and \U$12364 ( \12741 , \10548 , RIae767a8_49);
and \U$12365 ( \12742 , RIae76898_51, \10546 );
nor \U$12366 ( \12743 , \12741 , \12742 );
and \U$12367 ( \12744 , \12743 , \10118 );
not \U$12368 ( \12745 , \12743 );
and \U$12369 ( \12746 , \12745 , \10421 );
nor \U$12370 ( \12747 , \12744 , \12746 );
xor \U$12371 ( \12748 , \12740 , \12747 );
and \U$12372 ( \12749 , \8966 , RIae762f8_39);
and \U$12373 ( \12750 , RIae76208_37, \8964 );
nor \U$12374 ( \12751 , \12749 , \12750 );
and \U$12375 ( \12752 , \12751 , \8789 );
not \U$12376 ( \12753 , \12751 );
and \U$12377 ( \12754 , \12753 , \8799 );
nor \U$12378 ( \12755 , \12752 , \12754 );
and \U$12379 ( \12756 , \12748 , \12755 );
and \U$12380 ( \12757 , \12740 , \12747 );
nor \U$12381 ( \12758 , \12756 , \12757 );
nand \U$12382 ( \12759 , \12733 , \12758 );
nand \U$12383 ( \12760 , \12730 , \12759 );
xor \U$12384 ( \12761 , \12684 , \12760 );
and \U$12385 ( \12762 , \2607 , RIae78788_117);
and \U$12386 ( \12763 , RIae78698_115, \2605 );
nor \U$12387 ( \12764 , \12762 , \12763 );
and \U$12388 ( \12765 , \12764 , \2397 );
not \U$12389 ( \12766 , \12764 );
and \U$12390 ( \12767 , \12766 , \2611 );
nor \U$12391 ( \12768 , \12765 , \12767 );
and \U$12392 ( \12769 , \2783 , RIae75b78_23);
and \U$12393 ( \12770 , RIae75a88_21, \2781 );
nor \U$12394 ( \12771 , \12769 , \12770 );
not \U$12395 ( \12772 , \12771 );
not \U$12396 ( \12773 , \2789 );
and \U$12397 ( \12774 , \12772 , \12773 );
and \U$12398 ( \12775 , \12771 , \3089 );
nor \U$12399 ( \12776 , \12774 , \12775 );
xor \U$12400 ( \12777 , \12768 , \12776 );
and \U$12401 ( \12778 , \3214 , RIae75998_19);
and \U$12402 ( \12779 , RIae758a8_17, \3212 );
nor \U$12403 ( \12780 , \12778 , \12779 );
not \U$12404 ( \12781 , \12780 );
not \U$12405 ( \12782 , \3218 );
and \U$12406 ( \12783 , \12781 , \12782 );
and \U$12407 ( \12784 , \12780 , \3218 );
nor \U$12408 ( \12785 , \12783 , \12784 );
and \U$12409 ( \12786 , \12777 , \12785 );
and \U$12410 ( \12787 , \12768 , \12776 );
or \U$12411 ( \12788 , \12786 , \12787 );
and \U$12412 ( \12789 , \3730 , RIae75f38_31);
and \U$12413 ( \12790 , RIae75e48_29, \3728 );
nor \U$12414 ( \12791 , \12789 , \12790 );
and \U$12415 ( \12792 , \12791 , \3422 );
not \U$12416 ( \12793 , \12791 );
and \U$12417 ( \12794 , \12793 , \3732 );
nor \U$12418 ( \12795 , \12792 , \12794 );
not \U$12419 ( \12796 , \12795 );
and \U$12420 ( \12797 , \4688 , RIae755d8_11);
and \U$12421 ( \12798 , RIae754e8_9, \4686 );
nor \U$12422 ( \12799 , \12797 , \12798 );
and \U$12423 ( \12800 , \12799 , \4482 );
not \U$12424 ( \12801 , \12799 );
and \U$12425 ( \12802 , \12801 , \4481 );
nor \U$12426 ( \12803 , \12800 , \12802 );
not \U$12427 ( \12804 , \12803 );
and \U$12428 ( \12805 , \12796 , \12804 );
and \U$12429 ( \12806 , \12803 , \12795 );
and \U$12430 ( \12807 , \4247 , RIae75c68_25);
and \U$12431 ( \12808 , RIae75d58_27, \4245 );
nor \U$12432 ( \12809 , \12807 , \12808 );
and \U$12433 ( \12810 , \12809 , \4251 );
not \U$12434 ( \12811 , \12809 );
and \U$12435 ( \12812 , \12811 , \3989 );
nor \U$12436 ( \12813 , \12810 , \12812 );
nor \U$12437 ( \12814 , \12806 , \12813 );
nor \U$12438 ( \12815 , \12805 , \12814 );
xor \U$12439 ( \12816 , \12788 , \12815 );
and \U$12440 ( \12817 , \6172 , RIae75308_5);
and \U$12441 ( \12818 , RIae753f8_7, \6170 );
nor \U$12442 ( \12819 , \12817 , \12818 );
and \U$12443 ( \12820 , \12819 , \6175 );
not \U$12444 ( \12821 , \12819 );
and \U$12445 ( \12822 , \12821 , \6176 );
nor \U$12446 ( \12823 , \12820 , \12822 );
and \U$12447 ( \12824 , \5399 , RIae757b8_15);
and \U$12448 ( \12825 , RIae756c8_13, \5397 );
nor \U$12449 ( \12826 , \12824 , \12825 );
and \U$12450 ( \12827 , \12826 , \5403 );
not \U$12451 ( \12828 , \12826 );
and \U$12452 ( \12829 , \12828 , \5016 );
nor \U$12453 ( \12830 , \12827 , \12829 );
xor \U$12454 ( \12831 , \12823 , \12830 );
and \U$12455 ( \12832 , \5896 , RIae75218_3);
and \U$12456 ( \12833 , RIae75128_1, \5894 );
nor \U$12457 ( \12834 , \12832 , \12833 );
and \U$12458 ( \12835 , \12834 , \5589 );
not \U$12459 ( \12836 , \12834 );
and \U$12460 ( \12837 , \12836 , \5590 );
nor \U$12461 ( \12838 , \12835 , \12837 );
and \U$12462 ( \12839 , \12831 , \12838 );
and \U$12463 ( \12840 , \12823 , \12830 );
or \U$12464 ( \12841 , \12839 , \12840 );
and \U$12465 ( \12842 , \12816 , \12841 );
and \U$12466 ( \12843 , \12788 , \12815 );
nor \U$12467 ( \12844 , \12842 , \12843 );
and \U$12468 ( \12845 , \12761 , \12844 );
and \U$12469 ( \12846 , \12684 , \12760 );
or \U$12470 ( \12847 , \12845 , \12846 );
xor \U$12471 ( \12848 , \12601 , \12847 );
not \U$12472 ( \12849 , \12396 );
not \U$12473 ( \12850 , \12390 );
or \U$12474 ( \12851 , \12849 , \12850 );
or \U$12475 ( \12852 , \12396 , \12390 );
nand \U$12476 ( \12853 , \12851 , \12852 );
xor \U$12477 ( \12854 , \12388 , \12853 );
not \U$12478 ( \12855 , \12329 );
xor \U$12479 ( \12856 , \12341 , \12318 );
not \U$12480 ( \12857 , \12856 );
or \U$12481 ( \12858 , \12855 , \12857 );
or \U$12482 ( \12859 , \12856 , \12329 );
nand \U$12483 ( \12860 , \12858 , \12859 );
xor \U$12484 ( \12861 , \12854 , \12860 );
not \U$12485 ( \12862 , \12412 );
xor \U$12486 ( \12863 , \12401 , \12417 );
not \U$12487 ( \12864 , \12863 );
or \U$12488 ( \12865 , \12862 , \12864 );
or \U$12489 ( \12866 , \12863 , \12412 );
nand \U$12490 ( \12867 , \12865 , \12866 );
and \U$12491 ( \12868 , \12861 , \12867 );
and \U$12492 ( \12869 , \12854 , \12860 );
or \U$12493 ( \12870 , \12868 , \12869 );
and \U$12494 ( \12871 , \12848 , \12870 );
and \U$12495 ( \12872 , \12601 , \12847 );
or \U$12496 ( \12873 , \12871 , \12872 );
nand \U$12497 ( \12874 , \12538 , \12873 );
nand \U$12498 ( \12875 , \12535 , \12874 );
xor \U$12499 ( \12876 , \12481 , \12875 );
xor \U$12500 ( \12877 , \11664 , \11666 );
xor \U$12501 ( \12878 , \12877 , \11669 );
xor \U$12502 ( \12879 , \12018 , \12025 );
xor \U$12503 ( \12880 , \12878 , \12879 );
and \U$12504 ( \12881 , \12876 , \12880 );
and \U$12505 ( \12882 , \12481 , \12875 );
or \U$12506 ( \12883 , \12881 , \12882 );
xor \U$12507 ( \12884 , \12030 , \12445 );
xor \U$12508 ( \12885 , \12884 , \12448 );
and \U$12509 ( \12886 , \12883 , \12885 );
and \U$12510 ( \12887 , \12464 , \12883 );
or \U$12511 ( \12888 , \12467 , \12886 , \12887 );
not \U$12512 ( \12889 , \12888 );
xnor \U$12513 ( \12890 , \12010 , \12451 );
not \U$12514 ( \12891 , \12890 );
not \U$12515 ( \12892 , \12013 );
and \U$12516 ( \12893 , \12891 , \12892 );
and \U$12517 ( \12894 , \12890 , \12013 );
nor \U$12518 ( \12895 , \12893 , \12894 );
nor \U$12519 ( \12896 , \12889 , \12895 );
and \U$12520 ( \12897 , \12462 , \12896 );
xor \U$12521 ( \12898 , \12896 , \12462 );
xor \U$12522 ( \12899 , \12166 , \12197 );
xor \U$12523 ( \12900 , \12899 , \12223 );
not \U$12524 ( \12901 , \12900 );
xor \U$12525 ( \12902 , \12628 , \12654 );
xor \U$12526 ( \12903 , \12902 , \12681 );
xor \U$12527 ( \12904 , \12573 , \12575 );
xor \U$12528 ( \12905 , \12904 , \12582 );
and \U$12529 ( \12906 , \12903 , \12905 );
xor \U$12530 ( \12907 , \12094 , \12101 );
xor \U$12531 ( \12908 , \12907 , \12109 );
xor \U$12532 ( \12909 , \12540 , \12545 );
xor \U$12533 ( \12910 , \12908 , \12909 );
xor \U$12534 ( \12911 , \12573 , \12575 );
xor \U$12535 ( \12912 , \12911 , \12582 );
and \U$12536 ( \12913 , \12910 , \12912 );
and \U$12537 ( \12914 , \12903 , \12910 );
or \U$12538 ( \12915 , \12906 , \12913 , \12914 );
not \U$12539 ( \12916 , \12915 );
or \U$12540 ( \12917 , \12901 , \12916 );
or \U$12541 ( \12918 , \12915 , \12900 );
nand \U$12542 ( \12919 , \12917 , \12918 );
not \U$12543 ( \12920 , \12919 );
not \U$12544 ( \12921 , \12483 );
not \U$12545 ( \12922 , \12491 );
or \U$12546 ( \12923 , \12921 , \12922 );
or \U$12547 ( \12924 , \12483 , \12491 );
nand \U$12548 ( \12925 , \12923 , \12924 );
not \U$12549 ( \12926 , \12925 );
not \U$12550 ( \12927 , \12485 );
and \U$12551 ( \12928 , \12926 , \12927 );
and \U$12552 ( \12929 , \12925 , \12485 );
nor \U$12553 ( \12930 , \12928 , \12929 );
not \U$12554 ( \12931 , \12930 );
and \U$12555 ( \12932 , \12920 , \12931 );
and \U$12556 ( \12933 , \12919 , \12930 );
nor \U$12557 ( \12934 , \12932 , \12933 );
and \U$12558 ( \12935 , \1593 , RIae78530_112);
and \U$12559 ( \12936 , RIae77c48_93, \1591 );
nor \U$12560 ( \12937 , \12935 , \12936 );
and \U$12561 ( \12938 , \12937 , \1488 );
not \U$12562 ( \12939 , \12937 );
and \U$12563 ( \12940 , \12939 , \1498 );
nor \U$12564 ( \12941 , \12938 , \12940 );
not \U$12565 ( \12942 , \12941 );
and \U$12566 ( \12943 , \2224 , RIae77e28_97);
and \U$12567 ( \12944 , RIae78968_121, \2222 );
nor \U$12568 ( \12945 , \12943 , \12944 );
and \U$12569 ( \12946 , \12945 , \2060 );
not \U$12570 ( \12947 , \12945 );
and \U$12571 ( \12948 , \12947 , \2061 );
nor \U$12572 ( \12949 , \12946 , \12948 );
not \U$12573 ( \12950 , \12949 );
and \U$12574 ( \12951 , \12942 , \12950 );
and \U$12575 ( \12952 , \12949 , \12941 );
and \U$12576 ( \12953 , \1939 , RIae77b58_91);
and \U$12577 ( \12954 , RIae77d38_95, \1937 );
nor \U$12578 ( \12955 , \12953 , \12954 );
and \U$12579 ( \12956 , \12955 , \1734 );
not \U$12580 ( \12957 , \12955 );
and \U$12581 ( \12958 , \12957 , \1735 );
nor \U$12582 ( \12959 , \12956 , \12958 );
nor \U$12583 ( \12960 , \12952 , \12959 );
nor \U$12584 ( \12961 , \12951 , \12960 );
and \U$12585 ( \12962 , \883 , RIae780f8_103);
and \U$12586 ( \12963 , RIae77f18_99, \881 );
nor \U$12587 ( \12964 , \12962 , \12963 );
not \U$12588 ( \12965 , \12964 );
not \U$12589 ( \12966 , \787 );
and \U$12590 ( \12967 , \12965 , \12966 );
and \U$12591 ( \12968 , \12964 , \787 );
nor \U$12592 ( \12969 , \12967 , \12968 );
not \U$12593 ( \12970 , \12969 );
and \U$12594 ( \12971 , \1376 , RIae785a8_113);
and \U$12595 ( \12972 , RIae783c8_109, \1374 );
nor \U$12596 ( \12973 , \12971 , \12972 );
and \U$12597 ( \12974 , \12973 , \1261 );
not \U$12598 ( \12975 , \12973 );
and \U$12599 ( \12976 , \12975 , \1380 );
nor \U$12600 ( \12977 , \12974 , \12976 );
not \U$12601 ( \12978 , \12977 );
and \U$12602 ( \12979 , \12970 , \12978 );
and \U$12603 ( \12980 , \12977 , \12969 );
and \U$12604 ( \12981 , \1138 , RIae78008_101);
and \U$12605 ( \12982 , RIae781e8_105, \1136 );
nor \U$12606 ( \12983 , \12981 , \12982 );
and \U$12607 ( \12984 , \12983 , \1142 );
not \U$12608 ( \12985 , \12983 );
and \U$12609 ( \12986 , \12985 , \1012 );
nor \U$12610 ( \12987 , \12984 , \12986 );
nor \U$12611 ( \12988 , \12980 , \12987 );
nor \U$12612 ( \12989 , \12979 , \12988 );
xor \U$12613 ( \12990 , \12961 , \12989 );
and \U$12614 ( \12991 , \558 , RIae77018_67);
and \U$12615 ( \12992 , RIae771f8_71, \556 );
nor \U$12616 ( \12993 , \12991 , \12992 );
and \U$12617 ( \12994 , \12993 , \504 );
not \U$12618 ( \12995 , \12993 );
and \U$12619 ( \12996 , \12995 , \562 );
nor \U$12620 ( \12997 , \12994 , \12996 );
and \U$12621 ( \12998 , \672 , RIae772e8_73);
and \U$12622 ( \12999 , RIae782d8_107, \670 );
nor \U$12623 ( \13000 , \12998 , \12999 );
and \U$12624 ( \13001 , \13000 , \588 );
not \U$12625 ( \13002 , \13000 );
and \U$12626 ( \13003 , \13002 , \587 );
nor \U$12627 ( \13004 , \13001 , \13003 );
xor \U$12628 ( \13005 , \12997 , \13004 );
not \U$12629 ( \13006 , \471 );
and \U$12630 ( \13007 , \514 , RIae76c58_59);
and \U$12631 ( \13008 , RIae77180_70, \512 );
nor \U$12632 ( \13009 , \13007 , \13008 );
not \U$12633 ( \13010 , \13009 );
or \U$12634 ( \13011 , \13006 , \13010 );
or \U$12635 ( \13012 , \13009 , \471 );
nand \U$12636 ( \13013 , \13011 , \13012 );
and \U$12637 ( \13014 , \13005 , \13013 );
and \U$12638 ( \13015 , \12997 , \13004 );
nor \U$12639 ( \13016 , \13014 , \13015 );
and \U$12640 ( \13017 , \12990 , \13016 );
and \U$12641 ( \13018 , \12961 , \12989 );
or \U$12642 ( \13019 , \13017 , \13018 );
and \U$12643 ( \13020 , \7633 , RIae764d8_43);
and \U$12644 ( \13021 , RIae766b8_47, \7631 );
nor \U$12645 ( \13022 , \13020 , \13021 );
and \U$12646 ( \13023 , \13022 , \7205 );
not \U$12647 ( \13024 , \13022 );
and \U$12648 ( \13025 , \13024 , \7206 );
nor \U$12649 ( \13026 , \13023 , \13025 );
and \U$12650 ( \13027 , \6941 , RIae753f8_7);
and \U$12651 ( \13028 , RIae763e8_41, \6939 );
nor \U$12652 ( \13029 , \13027 , \13028 );
and \U$12653 ( \13030 , \13029 , \6945 );
not \U$12654 ( \13031 , \13029 );
and \U$12655 ( \13032 , \13031 , \6314 );
nor \U$12656 ( \13033 , \13030 , \13032 );
xor \U$12657 ( \13034 , \13026 , \13033 );
and \U$12658 ( \13035 , \8371 , RIae765c8_45);
and \U$12659 ( \13036 , RIae76118_35, \8369 );
nor \U$12660 ( \13037 , \13035 , \13036 );
and \U$12661 ( \13038 , \13037 , \8019 );
not \U$12662 ( \13039 , \13037 );
and \U$12663 ( \13040 , \13039 , \8020 );
nor \U$12664 ( \13041 , \13038 , \13040 );
and \U$12665 ( \13042 , \13034 , \13041 );
and \U$12666 ( \13043 , \13026 , \13033 );
or \U$12667 ( \13044 , \13042 , \13043 );
and \U$12668 ( \13045 , \11470 , RIae76898_51);
and \U$12669 ( \13046 , RIae76b68_57, \11468 );
nor \U$12670 ( \13047 , \13045 , \13046 );
and \U$12671 ( \13048 , \13047 , \11474 );
not \U$12672 ( \13049 , \13047 );
and \U$12673 ( \13050 , \13049 , \10936 );
nor \U$12674 ( \13051 , \13048 , \13050 );
and \U$12675 ( \13052 , RIae7a7e0_186, RIae7a768_185);
not \U$12676 ( \13053 , RIae7a768_185);
nor \U$12677 ( \13054 , \13053 , RIae7a6f0_184);
not \U$12678 ( \13055 , RIae7a6f0_184);
nor \U$12679 ( \13056 , \13055 , RIae7a768_185);
or \U$12680 ( \13057 , \13054 , \13056 );
nor \U$12681 ( \13058 , RIae7a7e0_186, RIae7a768_185);
nor \U$12682 ( \13059 , \13052 , \13057 , \13058 );
nand \U$12683 ( \13060 , RIae78da0_130, \13059 );
and \U$12684 ( \13061 , \13060 , \12718 );
not \U$12685 ( \13062 , \13060 );
not \U$12686 ( \13063 , \12718 );
and \U$12687 ( \13064 , \13062 , \13063 );
nor \U$12688 ( \13065 , \13061 , \13064 );
xor \U$12689 ( \13066 , \13051 , \13065 );
and \U$12690 ( \13067 , \12180 , RIae78a58_123);
and \U$12691 ( \13068 , RIae78cb0_128, \12178 );
nor \U$12692 ( \13069 , \13067 , \13068 );
and \U$12693 ( \13070 , \13069 , \11827 );
not \U$12694 ( \13071 , \13069 );
and \U$12695 ( \13072 , \13071 , \12184 );
nor \U$12696 ( \13073 , \13070 , \13072 );
and \U$12697 ( \13074 , \13066 , \13073 );
and \U$12698 ( \13075 , \13051 , \13065 );
or \U$12699 ( \13076 , \13074 , \13075 );
xor \U$12700 ( \13077 , \13044 , \13076 );
and \U$12701 ( \13078 , \10548 , RIae76988_53);
and \U$12702 ( \13079 , RIae767a8_49, \10546 );
nor \U$12703 ( \13080 , \13078 , \13079 );
and \U$12704 ( \13081 , \13080 , \10118 );
not \U$12705 ( \13082 , \13080 );
and \U$12706 ( \13083 , \13082 , \10421 );
nor \U$12707 ( \13084 , \13081 , \13083 );
and \U$12708 ( \13085 , \8966 , RIae76028_33);
and \U$12709 ( \13086 , RIae762f8_39, \8964 );
nor \U$12710 ( \13087 , \13085 , \13086 );
and \U$12711 ( \13088 , \13087 , \8789 );
not \U$12712 ( \13089 , \13087 );
and \U$12713 ( \13090 , \13089 , \8799 );
nor \U$12714 ( \13091 , \13088 , \13090 );
xor \U$12715 ( \13092 , \13084 , \13091 );
and \U$12716 ( \13093 , \9760 , RIae76208_37);
and \U$12717 ( \13094 , RIae76a78_55, \9758 );
nor \U$12718 ( \13095 , \13093 , \13094 );
and \U$12719 ( \13096 , \13095 , \9272 );
not \U$12720 ( \13097 , \13095 );
and \U$12721 ( \13098 , \13097 , \9273 );
nor \U$12722 ( \13099 , \13096 , \13098 );
and \U$12723 ( \13100 , \13092 , \13099 );
and \U$12724 ( \13101 , \13084 , \13091 );
or \U$12725 ( \13102 , \13100 , \13101 );
and \U$12726 ( \13103 , \13077 , \13102 );
and \U$12727 ( \13104 , \13044 , \13076 );
or \U$12728 ( \13105 , \13103 , \13104 );
xor \U$12729 ( \13106 , \13019 , \13105 );
and \U$12730 ( \13107 , \5896 , RIae756c8_13);
and \U$12731 ( \13108 , RIae75218_3, \5894 );
nor \U$12732 ( \13109 , \13107 , \13108 );
and \U$12733 ( \13110 , \13109 , \5590 );
not \U$12734 ( \13111 , \13109 );
and \U$12735 ( \13112 , \13111 , \5589 );
nor \U$12736 ( \13113 , \13110 , \13112 );
and \U$12737 ( \13114 , \6172 , RIae75128_1);
and \U$12738 ( \13115 , RIae75308_5, \6170 );
nor \U$12739 ( \13116 , \13114 , \13115 );
and \U$12740 ( \13117 , \13116 , \6176 );
not \U$12741 ( \13118 , \13116 );
and \U$12742 ( \13119 , \13118 , \6175 );
nor \U$12743 ( \13120 , \13117 , \13119 );
xor \U$12744 ( \13121 , \13113 , \13120 );
and \U$12745 ( \13122 , \5399 , RIae754e8_9);
and \U$12746 ( \13123 , RIae757b8_15, \5397 );
nor \U$12747 ( \13124 , \13122 , \13123 );
and \U$12748 ( \13125 , \13124 , \5016 );
not \U$12749 ( \13126 , \13124 );
and \U$12750 ( \13127 , \13126 , \5403 );
nor \U$12751 ( \13128 , \13125 , \13127 );
and \U$12752 ( \13129 , \13121 , \13128 );
and \U$12753 ( \13130 , \13113 , \13120 );
nor \U$12754 ( \13131 , \13129 , \13130 );
not \U$12755 ( \13132 , \3089 );
and \U$12756 ( \13133 , \2783 , RIae78698_115);
and \U$12757 ( \13134 , RIae75b78_23, \2781 );
nor \U$12758 ( \13135 , \13133 , \13134 );
not \U$12759 ( \13136 , \13135 );
or \U$12760 ( \13137 , \13132 , \13136 );
or \U$12761 ( \13138 , \13135 , \3089 );
nand \U$12762 ( \13139 , \13137 , \13138 );
not \U$12763 ( \13140 , \2774 );
and \U$12764 ( \13141 , \3214 , RIae75a88_21);
and \U$12765 ( \13142 , RIae75998_19, \3212 );
nor \U$12766 ( \13143 , \13141 , \13142 );
not \U$12767 ( \13144 , \13143 );
or \U$12768 ( \13145 , \13140 , \13144 );
or \U$12769 ( \13146 , \13143 , \3218 );
nand \U$12770 ( \13147 , \13145 , \13146 );
xor \U$12771 ( \13148 , \13139 , \13147 );
and \U$12772 ( \13149 , \2607 , RIae78878_119);
and \U$12773 ( \13150 , RIae78788_117, \2605 );
nor \U$12774 ( \13151 , \13149 , \13150 );
and \U$12775 ( \13152 , \13151 , \2611 );
not \U$12776 ( \13153 , \13151 );
and \U$12777 ( \13154 , \13153 , \2397 );
nor \U$12778 ( \13155 , \13152 , \13154 );
and \U$12779 ( \13156 , \13148 , \13155 );
and \U$12780 ( \13157 , \13139 , \13147 );
nor \U$12781 ( \13158 , \13156 , \13157 );
xor \U$12782 ( \13159 , \13131 , \13158 );
and \U$12783 ( \13160 , \3730 , RIae758a8_17);
and \U$12784 ( \13161 , RIae75f38_31, \3728 );
nor \U$12785 ( \13162 , \13160 , \13161 );
and \U$12786 ( \13163 , \13162 , \3422 );
not \U$12787 ( \13164 , \13162 );
and \U$12788 ( \13165 , \13164 , \3732 );
nor \U$12789 ( \13166 , \13163 , \13165 );
not \U$12790 ( \13167 , \13166 );
and \U$12791 ( \13168 , \4247 , RIae75e48_29);
and \U$12792 ( \13169 , RIae75c68_25, \4245 );
nor \U$12793 ( \13170 , \13168 , \13169 );
and \U$12794 ( \13171 , \13170 , \4251 );
not \U$12795 ( \13172 , \13170 );
and \U$12796 ( \13173 , \13172 , \3989 );
nor \U$12797 ( \13174 , \13171 , \13173 );
not \U$12798 ( \13175 , \13174 );
and \U$12799 ( \13176 , \13167 , \13175 );
and \U$12800 ( \13177 , \13174 , \13166 );
and \U$12801 ( \13178 , \4688 , RIae75d58_27);
and \U$12802 ( \13179 , RIae755d8_11, \4686 );
nor \U$12803 ( \13180 , \13178 , \13179 );
and \U$12804 ( \13181 , \13180 , \4482 );
not \U$12805 ( \13182 , \13180 );
and \U$12806 ( \13183 , \13182 , \4481 );
nor \U$12807 ( \13184 , \13181 , \13183 );
nor \U$12808 ( \13185 , \13177 , \13184 );
nor \U$12809 ( \13186 , \13176 , \13185 );
and \U$12810 ( \13187 , \13159 , \13186 );
and \U$12811 ( \13188 , \13131 , \13158 );
or \U$12812 ( \13189 , \13187 , \13188 );
and \U$12813 ( \13190 , \13106 , \13189 );
and \U$12814 ( \13191 , \13019 , \13105 );
or \U$12815 ( \13192 , \13190 , \13191 );
not \U$12816 ( \13193 , \13192 );
xor \U$12817 ( \13194 , \12823 , \12830 );
xor \U$12818 ( \13195 , \13194 , \12838 );
xor \U$12819 ( \13196 , \12691 , \12698 );
xor \U$12820 ( \13197 , \13196 , \12706 );
or \U$12821 ( \13198 , \13195 , \13197 );
not \U$12822 ( \13199 , \13197 );
not \U$12823 ( \13200 , \13195 );
or \U$12824 ( \13201 , \13199 , \13200 );
not \U$12825 ( \13202 , \12795 );
xor \U$12826 ( \13203 , \12813 , \12803 );
not \U$12827 ( \13204 , \13203 );
or \U$12828 ( \13205 , \13202 , \13204 );
or \U$12829 ( \13206 , \13203 , \12795 );
nand \U$12830 ( \13207 , \13205 , \13206 );
nand \U$12831 ( \13208 , \13201 , \13207 );
nand \U$12832 ( \13209 , \13198 , \13208 );
not \U$12833 ( \13210 , \13209 );
xor \U$12834 ( \13211 , \12662 , \12669 );
xor \U$12835 ( \13212 , \13211 , \12678 );
and \U$12836 ( \13213 , \436 , RIae76e38_63);
and \U$12837 ( \13214 , RIae76d48_61, \434 );
nor \U$12838 ( \13215 , \13213 , \13214 );
not \U$12839 ( \13216 , \13215 );
not \U$12840 ( \13217 , \402 );
and \U$12841 ( \13218 , \13216 , \13217 );
and \U$12842 ( \13219 , \13215 , \400 );
nor \U$12843 ( \13220 , \13218 , \13219 );
nand \U$12844 ( \13221 , RIae77798_83, RIae78b48_125);
xor \U$12845 ( \13222 , \13220 , \13221 );
and \U$12846 ( \13223 , \384 , RIae77888_85);
and \U$12847 ( \13224 , RIae76f28_65, \382 );
nor \U$12848 ( \13225 , \13223 , \13224 );
not \U$12849 ( \13226 , \13225 );
not \U$12850 ( \13227 , \392 );
and \U$12851 ( \13228 , \13226 , \13227 );
and \U$12852 ( \13229 , \13225 , \388 );
nor \U$12853 ( \13230 , \13228 , \13229 );
and \U$12854 ( \13231 , \13222 , \13230 );
and \U$12855 ( \13232 , \13220 , \13221 );
or \U$12856 ( \13233 , \13231 , \13232 );
xor \U$12857 ( \13234 , \13212 , \13233 );
not \U$12858 ( \13235 , \12558 );
not \U$12859 ( \13236 , \12571 );
or \U$12860 ( \13237 , \13235 , \13236 );
or \U$12861 ( \13238 , \12558 , \12571 );
nand \U$12862 ( \13239 , \13237 , \13238 );
not \U$12863 ( \13240 , \13239 );
not \U$12864 ( \13241 , \12559 );
and \U$12865 ( \13242 , \13240 , \13241 );
and \U$12866 ( \13243 , \13239 , \12559 );
nor \U$12867 ( \13244 , \13242 , \13243 );
and \U$12868 ( \13245 , \13234 , \13244 );
and \U$12869 ( \13246 , \13212 , \13233 );
or \U$12870 ( \13247 , \13245 , \13246 );
or \U$12871 ( \13248 , \13210 , \13247 );
and \U$12872 ( \13249 , \13210 , \13247 );
not \U$12873 ( \13250 , \12615 );
not \U$12874 ( \13251 , \12626 );
or \U$12875 ( \13252 , \13250 , \13251 );
or \U$12876 ( \13253 , \12615 , \12626 );
nand \U$12877 ( \13254 , \13252 , \13253 );
not \U$12878 ( \13255 , \13254 );
not \U$12879 ( \13256 , \12608 );
and \U$12880 ( \13257 , \13255 , \13256 );
and \U$12881 ( \13258 , \13254 , \12608 );
nor \U$12882 ( \13259 , \13257 , \13258 );
xor \U$12883 ( \13260 , \12635 , \12642 );
xor \U$12884 ( \13261 , \13260 , \12651 );
xor \U$12885 ( \13262 , \13259 , \13261 );
xor \U$12886 ( \13263 , \12768 , \12776 );
xor \U$12887 ( \13264 , \13263 , \12785 );
and \U$12888 ( \13265 , \13262 , \13264 );
and \U$12889 ( \13266 , \13259 , \13261 );
or \U$12890 ( \13267 , \13265 , \13266 );
nor \U$12891 ( \13268 , \13249 , \13267 );
not \U$12892 ( \13269 , \13268 );
nand \U$12893 ( \13270 , \13248 , \13269 );
not \U$12894 ( \13271 , \13270 );
or \U$12895 ( \13272 , \13193 , \13271 );
or \U$12896 ( \13273 , \13270 , \13192 );
nand \U$12897 ( \13274 , \13272 , \13273 );
not \U$12898 ( \13275 , \13274 );
xor \U$12899 ( \13276 , \12173 , \12186 );
xor \U$12900 ( \13277 , \13276 , \12194 );
xor \U$12901 ( \13278 , \12205 , \12212 );
xor \U$12902 ( \13279 , \13278 , \12220 );
and \U$12903 ( \13280 , \13277 , \13279 );
not \U$12904 ( \13281 , \12588 );
not \U$12905 ( \13282 , \12596 );
or \U$12906 ( \13283 , \13281 , \13282 );
or \U$12907 ( \13284 , \12588 , \12596 );
nand \U$12908 ( \13285 , \13283 , \13284 );
not \U$12909 ( \13286 , \13285 );
not \U$12910 ( \13287 , \12590 );
and \U$12911 ( \13288 , \13286 , \13287 );
and \U$12912 ( \13289 , \13285 , \12590 );
nor \U$12913 ( \13290 , \13288 , \13289 );
xor \U$12914 ( \13291 , \12205 , \12212 );
xor \U$12915 ( \13292 , \13291 , \12220 );
and \U$12916 ( \13293 , \13290 , \13292 );
and \U$12917 ( \13294 , \13277 , \13290 );
or \U$12918 ( \13295 , \13280 , \13293 , \13294 );
not \U$12919 ( \13296 , \13295 );
and \U$12920 ( \13297 , \13275 , \13296 );
and \U$12921 ( \13298 , \13274 , \13295 );
nor \U$12922 ( \13299 , \13297 , \13298 );
or \U$12923 ( \13300 , \12934 , \13299 );
not \U$12924 ( \13301 , \13299 );
not \U$12925 ( \13302 , \12934 );
or \U$12926 ( \13303 , \13301 , \13302 );
xor \U$12927 ( \13304 , \12550 , \12585 );
xor \U$12928 ( \13305 , \13304 , \12598 );
xor \U$12929 ( \13306 , \12684 , \12760 );
xor \U$12930 ( \13307 , \13306 , \12844 );
xor \U$12931 ( \13308 , \12854 , \12860 );
xor \U$12932 ( \13309 , \13308 , \12867 );
xor \U$12933 ( \13310 , \13307 , \13309 );
xor \U$12934 ( \13311 , \13305 , \13310 );
nand \U$12935 ( \13312 , \13303 , \13311 );
nand \U$12936 ( \13313 , \13300 , \13312 );
xor \U$12937 ( \13314 , \12205 , \12212 );
xor \U$12938 ( \13315 , \13314 , \12220 );
xor \U$12939 ( \13316 , \13277 , \13290 );
xor \U$12940 ( \13317 , \13315 , \13316 );
not \U$12941 ( \13318 , \12758 );
not \U$12942 ( \13319 , \12729 );
or \U$12943 ( \13320 , \13318 , \13319 );
or \U$12944 ( \13321 , \12729 , \12758 );
nand \U$12945 ( \13322 , \13320 , \13321 );
not \U$12946 ( \13323 , \13322 );
not \U$12947 ( \13324 , \12709 );
and \U$12948 ( \13325 , \13323 , \13324 );
and \U$12949 ( \13326 , \13322 , \12709 );
nor \U$12950 ( \13327 , \13325 , \13326 );
or \U$12951 ( \13328 , \13317 , \13327 );
not \U$12952 ( \13329 , \13327 );
not \U$12953 ( \13330 , \13317 );
or \U$12954 ( \13331 , \13329 , \13330 );
xor \U$12955 ( \13332 , \12573 , \12575 );
xor \U$12956 ( \13333 , \13332 , \12582 );
xor \U$12957 ( \13334 , \12903 , \12910 );
xor \U$12958 ( \13335 , \13333 , \13334 );
nand \U$12959 ( \13336 , \13331 , \13335 );
nand \U$12960 ( \13337 , \13328 , \13336 );
not \U$12961 ( \13338 , \13337 );
xor \U$12962 ( \13339 , \13131 , \13158 );
xor \U$12963 ( \13340 , \13339 , \13186 );
xor \U$12964 ( \13341 , \13044 , \13076 );
xor \U$12965 ( \13342 , \13341 , \13102 );
xor \U$12966 ( \13343 , \13340 , \13342 );
xor \U$12967 ( \13344 , \12961 , \12989 );
xor \U$12968 ( \13345 , \13344 , \13016 );
and \U$12969 ( \13346 , \13343 , \13345 );
and \U$12970 ( \13347 , \13340 , \13342 );
or \U$12971 ( \13348 , \13346 , \13347 );
xor \U$12972 ( \13349 , \12788 , \12815 );
xor \U$12973 ( \13350 , \13349 , \12841 );
or \U$12974 ( \13351 , \13348 , \13350 );
not \U$12975 ( \13352 , \13350 );
not \U$12976 ( \13353 , \13348 );
or \U$12977 ( \13354 , \13352 , \13353 );
xor \U$12978 ( \13355 , \13259 , \13261 );
xor \U$12979 ( \13356 , \13355 , \13264 );
not \U$12980 ( \13357 , \13197 );
not \U$12981 ( \13358 , \13207 );
or \U$12982 ( \13359 , \13357 , \13358 );
or \U$12983 ( \13360 , \13197 , \13207 );
nand \U$12984 ( \13361 , \13359 , \13360 );
not \U$12985 ( \13362 , \13361 );
not \U$12986 ( \13363 , \13195 );
and \U$12987 ( \13364 , \13362 , \13363 );
and \U$12988 ( \13365 , \13361 , \13195 );
nor \U$12989 ( \13366 , \13364 , \13365 );
xor \U$12990 ( \13367 , \13356 , \13366 );
xor \U$12991 ( \13368 , \13212 , \13233 );
xor \U$12992 ( \13369 , \13368 , \13244 );
and \U$12993 ( \13370 , \13367 , \13369 );
and \U$12994 ( \13371 , \13356 , \13366 );
nor \U$12995 ( \13372 , \13370 , \13371 );
nand \U$12996 ( \13373 , \13354 , \13372 );
nand \U$12997 ( \13374 , \13351 , \13373 );
not \U$12998 ( \13375 , \13374 );
or \U$12999 ( \13376 , \13338 , \13375 );
or \U$13000 ( \13377 , \13374 , \13337 );
and \U$13001 ( \13378 , \4247 , RIae75f38_31);
and \U$13002 ( \13379 , RIae75e48_29, \4245 );
nor \U$13003 ( \13380 , \13378 , \13379 );
and \U$13004 ( \13381 , \13380 , \4251 );
not \U$13005 ( \13382 , \13380 );
and \U$13006 ( \13383 , \13382 , \3989 );
nor \U$13007 ( \13384 , \13381 , \13383 );
not \U$13008 ( \13385 , \13384 );
and \U$13009 ( \13386 , \5399 , RIae755d8_11);
and \U$13010 ( \13387 , RIae754e8_9, \5397 );
nor \U$13011 ( \13388 , \13386 , \13387 );
and \U$13012 ( \13389 , \13388 , \5403 );
not \U$13013 ( \13390 , \13388 );
and \U$13014 ( \13391 , \13390 , \5016 );
nor \U$13015 ( \13392 , \13389 , \13391 );
not \U$13016 ( \13393 , \13392 );
and \U$13017 ( \13394 , \13385 , \13393 );
and \U$13018 ( \13395 , \13392 , \13384 );
and \U$13019 ( \13396 , \4688 , RIae75c68_25);
and \U$13020 ( \13397 , RIae75d58_27, \4686 );
nor \U$13021 ( \13398 , \13396 , \13397 );
and \U$13022 ( \13399 , \13398 , \4482 );
not \U$13023 ( \13400 , \13398 );
and \U$13024 ( \13401 , \13400 , \4481 );
nor \U$13025 ( \13402 , \13399 , \13401 );
nor \U$13026 ( \13403 , \13395 , \13402 );
nor \U$13027 ( \13404 , \13394 , \13403 );
not \U$13028 ( \13405 , \13404 );
and \U$13029 ( \13406 , \5896 , RIae757b8_15);
and \U$13030 ( \13407 , RIae756c8_13, \5894 );
nor \U$13031 ( \13408 , \13406 , \13407 );
and \U$13032 ( \13409 , \13408 , \5589 );
not \U$13033 ( \13410 , \13408 );
and \U$13034 ( \13411 , \13410 , \5590 );
nor \U$13035 ( \13412 , \13409 , \13411 );
not \U$13036 ( \13413 , \13412 );
and \U$13037 ( \13414 , \6172 , RIae75218_3);
and \U$13038 ( \13415 , RIae75128_1, \6170 );
nor \U$13039 ( \13416 , \13414 , \13415 );
and \U$13040 ( \13417 , \13416 , \6175 );
not \U$13041 ( \13418 , \13416 );
and \U$13042 ( \13419 , \13418 , \6176 );
nor \U$13043 ( \13420 , \13417 , \13419 );
not \U$13044 ( \13421 , \13420 );
and \U$13045 ( \13422 , \13413 , \13421 );
and \U$13046 ( \13423 , \13420 , \13412 );
and \U$13047 ( \13424 , \6941 , RIae75308_5);
and \U$13048 ( \13425 , RIae753f8_7, \6939 );
nor \U$13049 ( \13426 , \13424 , \13425 );
and \U$13050 ( \13427 , \13426 , \6945 );
not \U$13051 ( \13428 , \13426 );
and \U$13052 ( \13429 , \13428 , \6314 );
nor \U$13053 ( \13430 , \13427 , \13429 );
nor \U$13054 ( \13431 , \13423 , \13430 );
nor \U$13055 ( \13432 , \13422 , \13431 );
not \U$13056 ( \13433 , \13432 );
and \U$13057 ( \13434 , \13405 , \13433 );
and \U$13058 ( \13435 , \13404 , \13432 );
and \U$13059 ( \13436 , \2783 , RIae78788_117);
and \U$13060 ( \13437 , RIae78698_115, \2781 );
nor \U$13061 ( \13438 , \13436 , \13437 );
not \U$13062 ( \13439 , \13438 );
not \U$13063 ( \13440 , \2789 );
and \U$13064 ( \13441 , \13439 , \13440 );
and \U$13065 ( \13442 , \13438 , \3089 );
nor \U$13066 ( \13443 , \13441 , \13442 );
not \U$13067 ( \13444 , \13443 );
and \U$13068 ( \13445 , \3214 , RIae75b78_23);
and \U$13069 ( \13446 , RIae75a88_21, \3212 );
nor \U$13070 ( \13447 , \13445 , \13446 );
not \U$13071 ( \13448 , \13447 );
not \U$13072 ( \13449 , \2774 );
and \U$13073 ( \13450 , \13448 , \13449 );
and \U$13074 ( \13451 , \13447 , \2774 );
nor \U$13075 ( \13452 , \13450 , \13451 );
not \U$13076 ( \13453 , \13452 );
and \U$13077 ( \13454 , \13444 , \13453 );
and \U$13078 ( \13455 , \13452 , \13443 );
and \U$13079 ( \13456 , \3730 , RIae75998_19);
and \U$13080 ( \13457 , RIae758a8_17, \3728 );
nor \U$13081 ( \13458 , \13456 , \13457 );
and \U$13082 ( \13459 , \13458 , \3422 );
not \U$13083 ( \13460 , \13458 );
and \U$13084 ( \13461 , \13460 , \3732 );
nor \U$13085 ( \13462 , \13459 , \13461 );
nor \U$13086 ( \13463 , \13455 , \13462 );
nor \U$13087 ( \13464 , \13454 , \13463 );
nor \U$13088 ( \13465 , \13435 , \13464 );
nor \U$13089 ( \13466 , \13434 , \13465 );
and \U$13090 ( \13467 , \8371 , RIae766b8_47);
and \U$13091 ( \13468 , RIae765c8_45, \8369 );
nor \U$13092 ( \13469 , \13467 , \13468 );
and \U$13093 ( \13470 , \13469 , \8020 );
not \U$13094 ( \13471 , \13469 );
and \U$13095 ( \13472 , \13471 , \8019 );
nor \U$13096 ( \13473 , \13470 , \13472 );
and \U$13097 ( \13474 , \7633 , RIae763e8_41);
and \U$13098 ( \13475 , RIae764d8_43, \7631 );
nor \U$13099 ( \13476 , \13474 , \13475 );
and \U$13100 ( \13477 , \13476 , \7206 );
not \U$13101 ( \13478 , \13476 );
and \U$13102 ( \13479 , \13478 , \7205 );
nor \U$13103 ( \13480 , \13477 , \13479 );
xor \U$13104 ( \13481 , \13473 , \13480 );
and \U$13105 ( \13482 , \8966 , RIae76118_35);
and \U$13106 ( \13483 , RIae76028_33, \8964 );
nor \U$13107 ( \13484 , \13482 , \13483 );
and \U$13108 ( \13485 , \13484 , \8799 );
not \U$13109 ( \13486 , \13484 );
and \U$13110 ( \13487 , \13486 , \8789 );
nor \U$13111 ( \13488 , \13485 , \13487 );
and \U$13112 ( \13489 , \13481 , \13488 );
and \U$13113 ( \13490 , \13473 , \13480 );
or \U$13114 ( \13491 , \13489 , \13490 );
and \U$13115 ( \13492 , \13059 , RIae78cb0_128);
and \U$13116 ( \13493 , RIae78da0_130, \13057 );
nor \U$13117 ( \13494 , \13492 , \13493 );
and \U$13118 ( \13495 , \13494 , \13063 );
not \U$13119 ( \13496 , \13494 );
and \U$13120 ( \13497 , \13496 , \12718 );
nor \U$13121 ( \13498 , \13495 , \13497 );
not \U$13122 ( \13499 , RIae7a8d0_188);
not \U$13123 ( \13500 , RIae7a858_187);
or \U$13124 ( \13501 , \13499 , \13500 );
nand \U$13125 ( \13502 , \13501 , RIae7a6f0_184);
xor \U$13126 ( \13503 , \13498 , \13502 );
and \U$13127 ( \13504 , \12180 , RIae76b68_57);
and \U$13128 ( \13505 , RIae78a58_123, \12178 );
nor \U$13129 ( \13506 , \13504 , \13505 );
and \U$13130 ( \13507 , \13506 , \12184 );
not \U$13131 ( \13508 , \13506 );
and \U$13132 ( \13509 , \13508 , \11827 );
nor \U$13133 ( \13510 , \13507 , \13509 );
and \U$13134 ( \13511 , \13503 , \13510 );
and \U$13135 ( \13512 , \13498 , \13502 );
or \U$13136 ( \13513 , \13511 , \13512 );
xor \U$13137 ( \13514 , \13491 , \13513 );
and \U$13138 ( \13515 , \11470 , RIae767a8_49);
and \U$13139 ( \13516 , RIae76898_51, \11468 );
nor \U$13140 ( \13517 , \13515 , \13516 );
and \U$13141 ( \13518 , \13517 , \10936 );
not \U$13142 ( \13519 , \13517 );
and \U$13143 ( \13520 , \13519 , \11474 );
nor \U$13144 ( \13521 , \13518 , \13520 );
and \U$13145 ( \13522 , \9760 , RIae762f8_39);
and \U$13146 ( \13523 , RIae76208_37, \9758 );
nor \U$13147 ( \13524 , \13522 , \13523 );
and \U$13148 ( \13525 , \13524 , \9273 );
not \U$13149 ( \13526 , \13524 );
and \U$13150 ( \13527 , \13526 , \9272 );
nor \U$13151 ( \13528 , \13525 , \13527 );
xor \U$13152 ( \13529 , \13521 , \13528 );
and \U$13153 ( \13530 , \10548 , RIae76a78_55);
and \U$13154 ( \13531 , RIae76988_53, \10546 );
nor \U$13155 ( \13532 , \13530 , \13531 );
and \U$13156 ( \13533 , \13532 , \10421 );
not \U$13157 ( \13534 , \13532 );
and \U$13158 ( \13535 , \13534 , \10118 );
nor \U$13159 ( \13536 , \13533 , \13535 );
and \U$13160 ( \13537 , \13529 , \13536 );
and \U$13161 ( \13538 , \13521 , \13528 );
or \U$13162 ( \13539 , \13537 , \13538 );
and \U$13163 ( \13540 , \13514 , \13539 );
and \U$13164 ( \13541 , \13491 , \13513 );
nor \U$13165 ( \13542 , \13540 , \13541 );
xor \U$13166 ( \13543 , \13466 , \13542 );
and \U$13167 ( \13544 , \558 , RIae77180_70);
and \U$13168 ( \13545 , RIae77018_67, \556 );
nor \U$13169 ( \13546 , \13544 , \13545 );
and \U$13170 ( \13547 , \13546 , \562 );
not \U$13171 ( \13548 , \13546 );
and \U$13172 ( \13549 , \13548 , \504 );
nor \U$13173 ( \13550 , \13547 , \13549 );
not \U$13174 ( \13551 , \13550 );
and \U$13175 ( \13552 , \883 , RIae782d8_107);
and \U$13176 ( \13553 , RIae780f8_103, \881 );
nor \U$13177 ( \13554 , \13552 , \13553 );
not \U$13178 ( \13555 , \13554 );
not \U$13179 ( \13556 , \789 );
and \U$13180 ( \13557 , \13555 , \13556 );
and \U$13181 ( \13558 , \13554 , \787 );
nor \U$13182 ( \13559 , \13557 , \13558 );
not \U$13183 ( \13560 , \13559 );
and \U$13184 ( \13561 , \13551 , \13560 );
and \U$13185 ( \13562 , \13559 , \13550 );
and \U$13186 ( \13563 , \672 , RIae771f8_71);
and \U$13187 ( \13564 , RIae772e8_73, \670 );
nor \U$13188 ( \13565 , \13563 , \13564 );
and \U$13189 ( \13566 , \13565 , \587 );
not \U$13190 ( \13567 , \13565 );
and \U$13191 ( \13568 , \13567 , \588 );
nor \U$13192 ( \13569 , \13566 , \13568 );
nor \U$13193 ( \13570 , \13562 , \13569 );
nor \U$13194 ( \13571 , \13561 , \13570 );
not \U$13195 ( \13572 , \13571 );
and \U$13196 ( \13573 , \1939 , RIae77c48_93);
and \U$13197 ( \13574 , RIae77b58_91, \1937 );
nor \U$13198 ( \13575 , \13573 , \13574 );
and \U$13199 ( \13576 , \13575 , \1734 );
not \U$13200 ( \13577 , \13575 );
and \U$13201 ( \13578 , \13577 , \1735 );
nor \U$13202 ( \13579 , \13576 , \13578 );
not \U$13203 ( \13580 , \13579 );
and \U$13204 ( \13581 , \2224 , RIae77d38_95);
and \U$13205 ( \13582 , RIae77e28_97, \2222 );
nor \U$13206 ( \13583 , \13581 , \13582 );
and \U$13207 ( \13584 , \13583 , \2060 );
not \U$13208 ( \13585 , \13583 );
and \U$13209 ( \13586 , \13585 , \2061 );
nor \U$13210 ( \13587 , \13584 , \13586 );
not \U$13211 ( \13588 , \13587 );
and \U$13212 ( \13589 , \13580 , \13588 );
and \U$13213 ( \13590 , \13587 , \13579 );
and \U$13214 ( \13591 , \2607 , RIae78968_121);
and \U$13215 ( \13592 , RIae78878_119, \2605 );
nor \U$13216 ( \13593 , \13591 , \13592 );
and \U$13217 ( \13594 , \13593 , \2397 );
not \U$13218 ( \13595 , \13593 );
and \U$13219 ( \13596 , \13595 , \2611 );
nor \U$13220 ( \13597 , \13594 , \13596 );
nor \U$13221 ( \13598 , \13590 , \13597 );
nor \U$13222 ( \13599 , \13589 , \13598 );
not \U$13223 ( \13600 , \13599 );
and \U$13224 ( \13601 , \13572 , \13600 );
and \U$13225 ( \13602 , \13571 , \13599 );
and \U$13226 ( \13603 , \1138 , RIae77f18_99);
and \U$13227 ( \13604 , RIae78008_101, \1136 );
nor \U$13228 ( \13605 , \13603 , \13604 );
and \U$13229 ( \13606 , \13605 , \1142 );
not \U$13230 ( \13607 , \13605 );
and \U$13231 ( \13608 , \13607 , \1012 );
nor \U$13232 ( \13609 , \13606 , \13608 );
not \U$13233 ( \13610 , \13609 );
and \U$13234 ( \13611 , \1376 , RIae781e8_105);
and \U$13235 ( \13612 , RIae785a8_113, \1374 );
nor \U$13236 ( \13613 , \13611 , \13612 );
and \U$13237 ( \13614 , \13613 , \1261 );
not \U$13238 ( \13615 , \13613 );
and \U$13239 ( \13616 , \13615 , \1380 );
nor \U$13240 ( \13617 , \13614 , \13616 );
not \U$13241 ( \13618 , \13617 );
and \U$13242 ( \13619 , \13610 , \13618 );
and \U$13243 ( \13620 , \13617 , \13609 );
and \U$13244 ( \13621 , \1593 , RIae783c8_109);
and \U$13245 ( \13622 , RIae78530_112, \1591 );
nor \U$13246 ( \13623 , \13621 , \13622 );
and \U$13247 ( \13624 , \13623 , \1488 );
not \U$13248 ( \13625 , \13623 );
and \U$13249 ( \13626 , \13625 , \1498 );
nor \U$13250 ( \13627 , \13624 , \13626 );
nor \U$13251 ( \13628 , \13620 , \13627 );
nor \U$13252 ( \13629 , \13619 , \13628 );
nor \U$13253 ( \13630 , \13602 , \13629 );
nor \U$13254 ( \13631 , \13601 , \13630 );
and \U$13255 ( \13632 , \13543 , \13631 );
and \U$13256 ( \13633 , \13466 , \13542 );
or \U$13257 ( \13634 , \13632 , \13633 );
xor \U$13258 ( \13635 , \12740 , \12747 );
xor \U$13259 ( \13636 , \13635 , \12755 );
xor \U$13260 ( \13637 , \12716 , \12718 );
xor \U$13261 ( \13638 , \13637 , \12726 );
xor \U$13262 ( \13639 , \13636 , \13638 );
xor \U$13263 ( \13640 , \13026 , \13033 );
xor \U$13264 ( \13641 , \13640 , \13041 );
not \U$13265 ( \13642 , \13641 );
xor \U$13266 ( \13643 , \13084 , \13091 );
xor \U$13267 ( \13644 , \13643 , \13099 );
not \U$13268 ( \13645 , \13644 );
and \U$13269 ( \13646 , \13642 , \13645 );
and \U$13270 ( \13647 , \13644 , \13641 );
xor \U$13271 ( \13648 , \13051 , \13065 );
xor \U$13272 ( \13649 , \13648 , \13073 );
nor \U$13273 ( \13650 , \13647 , \13649 );
nor \U$13274 ( \13651 , \13646 , \13650 );
and \U$13275 ( \13652 , \13639 , \13651 );
and \U$13276 ( \13653 , \13636 , \13638 );
or \U$13277 ( \13654 , \13652 , \13653 );
or \U$13278 ( \13655 , \13634 , \13654 );
not \U$13279 ( \13656 , \13654 );
not \U$13280 ( \13657 , \13634 );
or \U$13281 ( \13658 , \13656 , \13657 );
and \U$13282 ( \13659 , \384 , RIae77798_83);
and \U$13283 ( \13660 , RIae77888_85, \382 );
nor \U$13284 ( \13661 , \13659 , \13660 );
not \U$13285 ( \13662 , \13661 );
not \U$13286 ( \13663 , \388 );
and \U$13287 ( \13664 , \13662 , \13663 );
and \U$13288 ( \13665 , \13661 , \392 );
nor \U$13289 ( \13666 , \13664 , \13665 );
not \U$13290 ( \13667 , \13666 );
and \U$13291 ( \13668 , \514 , RIae76d48_61);
and \U$13292 ( \13669 , RIae76c58_59, \512 );
nor \U$13293 ( \13670 , \13668 , \13669 );
not \U$13294 ( \13671 , \13670 );
not \U$13295 ( \13672 , \469 );
and \U$13296 ( \13673 , \13671 , \13672 );
and \U$13297 ( \13674 , \13670 , \469 );
nor \U$13298 ( \13675 , \13673 , \13674 );
not \U$13299 ( \13676 , \13675 );
and \U$13300 ( \13677 , \13667 , \13676 );
and \U$13301 ( \13678 , \13675 , \13666 );
and \U$13302 ( \13679 , \436 , RIae76f28_65);
and \U$13303 ( \13680 , RIae76e38_63, \434 );
nor \U$13304 ( \13681 , \13679 , \13680 );
not \U$13305 ( \13682 , \13681 );
not \U$13306 ( \13683 , \402 );
and \U$13307 ( \13684 , \13682 , \13683 );
and \U$13308 ( \13685 , \13681 , \402 );
nor \U$13309 ( \13686 , \13684 , \13685 );
nor \U$13310 ( \13687 , \13678 , \13686 );
nor \U$13311 ( \13688 , \13677 , \13687 );
xor \U$13312 ( \13689 , \13220 , \13221 );
xor \U$13313 ( \13690 , \13689 , \13230 );
nand \U$13314 ( \13691 , \13688 , \13690 );
not \U$13315 ( \13692 , \13691 );
not \U$13316 ( \13693 , \13166 );
xor \U$13317 ( \13694 , \13174 , \13184 );
not \U$13318 ( \13695 , \13694 );
or \U$13319 ( \13696 , \13693 , \13695 );
or \U$13320 ( \13697 , \13694 , \13166 );
nand \U$13321 ( \13698 , \13696 , \13697 );
xor \U$13322 ( \13699 , \13139 , \13147 );
xor \U$13323 ( \13700 , \13699 , \13155 );
xor \U$13324 ( \13701 , \13698 , \13700 );
xor \U$13325 ( \13702 , \13113 , \13120 );
xor \U$13326 ( \13703 , \13702 , \13128 );
and \U$13327 ( \13704 , \13701 , \13703 );
and \U$13328 ( \13705 , \13698 , \13700 );
or \U$13329 ( \13706 , \13704 , \13705 );
not \U$13330 ( \13707 , \13706 );
or \U$13331 ( \13708 , \13692 , \13707 );
or \U$13332 ( \13709 , \13706 , \13691 );
xor \U$13333 ( \13710 , \12997 , \13004 );
xor \U$13334 ( \13711 , \13710 , \13013 );
not \U$13335 ( \13712 , \12969 );
xor \U$13336 ( \13713 , \12987 , \12977 );
not \U$13337 ( \13714 , \13713 );
or \U$13338 ( \13715 , \13712 , \13714 );
or \U$13339 ( \13716 , \13713 , \12969 );
nand \U$13340 ( \13717 , \13715 , \13716 );
xor \U$13341 ( \13718 , \13711 , \13717 );
not \U$13342 ( \13719 , \12941 );
xor \U$13343 ( \13720 , \12959 , \12949 );
not \U$13344 ( \13721 , \13720 );
or \U$13345 ( \13722 , \13719 , \13721 );
or \U$13346 ( \13723 , \13720 , \12941 );
nand \U$13347 ( \13724 , \13722 , \13723 );
and \U$13348 ( \13725 , \13718 , \13724 );
and \U$13349 ( \13726 , \13711 , \13717 );
or \U$13350 ( \13727 , \13725 , \13726 );
nand \U$13351 ( \13728 , \13709 , \13727 );
nand \U$13352 ( \13729 , \13708 , \13728 );
nand \U$13353 ( \13730 , \13658 , \13729 );
nand \U$13354 ( \13731 , \13655 , \13730 );
nand \U$13355 ( \13732 , \13377 , \13731 );
nand \U$13356 ( \13733 , \13376 , \13732 );
xor \U$13357 ( \13734 , \13313 , \13733 );
not \U$13358 ( \13735 , \12516 );
xor \U$13359 ( \13736 , \12527 , \12532 );
not \U$13360 ( \13737 , \13736 );
or \U$13361 ( \13738 , \13735 , \13737 );
or \U$13362 ( \13739 , \13736 , \12516 );
nand \U$13363 ( \13740 , \13738 , \13739 );
xor \U$13364 ( \13741 , \12601 , \12847 );
xor \U$13365 ( \13742 , \13741 , \12870 );
xor \U$13366 ( \13743 , \13740 , \13742 );
xor \U$13367 ( \13744 , \12032 , \12034 );
xor \U$13368 ( \13745 , \13744 , \12037 );
xor \U$13369 ( \13746 , \12493 , \12500 );
xor \U$13370 ( \13747 , \13745 , \13746 );
xor \U$13371 ( \13748 , \13743 , \13747 );
and \U$13372 ( \13749 , \13734 , \13748 );
and \U$13373 ( \13750 , \13313 , \13733 );
or \U$13374 ( \13751 , \13749 , \13750 );
not \U$13375 ( \13752 , \12873 );
not \U$13376 ( \13753 , \12534 );
or \U$13377 ( \13754 , \13752 , \13753 );
or \U$13378 ( \13755 , \12534 , \12873 );
nand \U$13379 ( \13756 , \13754 , \13755 );
not \U$13380 ( \13757 , \13756 );
not \U$13381 ( \13758 , \12506 );
and \U$13382 ( \13759 , \13757 , \13758 );
and \U$13383 ( \13760 , \13756 , \12506 );
nor \U$13384 ( \13761 , \13759 , \13760 );
not \U$13385 ( \13762 , \13761 );
xor \U$13386 ( \13763 , \12040 , \12042 );
xor \U$13387 ( \13764 , \13763 , \12057 );
xor \U$13388 ( \13765 , \12469 , \12476 );
xor \U$13389 ( \13766 , \13764 , \13765 );
not \U$13390 ( \13767 , \13766 );
or \U$13391 ( \13768 , \13762 , \13767 );
or \U$13392 ( \13769 , \13766 , \13761 );
nand \U$13393 ( \13770 , \13768 , \13769 );
xor \U$13394 ( \13771 , \13751 , \13770 );
or \U$13395 ( \13772 , \12930 , \12900 );
not \U$13396 ( \13773 , \12900 );
not \U$13397 ( \13774 , \12930 );
or \U$13398 ( \13775 , \13773 , \13774 );
nand \U$13399 ( \13776 , \13775 , \12915 );
nand \U$13400 ( \13777 , \13772 , \13776 );
or \U$13401 ( \13778 , \13192 , \13295 );
not \U$13402 ( \13779 , \13295 );
not \U$13403 ( \13780 , \13192 );
or \U$13404 ( \13781 , \13779 , \13780 );
nand \U$13405 ( \13782 , \13781 , \13270 );
nand \U$13406 ( \13783 , \13778 , \13782 );
xor \U$13407 ( \13784 , \13777 , \13783 );
xor \U$13408 ( \13785 , \12550 , \12585 );
xor \U$13409 ( \13786 , \13785 , \12598 );
and \U$13410 ( \13787 , \13307 , \13786 );
xor \U$13411 ( \13788 , \12550 , \12585 );
xor \U$13412 ( \13789 , \13788 , \12598 );
and \U$13413 ( \13790 , \13309 , \13789 );
and \U$13414 ( \13791 , \13307 , \13309 );
or \U$13415 ( \13792 , \13787 , \13790 , \13791 );
and \U$13416 ( \13793 , \13784 , \13792 );
and \U$13417 ( \13794 , \13777 , \13783 );
or \U$13418 ( \13795 , \13793 , \13794 );
xor \U$13419 ( \13796 , \12316 , \12361 );
xor \U$13420 ( \13797 , \13796 , \12422 );
xor \U$13421 ( \13798 , \13795 , \13797 );
xor \U$13422 ( \13799 , \13740 , \13742 );
and \U$13423 ( \13800 , \13799 , \13747 );
and \U$13424 ( \13801 , \13740 , \13742 );
or \U$13425 ( \13802 , \13800 , \13801 );
xor \U$13426 ( \13803 , \13798 , \13802 );
xor \U$13427 ( \13804 , \13771 , \13803 );
not \U$13428 ( \13805 , \13804 );
xor \U$13429 ( \13806 , \13313 , \13733 );
xor \U$13430 ( \13807 , \13806 , \13748 );
xor \U$13431 ( \13808 , \13777 , \13783 );
xor \U$13432 ( \13809 , \13808 , \13792 );
and \U$13433 ( \13810 , \13807 , \13809 );
not \U$13434 ( \13811 , \13807 );
not \U$13435 ( \13812 , \13809 );
and \U$13436 ( \13813 , \13811 , \13812 );
xor \U$13437 ( \13814 , \13466 , \13542 );
xor \U$13438 ( \13815 , \13814 , \13631 );
xor \U$13439 ( \13816 , \13636 , \13638 );
xor \U$13440 ( \13817 , \13816 , \13651 );
and \U$13441 ( \13818 , \13815 , \13817 );
xnor \U$13442 ( \13819 , \13706 , \13727 );
not \U$13443 ( \13820 , \13819 );
not \U$13444 ( \13821 , \13691 );
and \U$13445 ( \13822 , \13820 , \13821 );
and \U$13446 ( \13823 , \13819 , \13691 );
nor \U$13447 ( \13824 , \13822 , \13823 );
xor \U$13448 ( \13825 , \13636 , \13638 );
xor \U$13449 ( \13826 , \13825 , \13651 );
and \U$13450 ( \13827 , \13824 , \13826 );
and \U$13451 ( \13828 , \13815 , \13824 );
or \U$13452 ( \13829 , \13818 , \13827 , \13828 );
not \U$13453 ( \13830 , \13550 );
xor \U$13454 ( \13831 , \13569 , \13559 );
not \U$13455 ( \13832 , \13831 );
or \U$13456 ( \13833 , \13830 , \13832 );
or \U$13457 ( \13834 , \13831 , \13550 );
nand \U$13458 ( \13835 , \13833 , \13834 );
not \U$13459 ( \13836 , \13666 );
xor \U$13460 ( \13837 , \13686 , \13675 );
not \U$13461 ( \13838 , \13837 );
or \U$13462 ( \13839 , \13836 , \13838 );
or \U$13463 ( \13840 , \13837 , \13666 );
nand \U$13464 ( \13841 , \13839 , \13840 );
xor \U$13465 ( \13842 , \13835 , \13841 );
not \U$13466 ( \13843 , \13609 );
xor \U$13467 ( \13844 , \13617 , \13627 );
not \U$13468 ( \13845 , \13844 );
or \U$13469 ( \13846 , \13843 , \13845 );
or \U$13470 ( \13847 , \13844 , \13609 );
nand \U$13471 ( \13848 , \13846 , \13847 );
and \U$13472 ( \13849 , \13842 , \13848 );
and \U$13473 ( \13850 , \13835 , \13841 );
or \U$13474 ( \13851 , \13849 , \13850 );
nand \U$13475 ( \13852 , RIae77a68_89, RIae78b48_125);
not \U$13476 ( \13853 , \13852 );
not \U$13477 ( \13854 , RIae77978_87);
nor \U$13478 ( \13855 , \13854 , \491 );
xor \U$13479 ( \13856 , \13853 , \13855 );
not \U$13480 ( \13857 , \392 );
and \U$13481 ( \13858 , \384 , RIae77978_87);
and \U$13482 ( \13859 , RIae77798_83, \382 );
nor \U$13483 ( \13860 , \13858 , \13859 );
not \U$13484 ( \13861 , \13860 );
or \U$13485 ( \13862 , \13857 , \13861 );
or \U$13486 ( \13863 , \13860 , \392 );
nand \U$13487 ( \13864 , \13862 , \13863 );
not \U$13488 ( \13865 , \402 );
and \U$13489 ( \13866 , \436 , RIae77888_85);
and \U$13490 ( \13867 , RIae76f28_65, \434 );
nor \U$13491 ( \13868 , \13866 , \13867 );
not \U$13492 ( \13869 , \13868 );
or \U$13493 ( \13870 , \13865 , \13869 );
or \U$13494 ( \13871 , \13868 , \400 );
nand \U$13495 ( \13872 , \13870 , \13871 );
xor \U$13496 ( \13873 , \13864 , \13872 );
not \U$13497 ( \13874 , \469 );
and \U$13498 ( \13875 , \514 , RIae76e38_63);
and \U$13499 ( \13876 , RIae76d48_61, \512 );
nor \U$13500 ( \13877 , \13875 , \13876 );
not \U$13501 ( \13878 , \13877 );
or \U$13502 ( \13879 , \13874 , \13878 );
or \U$13503 ( \13880 , \13877 , \471 );
nand \U$13504 ( \13881 , \13879 , \13880 );
and \U$13505 ( \13882 , \13873 , \13881 );
and \U$13506 ( \13883 , \13864 , \13872 );
or \U$13507 ( \13884 , \13882 , \13883 );
and \U$13508 ( \13885 , \13856 , \13884 );
and \U$13509 ( \13886 , \13853 , \13855 );
or \U$13510 ( \13887 , \13885 , \13886 );
xor \U$13511 ( \13888 , \13851 , \13887 );
not \U$13512 ( \13889 , \13443 );
xor \U$13513 ( \13890 , \13452 , \13462 );
not \U$13514 ( \13891 , \13890 );
or \U$13515 ( \13892 , \13889 , \13891 );
or \U$13516 ( \13893 , \13890 , \13443 );
nand \U$13517 ( \13894 , \13892 , \13893 );
not \U$13518 ( \13895 , \13579 );
xor \U$13519 ( \13896 , \13587 , \13597 );
not \U$13520 ( \13897 , \13896 );
or \U$13521 ( \13898 , \13895 , \13897 );
or \U$13522 ( \13899 , \13896 , \13579 );
nand \U$13523 ( \13900 , \13898 , \13899 );
xor \U$13524 ( \13901 , \13894 , \13900 );
not \U$13525 ( \13902 , \13384 );
xor \U$13526 ( \13903 , \13402 , \13392 );
not \U$13527 ( \13904 , \13903 );
or \U$13528 ( \13905 , \13902 , \13904 );
or \U$13529 ( \13906 , \13903 , \13384 );
nand \U$13530 ( \13907 , \13905 , \13906 );
and \U$13531 ( \13908 , \13901 , \13907 );
and \U$13532 ( \13909 , \13894 , \13900 );
or \U$13533 ( \13910 , \13908 , \13909 );
and \U$13534 ( \13911 , \13888 , \13910 );
and \U$13535 ( \13912 , \13851 , \13887 );
nor \U$13536 ( \13913 , \13911 , \13912 );
and \U$13537 ( \13914 , \6941 , RIae75128_1);
and \U$13538 ( \13915 , RIae75308_5, \6939 );
nor \U$13539 ( \13916 , \13914 , \13915 );
and \U$13540 ( \13917 , \13916 , \6314 );
not \U$13541 ( \13918 , \13916 );
and \U$13542 ( \13919 , \13918 , \6945 );
nor \U$13543 ( \13920 , \13917 , \13919 );
and \U$13544 ( \13921 , \5896 , RIae754e8_9);
and \U$13545 ( \13922 , RIae757b8_15, \5894 );
nor \U$13546 ( \13923 , \13921 , \13922 );
and \U$13547 ( \13924 , \13923 , \5590 );
not \U$13548 ( \13925 , \13923 );
and \U$13549 ( \13926 , \13925 , \5589 );
nor \U$13550 ( \13927 , \13924 , \13926 );
xor \U$13551 ( \13928 , \13920 , \13927 );
and \U$13552 ( \13929 , \6172 , RIae756c8_13);
and \U$13553 ( \13930 , RIae75218_3, \6170 );
nor \U$13554 ( \13931 , \13929 , \13930 );
and \U$13555 ( \13932 , \13931 , \6176 );
not \U$13556 ( \13933 , \13931 );
and \U$13557 ( \13934 , \13933 , \6175 );
nor \U$13558 ( \13935 , \13932 , \13934 );
and \U$13559 ( \13936 , \13928 , \13935 );
and \U$13560 ( \13937 , \13920 , \13927 );
or \U$13561 ( \13938 , \13936 , \13937 );
and \U$13562 ( \13939 , \5399 , RIae75d58_27);
and \U$13563 ( \13940 , RIae755d8_11, \5397 );
nor \U$13564 ( \13941 , \13939 , \13940 );
and \U$13565 ( \13942 , \13941 , \5016 );
not \U$13566 ( \13943 , \13941 );
and \U$13567 ( \13944 , \13943 , \5403 );
nor \U$13568 ( \13945 , \13942 , \13944 );
and \U$13569 ( \13946 , \4247 , RIae758a8_17);
and \U$13570 ( \13947 , RIae75f38_31, \4245 );
nor \U$13571 ( \13948 , \13946 , \13947 );
and \U$13572 ( \13949 , \13948 , \3989 );
not \U$13573 ( \13950 , \13948 );
and \U$13574 ( \13951 , \13950 , \4251 );
nor \U$13575 ( \13952 , \13949 , \13951 );
xor \U$13576 ( \13953 , \13945 , \13952 );
and \U$13577 ( \13954 , \4688 , RIae75e48_29);
and \U$13578 ( \13955 , RIae75c68_25, \4686 );
nor \U$13579 ( \13956 , \13954 , \13955 );
and \U$13580 ( \13957 , \13956 , \4481 );
not \U$13581 ( \13958 , \13956 );
and \U$13582 ( \13959 , \13958 , \4482 );
nor \U$13583 ( \13960 , \13957 , \13959 );
and \U$13584 ( \13961 , \13953 , \13960 );
and \U$13585 ( \13962 , \13945 , \13952 );
or \U$13586 ( \13963 , \13961 , \13962 );
xor \U$13587 ( \13964 , \13938 , \13963 );
not \U$13588 ( \13965 , \2789 );
and \U$13589 ( \13966 , \2783 , RIae78878_119);
and \U$13590 ( \13967 , RIae78788_117, \2781 );
nor \U$13591 ( \13968 , \13966 , \13967 );
not \U$13592 ( \13969 , \13968 );
or \U$13593 ( \13970 , \13965 , \13969 );
or \U$13594 ( \13971 , \13968 , \3089 );
nand \U$13595 ( \13972 , \13970 , \13971 );
not \U$13596 ( \13973 , \3218 );
and \U$13597 ( \13974 , \3214 , RIae78698_115);
and \U$13598 ( \13975 , RIae75b78_23, \3212 );
nor \U$13599 ( \13976 , \13974 , \13975 );
not \U$13600 ( \13977 , \13976 );
or \U$13601 ( \13978 , \13973 , \13977 );
or \U$13602 ( \13979 , \13976 , \3218 );
nand \U$13603 ( \13980 , \13978 , \13979 );
xor \U$13604 ( \13981 , \13972 , \13980 );
and \U$13605 ( \13982 , \3730 , RIae75a88_21);
and \U$13606 ( \13983 , RIae75998_19, \3728 );
nor \U$13607 ( \13984 , \13982 , \13983 );
and \U$13608 ( \13985 , \13984 , \3732 );
not \U$13609 ( \13986 , \13984 );
and \U$13610 ( \13987 , \13986 , \3422 );
nor \U$13611 ( \13988 , \13985 , \13987 );
and \U$13612 ( \13989 , \13981 , \13988 );
and \U$13613 ( \13990 , \13972 , \13980 );
or \U$13614 ( \13991 , \13989 , \13990 );
and \U$13615 ( \13992 , \13964 , \13991 );
and \U$13616 ( \13993 , \13938 , \13963 );
or \U$13617 ( \13994 , \13992 , \13993 );
and \U$13618 ( \13995 , \10548 , RIae76208_37);
and \U$13619 ( \13996 , RIae76a78_55, \10546 );
nor \U$13620 ( \13997 , \13995 , \13996 );
and \U$13621 ( \13998 , \13997 , \10421 );
not \U$13622 ( \13999 , \13997 );
and \U$13623 ( \14000 , \13999 , \10118 );
nor \U$13624 ( \14001 , \13998 , \14000 );
and \U$13625 ( \14002 , \9760 , RIae76028_33);
and \U$13626 ( \14003 , RIae762f8_39, \9758 );
nor \U$13627 ( \14004 , \14002 , \14003 );
and \U$13628 ( \14005 , \14004 , \9273 );
not \U$13629 ( \14006 , \14004 );
and \U$13630 ( \14007 , \14006 , \9764 );
nor \U$13631 ( \14008 , \14005 , \14007 );
xor \U$13632 ( \14009 , \14001 , \14008 );
and \U$13633 ( \14010 , \11470 , RIae76988_53);
and \U$13634 ( \14011 , RIae767a8_49, \11468 );
nor \U$13635 ( \14012 , \14010 , \14011 );
and \U$13636 ( \14013 , \14012 , \10936 );
not \U$13637 ( \14014 , \14012 );
and \U$13638 ( \14015 , \14014 , \11474 );
nor \U$13639 ( \14016 , \14013 , \14015 );
and \U$13640 ( \14017 , \14009 , \14016 );
and \U$13641 ( \14018 , \14001 , \14008 );
or \U$13642 ( \14019 , \14017 , \14018 );
and \U$13643 ( \14020 , \8966 , RIae765c8_45);
and \U$13644 ( \14021 , RIae76118_35, \8964 );
nor \U$13645 ( \14022 , \14020 , \14021 );
and \U$13646 ( \14023 , \14022 , \8799 );
not \U$13647 ( \14024 , \14022 );
and \U$13648 ( \14025 , \14024 , \8789 );
nor \U$13649 ( \14026 , \14023 , \14025 );
and \U$13650 ( \14027 , \7633 , RIae753f8_7);
and \U$13651 ( \14028 , RIae763e8_41, \7631 );
nor \U$13652 ( \14029 , \14027 , \14028 );
and \U$13653 ( \14030 , \14029 , \7206 );
not \U$13654 ( \14031 , \14029 );
and \U$13655 ( \14032 , \14031 , \7205 );
nor \U$13656 ( \14033 , \14030 , \14032 );
xor \U$13657 ( \14034 , \14026 , \14033 );
and \U$13658 ( \14035 , \8371 , RIae764d8_43);
and \U$13659 ( \14036 , RIae766b8_47, \8369 );
nor \U$13660 ( \14037 , \14035 , \14036 );
and \U$13661 ( \14038 , \14037 , \8020 );
not \U$13662 ( \14039 , \14037 );
and \U$13663 ( \14040 , \14039 , \8019 );
nor \U$13664 ( \14041 , \14038 , \14040 );
and \U$13665 ( \14042 , \14034 , \14041 );
and \U$13666 ( \14043 , \14026 , \14033 );
or \U$13667 ( \14044 , \14042 , \14043 );
xor \U$13668 ( \14045 , \14019 , \14044 );
and \U$13669 ( \14046 , \12180 , RIae76898_51);
and \U$13670 ( \14047 , RIae76b68_57, \12178 );
nor \U$13671 ( \14048 , \14046 , \14047 );
and \U$13672 ( \14049 , \14048 , \12184 );
not \U$13673 ( \14050 , \14048 );
and \U$13674 ( \14051 , \14050 , \11827 );
nor \U$13675 ( \14052 , \14049 , \14051 );
and \U$13676 ( \14053 , RIae7a6f0_184, RIae7a858_187);
not \U$13677 ( \14054 , RIae7a8d0_188);
and \U$13678 ( \14055 , \14054 , RIae7a858_187);
nor \U$13679 ( \14056 , \14054 , RIae7a858_187);
or \U$13680 ( \14057 , \14055 , \14056 );
nor \U$13681 ( \14058 , RIae7a6f0_184, RIae7a858_187);
nor \U$13682 ( \14059 , \14053 , \14057 , \14058 );
nand \U$13683 ( \14060 , RIae78da0_130, \14059 );
and \U$13684 ( \14061 , \14060 , \13502 );
not \U$13685 ( \14062 , \14060 );
not \U$13686 ( \14063 , \13502 );
and \U$13687 ( \14064 , \14062 , \14063 );
nor \U$13688 ( \14065 , \14061 , \14064 );
xor \U$13689 ( \14066 , \14052 , \14065 );
and \U$13690 ( \14067 , \13059 , RIae78a58_123);
and \U$13691 ( \14068 , RIae78cb0_128, \13057 );
nor \U$13692 ( \14069 , \14067 , \14068 );
and \U$13693 ( \14070 , \14069 , \13063 );
not \U$13694 ( \14071 , \14069 );
and \U$13695 ( \14072 , \14071 , \12718 );
nor \U$13696 ( \14073 , \14070 , \14072 );
and \U$13697 ( \14074 , \14066 , \14073 );
and \U$13698 ( \14075 , \14052 , \14065 );
or \U$13699 ( \14076 , \14074 , \14075 );
and \U$13700 ( \14077 , \14045 , \14076 );
and \U$13701 ( \14078 , \14019 , \14044 );
or \U$13702 ( \14079 , \14077 , \14078 );
xor \U$13703 ( \14080 , \13994 , \14079 );
and \U$13704 ( \14081 , \1376 , RIae78008_101);
and \U$13705 ( \14082 , RIae781e8_105, \1374 );
nor \U$13706 ( \14083 , \14081 , \14082 );
and \U$13707 ( \14084 , \14083 , \1380 );
not \U$13708 ( \14085 , \14083 );
and \U$13709 ( \14086 , \14085 , \1261 );
nor \U$13710 ( \14087 , \14084 , \14086 );
and \U$13711 ( \14088 , \1138 , RIae780f8_103);
and \U$13712 ( \14089 , RIae77f18_99, \1136 );
nor \U$13713 ( \14090 , \14088 , \14089 );
and \U$13714 ( \14091 , \14090 , \1012 );
not \U$13715 ( \14092 , \14090 );
and \U$13716 ( \14093 , \14092 , \1142 );
nor \U$13717 ( \14094 , \14091 , \14093 );
xor \U$13718 ( \14095 , \14087 , \14094 );
and \U$13719 ( \14096 , \1593 , RIae785a8_113);
and \U$13720 ( \14097 , RIae783c8_109, \1591 );
nor \U$13721 ( \14098 , \14096 , \14097 );
and \U$13722 ( \14099 , \14098 , \1498 );
not \U$13723 ( \14100 , \14098 );
and \U$13724 ( \14101 , \14100 , \1488 );
nor \U$13725 ( \14102 , \14099 , \14101 );
and \U$13726 ( \14103 , \14095 , \14102 );
and \U$13727 ( \14104 , \14087 , \14094 );
or \U$13728 ( \14105 , \14103 , \14104 );
and \U$13729 ( \14106 , \672 , RIae77018_67);
and \U$13730 ( \14107 , RIae771f8_71, \670 );
nor \U$13731 ( \14108 , \14106 , \14107 );
and \U$13732 ( \14109 , \14108 , \588 );
not \U$13733 ( \14110 , \14108 );
and \U$13734 ( \14111 , \14110 , \587 );
nor \U$13735 ( \14112 , \14109 , \14111 );
and \U$13736 ( \14113 , \558 , RIae76c58_59);
and \U$13737 ( \14114 , RIae77180_70, \556 );
nor \U$13738 ( \14115 , \14113 , \14114 );
and \U$13739 ( \14116 , \14115 , \504 );
not \U$13740 ( \14117 , \14115 );
and \U$13741 ( \14118 , \14117 , \562 );
nor \U$13742 ( \14119 , \14116 , \14118 );
xor \U$13743 ( \14120 , \14112 , \14119 );
not \U$13744 ( \14121 , \787 );
and \U$13745 ( \14122 , \883 , RIae772e8_73);
and \U$13746 ( \14123 , RIae782d8_107, \881 );
nor \U$13747 ( \14124 , \14122 , \14123 );
not \U$13748 ( \14125 , \14124 );
or \U$13749 ( \14126 , \14121 , \14125 );
or \U$13750 ( \14127 , \14124 , \787 );
nand \U$13751 ( \14128 , \14126 , \14127 );
and \U$13752 ( \14129 , \14120 , \14128 );
and \U$13753 ( \14130 , \14112 , \14119 );
or \U$13754 ( \14131 , \14129 , \14130 );
xor \U$13755 ( \14132 , \14105 , \14131 );
and \U$13756 ( \14133 , \2607 , RIae77e28_97);
and \U$13757 ( \14134 , RIae78968_121, \2605 );
nor \U$13758 ( \14135 , \14133 , \14134 );
and \U$13759 ( \14136 , \14135 , \2611 );
not \U$13760 ( \14137 , \14135 );
and \U$13761 ( \14138 , \14137 , \2397 );
nor \U$13762 ( \14139 , \14136 , \14138 );
and \U$13763 ( \14140 , \1939 , RIae78530_112);
and \U$13764 ( \14141 , RIae77c48_93, \1937 );
nor \U$13765 ( \14142 , \14140 , \14141 );
and \U$13766 ( \14143 , \14142 , \1735 );
not \U$13767 ( \14144 , \14142 );
and \U$13768 ( \14145 , \14144 , \1734 );
nor \U$13769 ( \14146 , \14143 , \14145 );
xor \U$13770 ( \14147 , \14139 , \14146 );
and \U$13771 ( \14148 , \2224 , RIae77b58_91);
and \U$13772 ( \14149 , RIae77d38_95, \2222 );
nor \U$13773 ( \14150 , \14148 , \14149 );
and \U$13774 ( \14151 , \14150 , \2061 );
not \U$13775 ( \14152 , \14150 );
and \U$13776 ( \14153 , \14152 , \2060 );
nor \U$13777 ( \14154 , \14151 , \14153 );
and \U$13778 ( \14155 , \14147 , \14154 );
and \U$13779 ( \14156 , \14139 , \14146 );
or \U$13780 ( \14157 , \14155 , \14156 );
and \U$13781 ( \14158 , \14132 , \14157 );
and \U$13782 ( \14159 , \14105 , \14131 );
or \U$13783 ( \14160 , \14158 , \14159 );
and \U$13784 ( \14161 , \14080 , \14160 );
and \U$13785 ( \14162 , \13994 , \14079 );
nor \U$13786 ( \14163 , \14161 , \14162 );
xor \U$13787 ( \14164 , \13913 , \14163 );
not \U$13788 ( \14165 , \13644 );
xor \U$13789 ( \14166 , \13649 , \13641 );
not \U$13790 ( \14167 , \14166 );
or \U$13791 ( \14168 , \14165 , \14167 );
or \U$13792 ( \14169 , \14166 , \13644 );
nand \U$13793 ( \14170 , \14168 , \14169 );
xor \U$13794 ( \14171 , \13698 , \13700 );
xor \U$13795 ( \14172 , \14171 , \13703 );
xor \U$13796 ( \14173 , \14170 , \14172 );
not \U$13797 ( \14174 , \13412 );
xor \U$13798 ( \14175 , \13420 , \13430 );
not \U$13799 ( \14176 , \14175 );
or \U$13800 ( \14177 , \14174 , \14176 );
or \U$13801 ( \14178 , \14175 , \13412 );
nand \U$13802 ( \14179 , \14177 , \14178 );
xor \U$13803 ( \14180 , \13473 , \13480 );
xor \U$13804 ( \14181 , \14180 , \13488 );
and \U$13805 ( \14182 , \14179 , \14181 );
xor \U$13806 ( \14183 , \13521 , \13528 );
xor \U$13807 ( \14184 , \14183 , \13536 );
xor \U$13808 ( \14185 , \13473 , \13480 );
xor \U$13809 ( \14186 , \14185 , \13488 );
and \U$13810 ( \14187 , \14184 , \14186 );
and \U$13811 ( \14188 , \14179 , \14184 );
or \U$13812 ( \14189 , \14182 , \14187 , \14188 );
and \U$13813 ( \14190 , \14173 , \14189 );
and \U$13814 ( \14191 , \14170 , \14172 );
nor \U$13815 ( \14192 , \14190 , \14191 );
and \U$13816 ( \14193 , \14164 , \14192 );
and \U$13817 ( \14194 , \13913 , \14163 );
or \U$13818 ( \14195 , \14193 , \14194 );
xor \U$13819 ( \14196 , \13829 , \14195 );
not \U$13820 ( \14197 , \13599 );
xor \U$13821 ( \14198 , \13571 , \13629 );
not \U$13822 ( \14199 , \14198 );
or \U$13823 ( \14200 , \14197 , \14199 );
or \U$13824 ( \14201 , \14198 , \13599 );
nand \U$13825 ( \14202 , \14200 , \14201 );
xor \U$13826 ( \14203 , \13711 , \13717 );
xor \U$13827 ( \14204 , \14203 , \13724 );
and \U$13828 ( \14205 , \14202 , \14204 );
or \U$13829 ( \14206 , \13690 , \13688 );
nand \U$13830 ( \14207 , \14206 , \13691 );
xor \U$13831 ( \14208 , \13711 , \13717 );
xor \U$13832 ( \14209 , \14208 , \13724 );
and \U$13833 ( \14210 , \14207 , \14209 );
and \U$13834 ( \14211 , \14202 , \14207 );
or \U$13835 ( \14212 , \14205 , \14210 , \14211 );
not \U$13836 ( \14213 , \14212 );
xor \U$13837 ( \14214 , \13340 , \13342 );
xor \U$13838 ( \14215 , \14214 , \13345 );
and \U$13839 ( \14216 , \14213 , \14215 );
xor \U$13840 ( \14217 , \13356 , \13366 );
xor \U$13841 ( \14218 , \14217 , \13369 );
xor \U$13842 ( \14219 , \13340 , \13342 );
xor \U$13843 ( \14220 , \14219 , \13345 );
and \U$13844 ( \14221 , \14218 , \14220 );
and \U$13845 ( \14222 , \14213 , \14218 );
or \U$13846 ( \14223 , \14216 , \14221 , \14222 );
and \U$13847 ( \14224 , \14196 , \14223 );
and \U$13848 ( \14225 , \13829 , \14195 );
or \U$13849 ( \14226 , \14224 , \14225 );
not \U$13850 ( \14227 , \13209 );
not \U$13851 ( \14228 , \13267 );
or \U$13852 ( \14229 , \14227 , \14228 );
or \U$13853 ( \14230 , \13267 , \13209 );
nand \U$13854 ( \14231 , \14229 , \14230 );
not \U$13855 ( \14232 , \14231 );
not \U$13856 ( \14233 , \13247 );
and \U$13857 ( \14234 , \14232 , \14233 );
and \U$13858 ( \14235 , \14231 , \13247 );
nor \U$13859 ( \14236 , \14234 , \14235 );
xor \U$13860 ( \14237 , \13019 , \13105 );
xor \U$13861 ( \14238 , \14237 , \13189 );
xor \U$13862 ( \14239 , \14236 , \14238 );
xnor \U$13863 ( \14240 , \13327 , \13317 );
not \U$13864 ( \14241 , \14240 );
not \U$13865 ( \14242 , \13335 );
and \U$13866 ( \14243 , \14241 , \14242 );
and \U$13867 ( \14244 , \14240 , \13335 );
nor \U$13868 ( \14245 , \14243 , \14244 );
and \U$13869 ( \14246 , \14239 , \14245 );
and \U$13870 ( \14247 , \14236 , \14238 );
or \U$13871 ( \14248 , \14246 , \14247 );
xor \U$13872 ( \14249 , \14226 , \14248 );
xnor \U$13873 ( \14250 , \13299 , \12934 );
not \U$13874 ( \14251 , \14250 );
not \U$13875 ( \14252 , \13311 );
and \U$13876 ( \14253 , \14251 , \14252 );
and \U$13877 ( \14254 , \14250 , \13311 );
nor \U$13878 ( \14255 , \14253 , \14254 );
and \U$13879 ( \14256 , \14249 , \14255 );
and \U$13880 ( \14257 , \14226 , \14248 );
or \U$13881 ( \14258 , \14256 , \14257 );
nor \U$13882 ( \14259 , \13813 , \14258 );
nor \U$13883 ( \14260 , \13810 , \14259 );
not \U$13884 ( \14261 , \14260 );
and \U$13885 ( \14262 , \13805 , \14261 );
and \U$13886 ( \14263 , \13804 , \14260 );
nor \U$13887 ( \14264 , \14262 , \14263 );
not \U$13888 ( \14265 , \13634 );
not \U$13889 ( \14266 , \13729 );
or \U$13890 ( \14267 , \14265 , \14266 );
or \U$13891 ( \14268 , \13729 , \13634 );
nand \U$13892 ( \14269 , \14267 , \14268 );
not \U$13893 ( \14270 , \14269 );
not \U$13894 ( \14271 , \13654 );
and \U$13895 ( \14272 , \14270 , \14271 );
and \U$13896 ( \14273 , \14269 , \13654 );
nor \U$13897 ( \14274 , \14272 , \14273 );
xor \U$13898 ( \14275 , \14236 , \14238 );
xor \U$13899 ( \14276 , \14275 , \14245 );
and \U$13900 ( \14277 , \14274 , \14276 );
xor \U$13901 ( \14278 , \13829 , \14195 );
xor \U$13902 ( \14279 , \14278 , \14223 );
xor \U$13903 ( \14280 , \14236 , \14238 );
xor \U$13904 ( \14281 , \14280 , \14245 );
and \U$13905 ( \14282 , \14279 , \14281 );
and \U$13906 ( \14283 , \14274 , \14279 );
or \U$13907 ( \14284 , \14277 , \14282 , \14283 );
xnor \U$13908 ( \14285 , \13731 , \13374 );
not \U$13909 ( \14286 , \14285 );
not \U$13910 ( \14287 , \13337 );
and \U$13911 ( \14288 , \14286 , \14287 );
and \U$13912 ( \14289 , \14285 , \13337 );
nor \U$13913 ( \14290 , \14288 , \14289 );
xor \U$13914 ( \14291 , \14284 , \14290 );
xor \U$13915 ( \14292 , \14105 , \14131 );
xor \U$13916 ( \14293 , \14292 , \14157 );
xor \U$13917 ( \14294 , \14019 , \14044 );
xor \U$13918 ( \14295 , \14294 , \14076 );
and \U$13919 ( \14296 , \14293 , \14295 );
xor \U$13920 ( \14297 , \13938 , \13963 );
xor \U$13921 ( \14298 , \14297 , \13991 );
xor \U$13922 ( \14299 , \14019 , \14044 );
xor \U$13923 ( \14300 , \14299 , \14076 );
and \U$13924 ( \14301 , \14298 , \14300 );
and \U$13925 ( \14302 , \14293 , \14298 );
or \U$13926 ( \14303 , \14296 , \14301 , \14302 );
not \U$13927 ( \14304 , \13432 );
xor \U$13928 ( \14305 , \13464 , \13404 );
not \U$13929 ( \14306 , \14305 );
or \U$13930 ( \14307 , \14304 , \14306 );
or \U$13931 ( \14308 , \14305 , \13432 );
nand \U$13932 ( \14309 , \14307 , \14308 );
xor \U$13933 ( \14310 , \14303 , \14309 );
xor \U$13934 ( \14311 , \13853 , \13855 );
xor \U$13935 ( \14312 , \14311 , \13884 );
xor \U$13936 ( \14313 , \13894 , \13900 );
xor \U$13937 ( \14314 , \14313 , \13907 );
and \U$13938 ( \14315 , \14312 , \14314 );
xor \U$13939 ( \14316 , \13835 , \13841 );
xor \U$13940 ( \14317 , \14316 , \13848 );
xor \U$13941 ( \14318 , \13894 , \13900 );
xor \U$13942 ( \14319 , \14318 , \13907 );
and \U$13943 ( \14320 , \14317 , \14319 );
and \U$13944 ( \14321 , \14312 , \14317 );
or \U$13945 ( \14322 , \14315 , \14320 , \14321 );
and \U$13946 ( \14323 , \14310 , \14322 );
and \U$13947 ( \14324 , \14303 , \14309 );
or \U$13948 ( \14325 , \14323 , \14324 );
xor \U$13949 ( \14326 , \14052 , \14065 );
xor \U$13950 ( \14327 , \14326 , \14073 );
xor \U$13951 ( \14328 , \14026 , \14033 );
xor \U$13952 ( \14329 , \14328 , \14041 );
and \U$13953 ( \14330 , \14327 , \14329 );
xor \U$13954 ( \14331 , \14001 , \14008 );
xor \U$13955 ( \14332 , \14331 , \14016 );
xor \U$13956 ( \14333 , \14026 , \14033 );
xor \U$13957 ( \14334 , \14333 , \14041 );
and \U$13958 ( \14335 , \14332 , \14334 );
and \U$13959 ( \14336 , \14327 , \14332 );
or \U$13960 ( \14337 , \14330 , \14335 , \14336 );
xor \U$13961 ( \14338 , \13498 , \13502 );
xor \U$13962 ( \14339 , \14338 , \13510 );
xor \U$13963 ( \14340 , \14337 , \14339 );
xor \U$13964 ( \14341 , \13473 , \13480 );
xor \U$13965 ( \14342 , \14341 , \13488 );
xor \U$13966 ( \14343 , \14179 , \14184 );
xor \U$13967 ( \14344 , \14342 , \14343 );
and \U$13968 ( \14345 , \14340 , \14344 );
and \U$13969 ( \14346 , \14337 , \14339 );
or \U$13970 ( \14347 , \14345 , \14346 );
and \U$13971 ( \14348 , \2224 , RIae77c48_93);
and \U$13972 ( \14349 , RIae77b58_91, \2222 );
nor \U$13973 ( \14350 , \14348 , \14349 );
and \U$13974 ( \14351 , \14350 , \2061 );
not \U$13975 ( \14352 , \14350 );
and \U$13976 ( \14353 , \14352 , \2060 );
nor \U$13977 ( \14354 , \14351 , \14353 );
and \U$13978 ( \14355 , \2607 , RIae77d38_95);
and \U$13979 ( \14356 , RIae77e28_97, \2605 );
nor \U$13980 ( \14357 , \14355 , \14356 );
and \U$13981 ( \14358 , \14357 , \2611 );
not \U$13982 ( \14359 , \14357 );
and \U$13983 ( \14360 , \14359 , \2397 );
nor \U$13984 ( \14361 , \14358 , \14360 );
xor \U$13985 ( \14362 , \14354 , \14361 );
not \U$13986 ( \14363 , \3089 );
and \U$13987 ( \14364 , \2783 , RIae78968_121);
and \U$13988 ( \14365 , RIae78878_119, \2781 );
nor \U$13989 ( \14366 , \14364 , \14365 );
not \U$13990 ( \14367 , \14366 );
or \U$13991 ( \14368 , \14363 , \14367 );
or \U$13992 ( \14369 , \14366 , \3089 );
nand \U$13993 ( \14370 , \14368 , \14369 );
and \U$13994 ( \14371 , \14362 , \14370 );
and \U$13995 ( \14372 , \14354 , \14361 );
or \U$13996 ( \14373 , \14371 , \14372 );
and \U$13997 ( \14374 , \1939 , RIae783c8_109);
and \U$13998 ( \14375 , RIae78530_112, \1937 );
nor \U$13999 ( \14376 , \14374 , \14375 );
and \U$14000 ( \14377 , \14376 , \1735 );
not \U$14001 ( \14378 , \14376 );
and \U$14002 ( \14379 , \14378 , \1734 );
nor \U$14003 ( \14380 , \14377 , \14379 );
and \U$14004 ( \14381 , \1376 , RIae77f18_99);
and \U$14005 ( \14382 , RIae78008_101, \1374 );
nor \U$14006 ( \14383 , \14381 , \14382 );
and \U$14007 ( \14384 , \14383 , \1380 );
not \U$14008 ( \14385 , \14383 );
and \U$14009 ( \14386 , \14385 , \1261 );
nor \U$14010 ( \14387 , \14384 , \14386 );
xor \U$14011 ( \14388 , \14380 , \14387 );
and \U$14012 ( \14389 , \1593 , RIae781e8_105);
and \U$14013 ( \14390 , RIae785a8_113, \1591 );
nor \U$14014 ( \14391 , \14389 , \14390 );
and \U$14015 ( \14392 , \14391 , \1498 );
not \U$14016 ( \14393 , \14391 );
and \U$14017 ( \14394 , \14393 , \1488 );
nor \U$14018 ( \14395 , \14392 , \14394 );
and \U$14019 ( \14396 , \14388 , \14395 );
and \U$14020 ( \14397 , \14380 , \14387 );
or \U$14021 ( \14398 , \14396 , \14397 );
xor \U$14022 ( \14399 , \14373 , \14398 );
and \U$14023 ( \14400 , \672 , RIae77180_70);
and \U$14024 ( \14401 , RIae77018_67, \670 );
nor \U$14025 ( \14402 , \14400 , \14401 );
and \U$14026 ( \14403 , \14402 , \588 );
not \U$14027 ( \14404 , \14402 );
and \U$14028 ( \14405 , \14404 , \587 );
nor \U$14029 ( \14406 , \14403 , \14405 );
not \U$14030 ( \14407 , \787 );
and \U$14031 ( \14408 , \883 , RIae771f8_71);
and \U$14032 ( \14409 , RIae772e8_73, \881 );
nor \U$14033 ( \14410 , \14408 , \14409 );
not \U$14034 ( \14411 , \14410 );
or \U$14035 ( \14412 , \14407 , \14411 );
or \U$14036 ( \14413 , \14410 , \789 );
nand \U$14037 ( \14414 , \14412 , \14413 );
xor \U$14038 ( \14415 , \14406 , \14414 );
and \U$14039 ( \14416 , \1138 , RIae782d8_107);
and \U$14040 ( \14417 , RIae780f8_103, \1136 );
nor \U$14041 ( \14418 , \14416 , \14417 );
and \U$14042 ( \14419 , \14418 , \1012 );
not \U$14043 ( \14420 , \14418 );
and \U$14044 ( \14421 , \14420 , \1142 );
nor \U$14045 ( \14422 , \14419 , \14421 );
and \U$14046 ( \14423 , \14415 , \14422 );
and \U$14047 ( \14424 , \14406 , \14414 );
or \U$14048 ( \14425 , \14423 , \14424 );
and \U$14049 ( \14426 , \14399 , \14425 );
and \U$14050 ( \14427 , \14373 , \14398 );
or \U$14051 ( \14428 , \14426 , \14427 );
and \U$14052 ( \14429 , \12180 , RIae767a8_49);
and \U$14053 ( \14430 , RIae76898_51, \12178 );
nor \U$14054 ( \14431 , \14429 , \14430 );
and \U$14055 ( \14432 , \14431 , \12184 );
not \U$14056 ( \14433 , \14431 );
and \U$14057 ( \14434 , \14433 , \11827 );
nor \U$14058 ( \14435 , \14432 , \14434 );
and \U$14059 ( \14436 , \10548 , RIae762f8_39);
and \U$14060 ( \14437 , RIae76208_37, \10546 );
nor \U$14061 ( \14438 , \14436 , \14437 );
and \U$14062 ( \14439 , \14438 , \10421 );
not \U$14063 ( \14440 , \14438 );
and \U$14064 ( \14441 , \14440 , \10118 );
nor \U$14065 ( \14442 , \14439 , \14441 );
xor \U$14066 ( \14443 , \14435 , \14442 );
and \U$14067 ( \14444 , \11470 , RIae76a78_55);
and \U$14068 ( \14445 , RIae76988_53, \11468 );
nor \U$14069 ( \14446 , \14444 , \14445 );
and \U$14070 ( \14447 , \14446 , \10936 );
not \U$14071 ( \14448 , \14446 );
and \U$14072 ( \14449 , \14448 , \11474 );
nor \U$14073 ( \14450 , \14447 , \14449 );
and \U$14074 ( \14451 , \14443 , \14450 );
and \U$14075 ( \14452 , \14435 , \14442 );
or \U$14076 ( \14453 , \14451 , \14452 );
and \U$14077 ( \14454 , \13059 , RIae76b68_57);
and \U$14078 ( \14455 , RIae78a58_123, \13057 );
nor \U$14079 ( \14456 , \14454 , \14455 );
and \U$14080 ( \14457 , \14456 , \13063 );
not \U$14081 ( \14458 , \14456 );
and \U$14082 ( \14459 , \14458 , \12718 );
nor \U$14083 ( \14460 , \14457 , \14459 );
nand \U$14084 ( \14461 , RIae7aa38_191, RIae7a9c0_190);
and \U$14085 ( \14462 , \14461 , RIae7a8d0_188);
not \U$14086 ( \14463 , \14462 );
xor \U$14087 ( \14464 , \14460 , \14463 );
and \U$14088 ( \14465 , \14059 , RIae78cb0_128);
and \U$14089 ( \14466 , RIae78da0_130, \14057 );
nor \U$14090 ( \14467 , \14465 , \14466 );
and \U$14091 ( \14468 , \14467 , \13502 );
not \U$14092 ( \14469 , \14467 );
and \U$14093 ( \14470 , \14469 , \14063 );
nor \U$14094 ( \14471 , \14468 , \14470 );
and \U$14095 ( \14472 , \14464 , \14471 );
and \U$14096 ( \14473 , \14460 , \14463 );
or \U$14097 ( \14474 , \14472 , \14473 );
xor \U$14098 ( \14475 , \14453 , \14474 );
and \U$14099 ( \14476 , \8966 , RIae766b8_47);
and \U$14100 ( \14477 , RIae765c8_45, \8964 );
nor \U$14101 ( \14478 , \14476 , \14477 );
and \U$14102 ( \14479 , \14478 , \8799 );
not \U$14103 ( \14480 , \14478 );
and \U$14104 ( \14481 , \14480 , \8789 );
nor \U$14105 ( \14482 , \14479 , \14481 );
and \U$14106 ( \14483 , \8371 , RIae763e8_41);
and \U$14107 ( \14484 , RIae764d8_43, \8369 );
nor \U$14108 ( \14485 , \14483 , \14484 );
and \U$14109 ( \14486 , \14485 , \8020 );
not \U$14110 ( \14487 , \14485 );
and \U$14111 ( \14488 , \14487 , \8019 );
nor \U$14112 ( \14489 , \14486 , \14488 );
xor \U$14113 ( \14490 , \14482 , \14489 );
and \U$14114 ( \14491 , \9760 , RIae76118_35);
and \U$14115 ( \14492 , RIae76028_33, \9758 );
nor \U$14116 ( \14493 , \14491 , \14492 );
and \U$14117 ( \14494 , \14493 , \9273 );
not \U$14118 ( \14495 , \14493 );
and \U$14119 ( \14496 , \14495 , \9272 );
nor \U$14120 ( \14497 , \14494 , \14496 );
and \U$14121 ( \14498 , \14490 , \14497 );
and \U$14122 ( \14499 , \14482 , \14489 );
or \U$14123 ( \14500 , \14498 , \14499 );
and \U$14124 ( \14501 , \14475 , \14500 );
and \U$14125 ( \14502 , \14453 , \14474 );
or \U$14126 ( \14503 , \14501 , \14502 );
xor \U$14127 ( \14504 , \14428 , \14503 );
and \U$14128 ( \14505 , \5896 , RIae755d8_11);
and \U$14129 ( \14506 , RIae754e8_9, \5894 );
nor \U$14130 ( \14507 , \14505 , \14506 );
and \U$14131 ( \14508 , \14507 , \5590 );
not \U$14132 ( \14509 , \14507 );
and \U$14133 ( \14510 , \14509 , \5589 );
nor \U$14134 ( \14511 , \14508 , \14510 );
and \U$14135 ( \14512 , \4688 , RIae75f38_31);
and \U$14136 ( \14513 , RIae75e48_29, \4686 );
nor \U$14137 ( \14514 , \14512 , \14513 );
and \U$14138 ( \14515 , \14514 , \4481 );
not \U$14139 ( \14516 , \14514 );
and \U$14140 ( \14517 , \14516 , \4482 );
nor \U$14141 ( \14518 , \14515 , \14517 );
xor \U$14142 ( \14519 , \14511 , \14518 );
and \U$14143 ( \14520 , \5399 , RIae75c68_25);
and \U$14144 ( \14521 , RIae75d58_27, \5397 );
nor \U$14145 ( \14522 , \14520 , \14521 );
and \U$14146 ( \14523 , \14522 , \5016 );
not \U$14147 ( \14524 , \14522 );
and \U$14148 ( \14525 , \14524 , \5403 );
nor \U$14149 ( \14526 , \14523 , \14525 );
and \U$14150 ( \14527 , \14519 , \14526 );
and \U$14151 ( \14528 , \14511 , \14518 );
or \U$14152 ( \14529 , \14527 , \14528 );
and \U$14153 ( \14530 , \4247 , RIae75998_19);
and \U$14154 ( \14531 , RIae758a8_17, \4245 );
nor \U$14155 ( \14532 , \14530 , \14531 );
and \U$14156 ( \14533 , \14532 , \3989 );
not \U$14157 ( \14534 , \14532 );
and \U$14158 ( \14535 , \14534 , \4251 );
nor \U$14159 ( \14536 , \14533 , \14535 );
not \U$14160 ( \14537 , \2774 );
and \U$14161 ( \14538 , \3214 , RIae78788_117);
and \U$14162 ( \14539 , RIae78698_115, \3212 );
nor \U$14163 ( \14540 , \14538 , \14539 );
not \U$14164 ( \14541 , \14540 );
or \U$14165 ( \14542 , \14537 , \14541 );
or \U$14166 ( \14543 , \14540 , \3218 );
nand \U$14167 ( \14544 , \14542 , \14543 );
xor \U$14168 ( \14545 , \14536 , \14544 );
and \U$14169 ( \14546 , \3730 , RIae75b78_23);
and \U$14170 ( \14547 , RIae75a88_21, \3728 );
nor \U$14171 ( \14548 , \14546 , \14547 );
and \U$14172 ( \14549 , \14548 , \3732 );
not \U$14173 ( \14550 , \14548 );
and \U$14174 ( \14551 , \14550 , \3422 );
nor \U$14175 ( \14552 , \14549 , \14551 );
and \U$14176 ( \14553 , \14545 , \14552 );
and \U$14177 ( \14554 , \14536 , \14544 );
or \U$14178 ( \14555 , \14553 , \14554 );
xor \U$14179 ( \14556 , \14529 , \14555 );
and \U$14180 ( \14557 , \7633 , RIae75308_5);
and \U$14181 ( \14558 , RIae753f8_7, \7631 );
nor \U$14182 ( \14559 , \14557 , \14558 );
and \U$14183 ( \14560 , \14559 , \7206 );
not \U$14184 ( \14561 , \14559 );
and \U$14185 ( \14562 , \14561 , \7205 );
nor \U$14186 ( \14563 , \14560 , \14562 );
and \U$14187 ( \14564 , \6172 , RIae757b8_15);
and \U$14188 ( \14565 , RIae756c8_13, \6170 );
nor \U$14189 ( \14566 , \14564 , \14565 );
and \U$14190 ( \14567 , \14566 , \6176 );
not \U$14191 ( \14568 , \14566 );
and \U$14192 ( \14569 , \14568 , \6175 );
nor \U$14193 ( \14570 , \14567 , \14569 );
xor \U$14194 ( \14571 , \14563 , \14570 );
and \U$14195 ( \14572 , \6941 , RIae75218_3);
and \U$14196 ( \14573 , RIae75128_1, \6939 );
nor \U$14197 ( \14574 , \14572 , \14573 );
and \U$14198 ( \14575 , \14574 , \6314 );
not \U$14199 ( \14576 , \14574 );
and \U$14200 ( \14577 , \14576 , \6945 );
nor \U$14201 ( \14578 , \14575 , \14577 );
and \U$14202 ( \14579 , \14571 , \14578 );
and \U$14203 ( \14580 , \14563 , \14570 );
or \U$14204 ( \14581 , \14579 , \14580 );
and \U$14205 ( \14582 , \14556 , \14581 );
and \U$14206 ( \14583 , \14529 , \14555 );
or \U$14207 ( \14584 , \14582 , \14583 );
and \U$14208 ( \14585 , \14504 , \14584 );
and \U$14209 ( \14586 , \14428 , \14503 );
or \U$14210 ( \14587 , \14585 , \14586 );
xor \U$14211 ( \14588 , \14347 , \14587 );
xor \U$14212 ( \14589 , \14087 , \14094 );
xor \U$14213 ( \14590 , \14589 , \14102 );
xor \U$14214 ( \14591 , \14112 , \14119 );
xor \U$14215 ( \14592 , \14591 , \14128 );
and \U$14216 ( \14593 , \14590 , \14592 );
xor \U$14217 ( \14594 , \14139 , \14146 );
xor \U$14218 ( \14595 , \14594 , \14154 );
xor \U$14219 ( \14596 , \14112 , \14119 );
xor \U$14220 ( \14597 , \14596 , \14128 );
and \U$14221 ( \14598 , \14595 , \14597 );
and \U$14222 ( \14599 , \14590 , \14595 );
or \U$14223 ( \14600 , \14593 , \14598 , \14599 );
not \U$14224 ( \14601 , \402 );
and \U$14225 ( \14602 , \436 , RIae77798_83);
and \U$14226 ( \14603 , RIae77888_85, \434 );
nor \U$14227 ( \14604 , \14602 , \14603 );
not \U$14228 ( \14605 , \14604 );
or \U$14229 ( \14606 , \14601 , \14605 );
or \U$14230 ( \14607 , \14604 , \400 );
nand \U$14231 ( \14608 , \14606 , \14607 );
not \U$14232 ( \14609 , \469 );
and \U$14233 ( \14610 , \514 , RIae76f28_65);
and \U$14234 ( \14611 , RIae76e38_63, \512 );
nor \U$14235 ( \14612 , \14610 , \14611 );
not \U$14236 ( \14613 , \14612 );
or \U$14237 ( \14614 , \14609 , \14613 );
or \U$14238 ( \14615 , \14612 , \471 );
nand \U$14239 ( \14616 , \14614 , \14615 );
xor \U$14240 ( \14617 , \14608 , \14616 );
and \U$14241 ( \14618 , \558 , RIae76d48_61);
and \U$14242 ( \14619 , RIae76c58_59, \556 );
nor \U$14243 ( \14620 , \14618 , \14619 );
and \U$14244 ( \14621 , \14620 , \504 );
not \U$14245 ( \14622 , \14620 );
and \U$14246 ( \14623 , \14622 , \562 );
nor \U$14247 ( \14624 , \14621 , \14623 );
and \U$14248 ( \14625 , \14617 , \14624 );
and \U$14249 ( \14626 , \14608 , \14616 );
or \U$14250 ( \14627 , \14625 , \14626 );
xor \U$14251 ( \14628 , \14627 , \13852 );
xor \U$14252 ( \14629 , \13864 , \13872 );
xor \U$14253 ( \14630 , \14629 , \13881 );
and \U$14254 ( \14631 , \14628 , \14630 );
and \U$14255 ( \14632 , \14627 , \13852 );
or \U$14256 ( \14633 , \14631 , \14632 );
xor \U$14257 ( \14634 , \14600 , \14633 );
xor \U$14258 ( \14635 , \13972 , \13980 );
xor \U$14259 ( \14636 , \14635 , \13988 );
xor \U$14260 ( \14637 , \13945 , \13952 );
xor \U$14261 ( \14638 , \14637 , \13960 );
and \U$14262 ( \14639 , \14636 , \14638 );
xor \U$14263 ( \14640 , \13920 , \13927 );
xor \U$14264 ( \14641 , \14640 , \13935 );
xor \U$14265 ( \14642 , \13945 , \13952 );
xor \U$14266 ( \14643 , \14642 , \13960 );
and \U$14267 ( \14644 , \14641 , \14643 );
and \U$14268 ( \14645 , \14636 , \14641 );
or \U$14269 ( \14646 , \14639 , \14644 , \14645 );
and \U$14270 ( \14647 , \14634 , \14646 );
and \U$14271 ( \14648 , \14600 , \14633 );
or \U$14272 ( \14649 , \14647 , \14648 );
and \U$14273 ( \14650 , \14588 , \14649 );
and \U$14274 ( \14651 , \14347 , \14587 );
or \U$14275 ( \14652 , \14650 , \14651 );
and \U$14276 ( \14653 , \14325 , \14652 );
xor \U$14277 ( \14654 , \13711 , \13717 );
xor \U$14278 ( \14655 , \14654 , \13724 );
xor \U$14279 ( \14656 , \14202 , \14207 );
xor \U$14280 ( \14657 , \14655 , \14656 );
xor \U$14281 ( \14658 , \13491 , \13513 );
xor \U$14282 ( \14659 , \14658 , \13539 );
xor \U$14283 ( \14660 , \14657 , \14659 );
xor \U$14284 ( \14661 , \14170 , \14172 );
xor \U$14285 ( \14662 , \14661 , \14189 );
and \U$14286 ( \14663 , \14660 , \14662 );
and \U$14287 ( \14664 , \14657 , \14659 );
or \U$14288 ( \14665 , \14663 , \14664 );
or \U$14289 ( \14666 , \14325 , \14652 );
and \U$14290 ( \14667 , \14665 , \14666 );
nor \U$14291 ( \14668 , \14653 , \14667 );
not \U$14292 ( \14669 , \13348 );
not \U$14293 ( \14670 , \13372 );
or \U$14294 ( \14671 , \14669 , \14670 );
or \U$14295 ( \14672 , \13348 , \13372 );
nand \U$14296 ( \14673 , \14671 , \14672 );
not \U$14297 ( \14674 , \14673 );
not \U$14298 ( \14675 , \13350 );
and \U$14299 ( \14676 , \14674 , \14675 );
and \U$14300 ( \14677 , \14673 , \13350 );
nor \U$14301 ( \14678 , \14676 , \14677 );
xor \U$14302 ( \14679 , \14668 , \14678 );
xor \U$14303 ( \14680 , \13340 , \13342 );
xor \U$14304 ( \14681 , \14680 , \13345 );
xor \U$14305 ( \14682 , \14213 , \14218 );
xor \U$14306 ( \14683 , \14681 , \14682 );
not \U$14307 ( \14684 , \14683 );
xor \U$14308 ( \14685 , \13913 , \14163 );
xor \U$14309 ( \14686 , \14685 , \14192 );
not \U$14310 ( \14687 , \14686 );
and \U$14311 ( \14688 , \14684 , \14687 );
and \U$14312 ( \14689 , \14683 , \14686 );
xor \U$14313 ( \14690 , \13636 , \13638 );
xor \U$14314 ( \14691 , \14690 , \13651 );
xor \U$14315 ( \14692 , \13815 , \13824 );
xor \U$14316 ( \14693 , \14691 , \14692 );
nor \U$14317 ( \14694 , \14689 , \14693 );
nor \U$14318 ( \14695 , \14688 , \14694 );
and \U$14319 ( \14696 , \14679 , \14695 );
and \U$14320 ( \14697 , \14668 , \14678 );
or \U$14321 ( \14698 , \14696 , \14697 );
and \U$14322 ( \14699 , \14291 , \14698 );
and \U$14323 ( \14700 , \14284 , \14290 );
or \U$14324 ( \14701 , \14699 , \14700 );
not \U$14325 ( \14702 , \14701 );
not \U$14326 ( \14703 , \13807 );
not \U$14327 ( \14704 , \14258 );
not \U$14328 ( \14705 , \13809 );
and \U$14329 ( \14706 , \14704 , \14705 );
and \U$14330 ( \14707 , \14258 , \13809 );
nor \U$14331 ( \14708 , \14706 , \14707 );
not \U$14332 ( \14709 , \14708 );
or \U$14333 ( \14710 , \14703 , \14709 );
or \U$14334 ( \14711 , \14708 , \13807 );
nand \U$14335 ( \14712 , \14710 , \14711 );
nand \U$14336 ( \14713 , \14702 , \14712 );
or \U$14337 ( \14714 , \14264 , \14713 );
xnor \U$14338 ( \14715 , \14713 , \14264 );
xor \U$14339 ( \14716 , \14284 , \14290 );
xor \U$14340 ( \14717 , \14716 , \14698 );
xor \U$14341 ( \14718 , \14226 , \14248 );
xor \U$14342 ( \14719 , \14718 , \14255 );
or \U$14343 ( \14720 , \14717 , \14719 );
not \U$14344 ( \14721 , \14719 );
not \U$14345 ( \14722 , \14717 );
or \U$14346 ( \14723 , \14721 , \14722 );
xor \U$14347 ( \14724 , \14668 , \14678 );
xor \U$14348 ( \14725 , \14724 , \14695 );
xor \U$14349 ( \14726 , \14236 , \14238 );
xor \U$14350 ( \14727 , \14726 , \14245 );
xor \U$14351 ( \14728 , \14274 , \14279 );
xor \U$14352 ( \14729 , \14727 , \14728 );
or \U$14353 ( \14730 , \14725 , \14729 );
not \U$14354 ( \14731 , \14729 );
not \U$14355 ( \14732 , \14725 );
or \U$14356 ( \14733 , \14731 , \14732 );
xor \U$14357 ( \14734 , \14112 , \14119 );
xor \U$14358 ( \14735 , \14734 , \14128 );
xor \U$14359 ( \14736 , \14590 , \14595 );
xor \U$14360 ( \14737 , \14735 , \14736 );
xor \U$14361 ( \14738 , \14627 , \13852 );
xor \U$14362 ( \14739 , \14738 , \14630 );
and \U$14363 ( \14740 , \14737 , \14739 );
xor \U$14364 ( \14741 , \13945 , \13952 );
xor \U$14365 ( \14742 , \14741 , \13960 );
xor \U$14366 ( \14743 , \14636 , \14641 );
xor \U$14367 ( \14744 , \14742 , \14743 );
xor \U$14368 ( \14745 , \14627 , \13852 );
xor \U$14369 ( \14746 , \14745 , \14630 );
and \U$14370 ( \14747 , \14744 , \14746 );
and \U$14371 ( \14748 , \14737 , \14744 );
or \U$14372 ( \14749 , \14740 , \14747 , \14748 );
xor \U$14373 ( \14750 , \14453 , \14474 );
xor \U$14374 ( \14751 , \14750 , \14500 );
xor \U$14375 ( \14752 , \14529 , \14555 );
xor \U$14376 ( \14753 , \14752 , \14581 );
and \U$14377 ( \14754 , \14751 , \14753 );
xor \U$14378 ( \14755 , \14373 , \14398 );
xor \U$14379 ( \14756 , \14755 , \14425 );
xor \U$14380 ( \14757 , \14529 , \14555 );
xor \U$14381 ( \14758 , \14757 , \14581 );
and \U$14382 ( \14759 , \14756 , \14758 );
and \U$14383 ( \14760 , \14751 , \14756 );
or \U$14384 ( \14761 , \14754 , \14759 , \14760 );
xor \U$14385 ( \14762 , \14749 , \14761 );
xor \U$14386 ( \14763 , \14019 , \14044 );
xor \U$14387 ( \14764 , \14763 , \14076 );
xor \U$14388 ( \14765 , \14293 , \14298 );
xor \U$14389 ( \14766 , \14764 , \14765 );
and \U$14390 ( \14767 , \14762 , \14766 );
and \U$14391 ( \14768 , \14749 , \14761 );
or \U$14392 ( \14769 , \14767 , \14768 );
not \U$14393 ( \14770 , RIae773d8_75);
nor \U$14394 ( \14771 , \14770 , \491 );
xor \U$14395 ( \14772 , \14608 , \14616 );
xor \U$14396 ( \14773 , \14772 , \14624 );
and \U$14397 ( \14774 , \14771 , \14773 );
xor \U$14398 ( \14775 , \14406 , \14414 );
xor \U$14399 ( \14776 , \14775 , \14422 );
xor \U$14400 ( \14777 , \14608 , \14616 );
xor \U$14401 ( \14778 , \14777 , \14624 );
and \U$14402 ( \14779 , \14776 , \14778 );
and \U$14403 ( \14780 , \14771 , \14776 );
or \U$14404 ( \14781 , \14774 , \14779 , \14780 );
nand \U$14405 ( \14782 , RIae77720_82, RIae78b48_125);
and \U$14406 ( \14783 , \384 , RIae773d8_75);
and \U$14407 ( \14784 , RIae77a68_89, \382 );
nor \U$14408 ( \14785 , \14783 , \14784 );
not \U$14409 ( \14786 , \14785 );
not \U$14410 ( \14787 , \388 );
and \U$14411 ( \14788 , \14786 , \14787 );
and \U$14412 ( \14789 , \14785 , \388 );
nor \U$14413 ( \14790 , \14788 , \14789 );
nand \U$14414 ( \14791 , \14782 , \14790 );
not \U$14415 ( \14792 , \388 );
and \U$14416 ( \14793 , \384 , RIae77a68_89);
and \U$14417 ( \14794 , RIae77978_87, \382 );
nor \U$14418 ( \14795 , \14793 , \14794 );
not \U$14419 ( \14796 , \14795 );
or \U$14420 ( \14797 , \14792 , \14796 );
or \U$14421 ( \14798 , \14795 , \392 );
nand \U$14422 ( \14799 , \14797 , \14798 );
xor \U$14423 ( \14800 , \14791 , \14799 );
not \U$14424 ( \14801 , \402 );
and \U$14425 ( \14802 , \436 , RIae77978_87);
and \U$14426 ( \14803 , RIae77798_83, \434 );
nor \U$14427 ( \14804 , \14802 , \14803 );
not \U$14428 ( \14805 , \14804 );
or \U$14429 ( \14806 , \14801 , \14805 );
or \U$14430 ( \14807 , \14804 , \402 );
nand \U$14431 ( \14808 , \14806 , \14807 );
not \U$14432 ( \14809 , \469 );
and \U$14433 ( \14810 , \514 , RIae77888_85);
and \U$14434 ( \14811 , RIae76f28_65, \512 );
nor \U$14435 ( \14812 , \14810 , \14811 );
not \U$14436 ( \14813 , \14812 );
or \U$14437 ( \14814 , \14809 , \14813 );
or \U$14438 ( \14815 , \14812 , \469 );
nand \U$14439 ( \14816 , \14814 , \14815 );
xor \U$14440 ( \14817 , \14808 , \14816 );
and \U$14441 ( \14818 , \558 , RIae76e38_63);
and \U$14442 ( \14819 , RIae76d48_61, \556 );
nor \U$14443 ( \14820 , \14818 , \14819 );
and \U$14444 ( \14821 , \14820 , \504 );
not \U$14445 ( \14822 , \14820 );
and \U$14446 ( \14823 , \14822 , \562 );
nor \U$14447 ( \14824 , \14821 , \14823 );
and \U$14448 ( \14825 , \14817 , \14824 );
and \U$14449 ( \14826 , \14808 , \14816 );
or \U$14450 ( \14827 , \14825 , \14826 );
and \U$14451 ( \14828 , \14800 , \14827 );
and \U$14452 ( \14829 , \14791 , \14799 );
or \U$14453 ( \14830 , \14828 , \14829 );
xor \U$14454 ( \14831 , \14781 , \14830 );
xor \U$14455 ( \14832 , \14380 , \14387 );
xor \U$14456 ( \14833 , \14832 , \14395 );
xor \U$14457 ( \14834 , \14354 , \14361 );
xor \U$14458 ( \14835 , \14834 , \14370 );
xor \U$14459 ( \14836 , \14833 , \14835 );
xor \U$14460 ( \14837 , \14536 , \14544 );
xor \U$14461 ( \14838 , \14837 , \14552 );
and \U$14462 ( \14839 , \14836 , \14838 );
and \U$14463 ( \14840 , \14833 , \14835 );
or \U$14464 ( \14841 , \14839 , \14840 );
and \U$14465 ( \14842 , \14831 , \14841 );
and \U$14466 ( \14843 , \14781 , \14830 );
or \U$14467 ( \14844 , \14842 , \14843 );
and \U$14468 ( \14845 , \1376 , RIae780f8_103);
and \U$14469 ( \14846 , RIae77f18_99, \1374 );
nor \U$14470 ( \14847 , \14845 , \14846 );
and \U$14471 ( \14848 , \14847 , \1380 );
not \U$14472 ( \14849 , \14847 );
and \U$14473 ( \14850 , \14849 , \1261 );
nor \U$14474 ( \14851 , \14848 , \14850 );
and \U$14475 ( \14852 , \1593 , RIae78008_101);
and \U$14476 ( \14853 , RIae781e8_105, \1591 );
nor \U$14477 ( \14854 , \14852 , \14853 );
and \U$14478 ( \14855 , \14854 , \1498 );
not \U$14479 ( \14856 , \14854 );
and \U$14480 ( \14857 , \14856 , \1488 );
nor \U$14481 ( \14858 , \14855 , \14857 );
xor \U$14482 ( \14859 , \14851 , \14858 );
and \U$14483 ( \14860 , \1939 , RIae785a8_113);
and \U$14484 ( \14861 , RIae783c8_109, \1937 );
nor \U$14485 ( \14862 , \14860 , \14861 );
and \U$14486 ( \14863 , \14862 , \1735 );
not \U$14487 ( \14864 , \14862 );
and \U$14488 ( \14865 , \14864 , \1734 );
nor \U$14489 ( \14866 , \14863 , \14865 );
and \U$14490 ( \14867 , \14859 , \14866 );
and \U$14491 ( \14868 , \14851 , \14858 );
or \U$14492 ( \14869 , \14867 , \14868 );
and \U$14493 ( \14870 , \1138 , RIae772e8_73);
and \U$14494 ( \14871 , RIae782d8_107, \1136 );
nor \U$14495 ( \14872 , \14870 , \14871 );
and \U$14496 ( \14873 , \14872 , \1012 );
not \U$14497 ( \14874 , \14872 );
and \U$14498 ( \14875 , \14874 , \1142 );
nor \U$14499 ( \14876 , \14873 , \14875 );
and \U$14500 ( \14877 , \672 , RIae76c58_59);
and \U$14501 ( \14878 , RIae77180_70, \670 );
nor \U$14502 ( \14879 , \14877 , \14878 );
and \U$14503 ( \14880 , \14879 , \588 );
not \U$14504 ( \14881 , \14879 );
and \U$14505 ( \14882 , \14881 , \587 );
nor \U$14506 ( \14883 , \14880 , \14882 );
xor \U$14507 ( \14884 , \14876 , \14883 );
not \U$14508 ( \14885 , \787 );
and \U$14509 ( \14886 , \883 , RIae77018_67);
and \U$14510 ( \14887 , RIae771f8_71, \881 );
nor \U$14511 ( \14888 , \14886 , \14887 );
not \U$14512 ( \14889 , \14888 );
or \U$14513 ( \14890 , \14885 , \14889 );
or \U$14514 ( \14891 , \14888 , \787 );
nand \U$14515 ( \14892 , \14890 , \14891 );
and \U$14516 ( \14893 , \14884 , \14892 );
and \U$14517 ( \14894 , \14876 , \14883 );
or \U$14518 ( \14895 , \14893 , \14894 );
xor \U$14519 ( \14896 , \14869 , \14895 );
and \U$14520 ( \14897 , \2607 , RIae77b58_91);
and \U$14521 ( \14898 , RIae77d38_95, \2605 );
nor \U$14522 ( \14899 , \14897 , \14898 );
and \U$14523 ( \14900 , \14899 , \2611 );
not \U$14524 ( \14901 , \14899 );
and \U$14525 ( \14902 , \14901 , \2397 );
nor \U$14526 ( \14903 , \14900 , \14902 );
and \U$14527 ( \14904 , \2224 , RIae78530_112);
and \U$14528 ( \14905 , RIae77c48_93, \2222 );
nor \U$14529 ( \14906 , \14904 , \14905 );
and \U$14530 ( \14907 , \14906 , \2061 );
not \U$14531 ( \14908 , \14906 );
and \U$14532 ( \14909 , \14908 , \2060 );
nor \U$14533 ( \14910 , \14907 , \14909 );
xor \U$14534 ( \14911 , \14903 , \14910 );
not \U$14535 ( \14912 , \3089 );
and \U$14536 ( \14913 , \2783 , RIae77e28_97);
and \U$14537 ( \14914 , RIae78968_121, \2781 );
nor \U$14538 ( \14915 , \14913 , \14914 );
not \U$14539 ( \14916 , \14915 );
or \U$14540 ( \14917 , \14912 , \14916 );
or \U$14541 ( \14918 , \14915 , \3089 );
nand \U$14542 ( \14919 , \14917 , \14918 );
and \U$14543 ( \14920 , \14911 , \14919 );
and \U$14544 ( \14921 , \14903 , \14910 );
or \U$14545 ( \14922 , \14920 , \14921 );
and \U$14546 ( \14923 , \14896 , \14922 );
and \U$14547 ( \14924 , \14869 , \14895 );
or \U$14548 ( \14925 , \14923 , \14924 );
and \U$14549 ( \14926 , \8371 , RIae753f8_7);
and \U$14550 ( \14927 , RIae763e8_41, \8369 );
nor \U$14551 ( \14928 , \14926 , \14927 );
and \U$14552 ( \14929 , \14928 , \8020 );
not \U$14553 ( \14930 , \14928 );
and \U$14554 ( \14931 , \14930 , \8019 );
nor \U$14555 ( \14932 , \14929 , \14931 );
and \U$14556 ( \14933 , \8966 , RIae764d8_43);
and \U$14557 ( \14934 , RIae766b8_47, \8964 );
nor \U$14558 ( \14935 , \14933 , \14934 );
and \U$14559 ( \14936 , \14935 , \8799 );
not \U$14560 ( \14937 , \14935 );
and \U$14561 ( \14938 , \14937 , \8789 );
nor \U$14562 ( \14939 , \14936 , \14938 );
xor \U$14563 ( \14940 , \14932 , \14939 );
and \U$14564 ( \14941 , \9760 , RIae765c8_45);
and \U$14565 ( \14942 , RIae76118_35, \9758 );
nor \U$14566 ( \14943 , \14941 , \14942 );
and \U$14567 ( \14944 , \14943 , \9273 );
not \U$14568 ( \14945 , \14943 );
and \U$14569 ( \14946 , \14945 , \9272 );
nor \U$14570 ( \14947 , \14944 , \14946 );
and \U$14571 ( \14948 , \14940 , \14947 );
and \U$14572 ( \14949 , \14932 , \14939 );
or \U$14573 ( \14950 , \14948 , \14949 );
and \U$14574 ( \14951 , \13059 , RIae76898_51);
and \U$14575 ( \14952 , RIae76b68_57, \13057 );
nor \U$14576 ( \14953 , \14951 , \14952 );
and \U$14577 ( \14954 , \14953 , \13063 );
not \U$14578 ( \14955 , \14953 );
and \U$14579 ( \14956 , \14955 , \12718 );
nor \U$14580 ( \14957 , \14954 , \14956 );
and \U$14581 ( \14958 , RIae7a8d0_188, RIae7a9c0_190);
not \U$14582 ( \14959 , RIae7aa38_191);
and \U$14583 ( \14960 , \14959 , RIae7a9c0_190);
nor \U$14584 ( \14961 , \14959 , RIae7a9c0_190);
or \U$14585 ( \14962 , \14960 , \14961 );
nor \U$14586 ( \14963 , RIae7a8d0_188, RIae7a9c0_190);
nor \U$14587 ( \14964 , \14958 , \14962 , \14963 );
nand \U$14588 ( \14965 , RIae78da0_130, \14964 );
and \U$14589 ( \14966 , \14965 , \14463 );
not \U$14590 ( \14967 , \14965 );
and \U$14591 ( \14968 , \14967 , \14462 );
nor \U$14592 ( \14969 , \14966 , \14968 );
xor \U$14593 ( \14970 , \14957 , \14969 );
and \U$14594 ( \14971 , \14059 , RIae78a58_123);
and \U$14595 ( \14972 , RIae78cb0_128, \14057 );
nor \U$14596 ( \14973 , \14971 , \14972 );
and \U$14597 ( \14974 , \14973 , \13502 );
not \U$14598 ( \14975 , \14973 );
and \U$14599 ( \14976 , \14975 , \14063 );
nor \U$14600 ( \14977 , \14974 , \14976 );
and \U$14601 ( \14978 , \14970 , \14977 );
and \U$14602 ( \14979 , \14957 , \14969 );
or \U$14603 ( \14980 , \14978 , \14979 );
xor \U$14604 ( \14981 , \14950 , \14980 );
and \U$14605 ( \14982 , \10548 , RIae76028_33);
and \U$14606 ( \14983 , RIae762f8_39, \10546 );
nor \U$14607 ( \14984 , \14982 , \14983 );
and \U$14608 ( \14985 , \14984 , \10421 );
not \U$14609 ( \14986 , \14984 );
and \U$14610 ( \14987 , \14986 , \10118 );
nor \U$14611 ( \14988 , \14985 , \14987 );
and \U$14612 ( \14989 , \11470 , RIae76208_37);
and \U$14613 ( \14990 , RIae76a78_55, \11468 );
nor \U$14614 ( \14991 , \14989 , \14990 );
and \U$14615 ( \14992 , \14991 , \10936 );
not \U$14616 ( \14993 , \14991 );
and \U$14617 ( \14994 , \14993 , \11474 );
nor \U$14618 ( \14995 , \14992 , \14994 );
xor \U$14619 ( \14996 , \14988 , \14995 );
and \U$14620 ( \14997 , \12180 , RIae76988_53);
and \U$14621 ( \14998 , RIae767a8_49, \12178 );
nor \U$14622 ( \14999 , \14997 , \14998 );
and \U$14623 ( \15000 , \14999 , \12184 );
not \U$14624 ( \15001 , \14999 );
and \U$14625 ( \15002 , \15001 , \11827 );
nor \U$14626 ( \15003 , \15000 , \15002 );
and \U$14627 ( \15004 , \14996 , \15003 );
and \U$14628 ( \15005 , \14988 , \14995 );
or \U$14629 ( \15006 , \15004 , \15005 );
and \U$14630 ( \15007 , \14981 , \15006 );
and \U$14631 ( \15008 , \14950 , \14980 );
or \U$14632 ( \15009 , \15007 , \15008 );
xor \U$14633 ( \15010 , \14925 , \15009 );
and \U$14634 ( \15011 , \6172 , RIae754e8_9);
and \U$14635 ( \15012 , RIae757b8_15, \6170 );
nor \U$14636 ( \15013 , \15011 , \15012 );
and \U$14637 ( \15014 , \15013 , \6176 );
not \U$14638 ( \15015 , \15013 );
and \U$14639 ( \15016 , \15015 , \6175 );
nor \U$14640 ( \15017 , \15014 , \15016 );
and \U$14641 ( \15018 , \6941 , RIae756c8_13);
and \U$14642 ( \15019 , RIae75218_3, \6939 );
nor \U$14643 ( \15020 , \15018 , \15019 );
and \U$14644 ( \15021 , \15020 , \6314 );
not \U$14645 ( \15022 , \15020 );
and \U$14646 ( \15023 , \15022 , \6945 );
nor \U$14647 ( \15024 , \15021 , \15023 );
xor \U$14648 ( \15025 , \15017 , \15024 );
and \U$14649 ( \15026 , \7633 , RIae75128_1);
and \U$14650 ( \15027 , RIae75308_5, \7631 );
nor \U$14651 ( \15028 , \15026 , \15027 );
and \U$14652 ( \15029 , \15028 , \7206 );
not \U$14653 ( \15030 , \15028 );
and \U$14654 ( \15031 , \15030 , \7205 );
nor \U$14655 ( \15032 , \15029 , \15031 );
and \U$14656 ( \15033 , \15025 , \15032 );
and \U$14657 ( \15034 , \15017 , \15024 );
or \U$14658 ( \15035 , \15033 , \15034 );
and \U$14659 ( \15036 , \5399 , RIae75e48_29);
and \U$14660 ( \15037 , RIae75c68_25, \5397 );
nor \U$14661 ( \15038 , \15036 , \15037 );
and \U$14662 ( \15039 , \15038 , \5016 );
not \U$14663 ( \15040 , \15038 );
and \U$14664 ( \15041 , \15040 , \5403 );
nor \U$14665 ( \15042 , \15039 , \15041 );
and \U$14666 ( \15043 , \4688 , RIae758a8_17);
and \U$14667 ( \15044 , RIae75f38_31, \4686 );
nor \U$14668 ( \15045 , \15043 , \15044 );
and \U$14669 ( \15046 , \15045 , \4481 );
not \U$14670 ( \15047 , \15045 );
and \U$14671 ( \15048 , \15047 , \4482 );
nor \U$14672 ( \15049 , \15046 , \15048 );
xor \U$14673 ( \15050 , \15042 , \15049 );
and \U$14674 ( \15051 , \5896 , RIae75d58_27);
and \U$14675 ( \15052 , RIae755d8_11, \5894 );
nor \U$14676 ( \15053 , \15051 , \15052 );
and \U$14677 ( \15054 , \15053 , \5590 );
not \U$14678 ( \15055 , \15053 );
and \U$14679 ( \15056 , \15055 , \5589 );
nor \U$14680 ( \15057 , \15054 , \15056 );
and \U$14681 ( \15058 , \15050 , \15057 );
and \U$14682 ( \15059 , \15042 , \15049 );
or \U$14683 ( \15060 , \15058 , \15059 );
xor \U$14684 ( \15061 , \15035 , \15060 );
and \U$14685 ( \15062 , \4247 , RIae75a88_21);
and \U$14686 ( \15063 , RIae75998_19, \4245 );
nor \U$14687 ( \15064 , \15062 , \15063 );
and \U$14688 ( \15065 , \15064 , \3989 );
not \U$14689 ( \15066 , \15064 );
and \U$14690 ( \15067 , \15066 , \4251 );
nor \U$14691 ( \15068 , \15065 , \15067 );
not \U$14692 ( \15069 , \3218 );
and \U$14693 ( \15070 , \3214 , RIae78878_119);
and \U$14694 ( \15071 , RIae78788_117, \3212 );
nor \U$14695 ( \15072 , \15070 , \15071 );
not \U$14696 ( \15073 , \15072 );
or \U$14697 ( \15074 , \15069 , \15073 );
or \U$14698 ( \15075 , \15072 , \3218 );
nand \U$14699 ( \15076 , \15074 , \15075 );
xor \U$14700 ( \15077 , \15068 , \15076 );
and \U$14701 ( \15078 , \3730 , RIae78698_115);
and \U$14702 ( \15079 , RIae75b78_23, \3728 );
nor \U$14703 ( \15080 , \15078 , \15079 );
and \U$14704 ( \15081 , \15080 , \3732 );
not \U$14705 ( \15082 , \15080 );
and \U$14706 ( \15083 , \15082 , \3422 );
nor \U$14707 ( \15084 , \15081 , \15083 );
and \U$14708 ( \15085 , \15077 , \15084 );
and \U$14709 ( \15086 , \15068 , \15076 );
or \U$14710 ( \15087 , \15085 , \15086 );
and \U$14711 ( \15088 , \15061 , \15087 );
and \U$14712 ( \15089 , \15035 , \15060 );
or \U$14713 ( \15090 , \15088 , \15089 );
and \U$14714 ( \15091 , \15010 , \15090 );
and \U$14715 ( \15092 , \14925 , \15009 );
or \U$14716 ( \15093 , \15091 , \15092 );
xor \U$14717 ( \15094 , \14844 , \15093 );
xor \U$14718 ( \15095 , \14511 , \14518 );
xor \U$14719 ( \15096 , \15095 , \14526 );
xor \U$14720 ( \15097 , \14563 , \14570 );
xor \U$14721 ( \15098 , \15097 , \14578 );
and \U$14722 ( \15099 , \15096 , \15098 );
xor \U$14723 ( \15100 , \14482 , \14489 );
xor \U$14724 ( \15101 , \15100 , \14497 );
xor \U$14725 ( \15102 , \14563 , \14570 );
xor \U$14726 ( \15103 , \15102 , \14578 );
and \U$14727 ( \15104 , \15101 , \15103 );
and \U$14728 ( \15105 , \15096 , \15101 );
or \U$14729 ( \15106 , \15099 , \15104 , \15105 );
xor \U$14730 ( \15107 , \14435 , \14442 );
xor \U$14731 ( \15108 , \15107 , \14450 );
xor \U$14732 ( \15109 , \14460 , \14463 );
xor \U$14733 ( \15110 , \15109 , \14471 );
and \U$14734 ( \15111 , \15108 , \15110 );
xor \U$14735 ( \15112 , \15106 , \15111 );
xor \U$14736 ( \15113 , \14026 , \14033 );
xor \U$14737 ( \15114 , \15113 , \14041 );
xor \U$14738 ( \15115 , \14327 , \14332 );
xor \U$14739 ( \15116 , \15114 , \15115 );
and \U$14740 ( \15117 , \15112 , \15116 );
and \U$14741 ( \15118 , \15106 , \15111 );
or \U$14742 ( \15119 , \15117 , \15118 );
and \U$14743 ( \15120 , \15094 , \15119 );
and \U$14744 ( \15121 , \14844 , \15093 );
or \U$14745 ( \15122 , \15120 , \15121 );
xor \U$14746 ( \15123 , \14769 , \15122 );
xor \U$14747 ( \15124 , \14337 , \14339 );
xor \U$14748 ( \15125 , \15124 , \14344 );
xor \U$14749 ( \15126 , \14600 , \14633 );
xor \U$14750 ( \15127 , \15126 , \14646 );
and \U$14751 ( \15128 , \15125 , \15127 );
xor \U$14752 ( \15129 , \13894 , \13900 );
xor \U$14753 ( \15130 , \15129 , \13907 );
xor \U$14754 ( \15131 , \14312 , \14317 );
xor \U$14755 ( \15132 , \15130 , \15131 );
xor \U$14756 ( \15133 , \14600 , \14633 );
xor \U$14757 ( \15134 , \15133 , \14646 );
and \U$14758 ( \15135 , \15132 , \15134 );
and \U$14759 ( \15136 , \15125 , \15132 );
or \U$14760 ( \15137 , \15128 , \15135 , \15136 );
and \U$14761 ( \15138 , \15123 , \15137 );
and \U$14762 ( \15139 , \14769 , \15122 );
or \U$14763 ( \15140 , \15138 , \15139 );
xor \U$14764 ( \15141 , \13851 , \13887 );
xor \U$14765 ( \15142 , \15141 , \13910 );
xor \U$14766 ( \15143 , \13994 , \14079 );
xor \U$14767 ( \15144 , \15143 , \14160 );
xor \U$14768 ( \15145 , \15142 , \15144 );
xor \U$14769 ( \15146 , \14657 , \14659 );
xor \U$14770 ( \15147 , \15146 , \14662 );
and \U$14771 ( \15148 , \15145 , \15147 );
and \U$14772 ( \15149 , \15142 , \15144 );
or \U$14773 ( \15150 , \15148 , \15149 );
xor \U$14774 ( \15151 , \15140 , \15150 );
not \U$14775 ( \15152 , \14683 );
xor \U$14776 ( \15153 , \14686 , \14693 );
not \U$14777 ( \15154 , \15153 );
or \U$14778 ( \15155 , \15152 , \15154 );
or \U$14779 ( \15156 , \15153 , \14683 );
nand \U$14780 ( \15157 , \15155 , \15156 );
and \U$14781 ( \15158 , \15151 , \15157 );
and \U$14782 ( \15159 , \15140 , \15150 );
or \U$14783 ( \15160 , \15158 , \15159 );
nand \U$14784 ( \15161 , \14733 , \15160 );
nand \U$14785 ( \15162 , \14730 , \15161 );
nand \U$14786 ( \15163 , \14723 , \15162 );
nand \U$14787 ( \15164 , \14720 , \15163 );
not \U$14788 ( \15165 , \14701 );
not \U$14789 ( \15166 , \14712 );
or \U$14790 ( \15167 , \15165 , \15166 );
or \U$14791 ( \15168 , \14712 , \14701 );
nand \U$14792 ( \15169 , \15167 , \15168 );
and \U$14793 ( \15170 , \15164 , \15169 );
xor \U$14794 ( \15171 , \15169 , \15164 );
xor \U$14795 ( \15172 , \14781 , \14830 );
xor \U$14796 ( \15173 , \15172 , \14841 );
xor \U$14797 ( \15174 , \15106 , \15111 );
xor \U$14798 ( \15175 , \15174 , \15116 );
and \U$14799 ( \15176 , \15173 , \15175 );
xor \U$14800 ( \15177 , \14627 , \13852 );
xor \U$14801 ( \15178 , \15177 , \14630 );
xor \U$14802 ( \15179 , \14737 , \14744 );
xor \U$14803 ( \15180 , \15178 , \15179 );
xor \U$14804 ( \15181 , \15106 , \15111 );
xor \U$14805 ( \15182 , \15181 , \15116 );
and \U$14806 ( \15183 , \15180 , \15182 );
and \U$14807 ( \15184 , \15173 , \15180 );
or \U$14808 ( \15185 , \15176 , \15183 , \15184 );
xor \U$14809 ( \15186 , \14876 , \14883 );
xor \U$14810 ( \15187 , \15186 , \14892 );
xor \U$14811 ( \15188 , \14808 , \14816 );
xor \U$14812 ( \15189 , \15188 , \14824 );
and \U$14813 ( \15190 , \15187 , \15189 );
xor \U$14814 ( \15191 , \14851 , \14858 );
xor \U$14815 ( \15192 , \15191 , \14866 );
xor \U$14816 ( \15193 , \14808 , \14816 );
xor \U$14817 ( \15194 , \15193 , \14824 );
and \U$14818 ( \15195 , \15192 , \15194 );
and \U$14819 ( \15196 , \15187 , \15192 );
or \U$14820 ( \15197 , \15190 , \15195 , \15196 );
not \U$14821 ( \15198 , \400 );
and \U$14822 ( \15199 , \436 , RIae77a68_89);
and \U$14823 ( \15200 , RIae77978_87, \434 );
nor \U$14824 ( \15201 , \15199 , \15200 );
not \U$14825 ( \15202 , \15201 );
or \U$14826 ( \15203 , \15198 , \15202 );
or \U$14827 ( \15204 , \15201 , \400 );
nand \U$14828 ( \15205 , \15203 , \15204 );
not \U$14829 ( \15206 , RIae774c8_77);
nor \U$14830 ( \15207 , \15206 , \491 );
xor \U$14831 ( \15208 , \15205 , \15207 );
not \U$14832 ( \15209 , \392 );
and \U$14833 ( \15210 , \384 , RIae77720_82);
and \U$14834 ( \15211 , RIae773d8_75, \382 );
nor \U$14835 ( \15212 , \15210 , \15211 );
not \U$14836 ( \15213 , \15212 );
or \U$14837 ( \15214 , \15209 , \15213 );
or \U$14838 ( \15215 , \15212 , \392 );
nand \U$14839 ( \15216 , \15214 , \15215 );
and \U$14840 ( \15217 , \15208 , \15216 );
and \U$14841 ( \15218 , \15205 , \15207 );
or \U$14842 ( \15219 , \15217 , \15218 );
or \U$14843 ( \15220 , \14790 , \14782 );
nand \U$14844 ( \15221 , \15220 , \14791 );
xor \U$14845 ( \15222 , \15219 , \15221 );
and \U$14846 ( \15223 , \558 , RIae76f28_65);
and \U$14847 ( \15224 , RIae76e38_63, \556 );
nor \U$14848 ( \15225 , \15223 , \15224 );
and \U$14849 ( \15226 , \15225 , \562 );
not \U$14850 ( \15227 , \15225 );
and \U$14851 ( \15228 , \15227 , \504 );
nor \U$14852 ( \15229 , \15226 , \15228 );
and \U$14853 ( \15230 , \672 , RIae76d48_61);
and \U$14854 ( \15231 , RIae76c58_59, \670 );
nor \U$14855 ( \15232 , \15230 , \15231 );
and \U$14856 ( \15233 , \15232 , \587 );
not \U$14857 ( \15234 , \15232 );
and \U$14858 ( \15235 , \15234 , \588 );
nor \U$14859 ( \15236 , \15233 , \15235 );
xor \U$14860 ( \15237 , \15229 , \15236 );
and \U$14861 ( \15238 , \514 , RIae77798_83);
and \U$14862 ( \15239 , RIae77888_85, \512 );
nor \U$14863 ( \15240 , \15238 , \15239 );
not \U$14864 ( \15241 , \15240 );
not \U$14865 ( \15242 , \471 );
and \U$14866 ( \15243 , \15241 , \15242 );
and \U$14867 ( \15244 , \15240 , \469 );
nor \U$14868 ( \15245 , \15243 , \15244 );
and \U$14869 ( \15246 , \15237 , \15245 );
and \U$14870 ( \15247 , \15229 , \15236 );
nor \U$14871 ( \15248 , \15246 , \15247 );
and \U$14872 ( \15249 , \15222 , \15248 );
and \U$14873 ( \15250 , \15219 , \15221 );
or \U$14874 ( \15251 , \15249 , \15250 );
xor \U$14875 ( \15252 , \15197 , \15251 );
xor \U$14876 ( \15253 , \15042 , \15049 );
xor \U$14877 ( \15254 , \15253 , \15057 );
xor \U$14878 ( \15255 , \14903 , \14910 );
xor \U$14879 ( \15256 , \15255 , \14919 );
xor \U$14880 ( \15257 , \15254 , \15256 );
xor \U$14881 ( \15258 , \15068 , \15076 );
xor \U$14882 ( \15259 , \15258 , \15084 );
and \U$14883 ( \15260 , \15257 , \15259 );
and \U$14884 ( \15261 , \15254 , \15256 );
or \U$14885 ( \15262 , \15260 , \15261 );
and \U$14886 ( \15263 , \15252 , \15262 );
and \U$14887 ( \15264 , \15197 , \15251 );
or \U$14888 ( \15265 , \15263 , \15264 );
and \U$14889 ( \15266 , \6941 , RIae757b8_15);
and \U$14890 ( \15267 , RIae756c8_13, \6939 );
nor \U$14891 ( \15268 , \15266 , \15267 );
and \U$14892 ( \15269 , \15268 , \6945 );
not \U$14893 ( \15270 , \15268 );
and \U$14894 ( \15271 , \15270 , \6314 );
nor \U$14895 ( \15272 , \15269 , \15271 );
and \U$14896 ( \15273 , \7633 , RIae75218_3);
and \U$14897 ( \15274 , RIae75128_1, \7631 );
nor \U$14898 ( \15275 , \15273 , \15274 );
and \U$14899 ( \15276 , \15275 , \7205 );
not \U$14900 ( \15277 , \15275 );
and \U$14901 ( \15278 , \15277 , \7206 );
nor \U$14902 ( \15279 , \15276 , \15278 );
or \U$14903 ( \15280 , \15272 , \15279 );
not \U$14904 ( \15281 , \15279 );
not \U$14905 ( \15282 , \15272 );
or \U$14906 ( \15283 , \15281 , \15282 );
and \U$14907 ( \15284 , \8371 , RIae75308_5);
and \U$14908 ( \15285 , RIae753f8_7, \8369 );
nor \U$14909 ( \15286 , \15284 , \15285 );
and \U$14910 ( \15287 , \15286 , \8020 );
not \U$14911 ( \15288 , \15286 );
and \U$14912 ( \15289 , \15288 , \8019 );
nor \U$14913 ( \15290 , \15287 , \15289 );
nand \U$14914 ( \15291 , \15283 , \15290 );
nand \U$14915 ( \15292 , \15280 , \15291 );
and \U$14916 ( \15293 , \4688 , RIae75998_19);
and \U$14917 ( \15294 , RIae758a8_17, \4686 );
nor \U$14918 ( \15295 , \15293 , \15294 );
and \U$14919 ( \15296 , \15295 , \4481 );
not \U$14920 ( \15297 , \15295 );
and \U$14921 ( \15298 , \15297 , \4482 );
nor \U$14922 ( \15299 , \15296 , \15298 );
and \U$14923 ( \15300 , \3730 , RIae78788_117);
and \U$14924 ( \15301 , RIae78698_115, \3728 );
nor \U$14925 ( \15302 , \15300 , \15301 );
and \U$14926 ( \15303 , \15302 , \3732 );
not \U$14927 ( \15304 , \15302 );
and \U$14928 ( \15305 , \15304 , \3422 );
nor \U$14929 ( \15306 , \15303 , \15305 );
xor \U$14930 ( \15307 , \15299 , \15306 );
and \U$14931 ( \15308 , \4247 , RIae75b78_23);
and \U$14932 ( \15309 , RIae75a88_21, \4245 );
nor \U$14933 ( \15310 , \15308 , \15309 );
and \U$14934 ( \15311 , \15310 , \3989 );
not \U$14935 ( \15312 , \15310 );
and \U$14936 ( \15313 , \15312 , \4251 );
nor \U$14937 ( \15314 , \15311 , \15313 );
and \U$14938 ( \15315 , \15307 , \15314 );
and \U$14939 ( \15316 , \15299 , \15306 );
or \U$14940 ( \15317 , \15315 , \15316 );
xor \U$14941 ( \15318 , \15292 , \15317 );
and \U$14942 ( \15319 , \5896 , RIae75c68_25);
and \U$14943 ( \15320 , RIae75d58_27, \5894 );
nor \U$14944 ( \15321 , \15319 , \15320 );
and \U$14945 ( \15322 , \15321 , \5590 );
not \U$14946 ( \15323 , \15321 );
and \U$14947 ( \15324 , \15323 , \5589 );
nor \U$14948 ( \15325 , \15322 , \15324 );
and \U$14949 ( \15326 , \5399 , RIae75f38_31);
and \U$14950 ( \15327 , RIae75e48_29, \5397 );
nor \U$14951 ( \15328 , \15326 , \15327 );
and \U$14952 ( \15329 , \15328 , \5016 );
not \U$14953 ( \15330 , \15328 );
and \U$14954 ( \15331 , \15330 , \5403 );
nor \U$14955 ( \15332 , \15329 , \15331 );
xor \U$14956 ( \15333 , \15325 , \15332 );
and \U$14957 ( \15334 , \6172 , RIae755d8_11);
and \U$14958 ( \15335 , RIae754e8_9, \6170 );
nor \U$14959 ( \15336 , \15334 , \15335 );
and \U$14960 ( \15337 , \15336 , \6176 );
not \U$14961 ( \15338 , \15336 );
and \U$14962 ( \15339 , \15338 , \6175 );
nor \U$14963 ( \15340 , \15337 , \15339 );
and \U$14964 ( \15341 , \15333 , \15340 );
and \U$14965 ( \15342 , \15325 , \15332 );
or \U$14966 ( \15343 , \15341 , \15342 );
and \U$14967 ( \15344 , \15318 , \15343 );
and \U$14968 ( \15345 , \15292 , \15317 );
or \U$14969 ( \15346 , \15344 , \15345 );
not \U$14970 ( \15347 , \3218 );
and \U$14971 ( \15348 , \3214 , RIae78968_121);
and \U$14972 ( \15349 , RIae78878_119, \3212 );
nor \U$14973 ( \15350 , \15348 , \15349 );
not \U$14974 ( \15351 , \15350 );
or \U$14975 ( \15352 , \15347 , \15351 );
or \U$14976 ( \15353 , \15350 , \2774 );
nand \U$14977 ( \15354 , \15352 , \15353 );
and \U$14978 ( \15355 , \2607 , RIae77c48_93);
and \U$14979 ( \15356 , RIae77b58_91, \2605 );
nor \U$14980 ( \15357 , \15355 , \15356 );
and \U$14981 ( \15358 , \15357 , \2611 );
not \U$14982 ( \15359 , \15357 );
and \U$14983 ( \15360 , \15359 , \2397 );
nor \U$14984 ( \15361 , \15358 , \15360 );
xor \U$14985 ( \15362 , \15354 , \15361 );
not \U$14986 ( \15363 , \2789 );
and \U$14987 ( \15364 , \2783 , RIae77d38_95);
and \U$14988 ( \15365 , RIae77e28_97, \2781 );
nor \U$14989 ( \15366 , \15364 , \15365 );
not \U$14990 ( \15367 , \15366 );
or \U$14991 ( \15368 , \15363 , \15367 );
or \U$14992 ( \15369 , \15366 , \2789 );
nand \U$14993 ( \15370 , \15368 , \15369 );
and \U$14994 ( \15371 , \15362 , \15370 );
and \U$14995 ( \15372 , \15354 , \15361 );
or \U$14996 ( \15373 , \15371 , \15372 );
and \U$14997 ( \15374 , \2224 , RIae783c8_109);
and \U$14998 ( \15375 , RIae78530_112, \2222 );
nor \U$14999 ( \15376 , \15374 , \15375 );
and \U$15000 ( \15377 , \15376 , \2061 );
not \U$15001 ( \15378 , \15376 );
and \U$15002 ( \15379 , \15378 , \2060 );
nor \U$15003 ( \15380 , \15377 , \15379 );
and \U$15004 ( \15381 , \1593 , RIae77f18_99);
and \U$15005 ( \15382 , RIae78008_101, \1591 );
nor \U$15006 ( \15383 , \15381 , \15382 );
and \U$15007 ( \15384 , \15383 , \1498 );
not \U$15008 ( \15385 , \15383 );
and \U$15009 ( \15386 , \15385 , \1488 );
nor \U$15010 ( \15387 , \15384 , \15386 );
xor \U$15011 ( \15388 , \15380 , \15387 );
and \U$15012 ( \15389 , \1939 , RIae781e8_105);
and \U$15013 ( \15390 , RIae785a8_113, \1937 );
nor \U$15014 ( \15391 , \15389 , \15390 );
and \U$15015 ( \15392 , \15391 , \1735 );
not \U$15016 ( \15393 , \15391 );
and \U$15017 ( \15394 , \15393 , \1734 );
nor \U$15018 ( \15395 , \15392 , \15394 );
and \U$15019 ( \15396 , \15388 , \15395 );
and \U$15020 ( \15397 , \15380 , \15387 );
or \U$15021 ( \15398 , \15396 , \15397 );
xor \U$15022 ( \15399 , \15373 , \15398 );
and \U$15023 ( \15400 , \883 , RIae77180_70);
and \U$15024 ( \15401 , RIae77018_67, \881 );
nor \U$15025 ( \15402 , \15400 , \15401 );
not \U$15026 ( \15403 , \15402 );
not \U$15027 ( \15404 , \787 );
and \U$15028 ( \15405 , \15403 , \15404 );
and \U$15029 ( \15406 , \15402 , \789 );
nor \U$15030 ( \15407 , \15405 , \15406 );
and \U$15031 ( \15408 , \1138 , RIae771f8_71);
and \U$15032 ( \15409 , RIae772e8_73, \1136 );
nor \U$15033 ( \15410 , \15408 , \15409 );
and \U$15034 ( \15411 , \15410 , \1142 );
not \U$15035 ( \15412 , \15410 );
and \U$15036 ( \15413 , \15412 , \1012 );
nor \U$15037 ( \15414 , \15411 , \15413 );
or \U$15038 ( \15415 , \15407 , \15414 );
not \U$15039 ( \15416 , \15414 );
not \U$15040 ( \15417 , \15407 );
or \U$15041 ( \15418 , \15416 , \15417 );
and \U$15042 ( \15419 , \1376 , RIae782d8_107);
and \U$15043 ( \15420 , RIae780f8_103, \1374 );
nor \U$15044 ( \15421 , \15419 , \15420 );
and \U$15045 ( \15422 , \15421 , \1380 );
not \U$15046 ( \15423 , \15421 );
and \U$15047 ( \15424 , \15423 , \1261 );
nor \U$15048 ( \15425 , \15422 , \15424 );
nand \U$15049 ( \15426 , \15418 , \15425 );
nand \U$15050 ( \15427 , \15415 , \15426 );
and \U$15051 ( \15428 , \15399 , \15427 );
and \U$15052 ( \15429 , \15373 , \15398 );
or \U$15053 ( \15430 , \15428 , \15429 );
xor \U$15054 ( \15431 , \15346 , \15430 );
and \U$15055 ( \15432 , \8966 , RIae763e8_41);
and \U$15056 ( \15433 , RIae764d8_43, \8964 );
nor \U$15057 ( \15434 , \15432 , \15433 );
and \U$15058 ( \15435 , \15434 , \8789 );
not \U$15059 ( \15436 , \15434 );
and \U$15060 ( \15437 , \15436 , \8799 );
nor \U$15061 ( \15438 , \15435 , \15437 );
and \U$15062 ( \15439 , \9760 , RIae766b8_47);
and \U$15063 ( \15440 , RIae765c8_45, \9758 );
nor \U$15064 ( \15441 , \15439 , \15440 );
and \U$15065 ( \15442 , \15441 , \9272 );
not \U$15066 ( \15443 , \15441 );
and \U$15067 ( \15444 , \15443 , \9273 );
nor \U$15068 ( \15445 , \15442 , \15444 );
xor \U$15069 ( \15446 , \15438 , \15445 );
and \U$15070 ( \15447 , \10548 , RIae76118_35);
and \U$15071 ( \15448 , RIae76028_33, \10546 );
nor \U$15072 ( \15449 , \15447 , \15448 );
and \U$15073 ( \15450 , \15449 , \10118 );
not \U$15074 ( \15451 , \15449 );
and \U$15075 ( \15452 , \15451 , \10421 );
nor \U$15076 ( \15453 , \15450 , \15452 );
and \U$15077 ( \15454 , \15446 , \15453 );
and \U$15078 ( \15455 , \15438 , \15445 );
or \U$15079 ( \15456 , \15454 , \15455 );
and \U$15080 ( \15457 , \11470 , RIae762f8_39);
and \U$15081 ( \15458 , RIae76208_37, \11468 );
nor \U$15082 ( \15459 , \15457 , \15458 );
and \U$15083 ( \15460 , \15459 , \11474 );
not \U$15084 ( \15461 , \15459 );
and \U$15085 ( \15462 , \15461 , \10936 );
nor \U$15086 ( \15463 , \15460 , \15462 );
not \U$15087 ( \15464 , \15463 );
and \U$15088 ( \15465 , \13059 , RIae767a8_49);
and \U$15089 ( \15466 , RIae76898_51, \13057 );
nor \U$15090 ( \15467 , \15465 , \15466 );
and \U$15091 ( \15468 , \15467 , \12718 );
not \U$15092 ( \15469 , \15467 );
and \U$15093 ( \15470 , \15469 , \13063 );
nor \U$15094 ( \15471 , \15468 , \15470 );
not \U$15095 ( \15472 , \15471 );
and \U$15096 ( \15473 , \15464 , \15472 );
and \U$15097 ( \15474 , \15471 , \15463 );
and \U$15098 ( \15475 , \12180 , RIae76a78_55);
and \U$15099 ( \15476 , RIae76988_53, \12178 );
nor \U$15100 ( \15477 , \15475 , \15476 );
and \U$15101 ( \15478 , \15477 , \11827 );
not \U$15102 ( \15479 , \15477 );
and \U$15103 ( \15480 , \15479 , \12184 );
nor \U$15104 ( \15481 , \15478 , \15480 );
nor \U$15105 ( \15482 , \15474 , \15481 );
nor \U$15106 ( \15483 , \15473 , \15482 );
or \U$15107 ( \15484 , \15456 , \15483 );
not \U$15108 ( \15485 , \15456 );
not \U$15109 ( \15486 , \15483 );
or \U$15110 ( \15487 , \15485 , \15486 );
and \U$15111 ( \15488 , \14964 , RIae78cb0_128);
and \U$15112 ( \15489 , RIae78da0_130, \14962 );
nor \U$15113 ( \15490 , \15488 , \15489 );
and \U$15114 ( \15491 , \15490 , \14462 );
not \U$15115 ( \15492 , \15490 );
and \U$15116 ( \15493 , \15492 , \14463 );
nor \U$15117 ( \15494 , \15491 , \15493 );
or \U$15118 ( \15495 , \15494 , RIae7aa38_191);
and \U$15119 ( \15496 , \15494 , RIae7aa38_191);
and \U$15120 ( \15497 , \14059 , RIae76b68_57);
and \U$15121 ( \15498 , RIae78a58_123, \14057 );
nor \U$15122 ( \15499 , \15497 , \15498 );
and \U$15123 ( \15500 , \15499 , \14063 );
not \U$15124 ( \15501 , \15499 );
and \U$15125 ( \15502 , \15501 , \13502 );
nor \U$15126 ( \15503 , \15500 , \15502 );
nor \U$15127 ( \15504 , \15496 , \15503 );
not \U$15128 ( \15505 , \15504 );
nand \U$15129 ( \15506 , \15495 , \15505 );
nand \U$15130 ( \15507 , \15487 , \15506 );
nand \U$15131 ( \15508 , \15484 , \15507 );
and \U$15132 ( \15509 , \15431 , \15508 );
and \U$15133 ( \15510 , \15346 , \15430 );
or \U$15134 ( \15511 , \15509 , \15510 );
xor \U$15135 ( \15512 , \15265 , \15511 );
xor \U$15136 ( \15513 , \15017 , \15024 );
xor \U$15137 ( \15514 , \15513 , \15032 );
xor \U$15138 ( \15515 , \14932 , \14939 );
xor \U$15139 ( \15516 , \15515 , \14947 );
and \U$15140 ( \15517 , \15514 , \15516 );
xor \U$15141 ( \15518 , \14988 , \14995 );
xor \U$15142 ( \15519 , \15518 , \15003 );
xor \U$15143 ( \15520 , \14932 , \14939 );
xor \U$15144 ( \15521 , \15520 , \14947 );
and \U$15145 ( \15522 , \15519 , \15521 );
and \U$15146 ( \15523 , \15514 , \15519 );
or \U$15147 ( \15524 , \15517 , \15522 , \15523 );
xor \U$15148 ( \15525 , \15108 , \15110 );
xor \U$15149 ( \15526 , \15524 , \15525 );
xor \U$15150 ( \15527 , \14563 , \14570 );
xor \U$15151 ( \15528 , \15527 , \14578 );
xor \U$15152 ( \15529 , \15096 , \15101 );
xor \U$15153 ( \15530 , \15528 , \15529 );
and \U$15154 ( \15531 , \15526 , \15530 );
and \U$15155 ( \15532 , \15524 , \15525 );
or \U$15156 ( \15533 , \15531 , \15532 );
and \U$15157 ( \15534 , \15512 , \15533 );
and \U$15158 ( \15535 , \15265 , \15511 );
or \U$15159 ( \15536 , \15534 , \15535 );
xor \U$15160 ( \15537 , \15185 , \15536 );
xor \U$15161 ( \15538 , \14791 , \14799 );
xor \U$15162 ( \15539 , \15538 , \14827 );
xor \U$15163 ( \15540 , \14833 , \14835 );
xor \U$15164 ( \15541 , \15540 , \14838 );
and \U$15165 ( \15542 , \15539 , \15541 );
xor \U$15166 ( \15543 , \14608 , \14616 );
xor \U$15167 ( \15544 , \15543 , \14624 );
xor \U$15168 ( \15545 , \14771 , \14776 );
xor \U$15169 ( \15546 , \15544 , \15545 );
xor \U$15170 ( \15547 , \14833 , \14835 );
xor \U$15171 ( \15548 , \15547 , \14838 );
and \U$15172 ( \15549 , \15546 , \15548 );
and \U$15173 ( \15550 , \15539 , \15546 );
or \U$15174 ( \15551 , \15542 , \15549 , \15550 );
xor \U$15175 ( \15552 , \14950 , \14980 );
xor \U$15176 ( \15553 , \15552 , \15006 );
xor \U$15177 ( \15554 , \14869 , \14895 );
xor \U$15178 ( \15555 , \15554 , \14922 );
and \U$15179 ( \15556 , \15553 , \15555 );
xor \U$15180 ( \15557 , \15035 , \15060 );
xor \U$15181 ( \15558 , \15557 , \15087 );
xor \U$15182 ( \15559 , \14869 , \14895 );
xor \U$15183 ( \15560 , \15559 , \14922 );
and \U$15184 ( \15561 , \15558 , \15560 );
and \U$15185 ( \15562 , \15553 , \15558 );
or \U$15186 ( \15563 , \15556 , \15561 , \15562 );
xor \U$15187 ( \15564 , \15551 , \15563 );
xor \U$15188 ( \15565 , \14529 , \14555 );
xor \U$15189 ( \15566 , \15565 , \14581 );
xor \U$15190 ( \15567 , \14751 , \14756 );
xor \U$15191 ( \15568 , \15566 , \15567 );
and \U$15192 ( \15569 , \15564 , \15568 );
and \U$15193 ( \15570 , \15551 , \15563 );
or \U$15194 ( \15571 , \15569 , \15570 );
xor \U$15195 ( \15572 , \15537 , \15571 );
xor \U$15196 ( \15573 , \14808 , \14816 );
xor \U$15197 ( \15574 , \15573 , \14824 );
xor \U$15198 ( \15575 , \15187 , \15192 );
xor \U$15199 ( \15576 , \15574 , \15575 );
xor \U$15200 ( \15577 , \15254 , \15256 );
xor \U$15201 ( \15578 , \15577 , \15259 );
and \U$15202 ( \15579 , \15576 , \15578 );
xor \U$15203 ( \15580 , \14932 , \14939 );
xor \U$15204 ( \15581 , \15580 , \14947 );
xor \U$15205 ( \15582 , \15514 , \15519 );
xor \U$15206 ( \15583 , \15581 , \15582 );
xor \U$15207 ( \15584 , \15254 , \15256 );
xor \U$15208 ( \15585 , \15584 , \15259 );
and \U$15209 ( \15586 , \15583 , \15585 );
and \U$15210 ( \15587 , \15576 , \15583 );
or \U$15211 ( \15588 , \15579 , \15586 , \15587 );
xor \U$15212 ( \15589 , \15219 , \15221 );
xor \U$15213 ( \15590 , \15589 , \15248 );
xor \U$15214 ( \15591 , \15373 , \15398 );
xor \U$15215 ( \15592 , \15591 , \15427 );
xor \U$15216 ( \15593 , \15590 , \15592 );
xor \U$15217 ( \15594 , \15292 , \15317 );
xor \U$15218 ( \15595 , \15594 , \15343 );
and \U$15219 ( \15596 , \15593 , \15595 );
and \U$15220 ( \15597 , \15590 , \15592 );
or \U$15221 ( \15598 , \15596 , \15597 );
xor \U$15222 ( \15599 , \15588 , \15598 );
xor \U$15223 ( \15600 , \14869 , \14895 );
xor \U$15224 ( \15601 , \15600 , \14922 );
xor \U$15225 ( \15602 , \15553 , \15558 );
xor \U$15226 ( \15603 , \15601 , \15602 );
and \U$15227 ( \15604 , \15599 , \15603 );
and \U$15228 ( \15605 , \15588 , \15598 );
or \U$15229 ( \15606 , \15604 , \15605 );
and \U$15230 ( \15607 , \2224 , RIae785a8_113);
and \U$15231 ( \15608 , RIae783c8_109, \2222 );
nor \U$15232 ( \15609 , \15607 , \15608 );
and \U$15233 ( \15610 , \15609 , \2060 );
not \U$15234 ( \15611 , \15609 );
and \U$15235 ( \15612 , \15611 , \2061 );
nor \U$15236 ( \15613 , \15610 , \15612 );
and \U$15237 ( \15614 , \2607 , RIae78530_112);
and \U$15238 ( \15615 , RIae77c48_93, \2605 );
nor \U$15239 ( \15616 , \15614 , \15615 );
and \U$15240 ( \15617 , \15616 , \2397 );
not \U$15241 ( \15618 , \15616 );
and \U$15242 ( \15619 , \15618 , \2611 );
nor \U$15243 ( \15620 , \15617 , \15619 );
xor \U$15244 ( \15621 , \15613 , \15620 );
and \U$15245 ( \15622 , \1939 , RIae78008_101);
and \U$15246 ( \15623 , RIae781e8_105, \1937 );
nor \U$15247 ( \15624 , \15622 , \15623 );
and \U$15248 ( \15625 , \15624 , \1734 );
not \U$15249 ( \15626 , \15624 );
and \U$15250 ( \15627 , \15626 , \1735 );
nor \U$15251 ( \15628 , \15625 , \15627 );
and \U$15252 ( \15629 , \15621 , \15628 );
and \U$15253 ( \15630 , \15613 , \15620 );
nor \U$15254 ( \15631 , \15629 , \15630 );
and \U$15255 ( \15632 , \1138 , RIae77018_67);
and \U$15256 ( \15633 , RIae771f8_71, \1136 );
nor \U$15257 ( \15634 , \15632 , \15633 );
and \U$15258 ( \15635 , \15634 , \1142 );
not \U$15259 ( \15636 , \15634 );
and \U$15260 ( \15637 , \15636 , \1012 );
nor \U$15261 ( \15638 , \15635 , \15637 );
and \U$15262 ( \15639 , \1376 , RIae772e8_73);
and \U$15263 ( \15640 , RIae782d8_107, \1374 );
nor \U$15264 ( \15641 , \15639 , \15640 );
and \U$15265 ( \15642 , \15641 , \1261 );
not \U$15266 ( \15643 , \15641 );
and \U$15267 ( \15644 , \15643 , \1380 );
nor \U$15268 ( \15645 , \15642 , \15644 );
or \U$15269 ( \15646 , \15638 , \15645 );
not \U$15270 ( \15647 , \15645 );
not \U$15271 ( \15648 , \15638 );
or \U$15272 ( \15649 , \15647 , \15648 );
and \U$15273 ( \15650 , \1593 , RIae780f8_103);
and \U$15274 ( \15651 , RIae77f18_99, \1591 );
nor \U$15275 ( \15652 , \15650 , \15651 );
and \U$15276 ( \15653 , \15652 , \1498 );
not \U$15277 ( \15654 , \15652 );
and \U$15278 ( \15655 , \15654 , \1488 );
nor \U$15279 ( \15656 , \15653 , \15655 );
nand \U$15280 ( \15657 , \15649 , \15656 );
nand \U$15281 ( \15658 , \15646 , \15657 );
xor \U$15282 ( \15659 , \15631 , \15658 );
and \U$15283 ( \15660 , \2783 , RIae77b58_91);
and \U$15284 ( \15661 , RIae77d38_95, \2781 );
nor \U$15285 ( \15662 , \15660 , \15661 );
not \U$15286 ( \15663 , \15662 );
not \U$15287 ( \15664 , \3089 );
and \U$15288 ( \15665 , \15663 , \15664 );
and \U$15289 ( \15666 , \15662 , \2789 );
nor \U$15290 ( \15667 , \15665 , \15666 );
and \U$15291 ( \15668 , \3214 , RIae77e28_97);
and \U$15292 ( \15669 , RIae78968_121, \3212 );
nor \U$15293 ( \15670 , \15668 , \15669 );
not \U$15294 ( \15671 , \15670 );
not \U$15295 ( \15672 , \3218 );
and \U$15296 ( \15673 , \15671 , \15672 );
and \U$15297 ( \15674 , \15670 , \3218 );
nor \U$15298 ( \15675 , \15673 , \15674 );
or \U$15299 ( \15676 , \15667 , \15675 );
not \U$15300 ( \15677 , \15675 );
not \U$15301 ( \15678 , \15667 );
or \U$15302 ( \15679 , \15677 , \15678 );
and \U$15303 ( \15680 , \3730 , RIae78878_119);
and \U$15304 ( \15681 , RIae78788_117, \3728 );
nor \U$15305 ( \15682 , \15680 , \15681 );
and \U$15306 ( \15683 , \15682 , \3732 );
not \U$15307 ( \15684 , \15682 );
and \U$15308 ( \15685 , \15684 , \3422 );
nor \U$15309 ( \15686 , \15683 , \15685 );
nand \U$15310 ( \15687 , \15679 , \15686 );
nand \U$15311 ( \15688 , \15676 , \15687 );
and \U$15312 ( \15689 , \15659 , \15688 );
and \U$15313 ( \15690 , \15631 , \15658 );
or \U$15314 ( \15691 , \15689 , \15690 );
and \U$15315 ( \15692 , \12180 , RIae76208_37);
and \U$15316 ( \15693 , RIae76a78_55, \12178 );
nor \U$15317 ( \15694 , \15692 , \15693 );
and \U$15318 ( \15695 , \15694 , \11827 );
not \U$15319 ( \15696 , \15694 );
and \U$15320 ( \15697 , \15696 , \12184 );
nor \U$15321 ( \15698 , \15695 , \15697 );
and \U$15322 ( \15699 , \13059 , RIae76988_53);
and \U$15323 ( \15700 , RIae767a8_49, \13057 );
nor \U$15324 ( \15701 , \15699 , \15700 );
and \U$15325 ( \15702 , \15701 , \12718 );
not \U$15326 ( \15703 , \15701 );
and \U$15327 ( \15704 , \15703 , \13063 );
nor \U$15328 ( \15705 , \15702 , \15704 );
xor \U$15329 ( \15706 , \15698 , \15705 );
and \U$15330 ( \15707 , \14059 , RIae76898_51);
and \U$15331 ( \15708 , RIae76b68_57, \14057 );
nor \U$15332 ( \15709 , \15707 , \15708 );
and \U$15333 ( \15710 , \15709 , \14063 );
not \U$15334 ( \15711 , \15709 );
and \U$15335 ( \15712 , \15711 , \13502 );
nor \U$15336 ( \15713 , \15710 , \15712 );
and \U$15337 ( \15714 , \15706 , \15713 );
and \U$15338 ( \15715 , \15698 , \15705 );
or \U$15339 ( \15716 , \15714 , \15715 );
and \U$15340 ( \15717 , \14964 , RIae78a58_123);
and \U$15341 ( \15718 , RIae78cb0_128, \14962 );
nor \U$15342 ( \15719 , \15717 , \15718 );
and \U$15343 ( \15720 , \15719 , \14462 );
not \U$15344 ( \15721 , \15719 );
and \U$15345 ( \15722 , \15721 , \14463 );
nor \U$15346 ( \15723 , \15720 , \15722 );
not \U$15347 ( \15724 , \15723 );
not \U$15348 ( \15725 , RIae7aab0_192);
and \U$15349 ( \15726 , \15725 , RIae7aa38_191);
and \U$15350 ( \15727 , \15726 , RIae78da0_130);
nor \U$15351 ( \15728 , \15727 , \14959 );
nand \U$15352 ( \15729 , \15724 , \15728 );
or \U$15353 ( \15730 , \15716 , \15729 );
not \U$15354 ( \15731 , \15729 );
not \U$15355 ( \15732 , \15716 );
or \U$15356 ( \15733 , \15731 , \15732 );
and \U$15357 ( \15734 , \10548 , RIae765c8_45);
and \U$15358 ( \15735 , RIae76118_35, \10546 );
nor \U$15359 ( \15736 , \15734 , \15735 );
and \U$15360 ( \15737 , \15736 , \10118 );
not \U$15361 ( \15738 , \15736 );
and \U$15362 ( \15739 , \15738 , \10421 );
nor \U$15363 ( \15740 , \15737 , \15739 );
and \U$15364 ( \15741 , \11470 , RIae76028_33);
and \U$15365 ( \15742 , RIae762f8_39, \11468 );
nor \U$15366 ( \15743 , \15741 , \15742 );
and \U$15367 ( \15744 , \15743 , \11474 );
not \U$15368 ( \15745 , \15743 );
and \U$15369 ( \15746 , \15745 , \10936 );
nor \U$15370 ( \15747 , \15744 , \15746 );
xor \U$15371 ( \15748 , \15740 , \15747 );
and \U$15372 ( \15749 , \9760 , RIae764d8_43);
and \U$15373 ( \15750 , RIae766b8_47, \9758 );
nor \U$15374 ( \15751 , \15749 , \15750 );
and \U$15375 ( \15752 , \15751 , \9272 );
not \U$15376 ( \15753 , \15751 );
and \U$15377 ( \15754 , \15753 , \9273 );
nor \U$15378 ( \15755 , \15752 , \15754 );
and \U$15379 ( \15756 , \15748 , \15755 );
and \U$15380 ( \15757 , \15740 , \15747 );
nor \U$15381 ( \15758 , \15756 , \15757 );
nand \U$15382 ( \15759 , \15733 , \15758 );
nand \U$15383 ( \15760 , \15730 , \15759 );
xor \U$15384 ( \15761 , \15691 , \15760 );
and \U$15385 ( \15762 , \6172 , RIae75d58_27);
and \U$15386 ( \15763 , RIae755d8_11, \6170 );
nor \U$15387 ( \15764 , \15762 , \15763 );
and \U$15388 ( \15765 , \15764 , \6175 );
not \U$15389 ( \15766 , \15764 );
and \U$15390 ( \15767 , \15766 , \6176 );
nor \U$15391 ( \15768 , \15765 , \15767 );
and \U$15392 ( \15769 , \6941 , RIae754e8_9);
and \U$15393 ( \15770 , RIae757b8_15, \6939 );
nor \U$15394 ( \15771 , \15769 , \15770 );
and \U$15395 ( \15772 , \15771 , \6945 );
not \U$15396 ( \15773 , \15771 );
and \U$15397 ( \15774 , \15773 , \6314 );
nor \U$15398 ( \15775 , \15772 , \15774 );
xor \U$15399 ( \15776 , \15768 , \15775 );
and \U$15400 ( \15777 , \5896 , RIae75e48_29);
and \U$15401 ( \15778 , RIae75c68_25, \5894 );
nor \U$15402 ( \15779 , \15777 , \15778 );
and \U$15403 ( \15780 , \15779 , \5589 );
not \U$15404 ( \15781 , \15779 );
and \U$15405 ( \15782 , \15781 , \5590 );
nor \U$15406 ( \15783 , \15780 , \15782 );
and \U$15407 ( \15784 , \15776 , \15783 );
and \U$15408 ( \15785 , \15768 , \15775 );
nor \U$15409 ( \15786 , \15784 , \15785 );
and \U$15410 ( \15787 , \4688 , RIae75a88_21);
and \U$15411 ( \15788 , RIae75998_19, \4686 );
nor \U$15412 ( \15789 , \15787 , \15788 );
and \U$15413 ( \15790 , \15789 , \4482 );
not \U$15414 ( \15791 , \15789 );
and \U$15415 ( \15792 , \15791 , \4481 );
nor \U$15416 ( \15793 , \15790 , \15792 );
and \U$15417 ( \15794 , \5399 , RIae758a8_17);
and \U$15418 ( \15795 , RIae75f38_31, \5397 );
nor \U$15419 ( \15796 , \15794 , \15795 );
and \U$15420 ( \15797 , \15796 , \5403 );
not \U$15421 ( \15798 , \15796 );
and \U$15422 ( \15799 , \15798 , \5016 );
nor \U$15423 ( \15800 , \15797 , \15799 );
xor \U$15424 ( \15801 , \15793 , \15800 );
and \U$15425 ( \15802 , \4247 , RIae78698_115);
and \U$15426 ( \15803 , RIae75b78_23, \4245 );
nor \U$15427 ( \15804 , \15802 , \15803 );
and \U$15428 ( \15805 , \15804 , \4251 );
not \U$15429 ( \15806 , \15804 );
and \U$15430 ( \15807 , \15806 , \3989 );
nor \U$15431 ( \15808 , \15805 , \15807 );
and \U$15432 ( \15809 , \15801 , \15808 );
and \U$15433 ( \15810 , \15793 , \15800 );
nor \U$15434 ( \15811 , \15809 , \15810 );
xor \U$15435 ( \15812 , \15786 , \15811 );
and \U$15436 ( \15813 , \7633 , RIae756c8_13);
and \U$15437 ( \15814 , RIae75218_3, \7631 );
nor \U$15438 ( \15815 , \15813 , \15814 );
and \U$15439 ( \15816 , \15815 , \7205 );
not \U$15440 ( \15817 , \15815 );
and \U$15441 ( \15818 , \15817 , \7206 );
nor \U$15442 ( \15819 , \15816 , \15818 );
and \U$15443 ( \15820 , \8371 , RIae75128_1);
and \U$15444 ( \15821 , RIae75308_5, \8369 );
nor \U$15445 ( \15822 , \15820 , \15821 );
and \U$15446 ( \15823 , \15822 , \8019 );
not \U$15447 ( \15824 , \15822 );
and \U$15448 ( \15825 , \15824 , \8020 );
nor \U$15449 ( \15826 , \15823 , \15825 );
or \U$15450 ( \15827 , \15819 , \15826 );
not \U$15451 ( \15828 , \15826 );
not \U$15452 ( \15829 , \15819 );
or \U$15453 ( \15830 , \15828 , \15829 );
and \U$15454 ( \15831 , \8966 , RIae753f8_7);
and \U$15455 ( \15832 , RIae763e8_41, \8964 );
nor \U$15456 ( \15833 , \15831 , \15832 );
and \U$15457 ( \15834 , \15833 , \8799 );
not \U$15458 ( \15835 , \15833 );
and \U$15459 ( \15836 , \15835 , \8789 );
nor \U$15460 ( \15837 , \15834 , \15836 );
nand \U$15461 ( \15838 , \15830 , \15837 );
nand \U$15462 ( \15839 , \15827 , \15838 );
and \U$15463 ( \15840 , \15812 , \15839 );
and \U$15464 ( \15841 , \15786 , \15811 );
or \U$15465 ( \15842 , \15840 , \15841 );
and \U$15466 ( \15843 , \15761 , \15842 );
and \U$15467 ( \15844 , \15691 , \15760 );
or \U$15468 ( \15845 , \15843 , \15844 );
not \U$15469 ( \15846 , \15463 );
xor \U$15470 ( \15847 , \15481 , \15471 );
not \U$15471 ( \15848 , \15847 );
or \U$15472 ( \15849 , \15846 , \15848 );
or \U$15473 ( \15850 , \15847 , \15463 );
nand \U$15474 ( \15851 , \15849 , \15850 );
not \U$15475 ( \15852 , \15851 );
and \U$15476 ( \15853 , \15494 , RIae7aa38_191);
not \U$15477 ( \15854 , \15494 );
and \U$15478 ( \15855 , \15854 , \14959 );
nor \U$15479 ( \15856 , \15853 , \15855 );
not \U$15480 ( \15857 , \15856 );
not \U$15481 ( \15858 , \15503 );
and \U$15482 ( \15859 , \15857 , \15858 );
and \U$15483 ( \15860 , \15856 , \15503 );
nor \U$15484 ( \15861 , \15859 , \15860 );
nor \U$15485 ( \15862 , \15852 , \15861 );
xor \U$15486 ( \15863 , \14957 , \14969 );
xor \U$15487 ( \15864 , \15863 , \14977 );
xor \U$15488 ( \15865 , \15862 , \15864 );
not \U$15489 ( \15866 , \15279 );
not \U$15490 ( \15867 , \15290 );
or \U$15491 ( \15868 , \15866 , \15867 );
or \U$15492 ( \15869 , \15279 , \15290 );
nand \U$15493 ( \15870 , \15868 , \15869 );
not \U$15494 ( \15871 , \15870 );
not \U$15495 ( \15872 , \15272 );
and \U$15496 ( \15873 , \15871 , \15872 );
and \U$15497 ( \15874 , \15870 , \15272 );
nor \U$15498 ( \15875 , \15873 , \15874 );
xor \U$15499 ( \15876 , \15438 , \15445 );
xor \U$15500 ( \15877 , \15876 , \15453 );
or \U$15501 ( \15878 , \15875 , \15877 );
not \U$15502 ( \15879 , \15877 );
not \U$15503 ( \15880 , \15875 );
or \U$15504 ( \15881 , \15879 , \15880 );
xor \U$15505 ( \15882 , \15325 , \15332 );
xor \U$15506 ( \15883 , \15882 , \15340 );
nand \U$15507 ( \15884 , \15881 , \15883 );
nand \U$15508 ( \15885 , \15878 , \15884 );
and \U$15509 ( \15886 , \15865 , \15885 );
and \U$15510 ( \15887 , \15862 , \15864 );
or \U$15511 ( \15888 , \15886 , \15887 );
xor \U$15512 ( \15889 , \15845 , \15888 );
xor \U$15513 ( \15890 , \15229 , \15236 );
xor \U$15514 ( \15891 , \15890 , \15245 );
not \U$15515 ( \15892 , \15414 );
not \U$15516 ( \15893 , \15425 );
or \U$15517 ( \15894 , \15892 , \15893 );
or \U$15518 ( \15895 , \15414 , \15425 );
nand \U$15519 ( \15896 , \15894 , \15895 );
not \U$15520 ( \15897 , \15896 );
not \U$15521 ( \15898 , \15407 );
and \U$15522 ( \15899 , \15897 , \15898 );
and \U$15523 ( \15900 , \15896 , \15407 );
nor \U$15524 ( \15901 , \15899 , \15900 );
or \U$15525 ( \15902 , \15891 , \15901 );
not \U$15526 ( \15903 , \15901 );
not \U$15527 ( \15904 , \15891 );
or \U$15528 ( \15905 , \15903 , \15904 );
xor \U$15529 ( \15906 , \15205 , \15207 );
xor \U$15530 ( \15907 , \15906 , \15216 );
nand \U$15531 ( \15908 , \15905 , \15907 );
nand \U$15532 ( \15909 , \15902 , \15908 );
and \U$15533 ( \15910 , \384 , RIae774c8_77);
and \U$15534 ( \15911 , RIae77720_82, \382 );
nor \U$15535 ( \15912 , \15910 , \15911 );
not \U$15536 ( \15913 , \15912 );
not \U$15537 ( \15914 , \392 );
and \U$15538 ( \15915 , \15913 , \15914 );
and \U$15539 ( \15916 , \15912 , \392 );
nor \U$15540 ( \15917 , \15915 , \15916 );
and \U$15541 ( \15918 , \436 , RIae773d8_75);
and \U$15542 ( \15919 , RIae77a68_89, \434 );
nor \U$15543 ( \15920 , \15918 , \15919 );
not \U$15544 ( \15921 , \15920 );
not \U$15545 ( \15922 , \402 );
and \U$15546 ( \15923 , \15921 , \15922 );
and \U$15547 ( \15924 , \15920 , \400 );
nor \U$15548 ( \15925 , \15923 , \15924 );
or \U$15549 ( \15926 , \15917 , \15925 );
not \U$15550 ( \15927 , \15925 );
not \U$15551 ( \15928 , \15917 );
or \U$15552 ( \15929 , \15927 , \15928 );
not \U$15553 ( \15930 , \469 );
and \U$15554 ( \15931 , \514 , RIae77978_87);
and \U$15555 ( \15932 , RIae77798_83, \512 );
nor \U$15556 ( \15933 , \15931 , \15932 );
not \U$15557 ( \15934 , \15933 );
or \U$15558 ( \15935 , \15930 , \15934 );
or \U$15559 ( \15936 , \15933 , \471 );
nand \U$15560 ( \15937 , \15935 , \15936 );
nand \U$15561 ( \15938 , \15929 , \15937 );
nand \U$15562 ( \15939 , \15926 , \15938 );
and \U$15563 ( \15940 , \672 , RIae76e38_63);
and \U$15564 ( \15941 , RIae76d48_61, \670 );
nor \U$15565 ( \15942 , \15940 , \15941 );
and \U$15566 ( \15943 , \15942 , \587 );
not \U$15567 ( \15944 , \15942 );
and \U$15568 ( \15945 , \15944 , \588 );
nor \U$15569 ( \15946 , \15943 , \15945 );
and \U$15570 ( \15947 , \883 , RIae76c58_59);
and \U$15571 ( \15948 , RIae77180_70, \881 );
nor \U$15572 ( \15949 , \15947 , \15948 );
not \U$15573 ( \15950 , \15949 );
not \U$15574 ( \15951 , \789 );
and \U$15575 ( \15952 , \15950 , \15951 );
and \U$15576 ( \15953 , \15949 , \787 );
nor \U$15577 ( \15954 , \15952 , \15953 );
xor \U$15578 ( \15955 , \15946 , \15954 );
and \U$15579 ( \15956 , \558 , RIae77888_85);
and \U$15580 ( \15957 , RIae76f28_65, \556 );
nor \U$15581 ( \15958 , \15956 , \15957 );
and \U$15582 ( \15959 , \15958 , \562 );
not \U$15583 ( \15960 , \15958 );
and \U$15584 ( \15961 , \15960 , \504 );
nor \U$15585 ( \15962 , \15959 , \15961 );
and \U$15586 ( \15963 , \15955 , \15962 );
and \U$15587 ( \15964 , \15946 , \15954 );
nor \U$15588 ( \15965 , \15963 , \15964 );
nor \U$15589 ( \15966 , \15939 , \15965 );
not \U$15590 ( \15967 , \15966 );
xor \U$15591 ( \15968 , \15909 , \15967 );
xor \U$15592 ( \15969 , \15354 , \15361 );
xor \U$15593 ( \15970 , \15969 , \15370 );
xor \U$15594 ( \15971 , \15380 , \15387 );
xor \U$15595 ( \15972 , \15971 , \15395 );
and \U$15596 ( \15973 , \15970 , \15972 );
xor \U$15597 ( \15974 , \15299 , \15306 );
xor \U$15598 ( \15975 , \15974 , \15314 );
xor \U$15599 ( \15976 , \15380 , \15387 );
xor \U$15600 ( \15977 , \15976 , \15395 );
and \U$15601 ( \15978 , \15975 , \15977 );
and \U$15602 ( \15979 , \15970 , \15975 );
or \U$15603 ( \15980 , \15973 , \15978 , \15979 );
and \U$15604 ( \15981 , \15968 , \15980 );
and \U$15605 ( \15982 , \15909 , \15967 );
or \U$15606 ( \15983 , \15981 , \15982 );
and \U$15607 ( \15984 , \15889 , \15983 );
and \U$15608 ( \15985 , \15845 , \15888 );
or \U$15609 ( \15986 , \15984 , \15985 );
xor \U$15610 ( \15987 , \15606 , \15986 );
xor \U$15611 ( \15988 , \15197 , \15251 );
xor \U$15612 ( \15989 , \15988 , \15262 );
xor \U$15613 ( \15990 , \15524 , \15525 );
xor \U$15614 ( \15991 , \15990 , \15530 );
and \U$15615 ( \15992 , \15989 , \15991 );
xor \U$15616 ( \15993 , \14833 , \14835 );
xor \U$15617 ( \15994 , \15993 , \14838 );
xor \U$15618 ( \15995 , \15539 , \15546 );
xor \U$15619 ( \15996 , \15994 , \15995 );
xor \U$15620 ( \15997 , \15524 , \15525 );
xor \U$15621 ( \15998 , \15997 , \15530 );
and \U$15622 ( \15999 , \15996 , \15998 );
and \U$15623 ( \16000 , \15989 , \15996 );
or \U$15624 ( \16001 , \15992 , \15999 , \16000 );
and \U$15625 ( \16002 , \15987 , \16001 );
and \U$15626 ( \16003 , \15606 , \15986 );
or \U$15627 ( \16004 , \16002 , \16003 );
xor \U$15628 ( \16005 , \14844 , \15093 );
xor \U$15629 ( \16006 , \16005 , \15119 );
xor \U$15630 ( \16007 , \16004 , \16006 );
xor \U$15631 ( \16008 , \14925 , \15009 );
xor \U$15632 ( \16009 , \16008 , \15090 );
xor \U$15633 ( \16010 , \15551 , \15563 );
xor \U$15634 ( \16011 , \16010 , \15568 );
and \U$15635 ( \16012 , \16009 , \16011 );
xor \U$15636 ( \16013 , \15106 , \15111 );
xor \U$15637 ( \16014 , \16013 , \15116 );
xor \U$15638 ( \16015 , \15173 , \15180 );
xor \U$15639 ( \16016 , \16014 , \16015 );
xor \U$15640 ( \16017 , \15551 , \15563 );
xor \U$15641 ( \16018 , \16017 , \15568 );
and \U$15642 ( \16019 , \16016 , \16018 );
and \U$15643 ( \16020 , \16009 , \16016 );
or \U$15644 ( \16021 , \16012 , \16019 , \16020 );
xor \U$15645 ( \16022 , \16007 , \16021 );
and \U$15646 ( \16023 , \15572 , \16022 );
xor \U$15647 ( \16024 , \15606 , \15986 );
xor \U$15648 ( \16025 , \16024 , \16001 );
xor \U$15649 ( \16026 , \15551 , \15563 );
xor \U$15650 ( \16027 , \16026 , \15568 );
xor \U$15651 ( \16028 , \16009 , \16016 );
xor \U$15652 ( \16029 , \16027 , \16028 );
and \U$15653 ( \16030 , \16025 , \16029 );
xor \U$15654 ( \16031 , \14749 , \14761 );
xor \U$15655 ( \16032 , \16031 , \14766 );
xor \U$15656 ( \16033 , \14428 , \14503 );
xor \U$15657 ( \16034 , \16033 , \14584 );
xor \U$15658 ( \16035 , \14600 , \14633 );
xor \U$15659 ( \16036 , \16035 , \14646 );
xor \U$15660 ( \16037 , \15125 , \15132 );
xor \U$15661 ( \16038 , \16036 , \16037 );
xor \U$15662 ( \16039 , \16034 , \16038 );
xor \U$15663 ( \16040 , \16032 , \16039 );
xor \U$15664 ( \16041 , \16030 , \16040 );
xor \U$15665 ( \16042 , \15786 , \15811 );
xor \U$15666 ( \16043 , \16042 , \15839 );
xor \U$15667 ( \16044 , \15631 , \15658 );
xor \U$15668 ( \16045 , \16044 , \15688 );
and \U$15669 ( \16046 , \16043 , \16045 );
not \U$15670 ( \16047 , \16045 );
not \U$15671 ( \16048 , \16043 );
and \U$15672 ( \16049 , \16047 , \16048 );
not \U$15673 ( \16050 , \15758 );
not \U$15674 ( \16051 , \15716 );
or \U$15675 ( \16052 , \16050 , \16051 );
or \U$15676 ( \16053 , \15716 , \15758 );
nand \U$15677 ( \16054 , \16052 , \16053 );
not \U$15678 ( \16055 , \16054 );
not \U$15679 ( \16056 , \15729 );
and \U$15680 ( \16057 , \16055 , \16056 );
and \U$15681 ( \16058 , \16054 , \15729 );
nor \U$15682 ( \16059 , \16057 , \16058 );
nor \U$15683 ( \16060 , \16049 , \16059 );
nor \U$15684 ( \16061 , \16046 , \16060 );
not \U$15685 ( \16062 , \15506 );
not \U$15686 ( \16063 , \15483 );
or \U$15687 ( \16064 , \16062 , \16063 );
or \U$15688 ( \16065 , \15483 , \15506 );
nand \U$15689 ( \16066 , \16064 , \16065 );
not \U$15690 ( \16067 , \16066 );
not \U$15691 ( \16068 , \15456 );
and \U$15692 ( \16069 , \16067 , \16068 );
and \U$15693 ( \16070 , \16066 , \15456 );
nor \U$15694 ( \16071 , \16069 , \16070 );
or \U$15695 ( \16072 , \16061 , \16071 );
not \U$15696 ( \16073 , \16071 );
not \U$15697 ( \16074 , \16061 );
or \U$15698 ( \16075 , \16073 , \16074 );
not \U$15699 ( \16076 , \15891 );
not \U$15700 ( \16077 , \15907 );
or \U$15701 ( \16078 , \16076 , \16077 );
or \U$15702 ( \16079 , \15907 , \15891 );
nand \U$15703 ( \16080 , \16078 , \16079 );
not \U$15704 ( \16081 , \16080 );
not \U$15705 ( \16082 , \15901 );
and \U$15706 ( \16083 , \16081 , \16082 );
and \U$15707 ( \16084 , \16080 , \15901 );
nor \U$15708 ( \16085 , \16083 , \16084 );
and \U$15709 ( \16086 , \15939 , \15965 );
nor \U$15710 ( \16087 , \16086 , \15966 );
or \U$15711 ( \16088 , \16085 , \16087 );
not \U$15712 ( \16089 , \16087 );
not \U$15713 ( \16090 , \16085 );
or \U$15714 ( \16091 , \16089 , \16090 );
xor \U$15715 ( \16092 , \15380 , \15387 );
xor \U$15716 ( \16093 , \16092 , \15395 );
xor \U$15717 ( \16094 , \15970 , \15975 );
xor \U$15718 ( \16095 , \16093 , \16094 );
nand \U$15719 ( \16096 , \16091 , \16095 );
nand \U$15720 ( \16097 , \16088 , \16096 );
nand \U$15721 ( \16098 , \16075 , \16097 );
nand \U$15722 ( \16099 , \16072 , \16098 );
not \U$15723 ( \16100 , \2774 );
and \U$15724 ( \16101 , \3214 , RIae77d38_95);
and \U$15725 ( \16102 , RIae77e28_97, \3212 );
nor \U$15726 ( \16103 , \16101 , \16102 );
not \U$15727 ( \16104 , \16103 );
or \U$15728 ( \16105 , \16100 , \16104 );
or \U$15729 ( \16106 , \16103 , \3218 );
nand \U$15730 ( \16107 , \16105 , \16106 );
and \U$15731 ( \16108 , \2607 , RIae783c8_109);
and \U$15732 ( \16109 , RIae78530_112, \2605 );
nor \U$15733 ( \16110 , \16108 , \16109 );
and \U$15734 ( \16111 , \16110 , \2611 );
not \U$15735 ( \16112 , \16110 );
and \U$15736 ( \16113 , \16112 , \2397 );
nor \U$15737 ( \16114 , \16111 , \16113 );
xor \U$15738 ( \16115 , \16107 , \16114 );
not \U$15739 ( \16116 , \2789 );
and \U$15740 ( \16117 , \2783 , RIae77c48_93);
and \U$15741 ( \16118 , RIae77b58_91, \2781 );
nor \U$15742 ( \16119 , \16117 , \16118 );
not \U$15743 ( \16120 , \16119 );
or \U$15744 ( \16121 , \16116 , \16120 );
or \U$15745 ( \16122 , \16119 , \2789 );
nand \U$15746 ( \16123 , \16121 , \16122 );
and \U$15747 ( \16124 , \16115 , \16123 );
and \U$15748 ( \16125 , \16107 , \16114 );
or \U$15749 ( \16126 , \16124 , \16125 );
and \U$15750 ( \16127 , \2224 , RIae781e8_105);
and \U$15751 ( \16128 , RIae785a8_113, \2222 );
nor \U$15752 ( \16129 , \16127 , \16128 );
and \U$15753 ( \16130 , \16129 , \2061 );
not \U$15754 ( \16131 , \16129 );
and \U$15755 ( \16132 , \16131 , \2060 );
nor \U$15756 ( \16133 , \16130 , \16132 );
and \U$15757 ( \16134 , \1593 , RIae782d8_107);
and \U$15758 ( \16135 , RIae780f8_103, \1591 );
nor \U$15759 ( \16136 , \16134 , \16135 );
and \U$15760 ( \16137 , \16136 , \1498 );
not \U$15761 ( \16138 , \16136 );
and \U$15762 ( \16139 , \16138 , \1488 );
nor \U$15763 ( \16140 , \16137 , \16139 );
xor \U$15764 ( \16141 , \16133 , \16140 );
and \U$15765 ( \16142 , \1939 , RIae77f18_99);
and \U$15766 ( \16143 , RIae78008_101, \1937 );
nor \U$15767 ( \16144 , \16142 , \16143 );
and \U$15768 ( \16145 , \16144 , \1735 );
not \U$15769 ( \16146 , \16144 );
and \U$15770 ( \16147 , \16146 , \1734 );
nor \U$15771 ( \16148 , \16145 , \16147 );
and \U$15772 ( \16149 , \16141 , \16148 );
and \U$15773 ( \16150 , \16133 , \16140 );
or \U$15774 ( \16151 , \16149 , \16150 );
xor \U$15775 ( \16152 , \16126 , \16151 );
and \U$15776 ( \16153 , \1376 , RIae771f8_71);
and \U$15777 ( \16154 , RIae772e8_73, \1374 );
nor \U$15778 ( \16155 , \16153 , \16154 );
and \U$15779 ( \16156 , \16155 , \1380 );
not \U$15780 ( \16157 , \16155 );
and \U$15781 ( \16158 , \16157 , \1261 );
nor \U$15782 ( \16159 , \16156 , \16158 );
not \U$15783 ( \16160 , \787 );
and \U$15784 ( \16161 , \883 , RIae76d48_61);
and \U$15785 ( \16162 , RIae76c58_59, \881 );
nor \U$15786 ( \16163 , \16161 , \16162 );
not \U$15787 ( \16164 , \16163 );
or \U$15788 ( \16165 , \16160 , \16164 );
or \U$15789 ( \16166 , \16163 , \787 );
nand \U$15790 ( \16167 , \16165 , \16166 );
xor \U$15791 ( \16168 , \16159 , \16167 );
and \U$15792 ( \16169 , \1138 , RIae77180_70);
and \U$15793 ( \16170 , RIae77018_67, \1136 );
nor \U$15794 ( \16171 , \16169 , \16170 );
and \U$15795 ( \16172 , \16171 , \1012 );
not \U$15796 ( \16173 , \16171 );
and \U$15797 ( \16174 , \16173 , \1142 );
nor \U$15798 ( \16175 , \16172 , \16174 );
and \U$15799 ( \16176 , \16168 , \16175 );
and \U$15800 ( \16177 , \16159 , \16167 );
or \U$15801 ( \16178 , \16176 , \16177 );
and \U$15802 ( \16179 , \16152 , \16178 );
and \U$15803 ( \16180 , \16126 , \16151 );
nor \U$15804 ( \16181 , \16179 , \16180 );
not \U$15805 ( \16182 , \16181 );
and \U$15806 ( \16183 , \6941 , RIae755d8_11);
and \U$15807 ( \16184 , RIae754e8_9, \6939 );
nor \U$15808 ( \16185 , \16183 , \16184 );
and \U$15809 ( \16186 , \16185 , \6945 );
not \U$15810 ( \16187 , \16185 );
and \U$15811 ( \16188 , \16187 , \6314 );
nor \U$15812 ( \16189 , \16186 , \16188 );
not \U$15813 ( \16190 , \16189 );
and \U$15814 ( \16191 , \7633 , RIae757b8_15);
and \U$15815 ( \16192 , RIae756c8_13, \7631 );
nor \U$15816 ( \16193 , \16191 , \16192 );
and \U$15817 ( \16194 , \16193 , \7205 );
not \U$15818 ( \16195 , \16193 );
and \U$15819 ( \16196 , \16195 , \7206 );
nor \U$15820 ( \16197 , \16194 , \16196 );
not \U$15821 ( \16198 , \16197 );
and \U$15822 ( \16199 , \16190 , \16198 );
and \U$15823 ( \16200 , \16197 , \16189 );
and \U$15824 ( \16201 , \8371 , RIae75218_3);
and \U$15825 ( \16202 , RIae75128_1, \8369 );
nor \U$15826 ( \16203 , \16201 , \16202 );
and \U$15827 ( \16204 , \16203 , \8019 );
not \U$15828 ( \16205 , \16203 );
and \U$15829 ( \16206 , \16205 , \8020 );
nor \U$15830 ( \16207 , \16204 , \16206 );
nor \U$15831 ( \16208 , \16200 , \16207 );
nor \U$15832 ( \16209 , \16199 , \16208 );
and \U$15833 ( \16210 , \5399 , RIae75998_19);
and \U$15834 ( \16211 , RIae758a8_17, \5397 );
nor \U$15835 ( \16212 , \16210 , \16211 );
and \U$15836 ( \16213 , \16212 , \5403 );
not \U$15837 ( \16214 , \16212 );
and \U$15838 ( \16215 , \16214 , \5016 );
nor \U$15839 ( \16216 , \16213 , \16215 );
not \U$15840 ( \16217 , \16216 );
and \U$15841 ( \16218 , \5896 , RIae75f38_31);
and \U$15842 ( \16219 , RIae75e48_29, \5894 );
nor \U$15843 ( \16220 , \16218 , \16219 );
and \U$15844 ( \16221 , \16220 , \5589 );
not \U$15845 ( \16222 , \16220 );
and \U$15846 ( \16223 , \16222 , \5590 );
nor \U$15847 ( \16224 , \16221 , \16223 );
not \U$15848 ( \16225 , \16224 );
and \U$15849 ( \16226 , \16217 , \16225 );
and \U$15850 ( \16227 , \16224 , \16216 );
and \U$15851 ( \16228 , \6172 , RIae75c68_25);
and \U$15852 ( \16229 , RIae75d58_27, \6170 );
nor \U$15853 ( \16230 , \16228 , \16229 );
and \U$15854 ( \16231 , \16230 , \6175 );
not \U$15855 ( \16232 , \16230 );
and \U$15856 ( \16233 , \16232 , \6176 );
nor \U$15857 ( \16234 , \16231 , \16233 );
nor \U$15858 ( \16235 , \16227 , \16234 );
nor \U$15859 ( \16236 , \16226 , \16235 );
xor \U$15860 ( \16237 , \16209 , \16236 );
and \U$15861 ( \16238 , \3730 , RIae78968_121);
and \U$15862 ( \16239 , RIae78878_119, \3728 );
nor \U$15863 ( \16240 , \16238 , \16239 );
and \U$15864 ( \16241 , \16240 , \3422 );
not \U$15865 ( \16242 , \16240 );
and \U$15866 ( \16243 , \16242 , \3732 );
nor \U$15867 ( \16244 , \16241 , \16243 );
not \U$15868 ( \16245 , \16244 );
and \U$15869 ( \16246 , \4247 , RIae78788_117);
and \U$15870 ( \16247 , RIae78698_115, \4245 );
nor \U$15871 ( \16248 , \16246 , \16247 );
and \U$15872 ( \16249 , \16248 , \4251 );
not \U$15873 ( \16250 , \16248 );
and \U$15874 ( \16251 , \16250 , \3989 );
nor \U$15875 ( \16252 , \16249 , \16251 );
not \U$15876 ( \16253 , \16252 );
and \U$15877 ( \16254 , \16245 , \16253 );
and \U$15878 ( \16255 , \16252 , \16244 );
and \U$15879 ( \16256 , \4688 , RIae75b78_23);
and \U$15880 ( \16257 , RIae75a88_21, \4686 );
nor \U$15881 ( \16258 , \16256 , \16257 );
and \U$15882 ( \16259 , \16258 , \4482 );
not \U$15883 ( \16260 , \16258 );
and \U$15884 ( \16261 , \16260 , \4481 );
nor \U$15885 ( \16262 , \16259 , \16261 );
nor \U$15886 ( \16263 , \16255 , \16262 );
nor \U$15887 ( \16264 , \16254 , \16263 );
and \U$15888 ( \16265 , \16237 , \16264 );
and \U$15889 ( \16266 , \16209 , \16236 );
or \U$15890 ( \16267 , \16265 , \16266 );
not \U$15891 ( \16268 , \16267 );
and \U$15892 ( \16269 , \16182 , \16268 );
and \U$15893 ( \16270 , \16181 , \16267 );
and \U$15894 ( \16271 , \13059 , RIae76a78_55);
and \U$15895 ( \16272 , RIae76988_53, \13057 );
nor \U$15896 ( \16273 , \16271 , \16272 );
and \U$15897 ( \16274 , \16273 , \13063 );
not \U$15898 ( \16275 , \16273 );
and \U$15899 ( \16276 , \16275 , \12718 );
nor \U$15900 ( \16277 , \16274 , \16276 );
and \U$15901 ( \16278 , \11470 , RIae76118_35);
and \U$15902 ( \16279 , RIae76028_33, \11468 );
nor \U$15903 ( \16280 , \16278 , \16279 );
and \U$15904 ( \16281 , \16280 , \10936 );
not \U$15905 ( \16282 , \16280 );
and \U$15906 ( \16283 , \16282 , \11474 );
nor \U$15907 ( \16284 , \16281 , \16283 );
xor \U$15908 ( \16285 , \16277 , \16284 );
and \U$15909 ( \16286 , \12180 , RIae762f8_39);
and \U$15910 ( \16287 , RIae76208_37, \12178 );
nor \U$15911 ( \16288 , \16286 , \16287 );
and \U$15912 ( \16289 , \16288 , \12184 );
not \U$15913 ( \16290 , \16288 );
and \U$15914 ( \16291 , \16290 , \11827 );
nor \U$15915 ( \16292 , \16289 , \16291 );
and \U$15916 ( \16293 , \16285 , \16292 );
and \U$15917 ( \16294 , \16277 , \16284 );
or \U$15918 ( \16295 , \16293 , \16294 );
and \U$15919 ( \16296 , \10548 , RIae766b8_47);
and \U$15920 ( \16297 , RIae765c8_45, \10546 );
nor \U$15921 ( \16298 , \16296 , \16297 );
and \U$15922 ( \16299 , \16298 , \10421 );
not \U$15923 ( \16300 , \16298 );
and \U$15924 ( \16301 , \16300 , \10118 );
nor \U$15925 ( \16302 , \16299 , \16301 );
and \U$15926 ( \16303 , \8966 , RIae75308_5);
and \U$15927 ( \16304 , RIae753f8_7, \8964 );
nor \U$15928 ( \16305 , \16303 , \16304 );
and \U$15929 ( \16306 , \16305 , \8799 );
not \U$15930 ( \16307 , \16305 );
and \U$15931 ( \16308 , \16307 , \8789 );
nor \U$15932 ( \16309 , \16306 , \16308 );
xor \U$15933 ( \16310 , \16302 , \16309 );
and \U$15934 ( \16311 , \9760 , RIae763e8_41);
and \U$15935 ( \16312 , RIae764d8_43, \9758 );
nor \U$15936 ( \16313 , \16311 , \16312 );
and \U$15937 ( \16314 , \16313 , \9273 );
not \U$15938 ( \16315 , \16313 );
and \U$15939 ( \16316 , \16315 , \9764 );
nor \U$15940 ( \16317 , \16314 , \16316 );
and \U$15941 ( \16318 , \16310 , \16317 );
and \U$15942 ( \16319 , \16302 , \16309 );
or \U$15943 ( \16320 , \16318 , \16319 );
xor \U$15944 ( \16321 , \16295 , \16320 );
and \U$15945 ( \16322 , \14059 , RIae767a8_49);
and \U$15946 ( \16323 , RIae76898_51, \14057 );
nor \U$15947 ( \16324 , \16322 , \16323 );
and \U$15948 ( \16325 , \16324 , \14063 );
not \U$15949 ( \16326 , \16324 );
and \U$15950 ( \16327 , \16326 , \13502 );
nor \U$15951 ( \16328 , \16325 , \16327 );
and \U$15952 ( \16329 , \15726 , RIae78cb0_128);
and \U$15953 ( \16330 , RIae7aab0_192, RIae78da0_130);
nor \U$15954 ( \16331 , \16329 , \16330 );
and \U$15955 ( \16332 , \16331 , RIae7aa38_191);
not \U$15956 ( \16333 , \16331 );
and \U$15957 ( \16334 , \16333 , \14959 );
nor \U$15958 ( \16335 , \16332 , \16334 );
or \U$15959 ( \16336 , \16328 , \16335 );
not \U$15960 ( \16337 , \16335 );
not \U$15961 ( \16338 , \16328 );
or \U$15962 ( \16339 , \16337 , \16338 );
and \U$15963 ( \16340 , \14964 , RIae76b68_57);
and \U$15964 ( \16341 , RIae78a58_123, \14962 );
nor \U$15965 ( \16342 , \16340 , \16341 );
and \U$15966 ( \16343 , \16342 , \14463 );
not \U$15967 ( \16344 , \16342 );
and \U$15968 ( \16345 , \16344 , \14462 );
nor \U$15969 ( \16346 , \16343 , \16345 );
nand \U$15970 ( \16347 , \16339 , \16346 );
nand \U$15971 ( \16348 , \16336 , \16347 );
and \U$15972 ( \16349 , \16321 , \16348 );
and \U$15973 ( \16350 , \16295 , \16320 );
nor \U$15974 ( \16351 , \16349 , \16350 );
nor \U$15975 ( \16352 , \16270 , \16351 );
nor \U$15976 ( \16353 , \16269 , \16352 );
not \U$15977 ( \16354 , \15645 );
not \U$15978 ( \16355 , \15656 );
or \U$15979 ( \16356 , \16354 , \16355 );
or \U$15980 ( \16357 , \15645 , \15656 );
nand \U$15981 ( \16358 , \16356 , \16357 );
not \U$15982 ( \16359 , \16358 );
not \U$15983 ( \16360 , \15638 );
and \U$15984 ( \16361 , \16359 , \16360 );
and \U$15985 ( \16362 , \16358 , \15638 );
nor \U$15986 ( \16363 , \16361 , \16362 );
not \U$15987 ( \16364 , \16363 );
xor \U$15988 ( \16365 , \15613 , \15620 );
xor \U$15989 ( \16366 , \16365 , \15628 );
not \U$15990 ( \16367 , \16366 );
and \U$15991 ( \16368 , \16364 , \16367 );
and \U$15992 ( \16369 , \16366 , \16363 );
xor \U$15993 ( \16370 , \15946 , \15954 );
xor \U$15994 ( \16371 , \16370 , \15962 );
nor \U$15995 ( \16372 , \16369 , \16371 );
nor \U$15996 ( \16373 , \16368 , \16372 );
and \U$15997 ( \16374 , \514 , RIae77a68_89);
and \U$15998 ( \16375 , RIae77978_87, \512 );
nor \U$15999 ( \16376 , \16374 , \16375 );
not \U$16000 ( \16377 , \16376 );
not \U$16001 ( \16378 , \471 );
and \U$16002 ( \16379 , \16377 , \16378 );
and \U$16003 ( \16380 , \16376 , \469 );
nor \U$16004 ( \16381 , \16379 , \16380 );
not \U$16005 ( \16382 , \16381 );
and \U$16006 ( \16383 , \558 , RIae77798_83);
and \U$16007 ( \16384 , RIae77888_85, \556 );
nor \U$16008 ( \16385 , \16383 , \16384 );
and \U$16009 ( \16386 , \16385 , \562 );
not \U$16010 ( \16387 , \16385 );
and \U$16011 ( \16388 , \16387 , \504 );
nor \U$16012 ( \16389 , \16386 , \16388 );
not \U$16013 ( \16390 , \16389 );
and \U$16014 ( \16391 , \16382 , \16390 );
and \U$16015 ( \16392 , \16389 , \16381 );
and \U$16016 ( \16393 , \672 , RIae76f28_65);
and \U$16017 ( \16394 , RIae76e38_63, \670 );
nor \U$16018 ( \16395 , \16393 , \16394 );
and \U$16019 ( \16396 , \16395 , \587 );
not \U$16020 ( \16397 , \16395 );
and \U$16021 ( \16398 , \16397 , \588 );
nor \U$16022 ( \16399 , \16396 , \16398 );
nor \U$16023 ( \16400 , \16392 , \16399 );
nor \U$16024 ( \16401 , \16391 , \16400 );
nand \U$16025 ( \16402 , RIae775b8_79, RIae78b48_125);
xor \U$16026 ( \16403 , \16401 , \16402 );
not \U$16027 ( \16404 , \15925 );
not \U$16028 ( \16405 , \15937 );
or \U$16029 ( \16406 , \16404 , \16405 );
or \U$16030 ( \16407 , \15925 , \15937 );
nand \U$16031 ( \16408 , \16406 , \16407 );
not \U$16032 ( \16409 , \16408 );
not \U$16033 ( \16410 , \15917 );
and \U$16034 ( \16411 , \16409 , \16410 );
and \U$16035 ( \16412 , \16408 , \15917 );
nor \U$16036 ( \16413 , \16411 , \16412 );
and \U$16037 ( \16414 , \16403 , \16413 );
and \U$16038 ( \16415 , \16401 , \16402 );
or \U$16039 ( \16416 , \16414 , \16415 );
xor \U$16040 ( \16417 , \16373 , \16416 );
not \U$16041 ( \16418 , \15675 );
not \U$16042 ( \16419 , \15686 );
or \U$16043 ( \16420 , \16418 , \16419 );
or \U$16044 ( \16421 , \15675 , \15686 );
nand \U$16045 ( \16422 , \16420 , \16421 );
not \U$16046 ( \16423 , \16422 );
not \U$16047 ( \16424 , \15667 );
and \U$16048 ( \16425 , \16423 , \16424 );
and \U$16049 ( \16426 , \16422 , \15667 );
nor \U$16050 ( \16427 , \16425 , \16426 );
xor \U$16051 ( \16428 , \15793 , \15800 );
xor \U$16052 ( \16429 , \16428 , \15808 );
xor \U$16053 ( \16430 , \16427 , \16429 );
xor \U$16054 ( \16431 , \15768 , \15775 );
xor \U$16055 ( \16432 , \16431 , \15783 );
and \U$16056 ( \16433 , \16430 , \16432 );
and \U$16057 ( \16434 , \16427 , \16429 );
or \U$16058 ( \16435 , \16433 , \16434 );
and \U$16059 ( \16436 , \16417 , \16435 );
and \U$16060 ( \16437 , \16373 , \16416 );
or \U$16061 ( \16438 , \16436 , \16437 );
xor \U$16062 ( \16439 , \16353 , \16438 );
xor \U$16063 ( \16440 , \15740 , \15747 );
xor \U$16064 ( \16441 , \16440 , \15755 );
not \U$16065 ( \16442 , \15826 );
not \U$16066 ( \16443 , \15837 );
or \U$16067 ( \16444 , \16442 , \16443 );
or \U$16068 ( \16445 , \15826 , \15837 );
nand \U$16069 ( \16446 , \16444 , \16445 );
not \U$16070 ( \16447 , \16446 );
not \U$16071 ( \16448 , \15819 );
and \U$16072 ( \16449 , \16447 , \16448 );
and \U$16073 ( \16450 , \16446 , \15819 );
nor \U$16074 ( \16451 , \16449 , \16450 );
xor \U$16075 ( \16452 , \16441 , \16451 );
xor \U$16076 ( \16453 , \15698 , \15705 );
xor \U$16077 ( \16454 , \16453 , \15713 );
and \U$16078 ( \16455 , \16452 , \16454 );
and \U$16079 ( \16456 , \16441 , \16451 );
or \U$16080 ( \16457 , \16455 , \16456 );
not \U$16081 ( \16458 , \15861 );
not \U$16082 ( \16459 , \15851 );
and \U$16083 ( \16460 , \16458 , \16459 );
and \U$16084 ( \16461 , \15861 , \15851 );
nor \U$16085 ( \16462 , \16460 , \16461 );
xor \U$16086 ( \16463 , \16457 , \16462 );
not \U$16087 ( \16464 , \15877 );
not \U$16088 ( \16465 , \15883 );
or \U$16089 ( \16466 , \16464 , \16465 );
or \U$16090 ( \16467 , \15877 , \15883 );
nand \U$16091 ( \16468 , \16466 , \16467 );
not \U$16092 ( \16469 , \16468 );
not \U$16093 ( \16470 , \15875 );
and \U$16094 ( \16471 , \16469 , \16470 );
and \U$16095 ( \16472 , \16468 , \15875 );
nor \U$16096 ( \16473 , \16471 , \16472 );
and \U$16097 ( \16474 , \16463 , \16473 );
and \U$16098 ( \16475 , \16457 , \16462 );
or \U$16099 ( \16476 , \16474 , \16475 );
and \U$16100 ( \16477 , \16439 , \16476 );
and \U$16101 ( \16478 , \16353 , \16438 );
nor \U$16102 ( \16479 , \16477 , \16478 );
xor \U$16103 ( \16480 , \16099 , \16479 );
xor \U$16104 ( \16481 , \15862 , \15864 );
xor \U$16105 ( \16482 , \16481 , \15885 );
xor \U$16106 ( \16483 , \15590 , \15592 );
xor \U$16107 ( \16484 , \16483 , \15595 );
and \U$16108 ( \16485 , \16482 , \16484 );
xor \U$16109 ( \16486 , \15254 , \15256 );
xor \U$16110 ( \16487 , \16486 , \15259 );
xor \U$16111 ( \16488 , \15576 , \15583 );
xor \U$16112 ( \16489 , \16487 , \16488 );
xor \U$16113 ( \16490 , \15590 , \15592 );
xor \U$16114 ( \16491 , \16490 , \15595 );
and \U$16115 ( \16492 , \16489 , \16491 );
and \U$16116 ( \16493 , \16482 , \16489 );
or \U$16117 ( \16494 , \16485 , \16492 , \16493 );
and \U$16118 ( \16495 , \16480 , \16494 );
and \U$16119 ( \16496 , \16099 , \16479 );
or \U$16120 ( \16497 , \16495 , \16496 );
xor \U$16121 ( \16498 , \15265 , \15511 );
xor \U$16122 ( \16499 , \16498 , \15533 );
xor \U$16123 ( \16500 , \16497 , \16499 );
xor \U$16124 ( \16501 , \15346 , \15430 );
xor \U$16125 ( \16502 , \16501 , \15508 );
xor \U$16126 ( \16503 , \15588 , \15598 );
xor \U$16127 ( \16504 , \16503 , \15603 );
and \U$16128 ( \16505 , \16502 , \16504 );
xor \U$16129 ( \16506 , \15524 , \15525 );
xor \U$16130 ( \16507 , \16506 , \15530 );
xor \U$16131 ( \16508 , \15989 , \15996 );
xor \U$16132 ( \16509 , \16507 , \16508 );
xor \U$16133 ( \16510 , \15588 , \15598 );
xor \U$16134 ( \16511 , \16510 , \15603 );
and \U$16135 ( \16512 , \16509 , \16511 );
and \U$16136 ( \16513 , \16502 , \16509 );
or \U$16137 ( \16514 , \16505 , \16512 , \16513 );
and \U$16138 ( \16515 , \16500 , \16514 );
and \U$16139 ( \16516 , \16497 , \16499 );
or \U$16140 ( \16517 , \16515 , \16516 );
and \U$16141 ( \16518 , \16041 , \16517 );
and \U$16142 ( \16519 , \16030 , \16040 );
or \U$16143 ( \16520 , \16518 , \16519 );
xor \U$16144 ( \16521 , \16023 , \16520 );
xor \U$16145 ( \16522 , \15142 , \15144 );
xor \U$16146 ( \16523 , \16522 , \15147 );
xor \U$16147 ( \16524 , \14347 , \14587 );
xor \U$16148 ( \16525 , \16524 , \14649 );
xor \U$16149 ( \16526 , \16523 , \16525 );
xor \U$16150 ( \16527 , \14769 , \15122 );
xor \U$16151 ( \16528 , \16527 , \15137 );
xor \U$16152 ( \16529 , \16526 , \16528 );
xor \U$16153 ( \16530 , \16004 , \16006 );
and \U$16154 ( \16531 , \16530 , \16021 );
and \U$16155 ( \16532 , \16004 , \16006 );
or \U$16156 ( \16533 , \16531 , \16532 );
xor \U$16157 ( \16534 , \15185 , \15536 );
and \U$16158 ( \16535 , \16534 , \15571 );
and \U$16159 ( \16536 , \15185 , \15536 );
or \U$16160 ( \16537 , \16535 , \16536 );
xor \U$16161 ( \16538 , \14303 , \14309 );
xor \U$16162 ( \16539 , \16538 , \14322 );
xor \U$16163 ( \16540 , \16537 , \16539 );
xor \U$16164 ( \16541 , \14749 , \14761 );
xor \U$16165 ( \16542 , \16541 , \14766 );
and \U$16166 ( \16543 , \16034 , \16542 );
xor \U$16167 ( \16544 , \14749 , \14761 );
xor \U$16168 ( \16545 , \16544 , \14766 );
and \U$16169 ( \16546 , \16038 , \16545 );
and \U$16170 ( \16547 , \16034 , \16038 );
or \U$16171 ( \16548 , \16543 , \16546 , \16547 );
xor \U$16172 ( \16549 , \16540 , \16548 );
xor \U$16173 ( \16550 , \16533 , \16549 );
xor \U$16174 ( \16551 , \16529 , \16550 );
and \U$16175 ( \16552 , \16521 , \16551 );
and \U$16176 ( \16553 , \16023 , \16520 );
or \U$16177 ( \16554 , \16552 , \16553 );
not \U$16178 ( \16555 , \16554 );
xor \U$16179 ( \16556 , \16523 , \16525 );
xor \U$16180 ( \16557 , \16556 , \16528 );
and \U$16181 ( \16558 , \16533 , \16557 );
xor \U$16182 ( \16559 , \16523 , \16525 );
xor \U$16183 ( \16560 , \16559 , \16528 );
and \U$16184 ( \16561 , \16549 , \16560 );
and \U$16185 ( \16562 , \16533 , \16549 );
or \U$16186 ( \16563 , \16558 , \16561 , \16562 );
xor \U$16187 ( \16564 , \15140 , \15150 );
xor \U$16188 ( \16565 , \16564 , \15157 );
xor \U$16189 ( \16566 , \16563 , \16565 );
xor \U$16190 ( \16567 , \16537 , \16539 );
and \U$16191 ( \16568 , \16567 , \16548 );
and \U$16192 ( \16569 , \16537 , \16539 );
or \U$16193 ( \16570 , \16568 , \16569 );
not \U$16194 ( \16571 , \14665 );
xnor \U$16195 ( \16572 , \14652 , \14325 );
not \U$16196 ( \16573 , \16572 );
or \U$16197 ( \16574 , \16571 , \16573 );
or \U$16198 ( \16575 , \16572 , \14665 );
nand \U$16199 ( \16576 , \16574 , \16575 );
xor \U$16200 ( \16577 , \16570 , \16576 );
xor \U$16201 ( \16578 , \16523 , \16525 );
and \U$16202 ( \16579 , \16578 , \16528 );
and \U$16203 ( \16580 , \16523 , \16525 );
or \U$16204 ( \16581 , \16579 , \16580 );
xor \U$16205 ( \16582 , \16577 , \16581 );
xor \U$16206 ( \16583 , \16566 , \16582 );
not \U$16207 ( \16584 , \16583 );
or \U$16208 ( \16585 , \16555 , \16584 );
xor \U$16209 ( \16586 , \16023 , \16520 );
xor \U$16210 ( \16587 , \16586 , \16551 );
xor \U$16211 ( \16588 , \15572 , \16022 );
not \U$16212 ( \16589 , \16588 );
xor \U$16213 ( \16590 , \16030 , \16040 );
xor \U$16214 ( \16591 , \16590 , \16517 );
not \U$16215 ( \16592 , \16591 );
or \U$16216 ( \16593 , \16589 , \16592 );
or \U$16217 ( \16594 , \16591 , \16588 );
xor \U$16218 ( \16595 , \16025 , \16029 );
xor \U$16219 ( \16596 , \15691 , \15760 );
xor \U$16220 ( \16597 , \16596 , \15842 );
xor \U$16221 ( \16598 , \15909 , \15967 );
xor \U$16222 ( \16599 , \16598 , \15980 );
and \U$16223 ( \16600 , \16597 , \16599 );
xor \U$16224 ( \16601 , \15590 , \15592 );
xor \U$16225 ( \16602 , \16601 , \15595 );
xor \U$16226 ( \16603 , \16482 , \16489 );
xor \U$16227 ( \16604 , \16602 , \16603 );
xor \U$16228 ( \16605 , \15909 , \15967 );
xor \U$16229 ( \16606 , \16605 , \15980 );
and \U$16230 ( \16607 , \16604 , \16606 );
and \U$16231 ( \16608 , \16597 , \16604 );
or \U$16232 ( \16609 , \16600 , \16607 , \16608 );
xor \U$16233 ( \16610 , \15845 , \15888 );
xor \U$16234 ( \16611 , \16610 , \15983 );
xor \U$16235 ( \16612 , \16609 , \16611 );
and \U$16236 ( \16613 , \3730 , RIae77e28_97);
and \U$16237 ( \16614 , RIae78968_121, \3728 );
nor \U$16238 ( \16615 , \16613 , \16614 );
and \U$16239 ( \16616 , \16615 , \3732 );
not \U$16240 ( \16617 , \16615 );
and \U$16241 ( \16618 , \16617 , \3422 );
nor \U$16242 ( \16619 , \16616 , \16618 );
not \U$16243 ( \16620 , \3089 );
and \U$16244 ( \16621 , \2783 , RIae78530_112);
and \U$16245 ( \16622 , RIae77c48_93, \2781 );
nor \U$16246 ( \16623 , \16621 , \16622 );
not \U$16247 ( \16624 , \16623 );
or \U$16248 ( \16625 , \16620 , \16624 );
or \U$16249 ( \16626 , \16623 , \3089 );
nand \U$16250 ( \16627 , \16625 , \16626 );
xor \U$16251 ( \16628 , \16619 , \16627 );
not \U$16252 ( \16629 , \2774 );
and \U$16253 ( \16630 , \3214 , RIae77b58_91);
and \U$16254 ( \16631 , RIae77d38_95, \3212 );
nor \U$16255 ( \16632 , \16630 , \16631 );
not \U$16256 ( \16633 , \16632 );
or \U$16257 ( \16634 , \16629 , \16633 );
or \U$16258 ( \16635 , \16632 , \3218 );
nand \U$16259 ( \16636 , \16634 , \16635 );
and \U$16260 ( \16637 , \16628 , \16636 );
and \U$16261 ( \16638 , \16619 , \16627 );
or \U$16262 ( \16639 , \16637 , \16638 );
and \U$16263 ( \16640 , \1939 , RIae780f8_103);
and \U$16264 ( \16641 , RIae77f18_99, \1937 );
nor \U$16265 ( \16642 , \16640 , \16641 );
and \U$16266 ( \16643 , \16642 , \1735 );
not \U$16267 ( \16644 , \16642 );
and \U$16268 ( \16645 , \16644 , \1734 );
nor \U$16269 ( \16646 , \16643 , \16645 );
and \U$16270 ( \16647 , \2224 , RIae78008_101);
and \U$16271 ( \16648 , RIae781e8_105, \2222 );
nor \U$16272 ( \16649 , \16647 , \16648 );
and \U$16273 ( \16650 , \16649 , \2061 );
not \U$16274 ( \16651 , \16649 );
and \U$16275 ( \16652 , \16651 , \2060 );
nor \U$16276 ( \16653 , \16650 , \16652 );
xor \U$16277 ( \16654 , \16646 , \16653 );
and \U$16278 ( \16655 , \2607 , RIae785a8_113);
and \U$16279 ( \16656 , RIae783c8_109, \2605 );
nor \U$16280 ( \16657 , \16655 , \16656 );
and \U$16281 ( \16658 , \16657 , \2611 );
not \U$16282 ( \16659 , \16657 );
and \U$16283 ( \16660 , \16659 , \2397 );
nor \U$16284 ( \16661 , \16658 , \16660 );
and \U$16285 ( \16662 , \16654 , \16661 );
and \U$16286 ( \16663 , \16646 , \16653 );
or \U$16287 ( \16664 , \16662 , \16663 );
xor \U$16288 ( \16665 , \16639 , \16664 );
and \U$16289 ( \16666 , \1593 , RIae772e8_73);
and \U$16290 ( \16667 , RIae782d8_107, \1591 );
nor \U$16291 ( \16668 , \16666 , \16667 );
and \U$16292 ( \16669 , \16668 , \1498 );
not \U$16293 ( \16670 , \16668 );
and \U$16294 ( \16671 , \16670 , \1488 );
nor \U$16295 ( \16672 , \16669 , \16671 );
and \U$16296 ( \16673 , \1138 , RIae76c58_59);
and \U$16297 ( \16674 , RIae77180_70, \1136 );
nor \U$16298 ( \16675 , \16673 , \16674 );
and \U$16299 ( \16676 , \16675 , \1012 );
not \U$16300 ( \16677 , \16675 );
and \U$16301 ( \16678 , \16677 , \1142 );
nor \U$16302 ( \16679 , \16676 , \16678 );
xor \U$16303 ( \16680 , \16672 , \16679 );
and \U$16304 ( \16681 , \1376 , RIae77018_67);
and \U$16305 ( \16682 , RIae771f8_71, \1374 );
nor \U$16306 ( \16683 , \16681 , \16682 );
and \U$16307 ( \16684 , \16683 , \1380 );
not \U$16308 ( \16685 , \16683 );
and \U$16309 ( \16686 , \16685 , \1261 );
nor \U$16310 ( \16687 , \16684 , \16686 );
and \U$16311 ( \16688 , \16680 , \16687 );
and \U$16312 ( \16689 , \16672 , \16679 );
or \U$16313 ( \16690 , \16688 , \16689 );
and \U$16314 ( \16691 , \16665 , \16690 );
and \U$16315 ( \16692 , \16639 , \16664 );
or \U$16316 ( \16693 , \16691 , \16692 );
and \U$16317 ( \16694 , \10548 , RIae764d8_43);
and \U$16318 ( \16695 , RIae766b8_47, \10546 );
nor \U$16319 ( \16696 , \16694 , \16695 );
and \U$16320 ( \16697 , \16696 , \10421 );
not \U$16321 ( \16698 , \16696 );
and \U$16322 ( \16699 , \16698 , \10118 );
nor \U$16323 ( \16700 , \16697 , \16699 );
and \U$16324 ( \16701 , \9760 , RIae753f8_7);
and \U$16325 ( \16702 , RIae763e8_41, \9758 );
nor \U$16326 ( \16703 , \16701 , \16702 );
and \U$16327 ( \16704 , \16703 , \9273 );
not \U$16328 ( \16705 , \16703 );
and \U$16329 ( \16706 , \16705 , \9272 );
nor \U$16330 ( \16707 , \16704 , \16706 );
xor \U$16331 ( \16708 , \16700 , \16707 );
and \U$16332 ( \16709 , \11470 , RIae765c8_45);
and \U$16333 ( \16710 , RIae76118_35, \11468 );
nor \U$16334 ( \16711 , \16709 , \16710 );
and \U$16335 ( \16712 , \16711 , \10936 );
not \U$16336 ( \16713 , \16711 );
and \U$16337 ( \16714 , \16713 , \11474 );
nor \U$16338 ( \16715 , \16712 , \16714 );
and \U$16339 ( \16716 , \16708 , \16715 );
and \U$16340 ( \16717 , \16700 , \16707 );
or \U$16341 ( \16718 , \16716 , \16717 );
and \U$16342 ( \16719 , \15726 , RIae78a58_123);
and \U$16343 ( \16720 , RIae7aab0_192, RIae78cb0_128);
nor \U$16344 ( \16721 , \16719 , \16720 );
and \U$16345 ( \16722 , \16721 , \14959 );
not \U$16346 ( \16723 , \16721 );
and \U$16347 ( \16724 , \16723 , RIae7aa38_191);
nor \U$16348 ( \16725 , \16722 , \16724 );
xor \U$16349 ( \16726 , \16725 , \388 );
and \U$16350 ( \16727 , \14964 , RIae76898_51);
and \U$16351 ( \16728 , RIae76b68_57, \14962 );
nor \U$16352 ( \16729 , \16727 , \16728 );
and \U$16353 ( \16730 , \16729 , \14463 );
not \U$16354 ( \16731 , \16729 );
and \U$16355 ( \16732 , \16731 , \14462 );
nor \U$16356 ( \16733 , \16730 , \16732 );
and \U$16357 ( \16734 , \16726 , \16733 );
and \U$16358 ( \16735 , \16725 , \388 );
or \U$16359 ( \16736 , \16734 , \16735 );
xor \U$16360 ( \16737 , \16718 , \16736 );
and \U$16361 ( \16738 , \12180 , RIae76028_33);
and \U$16362 ( \16739 , RIae762f8_39, \12178 );
nor \U$16363 ( \16740 , \16738 , \16739 );
and \U$16364 ( \16741 , \16740 , \12184 );
not \U$16365 ( \16742 , \16740 );
and \U$16366 ( \16743 , \16742 , \11827 );
nor \U$16367 ( \16744 , \16741 , \16743 );
and \U$16368 ( \16745 , \13059 , RIae76208_37);
and \U$16369 ( \16746 , RIae76a78_55, \13057 );
nor \U$16370 ( \16747 , \16745 , \16746 );
and \U$16371 ( \16748 , \16747 , \13063 );
not \U$16372 ( \16749 , \16747 );
and \U$16373 ( \16750 , \16749 , \12718 );
nor \U$16374 ( \16751 , \16748 , \16750 );
xor \U$16375 ( \16752 , \16744 , \16751 );
and \U$16376 ( \16753 , \14059 , RIae76988_53);
and \U$16377 ( \16754 , RIae767a8_49, \14057 );
nor \U$16378 ( \16755 , \16753 , \16754 );
and \U$16379 ( \16756 , \16755 , \13502 );
not \U$16380 ( \16757 , \16755 );
and \U$16381 ( \16758 , \16757 , \14063 );
nor \U$16382 ( \16759 , \16756 , \16758 );
and \U$16383 ( \16760 , \16752 , \16759 );
and \U$16384 ( \16761 , \16744 , \16751 );
or \U$16385 ( \16762 , \16760 , \16761 );
and \U$16386 ( \16763 , \16737 , \16762 );
and \U$16387 ( \16764 , \16718 , \16736 );
or \U$16388 ( \16765 , \16763 , \16764 );
xor \U$16389 ( \16766 , \16693 , \16765 );
and \U$16390 ( \16767 , \7633 , RIae754e8_9);
and \U$16391 ( \16768 , RIae757b8_15, \7631 );
nor \U$16392 ( \16769 , \16767 , \16768 );
and \U$16393 ( \16770 , \16769 , \7206 );
not \U$16394 ( \16771 , \16769 );
and \U$16395 ( \16772 , \16771 , \7205 );
nor \U$16396 ( \16773 , \16770 , \16772 );
and \U$16397 ( \16774 , \8371 , RIae756c8_13);
and \U$16398 ( \16775 , RIae75218_3, \8369 );
nor \U$16399 ( \16776 , \16774 , \16775 );
and \U$16400 ( \16777 , \16776 , \8020 );
not \U$16401 ( \16778 , \16776 );
and \U$16402 ( \16779 , \16778 , \8019 );
nor \U$16403 ( \16780 , \16777 , \16779 );
xor \U$16404 ( \16781 , \16773 , \16780 );
and \U$16405 ( \16782 , \8966 , RIae75128_1);
and \U$16406 ( \16783 , RIae75308_5, \8964 );
nor \U$16407 ( \16784 , \16782 , \16783 );
and \U$16408 ( \16785 , \16784 , \8799 );
not \U$16409 ( \16786 , \16784 );
and \U$16410 ( \16787 , \16786 , \8789 );
nor \U$16411 ( \16788 , \16785 , \16787 );
and \U$16412 ( \16789 , \16781 , \16788 );
and \U$16413 ( \16790 , \16773 , \16780 );
or \U$16414 ( \16791 , \16789 , \16790 );
and \U$16415 ( \16792 , \4247 , RIae78878_119);
and \U$16416 ( \16793 , RIae78788_117, \4245 );
nor \U$16417 ( \16794 , \16792 , \16793 );
and \U$16418 ( \16795 , \16794 , \3989 );
not \U$16419 ( \16796 , \16794 );
and \U$16420 ( \16797 , \16796 , \4251 );
nor \U$16421 ( \16798 , \16795 , \16797 );
and \U$16422 ( \16799 , \4688 , RIae78698_115);
and \U$16423 ( \16800 , RIae75b78_23, \4686 );
nor \U$16424 ( \16801 , \16799 , \16800 );
and \U$16425 ( \16802 , \16801 , \4481 );
not \U$16426 ( \16803 , \16801 );
and \U$16427 ( \16804 , \16803 , \4482 );
nor \U$16428 ( \16805 , \16802 , \16804 );
xor \U$16429 ( \16806 , \16798 , \16805 );
and \U$16430 ( \16807 , \5399 , RIae75a88_21);
and \U$16431 ( \16808 , RIae75998_19, \5397 );
nor \U$16432 ( \16809 , \16807 , \16808 );
and \U$16433 ( \16810 , \16809 , \5016 );
not \U$16434 ( \16811 , \16809 );
and \U$16435 ( \16812 , \16811 , \5403 );
nor \U$16436 ( \16813 , \16810 , \16812 );
and \U$16437 ( \16814 , \16806 , \16813 );
and \U$16438 ( \16815 , \16798 , \16805 );
or \U$16439 ( \16816 , \16814 , \16815 );
xor \U$16440 ( \16817 , \16791 , \16816 );
and \U$16441 ( \16818 , \6172 , RIae75e48_29);
and \U$16442 ( \16819 , RIae75c68_25, \6170 );
nor \U$16443 ( \16820 , \16818 , \16819 );
and \U$16444 ( \16821 , \16820 , \6176 );
not \U$16445 ( \16822 , \16820 );
and \U$16446 ( \16823 , \16822 , \6175 );
nor \U$16447 ( \16824 , \16821 , \16823 );
and \U$16448 ( \16825 , \5896 , RIae758a8_17);
and \U$16449 ( \16826 , RIae75f38_31, \5894 );
nor \U$16450 ( \16827 , \16825 , \16826 );
and \U$16451 ( \16828 , \16827 , \5590 );
not \U$16452 ( \16829 , \16827 );
and \U$16453 ( \16830 , \16829 , \5589 );
nor \U$16454 ( \16831 , \16828 , \16830 );
xor \U$16455 ( \16832 , \16824 , \16831 );
and \U$16456 ( \16833 , \6941 , RIae75d58_27);
and \U$16457 ( \16834 , RIae755d8_11, \6939 );
nor \U$16458 ( \16835 , \16833 , \16834 );
and \U$16459 ( \16836 , \16835 , \6314 );
not \U$16460 ( \16837 , \16835 );
and \U$16461 ( \16838 , \16837 , \6945 );
nor \U$16462 ( \16839 , \16836 , \16838 );
and \U$16463 ( \16840 , \16832 , \16839 );
and \U$16464 ( \16841 , \16824 , \16831 );
or \U$16465 ( \16842 , \16840 , \16841 );
and \U$16466 ( \16843 , \16817 , \16842 );
and \U$16467 ( \16844 , \16791 , \16816 );
or \U$16468 ( \16845 , \16843 , \16844 );
and \U$16469 ( \16846 , \16766 , \16845 );
and \U$16470 ( \16847 , \16693 , \16765 );
nor \U$16471 ( \16848 , \16846 , \16847 );
not \U$16472 ( \16849 , \16335 );
not \U$16473 ( \16850 , \16346 );
or \U$16474 ( \16851 , \16849 , \16850 );
or \U$16475 ( \16852 , \16346 , \16335 );
nand \U$16476 ( \16853 , \16851 , \16852 );
not \U$16477 ( \16854 , \16853 );
not \U$16478 ( \16855 , \16328 );
and \U$16479 ( \16856 , \16854 , \16855 );
and \U$16480 ( \16857 , \16853 , \16328 );
nor \U$16481 ( \16858 , \16856 , \16857 );
not \U$16482 ( \16859 , \16858 );
xor \U$16483 ( \16860 , \16277 , \16284 );
xor \U$16484 ( \16861 , \16860 , \16292 );
nand \U$16485 ( \16862 , \16859 , \16861 );
not \U$16486 ( \16863 , \15723 );
not \U$16487 ( \16864 , \15728 );
and \U$16488 ( \16865 , \16863 , \16864 );
and \U$16489 ( \16866 , \15723 , \15728 );
nor \U$16490 ( \16867 , \16865 , \16866 );
xor \U$16491 ( \16868 , \16862 , \16867 );
not \U$16492 ( \16869 , \16216 );
xor \U$16493 ( \16870 , \16224 , \16234 );
not \U$16494 ( \16871 , \16870 );
or \U$16495 ( \16872 , \16869 , \16871 );
or \U$16496 ( \16873 , \16870 , \16216 );
nand \U$16497 ( \16874 , \16872 , \16873 );
not \U$16498 ( \16875 , \16189 );
xor \U$16499 ( \16876 , \16197 , \16207 );
not \U$16500 ( \16877 , \16876 );
or \U$16501 ( \16878 , \16875 , \16877 );
or \U$16502 ( \16879 , \16876 , \16189 );
nand \U$16503 ( \16880 , \16878 , \16879 );
xor \U$16504 ( \16881 , \16874 , \16880 );
xor \U$16505 ( \16882 , \16302 , \16309 );
xor \U$16506 ( \16883 , \16882 , \16317 );
and \U$16507 ( \16884 , \16881 , \16883 );
and \U$16508 ( \16885 , \16874 , \16880 );
nor \U$16509 ( \16886 , \16884 , \16885 );
and \U$16510 ( \16887 , \16868 , \16886 );
and \U$16511 ( \16888 , \16862 , \16867 );
or \U$16512 ( \16889 , \16887 , \16888 );
xor \U$16513 ( \16890 , \16848 , \16889 );
not \U$16514 ( \16891 , \16381 );
xor \U$16515 ( \16892 , \16389 , \16399 );
not \U$16516 ( \16893 , \16892 );
or \U$16517 ( \16894 , \16891 , \16893 );
or \U$16518 ( \16895 , \16892 , \16381 );
nand \U$16519 ( \16896 , \16894 , \16895 );
not \U$16520 ( \16897 , \388 );
and \U$16521 ( \16898 , \384 , RIae775b8_79);
and \U$16522 ( \16899 , RIae774c8_77, \382 );
nor \U$16523 ( \16900 , \16898 , \16899 );
not \U$16524 ( \16901 , \16900 );
or \U$16525 ( \16902 , \16897 , \16901 );
or \U$16526 ( \16903 , \16900 , \388 );
nand \U$16527 ( \16904 , \16902 , \16903 );
xor \U$16528 ( \16905 , \16896 , \16904 );
xor \U$16529 ( \16906 , \16159 , \16167 );
xor \U$16530 ( \16907 , \16906 , \16175 );
and \U$16531 ( \16908 , \16905 , \16907 );
and \U$16532 ( \16909 , \16896 , \16904 );
or \U$16533 ( \16910 , \16908 , \16909 );
not \U$16534 ( \16911 , \402 );
and \U$16535 ( \16912 , \436 , RIae774c8_77);
and \U$16536 ( \16913 , RIae77720_82, \434 );
nor \U$16537 ( \16914 , \16912 , \16913 );
not \U$16538 ( \16915 , \16914 );
or \U$16539 ( \16916 , \16911 , \16915 );
or \U$16540 ( \16917 , \16914 , \402 );
nand \U$16541 ( \16918 , \16916 , \16917 );
nand \U$16542 ( \16919 , RIae775b8_79, \382 );
not \U$16543 ( \16920 , \16919 );
not \U$16544 ( \16921 , \388 );
or \U$16545 ( \16922 , \16920 , \16921 );
or \U$16546 ( \16923 , \388 , \16919 );
nand \U$16547 ( \16924 , \16922 , \16923 );
xor \U$16548 ( \16925 , \16918 , \16924 );
not \U$16549 ( \16926 , \471 );
and \U$16550 ( \16927 , \514 , RIae773d8_75);
and \U$16551 ( \16928 , RIae77a68_89, \512 );
nor \U$16552 ( \16929 , \16927 , \16928 );
not \U$16553 ( \16930 , \16929 );
or \U$16554 ( \16931 , \16926 , \16930 );
or \U$16555 ( \16932 , \16929 , \469 );
nand \U$16556 ( \16933 , \16931 , \16932 );
and \U$16557 ( \16934 , \16925 , \16933 );
and \U$16558 ( \16935 , \16918 , \16924 );
or \U$16559 ( \16936 , \16934 , \16935 );
not \U$16560 ( \16937 , \400 );
and \U$16561 ( \16938 , \436 , RIae77720_82);
and \U$16562 ( \16939 , RIae773d8_75, \434 );
nor \U$16563 ( \16940 , \16938 , \16939 );
not \U$16564 ( \16941 , \16940 );
or \U$16565 ( \16942 , \16937 , \16941 );
or \U$16566 ( \16943 , \16940 , \402 );
nand \U$16567 ( \16944 , \16942 , \16943 );
xor \U$16568 ( \16945 , \16936 , \16944 );
and \U$16569 ( \16946 , \558 , RIae77978_87);
and \U$16570 ( \16947 , RIae77798_83, \556 );
nor \U$16571 ( \16948 , \16946 , \16947 );
and \U$16572 ( \16949 , \16948 , \504 );
not \U$16573 ( \16950 , \16948 );
and \U$16574 ( \16951 , \16950 , \562 );
nor \U$16575 ( \16952 , \16949 , \16951 );
and \U$16576 ( \16953 , \672 , RIae77888_85);
and \U$16577 ( \16954 , RIae76f28_65, \670 );
nor \U$16578 ( \16955 , \16953 , \16954 );
and \U$16579 ( \16956 , \16955 , \588 );
not \U$16580 ( \16957 , \16955 );
and \U$16581 ( \16958 , \16957 , \587 );
nor \U$16582 ( \16959 , \16956 , \16958 );
xor \U$16583 ( \16960 , \16952 , \16959 );
not \U$16584 ( \16961 , \787 );
and \U$16585 ( \16962 , \883 , RIae76e38_63);
and \U$16586 ( \16963 , RIae76d48_61, \881 );
nor \U$16587 ( \16964 , \16962 , \16963 );
not \U$16588 ( \16965 , \16964 );
or \U$16589 ( \16966 , \16961 , \16965 );
or \U$16590 ( \16967 , \16964 , \787 );
nand \U$16591 ( \16968 , \16966 , \16967 );
and \U$16592 ( \16969 , \16960 , \16968 );
and \U$16593 ( \16970 , \16952 , \16959 );
or \U$16594 ( \16971 , \16969 , \16970 );
and \U$16595 ( \16972 , \16945 , \16971 );
and \U$16596 ( \16973 , \16936 , \16944 );
or \U$16597 ( \16974 , \16972 , \16973 );
xor \U$16598 ( \16975 , \16910 , \16974 );
xor \U$16599 ( \16976 , \16133 , \16140 );
xor \U$16600 ( \16977 , \16976 , \16148 );
xor \U$16601 ( \16978 , \16107 , \16114 );
xor \U$16602 ( \16979 , \16978 , \16123 );
xor \U$16603 ( \16980 , \16977 , \16979 );
not \U$16604 ( \16981 , \16244 );
xor \U$16605 ( \16982 , \16252 , \16262 );
not \U$16606 ( \16983 , \16982 );
or \U$16607 ( \16984 , \16981 , \16983 );
or \U$16608 ( \16985 , \16982 , \16244 );
nand \U$16609 ( \16986 , \16984 , \16985 );
and \U$16610 ( \16987 , \16980 , \16986 );
and \U$16611 ( \16988 , \16977 , \16979 );
or \U$16612 ( \16989 , \16987 , \16988 );
and \U$16613 ( \16990 , \16975 , \16989 );
and \U$16614 ( \16991 , \16910 , \16974 );
nor \U$16615 ( \16992 , \16990 , \16991 );
and \U$16616 ( \16993 , \16890 , \16992 );
and \U$16617 ( \16994 , \16848 , \16889 );
or \U$16618 ( \16995 , \16993 , \16994 );
not \U$16619 ( \16996 , \16059 );
xor \U$16620 ( \16997 , \16043 , \16045 );
not \U$16621 ( \16998 , \16997 );
or \U$16622 ( \16999 , \16996 , \16998 );
or \U$16623 ( \17000 , \16997 , \16059 );
nand \U$16624 ( \17001 , \16999 , \17000 );
xor \U$16625 ( \17002 , \16209 , \16236 );
xor \U$16626 ( \17003 , \17002 , \16264 );
xor \U$16627 ( \17004 , \16401 , \16402 );
xor \U$16628 ( \17005 , \17004 , \16413 );
or \U$16629 ( \17006 , \17003 , \17005 );
not \U$16630 ( \17007 , \17005 );
not \U$16631 ( \17008 , \17003 );
or \U$16632 ( \17009 , \17007 , \17008 );
xor \U$16633 ( \17010 , \16126 , \16151 );
xor \U$16634 ( \17011 , \17010 , \16178 );
nand \U$16635 ( \17012 , \17009 , \17011 );
nand \U$16636 ( \17013 , \17006 , \17012 );
xor \U$16637 ( \17014 , \17001 , \17013 );
xor \U$16638 ( \17015 , \16427 , \16429 );
xor \U$16639 ( \17016 , \17015 , \16432 );
xor \U$16640 ( \17017 , \16441 , \16451 );
xor \U$16641 ( \17018 , \17017 , \16454 );
or \U$16642 ( \17019 , \17016 , \17018 );
not \U$16643 ( \17020 , \17018 );
not \U$16644 ( \17021 , \17016 );
or \U$16645 ( \17022 , \17020 , \17021 );
not \U$16646 ( \17023 , \16363 );
xor \U$16647 ( \17024 , \16371 , \16366 );
not \U$16648 ( \17025 , \17024 );
or \U$16649 ( \17026 , \17023 , \17025 );
or \U$16650 ( \17027 , \17024 , \16363 );
nand \U$16651 ( \17028 , \17026 , \17027 );
nand \U$16652 ( \17029 , \17022 , \17028 );
nand \U$16653 ( \17030 , \17019 , \17029 );
and \U$16654 ( \17031 , \17014 , \17030 );
and \U$16655 ( \17032 , \17001 , \17013 );
nor \U$16656 ( \17033 , \17031 , \17032 );
xor \U$16657 ( \17034 , \16995 , \17033 );
xor \U$16658 ( \17035 , \16457 , \16462 );
xor \U$16659 ( \17036 , \17035 , \16473 );
not \U$16660 ( \17037 , \17036 );
xor \U$16661 ( \17038 , \16373 , \16416 );
xor \U$16662 ( \17039 , \17038 , \16435 );
not \U$16663 ( \17040 , \17039 );
and \U$16664 ( \17041 , \17037 , \17040 );
and \U$16665 ( \17042 , \17036 , \17039 );
not \U$16666 ( \17043 , \16095 );
not \U$16667 ( \17044 , \16085 );
or \U$16668 ( \17045 , \17043 , \17044 );
or \U$16669 ( \17046 , \16085 , \16095 );
nand \U$16670 ( \17047 , \17045 , \17046 );
not \U$16671 ( \17048 , \17047 );
not \U$16672 ( \17049 , \16087 );
and \U$16673 ( \17050 , \17048 , \17049 );
and \U$16674 ( \17051 , \17047 , \16087 );
nor \U$16675 ( \17052 , \17050 , \17051 );
nor \U$16676 ( \17053 , \17042 , \17052 );
nor \U$16677 ( \17054 , \17041 , \17053 );
and \U$16678 ( \17055 , \17034 , \17054 );
and \U$16679 ( \17056 , \16995 , \17033 );
nor \U$16680 ( \17057 , \17055 , \17056 );
and \U$16681 ( \17058 , \16612 , \17057 );
and \U$16682 ( \17059 , \16609 , \16611 );
or \U$16683 ( \17060 , \17058 , \17059 );
xor \U$16684 ( \17061 , \16595 , \17060 );
xor \U$16685 ( \17062 , \16497 , \16499 );
xor \U$16686 ( \17063 , \17062 , \16514 );
and \U$16687 ( \17064 , \17061 , \17063 );
and \U$16688 ( \17065 , \16595 , \17060 );
or \U$16689 ( \17066 , \17064 , \17065 );
nand \U$16690 ( \17067 , \16594 , \17066 );
nand \U$16691 ( \17068 , \16593 , \17067 );
and \U$16692 ( \17069 , \16587 , \17068 );
xor \U$16693 ( \17070 , \17068 , \16587 );
xor \U$16694 ( \17071 , \16910 , \16974 );
xor \U$16695 ( \17072 , \17071 , \16989 );
xor \U$16696 ( \17073 , \16693 , \16765 );
xor \U$16697 ( \17074 , \17073 , \16845 );
and \U$16698 ( \17075 , \17072 , \17074 );
not \U$16699 ( \17076 , \17072 );
not \U$16700 ( \17077 , \17074 );
and \U$16701 ( \17078 , \17076 , \17077 );
not \U$16702 ( \17079 , \17003 );
not \U$16703 ( \17080 , \17011 );
or \U$16704 ( \17081 , \17079 , \17080 );
or \U$16705 ( \17082 , \17003 , \17011 );
nand \U$16706 ( \17083 , \17081 , \17082 );
not \U$16707 ( \17084 , \17083 );
not \U$16708 ( \17085 , \17005 );
and \U$16709 ( \17086 , \17084 , \17085 );
and \U$16710 ( \17087 , \17083 , \17005 );
nor \U$16711 ( \17088 , \17086 , \17087 );
xor \U$16712 ( \17089 , \16862 , \16867 );
xor \U$16713 ( \17090 , \17089 , \16886 );
xor \U$16714 ( \17091 , \17088 , \17090 );
not \U$16715 ( \17092 , \17018 );
not \U$16716 ( \17093 , \17028 );
or \U$16717 ( \17094 , \17092 , \17093 );
or \U$16718 ( \17095 , \17018 , \17028 );
nand \U$16719 ( \17096 , \17094 , \17095 );
not \U$16720 ( \17097 , \17096 );
not \U$16721 ( \17098 , \17016 );
and \U$16722 ( \17099 , \17097 , \17098 );
and \U$16723 ( \17100 , \17096 , \17016 );
nor \U$16724 ( \17101 , \17099 , \17100 );
xor \U$16725 ( \17102 , \17091 , \17101 );
nor \U$16726 ( \17103 , \17078 , \17102 );
nor \U$16727 ( \17104 , \17075 , \17103 );
xor \U$16728 ( \17105 , \16848 , \16889 );
xor \U$16729 ( \17106 , \17105 , \16992 );
xor \U$16730 ( \17107 , \17104 , \17106 );
xor \U$16731 ( \17108 , \16798 , \16805 );
xor \U$16732 ( \17109 , \17108 , \16813 );
xor \U$16733 ( \17110 , \16824 , \16831 );
xor \U$16734 ( \17111 , \17110 , \16839 );
and \U$16735 ( \17112 , \17109 , \17111 );
xor \U$16736 ( \17113 , \16773 , \16780 );
xor \U$16737 ( \17114 , \17113 , \16788 );
xor \U$16738 ( \17115 , \16824 , \16831 );
xor \U$16739 ( \17116 , \17115 , \16839 );
and \U$16740 ( \17117 , \17114 , \17116 );
and \U$16741 ( \17118 , \17109 , \17114 );
or \U$16742 ( \17119 , \17112 , \17117 , \17118 );
not \U$16743 ( \17120 , \469 );
and \U$16744 ( \17121 , \514 , RIae77720_82);
and \U$16745 ( \17122 , RIae773d8_75, \512 );
nor \U$16746 ( \17123 , \17121 , \17122 );
not \U$16747 ( \17124 , \17123 );
or \U$16748 ( \17125 , \17120 , \17124 );
or \U$16749 ( \17126 , \17123 , \469 );
nand \U$16750 ( \17127 , \17125 , \17126 );
and \U$16751 ( \17128 , \558 , RIae77a68_89);
and \U$16752 ( \17129 , RIae77978_87, \556 );
nor \U$16753 ( \17130 , \17128 , \17129 );
and \U$16754 ( \17131 , \17130 , \504 );
not \U$16755 ( \17132 , \17130 );
and \U$16756 ( \17133 , \17132 , \562 );
nor \U$16757 ( \17134 , \17131 , \17133 );
xor \U$16758 ( \17135 , \17127 , \17134 );
and \U$16759 ( \17136 , \672 , RIae77798_83);
and \U$16760 ( \17137 , RIae77888_85, \670 );
nor \U$16761 ( \17138 , \17136 , \17137 );
and \U$16762 ( \17139 , \17138 , \588 );
not \U$16763 ( \17140 , \17138 );
and \U$16764 ( \17141 , \17140 , \587 );
nor \U$16765 ( \17142 , \17139 , \17141 );
and \U$16766 ( \17143 , \17135 , \17142 );
and \U$16767 ( \17144 , \17127 , \17134 );
or \U$16768 ( \17145 , \17143 , \17144 );
xor \U$16769 ( \17146 , \16918 , \16924 );
xor \U$16770 ( \17147 , \17146 , \16933 );
and \U$16771 ( \17148 , \17145 , \17147 );
xor \U$16772 ( \17149 , \16952 , \16959 );
xor \U$16773 ( \17150 , \17149 , \16968 );
xor \U$16774 ( \17151 , \16918 , \16924 );
xor \U$16775 ( \17152 , \17151 , \16933 );
and \U$16776 ( \17153 , \17150 , \17152 );
and \U$16777 ( \17154 , \17145 , \17150 );
or \U$16778 ( \17155 , \17148 , \17153 , \17154 );
xor \U$16779 ( \17156 , \17119 , \17155 );
xor \U$16780 ( \17157 , \16672 , \16679 );
xor \U$16781 ( \17158 , \17157 , \16687 );
xor \U$16782 ( \17159 , \16646 , \16653 );
xor \U$16783 ( \17160 , \17159 , \16661 );
and \U$16784 ( \17161 , \17158 , \17160 );
xor \U$16785 ( \17162 , \16619 , \16627 );
xor \U$16786 ( \17163 , \17162 , \16636 );
xor \U$16787 ( \17164 , \16646 , \16653 );
xor \U$16788 ( \17165 , \17164 , \16661 );
and \U$16789 ( \17166 , \17163 , \17165 );
and \U$16790 ( \17167 , \17158 , \17163 );
or \U$16791 ( \17168 , \17161 , \17166 , \17167 );
xor \U$16792 ( \17169 , \17156 , \17168 );
and \U$16793 ( \17170 , \7633 , RIae755d8_11);
and \U$16794 ( \17171 , RIae754e8_9, \7631 );
nor \U$16795 ( \17172 , \17170 , \17171 );
and \U$16796 ( \17173 , \17172 , \7206 );
not \U$16797 ( \17174 , \17172 );
and \U$16798 ( \17175 , \17174 , \7205 );
nor \U$16799 ( \17176 , \17173 , \17175 );
and \U$16800 ( \17177 , \6941 , RIae75c68_25);
and \U$16801 ( \17178 , RIae75d58_27, \6939 );
nor \U$16802 ( \17179 , \17177 , \17178 );
and \U$16803 ( \17180 , \17179 , \6314 );
not \U$16804 ( \17181 , \17179 );
and \U$16805 ( \17182 , \17181 , \6945 );
nor \U$16806 ( \17183 , \17180 , \17182 );
xor \U$16807 ( \17184 , \17176 , \17183 );
and \U$16808 ( \17185 , \8371 , RIae757b8_15);
and \U$16809 ( \17186 , RIae756c8_13, \8369 );
nor \U$16810 ( \17187 , \17185 , \17186 );
and \U$16811 ( \17188 , \17187 , \8020 );
not \U$16812 ( \17189 , \17187 );
and \U$16813 ( \17190 , \17189 , \8019 );
nor \U$16814 ( \17191 , \17188 , \17190 );
and \U$16815 ( \17192 , \17184 , \17191 );
and \U$16816 ( \17193 , \17176 , \17183 );
or \U$16817 ( \17194 , \17192 , \17193 );
and \U$16818 ( \17195 , \5399 , RIae75b78_23);
and \U$16819 ( \17196 , RIae75a88_21, \5397 );
nor \U$16820 ( \17197 , \17195 , \17196 );
and \U$16821 ( \17198 , \17197 , \5016 );
not \U$16822 ( \17199 , \17197 );
and \U$16823 ( \17200 , \17199 , \5403 );
nor \U$16824 ( \17201 , \17198 , \17200 );
and \U$16825 ( \17202 , \5896 , RIae75998_19);
and \U$16826 ( \17203 , RIae758a8_17, \5894 );
nor \U$16827 ( \17204 , \17202 , \17203 );
and \U$16828 ( \17205 , \17204 , \5590 );
not \U$16829 ( \17206 , \17204 );
and \U$16830 ( \17207 , \17206 , \5589 );
nor \U$16831 ( \17208 , \17205 , \17207 );
xor \U$16832 ( \17209 , \17201 , \17208 );
and \U$16833 ( \17210 , \6172 , RIae75f38_31);
and \U$16834 ( \17211 , RIae75e48_29, \6170 );
nor \U$16835 ( \17212 , \17210 , \17211 );
and \U$16836 ( \17213 , \17212 , \6176 );
not \U$16837 ( \17214 , \17212 );
and \U$16838 ( \17215 , \17214 , \6175 );
nor \U$16839 ( \17216 , \17213 , \17215 );
and \U$16840 ( \17217 , \17209 , \17216 );
and \U$16841 ( \17218 , \17201 , \17208 );
or \U$16842 ( \17219 , \17217 , \17218 );
xor \U$16843 ( \17220 , \17194 , \17219 );
and \U$16844 ( \17221 , \3730 , RIae77d38_95);
and \U$16845 ( \17222 , RIae77e28_97, \3728 );
nor \U$16846 ( \17223 , \17221 , \17222 );
and \U$16847 ( \17224 , \17223 , \3732 );
not \U$16848 ( \17225 , \17223 );
and \U$16849 ( \17226 , \17225 , \3422 );
nor \U$16850 ( \17227 , \17224 , \17226 );
and \U$16851 ( \17228 , \4247 , RIae78968_121);
and \U$16852 ( \17229 , RIae78878_119, \4245 );
nor \U$16853 ( \17230 , \17228 , \17229 );
and \U$16854 ( \17231 , \17230 , \3989 );
not \U$16855 ( \17232 , \17230 );
and \U$16856 ( \17233 , \17232 , \4251 );
nor \U$16857 ( \17234 , \17231 , \17233 );
xor \U$16858 ( \17235 , \17227 , \17234 );
and \U$16859 ( \17236 , \4688 , RIae78788_117);
and \U$16860 ( \17237 , RIae78698_115, \4686 );
nor \U$16861 ( \17238 , \17236 , \17237 );
and \U$16862 ( \17239 , \17238 , \4481 );
not \U$16863 ( \17240 , \17238 );
and \U$16864 ( \17241 , \17240 , \4482 );
nor \U$16865 ( \17242 , \17239 , \17241 );
and \U$16866 ( \17243 , \17235 , \17242 );
and \U$16867 ( \17244 , \17227 , \17234 );
or \U$16868 ( \17245 , \17243 , \17244 );
and \U$16869 ( \17246 , \17220 , \17245 );
and \U$16870 ( \17247 , \17194 , \17219 );
or \U$16871 ( \17248 , \17246 , \17247 );
and \U$16872 ( \17249 , \11470 , RIae766b8_47);
and \U$16873 ( \17250 , RIae765c8_45, \11468 );
nor \U$16874 ( \17251 , \17249 , \17250 );
and \U$16875 ( \17252 , \17251 , \10936 );
not \U$16876 ( \17253 , \17251 );
and \U$16877 ( \17254 , \17253 , \11474 );
nor \U$16878 ( \17255 , \17252 , \17254 );
and \U$16879 ( \17256 , \12180 , RIae76118_35);
and \U$16880 ( \17257 , RIae76028_33, \12178 );
nor \U$16881 ( \17258 , \17256 , \17257 );
and \U$16882 ( \17259 , \17258 , \12184 );
not \U$16883 ( \17260 , \17258 );
and \U$16884 ( \17261 , \17260 , \11827 );
nor \U$16885 ( \17262 , \17259 , \17261 );
xor \U$16886 ( \17263 , \17255 , \17262 );
and \U$16887 ( \17264 , \13059 , RIae762f8_39);
and \U$16888 ( \17265 , RIae76208_37, \13057 );
nor \U$16889 ( \17266 , \17264 , \17265 );
and \U$16890 ( \17267 , \17266 , \13063 );
not \U$16891 ( \17268 , \17266 );
and \U$16892 ( \17269 , \17268 , \12718 );
nor \U$16893 ( \17270 , \17267 , \17269 );
and \U$16894 ( \17271 , \17263 , \17270 );
and \U$16895 ( \17272 , \17255 , \17262 );
or \U$16896 ( \17273 , \17271 , \17272 );
and \U$16897 ( \17274 , \14964 , RIae767a8_49);
and \U$16898 ( \17275 , RIae76898_51, \14962 );
nor \U$16899 ( \17276 , \17274 , \17275 );
and \U$16900 ( \17277 , \17276 , \14463 );
not \U$16901 ( \17278 , \17276 );
and \U$16902 ( \17279 , \17278 , \14462 );
nor \U$16903 ( \17280 , \17277 , \17279 );
and \U$16904 ( \17281 , \15726 , RIae76b68_57);
and \U$16905 ( \17282 , RIae7aab0_192, RIae78a58_123);
nor \U$16906 ( \17283 , \17281 , \17282 );
and \U$16907 ( \17284 , \17283 , \14959 );
not \U$16908 ( \17285 , \17283 );
and \U$16909 ( \17286 , \17285 , RIae7aa38_191);
nor \U$16910 ( \17287 , \17284 , \17286 );
xor \U$16911 ( \17288 , \17280 , \17287 );
and \U$16912 ( \17289 , \14059 , RIae76a78_55);
and \U$16913 ( \17290 , RIae76988_53, \14057 );
nor \U$16914 ( \17291 , \17289 , \17290 );
and \U$16915 ( \17292 , \17291 , \13502 );
not \U$16916 ( \17293 , \17291 );
and \U$16917 ( \17294 , \17293 , \14063 );
nor \U$16918 ( \17295 , \17292 , \17294 );
and \U$16919 ( \17296 , \17288 , \17295 );
and \U$16920 ( \17297 , \17280 , \17287 );
or \U$16921 ( \17298 , \17296 , \17297 );
xor \U$16922 ( \17299 , \17273 , \17298 );
and \U$16923 ( \17300 , \10548 , RIae763e8_41);
and \U$16924 ( \17301 , RIae764d8_43, \10546 );
nor \U$16925 ( \17302 , \17300 , \17301 );
and \U$16926 ( \17303 , \17302 , \10421 );
not \U$16927 ( \17304 , \17302 );
and \U$16928 ( \17305 , \17304 , \10118 );
nor \U$16929 ( \17306 , \17303 , \17305 );
and \U$16930 ( \17307 , \8966 , RIae75218_3);
and \U$16931 ( \17308 , RIae75128_1, \8964 );
nor \U$16932 ( \17309 , \17307 , \17308 );
and \U$16933 ( \17310 , \17309 , \8799 );
not \U$16934 ( \17311 , \17309 );
and \U$16935 ( \17312 , \17311 , \8789 );
nor \U$16936 ( \17313 , \17310 , \17312 );
xor \U$16937 ( \17314 , \17306 , \17313 );
and \U$16938 ( \17315 , \9760 , RIae75308_5);
and \U$16939 ( \17316 , RIae753f8_7, \9758 );
nor \U$16940 ( \17317 , \17315 , \17316 );
and \U$16941 ( \17318 , \17317 , \9273 );
not \U$16942 ( \17319 , \17317 );
and \U$16943 ( \17320 , \17319 , \9764 );
nor \U$16944 ( \17321 , \17318 , \17320 );
and \U$16945 ( \17322 , \17314 , \17321 );
and \U$16946 ( \17323 , \17306 , \17313 );
or \U$16947 ( \17324 , \17322 , \17323 );
and \U$16948 ( \17325 , \17299 , \17324 );
and \U$16949 ( \17326 , \17273 , \17298 );
or \U$16950 ( \17327 , \17325 , \17326 );
xor \U$16951 ( \17328 , \17248 , \17327 );
and \U$16952 ( \17329 , \1593 , RIae771f8_71);
and \U$16953 ( \17330 , RIae772e8_73, \1591 );
nor \U$16954 ( \17331 , \17329 , \17330 );
and \U$16955 ( \17332 , \17331 , \1498 );
not \U$16956 ( \17333 , \17331 );
and \U$16957 ( \17334 , \17333 , \1488 );
nor \U$16958 ( \17335 , \17332 , \17334 );
and \U$16959 ( \17336 , \1939 , RIae782d8_107);
and \U$16960 ( \17337 , RIae780f8_103, \1937 );
nor \U$16961 ( \17338 , \17336 , \17337 );
and \U$16962 ( \17339 , \17338 , \1735 );
not \U$16963 ( \17340 , \17338 );
and \U$16964 ( \17341 , \17340 , \1734 );
nor \U$16965 ( \17342 , \17339 , \17341 );
xor \U$16966 ( \17343 , \17335 , \17342 );
and \U$16967 ( \17344 , \2224 , RIae77f18_99);
and \U$16968 ( \17345 , RIae78008_101, \2222 );
nor \U$16969 ( \17346 , \17344 , \17345 );
and \U$16970 ( \17347 , \17346 , \2061 );
not \U$16971 ( \17348 , \17346 );
and \U$16972 ( \17349 , \17348 , \2060 );
nor \U$16973 ( \17350 , \17347 , \17349 );
and \U$16974 ( \17351 , \17343 , \17350 );
and \U$16975 ( \17352 , \17335 , \17342 );
or \U$16976 ( \17353 , \17351 , \17352 );
and \U$16977 ( \17354 , \1376 , RIae77180_70);
and \U$16978 ( \17355 , RIae77018_67, \1374 );
nor \U$16979 ( \17356 , \17354 , \17355 );
and \U$16980 ( \17357 , \17356 , \1380 );
not \U$16981 ( \17358 , \17356 );
and \U$16982 ( \17359 , \17358 , \1261 );
nor \U$16983 ( \17360 , \17357 , \17359 );
not \U$16984 ( \17361 , \789 );
and \U$16985 ( \17362 , \883 , RIae76f28_65);
and \U$16986 ( \17363 , RIae76e38_63, \881 );
nor \U$16987 ( \17364 , \17362 , \17363 );
not \U$16988 ( \17365 , \17364 );
or \U$16989 ( \17366 , \17361 , \17365 );
or \U$16990 ( \17367 , \17364 , \787 );
nand \U$16991 ( \17368 , \17366 , \17367 );
xor \U$16992 ( \17369 , \17360 , \17368 );
and \U$16993 ( \17370 , \1138 , RIae76d48_61);
and \U$16994 ( \17371 , RIae76c58_59, \1136 );
nor \U$16995 ( \17372 , \17370 , \17371 );
and \U$16996 ( \17373 , \17372 , \1012 );
not \U$16997 ( \17374 , \17372 );
and \U$16998 ( \17375 , \17374 , \1142 );
nor \U$16999 ( \17376 , \17373 , \17375 );
and \U$17000 ( \17377 , \17369 , \17376 );
and \U$17001 ( \17378 , \17360 , \17368 );
or \U$17002 ( \17379 , \17377 , \17378 );
xor \U$17003 ( \17380 , \17353 , \17379 );
not \U$17004 ( \17381 , \3218 );
and \U$17005 ( \17382 , \3214 , RIae77c48_93);
and \U$17006 ( \17383 , RIae77b58_91, \3212 );
nor \U$17007 ( \17384 , \17382 , \17383 );
not \U$17008 ( \17385 , \17384 );
or \U$17009 ( \17386 , \17381 , \17385 );
or \U$17010 ( \17387 , \17384 , \3218 );
nand \U$17011 ( \17388 , \17386 , \17387 );
and \U$17012 ( \17389 , \2607 , RIae781e8_105);
and \U$17013 ( \17390 , RIae785a8_113, \2605 );
nor \U$17014 ( \17391 , \17389 , \17390 );
and \U$17015 ( \17392 , \17391 , \2611 );
not \U$17016 ( \17393 , \17391 );
and \U$17017 ( \17394 , \17393 , \2397 );
nor \U$17018 ( \17395 , \17392 , \17394 );
xor \U$17019 ( \17396 , \17388 , \17395 );
not \U$17020 ( \17397 , \3089 );
and \U$17021 ( \17398 , \2783 , RIae783c8_109);
and \U$17022 ( \17399 , RIae78530_112, \2781 );
nor \U$17023 ( \17400 , \17398 , \17399 );
not \U$17024 ( \17401 , \17400 );
or \U$17025 ( \17402 , \17397 , \17401 );
or \U$17026 ( \17403 , \17400 , \3089 );
nand \U$17027 ( \17404 , \17402 , \17403 );
and \U$17028 ( \17405 , \17396 , \17404 );
and \U$17029 ( \17406 , \17388 , \17395 );
or \U$17030 ( \17407 , \17405 , \17406 );
and \U$17031 ( \17408 , \17380 , \17407 );
and \U$17032 ( \17409 , \17353 , \17379 );
or \U$17033 ( \17410 , \17408 , \17409 );
xor \U$17034 ( \17411 , \17328 , \17410 );
xor \U$17035 ( \17412 , \17169 , \17411 );
xor \U$17036 ( \17413 , \16725 , \388 );
xor \U$17037 ( \17414 , \17413 , \16733 );
xor \U$17038 ( \17415 , \16700 , \16707 );
xor \U$17039 ( \17416 , \17415 , \16715 );
xor \U$17040 ( \17417 , \17414 , \17416 );
xor \U$17041 ( \17418 , \16744 , \16751 );
xor \U$17042 ( \17419 , \17418 , \16759 );
and \U$17043 ( \17420 , \17417 , \17419 );
and \U$17044 ( \17421 , \17414 , \17416 );
or \U$17045 ( \17422 , \17420 , \17421 );
not \U$17046 ( \17423 , \16861 );
not \U$17047 ( \17424 , \16858 );
or \U$17048 ( \17425 , \17423 , \17424 );
or \U$17049 ( \17426 , \16858 , \16861 );
nand \U$17050 ( \17427 , \17425 , \17426 );
xor \U$17051 ( \17428 , \17422 , \17427 );
xor \U$17052 ( \17429 , \16874 , \16880 );
xor \U$17053 ( \17430 , \17429 , \16883 );
xor \U$17054 ( \17431 , \17428 , \17430 );
and \U$17055 ( \17432 , \17412 , \17431 );
and \U$17056 ( \17433 , \17169 , \17411 );
or \U$17057 ( \17434 , \17432 , \17433 );
xor \U$17058 ( \17435 , \17388 , \17395 );
xor \U$17059 ( \17436 , \17435 , \17404 );
xor \U$17060 ( \17437 , \17201 , \17208 );
xor \U$17061 ( \17438 , \17437 , \17216 );
and \U$17062 ( \17439 , \17436 , \17438 );
xor \U$17063 ( \17440 , \17227 , \17234 );
xor \U$17064 ( \17441 , \17440 , \17242 );
xor \U$17065 ( \17442 , \17201 , \17208 );
xor \U$17066 ( \17443 , \17442 , \17216 );
and \U$17067 ( \17444 , \17441 , \17443 );
and \U$17068 ( \17445 , \17436 , \17441 );
or \U$17069 ( \17446 , \17439 , \17444 , \17445 );
nand \U$17070 ( \17447 , RIae775b8_79, \434 );
not \U$17071 ( \17448 , \17447 );
not \U$17072 ( \17449 , \400 );
or \U$17073 ( \17450 , \17448 , \17449 );
or \U$17074 ( \17451 , \400 , \17447 );
nand \U$17075 ( \17452 , \17450 , \17451 );
not \U$17076 ( \17453 , \471 );
and \U$17077 ( \17454 , \514 , RIae774c8_77);
and \U$17078 ( \17455 , RIae77720_82, \512 );
nor \U$17079 ( \17456 , \17454 , \17455 );
not \U$17080 ( \17457 , \17456 );
or \U$17081 ( \17458 , \17453 , \17457 );
or \U$17082 ( \17459 , \17456 , \471 );
nand \U$17083 ( \17460 , \17458 , \17459 );
and \U$17084 ( \17461 , \17452 , \17460 );
not \U$17085 ( \17462 , \402 );
and \U$17086 ( \17463 , \436 , RIae775b8_79);
and \U$17087 ( \17464 , RIae774c8_77, \434 );
nor \U$17088 ( \17465 , \17463 , \17464 );
not \U$17089 ( \17466 , \17465 );
or \U$17090 ( \17467 , \17462 , \17466 );
or \U$17091 ( \17468 , \17465 , \402 );
nand \U$17092 ( \17469 , \17467 , \17468 );
xor \U$17093 ( \17470 , \17461 , \17469 );
not \U$17094 ( \17471 , \789 );
and \U$17095 ( \17472 , \883 , RIae77888_85);
and \U$17096 ( \17473 , RIae76f28_65, \881 );
nor \U$17097 ( \17474 , \17472 , \17473 );
not \U$17098 ( \17475 , \17474 );
or \U$17099 ( \17476 , \17471 , \17475 );
or \U$17100 ( \17477 , \17474 , \789 );
nand \U$17101 ( \17478 , \17476 , \17477 );
and \U$17102 ( \17479 , \558 , RIae773d8_75);
and \U$17103 ( \17480 , RIae77a68_89, \556 );
nor \U$17104 ( \17481 , \17479 , \17480 );
and \U$17105 ( \17482 , \17481 , \504 );
not \U$17106 ( \17483 , \17481 );
and \U$17107 ( \17484 , \17483 , \562 );
nor \U$17108 ( \17485 , \17482 , \17484 );
xor \U$17109 ( \17486 , \17478 , \17485 );
and \U$17110 ( \17487 , \672 , RIae77978_87);
and \U$17111 ( \17488 , RIae77798_83, \670 );
nor \U$17112 ( \17489 , \17487 , \17488 );
and \U$17113 ( \17490 , \17489 , \588 );
not \U$17114 ( \17491 , \17489 );
and \U$17115 ( \17492 , \17491 , \587 );
nor \U$17116 ( \17493 , \17490 , \17492 );
and \U$17117 ( \17494 , \17486 , \17493 );
and \U$17118 ( \17495 , \17478 , \17485 );
or \U$17119 ( \17496 , \17494 , \17495 );
and \U$17120 ( \17497 , \17470 , \17496 );
and \U$17121 ( \17498 , \17461 , \17469 );
or \U$17122 ( \17499 , \17497 , \17498 );
xor \U$17123 ( \17500 , \17446 , \17499 );
xor \U$17124 ( \17501 , \17127 , \17134 );
xor \U$17125 ( \17502 , \17501 , \17142 );
xor \U$17126 ( \17503 , \17360 , \17368 );
xor \U$17127 ( \17504 , \17503 , \17376 );
xor \U$17128 ( \17505 , \17502 , \17504 );
xor \U$17129 ( \17506 , \17335 , \17342 );
xor \U$17130 ( \17507 , \17506 , \17350 );
and \U$17131 ( \17508 , \17505 , \17507 );
and \U$17132 ( \17509 , \17502 , \17504 );
or \U$17133 ( \17510 , \17508 , \17509 );
and \U$17134 ( \17511 , \17500 , \17510 );
and \U$17135 ( \17512 , \17446 , \17499 );
or \U$17136 ( \17513 , \17511 , \17512 );
and \U$17137 ( \17514 , \3730 , RIae77b58_91);
and \U$17138 ( \17515 , RIae77d38_95, \3728 );
nor \U$17139 ( \17516 , \17514 , \17515 );
and \U$17140 ( \17517 , \17516 , \3732 );
not \U$17141 ( \17518 , \17516 );
and \U$17142 ( \17519 , \17518 , \3422 );
nor \U$17143 ( \17520 , \17517 , \17519 );
not \U$17144 ( \17521 , \3089 );
and \U$17145 ( \17522 , \2783 , RIae785a8_113);
and \U$17146 ( \17523 , RIae783c8_109, \2781 );
nor \U$17147 ( \17524 , \17522 , \17523 );
not \U$17148 ( \17525 , \17524 );
or \U$17149 ( \17526 , \17521 , \17525 );
or \U$17150 ( \17527 , \17524 , \3089 );
nand \U$17151 ( \17528 , \17526 , \17527 );
xor \U$17152 ( \17529 , \17520 , \17528 );
not \U$17153 ( \17530 , \2774 );
and \U$17154 ( \17531 , \3214 , RIae78530_112);
and \U$17155 ( \17532 , RIae77c48_93, \3212 );
nor \U$17156 ( \17533 , \17531 , \17532 );
not \U$17157 ( \17534 , \17533 );
or \U$17158 ( \17535 , \17530 , \17534 );
or \U$17159 ( \17536 , \17533 , \2774 );
nand \U$17160 ( \17537 , \17535 , \17536 );
and \U$17161 ( \17538 , \17529 , \17537 );
and \U$17162 ( \17539 , \17520 , \17528 );
or \U$17163 ( \17540 , \17538 , \17539 );
and \U$17164 ( \17541 , \1593 , RIae77018_67);
and \U$17165 ( \17542 , RIae771f8_71, \1591 );
nor \U$17166 ( \17543 , \17541 , \17542 );
and \U$17167 ( \17544 , \17543 , \1498 );
not \U$17168 ( \17545 , \17543 );
and \U$17169 ( \17546 , \17545 , \1488 );
nor \U$17170 ( \17547 , \17544 , \17546 );
and \U$17171 ( \17548 , \1138 , RIae76e38_63);
and \U$17172 ( \17549 , RIae76d48_61, \1136 );
nor \U$17173 ( \17550 , \17548 , \17549 );
and \U$17174 ( \17551 , \17550 , \1012 );
not \U$17175 ( \17552 , \17550 );
and \U$17176 ( \17553 , \17552 , \1142 );
nor \U$17177 ( \17554 , \17551 , \17553 );
xor \U$17178 ( \17555 , \17547 , \17554 );
and \U$17179 ( \17556 , \1376 , RIae76c58_59);
and \U$17180 ( \17557 , RIae77180_70, \1374 );
nor \U$17181 ( \17558 , \17556 , \17557 );
and \U$17182 ( \17559 , \17558 , \1380 );
not \U$17183 ( \17560 , \17558 );
and \U$17184 ( \17561 , \17560 , \1261 );
nor \U$17185 ( \17562 , \17559 , \17561 );
and \U$17186 ( \17563 , \17555 , \17562 );
and \U$17187 ( \17564 , \17547 , \17554 );
or \U$17188 ( \17565 , \17563 , \17564 );
xor \U$17189 ( \17566 , \17540 , \17565 );
and \U$17190 ( \17567 , \2224 , RIae780f8_103);
and \U$17191 ( \17568 , RIae77f18_99, \2222 );
nor \U$17192 ( \17569 , \17567 , \17568 );
and \U$17193 ( \17570 , \17569 , \2061 );
not \U$17194 ( \17571 , \17569 );
and \U$17195 ( \17572 , \17571 , \2060 );
nor \U$17196 ( \17573 , \17570 , \17572 );
and \U$17197 ( \17574 , \1939 , RIae772e8_73);
and \U$17198 ( \17575 , RIae782d8_107, \1937 );
nor \U$17199 ( \17576 , \17574 , \17575 );
and \U$17200 ( \17577 , \17576 , \1735 );
not \U$17201 ( \17578 , \17576 );
and \U$17202 ( \17579 , \17578 , \1734 );
nor \U$17203 ( \17580 , \17577 , \17579 );
xor \U$17204 ( \17581 , \17573 , \17580 );
and \U$17205 ( \17582 , \2607 , RIae78008_101);
and \U$17206 ( \17583 , RIae781e8_105, \2605 );
nor \U$17207 ( \17584 , \17582 , \17583 );
and \U$17208 ( \17585 , \17584 , \2611 );
not \U$17209 ( \17586 , \17584 );
and \U$17210 ( \17587 , \17586 , \2397 );
nor \U$17211 ( \17588 , \17585 , \17587 );
and \U$17212 ( \17589 , \17581 , \17588 );
and \U$17213 ( \17590 , \17573 , \17580 );
or \U$17214 ( \17591 , \17589 , \17590 );
and \U$17215 ( \17592 , \17566 , \17591 );
and \U$17216 ( \17593 , \17540 , \17565 );
or \U$17217 ( \17594 , \17592 , \17593 );
and \U$17218 ( \17595 , \9760 , RIae75128_1);
and \U$17219 ( \17596 , RIae75308_5, \9758 );
nor \U$17220 ( \17597 , \17595 , \17596 );
and \U$17221 ( \17598 , \17597 , \9273 );
not \U$17222 ( \17599 , \17597 );
and \U$17223 ( \17600 , \17599 , \9764 );
nor \U$17224 ( \17601 , \17598 , \17600 );
and \U$17225 ( \17602 , \10548 , RIae753f8_7);
and \U$17226 ( \17603 , RIae763e8_41, \10546 );
nor \U$17227 ( \17604 , \17602 , \17603 );
and \U$17228 ( \17605 , \17604 , \10421 );
not \U$17229 ( \17606 , \17604 );
and \U$17230 ( \17607 , \17606 , \10118 );
nor \U$17231 ( \17608 , \17605 , \17607 );
xor \U$17232 ( \17609 , \17601 , \17608 );
and \U$17233 ( \17610 , \11470 , RIae764d8_43);
and \U$17234 ( \17611 , RIae766b8_47, \11468 );
nor \U$17235 ( \17612 , \17610 , \17611 );
and \U$17236 ( \17613 , \17612 , \10936 );
not \U$17237 ( \17614 , \17612 );
and \U$17238 ( \17615 , \17614 , \11474 );
nor \U$17239 ( \17616 , \17613 , \17615 );
and \U$17240 ( \17617 , \17609 , \17616 );
and \U$17241 ( \17618 , \17601 , \17608 );
or \U$17242 ( \17619 , \17617 , \17618 );
and \U$17243 ( \17620 , \15726 , RIae76898_51);
and \U$17244 ( \17621 , RIae7aab0_192, RIae76b68_57);
nor \U$17245 ( \17622 , \17620 , \17621 );
and \U$17246 ( \17623 , \17622 , \14959 );
not \U$17247 ( \17624 , \17622 );
and \U$17248 ( \17625 , \17624 , RIae7aa38_191);
nor \U$17249 ( \17626 , \17623 , \17625 );
xor \U$17250 ( \17627 , \17626 , \400 );
and \U$17251 ( \17628 , \14964 , RIae76988_53);
and \U$17252 ( \17629 , RIae767a8_49, \14962 );
nor \U$17253 ( \17630 , \17628 , \17629 );
and \U$17254 ( \17631 , \17630 , \14463 );
not \U$17255 ( \17632 , \17630 );
and \U$17256 ( \17633 , \17632 , \14462 );
nor \U$17257 ( \17634 , \17631 , \17633 );
and \U$17258 ( \17635 , \17627 , \17634 );
and \U$17259 ( \17636 , \17626 , \400 );
or \U$17260 ( \17637 , \17635 , \17636 );
xor \U$17261 ( \17638 , \17619 , \17637 );
and \U$17262 ( \17639 , \14059 , RIae76208_37);
and \U$17263 ( \17640 , RIae76a78_55, \14057 );
nor \U$17264 ( \17641 , \17639 , \17640 );
and \U$17265 ( \17642 , \17641 , \13502 );
not \U$17266 ( \17643 , \17641 );
and \U$17267 ( \17644 , \17643 , \14063 );
nor \U$17268 ( \17645 , \17642 , \17644 );
and \U$17269 ( \17646 , \12180 , RIae765c8_45);
and \U$17270 ( \17647 , RIae76118_35, \12178 );
nor \U$17271 ( \17648 , \17646 , \17647 );
and \U$17272 ( \17649 , \17648 , \12184 );
not \U$17273 ( \17650 , \17648 );
and \U$17274 ( \17651 , \17650 , \11827 );
nor \U$17275 ( \17652 , \17649 , \17651 );
xor \U$17276 ( \17653 , \17645 , \17652 );
and \U$17277 ( \17654 , \13059 , RIae76028_33);
and \U$17278 ( \17655 , RIae762f8_39, \13057 );
nor \U$17279 ( \17656 , \17654 , \17655 );
and \U$17280 ( \17657 , \17656 , \13063 );
not \U$17281 ( \17658 , \17656 );
and \U$17282 ( \17659 , \17658 , \12718 );
nor \U$17283 ( \17660 , \17657 , \17659 );
and \U$17284 ( \17661 , \17653 , \17660 );
and \U$17285 ( \17662 , \17645 , \17652 );
or \U$17286 ( \17663 , \17661 , \17662 );
and \U$17287 ( \17664 , \17638 , \17663 );
and \U$17288 ( \17665 , \17619 , \17637 );
or \U$17289 ( \17666 , \17664 , \17665 );
xor \U$17290 ( \17667 , \17594 , \17666 );
and \U$17291 ( \17668 , \8371 , RIae754e8_9);
and \U$17292 ( \17669 , RIae757b8_15, \8369 );
nor \U$17293 ( \17670 , \17668 , \17669 );
and \U$17294 ( \17671 , \17670 , \8020 );
not \U$17295 ( \17672 , \17670 );
and \U$17296 ( \17673 , \17672 , \8019 );
nor \U$17297 ( \17674 , \17671 , \17673 );
and \U$17298 ( \17675 , \7633 , RIae75d58_27);
and \U$17299 ( \17676 , RIae755d8_11, \7631 );
nor \U$17300 ( \17677 , \17675 , \17676 );
and \U$17301 ( \17678 , \17677 , \7206 );
not \U$17302 ( \17679 , \17677 );
and \U$17303 ( \17680 , \17679 , \7205 );
nor \U$17304 ( \17681 , \17678 , \17680 );
xor \U$17305 ( \17682 , \17674 , \17681 );
and \U$17306 ( \17683 , \8966 , RIae756c8_13);
and \U$17307 ( \17684 , RIae75218_3, \8964 );
nor \U$17308 ( \17685 , \17683 , \17684 );
and \U$17309 ( \17686 , \17685 , \8799 );
not \U$17310 ( \17687 , \17685 );
and \U$17311 ( \17688 , \17687 , \8789 );
nor \U$17312 ( \17689 , \17686 , \17688 );
and \U$17313 ( \17690 , \17682 , \17689 );
and \U$17314 ( \17691 , \17674 , \17681 );
or \U$17315 ( \17692 , \17690 , \17691 );
and \U$17316 ( \17693 , \5896 , RIae75a88_21);
and \U$17317 ( \17694 , RIae75998_19, \5894 );
nor \U$17318 ( \17695 , \17693 , \17694 );
and \U$17319 ( \17696 , \17695 , \5590 );
not \U$17320 ( \17697 , \17695 );
and \U$17321 ( \17698 , \17697 , \5589 );
nor \U$17322 ( \17699 , \17696 , \17698 );
and \U$17323 ( \17700 , \6172 , RIae758a8_17);
and \U$17324 ( \17701 , RIae75f38_31, \6170 );
nor \U$17325 ( \17702 , \17700 , \17701 );
and \U$17326 ( \17703 , \17702 , \6176 );
not \U$17327 ( \17704 , \17702 );
and \U$17328 ( \17705 , \17704 , \6175 );
nor \U$17329 ( \17706 , \17703 , \17705 );
xor \U$17330 ( \17707 , \17699 , \17706 );
and \U$17331 ( \17708 , \6941 , RIae75e48_29);
and \U$17332 ( \17709 , RIae75c68_25, \6939 );
nor \U$17333 ( \17710 , \17708 , \17709 );
and \U$17334 ( \17711 , \17710 , \6314 );
not \U$17335 ( \17712 , \17710 );
and \U$17336 ( \17713 , \17712 , \6945 );
nor \U$17337 ( \17714 , \17711 , \17713 );
and \U$17338 ( \17715 , \17707 , \17714 );
and \U$17339 ( \17716 , \17699 , \17706 );
or \U$17340 ( \17717 , \17715 , \17716 );
xor \U$17341 ( \17718 , \17692 , \17717 );
and \U$17342 ( \17719 , \5399 , RIae78698_115);
and \U$17343 ( \17720 , RIae75b78_23, \5397 );
nor \U$17344 ( \17721 , \17719 , \17720 );
and \U$17345 ( \17722 , \17721 , \5016 );
not \U$17346 ( \17723 , \17721 );
and \U$17347 ( \17724 , \17723 , \5403 );
nor \U$17348 ( \17725 , \17722 , \17724 );
and \U$17349 ( \17726 , \4247 , RIae77e28_97);
and \U$17350 ( \17727 , RIae78968_121, \4245 );
nor \U$17351 ( \17728 , \17726 , \17727 );
and \U$17352 ( \17729 , \17728 , \3989 );
not \U$17353 ( \17730 , \17728 );
and \U$17354 ( \17731 , \17730 , \4251 );
nor \U$17355 ( \17732 , \17729 , \17731 );
xor \U$17356 ( \17733 , \17725 , \17732 );
and \U$17357 ( \17734 , \4688 , RIae78878_119);
and \U$17358 ( \17735 , RIae78788_117, \4686 );
nor \U$17359 ( \17736 , \17734 , \17735 );
and \U$17360 ( \17737 , \17736 , \4481 );
not \U$17361 ( \17738 , \17736 );
and \U$17362 ( \17739 , \17738 , \4482 );
nor \U$17363 ( \17740 , \17737 , \17739 );
and \U$17364 ( \17741 , \17733 , \17740 );
and \U$17365 ( \17742 , \17725 , \17732 );
or \U$17366 ( \17743 , \17741 , \17742 );
and \U$17367 ( \17744 , \17718 , \17743 );
and \U$17368 ( \17745 , \17692 , \17717 );
or \U$17369 ( \17746 , \17744 , \17745 );
and \U$17370 ( \17747 , \17667 , \17746 );
and \U$17371 ( \17748 , \17594 , \17666 );
or \U$17372 ( \17749 , \17747 , \17748 );
xor \U$17373 ( \17750 , \17513 , \17749 );
xor \U$17374 ( \17751 , \17176 , \17183 );
xor \U$17375 ( \17752 , \17751 , \17191 );
xor \U$17376 ( \17753 , \17255 , \17262 );
xor \U$17377 ( \17754 , \17753 , \17270 );
and \U$17378 ( \17755 , \17752 , \17754 );
xor \U$17379 ( \17756 , \17306 , \17313 );
xor \U$17380 ( \17757 , \17756 , \17321 );
xor \U$17381 ( \17758 , \17255 , \17262 );
xor \U$17382 ( \17759 , \17758 , \17270 );
and \U$17383 ( \17760 , \17757 , \17759 );
and \U$17384 ( \17761 , \17752 , \17757 );
or \U$17385 ( \17762 , \17755 , \17760 , \17761 );
xor \U$17386 ( \17763 , \17414 , \17416 );
xor \U$17387 ( \17764 , \17763 , \17419 );
and \U$17388 ( \17765 , \17762 , \17764 );
xor \U$17389 ( \17766 , \16824 , \16831 );
xor \U$17390 ( \17767 , \17766 , \16839 );
xor \U$17391 ( \17768 , \17109 , \17114 );
xor \U$17392 ( \17769 , \17767 , \17768 );
xor \U$17393 ( \17770 , \17414 , \17416 );
xor \U$17394 ( \17771 , \17770 , \17419 );
and \U$17395 ( \17772 , \17769 , \17771 );
and \U$17396 ( \17773 , \17762 , \17769 );
or \U$17397 ( \17774 , \17765 , \17772 , \17773 );
and \U$17398 ( \17775 , \17750 , \17774 );
and \U$17399 ( \17776 , \17513 , \17749 );
or \U$17400 ( \17777 , \17775 , \17776 );
xor \U$17401 ( \17778 , \17434 , \17777 );
xor \U$17402 ( \17779 , \16646 , \16653 );
xor \U$17403 ( \17780 , \17779 , \16661 );
xor \U$17404 ( \17781 , \17158 , \17163 );
xor \U$17405 ( \17782 , \17780 , \17781 );
xor \U$17406 ( \17783 , \17353 , \17379 );
xor \U$17407 ( \17784 , \17783 , \17407 );
xor \U$17408 ( \17785 , \17782 , \17784 );
xor \U$17409 ( \17786 , \16918 , \16924 );
xor \U$17410 ( \17787 , \17786 , \16933 );
xor \U$17411 ( \17788 , \17145 , \17150 );
xor \U$17412 ( \17789 , \17787 , \17788 );
and \U$17413 ( \17790 , \17785 , \17789 );
and \U$17414 ( \17791 , \17782 , \17784 );
or \U$17415 ( \17792 , \17790 , \17791 );
xor \U$17416 ( \17793 , \16639 , \16664 );
xor \U$17417 ( \17794 , \17793 , \16690 );
xor \U$17418 ( \17795 , \16718 , \16736 );
xor \U$17419 ( \17796 , \17795 , \16762 );
xor \U$17420 ( \17797 , \17794 , \17796 );
xor \U$17421 ( \17798 , \16791 , \16816 );
xor \U$17422 ( \17799 , \17798 , \16842 );
xor \U$17423 ( \17800 , \17797 , \17799 );
and \U$17424 ( \17801 , \17792 , \17800 );
xor \U$17425 ( \17802 , \16977 , \16979 );
xor \U$17426 ( \17803 , \17802 , \16986 );
xor \U$17427 ( \17804 , \16936 , \16944 );
xor \U$17428 ( \17805 , \17804 , \16971 );
xor \U$17429 ( \17806 , \16896 , \16904 );
xor \U$17430 ( \17807 , \17806 , \16907 );
xor \U$17431 ( \17808 , \17805 , \17807 );
xor \U$17432 ( \17809 , \17803 , \17808 );
xor \U$17433 ( \17810 , \17794 , \17796 );
xor \U$17434 ( \17811 , \17810 , \17799 );
and \U$17435 ( \17812 , \17809 , \17811 );
and \U$17436 ( \17813 , \17792 , \17809 );
or \U$17437 ( \17814 , \17801 , \17812 , \17813 );
and \U$17438 ( \17815 , \17778 , \17814 );
and \U$17439 ( \17816 , \17434 , \17777 );
nor \U$17440 ( \17817 , \17815 , \17816 );
and \U$17441 ( \17818 , \17107 , \17817 );
and \U$17442 ( \17819 , \17104 , \17106 );
or \U$17443 ( \17820 , \17818 , \17819 );
not \U$17444 ( \17821 , \17820 );
not \U$17445 ( \17822 , \16097 );
not \U$17446 ( \17823 , \16061 );
or \U$17447 ( \17824 , \17822 , \17823 );
or \U$17448 ( \17825 , \16061 , \16097 );
nand \U$17449 ( \17826 , \17824 , \17825 );
not \U$17450 ( \17827 , \17826 );
not \U$17451 ( \17828 , \16071 );
and \U$17452 ( \17829 , \17827 , \17828 );
and \U$17453 ( \17830 , \17826 , \16071 );
nor \U$17454 ( \17831 , \17829 , \17830 );
not \U$17455 ( \17832 , \17831 );
xor \U$17456 ( \17833 , \17794 , \17796 );
and \U$17457 ( \17834 , \17833 , \17799 );
and \U$17458 ( \17835 , \17794 , \17796 );
or \U$17459 ( \17836 , \17834 , \17835 );
xor \U$17460 ( \17837 , \16295 , \16320 );
xor \U$17461 ( \17838 , \17837 , \16348 );
xor \U$17462 ( \17839 , \17836 , \17838 );
xor \U$17463 ( \17840 , \16977 , \16979 );
xor \U$17464 ( \17841 , \17840 , \16986 );
and \U$17465 ( \17842 , \17805 , \17841 );
xor \U$17466 ( \17843 , \16977 , \16979 );
xor \U$17467 ( \17844 , \17843 , \16986 );
and \U$17468 ( \17845 , \17807 , \17844 );
and \U$17469 ( \17846 , \17805 , \17807 );
or \U$17470 ( \17847 , \17842 , \17845 , \17846 );
and \U$17471 ( \17848 , \17839 , \17847 );
and \U$17472 ( \17849 , \17836 , \17838 );
or \U$17473 ( \17850 , \17848 , \17849 );
xor \U$17474 ( \17851 , \17119 , \17155 );
and \U$17475 ( \17852 , \17851 , \17168 );
and \U$17476 ( \17853 , \17119 , \17155 );
or \U$17477 ( \17854 , \17852 , \17853 );
xor \U$17478 ( \17855 , \17248 , \17327 );
and \U$17479 ( \17856 , \17855 , \17410 );
and \U$17480 ( \17857 , \17248 , \17327 );
or \U$17481 ( \17858 , \17856 , \17857 );
xor \U$17482 ( \17859 , \17854 , \17858 );
xor \U$17483 ( \17860 , \17422 , \17427 );
and \U$17484 ( \17861 , \17860 , \17430 );
and \U$17485 ( \17862 , \17422 , \17427 );
or \U$17486 ( \17863 , \17861 , \17862 );
and \U$17487 ( \17864 , \17859 , \17863 );
and \U$17488 ( \17865 , \17854 , \17858 );
or \U$17489 ( \17866 , \17864 , \17865 );
and \U$17490 ( \17867 , \17850 , \17866 );
not \U$17491 ( \17868 , \17850 );
not \U$17492 ( \17869 , \17866 );
and \U$17493 ( \17870 , \17868 , \17869 );
xor \U$17494 ( \17871 , \17088 , \17090 );
and \U$17495 ( \17872 , \17871 , \17101 );
and \U$17496 ( \17873 , \17088 , \17090 );
or \U$17497 ( \17874 , \17872 , \17873 );
nor \U$17498 ( \17875 , \17870 , \17874 );
nor \U$17499 ( \17876 , \17867 , \17875 );
xor \U$17500 ( \17877 , \17001 , \17013 );
xor \U$17501 ( \17878 , \17877 , \17030 );
not \U$17502 ( \17879 , \16181 );
xor \U$17503 ( \17880 , \16351 , \16267 );
not \U$17504 ( \17881 , \17880 );
or \U$17505 ( \17882 , \17879 , \17881 );
or \U$17506 ( \17883 , \17880 , \16181 );
nand \U$17507 ( \17884 , \17882 , \17883 );
xor \U$17508 ( \17885 , \17878 , \17884 );
not \U$17509 ( \17886 , \17036 );
xor \U$17510 ( \17887 , \17039 , \17052 );
not \U$17511 ( \17888 , \17887 );
or \U$17512 ( \17889 , \17886 , \17888 );
or \U$17513 ( \17890 , \17887 , \17036 );
nand \U$17514 ( \17891 , \17889 , \17890 );
and \U$17515 ( \17892 , \17885 , \17891 );
and \U$17516 ( \17893 , \17878 , \17884 );
nor \U$17517 ( \17894 , \17892 , \17893 );
xor \U$17518 ( \17895 , \17876 , \17894 );
not \U$17519 ( \17896 , \17895 );
or \U$17520 ( \17897 , \17832 , \17896 );
or \U$17521 ( \17898 , \17895 , \17831 );
nand \U$17522 ( \17899 , \17897 , \17898 );
not \U$17523 ( \17900 , \17899 );
or \U$17524 ( \17901 , \17821 , \17900 );
or \U$17525 ( \17902 , \17899 , \17820 );
nand \U$17526 ( \17903 , \17901 , \17902 );
not \U$17527 ( \17904 , \17903 );
xor \U$17528 ( \17905 , \16353 , \16438 );
xor \U$17529 ( \17906 , \17905 , \16476 );
xor \U$17530 ( \17907 , \16995 , \17033 );
xor \U$17531 ( \17908 , \17907 , \17054 );
xnor \U$17532 ( \17909 , \17906 , \17908 );
not \U$17533 ( \17910 , \17909 );
xor \U$17534 ( \17911 , \15909 , \15967 );
xor \U$17535 ( \17912 , \17911 , \15980 );
xor \U$17536 ( \17913 , \16597 , \16604 );
xor \U$17537 ( \17914 , \17912 , \17913 );
not \U$17538 ( \17915 , \17914 );
and \U$17539 ( \17916 , \17910 , \17915 );
and \U$17540 ( \17917 , \17909 , \17914 );
nor \U$17541 ( \17918 , \17916 , \17917 );
not \U$17542 ( \17919 , \17918 );
and \U$17543 ( \17920 , \17904 , \17919 );
and \U$17544 ( \17921 , \17903 , \17918 );
nor \U$17545 ( \17922 , \17920 , \17921 );
not \U$17546 ( \17923 , \17922 );
xor \U$17547 ( \17924 , \17104 , \17106 );
xor \U$17548 ( \17925 , \17924 , \17817 );
not \U$17549 ( \17926 , \17925 );
not \U$17550 ( \17927 , \17874 );
xor \U$17551 ( \17928 , \17866 , \17850 );
not \U$17552 ( \17929 , \17928 );
or \U$17553 ( \17930 , \17927 , \17929 );
or \U$17554 ( \17931 , \17928 , \17874 );
nand \U$17555 ( \17932 , \17930 , \17931 );
nand \U$17556 ( \17933 , \17926 , \17932 );
not \U$17557 ( \17934 , \17933 );
xor \U$17558 ( \17935 , \17074 , \17072 );
not \U$17559 ( \17936 , \17935 );
not \U$17560 ( \17937 , \17102 );
or \U$17561 ( \17938 , \17936 , \17937 );
or \U$17562 ( \17939 , \17102 , \17935 );
nand \U$17563 ( \17940 , \17938 , \17939 );
xor \U$17564 ( \17941 , \17854 , \17858 );
xor \U$17565 ( \17942 , \17941 , \17863 );
xor \U$17566 ( \17943 , \17940 , \17942 );
xor \U$17567 ( \17944 , \17434 , \17777 );
xor \U$17568 ( \17945 , \17944 , \17814 );
and \U$17569 ( \17946 , \17943 , \17945 );
and \U$17570 ( \17947 , \17940 , \17942 );
or \U$17571 ( \17948 , \17946 , \17947 );
xor \U$17572 ( \17949 , \17878 , \17884 );
xor \U$17573 ( \17950 , \17949 , \17891 );
xor \U$17574 ( \17951 , \17948 , \17950 );
xor \U$17575 ( \17952 , \17540 , \17565 );
xor \U$17576 ( \17953 , \17952 , \17591 );
xor \U$17577 ( \17954 , \17619 , \17637 );
xor \U$17578 ( \17955 , \17954 , \17663 );
and \U$17579 ( \17956 , \17953 , \17955 );
xor \U$17580 ( \17957 , \17692 , \17717 );
xor \U$17581 ( \17958 , \17957 , \17743 );
xor \U$17582 ( \17959 , \17619 , \17637 );
xor \U$17583 ( \17960 , \17959 , \17663 );
and \U$17584 ( \17961 , \17958 , \17960 );
and \U$17585 ( \17962 , \17953 , \17958 );
or \U$17586 ( \17963 , \17956 , \17961 , \17962 );
xor \U$17587 ( \17964 , \17194 , \17219 );
xor \U$17588 ( \17965 , \17964 , \17245 );
xor \U$17589 ( \17966 , \17963 , \17965 );
xor \U$17590 ( \17967 , \17461 , \17469 );
xor \U$17591 ( \17968 , \17967 , \17496 );
xor \U$17592 ( \17969 , \17502 , \17504 );
xor \U$17593 ( \17970 , \17969 , \17507 );
and \U$17594 ( \17971 , \17968 , \17970 );
xor \U$17595 ( \17972 , \17201 , \17208 );
xor \U$17596 ( \17973 , \17972 , \17216 );
xor \U$17597 ( \17974 , \17436 , \17441 );
xor \U$17598 ( \17975 , \17973 , \17974 );
xor \U$17599 ( \17976 , \17502 , \17504 );
xor \U$17600 ( \17977 , \17976 , \17507 );
and \U$17601 ( \17978 , \17975 , \17977 );
and \U$17602 ( \17979 , \17968 , \17975 );
or \U$17603 ( \17980 , \17971 , \17978 , \17979 );
and \U$17604 ( \17981 , \17966 , \17980 );
and \U$17605 ( \17982 , \17963 , \17965 );
or \U$17606 ( \17983 , \17981 , \17982 );
xor \U$17607 ( \17984 , \17626 , \400 );
xor \U$17608 ( \17985 , \17984 , \17634 );
xor \U$17609 ( \17986 , \17645 , \17652 );
xor \U$17610 ( \17987 , \17986 , \17660 );
and \U$17611 ( \17988 , \17985 , \17987 );
xor \U$17612 ( \17989 , \17601 , \17608 );
xor \U$17613 ( \17990 , \17989 , \17616 );
xor \U$17614 ( \17991 , \17645 , \17652 );
xor \U$17615 ( \17992 , \17991 , \17660 );
and \U$17616 ( \17993 , \17990 , \17992 );
and \U$17617 ( \17994 , \17985 , \17990 );
or \U$17618 ( \17995 , \17988 , \17993 , \17994 );
xor \U$17619 ( \17996 , \17280 , \17287 );
xor \U$17620 ( \17997 , \17996 , \17295 );
xor \U$17621 ( \17998 , \17995 , \17997 );
xor \U$17622 ( \17999 , \17255 , \17262 );
xor \U$17623 ( \18000 , \17999 , \17270 );
xor \U$17624 ( \18001 , \17752 , \17757 );
xor \U$17625 ( \18002 , \18000 , \18001 );
and \U$17626 ( \18003 , \17998 , \18002 );
and \U$17627 ( \18004 , \17995 , \17997 );
or \U$17628 ( \18005 , \18003 , \18004 );
and \U$17629 ( \18006 , \1939 , RIae771f8_71);
and \U$17630 ( \18007 , RIae772e8_73, \1937 );
nor \U$17631 ( \18008 , \18006 , \18007 );
and \U$17632 ( \18009 , \18008 , \1735 );
not \U$17633 ( \18010 , \18008 );
and \U$17634 ( \18011 , \18010 , \1734 );
nor \U$17635 ( \18012 , \18009 , \18011 );
and \U$17636 ( \18013 , \1593 , RIae77180_70);
and \U$17637 ( \18014 , RIae77018_67, \1591 );
nor \U$17638 ( \18015 , \18013 , \18014 );
and \U$17639 ( \18016 , \18015 , \1498 );
not \U$17640 ( \18017 , \18015 );
and \U$17641 ( \18018 , \18017 , \1488 );
nor \U$17642 ( \18019 , \18016 , \18018 );
xor \U$17643 ( \18020 , \18012 , \18019 );
and \U$17644 ( \18021 , \2224 , RIae782d8_107);
and \U$17645 ( \18022 , RIae780f8_103, \2222 );
nor \U$17646 ( \18023 , \18021 , \18022 );
and \U$17647 ( \18024 , \18023 , \2061 );
not \U$17648 ( \18025 , \18023 );
and \U$17649 ( \18026 , \18025 , \2060 );
nor \U$17650 ( \18027 , \18024 , \18026 );
and \U$17651 ( \18028 , \18020 , \18027 );
and \U$17652 ( \18029 , \18012 , \18019 );
or \U$17653 ( \18030 , \18028 , \18029 );
and \U$17654 ( \18031 , \1138 , RIae76f28_65);
and \U$17655 ( \18032 , RIae76e38_63, \1136 );
nor \U$17656 ( \18033 , \18031 , \18032 );
and \U$17657 ( \18034 , \18033 , \1012 );
not \U$17658 ( \18035 , \18033 );
and \U$17659 ( \18036 , \18035 , \1142 );
nor \U$17660 ( \18037 , \18034 , \18036 );
not \U$17661 ( \18038 , \789 );
and \U$17662 ( \18039 , \883 , RIae77798_83);
and \U$17663 ( \18040 , RIae77888_85, \881 );
nor \U$17664 ( \18041 , \18039 , \18040 );
not \U$17665 ( \18042 , \18041 );
or \U$17666 ( \18043 , \18038 , \18042 );
or \U$17667 ( \18044 , \18041 , \787 );
nand \U$17668 ( \18045 , \18043 , \18044 );
xor \U$17669 ( \18046 , \18037 , \18045 );
and \U$17670 ( \18047 , \1376 , RIae76d48_61);
and \U$17671 ( \18048 , RIae76c58_59, \1374 );
nor \U$17672 ( \18049 , \18047 , \18048 );
and \U$17673 ( \18050 , \18049 , \1380 );
not \U$17674 ( \18051 , \18049 );
and \U$17675 ( \18052 , \18051 , \1261 );
nor \U$17676 ( \18053 , \18050 , \18052 );
and \U$17677 ( \18054 , \18046 , \18053 );
and \U$17678 ( \18055 , \18037 , \18045 );
or \U$17679 ( \18056 , \18054 , \18055 );
xor \U$17680 ( \18057 , \18030 , \18056 );
not \U$17681 ( \18058 , \3218 );
and \U$17682 ( \18059 , \3214 , RIae783c8_109);
and \U$17683 ( \18060 , RIae78530_112, \3212 );
nor \U$17684 ( \18061 , \18059 , \18060 );
not \U$17685 ( \18062 , \18061 );
or \U$17686 ( \18063 , \18058 , \18062 );
or \U$17687 ( \18064 , \18061 , \2774 );
nand \U$17688 ( \18065 , \18063 , \18064 );
and \U$17689 ( \18066 , \2607 , RIae77f18_99);
and \U$17690 ( \18067 , RIae78008_101, \2605 );
nor \U$17691 ( \18068 , \18066 , \18067 );
and \U$17692 ( \18069 , \18068 , \2611 );
not \U$17693 ( \18070 , \18068 );
and \U$17694 ( \18071 , \18070 , \2397 );
nor \U$17695 ( \18072 , \18069 , \18071 );
xor \U$17696 ( \18073 , \18065 , \18072 );
not \U$17697 ( \18074 , \3089 );
and \U$17698 ( \18075 , \2783 , RIae781e8_105);
and \U$17699 ( \18076 , RIae785a8_113, \2781 );
nor \U$17700 ( \18077 , \18075 , \18076 );
not \U$17701 ( \18078 , \18077 );
or \U$17702 ( \18079 , \18074 , \18078 );
or \U$17703 ( \18080 , \18077 , \3089 );
nand \U$17704 ( \18081 , \18079 , \18080 );
and \U$17705 ( \18082 , \18073 , \18081 );
and \U$17706 ( \18083 , \18065 , \18072 );
or \U$17707 ( \18084 , \18082 , \18083 );
and \U$17708 ( \18085 , \18057 , \18084 );
and \U$17709 ( \18086 , \18030 , \18056 );
or \U$17710 ( \18087 , \18085 , \18086 );
and \U$17711 ( \18088 , \10548 , RIae75308_5);
and \U$17712 ( \18089 , RIae753f8_7, \10546 );
nor \U$17713 ( \18090 , \18088 , \18089 );
and \U$17714 ( \18091 , \18090 , \10421 );
not \U$17715 ( \18092 , \18090 );
and \U$17716 ( \18093 , \18092 , \10118 );
nor \U$17717 ( \18094 , \18091 , \18093 );
and \U$17718 ( \18095 , \8966 , RIae757b8_15);
and \U$17719 ( \18096 , RIae756c8_13, \8964 );
nor \U$17720 ( \18097 , \18095 , \18096 );
and \U$17721 ( \18098 , \18097 , \8799 );
not \U$17722 ( \18099 , \18097 );
and \U$17723 ( \18100 , \18099 , \8789 );
nor \U$17724 ( \18101 , \18098 , \18100 );
xor \U$17725 ( \18102 , \18094 , \18101 );
and \U$17726 ( \18103 , \9760 , RIae75218_3);
and \U$17727 ( \18104 , RIae75128_1, \9758 );
nor \U$17728 ( \18105 , \18103 , \18104 );
and \U$17729 ( \18106 , \18105 , \9273 );
not \U$17730 ( \18107 , \18105 );
and \U$17731 ( \18108 , \18107 , \9764 );
nor \U$17732 ( \18109 , \18106 , \18108 );
and \U$17733 ( \18110 , \18102 , \18109 );
and \U$17734 ( \18111 , \18094 , \18101 );
or \U$17735 ( \18112 , \18110 , \18111 );
and \U$17736 ( \18113 , \14059 , RIae762f8_39);
and \U$17737 ( \18114 , RIae76208_37, \14057 );
nor \U$17738 ( \18115 , \18113 , \18114 );
and \U$17739 ( \18116 , \18115 , \13502 );
not \U$17740 ( \18117 , \18115 );
and \U$17741 ( \18118 , \18117 , \14063 );
nor \U$17742 ( \18119 , \18116 , \18118 );
and \U$17743 ( \18120 , \15726 , RIae767a8_49);
and \U$17744 ( \18121 , RIae7aab0_192, RIae76898_51);
nor \U$17745 ( \18122 , \18120 , \18121 );
and \U$17746 ( \18123 , \18122 , \14959 );
not \U$17747 ( \18124 , \18122 );
and \U$17748 ( \18125 , \18124 , RIae7aa38_191);
nor \U$17749 ( \18126 , \18123 , \18125 );
xor \U$17750 ( \18127 , \18119 , \18126 );
and \U$17751 ( \18128 , \14964 , RIae76a78_55);
and \U$17752 ( \18129 , RIae76988_53, \14962 );
nor \U$17753 ( \18130 , \18128 , \18129 );
and \U$17754 ( \18131 , \18130 , \14463 );
not \U$17755 ( \18132 , \18130 );
and \U$17756 ( \18133 , \18132 , \14462 );
nor \U$17757 ( \18134 , \18131 , \18133 );
and \U$17758 ( \18135 , \18127 , \18134 );
and \U$17759 ( \18136 , \18119 , \18126 );
or \U$17760 ( \18137 , \18135 , \18136 );
xor \U$17761 ( \18138 , \18112 , \18137 );
and \U$17762 ( \18139 , \11470 , RIae763e8_41);
and \U$17763 ( \18140 , RIae764d8_43, \11468 );
nor \U$17764 ( \18141 , \18139 , \18140 );
and \U$17765 ( \18142 , \18141 , \10936 );
not \U$17766 ( \18143 , \18141 );
and \U$17767 ( \18144 , \18143 , \11474 );
nor \U$17768 ( \18145 , \18142 , \18144 );
and \U$17769 ( \18146 , \12180 , RIae766b8_47);
and \U$17770 ( \18147 , RIae765c8_45, \12178 );
nor \U$17771 ( \18148 , \18146 , \18147 );
and \U$17772 ( \18149 , \18148 , \12184 );
not \U$17773 ( \18150 , \18148 );
and \U$17774 ( \18151 , \18150 , \11827 );
nor \U$17775 ( \18152 , \18149 , \18151 );
xor \U$17776 ( \18153 , \18145 , \18152 );
and \U$17777 ( \18154 , \13059 , RIae76118_35);
and \U$17778 ( \18155 , RIae76028_33, \13057 );
nor \U$17779 ( \18156 , \18154 , \18155 );
and \U$17780 ( \18157 , \18156 , \13063 );
not \U$17781 ( \18158 , \18156 );
and \U$17782 ( \18159 , \18158 , \12718 );
nor \U$17783 ( \18160 , \18157 , \18159 );
and \U$17784 ( \18161 , \18153 , \18160 );
and \U$17785 ( \18162 , \18145 , \18152 );
or \U$17786 ( \18163 , \18161 , \18162 );
and \U$17787 ( \18164 , \18138 , \18163 );
and \U$17788 ( \18165 , \18112 , \18137 );
or \U$17789 ( \18166 , \18164 , \18165 );
xor \U$17790 ( \18167 , \18087 , \18166 );
and \U$17791 ( \18168 , \7633 , RIae75c68_25);
and \U$17792 ( \18169 , RIae75d58_27, \7631 );
nor \U$17793 ( \18170 , \18168 , \18169 );
and \U$17794 ( \18171 , \18170 , \7206 );
not \U$17795 ( \18172 , \18170 );
and \U$17796 ( \18173 , \18172 , \7205 );
nor \U$17797 ( \18174 , \18171 , \18173 );
and \U$17798 ( \18175 , \6941 , RIae75f38_31);
and \U$17799 ( \18176 , RIae75e48_29, \6939 );
nor \U$17800 ( \18177 , \18175 , \18176 );
and \U$17801 ( \18178 , \18177 , \6314 );
not \U$17802 ( \18179 , \18177 );
and \U$17803 ( \18180 , \18179 , \6945 );
nor \U$17804 ( \18181 , \18178 , \18180 );
xor \U$17805 ( \18182 , \18174 , \18181 );
and \U$17806 ( \18183 , \8371 , RIae755d8_11);
and \U$17807 ( \18184 , RIae754e8_9, \8369 );
nor \U$17808 ( \18185 , \18183 , \18184 );
and \U$17809 ( \18186 , \18185 , \8020 );
not \U$17810 ( \18187 , \18185 );
and \U$17811 ( \18188 , \18187 , \8019 );
nor \U$17812 ( \18189 , \18186 , \18188 );
and \U$17813 ( \18190 , \18182 , \18189 );
and \U$17814 ( \18191 , \18174 , \18181 );
or \U$17815 ( \18192 , \18190 , \18191 );
and \U$17816 ( \18193 , \4688 , RIae78968_121);
and \U$17817 ( \18194 , RIae78878_119, \4686 );
nor \U$17818 ( \18195 , \18193 , \18194 );
and \U$17819 ( \18196 , \18195 , \4481 );
not \U$17820 ( \18197 , \18195 );
and \U$17821 ( \18198 , \18197 , \4482 );
nor \U$17822 ( \18199 , \18196 , \18198 );
and \U$17823 ( \18200 , \3730 , RIae77c48_93);
and \U$17824 ( \18201 , RIae77b58_91, \3728 );
nor \U$17825 ( \18202 , \18200 , \18201 );
and \U$17826 ( \18203 , \18202 , \3732 );
not \U$17827 ( \18204 , \18202 );
and \U$17828 ( \18205 , \18204 , \3422 );
nor \U$17829 ( \18206 , \18203 , \18205 );
xor \U$17830 ( \18207 , \18199 , \18206 );
and \U$17831 ( \18208 , \4247 , RIae77d38_95);
and \U$17832 ( \18209 , RIae77e28_97, \4245 );
nor \U$17833 ( \18210 , \18208 , \18209 );
and \U$17834 ( \18211 , \18210 , \3989 );
not \U$17835 ( \18212 , \18210 );
and \U$17836 ( \18213 , \18212 , \4251 );
nor \U$17837 ( \18214 , \18211 , \18213 );
and \U$17838 ( \18215 , \18207 , \18214 );
and \U$17839 ( \18216 , \18199 , \18206 );
or \U$17840 ( \18217 , \18215 , \18216 );
xor \U$17841 ( \18218 , \18192 , \18217 );
and \U$17842 ( \18219 , \5399 , RIae78788_117);
and \U$17843 ( \18220 , RIae78698_115, \5397 );
nor \U$17844 ( \18221 , \18219 , \18220 );
and \U$17845 ( \18222 , \18221 , \5016 );
not \U$17846 ( \18223 , \18221 );
and \U$17847 ( \18224 , \18223 , \5403 );
nor \U$17848 ( \18225 , \18222 , \18224 );
and \U$17849 ( \18226 , \5896 , RIae75b78_23);
and \U$17850 ( \18227 , RIae75a88_21, \5894 );
nor \U$17851 ( \18228 , \18226 , \18227 );
and \U$17852 ( \18229 , \18228 , \5590 );
not \U$17853 ( \18230 , \18228 );
and \U$17854 ( \18231 , \18230 , \5589 );
nor \U$17855 ( \18232 , \18229 , \18231 );
xor \U$17856 ( \18233 , \18225 , \18232 );
and \U$17857 ( \18234 , \6172 , RIae75998_19);
and \U$17858 ( \18235 , RIae758a8_17, \6170 );
nor \U$17859 ( \18236 , \18234 , \18235 );
and \U$17860 ( \18237 , \18236 , \6176 );
not \U$17861 ( \18238 , \18236 );
and \U$17862 ( \18239 , \18238 , \6175 );
nor \U$17863 ( \18240 , \18237 , \18239 );
and \U$17864 ( \18241 , \18233 , \18240 );
and \U$17865 ( \18242 , \18225 , \18232 );
or \U$17866 ( \18243 , \18241 , \18242 );
and \U$17867 ( \18244 , \18218 , \18243 );
and \U$17868 ( \18245 , \18192 , \18217 );
or \U$17869 ( \18246 , \18244 , \18245 );
and \U$17870 ( \18247 , \18167 , \18246 );
and \U$17871 ( \18248 , \18087 , \18166 );
or \U$17872 ( \18249 , \18247 , \18248 );
xor \U$17873 ( \18250 , \18005 , \18249 );
xor \U$17874 ( \18251 , \17520 , \17528 );
xor \U$17875 ( \18252 , \18251 , \17537 );
xor \U$17876 ( \18253 , \17547 , \17554 );
xor \U$17877 ( \18254 , \18253 , \17562 );
xor \U$17878 ( \18255 , \18252 , \18254 );
xor \U$17879 ( \18256 , \17573 , \17580 );
xor \U$17880 ( \18257 , \18256 , \17588 );
and \U$17881 ( \18258 , \18255 , \18257 );
and \U$17882 ( \18259 , \18252 , \18254 );
or \U$17883 ( \18260 , \18258 , \18259 );
and \U$17884 ( \18261 , \672 , RIae77a68_89);
and \U$17885 ( \18262 , RIae77978_87, \670 );
nor \U$17886 ( \18263 , \18261 , \18262 );
and \U$17887 ( \18264 , \18263 , \588 );
not \U$17888 ( \18265 , \18263 );
and \U$17889 ( \18266 , \18265 , \587 );
nor \U$17890 ( \18267 , \18264 , \18266 );
not \U$17891 ( \18268 , \469 );
and \U$17892 ( \18269 , \514 , RIae775b8_79);
and \U$17893 ( \18270 , RIae774c8_77, \512 );
nor \U$17894 ( \18271 , \18269 , \18270 );
not \U$17895 ( \18272 , \18271 );
or \U$17896 ( \18273 , \18268 , \18272 );
or \U$17897 ( \18274 , \18271 , \471 );
nand \U$17898 ( \18275 , \18273 , \18274 );
xor \U$17899 ( \18276 , \18267 , \18275 );
and \U$17900 ( \18277 , \558 , RIae77720_82);
and \U$17901 ( \18278 , RIae773d8_75, \556 );
nor \U$17902 ( \18279 , \18277 , \18278 );
and \U$17903 ( \18280 , \18279 , \504 );
not \U$17904 ( \18281 , \18279 );
and \U$17905 ( \18282 , \18281 , \562 );
nor \U$17906 ( \18283 , \18280 , \18282 );
and \U$17907 ( \18284 , \18276 , \18283 );
and \U$17908 ( \18285 , \18267 , \18275 );
or \U$17909 ( \18286 , \18284 , \18285 );
xor \U$17910 ( \18287 , \17452 , \17460 );
xor \U$17911 ( \18288 , \18286 , \18287 );
xor \U$17912 ( \18289 , \17478 , \17485 );
xor \U$17913 ( \18290 , \18289 , \17493 );
and \U$17914 ( \18291 , \18288 , \18290 );
and \U$17915 ( \18292 , \18286 , \18287 );
or \U$17916 ( \18293 , \18291 , \18292 );
xor \U$17917 ( \18294 , \18260 , \18293 );
xor \U$17918 ( \18295 , \17699 , \17706 );
xor \U$17919 ( \18296 , \18295 , \17714 );
xor \U$17920 ( \18297 , \17725 , \17732 );
xor \U$17921 ( \18298 , \18297 , \17740 );
and \U$17922 ( \18299 , \18296 , \18298 );
xor \U$17923 ( \18300 , \17674 , \17681 );
xor \U$17924 ( \18301 , \18300 , \17689 );
xor \U$17925 ( \18302 , \17725 , \17732 );
xor \U$17926 ( \18303 , \18302 , \17740 );
and \U$17927 ( \18304 , \18301 , \18303 );
and \U$17928 ( \18305 , \18296 , \18301 );
or \U$17929 ( \18306 , \18299 , \18304 , \18305 );
and \U$17930 ( \18307 , \18294 , \18306 );
and \U$17931 ( \18308 , \18260 , \18293 );
or \U$17932 ( \18309 , \18307 , \18308 );
and \U$17933 ( \18310 , \18250 , \18309 );
and \U$17934 ( \18311 , \18005 , \18249 );
or \U$17935 ( \18312 , \18310 , \18311 );
xor \U$17936 ( \18313 , \17983 , \18312 );
xor \U$17937 ( \18314 , \17273 , \17298 );
xor \U$17938 ( \18315 , \18314 , \17324 );
xor \U$17939 ( \18316 , \17782 , \17784 );
xor \U$17940 ( \18317 , \18316 , \17789 );
and \U$17941 ( \18318 , \18315 , \18317 );
xor \U$17942 ( \18319 , \17414 , \17416 );
xor \U$17943 ( \18320 , \18319 , \17419 );
xor \U$17944 ( \18321 , \17762 , \17769 );
xor \U$17945 ( \18322 , \18320 , \18321 );
xor \U$17946 ( \18323 , \17782 , \17784 );
xor \U$17947 ( \18324 , \18323 , \17789 );
and \U$17948 ( \18325 , \18322 , \18324 );
and \U$17949 ( \18326 , \18315 , \18322 );
or \U$17950 ( \18327 , \18318 , \18325 , \18326 );
and \U$17951 ( \18328 , \18313 , \18327 );
and \U$17952 ( \18329 , \17983 , \18312 );
or \U$17953 ( \18330 , \18328 , \18329 );
xor \U$17954 ( \18331 , \17836 , \17838 );
xor \U$17955 ( \18332 , \18331 , \17847 );
xor \U$17956 ( \18333 , \18330 , \18332 );
xor \U$17957 ( \18334 , \17513 , \17749 );
xor \U$17958 ( \18335 , \18334 , \17774 );
xor \U$17959 ( \18336 , \17169 , \17411 );
xor \U$17960 ( \18337 , \18336 , \17431 );
and \U$17961 ( \18338 , \18335 , \18337 );
xor \U$17962 ( \18339 , \17794 , \17796 );
xor \U$17963 ( \18340 , \18339 , \17799 );
xor \U$17964 ( \18341 , \17792 , \17809 );
xor \U$17965 ( \18342 , \18340 , \18341 );
xor \U$17966 ( \18343 , \17169 , \17411 );
xor \U$17967 ( \18344 , \18343 , \17431 );
and \U$17968 ( \18345 , \18342 , \18344 );
and \U$17969 ( \18346 , \18335 , \18342 );
or \U$17970 ( \18347 , \18338 , \18345 , \18346 );
and \U$17971 ( \18348 , \18333 , \18347 );
and \U$17972 ( \18349 , \18330 , \18332 );
or \U$17973 ( \18350 , \18348 , \18349 );
and \U$17974 ( \18351 , \17951 , \18350 );
and \U$17975 ( \18352 , \17948 , \17950 );
or \U$17976 ( \18353 , \18351 , \18352 );
not \U$17977 ( \18354 , \18353 );
or \U$17978 ( \18355 , \17934 , \18354 );
or \U$17979 ( \18356 , \18353 , \17933 );
nand \U$17980 ( \18357 , \18355 , \18356 );
not \U$17981 ( \18358 , \18357 );
or \U$17982 ( \18359 , \17923 , \18358 );
or \U$17983 ( \18360 , \18357 , \17922 );
nand \U$17984 ( \18361 , \18359 , \18360 );
xor \U$17985 ( \18362 , \18087 , \18166 );
xor \U$17986 ( \18363 , \18362 , \18246 );
xor \U$17987 ( \18364 , \17995 , \17997 );
xor \U$17988 ( \18365 , \18364 , \18002 );
and \U$17989 ( \18366 , \18363 , \18365 );
xor \U$17990 ( \18367 , \18260 , \18293 );
xor \U$17991 ( \18368 , \18367 , \18306 );
xor \U$17992 ( \18369 , \17995 , \17997 );
xor \U$17993 ( \18370 , \18369 , \18002 );
and \U$17994 ( \18371 , \18368 , \18370 );
and \U$17995 ( \18372 , \18363 , \18368 );
or \U$17996 ( \18373 , \18366 , \18371 , \18372 );
xor \U$17997 ( \18374 , \18065 , \18072 );
xor \U$17998 ( \18375 , \18374 , \18081 );
xor \U$17999 ( \18376 , \18012 , \18019 );
xor \U$18000 ( \18377 , \18376 , \18027 );
xor \U$18001 ( \18378 , \18375 , \18377 );
xor \U$18002 ( \18379 , \18199 , \18206 );
xor \U$18003 ( \18380 , \18379 , \18214 );
and \U$18004 ( \18381 , \18378 , \18380 );
and \U$18005 ( \18382 , \18375 , \18377 );
or \U$18006 ( \18383 , \18381 , \18382 );
and \U$18007 ( \18384 , \558 , RIae774c8_77);
and \U$18008 ( \18385 , RIae77720_82, \556 );
nor \U$18009 ( \18386 , \18384 , \18385 );
and \U$18010 ( \18387 , \18386 , \504 );
not \U$18011 ( \18388 , \18386 );
and \U$18012 ( \18389 , \18388 , \562 );
nor \U$18013 ( \18390 , \18387 , \18389 );
and \U$18014 ( \18391 , \672 , RIae773d8_75);
and \U$18015 ( \18392 , RIae77a68_89, \670 );
nor \U$18016 ( \18393 , \18391 , \18392 );
and \U$18017 ( \18394 , \18393 , \588 );
not \U$18018 ( \18395 , \18393 );
and \U$18019 ( \18396 , \18395 , \587 );
nor \U$18020 ( \18397 , \18394 , \18396 );
xor \U$18021 ( \18398 , \18390 , \18397 );
not \U$18022 ( \18399 , \787 );
and \U$18023 ( \18400 , \883 , RIae77978_87);
and \U$18024 ( \18401 , RIae77798_83, \881 );
nor \U$18025 ( \18402 , \18400 , \18401 );
not \U$18026 ( \18403 , \18402 );
or \U$18027 ( \18404 , \18399 , \18403 );
or \U$18028 ( \18405 , \18402 , \789 );
nand \U$18029 ( \18406 , \18404 , \18405 );
and \U$18030 ( \18407 , \18398 , \18406 );
and \U$18031 ( \18408 , \18390 , \18397 );
or \U$18032 ( \18409 , \18407 , \18408 );
xor \U$18033 ( \18410 , \18267 , \18275 );
xor \U$18034 ( \18411 , \18410 , \18283 );
and \U$18035 ( \18412 , \18409 , \18411 );
xor \U$18036 ( \18413 , \18037 , \18045 );
xor \U$18037 ( \18414 , \18413 , \18053 );
xor \U$18038 ( \18415 , \18267 , \18275 );
xor \U$18039 ( \18416 , \18415 , \18283 );
and \U$18040 ( \18417 , \18414 , \18416 );
and \U$18041 ( \18418 , \18409 , \18414 );
or \U$18042 ( \18419 , \18412 , \18417 , \18418 );
xor \U$18043 ( \18420 , \18383 , \18419 );
xor \U$18044 ( \18421 , \18225 , \18232 );
xor \U$18045 ( \18422 , \18421 , \18240 );
xor \U$18046 ( \18423 , \18174 , \18181 );
xor \U$18047 ( \18424 , \18423 , \18189 );
and \U$18048 ( \18425 , \18422 , \18424 );
xor \U$18049 ( \18426 , \18094 , \18101 );
xor \U$18050 ( \18427 , \18426 , \18109 );
xor \U$18051 ( \18428 , \18174 , \18181 );
xor \U$18052 ( \18429 , \18428 , \18189 );
and \U$18053 ( \18430 , \18427 , \18429 );
and \U$18054 ( \18431 , \18422 , \18427 );
or \U$18055 ( \18432 , \18425 , \18430 , \18431 );
and \U$18056 ( \18433 , \18420 , \18432 );
and \U$18057 ( \18434 , \18383 , \18419 );
or \U$18058 ( \18435 , \18433 , \18434 );
and \U$18059 ( \18436 , \5896 , RIae78698_115);
and \U$18060 ( \18437 , RIae75b78_23, \5894 );
nor \U$18061 ( \18438 , \18436 , \18437 );
and \U$18062 ( \18439 , \18438 , \5589 );
not \U$18063 ( \18440 , \18438 );
and \U$18064 ( \18441 , \18440 , \5590 );
nor \U$18065 ( \18442 , \18439 , \18441 );
not \U$18066 ( \18443 , \18442 );
and \U$18067 ( \18444 , \6941 , RIae758a8_17);
and \U$18068 ( \18445 , RIae75f38_31, \6939 );
nor \U$18069 ( \18446 , \18444 , \18445 );
and \U$18070 ( \18447 , \18446 , \6945 );
not \U$18071 ( \18448 , \18446 );
and \U$18072 ( \18449 , \18448 , \6314 );
nor \U$18073 ( \18450 , \18447 , \18449 );
not \U$18074 ( \18451 , \18450 );
and \U$18075 ( \18452 , \18443 , \18451 );
and \U$18076 ( \18453 , \18450 , \18442 );
and \U$18077 ( \18454 , \6172 , RIae75a88_21);
and \U$18078 ( \18455 , RIae75998_19, \6170 );
nor \U$18079 ( \18456 , \18454 , \18455 );
and \U$18080 ( \18457 , \18456 , \6175 );
not \U$18081 ( \18458 , \18456 );
and \U$18082 ( \18459 , \18458 , \6176 );
nor \U$18083 ( \18460 , \18457 , \18459 );
nor \U$18084 ( \18461 , \18453 , \18460 );
nor \U$18085 ( \18462 , \18452 , \18461 );
and \U$18086 ( \18463 , \7633 , RIae75e48_29);
and \U$18087 ( \18464 , RIae75c68_25, \7631 );
nor \U$18088 ( \18465 , \18463 , \18464 );
and \U$18089 ( \18466 , \18465 , \7205 );
not \U$18090 ( \18467 , \18465 );
and \U$18091 ( \18468 , \18467 , \7206 );
nor \U$18092 ( \18469 , \18466 , \18468 );
not \U$18093 ( \18470 , \18469 );
and \U$18094 ( \18471 , \8966 , RIae754e8_9);
and \U$18095 ( \18472 , RIae757b8_15, \8964 );
nor \U$18096 ( \18473 , \18471 , \18472 );
and \U$18097 ( \18474 , \18473 , \8789 );
not \U$18098 ( \18475 , \18473 );
and \U$18099 ( \18476 , \18475 , \8799 );
nor \U$18100 ( \18477 , \18474 , \18476 );
not \U$18101 ( \18478 , \18477 );
and \U$18102 ( \18479 , \18470 , \18478 );
and \U$18103 ( \18480 , \18477 , \18469 );
and \U$18104 ( \18481 , \8371 , RIae75d58_27);
and \U$18105 ( \18482 , RIae755d8_11, \8369 );
nor \U$18106 ( \18483 , \18481 , \18482 );
and \U$18107 ( \18484 , \18483 , \8019 );
not \U$18108 ( \18485 , \18483 );
and \U$18109 ( \18486 , \18485 , \8020 );
nor \U$18110 ( \18487 , \18484 , \18486 );
nor \U$18111 ( \18488 , \18480 , \18487 );
nor \U$18112 ( \18489 , \18479 , \18488 );
or \U$18113 ( \18490 , \18462 , \18489 );
not \U$18114 ( \18491 , \18462 );
not \U$18115 ( \18492 , \18489 );
or \U$18116 ( \18493 , \18491 , \18492 );
and \U$18117 ( \18494 , \4688 , RIae77e28_97);
and \U$18118 ( \18495 , RIae78968_121, \4686 );
nor \U$18119 ( \18496 , \18494 , \18495 );
and \U$18120 ( \18497 , \18496 , \4481 );
not \U$18121 ( \18498 , \18496 );
and \U$18122 ( \18499 , \18498 , \4482 );
nor \U$18123 ( \18500 , \18497 , \18499 );
and \U$18124 ( \18501 , \4247 , RIae77b58_91);
and \U$18125 ( \18502 , RIae77d38_95, \4245 );
nor \U$18126 ( \18503 , \18501 , \18502 );
and \U$18127 ( \18504 , \18503 , \3989 );
not \U$18128 ( \18505 , \18503 );
and \U$18129 ( \18506 , \18505 , \4251 );
nor \U$18130 ( \18507 , \18504 , \18506 );
xor \U$18131 ( \18508 , \18500 , \18507 );
and \U$18132 ( \18509 , \5399 , RIae78878_119);
and \U$18133 ( \18510 , RIae78788_117, \5397 );
nor \U$18134 ( \18511 , \18509 , \18510 );
and \U$18135 ( \18512 , \18511 , \5016 );
not \U$18136 ( \18513 , \18511 );
and \U$18137 ( \18514 , \18513 , \5403 );
nor \U$18138 ( \18515 , \18512 , \18514 );
and \U$18139 ( \18516 , \18508 , \18515 );
and \U$18140 ( \18517 , \18500 , \18507 );
or \U$18141 ( \18518 , \18516 , \18517 );
nand \U$18142 ( \18519 , \18493 , \18518 );
nand \U$18143 ( \18520 , \18490 , \18519 );
and \U$18144 ( \18521 , \9760 , RIae756c8_13);
and \U$18145 ( \18522 , RIae75218_3, \9758 );
nor \U$18146 ( \18523 , \18521 , \18522 );
and \U$18147 ( \18524 , \18523 , \9273 );
not \U$18148 ( \18525 , \18523 );
and \U$18149 ( \18526 , \18525 , \9764 );
nor \U$18150 ( \18527 , \18524 , \18526 );
and \U$18151 ( \18528 , \10548 , RIae75128_1);
and \U$18152 ( \18529 , RIae75308_5, \10546 );
nor \U$18153 ( \18530 , \18528 , \18529 );
and \U$18154 ( \18531 , \18530 , \10421 );
not \U$18155 ( \18532 , \18530 );
and \U$18156 ( \18533 , \18532 , \10118 );
nor \U$18157 ( \18534 , \18531 , \18533 );
xor \U$18158 ( \18535 , \18527 , \18534 );
and \U$18159 ( \18536 , \11470 , RIae753f8_7);
and \U$18160 ( \18537 , RIae763e8_41, \11468 );
nor \U$18161 ( \18538 , \18536 , \18537 );
and \U$18162 ( \18539 , \18538 , \10936 );
not \U$18163 ( \18540 , \18538 );
and \U$18164 ( \18541 , \18540 , \11474 );
nor \U$18165 ( \18542 , \18539 , \18541 );
and \U$18166 ( \18543 , \18535 , \18542 );
and \U$18167 ( \18544 , \18527 , \18534 );
or \U$18168 ( \18545 , \18543 , \18544 );
and \U$18169 ( \18546 , \15726 , RIae76988_53);
and \U$18170 ( \18547 , RIae7aab0_192, RIae767a8_49);
nor \U$18171 ( \18548 , \18546 , \18547 );
and \U$18172 ( \18549 , \18548 , \14959 );
not \U$18173 ( \18550 , \18548 );
and \U$18174 ( \18551 , \18550 , RIae7aa38_191);
nor \U$18175 ( \18552 , \18549 , \18551 );
xor \U$18176 ( \18553 , \18552 , \471 );
and \U$18177 ( \18554 , \14964 , RIae76208_37);
and \U$18178 ( \18555 , RIae76a78_55, \14962 );
nor \U$18179 ( \18556 , \18554 , \18555 );
and \U$18180 ( \18557 , \18556 , \14463 );
not \U$18181 ( \18558 , \18556 );
and \U$18182 ( \18559 , \18558 , \14462 );
nor \U$18183 ( \18560 , \18557 , \18559 );
and \U$18184 ( \18561 , \18553 , \18560 );
and \U$18185 ( \18562 , \18552 , \471 );
or \U$18186 ( \18563 , \18561 , \18562 );
xor \U$18187 ( \18564 , \18545 , \18563 );
and \U$18188 ( \18565 , \12180 , RIae764d8_43);
and \U$18189 ( \18566 , RIae766b8_47, \12178 );
nor \U$18190 ( \18567 , \18565 , \18566 );
and \U$18191 ( \18568 , \18567 , \12184 );
not \U$18192 ( \18569 , \18567 );
and \U$18193 ( \18570 , \18569 , \11827 );
nor \U$18194 ( \18571 , \18568 , \18570 );
and \U$18195 ( \18572 , \13059 , RIae765c8_45);
and \U$18196 ( \18573 , RIae76118_35, \13057 );
nor \U$18197 ( \18574 , \18572 , \18573 );
and \U$18198 ( \18575 , \18574 , \13063 );
not \U$18199 ( \18576 , \18574 );
and \U$18200 ( \18577 , \18576 , \12718 );
nor \U$18201 ( \18578 , \18575 , \18577 );
xor \U$18202 ( \18579 , \18571 , \18578 );
and \U$18203 ( \18580 , \14059 , RIae76028_33);
and \U$18204 ( \18581 , RIae762f8_39, \14057 );
nor \U$18205 ( \18582 , \18580 , \18581 );
and \U$18206 ( \18583 , \18582 , \13502 );
not \U$18207 ( \18584 , \18582 );
and \U$18208 ( \18585 , \18584 , \14063 );
nor \U$18209 ( \18586 , \18583 , \18585 );
and \U$18210 ( \18587 , \18579 , \18586 );
and \U$18211 ( \18588 , \18571 , \18578 );
or \U$18212 ( \18589 , \18587 , \18588 );
and \U$18213 ( \18590 , \18564 , \18589 );
and \U$18214 ( \18591 , \18545 , \18563 );
or \U$18215 ( \18592 , \18590 , \18591 );
xor \U$18216 ( \18593 , \18520 , \18592 );
and \U$18217 ( \18594 , \2224 , RIae772e8_73);
and \U$18218 ( \18595 , RIae782d8_107, \2222 );
nor \U$18219 ( \18596 , \18594 , \18595 );
and \U$18220 ( \18597 , \18596 , \2061 );
not \U$18221 ( \18598 , \18596 );
and \U$18222 ( \18599 , \18598 , \2060 );
nor \U$18223 ( \18600 , \18597 , \18599 );
and \U$18224 ( \18601 , \1939 , RIae77018_67);
and \U$18225 ( \18602 , RIae771f8_71, \1937 );
nor \U$18226 ( \18603 , \18601 , \18602 );
and \U$18227 ( \18604 , \18603 , \1735 );
not \U$18228 ( \18605 , \18603 );
and \U$18229 ( \18606 , \18605 , \1734 );
nor \U$18230 ( \18607 , \18604 , \18606 );
xor \U$18231 ( \18608 , \18600 , \18607 );
and \U$18232 ( \18609 , \2607 , RIae780f8_103);
and \U$18233 ( \18610 , RIae77f18_99, \2605 );
nor \U$18234 ( \18611 , \18609 , \18610 );
and \U$18235 ( \18612 , \18611 , \2611 );
not \U$18236 ( \18613 , \18611 );
and \U$18237 ( \18614 , \18613 , \2397 );
nor \U$18238 ( \18615 , \18612 , \18614 );
and \U$18239 ( \18616 , \18608 , \18615 );
and \U$18240 ( \18617 , \18600 , \18607 );
or \U$18241 ( \18618 , \18616 , \18617 );
and \U$18242 ( \18619 , \1138 , RIae77888_85);
and \U$18243 ( \18620 , RIae76f28_65, \1136 );
nor \U$18244 ( \18621 , \18619 , \18620 );
and \U$18245 ( \18622 , \18621 , \1012 );
not \U$18246 ( \18623 , \18621 );
and \U$18247 ( \18624 , \18623 , \1142 );
nor \U$18248 ( \18625 , \18622 , \18624 );
and \U$18249 ( \18626 , \1376 , RIae76e38_63);
and \U$18250 ( \18627 , RIae76d48_61, \1374 );
nor \U$18251 ( \18628 , \18626 , \18627 );
and \U$18252 ( \18629 , \18628 , \1380 );
not \U$18253 ( \18630 , \18628 );
and \U$18254 ( \18631 , \18630 , \1261 );
nor \U$18255 ( \18632 , \18629 , \18631 );
xor \U$18256 ( \18633 , \18625 , \18632 );
and \U$18257 ( \18634 , \1593 , RIae76c58_59);
and \U$18258 ( \18635 , RIae77180_70, \1591 );
nor \U$18259 ( \18636 , \18634 , \18635 );
and \U$18260 ( \18637 , \18636 , \1498 );
not \U$18261 ( \18638 , \18636 );
and \U$18262 ( \18639 , \18638 , \1488 );
nor \U$18263 ( \18640 , \18637 , \18639 );
and \U$18264 ( \18641 , \18633 , \18640 );
and \U$18265 ( \18642 , \18625 , \18632 );
or \U$18266 ( \18643 , \18641 , \18642 );
xor \U$18267 ( \18644 , \18618 , \18643 );
not \U$18268 ( \18645 , \3218 );
and \U$18269 ( \18646 , \3214 , RIae785a8_113);
and \U$18270 ( \18647 , RIae783c8_109, \3212 );
nor \U$18271 ( \18648 , \18646 , \18647 );
not \U$18272 ( \18649 , \18648 );
or \U$18273 ( \18650 , \18645 , \18649 );
or \U$18274 ( \18651 , \18648 , \3218 );
nand \U$18275 ( \18652 , \18650 , \18651 );
not \U$18276 ( \18653 , \2789 );
and \U$18277 ( \18654 , \2783 , RIae78008_101);
and \U$18278 ( \18655 , RIae781e8_105, \2781 );
nor \U$18279 ( \18656 , \18654 , \18655 );
not \U$18280 ( \18657 , \18656 );
or \U$18281 ( \18658 , \18653 , \18657 );
or \U$18282 ( \18659 , \18656 , \3089 );
nand \U$18283 ( \18660 , \18658 , \18659 );
xor \U$18284 ( \18661 , \18652 , \18660 );
and \U$18285 ( \18662 , \3730 , RIae78530_112);
and \U$18286 ( \18663 , RIae77c48_93, \3728 );
nor \U$18287 ( \18664 , \18662 , \18663 );
and \U$18288 ( \18665 , \18664 , \3732 );
not \U$18289 ( \18666 , \18664 );
and \U$18290 ( \18667 , \18666 , \3422 );
nor \U$18291 ( \18668 , \18665 , \18667 );
and \U$18292 ( \18669 , \18661 , \18668 );
and \U$18293 ( \18670 , \18652 , \18660 );
or \U$18294 ( \18671 , \18669 , \18670 );
and \U$18295 ( \18672 , \18644 , \18671 );
and \U$18296 ( \18673 , \18618 , \18643 );
or \U$18297 ( \18674 , \18672 , \18673 );
and \U$18298 ( \18675 , \18593 , \18674 );
and \U$18299 ( \18676 , \18520 , \18592 );
or \U$18300 ( \18677 , \18675 , \18676 );
xor \U$18301 ( \18678 , \18435 , \18677 );
xor \U$18302 ( \18679 , \17725 , \17732 );
xor \U$18303 ( \18680 , \18679 , \17740 );
xor \U$18304 ( \18681 , \18296 , \18301 );
xor \U$18305 ( \18682 , \18680 , \18681 );
xor \U$18306 ( \18683 , \18252 , \18254 );
xor \U$18307 ( \18684 , \18683 , \18257 );
and \U$18308 ( \18685 , \18682 , \18684 );
xor \U$18309 ( \18686 , \17645 , \17652 );
xor \U$18310 ( \18687 , \18686 , \17660 );
xor \U$18311 ( \18688 , \17985 , \17990 );
xor \U$18312 ( \18689 , \18687 , \18688 );
xor \U$18313 ( \18690 , \18252 , \18254 );
xor \U$18314 ( \18691 , \18690 , \18257 );
and \U$18315 ( \18692 , \18689 , \18691 );
and \U$18316 ( \18693 , \18682 , \18689 );
or \U$18317 ( \18694 , \18685 , \18692 , \18693 );
and \U$18318 ( \18695 , \18678 , \18694 );
and \U$18319 ( \18696 , \18435 , \18677 );
or \U$18320 ( \18697 , \18695 , \18696 );
xor \U$18321 ( \18698 , \18373 , \18697 );
xor \U$18322 ( \18699 , \17619 , \17637 );
xor \U$18323 ( \18700 , \18699 , \17663 );
xor \U$18324 ( \18701 , \17953 , \17958 );
xor \U$18325 ( \18702 , \18700 , \18701 );
xor \U$18326 ( \18703 , \18030 , \18056 );
xor \U$18327 ( \18704 , \18703 , \18084 );
xor \U$18328 ( \18705 , \18192 , \18217 );
xor \U$18329 ( \18706 , \18705 , \18243 );
and \U$18330 ( \18707 , \18704 , \18706 );
xor \U$18331 ( \18708 , \18286 , \18287 );
xor \U$18332 ( \18709 , \18708 , \18290 );
xor \U$18333 ( \18710 , \18192 , \18217 );
xor \U$18334 ( \18711 , \18710 , \18243 );
and \U$18335 ( \18712 , \18709 , \18711 );
and \U$18336 ( \18713 , \18704 , \18709 );
or \U$18337 ( \18714 , \18707 , \18712 , \18713 );
xor \U$18338 ( \18715 , \18702 , \18714 );
xor \U$18339 ( \18716 , \17502 , \17504 );
xor \U$18340 ( \18717 , \18716 , \17507 );
xor \U$18341 ( \18718 , \17968 , \17975 );
xor \U$18342 ( \18719 , \18717 , \18718 );
and \U$18343 ( \18720 , \18715 , \18719 );
and \U$18344 ( \18721 , \18702 , \18714 );
or \U$18345 ( \18722 , \18720 , \18721 );
and \U$18346 ( \18723 , \18698 , \18722 );
and \U$18347 ( \18724 , \18373 , \18697 );
or \U$18348 ( \18725 , \18723 , \18724 );
xor \U$18349 ( \18726 , \17446 , \17499 );
xor \U$18350 ( \18727 , \18726 , \17510 );
xor \U$18351 ( \18728 , \17594 , \17666 );
xor \U$18352 ( \18729 , \18728 , \17746 );
xor \U$18353 ( \18730 , \18727 , \18729 );
xor \U$18354 ( \18731 , \17782 , \17784 );
xor \U$18355 ( \18732 , \18731 , \17789 );
xor \U$18356 ( \18733 , \18315 , \18322 );
xor \U$18357 ( \18734 , \18732 , \18733 );
and \U$18358 ( \18735 , \18730 , \18734 );
and \U$18359 ( \18736 , \18727 , \18729 );
or \U$18360 ( \18737 , \18735 , \18736 );
xor \U$18361 ( \18738 , \18725 , \18737 );
xor \U$18362 ( \18739 , \17169 , \17411 );
xor \U$18363 ( \18740 , \18739 , \17431 );
xor \U$18364 ( \18741 , \18335 , \18342 );
xor \U$18365 ( \18742 , \18740 , \18741 );
and \U$18366 ( \18743 , \18738 , \18742 );
and \U$18367 ( \18744 , \18725 , \18737 );
or \U$18368 ( \18745 , \18743 , \18744 );
xor \U$18369 ( \18746 , \18330 , \18332 );
xor \U$18370 ( \18747 , \18746 , \18347 );
and \U$18371 ( \18748 , \18745 , \18747 );
xor \U$18372 ( \18749 , \17940 , \17942 );
xor \U$18373 ( \18750 , \18749 , \17945 );
xor \U$18374 ( \18751 , \18330 , \18332 );
xor \U$18375 ( \18752 , \18751 , \18347 );
and \U$18376 ( \18753 , \18750 , \18752 );
and \U$18377 ( \18754 , \18745 , \18750 );
or \U$18378 ( \18755 , \18748 , \18753 , \18754 );
not \U$18379 ( \18756 , \17932 );
not \U$18380 ( \18757 , \17925 );
or \U$18381 ( \18758 , \18756 , \18757 );
or \U$18382 ( \18759 , \17925 , \17932 );
nand \U$18383 ( \18760 , \18758 , \18759 );
xor \U$18384 ( \18761 , \18755 , \18760 );
xor \U$18385 ( \18762 , \17948 , \17950 );
xor \U$18386 ( \18763 , \18762 , \18350 );
and \U$18387 ( \18764 , \18761 , \18763 );
and \U$18388 ( \18765 , \18755 , \18760 );
or \U$18389 ( \18766 , \18764 , \18765 );
and \U$18390 ( \18767 , \18361 , \18766 );
xor \U$18391 ( \18768 , \18766 , \18361 );
xor \U$18392 ( \18769 , \18755 , \18760 );
xor \U$18393 ( \18770 , \18769 , \18763 );
not \U$18394 ( \18771 , \18770 );
xor \U$18395 ( \18772 , \17983 , \18312 );
xor \U$18396 ( \18773 , \18772 , \18327 );
xor \U$18397 ( \18774 , \18005 , \18249 );
xor \U$18398 ( \18775 , \18774 , \18309 );
xor \U$18399 ( \18776 , \18727 , \18729 );
xor \U$18400 ( \18777 , \18776 , \18734 );
and \U$18401 ( \18778 , \18775 , \18777 );
xor \U$18402 ( \18779 , \18373 , \18697 );
xor \U$18403 ( \18780 , \18779 , \18722 );
xor \U$18404 ( \18781 , \18727 , \18729 );
xor \U$18405 ( \18782 , \18781 , \18734 );
and \U$18406 ( \18783 , \18780 , \18782 );
and \U$18407 ( \18784 , \18775 , \18780 );
or \U$18408 ( \18785 , \18778 , \18783 , \18784 );
xor \U$18409 ( \18786 , \18773 , \18785 );
xor \U$18410 ( \18787 , \18520 , \18592 );
xor \U$18411 ( \18788 , \18787 , \18674 );
xor \U$18412 ( \18789 , \18383 , \18419 );
xor \U$18413 ( \18790 , \18789 , \18432 );
and \U$18414 ( \18791 , \18788 , \18790 );
xor \U$18415 ( \18792 , \18252 , \18254 );
xor \U$18416 ( \18793 , \18792 , \18257 );
xor \U$18417 ( \18794 , \18682 , \18689 );
xor \U$18418 ( \18795 , \18793 , \18794 );
xor \U$18419 ( \18796 , \18383 , \18419 );
xor \U$18420 ( \18797 , \18796 , \18432 );
and \U$18421 ( \18798 , \18795 , \18797 );
and \U$18422 ( \18799 , \18788 , \18795 );
or \U$18423 ( \18800 , \18791 , \18798 , \18799 );
xor \U$18424 ( \18801 , \18145 , \18152 );
xor \U$18425 ( \18802 , \18801 , \18160 );
xor \U$18426 ( \18803 , \18119 , \18126 );
xor \U$18427 ( \18804 , \18803 , \18134 );
xor \U$18428 ( \18805 , \18802 , \18804 );
xor \U$18429 ( \18806 , \18174 , \18181 );
xor \U$18430 ( \18807 , \18806 , \18189 );
xor \U$18431 ( \18808 , \18422 , \18427 );
xor \U$18432 ( \18809 , \18807 , \18808 );
and \U$18433 ( \18810 , \18805 , \18809 );
and \U$18434 ( \18811 , \18802 , \18804 );
or \U$18435 ( \18812 , \18810 , \18811 );
and \U$18436 ( \18813 , \1138 , RIae77798_83);
and \U$18437 ( \18814 , RIae77888_85, \1136 );
nor \U$18438 ( \18815 , \18813 , \18814 );
and \U$18439 ( \18816 , \18815 , \1012 );
not \U$18440 ( \18817 , \18815 );
and \U$18441 ( \18818 , \18817 , \1142 );
nor \U$18442 ( \18819 , \18816 , \18818 );
and \U$18443 ( \18820 , \1376 , RIae76f28_65);
and \U$18444 ( \18821 , RIae76e38_63, \1374 );
nor \U$18445 ( \18822 , \18820 , \18821 );
and \U$18446 ( \18823 , \18822 , \1380 );
not \U$18447 ( \18824 , \18822 );
and \U$18448 ( \18825 , \18824 , \1261 );
nor \U$18449 ( \18826 , \18823 , \18825 );
xor \U$18450 ( \18827 , \18819 , \18826 );
not \U$18451 ( \18828 , \789 );
and \U$18452 ( \18829 , \883 , RIae77a68_89);
and \U$18453 ( \18830 , RIae77978_87, \881 );
nor \U$18454 ( \18831 , \18829 , \18830 );
not \U$18455 ( \18832 , \18831 );
or \U$18456 ( \18833 , \18828 , \18832 );
or \U$18457 ( \18834 , \18831 , \787 );
nand \U$18458 ( \18835 , \18833 , \18834 );
and \U$18459 ( \18836 , \18827 , \18835 );
and \U$18460 ( \18837 , \18819 , \18826 );
nor \U$18461 ( \18838 , \18836 , \18837 );
and \U$18462 ( \18839 , \1939 , RIae77180_70);
and \U$18463 ( \18840 , RIae77018_67, \1937 );
nor \U$18464 ( \18841 , \18839 , \18840 );
and \U$18465 ( \18842 , \18841 , \1735 );
not \U$18466 ( \18843 , \18841 );
and \U$18467 ( \18844 , \18843 , \1734 );
nor \U$18468 ( \18845 , \18842 , \18844 );
and \U$18469 ( \18846 , \2224 , RIae771f8_71);
and \U$18470 ( \18847 , RIae772e8_73, \2222 );
nor \U$18471 ( \18848 , \18846 , \18847 );
and \U$18472 ( \18849 , \18848 , \2061 );
not \U$18473 ( \18850 , \18848 );
and \U$18474 ( \18851 , \18850 , \2060 );
nor \U$18475 ( \18852 , \18849 , \18851 );
xor \U$18476 ( \18853 , \18845 , \18852 );
and \U$18477 ( \18854 , \1593 , RIae76d48_61);
and \U$18478 ( \18855 , RIae76c58_59, \1591 );
nor \U$18479 ( \18856 , \18854 , \18855 );
and \U$18480 ( \18857 , \18856 , \1498 );
not \U$18481 ( \18858 , \18856 );
and \U$18482 ( \18859 , \18858 , \1488 );
nor \U$18483 ( \18860 , \18857 , \18859 );
and \U$18484 ( \18861 , \18853 , \18860 );
and \U$18485 ( \18862 , \18845 , \18852 );
nor \U$18486 ( \18863 , \18861 , \18862 );
xor \U$18487 ( \18864 , \18838 , \18863 );
and \U$18488 ( \18865 , \2607 , RIae782d8_107);
and \U$18489 ( \18866 , RIae780f8_103, \2605 );
nor \U$18490 ( \18867 , \18865 , \18866 );
and \U$18491 ( \18868 , \18867 , \2397 );
not \U$18492 ( \18869 , \18867 );
and \U$18493 ( \18870 , \18869 , \2611 );
nor \U$18494 ( \18871 , \18868 , \18870 );
not \U$18495 ( \18872 , \18871 );
and \U$18496 ( \18873 , \3214 , RIae781e8_105);
and \U$18497 ( \18874 , RIae785a8_113, \3212 );
nor \U$18498 ( \18875 , \18873 , \18874 );
not \U$18499 ( \18876 , \18875 );
not \U$18500 ( \18877 , \3218 );
and \U$18501 ( \18878 , \18876 , \18877 );
and \U$18502 ( \18879 , \18875 , \3218 );
nor \U$18503 ( \18880 , \18878 , \18879 );
not \U$18504 ( \18881 , \18880 );
and \U$18505 ( \18882 , \18872 , \18881 );
and \U$18506 ( \18883 , \18880 , \18871 );
and \U$18507 ( \18884 , \2783 , RIae77f18_99);
and \U$18508 ( \18885 , RIae78008_101, \2781 );
nor \U$18509 ( \18886 , \18884 , \18885 );
not \U$18510 ( \18887 , \18886 );
not \U$18511 ( \18888 , \2789 );
and \U$18512 ( \18889 , \18887 , \18888 );
and \U$18513 ( \18890 , \18886 , \3089 );
nor \U$18514 ( \18891 , \18889 , \18890 );
nor \U$18515 ( \18892 , \18883 , \18891 );
nor \U$18516 ( \18893 , \18882 , \18892 );
and \U$18517 ( \18894 , \18864 , \18893 );
and \U$18518 ( \18895 , \18838 , \18863 );
nor \U$18519 ( \18896 , \18894 , \18895 );
and \U$18520 ( \18897 , \9760 , RIae757b8_15);
and \U$18521 ( \18898 , RIae756c8_13, \9758 );
nor \U$18522 ( \18899 , \18897 , \18898 );
and \U$18523 ( \18900 , \18899 , \9273 );
not \U$18524 ( \18901 , \18899 );
and \U$18525 ( \18902 , \18901 , \9764 );
nor \U$18526 ( \18903 , \18900 , \18902 );
and \U$18527 ( \18904 , \10548 , RIae75218_3);
and \U$18528 ( \18905 , RIae75128_1, \10546 );
nor \U$18529 ( \18906 , \18904 , \18905 );
and \U$18530 ( \18907 , \18906 , \10421 );
not \U$18531 ( \18908 , \18906 );
and \U$18532 ( \18909 , \18908 , \10118 );
nor \U$18533 ( \18910 , \18907 , \18909 );
xor \U$18534 ( \18911 , \18903 , \18910 );
and \U$18535 ( \18912 , \8966 , RIae755d8_11);
and \U$18536 ( \18913 , RIae754e8_9, \8964 );
nor \U$18537 ( \18914 , \18912 , \18913 );
and \U$18538 ( \18915 , \18914 , \8799 );
not \U$18539 ( \18916 , \18914 );
and \U$18540 ( \18917 , \18916 , \8789 );
nor \U$18541 ( \18918 , \18915 , \18917 );
and \U$18542 ( \18919 , \18911 , \18918 );
and \U$18543 ( \18920 , \18903 , \18910 );
nor \U$18544 ( \18921 , \18919 , \18920 );
and \U$18545 ( \18922 , \14964 , RIae762f8_39);
and \U$18546 ( \18923 , RIae76208_37, \14962 );
nor \U$18547 ( \18924 , \18922 , \18923 );
and \U$18548 ( \18925 , \18924 , \14463 );
not \U$18549 ( \18926 , \18924 );
and \U$18550 ( \18927 , \18926 , \14462 );
nor \U$18551 ( \18928 , \18925 , \18927 );
and \U$18552 ( \18929 , \15726 , RIae76a78_55);
and \U$18553 ( \18930 , RIae7aab0_192, RIae76988_53);
nor \U$18554 ( \18931 , \18929 , \18930 );
and \U$18555 ( \18932 , \18931 , \14959 );
not \U$18556 ( \18933 , \18931 );
and \U$18557 ( \18934 , \18933 , RIae7aa38_191);
nor \U$18558 ( \18935 , \18932 , \18934 );
xor \U$18559 ( \18936 , \18928 , \18935 );
and \U$18560 ( \18937 , \14059 , RIae76118_35);
and \U$18561 ( \18938 , RIae76028_33, \14057 );
nor \U$18562 ( \18939 , \18937 , \18938 );
and \U$18563 ( \18940 , \18939 , \13502 );
not \U$18564 ( \18941 , \18939 );
and \U$18565 ( \18942 , \18941 , \14063 );
nor \U$18566 ( \18943 , \18940 , \18942 );
and \U$18567 ( \18944 , \18936 , \18943 );
and \U$18568 ( \18945 , \18928 , \18935 );
nor \U$18569 ( \18946 , \18944 , \18945 );
or \U$18570 ( \18947 , \18921 , \18946 );
not \U$18571 ( \18948 , \18946 );
not \U$18572 ( \18949 , \18921 );
or \U$18573 ( \18950 , \18948 , \18949 );
and \U$18574 ( \18951 , \13059 , RIae766b8_47);
and \U$18575 ( \18952 , RIae765c8_45, \13057 );
nor \U$18576 ( \18953 , \18951 , \18952 );
and \U$18577 ( \18954 , \18953 , \13063 );
not \U$18578 ( \18955 , \18953 );
and \U$18579 ( \18956 , \18955 , \12718 );
nor \U$18580 ( \18957 , \18954 , \18956 );
and \U$18581 ( \18958 , \11470 , RIae75308_5);
and \U$18582 ( \18959 , RIae753f8_7, \11468 );
nor \U$18583 ( \18960 , \18958 , \18959 );
and \U$18584 ( \18961 , \18960 , \10936 );
not \U$18585 ( \18962 , \18960 );
and \U$18586 ( \18963 , \18962 , \11474 );
nor \U$18587 ( \18964 , \18961 , \18963 );
xor \U$18588 ( \18965 , \18957 , \18964 );
and \U$18589 ( \18966 , \12180 , RIae763e8_41);
and \U$18590 ( \18967 , RIae764d8_43, \12178 );
nor \U$18591 ( \18968 , \18966 , \18967 );
and \U$18592 ( \18969 , \18968 , \12184 );
not \U$18593 ( \18970 , \18968 );
and \U$18594 ( \18971 , \18970 , \11827 );
nor \U$18595 ( \18972 , \18969 , \18971 );
and \U$18596 ( \18973 , \18965 , \18972 );
and \U$18597 ( \18974 , \18957 , \18964 );
or \U$18598 ( \18975 , \18973 , \18974 );
nand \U$18599 ( \18976 , \18950 , \18975 );
nand \U$18600 ( \18977 , \18947 , \18976 );
xor \U$18601 ( \18978 , \18896 , \18977 );
and \U$18602 ( \18979 , \5896 , RIae78788_117);
and \U$18603 ( \18980 , RIae78698_115, \5894 );
nor \U$18604 ( \18981 , \18979 , \18980 );
and \U$18605 ( \18982 , \18981 , \5590 );
not \U$18606 ( \18983 , \18981 );
and \U$18607 ( \18984 , \18983 , \5589 );
nor \U$18608 ( \18985 , \18982 , \18984 );
and \U$18609 ( \18986 , \6172 , RIae75b78_23);
and \U$18610 ( \18987 , RIae75a88_21, \6170 );
nor \U$18611 ( \18988 , \18986 , \18987 );
and \U$18612 ( \18989 , \18988 , \6176 );
not \U$18613 ( \18990 , \18988 );
and \U$18614 ( \18991 , \18990 , \6175 );
nor \U$18615 ( \18992 , \18989 , \18991 );
xor \U$18616 ( \18993 , \18985 , \18992 );
and \U$18617 ( \18994 , \5399 , RIae78968_121);
and \U$18618 ( \18995 , RIae78878_119, \5397 );
nor \U$18619 ( \18996 , \18994 , \18995 );
and \U$18620 ( \18997 , \18996 , \5016 );
not \U$18621 ( \18998 , \18996 );
and \U$18622 ( \18999 , \18998 , \5403 );
nor \U$18623 ( \19000 , \18997 , \18999 );
and \U$18624 ( \19001 , \18993 , \19000 );
and \U$18625 ( \19002 , \18985 , \18992 );
nor \U$18626 ( \19003 , \19001 , \19002 );
and \U$18627 ( \19004 , \7633 , RIae75f38_31);
and \U$18628 ( \19005 , RIae75e48_29, \7631 );
nor \U$18629 ( \19006 , \19004 , \19005 );
and \U$18630 ( \19007 , \19006 , \7206 );
not \U$18631 ( \19008 , \19006 );
and \U$18632 ( \19009 , \19008 , \7205 );
nor \U$18633 ( \19010 , \19007 , \19009 );
and \U$18634 ( \19011 , \8371 , RIae75c68_25);
and \U$18635 ( \19012 , RIae75d58_27, \8369 );
nor \U$18636 ( \19013 , \19011 , \19012 );
and \U$18637 ( \19014 , \19013 , \8020 );
not \U$18638 ( \19015 , \19013 );
and \U$18639 ( \19016 , \19015 , \8019 );
nor \U$18640 ( \19017 , \19014 , \19016 );
xor \U$18641 ( \19018 , \19010 , \19017 );
and \U$18642 ( \19019 , \6941 , RIae75998_19);
and \U$18643 ( \19020 , RIae758a8_17, \6939 );
nor \U$18644 ( \19021 , \19019 , \19020 );
and \U$18645 ( \19022 , \19021 , \6314 );
not \U$18646 ( \19023 , \19021 );
and \U$18647 ( \19024 , \19023 , \6945 );
nor \U$18648 ( \19025 , \19022 , \19024 );
and \U$18649 ( \19026 , \19018 , \19025 );
and \U$18650 ( \19027 , \19010 , \19017 );
nor \U$18651 ( \19028 , \19026 , \19027 );
or \U$18652 ( \19029 , \19003 , \19028 );
not \U$18653 ( \19030 , \19003 );
not \U$18654 ( \19031 , \19028 );
or \U$18655 ( \19032 , \19030 , \19031 );
and \U$18656 ( \19033 , \3730 , RIae783c8_109);
and \U$18657 ( \19034 , RIae78530_112, \3728 );
nor \U$18658 ( \19035 , \19033 , \19034 );
and \U$18659 ( \19036 , \19035 , \3732 );
not \U$18660 ( \19037 , \19035 );
and \U$18661 ( \19038 , \19037 , \3422 );
nor \U$18662 ( \19039 , \19036 , \19038 );
and \U$18663 ( \19040 , \4247 , RIae77c48_93);
and \U$18664 ( \19041 , RIae77b58_91, \4245 );
nor \U$18665 ( \19042 , \19040 , \19041 );
and \U$18666 ( \19043 , \19042 , \3989 );
not \U$18667 ( \19044 , \19042 );
and \U$18668 ( \19045 , \19044 , \4251 );
nor \U$18669 ( \19046 , \19043 , \19045 );
xor \U$18670 ( \19047 , \19039 , \19046 );
and \U$18671 ( \19048 , \4688 , RIae77d38_95);
and \U$18672 ( \19049 , RIae77e28_97, \4686 );
nor \U$18673 ( \19050 , \19048 , \19049 );
and \U$18674 ( \19051 , \19050 , \4481 );
not \U$18675 ( \19052 , \19050 );
and \U$18676 ( \19053 , \19052 , \4482 );
nor \U$18677 ( \19054 , \19051 , \19053 );
and \U$18678 ( \19055 , \19047 , \19054 );
and \U$18679 ( \19056 , \19039 , \19046 );
or \U$18680 ( \19057 , \19055 , \19056 );
nand \U$18681 ( \19058 , \19032 , \19057 );
nand \U$18682 ( \19059 , \19029 , \19058 );
and \U$18683 ( \19060 , \18978 , \19059 );
and \U$18684 ( \19061 , \18896 , \18977 );
or \U$18685 ( \19062 , \19060 , \19061 );
xor \U$18686 ( \19063 , \18812 , \19062 );
xor \U$18687 ( \19064 , \18652 , \18660 );
xor \U$18688 ( \19065 , \19064 , \18668 );
xor \U$18689 ( \19066 , \18600 , \18607 );
xor \U$18690 ( \19067 , \19066 , \18615 );
xor \U$18691 ( \19068 , \19065 , \19067 );
xor \U$18692 ( \19069 , \18500 , \18507 );
xor \U$18693 ( \19070 , \19069 , \18515 );
and \U$18694 ( \19071 , \19068 , \19070 );
and \U$18695 ( \19072 , \19065 , \19067 );
or \U$18696 ( \19073 , \19071 , \19072 );
nand \U$18697 ( \19074 , RIae775b8_79, \512 );
not \U$18698 ( \19075 , \19074 );
not \U$18699 ( \19076 , \469 );
or \U$18700 ( \19077 , \19075 , \19076 );
or \U$18701 ( \19078 , \469 , \19074 );
nand \U$18702 ( \19079 , \19077 , \19078 );
xor \U$18703 ( \19080 , \18390 , \18397 );
xor \U$18704 ( \19081 , \19080 , \18406 );
and \U$18705 ( \19082 , \19079 , \19081 );
xor \U$18706 ( \19083 , \18625 , \18632 );
xor \U$18707 ( \19084 , \19083 , \18640 );
xor \U$18708 ( \19085 , \18390 , \18397 );
xor \U$18709 ( \19086 , \19085 , \18406 );
and \U$18710 ( \19087 , \19084 , \19086 );
and \U$18711 ( \19088 , \19079 , \19084 );
or \U$18712 ( \19089 , \19082 , \19087 , \19088 );
xor \U$18713 ( \19090 , \19073 , \19089 );
not \U$18714 ( \19091 , \18442 );
xor \U$18715 ( \19092 , \18460 , \18450 );
not \U$18716 ( \19093 , \19092 );
or \U$18717 ( \19094 , \19091 , \19093 );
or \U$18718 ( \19095 , \19092 , \18442 );
nand \U$18719 ( \19096 , \19094 , \19095 );
not \U$18720 ( \19097 , \18469 );
xor \U$18721 ( \19098 , \18487 , \18477 );
not \U$18722 ( \19099 , \19098 );
or \U$18723 ( \19100 , \19097 , \19099 );
or \U$18724 ( \19101 , \19098 , \18469 );
nand \U$18725 ( \19102 , \19100 , \19101 );
xor \U$18726 ( \19103 , \19096 , \19102 );
xor \U$18727 ( \19104 , \18527 , \18534 );
xor \U$18728 ( \19105 , \19104 , \18542 );
and \U$18729 ( \19106 , \19103 , \19105 );
and \U$18730 ( \19107 , \19096 , \19102 );
or \U$18731 ( \19108 , \19106 , \19107 );
and \U$18732 ( \19109 , \19090 , \19108 );
and \U$18733 ( \19110 , \19073 , \19089 );
or \U$18734 ( \19111 , \19109 , \19110 );
and \U$18735 ( \19112 , \19063 , \19111 );
and \U$18736 ( \19113 , \18812 , \19062 );
or \U$18737 ( \19114 , \19112 , \19113 );
xor \U$18738 ( \19115 , \18800 , \19114 );
xor \U$18739 ( \19116 , \18618 , \18643 );
xor \U$18740 ( \19117 , \19116 , \18671 );
xor \U$18741 ( \19118 , \18375 , \18377 );
xor \U$18742 ( \19119 , \19118 , \18380 );
and \U$18743 ( \19120 , \19117 , \19119 );
xor \U$18744 ( \19121 , \18267 , \18275 );
xor \U$18745 ( \19122 , \19121 , \18283 );
xor \U$18746 ( \19123 , \18409 , \18414 );
xor \U$18747 ( \19124 , \19122 , \19123 );
xor \U$18748 ( \19125 , \18375 , \18377 );
xor \U$18749 ( \19126 , \19125 , \18380 );
and \U$18750 ( \19127 , \19124 , \19126 );
and \U$18751 ( \19128 , \19117 , \19124 );
or \U$18752 ( \19129 , \19120 , \19127 , \19128 );
xor \U$18753 ( \19130 , \18112 , \18137 );
xor \U$18754 ( \19131 , \19130 , \18163 );
xor \U$18755 ( \19132 , \19129 , \19131 );
xor \U$18756 ( \19133 , \18192 , \18217 );
xor \U$18757 ( \19134 , \19133 , \18243 );
xor \U$18758 ( \19135 , \18704 , \18709 );
xor \U$18759 ( \19136 , \19134 , \19135 );
and \U$18760 ( \19137 , \19132 , \19136 );
and \U$18761 ( \19138 , \19129 , \19131 );
or \U$18762 ( \19139 , \19137 , \19138 );
and \U$18763 ( \19140 , \19115 , \19139 );
and \U$18764 ( \19141 , \18800 , \19114 );
or \U$18765 ( \19142 , \19140 , \19141 );
xor \U$18766 ( \19143 , \17963 , \17965 );
xor \U$18767 ( \19144 , \19143 , \17980 );
xor \U$18768 ( \19145 , \19142 , \19144 );
xor \U$18769 ( \19146 , \18435 , \18677 );
xor \U$18770 ( \19147 , \19146 , \18694 );
xor \U$18771 ( \19148 , \18702 , \18714 );
xor \U$18772 ( \19149 , \19148 , \18719 );
and \U$18773 ( \19150 , \19147 , \19149 );
xor \U$18774 ( \19151 , \17995 , \17997 );
xor \U$18775 ( \19152 , \19151 , \18002 );
xor \U$18776 ( \19153 , \18363 , \18368 );
xor \U$18777 ( \19154 , \19152 , \19153 );
xor \U$18778 ( \19155 , \18702 , \18714 );
xor \U$18779 ( \19156 , \19155 , \18719 );
and \U$18780 ( \19157 , \19154 , \19156 );
and \U$18781 ( \19158 , \19147 , \19154 );
or \U$18782 ( \19159 , \19150 , \19157 , \19158 );
and \U$18783 ( \19160 , \19145 , \19159 );
and \U$18784 ( \19161 , \19142 , \19144 );
or \U$18785 ( \19162 , \19160 , \19161 );
and \U$18786 ( \19163 , \18786 , \19162 );
and \U$18787 ( \19164 , \18773 , \18785 );
nor \U$18788 ( \19165 , \19163 , \19164 );
not \U$18789 ( \19166 , \19165 );
xor \U$18790 ( \19167 , \18330 , \18332 );
xor \U$18791 ( \19168 , \19167 , \18347 );
xor \U$18792 ( \19169 , \18745 , \18750 );
xor \U$18793 ( \19170 , \19168 , \19169 );
nand \U$18794 ( \19171 , \19166 , \19170 );
or \U$18795 ( \19172 , \18771 , \19171 );
and \U$18796 ( \19173 , \19171 , \18770 );
not \U$18797 ( \19174 , \19171 );
and \U$18798 ( \19175 , \19174 , \18771 );
nor \U$18799 ( \19176 , \19173 , \19175 );
xor \U$18800 ( \19177 , \18812 , \19062 );
xor \U$18801 ( \19178 , \19177 , \19111 );
xor \U$18802 ( \19179 , \19129 , \19131 );
xor \U$18803 ( \19180 , \19179 , \19136 );
and \U$18804 ( \19181 , \19178 , \19180 );
xor \U$18805 ( \19182 , \18383 , \18419 );
xor \U$18806 ( \19183 , \19182 , \18432 );
xor \U$18807 ( \19184 , \18788 , \18795 );
xor \U$18808 ( \19185 , \19183 , \19184 );
xor \U$18809 ( \19186 , \19129 , \19131 );
xor \U$18810 ( \19187 , \19186 , \19136 );
and \U$18811 ( \19188 , \19185 , \19187 );
and \U$18812 ( \19189 , \19178 , \19185 );
or \U$18813 ( \19190 , \19181 , \19188 , \19189 );
xor \U$18814 ( \19191 , \18545 , \18563 );
xor \U$18815 ( \19192 , \19191 , \18589 );
xor \U$18816 ( \19193 , \18802 , \18804 );
xor \U$18817 ( \19194 , \19193 , \18809 );
and \U$18818 ( \19195 , \19192 , \19194 );
xor \U$18819 ( \19196 , \18375 , \18377 );
xor \U$18820 ( \19197 , \19196 , \18380 );
xor \U$18821 ( \19198 , \19117 , \19124 );
xor \U$18822 ( \19199 , \19197 , \19198 );
xor \U$18823 ( \19200 , \18802 , \18804 );
xor \U$18824 ( \19201 , \19200 , \18809 );
and \U$18825 ( \19202 , \19199 , \19201 );
and \U$18826 ( \19203 , \19192 , \19199 );
or \U$18827 ( \19204 , \19195 , \19202 , \19203 );
and \U$18828 ( \19205 , \2607 , RIae772e8_73);
and \U$18829 ( \19206 , RIae782d8_107, \2605 );
nor \U$18830 ( \19207 , \19205 , \19206 );
and \U$18831 ( \19208 , \19207 , \2611 );
not \U$18832 ( \19209 , \19207 );
and \U$18833 ( \19210 , \19209 , \2397 );
nor \U$18834 ( \19211 , \19208 , \19210 );
and \U$18835 ( \19212 , \1939 , RIae76c58_59);
and \U$18836 ( \19213 , RIae77180_70, \1937 );
nor \U$18837 ( \19214 , \19212 , \19213 );
and \U$18838 ( \19215 , \19214 , \1735 );
not \U$18839 ( \19216 , \19214 );
and \U$18840 ( \19217 , \19216 , \1734 );
nor \U$18841 ( \19218 , \19215 , \19217 );
xor \U$18842 ( \19219 , \19211 , \19218 );
and \U$18843 ( \19220 , \2224 , RIae77018_67);
and \U$18844 ( \19221 , RIae771f8_71, \2222 );
nor \U$18845 ( \19222 , \19220 , \19221 );
and \U$18846 ( \19223 , \19222 , \2061 );
not \U$18847 ( \19224 , \19222 );
and \U$18848 ( \19225 , \19224 , \2060 );
nor \U$18849 ( \19226 , \19223 , \19225 );
and \U$18850 ( \19227 , \19219 , \19226 );
and \U$18851 ( \19228 , \19211 , \19218 );
or \U$18852 ( \19229 , \19227 , \19228 );
and \U$18853 ( \19230 , \1376 , RIae77888_85);
and \U$18854 ( \19231 , RIae76f28_65, \1374 );
nor \U$18855 ( \19232 , \19230 , \19231 );
and \U$18856 ( \19233 , \19232 , \1261 );
not \U$18857 ( \19234 , \19232 );
and \U$18858 ( \19235 , \19234 , \1380 );
nor \U$18859 ( \19236 , \19233 , \19235 );
and \U$18860 ( \19237 , \1593 , RIae76e38_63);
and \U$18861 ( \19238 , RIae76d48_61, \1591 );
nor \U$18862 ( \19239 , \19237 , \19238 );
and \U$18863 ( \19240 , \19239 , \1488 );
not \U$18864 ( \19241 , \19239 );
and \U$18865 ( \19242 , \19241 , \1498 );
nor \U$18866 ( \19243 , \19240 , \19242 );
xor \U$18867 ( \19244 , \19236 , \19243 );
and \U$18868 ( \19245 , \1138 , RIae77978_87);
and \U$18869 ( \19246 , RIae77798_83, \1136 );
nor \U$18870 ( \19247 , \19245 , \19246 );
and \U$18871 ( \19248 , \19247 , \1142 );
not \U$18872 ( \19249 , \19247 );
and \U$18873 ( \19250 , \19249 , \1012 );
nor \U$18874 ( \19251 , \19248 , \19250 );
and \U$18875 ( \19252 , \19244 , \19251 );
and \U$18876 ( \19253 , \19236 , \19243 );
nor \U$18877 ( \19254 , \19252 , \19253 );
xor \U$18878 ( \19255 , \19229 , \19254 );
and \U$18879 ( \19256 , \3730 , RIae785a8_113);
and \U$18880 ( \19257 , RIae783c8_109, \3728 );
nor \U$18881 ( \19258 , \19256 , \19257 );
and \U$18882 ( \19259 , \19258 , \3732 );
not \U$18883 ( \19260 , \19258 );
and \U$18884 ( \19261 , \19260 , \3422 );
nor \U$18885 ( \19262 , \19259 , \19261 );
not \U$18886 ( \19263 , \3089 );
and \U$18887 ( \19264 , \2783 , RIae780f8_103);
and \U$18888 ( \19265 , RIae77f18_99, \2781 );
nor \U$18889 ( \19266 , \19264 , \19265 );
not \U$18890 ( \19267 , \19266 );
or \U$18891 ( \19268 , \19263 , \19267 );
or \U$18892 ( \19269 , \19266 , \2789 );
nand \U$18893 ( \19270 , \19268 , \19269 );
xor \U$18894 ( \19271 , \19262 , \19270 );
not \U$18895 ( \19272 , \2774 );
and \U$18896 ( \19273 , \3214 , RIae78008_101);
and \U$18897 ( \19274 , RIae781e8_105, \3212 );
nor \U$18898 ( \19275 , \19273 , \19274 );
not \U$18899 ( \19276 , \19275 );
or \U$18900 ( \19277 , \19272 , \19276 );
or \U$18901 ( \19278 , \19275 , \3218 );
nand \U$18902 ( \19279 , \19277 , \19278 );
and \U$18903 ( \19280 , \19271 , \19279 );
and \U$18904 ( \19281 , \19262 , \19270 );
or \U$18905 ( \19282 , \19280 , \19281 );
and \U$18906 ( \19283 , \19255 , \19282 );
and \U$18907 ( \19284 , \19229 , \19254 );
or \U$18908 ( \19285 , \19283 , \19284 );
and \U$18909 ( \19286 , \9760 , RIae754e8_9);
and \U$18910 ( \19287 , RIae757b8_15, \9758 );
nor \U$18911 ( \19288 , \19286 , \19287 );
and \U$18912 ( \19289 , \19288 , \9273 );
not \U$18913 ( \19290 , \19288 );
and \U$18914 ( \19291 , \19290 , \9764 );
nor \U$18915 ( \19292 , \19289 , \19291 );
and \U$18916 ( \19293 , \10548 , RIae756c8_13);
and \U$18917 ( \19294 , RIae75218_3, \10546 );
nor \U$18918 ( \19295 , \19293 , \19294 );
and \U$18919 ( \19296 , \19295 , \10421 );
not \U$18920 ( \19297 , \19295 );
and \U$18921 ( \19298 , \19297 , \10118 );
nor \U$18922 ( \19299 , \19296 , \19298 );
xor \U$18923 ( \19300 , \19292 , \19299 );
and \U$18924 ( \19301 , \11470 , RIae75128_1);
and \U$18925 ( \19302 , RIae75308_5, \11468 );
nor \U$18926 ( \19303 , \19301 , \19302 );
and \U$18927 ( \19304 , \19303 , \10936 );
not \U$18928 ( \19305 , \19303 );
and \U$18929 ( \19306 , \19305 , \11474 );
nor \U$18930 ( \19307 , \19304 , \19306 );
and \U$18931 ( \19308 , \19300 , \19307 );
and \U$18932 ( \19309 , \19292 , \19299 );
or \U$18933 ( \19310 , \19308 , \19309 );
and \U$18934 ( \19311 , \15726 , RIae76208_37);
and \U$18935 ( \19312 , RIae7aab0_192, RIae76a78_55);
nor \U$18936 ( \19313 , \19311 , \19312 );
and \U$18937 ( \19314 , \19313 , \14959 );
not \U$18938 ( \19315 , \19313 );
and \U$18939 ( \19316 , \19315 , RIae7aa38_191);
nor \U$18940 ( \19317 , \19314 , \19316 );
xor \U$18941 ( \19318 , \19317 , \562 );
and \U$18942 ( \19319 , \14964 , RIae76028_33);
and \U$18943 ( \19320 , RIae762f8_39, \14962 );
nor \U$18944 ( \19321 , \19319 , \19320 );
and \U$18945 ( \19322 , \19321 , \14463 );
not \U$18946 ( \19323 , \19321 );
and \U$18947 ( \19324 , \19323 , \14462 );
nor \U$18948 ( \19325 , \19322 , \19324 );
and \U$18949 ( \19326 , \19318 , \19325 );
and \U$18950 ( \19327 , \19317 , \562 );
or \U$18951 ( \19328 , \19326 , \19327 );
xor \U$18952 ( \19329 , \19310 , \19328 );
and \U$18953 ( \19330 , \13059 , RIae764d8_43);
and \U$18954 ( \19331 , RIae766b8_47, \13057 );
nor \U$18955 ( \19332 , \19330 , \19331 );
and \U$18956 ( \19333 , \19332 , \13063 );
not \U$18957 ( \19334 , \19332 );
and \U$18958 ( \19335 , \19334 , \12718 );
nor \U$18959 ( \19336 , \19333 , \19335 );
and \U$18960 ( \19337 , \12180 , RIae753f8_7);
and \U$18961 ( \19338 , RIae763e8_41, \12178 );
nor \U$18962 ( \19339 , \19337 , \19338 );
and \U$18963 ( \19340 , \19339 , \12184 );
not \U$18964 ( \19341 , \19339 );
and \U$18965 ( \19342 , \19341 , \11827 );
nor \U$18966 ( \19343 , \19340 , \19342 );
xor \U$18967 ( \19344 , \19336 , \19343 );
and \U$18968 ( \19345 , \14059 , RIae765c8_45);
and \U$18969 ( \19346 , RIae76118_35, \14057 );
nor \U$18970 ( \19347 , \19345 , \19346 );
and \U$18971 ( \19348 , \19347 , \13502 );
not \U$18972 ( \19349 , \19347 );
and \U$18973 ( \19350 , \19349 , \14063 );
nor \U$18974 ( \19351 , \19348 , \19350 );
and \U$18975 ( \19352 , \19344 , \19351 );
and \U$18976 ( \19353 , \19336 , \19343 );
or \U$18977 ( \19354 , \19352 , \19353 );
and \U$18978 ( \19355 , \19329 , \19354 );
and \U$18979 ( \19356 , \19310 , \19328 );
or \U$18980 ( \19357 , \19355 , \19356 );
xor \U$18981 ( \19358 , \19285 , \19357 );
and \U$18982 ( \19359 , \8371 , RIae75e48_29);
and \U$18983 ( \19360 , RIae75c68_25, \8369 );
nor \U$18984 ( \19361 , \19359 , \19360 );
and \U$18985 ( \19362 , \19361 , \8020 );
not \U$18986 ( \19363 , \19361 );
and \U$18987 ( \19364 , \19363 , \8019 );
nor \U$18988 ( \19365 , \19362 , \19364 );
and \U$18989 ( \19366 , \7633 , RIae758a8_17);
and \U$18990 ( \19367 , RIae75f38_31, \7631 );
nor \U$18991 ( \19368 , \19366 , \19367 );
and \U$18992 ( \19369 , \19368 , \7206 );
not \U$18993 ( \19370 , \19368 );
and \U$18994 ( \19371 , \19370 , \7205 );
nor \U$18995 ( \19372 , \19369 , \19371 );
xor \U$18996 ( \19373 , \19365 , \19372 );
and \U$18997 ( \19374 , \8966 , RIae75d58_27);
and \U$18998 ( \19375 , RIae755d8_11, \8964 );
nor \U$18999 ( \19376 , \19374 , \19375 );
and \U$19000 ( \19377 , \19376 , \8799 );
not \U$19001 ( \19378 , \19376 );
and \U$19002 ( \19379 , \19378 , \8789 );
nor \U$19003 ( \19380 , \19377 , \19379 );
and \U$19004 ( \19381 , \19373 , \19380 );
and \U$19005 ( \19382 , \19365 , \19372 );
or \U$19006 ( \19383 , \19381 , \19382 );
and \U$19007 ( \19384 , \4247 , RIae78530_112);
and \U$19008 ( \19385 , RIae77c48_93, \4245 );
nor \U$19009 ( \19386 , \19384 , \19385 );
and \U$19010 ( \19387 , \19386 , \3989 );
not \U$19011 ( \19388 , \19386 );
and \U$19012 ( \19389 , \19388 , \4251 );
nor \U$19013 ( \19390 , \19387 , \19389 );
and \U$19014 ( \19391 , \4688 , RIae77b58_91);
and \U$19015 ( \19392 , RIae77d38_95, \4686 );
nor \U$19016 ( \19393 , \19391 , \19392 );
and \U$19017 ( \19394 , \19393 , \4481 );
not \U$19018 ( \19395 , \19393 );
and \U$19019 ( \19396 , \19395 , \4482 );
nor \U$19020 ( \19397 , \19394 , \19396 );
xor \U$19021 ( \19398 , \19390 , \19397 );
and \U$19022 ( \19399 , \5399 , RIae77e28_97);
and \U$19023 ( \19400 , RIae78968_121, \5397 );
nor \U$19024 ( \19401 , \19399 , \19400 );
and \U$19025 ( \19402 , \19401 , \5016 );
not \U$19026 ( \19403 , \19401 );
and \U$19027 ( \19404 , \19403 , \5403 );
nor \U$19028 ( \19405 , \19402 , \19404 );
and \U$19029 ( \19406 , \19398 , \19405 );
and \U$19030 ( \19407 , \19390 , \19397 );
or \U$19031 ( \19408 , \19406 , \19407 );
xor \U$19032 ( \19409 , \19383 , \19408 );
and \U$19033 ( \19410 , \6941 , RIae75a88_21);
and \U$19034 ( \19411 , RIae75998_19, \6939 );
nor \U$19035 ( \19412 , \19410 , \19411 );
and \U$19036 ( \19413 , \19412 , \6314 );
not \U$19037 ( \19414 , \19412 );
and \U$19038 ( \19415 , \19414 , \6945 );
nor \U$19039 ( \19416 , \19413 , \19415 );
and \U$19040 ( \19417 , \5896 , RIae78878_119);
and \U$19041 ( \19418 , RIae78788_117, \5894 );
nor \U$19042 ( \19419 , \19417 , \19418 );
and \U$19043 ( \19420 , \19419 , \5590 );
not \U$19044 ( \19421 , \19419 );
and \U$19045 ( \19422 , \19421 , \5589 );
nor \U$19046 ( \19423 , \19420 , \19422 );
xor \U$19047 ( \19424 , \19416 , \19423 );
and \U$19048 ( \19425 , \6172 , RIae78698_115);
and \U$19049 ( \19426 , RIae75b78_23, \6170 );
nor \U$19050 ( \19427 , \19425 , \19426 );
and \U$19051 ( \19428 , \19427 , \6176 );
not \U$19052 ( \19429 , \19427 );
and \U$19053 ( \19430 , \19429 , \6175 );
nor \U$19054 ( \19431 , \19428 , \19430 );
and \U$19055 ( \19432 , \19424 , \19431 );
and \U$19056 ( \19433 , \19416 , \19423 );
or \U$19057 ( \19434 , \19432 , \19433 );
and \U$19058 ( \19435 , \19409 , \19434 );
and \U$19059 ( \19436 , \19383 , \19408 );
or \U$19060 ( \19437 , \19435 , \19436 );
and \U$19061 ( \19438 , \19358 , \19437 );
and \U$19062 ( \19439 , \19285 , \19357 );
or \U$19063 ( \19440 , \19438 , \19439 );
xor \U$19064 ( \19441 , \18552 , \471 );
xor \U$19065 ( \19442 , \19441 , \18560 );
xor \U$19066 ( \19443 , \18571 , \18578 );
xor \U$19067 ( \19444 , \19443 , \18586 );
and \U$19068 ( \19445 , \19442 , \19444 );
xor \U$19069 ( \19446 , \18928 , \18935 );
xor \U$19070 ( \19447 , \19446 , \18943 );
xor \U$19071 ( \19448 , \18903 , \18910 );
xor \U$19072 ( \19449 , \19448 , \18918 );
xor \U$19073 ( \19450 , \19447 , \19449 );
xor \U$19074 ( \19451 , \18957 , \18964 );
xor \U$19075 ( \19452 , \19451 , \18972 );
and \U$19076 ( \19453 , \19450 , \19452 );
and \U$19077 ( \19454 , \19447 , \19449 );
or \U$19078 ( \19455 , \19453 , \19454 );
xor \U$19079 ( \19456 , \18571 , \18578 );
xor \U$19080 ( \19457 , \19456 , \18586 );
and \U$19081 ( \19458 , \19455 , \19457 );
and \U$19082 ( \19459 , \19442 , \19455 );
or \U$19083 ( \19460 , \19445 , \19458 , \19459 );
xor \U$19084 ( \19461 , \19440 , \19460 );
xor \U$19085 ( \19462 , \18819 , \18826 );
xor \U$19086 ( \19463 , \19462 , \18835 );
xor \U$19087 ( \19464 , \18845 , \18852 );
xor \U$19088 ( \19465 , \19464 , \18860 );
xor \U$19089 ( \19466 , \19463 , \19465 );
not \U$19090 ( \19467 , \18871 );
xor \U$19091 ( \19468 , \18891 , \18880 );
not \U$19092 ( \19469 , \19468 );
or \U$19093 ( \19470 , \19467 , \19469 );
or \U$19094 ( \19471 , \19468 , \18871 );
nand \U$19095 ( \19472 , \19470 , \19471 );
and \U$19096 ( \19473 , \19466 , \19472 );
and \U$19097 ( \19474 , \19463 , \19465 );
or \U$19098 ( \19475 , \19473 , \19474 );
and \U$19099 ( \19476 , \672 , RIae77720_82);
and \U$19100 ( \19477 , RIae773d8_75, \670 );
nor \U$19101 ( \19478 , \19476 , \19477 );
and \U$19102 ( \19479 , \19478 , \588 );
not \U$19103 ( \19480 , \19478 );
and \U$19104 ( \19481 , \19480 , \587 );
nor \U$19105 ( \19482 , \19479 , \19481 );
and \U$19106 ( \19483 , \558 , RIae775b8_79);
and \U$19107 ( \19484 , RIae774c8_77, \556 );
nor \U$19108 ( \19485 , \19483 , \19484 );
and \U$19109 ( \19486 , \19485 , \504 );
not \U$19110 ( \19487 , \19485 );
and \U$19111 ( \19488 , \19487 , \562 );
nor \U$19112 ( \19489 , \19486 , \19488 );
xor \U$19113 ( \19490 , \19482 , \19489 );
nand \U$19114 ( \19491 , RIae775b8_79, \556 );
and \U$19115 ( \19492 , \19491 , \504 );
not \U$19116 ( \19493 , \19491 );
and \U$19117 ( \19494 , \19493 , \562 );
nor \U$19118 ( \19495 , \19492 , \19494 );
not \U$19119 ( \19496 , \19495 );
and \U$19120 ( \19497 , \672 , RIae774c8_77);
and \U$19121 ( \19498 , RIae77720_82, \670 );
nor \U$19122 ( \19499 , \19497 , \19498 );
and \U$19123 ( \19500 , \19499 , \588 );
not \U$19124 ( \19501 , \19499 );
and \U$19125 ( \19502 , \19501 , \587 );
nor \U$19126 ( \19503 , \19500 , \19502 );
not \U$19127 ( \19504 , \19503 );
or \U$19128 ( \19505 , \19496 , \19504 );
or \U$19129 ( \19506 , \19503 , \19495 );
not \U$19130 ( \19507 , \787 );
and \U$19131 ( \19508 , \883 , RIae773d8_75);
and \U$19132 ( \19509 , RIae77a68_89, \881 );
nor \U$19133 ( \19510 , \19508 , \19509 );
not \U$19134 ( \19511 , \19510 );
or \U$19135 ( \19512 , \19507 , \19511 );
or \U$19136 ( \19513 , \19510 , \789 );
nand \U$19137 ( \19514 , \19512 , \19513 );
nand \U$19138 ( \19515 , \19506 , \19514 );
nand \U$19139 ( \19516 , \19505 , \19515 );
and \U$19140 ( \19517 , \19490 , \19516 );
and \U$19141 ( \19518 , \19482 , \19489 );
or \U$19142 ( \19519 , \19517 , \19518 );
xor \U$19143 ( \19520 , \19475 , \19519 );
xor \U$19144 ( \19521 , \18985 , \18992 );
xor \U$19145 ( \19522 , \19521 , \19000 );
xor \U$19146 ( \19523 , \19039 , \19046 );
xor \U$19147 ( \19524 , \19523 , \19054 );
and \U$19148 ( \19525 , \19522 , \19524 );
xor \U$19149 ( \19526 , \19010 , \19017 );
xor \U$19150 ( \19527 , \19526 , \19025 );
xor \U$19151 ( \19528 , \19039 , \19046 );
xor \U$19152 ( \19529 , \19528 , \19054 );
and \U$19153 ( \19530 , \19527 , \19529 );
and \U$19154 ( \19531 , \19522 , \19527 );
or \U$19155 ( \19532 , \19525 , \19530 , \19531 );
and \U$19156 ( \19533 , \19520 , \19532 );
and \U$19157 ( \19534 , \19475 , \19519 );
or \U$19158 ( \19535 , \19533 , \19534 );
and \U$19159 ( \19536 , \19461 , \19535 );
and \U$19160 ( \19537 , \19440 , \19460 );
or \U$19161 ( \19538 , \19536 , \19537 );
xor \U$19162 ( \19539 , \19204 , \19538 );
not \U$19163 ( \19540 , \18975 );
not \U$19164 ( \19541 , \18946 );
or \U$19165 ( \19542 , \19540 , \19541 );
or \U$19166 ( \19543 , \18946 , \18975 );
nand \U$19167 ( \19544 , \19542 , \19543 );
not \U$19168 ( \19545 , \19544 );
not \U$19169 ( \19546 , \18921 );
and \U$19170 ( \19547 , \19545 , \19546 );
and \U$19171 ( \19548 , \19544 , \18921 );
nor \U$19172 ( \19549 , \19547 , \19548 );
not \U$19173 ( \19550 , \19549 );
xor \U$19174 ( \19551 , \18838 , \18863 );
xor \U$19175 ( \19552 , \19551 , \18893 );
not \U$19176 ( \19553 , \19552 );
and \U$19177 ( \19554 , \19550 , \19553 );
and \U$19178 ( \19555 , \19549 , \19552 );
not \U$19179 ( \19556 , \19057 );
not \U$19180 ( \19557 , \19003 );
or \U$19181 ( \19558 , \19556 , \19557 );
or \U$19182 ( \19559 , \19003 , \19057 );
nand \U$19183 ( \19560 , \19558 , \19559 );
not \U$19184 ( \19561 , \19560 );
not \U$19185 ( \19562 , \19028 );
and \U$19186 ( \19563 , \19561 , \19562 );
and \U$19187 ( \19564 , \19560 , \19028 );
nor \U$19188 ( \19565 , \19563 , \19564 );
nor \U$19189 ( \19566 , \19555 , \19565 );
nor \U$19190 ( \19567 , \19554 , \19566 );
not \U$19191 ( \19568 , \18518 );
not \U$19192 ( \19569 , \18462 );
or \U$19193 ( \19570 , \19568 , \19569 );
or \U$19194 ( \19571 , \18462 , \18518 );
nand \U$19195 ( \19572 , \19570 , \19571 );
not \U$19196 ( \19573 , \19572 );
not \U$19197 ( \19574 , \18489 );
and \U$19198 ( \19575 , \19573 , \19574 );
and \U$19199 ( \19576 , \19572 , \18489 );
nor \U$19200 ( \19577 , \19575 , \19576 );
or \U$19201 ( \19578 , \19567 , \19577 );
not \U$19202 ( \19579 , \19577 );
not \U$19203 ( \19580 , \19567 );
or \U$19204 ( \19581 , \19579 , \19580 );
xor \U$19205 ( \19582 , \18390 , \18397 );
xor \U$19206 ( \19583 , \19582 , \18406 );
xor \U$19207 ( \19584 , \19079 , \19084 );
xor \U$19208 ( \19585 , \19583 , \19584 );
xor \U$19209 ( \19586 , \19065 , \19067 );
xor \U$19210 ( \19587 , \19586 , \19070 );
and \U$19211 ( \19588 , \19585 , \19587 );
xor \U$19212 ( \19589 , \19096 , \19102 );
xor \U$19213 ( \19590 , \19589 , \19105 );
xor \U$19214 ( \19591 , \19065 , \19067 );
xor \U$19215 ( \19592 , \19591 , \19070 );
and \U$19216 ( \19593 , \19590 , \19592 );
and \U$19217 ( \19594 , \19585 , \19590 );
or \U$19218 ( \19595 , \19588 , \19593 , \19594 );
nand \U$19219 ( \19596 , \19581 , \19595 );
nand \U$19220 ( \19597 , \19578 , \19596 );
and \U$19221 ( \19598 , \19539 , \19597 );
and \U$19222 ( \19599 , \19204 , \19538 );
or \U$19223 ( \19600 , \19598 , \19599 );
xor \U$19224 ( \19601 , \19190 , \19600 );
xor \U$19225 ( \19602 , \18702 , \18714 );
xor \U$19226 ( \19603 , \19602 , \18719 );
xor \U$19227 ( \19604 , \19147 , \19154 );
xor \U$19228 ( \19605 , \19603 , \19604 );
xor \U$19229 ( \19606 , \19601 , \19605 );
xor \U$19230 ( \19607 , \19475 , \19519 );
xor \U$19231 ( \19608 , \19607 , \19532 );
xor \U$19232 ( \19609 , \19285 , \19357 );
xor \U$19233 ( \19610 , \19609 , \19437 );
xor \U$19234 ( \19611 , \19608 , \19610 );
xor \U$19235 ( \19612 , \18571 , \18578 );
xor \U$19236 ( \19613 , \19612 , \18586 );
xor \U$19237 ( \19614 , \19442 , \19455 );
xor \U$19238 ( \19615 , \19613 , \19614 );
and \U$19239 ( \19616 , \19611 , \19615 );
and \U$19240 ( \19617 , \19608 , \19610 );
or \U$19241 ( \19618 , \19616 , \19617 );
xor \U$19242 ( \19619 , \19262 , \19270 );
xor \U$19243 ( \19620 , \19619 , \19279 );
xor \U$19244 ( \19621 , \19390 , \19397 );
xor \U$19245 ( \19622 , \19621 , \19405 );
xor \U$19246 ( \19623 , \19620 , \19622 );
xor \U$19247 ( \19624 , \19416 , \19423 );
xor \U$19248 ( \19625 , \19624 , \19431 );
and \U$19249 ( \19626 , \19623 , \19625 );
and \U$19250 ( \19627 , \19620 , \19622 );
or \U$19251 ( \19628 , \19626 , \19627 );
xnor \U$19252 ( \19629 , \19514 , \19503 );
not \U$19253 ( \19630 , \19629 );
not \U$19254 ( \19631 , \19495 );
and \U$19255 ( \19632 , \19630 , \19631 );
and \U$19256 ( \19633 , \19629 , \19495 );
nor \U$19257 ( \19634 , \19632 , \19633 );
xor \U$19258 ( \19635 , \19236 , \19243 );
xor \U$19259 ( \19636 , \19635 , \19251 );
or \U$19260 ( \19637 , \19634 , \19636 );
not \U$19261 ( \19638 , \19636 );
not \U$19262 ( \19639 , \19634 );
or \U$19263 ( \19640 , \19638 , \19639 );
xor \U$19264 ( \19641 , \19211 , \19218 );
xor \U$19265 ( \19642 , \19641 , \19226 );
nand \U$19266 ( \19643 , \19640 , \19642 );
nand \U$19267 ( \19644 , \19637 , \19643 );
xor \U$19268 ( \19645 , \19628 , \19644 );
xor \U$19269 ( \19646 , \19365 , \19372 );
xor \U$19270 ( \19647 , \19646 , \19380 );
xor \U$19271 ( \19648 , \19336 , \19343 );
xor \U$19272 ( \19649 , \19648 , \19351 );
and \U$19273 ( \19650 , \19647 , \19649 );
xor \U$19274 ( \19651 , \19292 , \19299 );
xor \U$19275 ( \19652 , \19651 , \19307 );
xor \U$19276 ( \19653 , \19336 , \19343 );
xor \U$19277 ( \19654 , \19653 , \19351 );
and \U$19278 ( \19655 , \19652 , \19654 );
and \U$19279 ( \19656 , \19647 , \19652 );
or \U$19280 ( \19657 , \19650 , \19655 , \19656 );
and \U$19281 ( \19658 , \19645 , \19657 );
and \U$19282 ( \19659 , \19628 , \19644 );
or \U$19283 ( \19660 , \19658 , \19659 );
and \U$19284 ( \19661 , \1138 , RIae77a68_89);
and \U$19285 ( \19662 , RIae77978_87, \1136 );
nor \U$19286 ( \19663 , \19661 , \19662 );
and \U$19287 ( \19664 , \19663 , \1012 );
not \U$19288 ( \19665 , \19663 );
and \U$19289 ( \19666 , \19665 , \1142 );
nor \U$19290 ( \19667 , \19664 , \19666 );
and \U$19291 ( \19668 , \1376 , RIae77798_83);
and \U$19292 ( \19669 , RIae77888_85, \1374 );
nor \U$19293 ( \19670 , \19668 , \19669 );
and \U$19294 ( \19671 , \19670 , \1380 );
not \U$19295 ( \19672 , \19670 );
and \U$19296 ( \19673 , \19672 , \1261 );
nor \U$19297 ( \19674 , \19671 , \19673 );
xor \U$19298 ( \19675 , \19667 , \19674 );
not \U$19299 ( \19676 , \789 );
and \U$19300 ( \19677 , \883 , RIae77720_82);
and \U$19301 ( \19678 , RIae773d8_75, \881 );
nor \U$19302 ( \19679 , \19677 , \19678 );
not \U$19303 ( \19680 , \19679 );
or \U$19304 ( \19681 , \19676 , \19680 );
or \U$19305 ( \19682 , \19679 , \789 );
nand \U$19306 ( \19683 , \19681 , \19682 );
and \U$19307 ( \19684 , \19675 , \19683 );
and \U$19308 ( \19685 , \19667 , \19674 );
nor \U$19309 ( \19686 , \19684 , \19685 );
and \U$19310 ( \19687 , \1593 , RIae76f28_65);
and \U$19311 ( \19688 , RIae76e38_63, \1591 );
nor \U$19312 ( \19689 , \19687 , \19688 );
and \U$19313 ( \19690 , \19689 , \1488 );
not \U$19314 ( \19691 , \19689 );
and \U$19315 ( \19692 , \19691 , \1498 );
nor \U$19316 ( \19693 , \19690 , \19692 );
and \U$19317 ( \19694 , \1939 , RIae76d48_61);
and \U$19318 ( \19695 , RIae76c58_59, \1937 );
nor \U$19319 ( \19696 , \19694 , \19695 );
and \U$19320 ( \19697 , \19696 , \1734 );
not \U$19321 ( \19698 , \19696 );
and \U$19322 ( \19699 , \19698 , \1735 );
nor \U$19323 ( \19700 , \19697 , \19699 );
xor \U$19324 ( \19701 , \19693 , \19700 );
and \U$19325 ( \19702 , \2224 , RIae77180_70);
and \U$19326 ( \19703 , RIae77018_67, \2222 );
nor \U$19327 ( \19704 , \19702 , \19703 );
and \U$19328 ( \19705 , \19704 , \2060 );
not \U$19329 ( \19706 , \19704 );
and \U$19330 ( \19707 , \19706 , \2061 );
nor \U$19331 ( \19708 , \19705 , \19707 );
and \U$19332 ( \19709 , \19701 , \19708 );
and \U$19333 ( \19710 , \19693 , \19700 );
or \U$19334 ( \19711 , \19709 , \19710 );
xor \U$19335 ( \19712 , \19686 , \19711 );
and \U$19336 ( \19713 , \3214 , RIae77f18_99);
and \U$19337 ( \19714 , RIae78008_101, \3212 );
nor \U$19338 ( \19715 , \19713 , \19714 );
not \U$19339 ( \19716 , \19715 );
not \U$19340 ( \19717 , \3218 );
and \U$19341 ( \19718 , \19716 , \19717 );
and \U$19342 ( \19719 , \19715 , \2774 );
nor \U$19343 ( \19720 , \19718 , \19719 );
and \U$19344 ( \19721 , \2607 , RIae771f8_71);
and \U$19345 ( \19722 , RIae772e8_73, \2605 );
nor \U$19346 ( \19723 , \19721 , \19722 );
and \U$19347 ( \19724 , \19723 , \2397 );
not \U$19348 ( \19725 , \19723 );
and \U$19349 ( \19726 , \19725 , \2611 );
nor \U$19350 ( \19727 , \19724 , \19726 );
xor \U$19351 ( \19728 , \19720 , \19727 );
and \U$19352 ( \19729 , \2783 , RIae782d8_107);
and \U$19353 ( \19730 , RIae780f8_103, \2781 );
nor \U$19354 ( \19731 , \19729 , \19730 );
not \U$19355 ( \19732 , \19731 );
not \U$19356 ( \19733 , \2789 );
and \U$19357 ( \19734 , \19732 , \19733 );
and \U$19358 ( \19735 , \19731 , \2789 );
nor \U$19359 ( \19736 , \19734 , \19735 );
and \U$19360 ( \19737 , \19728 , \19736 );
and \U$19361 ( \19738 , \19720 , \19727 );
or \U$19362 ( \19739 , \19737 , \19738 );
and \U$19363 ( \19740 , \19712 , \19739 );
and \U$19364 ( \19741 , \19686 , \19711 );
nor \U$19365 ( \19742 , \19740 , \19741 );
and \U$19366 ( \19743 , \14059 , RIae766b8_47);
and \U$19367 ( \19744 , RIae765c8_45, \14057 );
nor \U$19368 ( \19745 , \19743 , \19744 );
and \U$19369 ( \19746 , \19745 , \14063 );
not \U$19370 ( \19747 , \19745 );
and \U$19371 ( \19748 , \19747 , \13502 );
nor \U$19372 ( \19749 , \19746 , \19748 );
and \U$19373 ( \19750 , \15726 , RIae762f8_39);
and \U$19374 ( \19751 , RIae7aab0_192, RIae76208_37);
nor \U$19375 ( \19752 , \19750 , \19751 );
and \U$19376 ( \19753 , \19752 , RIae7aa38_191);
not \U$19377 ( \19754 , \19752 );
and \U$19378 ( \19755 , \19754 , \14959 );
nor \U$19379 ( \19756 , \19753 , \19755 );
xor \U$19380 ( \19757 , \19749 , \19756 );
and \U$19381 ( \19758 , \14964 , RIae76118_35);
and \U$19382 ( \19759 , RIae76028_33, \14962 );
nor \U$19383 ( \19760 , \19758 , \19759 );
and \U$19384 ( \19761 , \19760 , \14462 );
not \U$19385 ( \19762 , \19760 );
and \U$19386 ( \19763 , \19762 , \14463 );
nor \U$19387 ( \19764 , \19761 , \19763 );
and \U$19388 ( \19765 , \19757 , \19764 );
and \U$19389 ( \19766 , \19749 , \19756 );
or \U$19390 ( \19767 , \19765 , \19766 );
and \U$19391 ( \19768 , \8966 , RIae75c68_25);
and \U$19392 ( \19769 , RIae75d58_27, \8964 );
nor \U$19393 ( \19770 , \19768 , \19769 );
and \U$19394 ( \19771 , \19770 , \8789 );
not \U$19395 ( \19772 , \19770 );
and \U$19396 ( \19773 , \19772 , \8799 );
nor \U$19397 ( \19774 , \19771 , \19773 );
not \U$19398 ( \19775 , \19774 );
and \U$19399 ( \19776 , \10548 , RIae757b8_15);
and \U$19400 ( \19777 , RIae756c8_13, \10546 );
nor \U$19401 ( \19778 , \19776 , \19777 );
and \U$19402 ( \19779 , \19778 , \10118 );
not \U$19403 ( \19780 , \19778 );
and \U$19404 ( \19781 , \19780 , \10421 );
nor \U$19405 ( \19782 , \19779 , \19781 );
not \U$19406 ( \19783 , \19782 );
and \U$19407 ( \19784 , \19775 , \19783 );
and \U$19408 ( \19785 , \19782 , \19774 );
and \U$19409 ( \19786 , \9760 , RIae755d8_11);
and \U$19410 ( \19787 , RIae754e8_9, \9758 );
nor \U$19411 ( \19788 , \19786 , \19787 );
and \U$19412 ( \19789 , \19788 , \9272 );
not \U$19413 ( \19790 , \19788 );
and \U$19414 ( \19791 , \19790 , \9273 );
nor \U$19415 ( \19792 , \19789 , \19791 );
nor \U$19416 ( \19793 , \19785 , \19792 );
nor \U$19417 ( \19794 , \19784 , \19793 );
xor \U$19418 ( \19795 , \19767 , \19794 );
and \U$19419 ( \19796 , \13059 , RIae763e8_41);
and \U$19420 ( \19797 , RIae764d8_43, \13057 );
nor \U$19421 ( \19798 , \19796 , \19797 );
and \U$19422 ( \19799 , \19798 , \12718 );
not \U$19423 ( \19800 , \19798 );
and \U$19424 ( \19801 , \19800 , \13063 );
nor \U$19425 ( \19802 , \19799 , \19801 );
and \U$19426 ( \19803 , \11470 , RIae75218_3);
and \U$19427 ( \19804 , RIae75128_1, \11468 );
nor \U$19428 ( \19805 , \19803 , \19804 );
and \U$19429 ( \19806 , \19805 , \11474 );
not \U$19430 ( \19807 , \19805 );
and \U$19431 ( \19808 , \19807 , \10936 );
nor \U$19432 ( \19809 , \19806 , \19808 );
xor \U$19433 ( \19810 , \19802 , \19809 );
and \U$19434 ( \19811 , \12180 , RIae75308_5);
and \U$19435 ( \19812 , RIae753f8_7, \12178 );
nor \U$19436 ( \19813 , \19811 , \19812 );
and \U$19437 ( \19814 , \19813 , \11827 );
not \U$19438 ( \19815 , \19813 );
and \U$19439 ( \19816 , \19815 , \12184 );
nor \U$19440 ( \19817 , \19814 , \19816 );
and \U$19441 ( \19818 , \19810 , \19817 );
and \U$19442 ( \19819 , \19802 , \19809 );
or \U$19443 ( \19820 , \19818 , \19819 );
and \U$19444 ( \19821 , \19795 , \19820 );
and \U$19445 ( \19822 , \19767 , \19794 );
nor \U$19446 ( \19823 , \19821 , \19822 );
xor \U$19447 ( \19824 , \19742 , \19823 );
and \U$19448 ( \19825 , \3730 , RIae781e8_105);
and \U$19449 ( \19826 , RIae785a8_113, \3728 );
nor \U$19450 ( \19827 , \19825 , \19826 );
and \U$19451 ( \19828 , \19827 , \3422 );
not \U$19452 ( \19829 , \19827 );
and \U$19453 ( \19830 , \19829 , \3732 );
nor \U$19454 ( \19831 , \19828 , \19830 );
and \U$19455 ( \19832 , \4247 , RIae783c8_109);
and \U$19456 ( \19833 , RIae78530_112, \4245 );
nor \U$19457 ( \19834 , \19832 , \19833 );
and \U$19458 ( \19835 , \19834 , \4251 );
not \U$19459 ( \19836 , \19834 );
and \U$19460 ( \19837 , \19836 , \3989 );
nor \U$19461 ( \19838 , \19835 , \19837 );
xor \U$19462 ( \19839 , \19831 , \19838 );
and \U$19463 ( \19840 , \4688 , RIae77c48_93);
and \U$19464 ( \19841 , RIae77b58_91, \4686 );
nor \U$19465 ( \19842 , \19840 , \19841 );
and \U$19466 ( \19843 , \19842 , \4482 );
not \U$19467 ( \19844 , \19842 );
and \U$19468 ( \19845 , \19844 , \4481 );
nor \U$19469 ( \19846 , \19843 , \19845 );
and \U$19470 ( \19847 , \19839 , \19846 );
and \U$19471 ( \19848 , \19831 , \19838 );
or \U$19472 ( \19849 , \19847 , \19848 );
and \U$19473 ( \19850 , \6941 , RIae75b78_23);
and \U$19474 ( \19851 , RIae75a88_21, \6939 );
nor \U$19475 ( \19852 , \19850 , \19851 );
and \U$19476 ( \19853 , \19852 , \6945 );
not \U$19477 ( \19854 , \19852 );
and \U$19478 ( \19855 , \19854 , \6314 );
nor \U$19479 ( \19856 , \19853 , \19855 );
and \U$19480 ( \19857 , \7633 , RIae75998_19);
and \U$19481 ( \19858 , RIae758a8_17, \7631 );
nor \U$19482 ( \19859 , \19857 , \19858 );
and \U$19483 ( \19860 , \19859 , \7205 );
not \U$19484 ( \19861 , \19859 );
and \U$19485 ( \19862 , \19861 , \7206 );
nor \U$19486 ( \19863 , \19860 , \19862 );
xor \U$19487 ( \19864 , \19856 , \19863 );
and \U$19488 ( \19865 , \8371 , RIae75f38_31);
and \U$19489 ( \19866 , RIae75e48_29, \8369 );
nor \U$19490 ( \19867 , \19865 , \19866 );
and \U$19491 ( \19868 , \19867 , \8019 );
not \U$19492 ( \19869 , \19867 );
and \U$19493 ( \19870 , \19869 , \8020 );
nor \U$19494 ( \19871 , \19868 , \19870 );
and \U$19495 ( \19872 , \19864 , \19871 );
and \U$19496 ( \19873 , \19856 , \19863 );
or \U$19497 ( \19874 , \19872 , \19873 );
xor \U$19498 ( \19875 , \19849 , \19874 );
and \U$19499 ( \19876 , \5896 , RIae78968_121);
and \U$19500 ( \19877 , RIae78878_119, \5894 );
nor \U$19501 ( \19878 , \19876 , \19877 );
and \U$19502 ( \19879 , \19878 , \5589 );
not \U$19503 ( \19880 , \19878 );
and \U$19504 ( \19881 , \19880 , \5590 );
nor \U$19505 ( \19882 , \19879 , \19881 );
and \U$19506 ( \19883 , \5399 , RIae77d38_95);
and \U$19507 ( \19884 , RIae77e28_97, \5397 );
nor \U$19508 ( \19885 , \19883 , \19884 );
and \U$19509 ( \19886 , \19885 , \5403 );
not \U$19510 ( \19887 , \19885 );
and \U$19511 ( \19888 , \19887 , \5016 );
nor \U$19512 ( \19889 , \19886 , \19888 );
xor \U$19513 ( \19890 , \19882 , \19889 );
and \U$19514 ( \19891 , \6172 , RIae78788_117);
and \U$19515 ( \19892 , RIae78698_115, \6170 );
nor \U$19516 ( \19893 , \19891 , \19892 );
and \U$19517 ( \19894 , \19893 , \6175 );
not \U$19518 ( \19895 , \19893 );
and \U$19519 ( \19896 , \19895 , \6176 );
nor \U$19520 ( \19897 , \19894 , \19896 );
and \U$19521 ( \19898 , \19890 , \19897 );
and \U$19522 ( \19899 , \19882 , \19889 );
or \U$19523 ( \19900 , \19898 , \19899 );
and \U$19524 ( \19901 , \19875 , \19900 );
and \U$19525 ( \19902 , \19849 , \19874 );
nor \U$19526 ( \19903 , \19901 , \19902 );
and \U$19527 ( \19904 , \19824 , \19903 );
and \U$19528 ( \19905 , \19742 , \19823 );
or \U$19529 ( \19906 , \19904 , \19905 );
xor \U$19530 ( \19907 , \19660 , \19906 );
xor \U$19531 ( \19908 , \19463 , \19465 );
xor \U$19532 ( \19909 , \19908 , \19472 );
xor \U$19533 ( \19910 , \19447 , \19449 );
xor \U$19534 ( \19911 , \19910 , \19452 );
and \U$19535 ( \19912 , \19909 , \19911 );
xor \U$19536 ( \19913 , \19039 , \19046 );
xor \U$19537 ( \19914 , \19913 , \19054 );
xor \U$19538 ( \19915 , \19522 , \19527 );
xor \U$19539 ( \19916 , \19914 , \19915 );
xor \U$19540 ( \19917 , \19447 , \19449 );
xor \U$19541 ( \19918 , \19917 , \19452 );
and \U$19542 ( \19919 , \19916 , \19918 );
and \U$19543 ( \19920 , \19909 , \19916 );
or \U$19544 ( \19921 , \19912 , \19919 , \19920 );
and \U$19545 ( \19922 , \19907 , \19921 );
and \U$19546 ( \19923 , \19660 , \19906 );
or \U$19547 ( \19924 , \19922 , \19923 );
xor \U$19548 ( \19925 , \19618 , \19924 );
not \U$19549 ( \19926 , \19549 );
xor \U$19550 ( \19927 , \19552 , \19565 );
not \U$19551 ( \19928 , \19927 );
or \U$19552 ( \19929 , \19926 , \19928 );
or \U$19553 ( \19930 , \19927 , \19549 );
nand \U$19554 ( \19931 , \19929 , \19930 );
xor \U$19555 ( \19932 , \19482 , \19489 );
xor \U$19556 ( \19933 , \19932 , \19516 );
xor \U$19557 ( \19934 , \19229 , \19254 );
xor \U$19558 ( \19935 , \19934 , \19282 );
and \U$19559 ( \19936 , \19933 , \19935 );
xor \U$19560 ( \19937 , \19383 , \19408 );
xor \U$19561 ( \19938 , \19937 , \19434 );
xor \U$19562 ( \19939 , \19229 , \19254 );
xor \U$19563 ( \19940 , \19939 , \19282 );
and \U$19564 ( \19941 , \19938 , \19940 );
and \U$19565 ( \19942 , \19933 , \19938 );
or \U$19566 ( \19943 , \19936 , \19941 , \19942 );
xor \U$19567 ( \19944 , \19931 , \19943 );
xor \U$19568 ( \19945 , \19065 , \19067 );
xor \U$19569 ( \19946 , \19945 , \19070 );
xor \U$19570 ( \19947 , \19585 , \19590 );
xor \U$19571 ( \19948 , \19946 , \19947 );
and \U$19572 ( \19949 , \19944 , \19948 );
and \U$19573 ( \19950 , \19931 , \19943 );
or \U$19574 ( \19951 , \19949 , \19950 );
and \U$19575 ( \19952 , \19925 , \19951 );
and \U$19576 ( \19953 , \19618 , \19924 );
or \U$19577 ( \19954 , \19952 , \19953 );
xor \U$19578 ( \19955 , \19073 , \19089 );
xor \U$19579 ( \19956 , \19955 , \19108 );
xor \U$19580 ( \19957 , \18896 , \18977 );
xor \U$19581 ( \19958 , \19957 , \19059 );
xor \U$19582 ( \19959 , \19956 , \19958 );
xor \U$19583 ( \19960 , \18802 , \18804 );
xor \U$19584 ( \19961 , \19960 , \18809 );
xor \U$19585 ( \19962 , \19192 , \19199 );
xor \U$19586 ( \19963 , \19961 , \19962 );
and \U$19587 ( \19964 , \19959 , \19963 );
and \U$19588 ( \19965 , \19956 , \19958 );
or \U$19589 ( \19966 , \19964 , \19965 );
xor \U$19590 ( \19967 , \19954 , \19966 );
xor \U$19591 ( \19968 , \19129 , \19131 );
xor \U$19592 ( \19969 , \19968 , \19136 );
xor \U$19593 ( \19970 , \19178 , \19185 );
xor \U$19594 ( \19971 , \19969 , \19970 );
and \U$19595 ( \19972 , \19967 , \19971 );
and \U$19596 ( \19973 , \19954 , \19966 );
or \U$19597 ( \19974 , \19972 , \19973 );
xor \U$19598 ( \19975 , \19606 , \19974 );
xor \U$19599 ( \19976 , \18800 , \19114 );
xor \U$19600 ( \19977 , \19976 , \19139 );
and \U$19601 ( \19978 , \19975 , \19977 );
and \U$19602 ( \19979 , \19606 , \19974 );
nor \U$19603 ( \19980 , \19978 , \19979 );
not \U$19604 ( \19981 , \19980 );
xor \U$19605 ( \19982 , \19142 , \19144 );
xor \U$19606 ( \19983 , \19982 , \19159 );
xor \U$19607 ( \19984 , \19190 , \19600 );
and \U$19608 ( \19985 , \19984 , \19605 );
and \U$19609 ( \19986 , \19190 , \19600 );
or \U$19610 ( \19987 , \19985 , \19986 );
xor \U$19611 ( \19988 , \18727 , \18729 );
xor \U$19612 ( \19989 , \19988 , \18734 );
xor \U$19613 ( \19990 , \18775 , \18780 );
xor \U$19614 ( \19991 , \19989 , \19990 );
xor \U$19615 ( \19992 , \19987 , \19991 );
xor \U$19616 ( \19993 , \19983 , \19992 );
not \U$19617 ( \19994 , \19993 );
or \U$19618 ( \19995 , \19981 , \19994 );
or \U$19619 ( \19996 , \19993 , \19980 );
nand \U$19620 ( \19997 , \19995 , \19996 );
xor \U$19621 ( \19998 , \19606 , \19974 );
xor \U$19622 ( \19999 , \19998 , \19977 );
not \U$19623 ( \20000 , \19999 );
xor \U$19624 ( \20001 , \19204 , \19538 );
xor \U$19625 ( \20002 , \20001 , \19597 );
xor \U$19626 ( \20003 , \19440 , \19460 );
xor \U$19627 ( \20004 , \20003 , \19535 );
xor \U$19628 ( \20005 , \19956 , \19958 );
xor \U$19629 ( \20006 , \20005 , \19963 );
and \U$19630 ( \20007 , \20004 , \20006 );
xor \U$19631 ( \20008 , \19618 , \19924 );
xor \U$19632 ( \20009 , \20008 , \19951 );
xor \U$19633 ( \20010 , \19956 , \19958 );
xor \U$19634 ( \20011 , \20010 , \19963 );
and \U$19635 ( \20012 , \20009 , \20011 );
and \U$19636 ( \20013 , \20004 , \20009 );
or \U$19637 ( \20014 , \20007 , \20012 , \20013 );
xor \U$19638 ( \20015 , \20002 , \20014 );
xor \U$19639 ( \20016 , \19742 , \19823 );
xor \U$19640 ( \20017 , \20016 , \19903 );
xor \U$19641 ( \20018 , \19628 , \19644 );
xor \U$19642 ( \20019 , \20018 , \19657 );
and \U$19643 ( \20020 , \20017 , \20019 );
xor \U$19644 ( \20021 , \19447 , \19449 );
xor \U$19645 ( \20022 , \20021 , \19452 );
xor \U$19646 ( \20023 , \19909 , \19916 );
xor \U$19647 ( \20024 , \20022 , \20023 );
xor \U$19648 ( \20025 , \19628 , \19644 );
xor \U$19649 ( \20026 , \20025 , \19657 );
and \U$19650 ( \20027 , \20024 , \20026 );
and \U$19651 ( \20028 , \20017 , \20024 );
or \U$19652 ( \20029 , \20020 , \20027 , \20028 );
not \U$19653 ( \20030 , \20029 );
not \U$19654 ( \20031 , \20030 );
xor \U$19655 ( \20032 , \19229 , \19254 );
xor \U$19656 ( \20033 , \20032 , \19282 );
xor \U$19657 ( \20034 , \19933 , \19938 );
xor \U$19658 ( \20035 , \20033 , \20034 );
xor \U$19659 ( \20036 , \19310 , \19328 );
xor \U$19660 ( \20037 , \20036 , \19354 );
and \U$19661 ( \20038 , \20035 , \20037 );
not \U$19662 ( \20039 , \20035 );
not \U$19663 ( \20040 , \20037 );
and \U$19664 ( \20041 , \20039 , \20040 );
xor \U$19665 ( \20042 , \19849 , \19874 );
xor \U$19666 ( \20043 , \20042 , \19900 );
xor \U$19667 ( \20044 , \19686 , \19711 );
xor \U$19668 ( \20045 , \20044 , \19739 );
xor \U$19669 ( \20046 , \20043 , \20045 );
not \U$19670 ( \20047 , \19642 );
not \U$19671 ( \20048 , \19634 );
or \U$19672 ( \20049 , \20047 , \20048 );
or \U$19673 ( \20050 , \19634 , \19642 );
nand \U$19674 ( \20051 , \20049 , \20050 );
not \U$19675 ( \20052 , \20051 );
not \U$19676 ( \20053 , \19636 );
and \U$19677 ( \20054 , \20052 , \20053 );
and \U$19678 ( \20055 , \20051 , \19636 );
nor \U$19679 ( \20056 , \20054 , \20055 );
and \U$19680 ( \20057 , \20046 , \20056 );
and \U$19681 ( \20058 , \20043 , \20045 );
or \U$19682 ( \20059 , \20057 , \20058 );
nor \U$19683 ( \20060 , \20041 , \20059 );
nor \U$19684 ( \20061 , \20038 , \20060 );
not \U$19685 ( \20062 , \20061 );
and \U$19686 ( \20063 , \20031 , \20062 );
and \U$19687 ( \20064 , \20030 , \20061 );
xor \U$19688 ( \20065 , \19831 , \19838 );
xor \U$19689 ( \20066 , \20065 , \19846 );
xor \U$19690 ( \20067 , \19882 , \19889 );
xor \U$19691 ( \20068 , \20067 , \19897 );
xor \U$19692 ( \20069 , \20066 , \20068 );
xor \U$19693 ( \20070 , \19720 , \19727 );
xor \U$19694 ( \20071 , \20070 , \19736 );
and \U$19695 ( \20072 , \20069 , \20071 );
and \U$19696 ( \20073 , \20066 , \20068 );
nor \U$19697 ( \20074 , \20072 , \20073 );
xor \U$19698 ( \20075 , \19693 , \19700 );
xor \U$19699 ( \20076 , \20075 , \19708 );
and \U$19700 ( \20077 , \672 , RIae775b8_79);
and \U$19701 ( \20078 , RIae774c8_77, \670 );
nor \U$19702 ( \20079 , \20077 , \20078 );
and \U$19703 ( \20080 , \20079 , \587 );
not \U$19704 ( \20081 , \20079 );
and \U$19705 ( \20082 , \20081 , \588 );
nor \U$19706 ( \20083 , \20080 , \20082 );
or \U$19707 ( \20084 , \20076 , \20083 );
not \U$19708 ( \20085 , \20083 );
not \U$19709 ( \20086 , \20076 );
or \U$19710 ( \20087 , \20085 , \20086 );
xor \U$19711 ( \20088 , \19667 , \19674 );
xor \U$19712 ( \20089 , \20088 , \19683 );
nand \U$19713 ( \20090 , \20087 , \20089 );
nand \U$19714 ( \20091 , \20084 , \20090 );
xor \U$19715 ( \20092 , \20074 , \20091 );
xor \U$19716 ( \20093 , \19856 , \19863 );
xor \U$19717 ( \20094 , \20093 , \19871 );
xor \U$19718 ( \20095 , \19802 , \19809 );
xor \U$19719 ( \20096 , \20095 , \19817 );
or \U$19720 ( \20097 , \20094 , \20096 );
not \U$19721 ( \20098 , \20096 );
not \U$19722 ( \20099 , \20094 );
or \U$19723 ( \20100 , \20098 , \20099 );
not \U$19724 ( \20101 , \19774 );
xor \U$19725 ( \20102 , \19792 , \19782 );
not \U$19726 ( \20103 , \20102 );
or \U$19727 ( \20104 , \20101 , \20103 );
or \U$19728 ( \20105 , \20102 , \19774 );
nand \U$19729 ( \20106 , \20104 , \20105 );
nand \U$19730 ( \20107 , \20100 , \20106 );
nand \U$19731 ( \20108 , \20097 , \20107 );
and \U$19732 ( \20109 , \20092 , \20108 );
and \U$19733 ( \20110 , \20074 , \20091 );
or \U$19734 ( \20111 , \20109 , \20110 );
and \U$19735 ( \20112 , \5399 , RIae77b58_91);
and \U$19736 ( \20113 , RIae77d38_95, \5397 );
nor \U$19737 ( \20114 , \20112 , \20113 );
and \U$19738 ( \20115 , \20114 , \5403 );
not \U$19739 ( \20116 , \20114 );
and \U$19740 ( \20117 , \20116 , \5016 );
nor \U$19741 ( \20118 , \20115 , \20117 );
and \U$19742 ( \20119 , \4247 , RIae785a8_113);
and \U$19743 ( \20120 , RIae783c8_109, \4245 );
nor \U$19744 ( \20121 , \20119 , \20120 );
and \U$19745 ( \20122 , \20121 , \4251 );
not \U$19746 ( \20123 , \20121 );
and \U$19747 ( \20124 , \20123 , \3989 );
nor \U$19748 ( \20125 , \20122 , \20124 );
xor \U$19749 ( \20126 , \20118 , \20125 );
and \U$19750 ( \20127 , \4688 , RIae78530_112);
and \U$19751 ( \20128 , RIae77c48_93, \4686 );
nor \U$19752 ( \20129 , \20127 , \20128 );
and \U$19753 ( \20130 , \20129 , \4482 );
not \U$19754 ( \20131 , \20129 );
and \U$19755 ( \20132 , \20131 , \4481 );
nor \U$19756 ( \20133 , \20130 , \20132 );
and \U$19757 ( \20134 , \20126 , \20133 );
and \U$19758 ( \20135 , \20118 , \20125 );
or \U$19759 ( \20136 , \20134 , \20135 );
and \U$19760 ( \20137 , \7633 , RIae75a88_21);
and \U$19761 ( \20138 , RIae75998_19, \7631 );
nor \U$19762 ( \20139 , \20137 , \20138 );
and \U$19763 ( \20140 , \20139 , \7205 );
not \U$19764 ( \20141 , \20139 );
and \U$19765 ( \20142 , \20141 , \7206 );
nor \U$19766 ( \20143 , \20140 , \20142 );
not \U$19767 ( \20144 , \20143 );
and \U$19768 ( \20145 , \8966 , RIae75e48_29);
and \U$19769 ( \20146 , RIae75c68_25, \8964 );
nor \U$19770 ( \20147 , \20145 , \20146 );
and \U$19771 ( \20148 , \20147 , \8789 );
not \U$19772 ( \20149 , \20147 );
and \U$19773 ( \20150 , \20149 , \8799 );
nor \U$19774 ( \20151 , \20148 , \20150 );
not \U$19775 ( \20152 , \20151 );
and \U$19776 ( \20153 , \20144 , \20152 );
and \U$19777 ( \20154 , \20151 , \20143 );
and \U$19778 ( \20155 , \8371 , RIae758a8_17);
and \U$19779 ( \20156 , RIae75f38_31, \8369 );
nor \U$19780 ( \20157 , \20155 , \20156 );
and \U$19781 ( \20158 , \20157 , \8019 );
not \U$19782 ( \20159 , \20157 );
and \U$19783 ( \20160 , \20159 , \8020 );
nor \U$19784 ( \20161 , \20158 , \20160 );
nor \U$19785 ( \20162 , \20154 , \20161 );
nor \U$19786 ( \20163 , \20153 , \20162 );
or \U$19787 ( \20164 , \20136 , \20163 );
not \U$19788 ( \20165 , \20136 );
not \U$19789 ( \20166 , \20163 );
or \U$19790 ( \20167 , \20165 , \20166 );
and \U$19791 ( \20168 , \5896 , RIae77e28_97);
and \U$19792 ( \20169 , RIae78968_121, \5894 );
nor \U$19793 ( \20170 , \20168 , \20169 );
and \U$19794 ( \20171 , \20170 , \5590 );
not \U$19795 ( \20172 , \20170 );
and \U$19796 ( \20173 , \20172 , \5589 );
nor \U$19797 ( \20174 , \20171 , \20173 );
and \U$19798 ( \20175 , \6172 , RIae78878_119);
and \U$19799 ( \20176 , RIae78788_117, \6170 );
nor \U$19800 ( \20177 , \20175 , \20176 );
and \U$19801 ( \20178 , \20177 , \6176 );
not \U$19802 ( \20179 , \20177 );
and \U$19803 ( \20180 , \20179 , \6175 );
nor \U$19804 ( \20181 , \20178 , \20180 );
xor \U$19805 ( \20182 , \20174 , \20181 );
and \U$19806 ( \20183 , \6941 , RIae78698_115);
and \U$19807 ( \20184 , RIae75b78_23, \6939 );
nor \U$19808 ( \20185 , \20183 , \20184 );
and \U$19809 ( \20186 , \20185 , \6314 );
not \U$19810 ( \20187 , \20185 );
and \U$19811 ( \20188 , \20187 , \6945 );
nor \U$19812 ( \20189 , \20186 , \20188 );
and \U$19813 ( \20190 , \20182 , \20189 );
and \U$19814 ( \20191 , \20174 , \20181 );
or \U$19815 ( \20192 , \20190 , \20191 );
nand \U$19816 ( \20193 , \20167 , \20192 );
nand \U$19817 ( \20194 , \20164 , \20193 );
and \U$19818 ( \20195 , \12180 , RIae75128_1);
and \U$19819 ( \20196 , RIae75308_5, \12178 );
nor \U$19820 ( \20197 , \20195 , \20196 );
and \U$19821 ( \20198 , \20197 , \12184 );
not \U$19822 ( \20199 , \20197 );
and \U$19823 ( \20200 , \20199 , \11827 );
nor \U$19824 ( \20201 , \20198 , \20200 );
and \U$19825 ( \20202 , \13059 , RIae753f8_7);
and \U$19826 ( \20203 , RIae763e8_41, \13057 );
nor \U$19827 ( \20204 , \20202 , \20203 );
and \U$19828 ( \20205 , \20204 , \13063 );
not \U$19829 ( \20206 , \20204 );
and \U$19830 ( \20207 , \20206 , \12718 );
nor \U$19831 ( \20208 , \20205 , \20207 );
xor \U$19832 ( \20209 , \20201 , \20208 );
and \U$19833 ( \20210 , \14059 , RIae764d8_43);
and \U$19834 ( \20211 , RIae766b8_47, \14057 );
nor \U$19835 ( \20212 , \20210 , \20211 );
and \U$19836 ( \20213 , \20212 , \13502 );
not \U$19837 ( \20214 , \20212 );
and \U$19838 ( \20215 , \20214 , \14063 );
nor \U$19839 ( \20216 , \20213 , \20215 );
and \U$19840 ( \20217 , \20209 , \20216 );
and \U$19841 ( \20218 , \20201 , \20208 );
or \U$19842 ( \20219 , \20217 , \20218 );
and \U$19843 ( \20220 , \15726 , RIae76028_33);
and \U$19844 ( \20221 , RIae7aab0_192, RIae762f8_39);
nor \U$19845 ( \20222 , \20220 , \20221 );
and \U$19846 ( \20223 , \20222 , \14959 );
not \U$19847 ( \20224 , \20222 );
and \U$19848 ( \20225 , \20224 , RIae7aa38_191);
nor \U$19849 ( \20226 , \20223 , \20225 );
xor \U$19850 ( \20227 , \20226 , \587 );
and \U$19851 ( \20228 , \14964 , RIae765c8_45);
and \U$19852 ( \20229 , RIae76118_35, \14962 );
nor \U$19853 ( \20230 , \20228 , \20229 );
and \U$19854 ( \20231 , \20230 , \14463 );
not \U$19855 ( \20232 , \20230 );
and \U$19856 ( \20233 , \20232 , \14462 );
nor \U$19857 ( \20234 , \20231 , \20233 );
and \U$19858 ( \20235 , \20227 , \20234 );
and \U$19859 ( \20236 , \20226 , \587 );
or \U$19860 ( \20237 , \20235 , \20236 );
xor \U$19861 ( \20238 , \20219 , \20237 );
and \U$19862 ( \20239 , \9760 , RIae75d58_27);
and \U$19863 ( \20240 , RIae755d8_11, \9758 );
nor \U$19864 ( \20241 , \20239 , \20240 );
and \U$19865 ( \20242 , \20241 , \9273 );
not \U$19866 ( \20243 , \20241 );
and \U$19867 ( \20244 , \20243 , \9764 );
nor \U$19868 ( \20245 , \20242 , \20244 );
and \U$19869 ( \20246 , \10548 , RIae754e8_9);
and \U$19870 ( \20247 , RIae757b8_15, \10546 );
nor \U$19871 ( \20248 , \20246 , \20247 );
and \U$19872 ( \20249 , \20248 , \10421 );
not \U$19873 ( \20250 , \20248 );
and \U$19874 ( \20251 , \20250 , \10118 );
nor \U$19875 ( \20252 , \20249 , \20251 );
xor \U$19876 ( \20253 , \20245 , \20252 );
and \U$19877 ( \20254 , \11470 , RIae756c8_13);
and \U$19878 ( \20255 , RIae75218_3, \11468 );
nor \U$19879 ( \20256 , \20254 , \20255 );
and \U$19880 ( \20257 , \20256 , \10936 );
not \U$19881 ( \20258 , \20256 );
and \U$19882 ( \20259 , \20258 , \11474 );
nor \U$19883 ( \20260 , \20257 , \20259 );
and \U$19884 ( \20261 , \20253 , \20260 );
and \U$19885 ( \20262 , \20245 , \20252 );
or \U$19886 ( \20263 , \20261 , \20262 );
and \U$19887 ( \20264 , \20238 , \20263 );
and \U$19888 ( \20265 , \20219 , \20237 );
or \U$19889 ( \20266 , \20264 , \20265 );
xor \U$19890 ( \20267 , \20194 , \20266 );
and \U$19891 ( \20268 , \1138 , RIae773d8_75);
and \U$19892 ( \20269 , RIae77a68_89, \1136 );
nor \U$19893 ( \20270 , \20268 , \20269 );
and \U$19894 ( \20271 , \20270 , \1142 );
not \U$19895 ( \20272 , \20270 );
and \U$19896 ( \20273 , \20272 , \1012 );
nor \U$19897 ( \20274 , \20271 , \20273 );
not \U$19898 ( \20275 , \20274 );
and \U$19899 ( \20276 , \1593 , RIae77888_85);
and \U$19900 ( \20277 , RIae76f28_65, \1591 );
nor \U$19901 ( \20278 , \20276 , \20277 );
and \U$19902 ( \20279 , \20278 , \1488 );
not \U$19903 ( \20280 , \20278 );
and \U$19904 ( \20281 , \20280 , \1498 );
nor \U$19905 ( \20282 , \20279 , \20281 );
not \U$19906 ( \20283 , \20282 );
and \U$19907 ( \20284 , \20275 , \20283 );
and \U$19908 ( \20285 , \20282 , \20274 );
and \U$19909 ( \20286 , \1376 , RIae77978_87);
and \U$19910 ( \20287 , RIae77798_83, \1374 );
nor \U$19911 ( \20288 , \20286 , \20287 );
and \U$19912 ( \20289 , \20288 , \1261 );
not \U$19913 ( \20290 , \20288 );
and \U$19914 ( \20291 , \20290 , \1380 );
nor \U$19915 ( \20292 , \20289 , \20291 );
nor \U$19916 ( \20293 , \20285 , \20292 );
nor \U$19917 ( \20294 , \20284 , \20293 );
and \U$19918 ( \20295 , \3214 , RIae780f8_103);
and \U$19919 ( \20296 , RIae77f18_99, \3212 );
nor \U$19920 ( \20297 , \20295 , \20296 );
not \U$19921 ( \20298 , \20297 );
not \U$19922 ( \20299 , \2774 );
and \U$19923 ( \20300 , \20298 , \20299 );
and \U$19924 ( \20301 , \20297 , \3218 );
nor \U$19925 ( \20302 , \20300 , \20301 );
and \U$19926 ( \20303 , \2783 , RIae772e8_73);
and \U$19927 ( \20304 , RIae782d8_107, \2781 );
nor \U$19928 ( \20305 , \20303 , \20304 );
not \U$19929 ( \20306 , \20305 );
not \U$19930 ( \20307 , \3089 );
and \U$19931 ( \20308 , \20306 , \20307 );
and \U$19932 ( \20309 , \20305 , \3089 );
nor \U$19933 ( \20310 , \20308 , \20309 );
xor \U$19934 ( \20311 , \20302 , \20310 );
and \U$19935 ( \20312 , \3730 , RIae78008_101);
and \U$19936 ( \20313 , RIae781e8_105, \3728 );
nor \U$19937 ( \20314 , \20312 , \20313 );
and \U$19938 ( \20315 , \20314 , \3422 );
not \U$19939 ( \20316 , \20314 );
and \U$19940 ( \20317 , \20316 , \3732 );
nor \U$19941 ( \20318 , \20315 , \20317 );
and \U$19942 ( \20319 , \20311 , \20318 );
and \U$19943 ( \20320 , \20302 , \20310 );
or \U$19944 ( \20321 , \20319 , \20320 );
xor \U$19945 ( \20322 , \20294 , \20321 );
and \U$19946 ( \20323 , \2224 , RIae76c58_59);
and \U$19947 ( \20324 , RIae77180_70, \2222 );
nor \U$19948 ( \20325 , \20323 , \20324 );
and \U$19949 ( \20326 , \20325 , \2060 );
not \U$19950 ( \20327 , \20325 );
and \U$19951 ( \20328 , \20327 , \2061 );
nor \U$19952 ( \20329 , \20326 , \20328 );
and \U$19953 ( \20330 , \1939 , RIae76e38_63);
and \U$19954 ( \20331 , RIae76d48_61, \1937 );
nor \U$19955 ( \20332 , \20330 , \20331 );
and \U$19956 ( \20333 , \20332 , \1734 );
not \U$19957 ( \20334 , \20332 );
and \U$19958 ( \20335 , \20334 , \1735 );
nor \U$19959 ( \20336 , \20333 , \20335 );
xor \U$19960 ( \20337 , \20329 , \20336 );
and \U$19961 ( \20338 , \2607 , RIae77018_67);
and \U$19962 ( \20339 , RIae771f8_71, \2605 );
nor \U$19963 ( \20340 , \20338 , \20339 );
and \U$19964 ( \20341 , \20340 , \2397 );
not \U$19965 ( \20342 , \20340 );
and \U$19966 ( \20343 , \20342 , \2611 );
nor \U$19967 ( \20344 , \20341 , \20343 );
and \U$19968 ( \20345 , \20337 , \20344 );
and \U$19969 ( \20346 , \20329 , \20336 );
or \U$19970 ( \20347 , \20345 , \20346 );
and \U$19971 ( \20348 , \20322 , \20347 );
and \U$19972 ( \20349 , \20294 , \20321 );
nor \U$19973 ( \20350 , \20348 , \20349 );
and \U$19974 ( \20351 , \20267 , \20350 );
and \U$19975 ( \20352 , \20194 , \20266 );
or \U$19976 ( \20353 , \20351 , \20352 );
xor \U$19977 ( \20354 , \20111 , \20353 );
xor \U$19978 ( \20355 , \19317 , \562 );
xor \U$19979 ( \20356 , \20355 , \19325 );
xor \U$19980 ( \20357 , \19620 , \19622 );
xor \U$19981 ( \20358 , \20357 , \19625 );
and \U$19982 ( \20359 , \20356 , \20358 );
xor \U$19983 ( \20360 , \19336 , \19343 );
xor \U$19984 ( \20361 , \20360 , \19351 );
xor \U$19985 ( \20362 , \19647 , \19652 );
xor \U$19986 ( \20363 , \20361 , \20362 );
xor \U$19987 ( \20364 , \19620 , \19622 );
xor \U$19988 ( \20365 , \20364 , \19625 );
and \U$19989 ( \20366 , \20363 , \20365 );
and \U$19990 ( \20367 , \20356 , \20363 );
or \U$19991 ( \20368 , \20359 , \20366 , \20367 );
and \U$19992 ( \20369 , \20354 , \20368 );
and \U$19993 ( \20370 , \20111 , \20353 );
nor \U$19994 ( \20371 , \20369 , \20370 );
nor \U$19995 ( \20372 , \20064 , \20371 );
nor \U$19996 ( \20373 , \20063 , \20372 );
not \U$19997 ( \20374 , \19595 );
not \U$19998 ( \20375 , \19567 );
or \U$19999 ( \20376 , \20374 , \20375 );
or \U$20000 ( \20377 , \19567 , \19595 );
nand \U$20001 ( \20378 , \20376 , \20377 );
not \U$20002 ( \20379 , \20378 );
not \U$20003 ( \20380 , \19577 );
and \U$20004 ( \20381 , \20379 , \20380 );
and \U$20005 ( \20382 , \20378 , \19577 );
nor \U$20006 ( \20383 , \20381 , \20382 );
or \U$20007 ( \20384 , \20373 , \20383 );
not \U$20008 ( \20385 , \20383 );
not \U$20009 ( \20386 , \20373 );
or \U$20010 ( \20387 , \20385 , \20386 );
xor \U$20011 ( \20388 , \19660 , \19906 );
xor \U$20012 ( \20389 , \20388 , \19921 );
xor \U$20013 ( \20390 , \19608 , \19610 );
xor \U$20014 ( \20391 , \20390 , \19615 );
and \U$20015 ( \20392 , \20389 , \20391 );
xor \U$20016 ( \20393 , \19931 , \19943 );
xor \U$20017 ( \20394 , \20393 , \19948 );
xor \U$20018 ( \20395 , \19608 , \19610 );
xor \U$20019 ( \20396 , \20395 , \19615 );
and \U$20020 ( \20397 , \20394 , \20396 );
and \U$20021 ( \20398 , \20389 , \20394 );
or \U$20022 ( \20399 , \20392 , \20397 , \20398 );
nand \U$20023 ( \20400 , \20387 , \20399 );
nand \U$20024 ( \20401 , \20384 , \20400 );
and \U$20025 ( \20402 , \20015 , \20401 );
and \U$20026 ( \20403 , \20002 , \20014 );
nor \U$20027 ( \20404 , \20402 , \20403 );
nor \U$20028 ( \20405 , \20000 , \20404 );
and \U$20029 ( \20406 , \19997 , \20405 );
xor \U$20030 ( \20407 , \20405 , \19997 );
xor \U$20031 ( \20408 , \19767 , \19794 );
xor \U$20032 ( \20409 , \20408 , \19820 );
not \U$20033 ( \20410 , \20409 );
xor \U$20034 ( \20411 , \20294 , \20321 );
xor \U$20035 ( \20412 , \20411 , \20347 );
not \U$20036 ( \20413 , \20192 );
not \U$20037 ( \20414 , \20136 );
or \U$20038 ( \20415 , \20413 , \20414 );
or \U$20039 ( \20416 , \20136 , \20192 );
nand \U$20040 ( \20417 , \20415 , \20416 );
not \U$20041 ( \20418 , \20417 );
not \U$20042 ( \20419 , \20163 );
and \U$20043 ( \20420 , \20418 , \20419 );
and \U$20044 ( \20421 , \20417 , \20163 );
nor \U$20045 ( \20422 , \20420 , \20421 );
xor \U$20046 ( \20423 , \20412 , \20422 );
not \U$20047 ( \20424 , \20083 );
not \U$20048 ( \20425 , \20089 );
or \U$20049 ( \20426 , \20424 , \20425 );
or \U$20050 ( \20427 , \20089 , \20083 );
nand \U$20051 ( \20428 , \20426 , \20427 );
not \U$20052 ( \20429 , \20428 );
not \U$20053 ( \20430 , \20076 );
and \U$20054 ( \20431 , \20429 , \20430 );
and \U$20055 ( \20432 , \20428 , \20076 );
nor \U$20056 ( \20433 , \20431 , \20432 );
and \U$20057 ( \20434 , \20423 , \20433 );
and \U$20058 ( \20435 , \20412 , \20422 );
nor \U$20059 ( \20436 , \20434 , \20435 );
not \U$20060 ( \20437 , \20436 );
or \U$20061 ( \20438 , \20410 , \20437 );
or \U$20062 ( \20439 , \20436 , \20409 );
nand \U$20063 ( \20440 , \20438 , \20439 );
not \U$20064 ( \20441 , \20440 );
xor \U$20065 ( \20442 , \20043 , \20045 );
xor \U$20066 ( \20443 , \20442 , \20056 );
not \U$20067 ( \20444 , \20443 );
and \U$20068 ( \20445 , \20441 , \20444 );
and \U$20069 ( \20446 , \20440 , \20443 );
nor \U$20070 ( \20447 , \20445 , \20446 );
and \U$20071 ( \20448 , \4247 , RIae781e8_105);
and \U$20072 ( \20449 , RIae785a8_113, \4245 );
nor \U$20073 ( \20450 , \20448 , \20449 );
and \U$20074 ( \20451 , \20450 , \3989 );
not \U$20075 ( \20452 , \20450 );
and \U$20076 ( \20453 , \20452 , \4251 );
nor \U$20077 ( \20454 , \20451 , \20453 );
and \U$20078 ( \20455 , \4688 , RIae783c8_109);
and \U$20079 ( \20456 , RIae78530_112, \4686 );
nor \U$20080 ( \20457 , \20455 , \20456 );
and \U$20081 ( \20458 , \20457 , \4481 );
not \U$20082 ( \20459 , \20457 );
and \U$20083 ( \20460 , \20459 , \4482 );
nor \U$20084 ( \20461 , \20458 , \20460 );
xor \U$20085 ( \20462 , \20454 , \20461 );
and \U$20086 ( \20463 , \3730 , RIae77f18_99);
and \U$20087 ( \20464 , RIae78008_101, \3728 );
nor \U$20088 ( \20465 , \20463 , \20464 );
and \U$20089 ( \20466 , \20465 , \3732 );
not \U$20090 ( \20467 , \20465 );
and \U$20091 ( \20468 , \20467 , \3422 );
nor \U$20092 ( \20469 , \20466 , \20468 );
and \U$20093 ( \20470 , \20462 , \20469 );
and \U$20094 ( \20471 , \20454 , \20461 );
nor \U$20095 ( \20472 , \20470 , \20471 );
not \U$20096 ( \20473 , \20472 );
and \U$20097 ( \20474 , \7633 , RIae75b78_23);
and \U$20098 ( \20475 , RIae75a88_21, \7631 );
nor \U$20099 ( \20476 , \20474 , \20475 );
and \U$20100 ( \20477 , \20476 , \7206 );
not \U$20101 ( \20478 , \20476 );
and \U$20102 ( \20479 , \20478 , \7205 );
nor \U$20103 ( \20480 , \20477 , \20479 );
and \U$20104 ( \20481 , \8371 , RIae75998_19);
and \U$20105 ( \20482 , RIae758a8_17, \8369 );
nor \U$20106 ( \20483 , \20481 , \20482 );
and \U$20107 ( \20484 , \20483 , \8020 );
not \U$20108 ( \20485 , \20483 );
and \U$20109 ( \20486 , \20485 , \8019 );
nor \U$20110 ( \20487 , \20484 , \20486 );
xor \U$20111 ( \20488 , \20480 , \20487 );
and \U$20112 ( \20489 , \6941 , RIae78788_117);
and \U$20113 ( \20490 , RIae78698_115, \6939 );
nor \U$20114 ( \20491 , \20489 , \20490 );
and \U$20115 ( \20492 , \20491 , \6314 );
not \U$20116 ( \20493 , \20491 );
and \U$20117 ( \20494 , \20493 , \6945 );
nor \U$20118 ( \20495 , \20492 , \20494 );
and \U$20119 ( \20496 , \20488 , \20495 );
and \U$20120 ( \20497 , \20480 , \20487 );
nor \U$20121 ( \20498 , \20496 , \20497 );
not \U$20122 ( \20499 , \20498 );
and \U$20123 ( \20500 , \20473 , \20499 );
and \U$20124 ( \20501 , \20472 , \20498 );
and \U$20125 ( \20502 , \5399 , RIae77c48_93);
and \U$20126 ( \20503 , RIae77b58_91, \5397 );
nor \U$20127 ( \20504 , \20502 , \20503 );
and \U$20128 ( \20505 , \20504 , \5403 );
not \U$20129 ( \20506 , \20504 );
and \U$20130 ( \20507 , \20506 , \5016 );
nor \U$20131 ( \20508 , \20505 , \20507 );
not \U$20132 ( \20509 , \20508 );
and \U$20133 ( \20510 , \5896 , RIae77d38_95);
and \U$20134 ( \20511 , RIae77e28_97, \5894 );
nor \U$20135 ( \20512 , \20510 , \20511 );
and \U$20136 ( \20513 , \20512 , \5589 );
not \U$20137 ( \20514 , \20512 );
and \U$20138 ( \20515 , \20514 , \5590 );
nor \U$20139 ( \20516 , \20513 , \20515 );
not \U$20140 ( \20517 , \20516 );
and \U$20141 ( \20518 , \20509 , \20517 );
and \U$20142 ( \20519 , \20516 , \20508 );
and \U$20143 ( \20520 , \6172 , RIae78968_121);
and \U$20144 ( \20521 , RIae78878_119, \6170 );
nor \U$20145 ( \20522 , \20520 , \20521 );
and \U$20146 ( \20523 , \20522 , \6175 );
not \U$20147 ( \20524 , \20522 );
and \U$20148 ( \20525 , \20524 , \6176 );
nor \U$20149 ( \20526 , \20523 , \20525 );
nor \U$20150 ( \20527 , \20519 , \20526 );
nor \U$20151 ( \20528 , \20518 , \20527 );
nor \U$20152 ( \20529 , \20501 , \20528 );
nor \U$20153 ( \20530 , \20500 , \20529 );
and \U$20154 ( \20531 , \2607 , RIae77180_70);
and \U$20155 ( \20532 , RIae77018_67, \2605 );
nor \U$20156 ( \20533 , \20531 , \20532 );
and \U$20157 ( \20534 , \20533 , \2611 );
not \U$20158 ( \20535 , \20533 );
and \U$20159 ( \20536 , \20535 , \2397 );
nor \U$20160 ( \20537 , \20534 , \20536 );
not \U$20161 ( \20538 , \3089 );
and \U$20162 ( \20539 , \2783 , RIae771f8_71);
and \U$20163 ( \20540 , RIae772e8_73, \2781 );
nor \U$20164 ( \20541 , \20539 , \20540 );
not \U$20165 ( \20542 , \20541 );
or \U$20166 ( \20543 , \20538 , \20542 );
or \U$20167 ( \20544 , \20541 , \3089 );
nand \U$20168 ( \20545 , \20543 , \20544 );
xor \U$20169 ( \20546 , \20537 , \20545 );
not \U$20170 ( \20547 , \3218 );
and \U$20171 ( \20548 , \3214 , RIae782d8_107);
and \U$20172 ( \20549 , RIae780f8_103, \3212 );
nor \U$20173 ( \20550 , \20548 , \20549 );
not \U$20174 ( \20551 , \20550 );
or \U$20175 ( \20552 , \20547 , \20551 );
or \U$20176 ( \20553 , \20550 , \2774 );
nand \U$20177 ( \20554 , \20552 , \20553 );
and \U$20178 ( \20555 , \20546 , \20554 );
and \U$20179 ( \20556 , \20537 , \20545 );
or \U$20180 ( \20557 , \20555 , \20556 );
and \U$20181 ( \20558 , \1138 , RIae77720_82);
and \U$20182 ( \20559 , RIae773d8_75, \1136 );
nor \U$20183 ( \20560 , \20558 , \20559 );
and \U$20184 ( \20561 , \20560 , \1012 );
not \U$20185 ( \20562 , \20560 );
and \U$20186 ( \20563 , \20562 , \1142 );
nor \U$20187 ( \20564 , \20561 , \20563 );
not \U$20188 ( \20565 , \787 );
and \U$20189 ( \20566 , \883 , RIae775b8_79);
and \U$20190 ( \20567 , RIae774c8_77, \881 );
nor \U$20191 ( \20568 , \20566 , \20567 );
not \U$20192 ( \20569 , \20568 );
or \U$20193 ( \20570 , \20565 , \20569 );
or \U$20194 ( \20571 , \20568 , \789 );
nand \U$20195 ( \20572 , \20570 , \20571 );
xor \U$20196 ( \20573 , \20564 , \20572 );
and \U$20197 ( \20574 , \1376 , RIae77a68_89);
and \U$20198 ( \20575 , RIae77978_87, \1374 );
nor \U$20199 ( \20576 , \20574 , \20575 );
and \U$20200 ( \20577 , \20576 , \1380 );
not \U$20201 ( \20578 , \20576 );
and \U$20202 ( \20579 , \20578 , \1261 );
nor \U$20203 ( \20580 , \20577 , \20579 );
and \U$20204 ( \20581 , \20573 , \20580 );
and \U$20205 ( \20582 , \20564 , \20572 );
or \U$20206 ( \20583 , \20581 , \20582 );
xor \U$20207 ( \20584 , \20557 , \20583 );
and \U$20208 ( \20585 , \1939 , RIae76f28_65);
and \U$20209 ( \20586 , RIae76e38_63, \1937 );
nor \U$20210 ( \20587 , \20585 , \20586 );
and \U$20211 ( \20588 , \20587 , \1735 );
not \U$20212 ( \20589 , \20587 );
and \U$20213 ( \20590 , \20589 , \1734 );
nor \U$20214 ( \20591 , \20588 , \20590 );
and \U$20215 ( \20592 , \1593 , RIae77798_83);
and \U$20216 ( \20593 , RIae77888_85, \1591 );
nor \U$20217 ( \20594 , \20592 , \20593 );
and \U$20218 ( \20595 , \20594 , \1498 );
not \U$20219 ( \20596 , \20594 );
and \U$20220 ( \20597 , \20596 , \1488 );
nor \U$20221 ( \20598 , \20595 , \20597 );
xor \U$20222 ( \20599 , \20591 , \20598 );
and \U$20223 ( \20600 , \2224 , RIae76d48_61);
and \U$20224 ( \20601 , RIae76c58_59, \2222 );
nor \U$20225 ( \20602 , \20600 , \20601 );
and \U$20226 ( \20603 , \20602 , \2061 );
not \U$20227 ( \20604 , \20602 );
and \U$20228 ( \20605 , \20604 , \2060 );
nor \U$20229 ( \20606 , \20603 , \20605 );
and \U$20230 ( \20607 , \20599 , \20606 );
and \U$20231 ( \20608 , \20591 , \20598 );
or \U$20232 ( \20609 , \20607 , \20608 );
and \U$20233 ( \20610 , \20584 , \20609 );
and \U$20234 ( \20611 , \20557 , \20583 );
nor \U$20235 ( \20612 , \20610 , \20611 );
xor \U$20236 ( \20613 , \20530 , \20612 );
and \U$20237 ( \20614 , \13059 , RIae75308_5);
and \U$20238 ( \20615 , RIae753f8_7, \13057 );
nor \U$20239 ( \20616 , \20614 , \20615 );
and \U$20240 ( \20617 , \20616 , \13063 );
not \U$20241 ( \20618 , \20616 );
and \U$20242 ( \20619 , \20618 , \12718 );
nor \U$20243 ( \20620 , \20617 , \20619 );
and \U$20244 ( \20621 , \11470 , RIae757b8_15);
and \U$20245 ( \20622 , RIae756c8_13, \11468 );
nor \U$20246 ( \20623 , \20621 , \20622 );
and \U$20247 ( \20624 , \20623 , \10936 );
not \U$20248 ( \20625 , \20623 );
and \U$20249 ( \20626 , \20625 , \11474 );
nor \U$20250 ( \20627 , \20624 , \20626 );
xor \U$20251 ( \20628 , \20620 , \20627 );
and \U$20252 ( \20629 , \12180 , RIae75218_3);
and \U$20253 ( \20630 , RIae75128_1, \12178 );
nor \U$20254 ( \20631 , \20629 , \20630 );
and \U$20255 ( \20632 , \20631 , \12184 );
not \U$20256 ( \20633 , \20631 );
and \U$20257 ( \20634 , \20633 , \11827 );
nor \U$20258 ( \20635 , \20632 , \20634 );
and \U$20259 ( \20636 , \20628 , \20635 );
and \U$20260 ( \20637 , \20620 , \20627 );
or \U$20261 ( \20638 , \20636 , \20637 );
and \U$20262 ( \20639 , \8966 , RIae75f38_31);
and \U$20263 ( \20640 , RIae75e48_29, \8964 );
nor \U$20264 ( \20641 , \20639 , \20640 );
and \U$20265 ( \20642 , \20641 , \8799 );
not \U$20266 ( \20643 , \20641 );
and \U$20267 ( \20644 , \20643 , \8789 );
nor \U$20268 ( \20645 , \20642 , \20644 );
and \U$20269 ( \20646 , \9760 , RIae75c68_25);
and \U$20270 ( \20647 , RIae75d58_27, \9758 );
nor \U$20271 ( \20648 , \20646 , \20647 );
and \U$20272 ( \20649 , \20648 , \9273 );
not \U$20273 ( \20650 , \20648 );
and \U$20274 ( \20651 , \20650 , \9272 );
nor \U$20275 ( \20652 , \20649 , \20651 );
xor \U$20276 ( \20653 , \20645 , \20652 );
and \U$20277 ( \20654 , \10548 , RIae755d8_11);
and \U$20278 ( \20655 , RIae754e8_9, \10546 );
nor \U$20279 ( \20656 , \20654 , \20655 );
and \U$20280 ( \20657 , \20656 , \10421 );
not \U$20281 ( \20658 , \20656 );
and \U$20282 ( \20659 , \20658 , \10118 );
nor \U$20283 ( \20660 , \20657 , \20659 );
and \U$20284 ( \20661 , \20653 , \20660 );
and \U$20285 ( \20662 , \20645 , \20652 );
or \U$20286 ( \20663 , \20661 , \20662 );
xor \U$20287 ( \20664 , \20638 , \20663 );
and \U$20288 ( \20665 , \14964 , RIae766b8_47);
and \U$20289 ( \20666 , RIae765c8_45, \14962 );
nor \U$20290 ( \20667 , \20665 , \20666 );
and \U$20291 ( \20668 , \20667 , \14463 );
not \U$20292 ( \20669 , \20667 );
and \U$20293 ( \20670 , \20669 , \14462 );
nor \U$20294 ( \20671 , \20668 , \20670 );
and \U$20295 ( \20672 , \15726 , RIae76118_35);
and \U$20296 ( \20673 , RIae7aab0_192, RIae76028_33);
nor \U$20297 ( \20674 , \20672 , \20673 );
and \U$20298 ( \20675 , \20674 , \14959 );
not \U$20299 ( \20676 , \20674 );
and \U$20300 ( \20677 , \20676 , RIae7aa38_191);
nor \U$20301 ( \20678 , \20675 , \20677 );
xor \U$20302 ( \20679 , \20671 , \20678 );
and \U$20303 ( \20680 , \14059 , RIae763e8_41);
and \U$20304 ( \20681 , RIae764d8_43, \14057 );
nor \U$20305 ( \20682 , \20680 , \20681 );
and \U$20306 ( \20683 , \20682 , \13502 );
not \U$20307 ( \20684 , \20682 );
and \U$20308 ( \20685 , \20684 , \14063 );
nor \U$20309 ( \20686 , \20683 , \20685 );
and \U$20310 ( \20687 , \20679 , \20686 );
and \U$20311 ( \20688 , \20671 , \20678 );
or \U$20312 ( \20689 , \20687 , \20688 );
and \U$20313 ( \20690 , \20664 , \20689 );
and \U$20314 ( \20691 , \20638 , \20663 );
nor \U$20315 ( \20692 , \20690 , \20691 );
and \U$20316 ( \20693 , \20613 , \20692 );
and \U$20317 ( \20694 , \20530 , \20612 );
or \U$20318 ( \20695 , \20693 , \20694 );
xor \U$20319 ( \20696 , \20329 , \20336 );
xor \U$20320 ( \20697 , \20696 , \20344 );
not \U$20321 ( \20698 , \20697 );
xor \U$20322 ( \20699 , \20118 , \20125 );
xor \U$20323 ( \20700 , \20699 , \20133 );
not \U$20324 ( \20701 , \20700 );
and \U$20325 ( \20702 , \20698 , \20701 );
and \U$20326 ( \20703 , \20700 , \20697 );
xor \U$20327 ( \20704 , \20302 , \20310 );
xor \U$20328 ( \20705 , \20704 , \20318 );
nor \U$20329 ( \20706 , \20703 , \20705 );
nor \U$20330 ( \20707 , \20702 , \20706 );
nand \U$20331 ( \20708 , RIae775b8_79, \670 );
and \U$20332 ( \20709 , \20708 , \588 );
not \U$20333 ( \20710 , \20708 );
and \U$20334 ( \20711 , \20710 , \587 );
nor \U$20335 ( \20712 , \20709 , \20711 );
not \U$20336 ( \20713 , \787 );
and \U$20337 ( \20714 , \883 , RIae774c8_77);
and \U$20338 ( \20715 , RIae77720_82, \881 );
nor \U$20339 ( \20716 , \20714 , \20715 );
not \U$20340 ( \20717 , \20716 );
or \U$20341 ( \20718 , \20713 , \20717 );
or \U$20342 ( \20719 , \20716 , \789 );
nand \U$20343 ( \20720 , \20718 , \20719 );
xor \U$20344 ( \20721 , \20712 , \20720 );
not \U$20345 ( \20722 , \20274 );
xor \U$20346 ( \20723 , \20292 , \20282 );
not \U$20347 ( \20724 , \20723 );
or \U$20348 ( \20725 , \20722 , \20724 );
or \U$20349 ( \20726 , \20723 , \20274 );
nand \U$20350 ( \20727 , \20725 , \20726 );
and \U$20351 ( \20728 , \20721 , \20727 );
and \U$20352 ( \20729 , \20712 , \20720 );
nor \U$20353 ( \20730 , \20728 , \20729 );
xor \U$20354 ( \20731 , \20707 , \20730 );
xor \U$20355 ( \20732 , \20245 , \20252 );
xor \U$20356 ( \20733 , \20732 , \20260 );
xor \U$20357 ( \20734 , \20174 , \20181 );
xor \U$20358 ( \20735 , \20734 , \20189 );
and \U$20359 ( \20736 , \20733 , \20735 );
not \U$20360 ( \20737 , \20143 );
xor \U$20361 ( \20738 , \20161 , \20151 );
not \U$20362 ( \20739 , \20738 );
or \U$20363 ( \20740 , \20737 , \20739 );
or \U$20364 ( \20741 , \20738 , \20143 );
nand \U$20365 ( \20742 , \20740 , \20741 );
xor \U$20366 ( \20743 , \20174 , \20181 );
xor \U$20367 ( \20744 , \20743 , \20189 );
and \U$20368 ( \20745 , \20742 , \20744 );
and \U$20369 ( \20746 , \20733 , \20742 );
or \U$20370 ( \20747 , \20736 , \20745 , \20746 );
not \U$20371 ( \20748 , \20747 );
and \U$20372 ( \20749 , \20731 , \20748 );
and \U$20373 ( \20750 , \20707 , \20730 );
or \U$20374 ( \20751 , \20749 , \20750 );
xor \U$20375 ( \20752 , \20695 , \20751 );
xor \U$20376 ( \20753 , \20066 , \20068 );
xor \U$20377 ( \20754 , \20753 , \20071 );
xor \U$20378 ( \20755 , \19749 , \19756 );
xor \U$20379 ( \20756 , \20755 , \19764 );
xor \U$20380 ( \20757 , \20754 , \20756 );
not \U$20381 ( \20758 , \20094 );
not \U$20382 ( \20759 , \20106 );
or \U$20383 ( \20760 , \20758 , \20759 );
or \U$20384 ( \20761 , \20094 , \20106 );
nand \U$20385 ( \20762 , \20760 , \20761 );
not \U$20386 ( \20763 , \20762 );
not \U$20387 ( \20764 , \20096 );
and \U$20388 ( \20765 , \20763 , \20764 );
and \U$20389 ( \20766 , \20762 , \20096 );
nor \U$20390 ( \20767 , \20765 , \20766 );
and \U$20391 ( \20768 , \20757 , \20767 );
and \U$20392 ( \20769 , \20754 , \20756 );
or \U$20393 ( \20770 , \20768 , \20769 );
xor \U$20394 ( \20771 , \20752 , \20770 );
or \U$20395 ( \20772 , \20447 , \20771 );
not \U$20396 ( \20773 , \20771 );
not \U$20397 ( \20774 , \20447 );
or \U$20398 ( \20775 , \20773 , \20774 );
xor \U$20399 ( \20776 , \20074 , \20091 );
xor \U$20400 ( \20777 , \20776 , \20108 );
xor \U$20401 ( \20778 , \20194 , \20266 );
xor \U$20402 ( \20779 , \20778 , \20350 );
xor \U$20403 ( \20780 , \19620 , \19622 );
xor \U$20404 ( \20781 , \20780 , \19625 );
xor \U$20405 ( \20782 , \20356 , \20363 );
xor \U$20406 ( \20783 , \20781 , \20782 );
xor \U$20407 ( \20784 , \20779 , \20783 );
xor \U$20408 ( \20785 , \20777 , \20784 );
nand \U$20409 ( \20786 , \20775 , \20785 );
nand \U$20410 ( \20787 , \20772 , \20786 );
and \U$20411 ( \20788 , \1939 , RIae77888_85);
and \U$20412 ( \20789 , RIae76f28_65, \1937 );
nor \U$20413 ( \20790 , \20788 , \20789 );
and \U$20414 ( \20791 , \20790 , \1735 );
not \U$20415 ( \20792 , \20790 );
and \U$20416 ( \20793 , \20792 , \1734 );
nor \U$20417 ( \20794 , \20791 , \20793 );
and \U$20418 ( \20795 , \2224 , RIae76e38_63);
and \U$20419 ( \20796 , RIae76d48_61, \2222 );
nor \U$20420 ( \20797 , \20795 , \20796 );
and \U$20421 ( \20798 , \20797 , \2061 );
not \U$20422 ( \20799 , \20797 );
and \U$20423 ( \20800 , \20799 , \2060 );
nor \U$20424 ( \20801 , \20798 , \20800 );
xor \U$20425 ( \20802 , \20794 , \20801 );
and \U$20426 ( \20803 , \2607 , RIae76c58_59);
and \U$20427 ( \20804 , RIae77180_70, \2605 );
nor \U$20428 ( \20805 , \20803 , \20804 );
and \U$20429 ( \20806 , \20805 , \2611 );
not \U$20430 ( \20807 , \20805 );
and \U$20431 ( \20808 , \20807 , \2396 );
nor \U$20432 ( \20809 , \20806 , \20808 );
and \U$20433 ( \20810 , \20802 , \20809 );
and \U$20434 ( \20811 , \20794 , \20801 );
or \U$20435 ( \20812 , \20810 , \20811 );
and \U$20436 ( \20813 , \1138 , RIae774c8_77);
and \U$20437 ( \20814 , RIae77720_82, \1136 );
nor \U$20438 ( \20815 , \20813 , \20814 );
and \U$20439 ( \20816 , \20815 , \1012 );
not \U$20440 ( \20817 , \20815 );
and \U$20441 ( \20818 , \20817 , \1142 );
nor \U$20442 ( \20819 , \20816 , \20818 );
and \U$20443 ( \20820 , \1376 , RIae773d8_75);
and \U$20444 ( \20821 , RIae77a68_89, \1374 );
nor \U$20445 ( \20822 , \20820 , \20821 );
and \U$20446 ( \20823 , \20822 , \1380 );
not \U$20447 ( \20824 , \20822 );
and \U$20448 ( \20825 , \20824 , \1261 );
nor \U$20449 ( \20826 , \20823 , \20825 );
xor \U$20450 ( \20827 , \20819 , \20826 );
and \U$20451 ( \20828 , \1593 , RIae77978_87);
and \U$20452 ( \20829 , RIae77798_83, \1591 );
nor \U$20453 ( \20830 , \20828 , \20829 );
and \U$20454 ( \20831 , \20830 , \1498 );
not \U$20455 ( \20832 , \20830 );
and \U$20456 ( \20833 , \20832 , \1488 );
nor \U$20457 ( \20834 , \20831 , \20833 );
and \U$20458 ( \20835 , \20827 , \20834 );
and \U$20459 ( \20836 , \20819 , \20826 );
or \U$20460 ( \20837 , \20835 , \20836 );
xor \U$20461 ( \20838 , \20812 , \20837 );
and \U$20462 ( \20839 , \3730 , RIae780f8_103);
and \U$20463 ( \20840 , RIae77f18_99, \3728 );
nor \U$20464 ( \20841 , \20839 , \20840 );
and \U$20465 ( \20842 , \20841 , \3732 );
not \U$20466 ( \20843 , \20841 );
and \U$20467 ( \20844 , \20843 , \3422 );
nor \U$20468 ( \20845 , \20842 , \20844 );
not \U$20469 ( \20846 , \2789 );
and \U$20470 ( \20847 , \2783 , RIae77018_67);
and \U$20471 ( \20848 , RIae771f8_71, \2781 );
nor \U$20472 ( \20849 , \20847 , \20848 );
not \U$20473 ( \20850 , \20849 );
or \U$20474 ( \20851 , \20846 , \20850 );
or \U$20475 ( \20852 , \20849 , \3089 );
nand \U$20476 ( \20853 , \20851 , \20852 );
xor \U$20477 ( \20854 , \20845 , \20853 );
not \U$20478 ( \20855 , \2774 );
and \U$20479 ( \20856 , \3214 , RIae772e8_73);
and \U$20480 ( \20857 , RIae782d8_107, \3212 );
nor \U$20481 ( \20858 , \20856 , \20857 );
not \U$20482 ( \20859 , \20858 );
or \U$20483 ( \20860 , \20855 , \20859 );
or \U$20484 ( \20861 , \20858 , \3218 );
nand \U$20485 ( \20862 , \20860 , \20861 );
and \U$20486 ( \20863 , \20854 , \20862 );
and \U$20487 ( \20864 , \20845 , \20853 );
or \U$20488 ( \20865 , \20863 , \20864 );
and \U$20489 ( \20866 , \20838 , \20865 );
and \U$20490 ( \20867 , \20812 , \20837 );
or \U$20491 ( \20868 , \20866 , \20867 );
and \U$20492 ( \20869 , \9760 , RIae75e48_29);
and \U$20493 ( \20870 , RIae75c68_25, \9758 );
nor \U$20494 ( \20871 , \20869 , \20870 );
and \U$20495 ( \20872 , \20871 , \9273 );
not \U$20496 ( \20873 , \20871 );
and \U$20497 ( \20874 , \20873 , \9764 );
nor \U$20498 ( \20875 , \20872 , \20874 );
and \U$20499 ( \20876 , \10548 , RIae75d58_27);
and \U$20500 ( \20877 , RIae755d8_11, \10546 );
nor \U$20501 ( \20878 , \20876 , \20877 );
and \U$20502 ( \20879 , \20878 , \10421 );
not \U$20503 ( \20880 , \20878 );
and \U$20504 ( \20881 , \20880 , \10118 );
nor \U$20505 ( \20882 , \20879 , \20881 );
xor \U$20506 ( \20883 , \20875 , \20882 );
and \U$20507 ( \20884 , \11470 , RIae754e8_9);
and \U$20508 ( \20885 , RIae757b8_15, \11468 );
nor \U$20509 ( \20886 , \20884 , \20885 );
and \U$20510 ( \20887 , \20886 , \10936 );
not \U$20511 ( \20888 , \20886 );
and \U$20512 ( \20889 , \20888 , \11474 );
nor \U$20513 ( \20890 , \20887 , \20889 );
and \U$20514 ( \20891 , \20883 , \20890 );
and \U$20515 ( \20892 , \20875 , \20882 );
or \U$20516 ( \20893 , \20891 , \20892 );
and \U$20517 ( \20894 , \15726 , RIae765c8_45);
and \U$20518 ( \20895 , RIae7aab0_192, RIae76118_35);
nor \U$20519 ( \20896 , \20894 , \20895 );
and \U$20520 ( \20897 , \20896 , \14959 );
not \U$20521 ( \20898 , \20896 );
and \U$20522 ( \20899 , \20898 , RIae7aa38_191);
nor \U$20523 ( \20900 , \20897 , \20899 );
xor \U$20524 ( \20901 , \20900 , \789 );
and \U$20525 ( \20902 , \14964 , RIae764d8_43);
and \U$20526 ( \20903 , RIae766b8_47, \14962 );
nor \U$20527 ( \20904 , \20902 , \20903 );
and \U$20528 ( \20905 , \20904 , \14463 );
not \U$20529 ( \20906 , \20904 );
and \U$20530 ( \20907 , \20906 , \14462 );
nor \U$20531 ( \20908 , \20905 , \20907 );
and \U$20532 ( \20909 , \20901 , \20908 );
and \U$20533 ( \20910 , \20900 , \789 );
or \U$20534 ( \20911 , \20909 , \20910 );
xor \U$20535 ( \20912 , \20893 , \20911 );
and \U$20536 ( \20913 , \14059 , RIae753f8_7);
and \U$20537 ( \20914 , RIae763e8_41, \14057 );
nor \U$20538 ( \20915 , \20913 , \20914 );
and \U$20539 ( \20916 , \20915 , \13502 );
not \U$20540 ( \20917 , \20915 );
and \U$20541 ( \20918 , \20917 , \14063 );
nor \U$20542 ( \20919 , \20916 , \20918 );
and \U$20543 ( \20920 , \12180 , RIae756c8_13);
and \U$20544 ( \20921 , RIae75218_3, \12178 );
nor \U$20545 ( \20922 , \20920 , \20921 );
and \U$20546 ( \20923 , \20922 , \12184 );
not \U$20547 ( \20924 , \20922 );
and \U$20548 ( \20925 , \20924 , \11827 );
nor \U$20549 ( \20926 , \20923 , \20925 );
xor \U$20550 ( \20927 , \20919 , \20926 );
and \U$20551 ( \20928 , \13059 , RIae75128_1);
and \U$20552 ( \20929 , RIae75308_5, \13057 );
nor \U$20553 ( \20930 , \20928 , \20929 );
and \U$20554 ( \20931 , \20930 , \13063 );
not \U$20555 ( \20932 , \20930 );
and \U$20556 ( \20933 , \20932 , \12718 );
nor \U$20557 ( \20934 , \20931 , \20933 );
and \U$20558 ( \20935 , \20927 , \20934 );
and \U$20559 ( \20936 , \20919 , \20926 );
or \U$20560 ( \20937 , \20935 , \20936 );
and \U$20561 ( \20938 , \20912 , \20937 );
and \U$20562 ( \20939 , \20893 , \20911 );
or \U$20563 ( \20940 , \20938 , \20939 );
xor \U$20564 ( \20941 , \20868 , \20940 );
and \U$20565 ( \20942 , \8371 , RIae75a88_21);
and \U$20566 ( \20943 , RIae75998_19, \8369 );
nor \U$20567 ( \20944 , \20942 , \20943 );
and \U$20568 ( \20945 , \20944 , \8020 );
not \U$20569 ( \20946 , \20944 );
and \U$20570 ( \20947 , \20946 , \8019 );
nor \U$20571 ( \20948 , \20945 , \20947 );
and \U$20572 ( \20949 , \7633 , RIae78698_115);
and \U$20573 ( \20950 , RIae75b78_23, \7631 );
nor \U$20574 ( \20951 , \20949 , \20950 );
and \U$20575 ( \20952 , \20951 , \7206 );
not \U$20576 ( \20953 , \20951 );
and \U$20577 ( \20954 , \20953 , \7205 );
nor \U$20578 ( \20955 , \20952 , \20954 );
xor \U$20579 ( \20956 , \20948 , \20955 );
and \U$20580 ( \20957 , \8966 , RIae758a8_17);
and \U$20581 ( \20958 , RIae75f38_31, \8964 );
nor \U$20582 ( \20959 , \20957 , \20958 );
and \U$20583 ( \20960 , \20959 , \8799 );
not \U$20584 ( \20961 , \20959 );
and \U$20585 ( \20962 , \20961 , \8789 );
nor \U$20586 ( \20963 , \20960 , \20962 );
and \U$20587 ( \20964 , \20956 , \20963 );
and \U$20588 ( \20965 , \20948 , \20955 );
or \U$20589 ( \20966 , \20964 , \20965 );
and \U$20590 ( \20967 , \5399 , RIae78530_112);
and \U$20591 ( \20968 , RIae77c48_93, \5397 );
nor \U$20592 ( \20969 , \20967 , \20968 );
and \U$20593 ( \20970 , \20969 , \5016 );
not \U$20594 ( \20971 , \20969 );
and \U$20595 ( \20972 , \20971 , \5403 );
nor \U$20596 ( \20973 , \20970 , \20972 );
and \U$20597 ( \20974 , \4247 , RIae78008_101);
and \U$20598 ( \20975 , RIae781e8_105, \4245 );
nor \U$20599 ( \20976 , \20974 , \20975 );
and \U$20600 ( \20977 , \20976 , \3989 );
not \U$20601 ( \20978 , \20976 );
and \U$20602 ( \20979 , \20978 , \4251 );
nor \U$20603 ( \20980 , \20977 , \20979 );
xor \U$20604 ( \20981 , \20973 , \20980 );
and \U$20605 ( \20982 , \4688 , RIae785a8_113);
and \U$20606 ( \20983 , RIae783c8_109, \4686 );
nor \U$20607 ( \20984 , \20982 , \20983 );
and \U$20608 ( \20985 , \20984 , \4481 );
not \U$20609 ( \20986 , \20984 );
and \U$20610 ( \20987 , \20986 , \4482 );
nor \U$20611 ( \20988 , \20985 , \20987 );
and \U$20612 ( \20989 , \20981 , \20988 );
and \U$20613 ( \20990 , \20973 , \20980 );
or \U$20614 ( \20991 , \20989 , \20990 );
xor \U$20615 ( \20992 , \20966 , \20991 );
and \U$20616 ( \20993 , \6941 , RIae78878_119);
and \U$20617 ( \20994 , RIae78788_117, \6939 );
nor \U$20618 ( \20995 , \20993 , \20994 );
and \U$20619 ( \20996 , \20995 , \6314 );
not \U$20620 ( \20997 , \20995 );
and \U$20621 ( \20998 , \20997 , \6945 );
nor \U$20622 ( \20999 , \20996 , \20998 );
and \U$20623 ( \21000 , \5896 , RIae77b58_91);
and \U$20624 ( \21001 , RIae77d38_95, \5894 );
nor \U$20625 ( \21002 , \21000 , \21001 );
and \U$20626 ( \21003 , \21002 , \5590 );
not \U$20627 ( \21004 , \21002 );
and \U$20628 ( \21005 , \21004 , \5589 );
nor \U$20629 ( \21006 , \21003 , \21005 );
xor \U$20630 ( \21007 , \20999 , \21006 );
and \U$20631 ( \21008 , \6172 , RIae77e28_97);
and \U$20632 ( \21009 , RIae78968_121, \6170 );
nor \U$20633 ( \21010 , \21008 , \21009 );
and \U$20634 ( \21011 , \21010 , \6176 );
not \U$20635 ( \21012 , \21010 );
and \U$20636 ( \21013 , \21012 , \6175 );
nor \U$20637 ( \21014 , \21011 , \21013 );
and \U$20638 ( \21015 , \21007 , \21014 );
and \U$20639 ( \21016 , \20999 , \21006 );
or \U$20640 ( \21017 , \21015 , \21016 );
and \U$20641 ( \21018 , \20992 , \21017 );
and \U$20642 ( \21019 , \20966 , \20991 );
or \U$20643 ( \21020 , \21018 , \21019 );
and \U$20644 ( \21021 , \20941 , \21020 );
and \U$20645 ( \21022 , \20868 , \20940 );
or \U$20646 ( \21023 , \21021 , \21022 );
xor \U$20647 ( \21024 , \20201 , \20208 );
xor \U$20648 ( \21025 , \21024 , \20216 );
xor \U$20649 ( \21026 , \20226 , \587 );
xor \U$20650 ( \21027 , \21026 , \20234 );
and \U$20651 ( \21028 , \21025 , \21027 );
xor \U$20652 ( \21029 , \20174 , \20181 );
xor \U$20653 ( \21030 , \21029 , \20189 );
xor \U$20654 ( \21031 , \20733 , \20742 );
xor \U$20655 ( \21032 , \21030 , \21031 );
xor \U$20656 ( \21033 , \20226 , \587 );
xor \U$20657 ( \21034 , \21033 , \20234 );
and \U$20658 ( \21035 , \21032 , \21034 );
and \U$20659 ( \21036 , \21025 , \21032 );
or \U$20660 ( \21037 , \21028 , \21035 , \21036 );
xor \U$20661 ( \21038 , \21023 , \21037 );
xor \U$20662 ( \21039 , \20671 , \20678 );
xor \U$20663 ( \21040 , \21039 , \20686 );
xor \U$20664 ( \21041 , \20645 , \20652 );
xor \U$20665 ( \21042 , \21041 , \20660 );
and \U$20666 ( \21043 , \21040 , \21042 );
xor \U$20667 ( \21044 , \20620 , \20627 );
xor \U$20668 ( \21045 , \21044 , \20635 );
xor \U$20669 ( \21046 , \20645 , \20652 );
xor \U$20670 ( \21047 , \21046 , \20660 );
and \U$20671 ( \21048 , \21045 , \21047 );
and \U$20672 ( \21049 , \21040 , \21045 );
or \U$20673 ( \21050 , \21043 , \21048 , \21049 );
xor \U$20674 ( \21051 , \20591 , \20598 );
xor \U$20675 ( \21052 , \21051 , \20606 );
xor \U$20676 ( \21053 , \20564 , \20572 );
xor \U$20677 ( \21054 , \21053 , \20580 );
and \U$20678 ( \21055 , \21052 , \21054 );
xor \U$20679 ( \21056 , \20537 , \20545 );
xor \U$20680 ( \21057 , \21056 , \20554 );
xor \U$20681 ( \21058 , \20564 , \20572 );
xor \U$20682 ( \21059 , \21058 , \20580 );
and \U$20683 ( \21060 , \21057 , \21059 );
and \U$20684 ( \21061 , \21052 , \21057 );
or \U$20685 ( \21062 , \21055 , \21060 , \21061 );
xor \U$20686 ( \21063 , \21050 , \21062 );
xor \U$20687 ( \21064 , \20454 , \20461 );
xor \U$20688 ( \21065 , \21064 , \20469 );
not \U$20689 ( \21066 , \20508 );
xor \U$20690 ( \21067 , \20516 , \20526 );
not \U$20691 ( \21068 , \21067 );
or \U$20692 ( \21069 , \21066 , \21068 );
or \U$20693 ( \21070 , \21067 , \20508 );
nand \U$20694 ( \21071 , \21069 , \21070 );
xor \U$20695 ( \21072 , \21065 , \21071 );
xor \U$20696 ( \21073 , \20480 , \20487 );
xor \U$20697 ( \21074 , \21073 , \20495 );
and \U$20698 ( \21075 , \21072 , \21074 );
and \U$20699 ( \21076 , \21065 , \21071 );
or \U$20700 ( \21077 , \21075 , \21076 );
and \U$20701 ( \21078 , \21063 , \21077 );
and \U$20702 ( \21079 , \21050 , \21062 );
or \U$20703 ( \21080 , \21078 , \21079 );
and \U$20704 ( \21081 , \21038 , \21080 );
and \U$20705 ( \21082 , \21023 , \21037 );
or \U$20706 ( \21083 , \21081 , \21082 );
xor \U$20707 ( \21084 , \20219 , \20237 );
xor \U$20708 ( \21085 , \21084 , \20263 );
not \U$20709 ( \21086 , \21085 );
not \U$20710 ( \21087 , \20498 );
xor \U$20711 ( \21088 , \20472 , \20528 );
not \U$20712 ( \21089 , \21088 );
or \U$20713 ( \21090 , \21087 , \21089 );
or \U$20714 ( \21091 , \21088 , \20498 );
nand \U$20715 ( \21092 , \21090 , \21091 );
xor \U$20716 ( \21093 , \20638 , \20663 );
xor \U$20717 ( \21094 , \21093 , \20689 );
and \U$20718 ( \21095 , \21092 , \21094 );
not \U$20719 ( \21096 , \21095 );
or \U$20720 ( \21097 , \21086 , \21096 );
or \U$20721 ( \21098 , \21095 , \21085 );
xor \U$20722 ( \21099 , \20557 , \20583 );
xor \U$20723 ( \21100 , \21099 , \20609 );
xor \U$20724 ( \21101 , \20712 , \20720 );
xor \U$20725 ( \21102 , \21101 , \20727 );
xor \U$20726 ( \21103 , \21100 , \21102 );
not \U$20727 ( \21104 , \20697 );
xor \U$20728 ( \21105 , \20705 , \20700 );
not \U$20729 ( \21106 , \21105 );
or \U$20730 ( \21107 , \21104 , \21106 );
or \U$20731 ( \21108 , \21105 , \20697 );
nand \U$20732 ( \21109 , \21107 , \21108 );
and \U$20733 ( \21110 , \21103 , \21109 );
and \U$20734 ( \21111 , \21100 , \21102 );
or \U$20735 ( \21112 , \21110 , \21111 );
nand \U$20736 ( \21113 , \21098 , \21112 );
nand \U$20737 ( \21114 , \21097 , \21113 );
xor \U$20738 ( \21115 , \21083 , \21114 );
xor \U$20739 ( \21116 , \20707 , \20730 );
xor \U$20740 ( \21117 , \21116 , \20748 );
xor \U$20741 ( \21118 , \20412 , \20422 );
xor \U$20742 ( \21119 , \21118 , \20433 );
xor \U$20743 ( \21120 , \21117 , \21119 );
xor \U$20744 ( \21121 , \20754 , \20756 );
xor \U$20745 ( \21122 , \21121 , \20767 );
and \U$20746 ( \21123 , \21120 , \21122 );
and \U$20747 ( \21124 , \21117 , \21119 );
nor \U$20748 ( \21125 , \21123 , \21124 );
and \U$20749 ( \21126 , \21115 , \21125 );
and \U$20750 ( \21127 , \21083 , \21114 );
or \U$20751 ( \21128 , \21126 , \21127 );
xor \U$20752 ( \21129 , \20787 , \21128 );
not \U$20753 ( \21130 , \20037 );
not \U$20754 ( \21131 , \20059 );
or \U$20755 ( \21132 , \21130 , \21131 );
or \U$20756 ( \21133 , \20059 , \20037 );
nand \U$20757 ( \21134 , \21132 , \21133 );
xor \U$20758 ( \21135 , \20035 , \21134 );
xor \U$20759 ( \21136 , \20111 , \20353 );
xor \U$20760 ( \21137 , \21136 , \20368 );
xor \U$20761 ( \21138 , \21135 , \21137 );
xor \U$20762 ( \21139 , \19628 , \19644 );
xor \U$20763 ( \21140 , \21139 , \19657 );
xor \U$20764 ( \21141 , \20017 , \20024 );
xor \U$20765 ( \21142 , \21140 , \21141 );
xor \U$20766 ( \21143 , \21138 , \21142 );
and \U$20767 ( \21144 , \21129 , \21143 );
and \U$20768 ( \21145 , \20787 , \21128 );
or \U$20769 ( \21146 , \21144 , \21145 );
not \U$20770 ( \21147 , \20030 );
xor \U$20771 ( \21148 , \20371 , \20061 );
not \U$20772 ( \21149 , \21148 );
or \U$20773 ( \21150 , \21147 , \21149 );
or \U$20774 ( \21151 , \21148 , \20030 );
nand \U$20775 ( \21152 , \21150 , \21151 );
xor \U$20776 ( \21153 , \21146 , \21152 );
xor \U$20777 ( \21154 , \21135 , \21137 );
and \U$20778 ( \21155 , \21154 , \21142 );
and \U$20779 ( \21156 , \21135 , \21137 );
or \U$20780 ( \21157 , \21155 , \21156 );
or \U$20781 ( \21158 , \20443 , \20409 );
not \U$20782 ( \21159 , \20409 );
not \U$20783 ( \21160 , \20443 );
or \U$20784 ( \21161 , \21159 , \21160 );
nand \U$20785 ( \21162 , \21161 , \20436 );
nand \U$20786 ( \21163 , \21158 , \21162 );
xor \U$20787 ( \21164 , \20695 , \20751 );
and \U$20788 ( \21165 , \21164 , \20770 );
and \U$20789 ( \21166 , \20695 , \20751 );
nor \U$20790 ( \21167 , \21165 , \21166 );
xor \U$20791 ( \21168 , \21163 , \21167 );
xor \U$20792 ( \21169 , \20074 , \20091 );
xor \U$20793 ( \21170 , \21169 , \20108 );
and \U$20794 ( \21171 , \20779 , \21170 );
xor \U$20795 ( \21172 , \20074 , \20091 );
xor \U$20796 ( \21173 , \21172 , \20108 );
and \U$20797 ( \21174 , \20783 , \21173 );
and \U$20798 ( \21175 , \20779 , \20783 );
or \U$20799 ( \21176 , \21171 , \21174 , \21175 );
and \U$20800 ( \21177 , \21168 , \21176 );
and \U$20801 ( \21178 , \21163 , \21167 );
or \U$20802 ( \21179 , \21177 , \21178 );
xor \U$20803 ( \21180 , \21157 , \21179 );
xor \U$20804 ( \21181 , \19608 , \19610 );
xor \U$20805 ( \21182 , \21181 , \19615 );
xor \U$20806 ( \21183 , \20389 , \20394 );
xor \U$20807 ( \21184 , \21182 , \21183 );
xor \U$20808 ( \21185 , \21180 , \21184 );
xor \U$20809 ( \21186 , \21153 , \21185 );
not \U$20810 ( \21187 , \21186 );
xnor \U$20811 ( \21188 , \20771 , \20447 );
not \U$20812 ( \21189 , \21188 );
not \U$20813 ( \21190 , \20785 );
and \U$20814 ( \21191 , \21189 , \21190 );
and \U$20815 ( \21192 , \21188 , \20785 );
nor \U$20816 ( \21193 , \21191 , \21192 );
xnor \U$20817 ( \21194 , \21112 , \21095 );
not \U$20818 ( \21195 , \21194 );
not \U$20819 ( \21196 , \21085 );
and \U$20820 ( \21197 , \21195 , \21196 );
and \U$20821 ( \21198 , \21194 , \21085 );
nor \U$20822 ( \21199 , \21197 , \21198 );
xor \U$20823 ( \21200 , \20530 , \20612 );
xor \U$20824 ( \21201 , \21200 , \20692 );
xor \U$20825 ( \21202 , \21199 , \21201 );
xor \U$20826 ( \21203 , \21117 , \21119 );
xor \U$20827 ( \21204 , \21203 , \21122 );
and \U$20828 ( \21205 , \21202 , \21204 );
and \U$20829 ( \21206 , \21199 , \21201 );
or \U$20830 ( \21207 , \21205 , \21206 );
or \U$20831 ( \21208 , \21193 , \21207 );
not \U$20832 ( \21209 , \21207 );
not \U$20833 ( \21210 , \21193 );
or \U$20834 ( \21211 , \21209 , \21210 );
xor \U$20835 ( \21212 , \20868 , \20940 );
xor \U$20836 ( \21213 , \21212 , \21020 );
xor \U$20837 ( \21214 , \20226 , \587 );
xor \U$20838 ( \21215 , \21214 , \20234 );
xor \U$20839 ( \21216 , \21025 , \21032 );
xor \U$20840 ( \21217 , \21215 , \21216 );
xor \U$20841 ( \21218 , \21213 , \21217 );
xor \U$20842 ( \21219 , \21050 , \21062 );
xor \U$20843 ( \21220 , \21219 , \21077 );
and \U$20844 ( \21221 , \21218 , \21220 );
and \U$20845 ( \21222 , \21213 , \21217 );
or \U$20846 ( \21223 , \21221 , \21222 );
xor \U$20847 ( \21224 , \20845 , \20853 );
xor \U$20848 ( \21225 , \21224 , \20862 );
xor \U$20849 ( \21226 , \20999 , \21006 );
xor \U$20850 ( \21227 , \21226 , \21014 );
and \U$20851 ( \21228 , \21225 , \21227 );
xor \U$20852 ( \21229 , \20973 , \20980 );
xor \U$20853 ( \21230 , \21229 , \20988 );
xor \U$20854 ( \21231 , \20999 , \21006 );
xor \U$20855 ( \21232 , \21231 , \21014 );
and \U$20856 ( \21233 , \21230 , \21232 );
and \U$20857 ( \21234 , \21225 , \21230 );
or \U$20858 ( \21235 , \21228 , \21233 , \21234 );
nand \U$20859 ( \21236 , RIae775b8_79, \881 );
not \U$20860 ( \21237 , \21236 );
not \U$20861 ( \21238 , \787 );
or \U$20862 ( \21239 , \21237 , \21238 );
or \U$20863 ( \21240 , \787 , \21236 );
nand \U$20864 ( \21241 , \21239 , \21240 );
xor \U$20865 ( \21242 , \20794 , \20801 );
xor \U$20866 ( \21243 , \21242 , \20809 );
and \U$20867 ( \21244 , \21241 , \21243 );
xor \U$20868 ( \21245 , \20819 , \20826 );
xor \U$20869 ( \21246 , \21245 , \20834 );
xor \U$20870 ( \21247 , \20794 , \20801 );
xor \U$20871 ( \21248 , \21247 , \20809 );
and \U$20872 ( \21249 , \21246 , \21248 );
and \U$20873 ( \21250 , \21241 , \21246 );
or \U$20874 ( \21251 , \21244 , \21249 , \21250 );
xor \U$20875 ( \21252 , \21235 , \21251 );
xor \U$20876 ( \21253 , \20919 , \20926 );
xor \U$20877 ( \21254 , \21253 , \20934 );
xor \U$20878 ( \21255 , \20948 , \20955 );
xor \U$20879 ( \21256 , \21255 , \20963 );
xor \U$20880 ( \21257 , \21254 , \21256 );
xor \U$20881 ( \21258 , \20875 , \20882 );
xor \U$20882 ( \21259 , \21258 , \20890 );
and \U$20883 ( \21260 , \21257 , \21259 );
and \U$20884 ( \21261 , \21254 , \21256 );
or \U$20885 ( \21262 , \21260 , \21261 );
and \U$20886 ( \21263 , \21252 , \21262 );
and \U$20887 ( \21264 , \21235 , \21251 );
or \U$20888 ( \21265 , \21263 , \21264 );
and \U$20889 ( \21266 , \1939 , RIae77798_83);
and \U$20890 ( \21267 , RIae77888_85, \1937 );
nor \U$20891 ( \21268 , \21266 , \21267 );
and \U$20892 ( \21269 , \21268 , \1735 );
not \U$20893 ( \21270 , \21268 );
and \U$20894 ( \21271 , \21270 , \1734 );
nor \U$20895 ( \21272 , \21269 , \21271 );
and \U$20896 ( \21273 , \1593 , RIae77a68_89);
and \U$20897 ( \21274 , RIae77978_87, \1591 );
nor \U$20898 ( \21275 , \21273 , \21274 );
and \U$20899 ( \21276 , \21275 , \1498 );
not \U$20900 ( \21277 , \21275 );
and \U$20901 ( \21278 , \21277 , \1488 );
nor \U$20902 ( \21279 , \21276 , \21278 );
xor \U$20903 ( \21280 , \21272 , \21279 );
and \U$20904 ( \21281 , \2224 , RIae76f28_65);
and \U$20905 ( \21282 , RIae76e38_63, \2222 );
nor \U$20906 ( \21283 , \21281 , \21282 );
and \U$20907 ( \21284 , \21283 , \2061 );
not \U$20908 ( \21285 , \21283 );
and \U$20909 ( \21286 , \21285 , \2060 );
nor \U$20910 ( \21287 , \21284 , \21286 );
and \U$20911 ( \21288 , \21280 , \21287 );
and \U$20912 ( \21289 , \21272 , \21279 );
or \U$20913 ( \21290 , \21288 , \21289 );
and \U$20914 ( \21291 , \1376 , RIae77720_82);
and \U$20915 ( \21292 , RIae773d8_75, \1374 );
nor \U$20916 ( \21293 , \21291 , \21292 );
and \U$20917 ( \21294 , \21293 , \1380 );
not \U$20918 ( \21295 , \21293 );
and \U$20919 ( \21296 , \21295 , \1261 );
nor \U$20920 ( \21297 , \21294 , \21296 );
and \U$20921 ( \21298 , \1138 , RIae775b8_79);
and \U$20922 ( \21299 , RIae774c8_77, \1136 );
nor \U$20923 ( \21300 , \21298 , \21299 );
and \U$20924 ( \21301 , \21300 , \1012 );
not \U$20925 ( \21302 , \21300 );
and \U$20926 ( \21303 , \21302 , \1142 );
nor \U$20927 ( \21304 , \21301 , \21303 );
and \U$20928 ( \21305 , \21297 , \21304 );
xor \U$20929 ( \21306 , \21290 , \21305 );
not \U$20930 ( \21307 , \3218 );
and \U$20931 ( \21308 , \3214 , RIae771f8_71);
and \U$20932 ( \21309 , RIae772e8_73, \3212 );
nor \U$20933 ( \21310 , \21308 , \21309 );
not \U$20934 ( \21311 , \21310 );
or \U$20935 ( \21312 , \21307 , \21311 );
or \U$20936 ( \21313 , \21310 , \2774 );
nand \U$20937 ( \21314 , \21312 , \21313 );
and \U$20938 ( \21315 , \2607 , RIae76d48_61);
and \U$20939 ( \21316 , RIae76c58_59, \2605 );
nor \U$20940 ( \21317 , \21315 , \21316 );
and \U$20941 ( \21318 , \21317 , \2611 );
not \U$20942 ( \21319 , \21317 );
and \U$20943 ( \21320 , \21319 , \2397 );
nor \U$20944 ( \21321 , \21318 , \21320 );
xor \U$20945 ( \21322 , \21314 , \21321 );
not \U$20946 ( \21323 , \2789 );
and \U$20947 ( \21324 , \2783 , RIae77180_70);
and \U$20948 ( \21325 , RIae77018_67, \2781 );
nor \U$20949 ( \21326 , \21324 , \21325 );
not \U$20950 ( \21327 , \21326 );
or \U$20951 ( \21328 , \21323 , \21327 );
or \U$20952 ( \21329 , \21326 , \2789 );
nand \U$20953 ( \21330 , \21328 , \21329 );
and \U$20954 ( \21331 , \21322 , \21330 );
and \U$20955 ( \21332 , \21314 , \21321 );
or \U$20956 ( \21333 , \21331 , \21332 );
and \U$20957 ( \21334 , \21306 , \21333 );
and \U$20958 ( \21335 , \21290 , \21305 );
or \U$20959 ( \21336 , \21334 , \21335 );
and \U$20960 ( \21337 , \10548 , RIae75c68_25);
and \U$20961 ( \21338 , RIae75d58_27, \10546 );
nor \U$20962 ( \21339 , \21337 , \21338 );
and \U$20963 ( \21340 , \21339 , \10421 );
not \U$20964 ( \21341 , \21339 );
and \U$20965 ( \21342 , \21341 , \10118 );
nor \U$20966 ( \21343 , \21340 , \21342 );
and \U$20967 ( \21344 , \8966 , RIae75998_19);
and \U$20968 ( \21345 , RIae758a8_17, \8964 );
nor \U$20969 ( \21346 , \21344 , \21345 );
and \U$20970 ( \21347 , \21346 , \8799 );
not \U$20971 ( \21348 , \21346 );
and \U$20972 ( \21349 , \21348 , \8789 );
nor \U$20973 ( \21350 , \21347 , \21349 );
xor \U$20974 ( \21351 , \21343 , \21350 );
and \U$20975 ( \21352 , \9760 , RIae75f38_31);
and \U$20976 ( \21353 , RIae75e48_29, \9758 );
nor \U$20977 ( \21354 , \21352 , \21353 );
and \U$20978 ( \21355 , \21354 , \9273 );
not \U$20979 ( \21356 , \21354 );
and \U$20980 ( \21357 , \21356 , \9764 );
nor \U$20981 ( \21358 , \21355 , \21357 );
and \U$20982 ( \21359 , \21351 , \21358 );
and \U$20983 ( \21360 , \21343 , \21350 );
or \U$20984 ( \21361 , \21359 , \21360 );
and \U$20985 ( \21362 , \15726 , RIae766b8_47);
and \U$20986 ( \21363 , RIae7aab0_192, RIae765c8_45);
nor \U$20987 ( \21364 , \21362 , \21363 );
and \U$20988 ( \21365 , \21364 , RIae7aa38_191);
not \U$20989 ( \21366 , \21364 );
and \U$20990 ( \21367 , \21366 , \14959 );
nor \U$20991 ( \21368 , \21365 , \21367 );
and \U$20992 ( \21369 , \14964 , RIae763e8_41);
and \U$20993 ( \21370 , RIae764d8_43, \14962 );
nor \U$20994 ( \21371 , \21369 , \21370 );
and \U$20995 ( \21372 , \21371 , \14462 );
not \U$20996 ( \21373 , \21371 );
and \U$20997 ( \21374 , \21373 , \14463 );
nor \U$20998 ( \21375 , \21372 , \21374 );
xor \U$20999 ( \21376 , \21368 , \21375 );
and \U$21000 ( \21377 , \14059 , RIae75308_5);
and \U$21001 ( \21378 , RIae753f8_7, \14057 );
nor \U$21002 ( \21379 , \21377 , \21378 );
and \U$21003 ( \21380 , \21379 , \14063 );
not \U$21004 ( \21381 , \21379 );
and \U$21005 ( \21382 , \21381 , \13502 );
nor \U$21006 ( \21383 , \21380 , \21382 );
and \U$21007 ( \21384 , \21376 , \21383 );
and \U$21008 ( \21385 , \21368 , \21375 );
nor \U$21009 ( \21386 , \21384 , \21385 );
xor \U$21010 ( \21387 , \21361 , \21386 );
and \U$21011 ( \21388 , \11470 , RIae755d8_11);
and \U$21012 ( \21389 , RIae754e8_9, \11468 );
nor \U$21013 ( \21390 , \21388 , \21389 );
and \U$21014 ( \21391 , \21390 , \11474 );
not \U$21015 ( \21392 , \21390 );
and \U$21016 ( \21393 , \21392 , \10936 );
nor \U$21017 ( \21394 , \21391 , \21393 );
and \U$21018 ( \21395 , \12180 , RIae757b8_15);
and \U$21019 ( \21396 , RIae756c8_13, \12178 );
nor \U$21020 ( \21397 , \21395 , \21396 );
and \U$21021 ( \21398 , \21397 , \11827 );
not \U$21022 ( \21399 , \21397 );
and \U$21023 ( \21400 , \21399 , \12184 );
nor \U$21024 ( \21401 , \21398 , \21400 );
or \U$21025 ( \21402 , \21394 , \21401 );
not \U$21026 ( \21403 , \21401 );
not \U$21027 ( \21404 , \21394 );
or \U$21028 ( \21405 , \21403 , \21404 );
and \U$21029 ( \21406 , \13059 , RIae75218_3);
and \U$21030 ( \21407 , RIae75128_1, \13057 );
nor \U$21031 ( \21408 , \21406 , \21407 );
and \U$21032 ( \21409 , \21408 , \13063 );
not \U$21033 ( \21410 , \21408 );
and \U$21034 ( \21411 , \21410 , \12718 );
nor \U$21035 ( \21412 , \21409 , \21411 );
nand \U$21036 ( \21413 , \21405 , \21412 );
nand \U$21037 ( \21414 , \21402 , \21413 );
and \U$21038 ( \21415 , \21387 , \21414 );
and \U$21039 ( \21416 , \21361 , \21386 );
or \U$21040 ( \21417 , \21415 , \21416 );
xor \U$21041 ( \21418 , \21336 , \21417 );
and \U$21042 ( \21419 , \6172 , RIae77d38_95);
and \U$21043 ( \21420 , RIae77e28_97, \6170 );
nor \U$21044 ( \21421 , \21419 , \21420 );
and \U$21045 ( \21422 , \21421 , \6176 );
not \U$21046 ( \21423 , \21421 );
and \U$21047 ( \21424 , \21423 , \6175 );
nor \U$21048 ( \21425 , \21422 , \21424 );
and \U$21049 ( \21426 , \5399 , RIae783c8_109);
and \U$21050 ( \21427 , RIae78530_112, \5397 );
nor \U$21051 ( \21428 , \21426 , \21427 );
and \U$21052 ( \21429 , \21428 , \5016 );
not \U$21053 ( \21430 , \21428 );
and \U$21054 ( \21431 , \21430 , \5403 );
nor \U$21055 ( \21432 , \21429 , \21431 );
xor \U$21056 ( \21433 , \21425 , \21432 );
and \U$21057 ( \21434 , \5896 , RIae77c48_93);
and \U$21058 ( \21435 , RIae77b58_91, \5894 );
nor \U$21059 ( \21436 , \21434 , \21435 );
and \U$21060 ( \21437 , \21436 , \5590 );
not \U$21061 ( \21438 , \21436 );
and \U$21062 ( \21439 , \21438 , \5589 );
nor \U$21063 ( \21440 , \21437 , \21439 );
and \U$21064 ( \21441 , \21433 , \21440 );
and \U$21065 ( \21442 , \21425 , \21432 );
or \U$21066 ( \21443 , \21441 , \21442 );
and \U$21067 ( \21444 , \4688 , RIae781e8_105);
and \U$21068 ( \21445 , RIae785a8_113, \4686 );
nor \U$21069 ( \21446 , \21444 , \21445 );
and \U$21070 ( \21447 , \21446 , \4481 );
not \U$21071 ( \21448 , \21446 );
and \U$21072 ( \21449 , \21448 , \4482 );
nor \U$21073 ( \21450 , \21447 , \21449 );
and \U$21074 ( \21451 , \3730 , RIae782d8_107);
and \U$21075 ( \21452 , RIae780f8_103, \3728 );
nor \U$21076 ( \21453 , \21451 , \21452 );
and \U$21077 ( \21454 , \21453 , \3732 );
not \U$21078 ( \21455 , \21453 );
and \U$21079 ( \21456 , \21455 , \3422 );
nor \U$21080 ( \21457 , \21454 , \21456 );
xor \U$21081 ( \21458 , \21450 , \21457 );
and \U$21082 ( \21459 , \4247 , RIae77f18_99);
and \U$21083 ( \21460 , RIae78008_101, \4245 );
nor \U$21084 ( \21461 , \21459 , \21460 );
and \U$21085 ( \21462 , \21461 , \3989 );
not \U$21086 ( \21463 , \21461 );
and \U$21087 ( \21464 , \21463 , \4251 );
nor \U$21088 ( \21465 , \21462 , \21464 );
and \U$21089 ( \21466 , \21458 , \21465 );
and \U$21090 ( \21467 , \21450 , \21457 );
or \U$21091 ( \21468 , \21466 , \21467 );
xor \U$21092 ( \21469 , \21443 , \21468 );
and \U$21093 ( \21470 , \8371 , RIae75b78_23);
and \U$21094 ( \21471 , RIae75a88_21, \8369 );
nor \U$21095 ( \21472 , \21470 , \21471 );
and \U$21096 ( \21473 , \21472 , \8020 );
not \U$21097 ( \21474 , \21472 );
and \U$21098 ( \21475 , \21474 , \8019 );
nor \U$21099 ( \21476 , \21473 , \21475 );
and \U$21100 ( \21477 , \6941 , RIae78968_121);
and \U$21101 ( \21478 , RIae78878_119, \6939 );
nor \U$21102 ( \21479 , \21477 , \21478 );
and \U$21103 ( \21480 , \21479 , \6314 );
not \U$21104 ( \21481 , \21479 );
and \U$21105 ( \21482 , \21481 , \6945 );
nor \U$21106 ( \21483 , \21480 , \21482 );
xor \U$21107 ( \21484 , \21476 , \21483 );
and \U$21108 ( \21485 , \7633 , RIae78788_117);
and \U$21109 ( \21486 , RIae78698_115, \7631 );
nor \U$21110 ( \21487 , \21485 , \21486 );
and \U$21111 ( \21488 , \21487 , \7206 );
not \U$21112 ( \21489 , \21487 );
and \U$21113 ( \21490 , \21489 , \7205 );
nor \U$21114 ( \21491 , \21488 , \21490 );
and \U$21115 ( \21492 , \21484 , \21491 );
and \U$21116 ( \21493 , \21476 , \21483 );
or \U$21117 ( \21494 , \21492 , \21493 );
and \U$21118 ( \21495 , \21469 , \21494 );
and \U$21119 ( \21496 , \21443 , \21468 );
or \U$21120 ( \21497 , \21495 , \21496 );
and \U$21121 ( \21498 , \21418 , \21497 );
and \U$21122 ( \21499 , \21336 , \21417 );
or \U$21123 ( \21500 , \21498 , \21499 );
xor \U$21124 ( \21501 , \21265 , \21500 );
xor \U$21125 ( \21502 , \20645 , \20652 );
xor \U$21126 ( \21503 , \21502 , \20660 );
xor \U$21127 ( \21504 , \21040 , \21045 );
xor \U$21128 ( \21505 , \21503 , \21504 );
xor \U$21129 ( \21506 , \21065 , \21071 );
xor \U$21130 ( \21507 , \21506 , \21074 );
and \U$21131 ( \21508 , \21505 , \21507 );
xor \U$21132 ( \21509 , \20564 , \20572 );
xor \U$21133 ( \21510 , \21509 , \20580 );
xor \U$21134 ( \21511 , \21052 , \21057 );
xor \U$21135 ( \21512 , \21510 , \21511 );
xor \U$21136 ( \21513 , \21065 , \21071 );
xor \U$21137 ( \21514 , \21513 , \21074 );
and \U$21138 ( \21515 , \21512 , \21514 );
and \U$21139 ( \21516 , \21505 , \21512 );
or \U$21140 ( \21517 , \21508 , \21515 , \21516 );
and \U$21141 ( \21518 , \21501 , \21517 );
and \U$21142 ( \21519 , \21265 , \21500 );
or \U$21143 ( \21520 , \21518 , \21519 );
xor \U$21144 ( \21521 , \21223 , \21520 );
xor \U$21145 ( \21522 , \20812 , \20837 );
xor \U$21146 ( \21523 , \21522 , \20865 );
xor \U$21147 ( \21524 , \20893 , \20911 );
xor \U$21148 ( \21525 , \21524 , \20937 );
xor \U$21149 ( \21526 , \21523 , \21525 );
xor \U$21150 ( \21527 , \20966 , \20991 );
xor \U$21151 ( \21528 , \21527 , \21017 );
and \U$21152 ( \21529 , \21526 , \21528 );
and \U$21153 ( \21530 , \21523 , \21525 );
or \U$21154 ( \21531 , \21529 , \21530 );
xor \U$21155 ( \21532 , \21092 , \21094 );
xor \U$21156 ( \21533 , \21531 , \21532 );
xor \U$21157 ( \21534 , \21100 , \21102 );
xor \U$21158 ( \21535 , \21534 , \21109 );
and \U$21159 ( \21536 , \21533 , \21535 );
and \U$21160 ( \21537 , \21531 , \21532 );
or \U$21161 ( \21538 , \21536 , \21537 );
and \U$21162 ( \21539 , \21521 , \21538 );
and \U$21163 ( \21540 , \21223 , \21520 );
or \U$21164 ( \21541 , \21539 , \21540 );
nand \U$21165 ( \21542 , \21211 , \21541 );
nand \U$21166 ( \21543 , \21208 , \21542 );
xor \U$21167 ( \21544 , \21163 , \21167 );
xor \U$21168 ( \21545 , \21544 , \21176 );
and \U$21169 ( \21546 , \21543 , \21545 );
xor \U$21170 ( \21547 , \20787 , \21128 );
xor \U$21171 ( \21548 , \21547 , \21143 );
xor \U$21172 ( \21549 , \21163 , \21167 );
xor \U$21173 ( \21550 , \21549 , \21176 );
and \U$21174 ( \21551 , \21548 , \21550 );
and \U$21175 ( \21552 , \21543 , \21548 );
or \U$21176 ( \21553 , \21546 , \21551 , \21552 );
not \U$21177 ( \21554 , \21553 );
not \U$21178 ( \21555 , \21554 );
or \U$21179 ( \21556 , \21187 , \21555 );
or \U$21180 ( \21557 , \21186 , \21554 );
nand \U$21181 ( \21558 , \21556 , \21557 );
xor \U$21182 ( \21559 , \21163 , \21167 );
xor \U$21183 ( \21560 , \21559 , \21176 );
xor \U$21184 ( \21561 , \21543 , \21548 );
xor \U$21185 ( \21562 , \21560 , \21561 );
not \U$21186 ( \21563 , \21562 );
xor \U$21187 ( \21564 , \21083 , \21114 );
xor \U$21188 ( \21565 , \21564 , \21125 );
not \U$21189 ( \21566 , \21565 );
xor \U$21190 ( \21567 , \21199 , \21201 );
xor \U$21191 ( \21568 , \21567 , \21204 );
not \U$21192 ( \21569 , \21568 );
xor \U$21193 ( \21570 , \21223 , \21520 );
xor \U$21194 ( \21571 , \21570 , \21538 );
nand \U$21195 ( \21572 , \21569 , \21571 );
nand \U$21196 ( \21573 , \21566 , \21572 );
xor \U$21197 ( \21574 , \21368 , \21375 );
xor \U$21198 ( \21575 , \21574 , \21383 );
not \U$21199 ( \21576 , \21401 );
not \U$21200 ( \21577 , \21412 );
or \U$21201 ( \21578 , \21576 , \21577 );
or \U$21202 ( \21579 , \21401 , \21412 );
nand \U$21203 ( \21580 , \21578 , \21579 );
not \U$21204 ( \21581 , \21580 );
not \U$21205 ( \21582 , \21394 );
and \U$21206 ( \21583 , \21581 , \21582 );
and \U$21207 ( \21584 , \21580 , \21394 );
nor \U$21208 ( \21585 , \21583 , \21584 );
or \U$21209 ( \21586 , \21575 , \21585 );
not \U$21210 ( \21587 , \21585 );
not \U$21211 ( \21588 , \21575 );
or \U$21212 ( \21589 , \21587 , \21588 );
xor \U$21213 ( \21590 , \21343 , \21350 );
xor \U$21214 ( \21591 , \21590 , \21358 );
nand \U$21215 ( \21592 , \21589 , \21591 );
nand \U$21216 ( \21593 , \21586 , \21592 );
xor \U$21217 ( \21594 , \21297 , \21304 );
not \U$21218 ( \21595 , \21594 );
xor \U$21219 ( \21596 , \21314 , \21321 );
xor \U$21220 ( \21597 , \21596 , \21330 );
not \U$21221 ( \21598 , \21597 );
or \U$21222 ( \21599 , \21595 , \21598 );
or \U$21223 ( \21600 , \21597 , \21594 );
xor \U$21224 ( \21601 , \21272 , \21279 );
xor \U$21225 ( \21602 , \21601 , \21287 );
nand \U$21226 ( \21603 , \21600 , \21602 );
nand \U$21227 ( \21604 , \21599 , \21603 );
xor \U$21228 ( \21605 , \21593 , \21604 );
xor \U$21229 ( \21606 , \21450 , \21457 );
xor \U$21230 ( \21607 , \21606 , \21465 );
xor \U$21231 ( \21608 , \21425 , \21432 );
xor \U$21232 ( \21609 , \21608 , \21440 );
and \U$21233 ( \21610 , \21607 , \21609 );
xor \U$21234 ( \21611 , \21476 , \21483 );
xor \U$21235 ( \21612 , \21611 , \21491 );
xor \U$21236 ( \21613 , \21425 , \21432 );
xor \U$21237 ( \21614 , \21613 , \21440 );
and \U$21238 ( \21615 , \21612 , \21614 );
and \U$21239 ( \21616 , \21607 , \21612 );
or \U$21240 ( \21617 , \21610 , \21615 , \21616 );
and \U$21241 ( \21618 , \21605 , \21617 );
and \U$21242 ( \21619 , \21593 , \21604 );
or \U$21243 ( \21620 , \21618 , \21619 );
and \U$21244 ( \21621 , \2224 , RIae77888_85);
and \U$21245 ( \21622 , RIae76f28_65, \2222 );
nor \U$21246 ( \21623 , \21621 , \21622 );
and \U$21247 ( \21624 , \21623 , \2060 );
not \U$21248 ( \21625 , \21623 );
and \U$21249 ( \21626 , \21625 , \2061 );
nor \U$21250 ( \21627 , \21624 , \21626 );
and \U$21251 ( \21628 , \2607 , RIae76e38_63);
and \U$21252 ( \21629 , RIae76d48_61, \2605 );
nor \U$21253 ( \21630 , \21628 , \21629 );
and \U$21254 ( \21631 , \21630 , \2397 );
not \U$21255 ( \21632 , \21630 );
and \U$21256 ( \21633 , \21632 , \2611 );
nor \U$21257 ( \21634 , \21631 , \21633 );
xor \U$21258 ( \21635 , \21627 , \21634 );
and \U$21259 ( \21636 , \1939 , RIae77978_87);
and \U$21260 ( \21637 , RIae77798_83, \1937 );
nor \U$21261 ( \21638 , \21636 , \21637 );
and \U$21262 ( \21639 , \21638 , \1734 );
not \U$21263 ( \21640 , \21638 );
and \U$21264 ( \21641 , \21640 , \1735 );
nor \U$21265 ( \21642 , \21639 , \21641 );
and \U$21266 ( \21643 , \21635 , \21642 );
and \U$21267 ( \21644 , \21627 , \21634 );
nor \U$21268 ( \21645 , \21643 , \21644 );
and \U$21269 ( \21646 , \1376 , RIae774c8_77);
and \U$21270 ( \21647 , RIae77720_82, \1374 );
nor \U$21271 ( \21648 , \21646 , \21647 );
and \U$21272 ( \21649 , \21648 , \1380 );
not \U$21273 ( \21650 , \21648 );
and \U$21274 ( \21651 , \21650 , \1261 );
nor \U$21275 ( \21652 , \21649 , \21651 );
nand \U$21276 ( \21653 , RIae775b8_79, \1136 );
and \U$21277 ( \21654 , \21653 , \1012 );
not \U$21278 ( \21655 , \21653 );
and \U$21279 ( \21656 , \21655 , \1142 );
nor \U$21280 ( \21657 , \21654 , \21656 );
xor \U$21281 ( \21658 , \21652 , \21657 );
and \U$21282 ( \21659 , \1593 , RIae773d8_75);
and \U$21283 ( \21660 , RIae77a68_89, \1591 );
nor \U$21284 ( \21661 , \21659 , \21660 );
and \U$21285 ( \21662 , \21661 , \1498 );
not \U$21286 ( \21663 , \21661 );
and \U$21287 ( \21664 , \21663 , \1488 );
nor \U$21288 ( \21665 , \21662 , \21664 );
and \U$21289 ( \21666 , \21658 , \21665 );
and \U$21290 ( \21667 , \21652 , \21657 );
or \U$21291 ( \21668 , \21666 , \21667 );
xor \U$21292 ( \21669 , \21645 , \21668 );
and \U$21293 ( \21670 , \3214 , RIae77018_67);
and \U$21294 ( \21671 , RIae771f8_71, \3212 );
nor \U$21295 ( \21672 , \21670 , \21671 );
not \U$21296 ( \21673 , \21672 );
not \U$21297 ( \21674 , \2774 );
and \U$21298 ( \21675 , \21673 , \21674 );
and \U$21299 ( \21676 , \21672 , \2774 );
nor \U$21300 ( \21677 , \21675 , \21676 );
and \U$21301 ( \21678 , \3730 , RIae772e8_73);
and \U$21302 ( \21679 , RIae782d8_107, \3728 );
nor \U$21303 ( \21680 , \21678 , \21679 );
and \U$21304 ( \21681 , \21680 , \3422 );
not \U$21305 ( \21682 , \21680 );
and \U$21306 ( \21683 , \21682 , \3732 );
nor \U$21307 ( \21684 , \21681 , \21683 );
xor \U$21308 ( \21685 , \21677 , \21684 );
and \U$21309 ( \21686 , \2783 , RIae76c58_59);
and \U$21310 ( \21687 , RIae77180_70, \2781 );
nor \U$21311 ( \21688 , \21686 , \21687 );
not \U$21312 ( \21689 , \21688 );
not \U$21313 ( \21690 , \2789 );
and \U$21314 ( \21691 , \21689 , \21690 );
and \U$21315 ( \21692 , \21688 , \2789 );
nor \U$21316 ( \21693 , \21691 , \21692 );
and \U$21317 ( \21694 , \21685 , \21693 );
and \U$21318 ( \21695 , \21677 , \21684 );
nor \U$21319 ( \21696 , \21694 , \21695 );
and \U$21320 ( \21697 , \21669 , \21696 );
and \U$21321 ( \21698 , \21645 , \21668 );
or \U$21322 ( \21699 , \21697 , \21698 );
and \U$21323 ( \21700 , \9760 , RIae758a8_17);
and \U$21324 ( \21701 , RIae75f38_31, \9758 );
nor \U$21325 ( \21702 , \21700 , \21701 );
and \U$21326 ( \21703 , \21702 , \9273 );
not \U$21327 ( \21704 , \21702 );
and \U$21328 ( \21705 , \21704 , \9764 );
nor \U$21329 ( \21706 , \21703 , \21705 );
and \U$21330 ( \21707 , \10548 , RIae75e48_29);
and \U$21331 ( \21708 , RIae75c68_25, \10546 );
nor \U$21332 ( \21709 , \21707 , \21708 );
and \U$21333 ( \21710 , \21709 , \10421 );
not \U$21334 ( \21711 , \21709 );
and \U$21335 ( \21712 , \21711 , \10118 );
nor \U$21336 ( \21713 , \21710 , \21712 );
xor \U$21337 ( \21714 , \21706 , \21713 );
and \U$21338 ( \21715 , \11470 , RIae75d58_27);
and \U$21339 ( \21716 , RIae755d8_11, \11468 );
nor \U$21340 ( \21717 , \21715 , \21716 );
and \U$21341 ( \21718 , \21717 , \10936 );
not \U$21342 ( \21719 , \21717 );
and \U$21343 ( \21720 , \21719 , \11474 );
nor \U$21344 ( \21721 , \21718 , \21720 );
and \U$21345 ( \21722 , \21714 , \21721 );
and \U$21346 ( \21723 , \21706 , \21713 );
or \U$21347 ( \21724 , \21722 , \21723 );
and \U$21348 ( \21725 , \15726 , RIae764d8_43);
and \U$21349 ( \21726 , RIae7aab0_192, RIae766b8_47);
nor \U$21350 ( \21727 , \21725 , \21726 );
and \U$21351 ( \21728 , \21727 , \14959 );
not \U$21352 ( \21729 , \21727 );
and \U$21353 ( \21730 , \21729 , RIae7aa38_191);
nor \U$21354 ( \21731 , \21728 , \21730 );
xor \U$21355 ( \21732 , \21731 , \1142 );
and \U$21356 ( \21733 , \14964 , RIae753f8_7);
and \U$21357 ( \21734 , RIae763e8_41, \14962 );
nor \U$21358 ( \21735 , \21733 , \21734 );
and \U$21359 ( \21736 , \21735 , \14463 );
not \U$21360 ( \21737 , \21735 );
and \U$21361 ( \21738 , \21737 , \14462 );
nor \U$21362 ( \21739 , \21736 , \21738 );
and \U$21363 ( \21740 , \21732 , \21739 );
and \U$21364 ( \21741 , \21731 , \1142 );
or \U$21365 ( \21742 , \21740 , \21741 );
xor \U$21366 ( \21743 , \21724 , \21742 );
and \U$21367 ( \21744 , \13059 , RIae756c8_13);
and \U$21368 ( \21745 , RIae75218_3, \13057 );
nor \U$21369 ( \21746 , \21744 , \21745 );
and \U$21370 ( \21747 , \21746 , \12718 );
not \U$21371 ( \21748 , \21746 );
and \U$21372 ( \21749 , \21748 , \13063 );
nor \U$21373 ( \21750 , \21747 , \21749 );
and \U$21374 ( \21751 , \14059 , RIae75128_1);
and \U$21375 ( \21752 , RIae75308_5, \14057 );
nor \U$21376 ( \21753 , \21751 , \21752 );
and \U$21377 ( \21754 , \21753 , \14063 );
not \U$21378 ( \21755 , \21753 );
and \U$21379 ( \21756 , \21755 , \13502 );
nor \U$21380 ( \21757 , \21754 , \21756 );
xor \U$21381 ( \21758 , \21750 , \21757 );
and \U$21382 ( \21759 , \12180 , RIae754e8_9);
and \U$21383 ( \21760 , RIae757b8_15, \12178 );
nor \U$21384 ( \21761 , \21759 , \21760 );
and \U$21385 ( \21762 , \21761 , \11827 );
not \U$21386 ( \21763 , \21761 );
and \U$21387 ( \21764 , \21763 , \12184 );
nor \U$21388 ( \21765 , \21762 , \21764 );
and \U$21389 ( \21766 , \21758 , \21765 );
and \U$21390 ( \21767 , \21750 , \21757 );
nor \U$21391 ( \21768 , \21766 , \21767 );
and \U$21392 ( \21769 , \21743 , \21768 );
and \U$21393 ( \21770 , \21724 , \21742 );
or \U$21394 ( \21771 , \21769 , \21770 );
xor \U$21395 ( \21772 , \21699 , \21771 );
and \U$21396 ( \21773 , \7633 , RIae78878_119);
and \U$21397 ( \21774 , RIae78788_117, \7631 );
nor \U$21398 ( \21775 , \21773 , \21774 );
and \U$21399 ( \21776 , \21775 , \7206 );
not \U$21400 ( \21777 , \21775 );
and \U$21401 ( \21778 , \21777 , \7205 );
nor \U$21402 ( \21779 , \21776 , \21778 );
and \U$21403 ( \21780 , \8371 , RIae78698_115);
and \U$21404 ( \21781 , RIae75b78_23, \8369 );
nor \U$21405 ( \21782 , \21780 , \21781 );
and \U$21406 ( \21783 , \21782 , \8020 );
not \U$21407 ( \21784 , \21782 );
and \U$21408 ( \21785 , \21784 , \8019 );
nor \U$21409 ( \21786 , \21783 , \21785 );
xor \U$21410 ( \21787 , \21779 , \21786 );
and \U$21411 ( \21788 , \8966 , RIae75a88_21);
and \U$21412 ( \21789 , RIae75998_19, \8964 );
nor \U$21413 ( \21790 , \21788 , \21789 );
and \U$21414 ( \21791 , \21790 , \8799 );
not \U$21415 ( \21792 , \21790 );
and \U$21416 ( \21793 , \21792 , \8789 );
nor \U$21417 ( \21794 , \21791 , \21793 );
and \U$21418 ( \21795 , \21787 , \21794 );
and \U$21419 ( \21796 , \21779 , \21786 );
or \U$21420 ( \21797 , \21795 , \21796 );
and \U$21421 ( \21798 , \4247 , RIae780f8_103);
and \U$21422 ( \21799 , RIae77f18_99, \4245 );
nor \U$21423 ( \21800 , \21798 , \21799 );
and \U$21424 ( \21801 , \21800 , \4251 );
not \U$21425 ( \21802 , \21800 );
and \U$21426 ( \21803 , \21802 , \3989 );
nor \U$21427 ( \21804 , \21801 , \21803 );
and \U$21428 ( \21805 , \5399 , RIae785a8_113);
and \U$21429 ( \21806 , RIae783c8_109, \5397 );
nor \U$21430 ( \21807 , \21805 , \21806 );
and \U$21431 ( \21808 , \21807 , \5403 );
not \U$21432 ( \21809 , \21807 );
and \U$21433 ( \21810 , \21809 , \5016 );
nor \U$21434 ( \21811 , \21808 , \21810 );
or \U$21435 ( \21812 , \21804 , \21811 );
not \U$21436 ( \21813 , \21811 );
not \U$21437 ( \21814 , \21804 );
or \U$21438 ( \21815 , \21813 , \21814 );
and \U$21439 ( \21816 , \4688 , RIae78008_101);
and \U$21440 ( \21817 , RIae781e8_105, \4686 );
nor \U$21441 ( \21818 , \21816 , \21817 );
and \U$21442 ( \21819 , \21818 , \4481 );
not \U$21443 ( \21820 , \21818 );
and \U$21444 ( \21821 , \21820 , \4482 );
nor \U$21445 ( \21822 , \21819 , \21821 );
nand \U$21446 ( \21823 , \21815 , \21822 );
nand \U$21447 ( \21824 , \21812 , \21823 );
xor \U$21448 ( \21825 , \21797 , \21824 );
and \U$21449 ( \21826 , \6941 , RIae77e28_97);
and \U$21450 ( \21827 , RIae78968_121, \6939 );
nor \U$21451 ( \21828 , \21826 , \21827 );
and \U$21452 ( \21829 , \21828 , \6314 );
not \U$21453 ( \21830 , \21828 );
and \U$21454 ( \21831 , \21830 , \6945 );
nor \U$21455 ( \21832 , \21829 , \21831 );
and \U$21456 ( \21833 , \5896 , RIae78530_112);
and \U$21457 ( \21834 , RIae77c48_93, \5894 );
nor \U$21458 ( \21835 , \21833 , \21834 );
and \U$21459 ( \21836 , \21835 , \5590 );
not \U$21460 ( \21837 , \21835 );
and \U$21461 ( \21838 , \21837 , \5589 );
nor \U$21462 ( \21839 , \21836 , \21838 );
xor \U$21463 ( \21840 , \21832 , \21839 );
and \U$21464 ( \21841 , \6172 , RIae77b58_91);
and \U$21465 ( \21842 , RIae77d38_95, \6170 );
nor \U$21466 ( \21843 , \21841 , \21842 );
and \U$21467 ( \21844 , \21843 , \6176 );
not \U$21468 ( \21845 , \21843 );
and \U$21469 ( \21846 , \21845 , \6175 );
nor \U$21470 ( \21847 , \21844 , \21846 );
and \U$21471 ( \21848 , \21840 , \21847 );
and \U$21472 ( \21849 , \21832 , \21839 );
or \U$21473 ( \21850 , \21848 , \21849 );
and \U$21474 ( \21851 , \21825 , \21850 );
and \U$21475 ( \21852 , \21797 , \21824 );
or \U$21476 ( \21853 , \21851 , \21852 );
and \U$21477 ( \21854 , \21772 , \21853 );
and \U$21478 ( \21855 , \21699 , \21771 );
or \U$21479 ( \21856 , \21854 , \21855 );
xor \U$21480 ( \21857 , \21620 , \21856 );
xor \U$21481 ( \21858 , \20900 , \789 );
xor \U$21482 ( \21859 , \21858 , \20908 );
xor \U$21483 ( \21860 , \21254 , \21256 );
xor \U$21484 ( \21861 , \21860 , \21259 );
and \U$21485 ( \21862 , \21859 , \21861 );
xor \U$21486 ( \21863 , \20999 , \21006 );
xor \U$21487 ( \21864 , \21863 , \21014 );
xor \U$21488 ( \21865 , \21225 , \21230 );
xor \U$21489 ( \21866 , \21864 , \21865 );
xor \U$21490 ( \21867 , \21254 , \21256 );
xor \U$21491 ( \21868 , \21867 , \21259 );
and \U$21492 ( \21869 , \21866 , \21868 );
and \U$21493 ( \21870 , \21859 , \21866 );
or \U$21494 ( \21871 , \21862 , \21869 , \21870 );
and \U$21495 ( \21872 , \21857 , \21871 );
and \U$21496 ( \21873 , \21620 , \21856 );
or \U$21497 ( \21874 , \21872 , \21873 );
xor \U$21498 ( \21875 , \21336 , \21417 );
xor \U$21499 ( \21876 , \21875 , \21497 );
xor \U$21500 ( \21877 , \21235 , \21251 );
xor \U$21501 ( \21878 , \21877 , \21262 );
and \U$21502 ( \21879 , \21876 , \21878 );
xor \U$21503 ( \21880 , \21874 , \21879 );
xor \U$21504 ( \21881 , \21290 , \21305 );
xor \U$21505 ( \21882 , \21881 , \21333 );
xor \U$21506 ( \21883 , \21443 , \21468 );
xor \U$21507 ( \21884 , \21883 , \21494 );
and \U$21508 ( \21885 , \21882 , \21884 );
xor \U$21509 ( \21886 , \20794 , \20801 );
xor \U$21510 ( \21887 , \21886 , \20809 );
xor \U$21511 ( \21888 , \21241 , \21246 );
xor \U$21512 ( \21889 , \21887 , \21888 );
xor \U$21513 ( \21890 , \21443 , \21468 );
xor \U$21514 ( \21891 , \21890 , \21494 );
and \U$21515 ( \21892 , \21889 , \21891 );
and \U$21516 ( \21893 , \21882 , \21889 );
or \U$21517 ( \21894 , \21885 , \21892 , \21893 );
xor \U$21518 ( \21895 , \21523 , \21525 );
xor \U$21519 ( \21896 , \21895 , \21528 );
and \U$21520 ( \21897 , \21894 , \21896 );
xor \U$21521 ( \21898 , \21065 , \21071 );
xor \U$21522 ( \21899 , \21898 , \21074 );
xor \U$21523 ( \21900 , \21505 , \21512 );
xor \U$21524 ( \21901 , \21899 , \21900 );
xor \U$21525 ( \21902 , \21523 , \21525 );
xor \U$21526 ( \21903 , \21902 , \21528 );
and \U$21527 ( \21904 , \21901 , \21903 );
and \U$21528 ( \21905 , \21894 , \21901 );
or \U$21529 ( \21906 , \21897 , \21904 , \21905 );
and \U$21530 ( \21907 , \21880 , \21906 );
and \U$21531 ( \21908 , \21874 , \21879 );
or \U$21532 ( \21909 , \21907 , \21908 );
xor \U$21533 ( \21910 , \21023 , \21037 );
xor \U$21534 ( \21911 , \21910 , \21080 );
xor \U$21535 ( \21912 , \21909 , \21911 );
xor \U$21536 ( \21913 , \21265 , \21500 );
xor \U$21537 ( \21914 , \21913 , \21517 );
xor \U$21538 ( \21915 , \21213 , \21217 );
xor \U$21539 ( \21916 , \21915 , \21220 );
and \U$21540 ( \21917 , \21914 , \21916 );
xor \U$21541 ( \21918 , \21531 , \21532 );
xor \U$21542 ( \21919 , \21918 , \21535 );
xor \U$21543 ( \21920 , \21213 , \21217 );
xor \U$21544 ( \21921 , \21920 , \21220 );
and \U$21545 ( \21922 , \21919 , \21921 );
and \U$21546 ( \21923 , \21914 , \21919 );
or \U$21547 ( \21924 , \21917 , \21922 , \21923 );
and \U$21548 ( \21925 , \21912 , \21924 );
and \U$21549 ( \21926 , \21909 , \21911 );
or \U$21550 ( \21927 , \21925 , \21926 );
and \U$21551 ( \21928 , \21573 , \21927 );
not \U$21552 ( \21929 , \21572 );
and \U$21553 ( \21930 , \21565 , \21929 );
nor \U$21554 ( \21931 , \21928 , \21930 );
nor \U$21555 ( \21932 , \21563 , \21931 );
and \U$21556 ( \21933 , \21558 , \21932 );
xor \U$21557 ( \21934 , \21932 , \21558 );
not \U$21558 ( \21935 , \21562 );
not \U$21559 ( \21936 , \21931 );
and \U$21560 ( \21937 , \21935 , \21936 );
and \U$21561 ( \21938 , \21562 , \21931 );
nor \U$21562 ( \21939 , \21937 , \21938 );
not \U$21563 ( \21940 , \21541 );
not \U$21564 ( \21941 , \21207 );
or \U$21565 ( \21942 , \21940 , \21941 );
or \U$21566 ( \21943 , \21207 , \21541 );
nand \U$21567 ( \21944 , \21942 , \21943 );
not \U$21568 ( \21945 , \21944 );
not \U$21569 ( \21946 , \21193 );
and \U$21570 ( \21947 , \21945 , \21946 );
and \U$21571 ( \21948 , \21944 , \21193 );
nor \U$21572 ( \21949 , \21947 , \21948 );
not \U$21573 ( \21950 , \21949 );
not \U$21574 ( \21951 , \21565 );
not \U$21575 ( \21952 , \21927 );
not \U$21576 ( \21953 , \21572 );
and \U$21577 ( \21954 , \21952 , \21953 );
and \U$21578 ( \21955 , \21927 , \21572 );
nor \U$21579 ( \21956 , \21954 , \21955 );
not \U$21580 ( \21957 , \21956 );
or \U$21581 ( \21958 , \21951 , \21957 );
or \U$21582 ( \21959 , \21956 , \21565 );
nand \U$21583 ( \21960 , \21958 , \21959 );
nand \U$21584 ( \21961 , \21950 , \21960 );
or \U$21585 ( \21962 , \21939 , \21961 );
xnor \U$21586 ( \21963 , \21961 , \21939 );
xor \U$21587 ( \21964 , \21699 , \21771 );
xor \U$21588 ( \21965 , \21964 , \21853 );
xor \U$21589 ( \21966 , \21593 , \21604 );
xor \U$21590 ( \21967 , \21966 , \21617 );
and \U$21591 ( \21968 , \21965 , \21967 );
xor \U$21592 ( \21969 , \21254 , \21256 );
xor \U$21593 ( \21970 , \21969 , \21259 );
xor \U$21594 ( \21971 , \21859 , \21866 );
xor \U$21595 ( \21972 , \21970 , \21971 );
xor \U$21596 ( \21973 , \21593 , \21604 );
xor \U$21597 ( \21974 , \21973 , \21617 );
and \U$21598 ( \21975 , \21972 , \21974 );
and \U$21599 ( \21976 , \21965 , \21972 );
or \U$21600 ( \21977 , \21968 , \21975 , \21976 );
and \U$21601 ( \21978 , \2607 , RIae76f28_65);
and \U$21602 ( \21979 , RIae76e38_63, \2605 );
nor \U$21603 ( \21980 , \21978 , \21979 );
and \U$21604 ( \21981 , \21980 , \2611 );
not \U$21605 ( \21982 , \21980 );
and \U$21606 ( \21983 , \21982 , \2397 );
nor \U$21607 ( \21984 , \21981 , \21983 );
not \U$21608 ( \21985 , \3089 );
and \U$21609 ( \21986 , \2783 , RIae76d48_61);
and \U$21610 ( \21987 , RIae76c58_59, \2781 );
nor \U$21611 ( \21988 , \21986 , \21987 );
not \U$21612 ( \21989 , \21988 );
or \U$21613 ( \21990 , \21985 , \21989 );
or \U$21614 ( \21991 , \21988 , \3089 );
nand \U$21615 ( \21992 , \21990 , \21991 );
xor \U$21616 ( \21993 , \21984 , \21992 );
not \U$21617 ( \21994 , \2774 );
and \U$21618 ( \21995 , \3214 , RIae77180_70);
and \U$21619 ( \21996 , RIae77018_67, \3212 );
nor \U$21620 ( \21997 , \21995 , \21996 );
not \U$21621 ( \21998 , \21997 );
or \U$21622 ( \21999 , \21994 , \21998 );
or \U$21623 ( \22000 , \21997 , \2774 );
nand \U$21624 ( \22001 , \21999 , \22000 );
and \U$21625 ( \22002 , \21993 , \22001 );
and \U$21626 ( \22003 , \21984 , \21992 );
or \U$21627 ( \22004 , \22002 , \22003 );
and \U$21628 ( \22005 , \2224 , RIae77798_83);
and \U$21629 ( \22006 , RIae77888_85, \2222 );
nor \U$21630 ( \22007 , \22005 , \22006 );
and \U$21631 ( \22008 , \22007 , \2061 );
not \U$21632 ( \22009 , \22007 );
and \U$21633 ( \22010 , \22009 , \2060 );
nor \U$21634 ( \22011 , \22008 , \22010 );
and \U$21635 ( \22012 , \1593 , RIae77720_82);
and \U$21636 ( \22013 , RIae773d8_75, \1591 );
nor \U$21637 ( \22014 , \22012 , \22013 );
and \U$21638 ( \22015 , \22014 , \1498 );
not \U$21639 ( \22016 , \22014 );
and \U$21640 ( \22017 , \22016 , \1488 );
nor \U$21641 ( \22018 , \22015 , \22017 );
xor \U$21642 ( \22019 , \22011 , \22018 );
and \U$21643 ( \22020 , \1939 , RIae77a68_89);
and \U$21644 ( \22021 , RIae77978_87, \1937 );
nor \U$21645 ( \22022 , \22020 , \22021 );
and \U$21646 ( \22023 , \22022 , \1735 );
not \U$21647 ( \22024 , \22022 );
and \U$21648 ( \22025 , \22024 , \1734 );
nor \U$21649 ( \22026 , \22023 , \22025 );
and \U$21650 ( \22027 , \22019 , \22026 );
and \U$21651 ( \22028 , \22011 , \22018 );
or \U$21652 ( \22029 , \22027 , \22028 );
xor \U$21653 ( \22030 , \22004 , \22029 );
xor \U$21654 ( \22031 , \21652 , \21657 );
xor \U$21655 ( \22032 , \22031 , \21665 );
and \U$21656 ( \22033 , \22030 , \22032 );
and \U$21657 ( \22034 , \22004 , \22029 );
or \U$21658 ( \22035 , \22033 , \22034 );
and \U$21659 ( \22036 , \12180 , RIae755d8_11);
and \U$21660 ( \22037 , RIae754e8_9, \12178 );
nor \U$21661 ( \22038 , \22036 , \22037 );
and \U$21662 ( \22039 , \22038 , \12184 );
not \U$21663 ( \22040 , \22038 );
and \U$21664 ( \22041 , \22040 , \11827 );
nor \U$21665 ( \22042 , \22039 , \22041 );
and \U$21666 ( \22043 , \11470 , RIae75c68_25);
and \U$21667 ( \22044 , RIae75d58_27, \11468 );
nor \U$21668 ( \22045 , \22043 , \22044 );
and \U$21669 ( \22046 , \22045 , \10936 );
not \U$21670 ( \22047 , \22045 );
and \U$21671 ( \22048 , \22047 , \11474 );
nor \U$21672 ( \22049 , \22046 , \22048 );
xor \U$21673 ( \22050 , \22042 , \22049 );
and \U$21674 ( \22051 , \13059 , RIae757b8_15);
and \U$21675 ( \22052 , RIae756c8_13, \13057 );
nor \U$21676 ( \22053 , \22051 , \22052 );
and \U$21677 ( \22054 , \22053 , \13063 );
not \U$21678 ( \22055 , \22053 );
and \U$21679 ( \22056 , \22055 , \12718 );
nor \U$21680 ( \22057 , \22054 , \22056 );
and \U$21681 ( \22058 , \22050 , \22057 );
and \U$21682 ( \22059 , \22042 , \22049 );
or \U$21683 ( \22060 , \22058 , \22059 );
and \U$21684 ( \22061 , \14059 , RIae75218_3);
and \U$21685 ( \22062 , RIae75128_1, \14057 );
nor \U$21686 ( \22063 , \22061 , \22062 );
and \U$21687 ( \22064 , \22063 , \13502 );
not \U$21688 ( \22065 , \22063 );
and \U$21689 ( \22066 , \22065 , \14063 );
nor \U$21690 ( \22067 , \22064 , \22066 );
and \U$21691 ( \22068 , \15726 , RIae763e8_41);
and \U$21692 ( \22069 , RIae7aab0_192, RIae764d8_43);
nor \U$21693 ( \22070 , \22068 , \22069 );
and \U$21694 ( \22071 , \22070 , \14959 );
not \U$21695 ( \22072 , \22070 );
and \U$21696 ( \22073 , \22072 , RIae7aa38_191);
nor \U$21697 ( \22074 , \22071 , \22073 );
xor \U$21698 ( \22075 , \22067 , \22074 );
and \U$21699 ( \22076 , \14964 , RIae75308_5);
and \U$21700 ( \22077 , RIae753f8_7, \14962 );
nor \U$21701 ( \22078 , \22076 , \22077 );
and \U$21702 ( \22079 , \22078 , \14463 );
not \U$21703 ( \22080 , \22078 );
and \U$21704 ( \22081 , \22080 , \14462 );
nor \U$21705 ( \22082 , \22079 , \22081 );
and \U$21706 ( \22083 , \22075 , \22082 );
and \U$21707 ( \22084 , \22067 , \22074 );
or \U$21708 ( \22085 , \22083 , \22084 );
xor \U$21709 ( \22086 , \22060 , \22085 );
and \U$21710 ( \22087 , \9760 , RIae75998_19);
and \U$21711 ( \22088 , RIae758a8_17, \9758 );
nor \U$21712 ( \22089 , \22087 , \22088 );
and \U$21713 ( \22090 , \22089 , \9273 );
not \U$21714 ( \22091 , \22089 );
and \U$21715 ( \22092 , \22091 , \9272 );
nor \U$21716 ( \22093 , \22090 , \22092 );
and \U$21717 ( \22094 , \8966 , RIae75b78_23);
and \U$21718 ( \22095 , RIae75a88_21, \8964 );
nor \U$21719 ( \22096 , \22094 , \22095 );
and \U$21720 ( \22097 , \22096 , \8799 );
not \U$21721 ( \22098 , \22096 );
and \U$21722 ( \22099 , \22098 , \8789 );
nor \U$21723 ( \22100 , \22097 , \22099 );
xor \U$21724 ( \22101 , \22093 , \22100 );
and \U$21725 ( \22102 , \10548 , RIae75f38_31);
and \U$21726 ( \22103 , RIae75e48_29, \10546 );
nor \U$21727 ( \22104 , \22102 , \22103 );
and \U$21728 ( \22105 , \22104 , \10421 );
not \U$21729 ( \22106 , \22104 );
and \U$21730 ( \22107 , \22106 , \10118 );
nor \U$21731 ( \22108 , \22105 , \22107 );
and \U$21732 ( \22109 , \22101 , \22108 );
and \U$21733 ( \22110 , \22093 , \22100 );
or \U$21734 ( \22111 , \22109 , \22110 );
and \U$21735 ( \22112 , \22086 , \22111 );
and \U$21736 ( \22113 , \22060 , \22085 );
or \U$21737 ( \22114 , \22112 , \22113 );
xor \U$21738 ( \22115 , \22035 , \22114 );
and \U$21739 ( \22116 , \5399 , RIae781e8_105);
and \U$21740 ( \22117 , RIae785a8_113, \5397 );
nor \U$21741 ( \22118 , \22116 , \22117 );
and \U$21742 ( \22119 , \22118 , \5016 );
not \U$21743 ( \22120 , \22118 );
and \U$21744 ( \22121 , \22120 , \5403 );
nor \U$21745 ( \22122 , \22119 , \22121 );
and \U$21746 ( \22123 , \5896 , RIae783c8_109);
and \U$21747 ( \22124 , RIae78530_112, \5894 );
nor \U$21748 ( \22125 , \22123 , \22124 );
and \U$21749 ( \22126 , \22125 , \5590 );
not \U$21750 ( \22127 , \22125 );
and \U$21751 ( \22128 , \22127 , \5589 );
nor \U$21752 ( \22129 , \22126 , \22128 );
xor \U$21753 ( \22130 , \22122 , \22129 );
and \U$21754 ( \22131 , \6172 , RIae77c48_93);
and \U$21755 ( \22132 , RIae77b58_91, \6170 );
nor \U$21756 ( \22133 , \22131 , \22132 );
and \U$21757 ( \22134 , \22133 , \6176 );
not \U$21758 ( \22135 , \22133 );
and \U$21759 ( \22136 , \22135 , \6175 );
nor \U$21760 ( \22137 , \22134 , \22136 );
and \U$21761 ( \22138 , \22130 , \22137 );
and \U$21762 ( \22139 , \22122 , \22129 );
or \U$21763 ( \22140 , \22138 , \22139 );
and \U$21764 ( \22141 , \3730 , RIae771f8_71);
and \U$21765 ( \22142 , RIae772e8_73, \3728 );
nor \U$21766 ( \22143 , \22141 , \22142 );
and \U$21767 ( \22144 , \22143 , \3732 );
not \U$21768 ( \22145 , \22143 );
and \U$21769 ( \22146 , \22145 , \3422 );
nor \U$21770 ( \22147 , \22144 , \22146 );
and \U$21771 ( \22148 , \4247 , RIae782d8_107);
and \U$21772 ( \22149 , RIae780f8_103, \4245 );
nor \U$21773 ( \22150 , \22148 , \22149 );
and \U$21774 ( \22151 , \22150 , \3989 );
not \U$21775 ( \22152 , \22150 );
and \U$21776 ( \22153 , \22152 , \4251 );
nor \U$21777 ( \22154 , \22151 , \22153 );
xor \U$21778 ( \22155 , \22147 , \22154 );
and \U$21779 ( \22156 , \4688 , RIae77f18_99);
and \U$21780 ( \22157 , RIae78008_101, \4686 );
nor \U$21781 ( \22158 , \22156 , \22157 );
and \U$21782 ( \22159 , \22158 , \4481 );
not \U$21783 ( \22160 , \22158 );
and \U$21784 ( \22161 , \22160 , \4482 );
nor \U$21785 ( \22162 , \22159 , \22161 );
and \U$21786 ( \22163 , \22155 , \22162 );
and \U$21787 ( \22164 , \22147 , \22154 );
or \U$21788 ( \22165 , \22163 , \22164 );
xor \U$21789 ( \22166 , \22140 , \22165 );
and \U$21790 ( \22167 , \8371 , RIae78788_117);
and \U$21791 ( \22168 , RIae78698_115, \8369 );
nor \U$21792 ( \22169 , \22167 , \22168 );
and \U$21793 ( \22170 , \22169 , \8020 );
not \U$21794 ( \22171 , \22169 );
and \U$21795 ( \22172 , \22171 , \8019 );
nor \U$21796 ( \22173 , \22170 , \22172 );
and \U$21797 ( \22174 , \6941 , RIae77d38_95);
and \U$21798 ( \22175 , RIae77e28_97, \6939 );
nor \U$21799 ( \22176 , \22174 , \22175 );
and \U$21800 ( \22177 , \22176 , \6314 );
not \U$21801 ( \22178 , \22176 );
and \U$21802 ( \22179 , \22178 , \6945 );
nor \U$21803 ( \22180 , \22177 , \22179 );
xor \U$21804 ( \22181 , \22173 , \22180 );
and \U$21805 ( \22182 , \7633 , RIae78968_121);
and \U$21806 ( \22183 , RIae78878_119, \7631 );
nor \U$21807 ( \22184 , \22182 , \22183 );
and \U$21808 ( \22185 , \22184 , \7206 );
not \U$21809 ( \22186 , \22184 );
and \U$21810 ( \22187 , \22186 , \7205 );
nor \U$21811 ( \22188 , \22185 , \22187 );
and \U$21812 ( \22189 , \22181 , \22188 );
and \U$21813 ( \22190 , \22173 , \22180 );
or \U$21814 ( \22191 , \22189 , \22190 );
and \U$21815 ( \22192 , \22166 , \22191 );
and \U$21816 ( \22193 , \22140 , \22165 );
or \U$21817 ( \22194 , \22192 , \22193 );
and \U$21818 ( \22195 , \22115 , \22194 );
and \U$21819 ( \22196 , \22035 , \22114 );
nor \U$21820 ( \22197 , \22195 , \22196 );
xor \U$21821 ( \22198 , \21779 , \21786 );
xor \U$21822 ( \22199 , \22198 , \21794 );
xor \U$21823 ( \22200 , \21832 , \21839 );
xor \U$21824 ( \22201 , \22200 , \21847 );
and \U$21825 ( \22202 , \22199 , \22201 );
xor \U$21826 ( \22203 , \21706 , \21713 );
xor \U$21827 ( \22204 , \22203 , \21721 );
xor \U$21828 ( \22205 , \21832 , \21839 );
xor \U$21829 ( \22206 , \22205 , \21847 );
and \U$21830 ( \22207 , \22204 , \22206 );
and \U$21831 ( \22208 , \22199 , \22204 );
or \U$21832 ( \22209 , \22202 , \22207 , \22208 );
not \U$21833 ( \22210 , \22209 );
xor \U$21834 ( \22211 , \21750 , \21757 );
xor \U$21835 ( \22212 , \22211 , \21765 );
not \U$21836 ( \22213 , \22212 );
xor \U$21837 ( \22214 , \21731 , \1142 );
xor \U$21838 ( \22215 , \22214 , \21739 );
nand \U$21839 ( \22216 , \22213 , \22215 );
xor \U$21840 ( \22217 , \22210 , \22216 );
xor \U$21841 ( \22218 , \21627 , \21634 );
xor \U$21842 ( \22219 , \22218 , \21642 );
not \U$21843 ( \22220 , \22219 );
not \U$21844 ( \22221 , \21811 );
not \U$21845 ( \22222 , \21822 );
or \U$21846 ( \22223 , \22221 , \22222 );
or \U$21847 ( \22224 , \21811 , \21822 );
nand \U$21848 ( \22225 , \22223 , \22224 );
not \U$21849 ( \22226 , \22225 );
not \U$21850 ( \22227 , \21804 );
and \U$21851 ( \22228 , \22226 , \22227 );
and \U$21852 ( \22229 , \22225 , \21804 );
nor \U$21853 ( \22230 , \22228 , \22229 );
not \U$21854 ( \22231 , \22230 );
and \U$21855 ( \22232 , \22220 , \22231 );
and \U$21856 ( \22233 , \22230 , \22219 );
xor \U$21857 ( \22234 , \21677 , \21684 );
xor \U$21858 ( \22235 , \22234 , \21693 );
nor \U$21859 ( \22236 , \22233 , \22235 );
nor \U$21860 ( \22237 , \22232 , \22236 );
and \U$21861 ( \22238 , \22217 , \22237 );
and \U$21862 ( \22239 , \22210 , \22216 );
or \U$21863 ( \22240 , \22238 , \22239 );
xor \U$21864 ( \22241 , \22197 , \22240 );
xor \U$21865 ( \22242 , \21425 , \21432 );
xor \U$21866 ( \22243 , \22242 , \21440 );
xor \U$21867 ( \22244 , \21607 , \21612 );
xor \U$21868 ( \22245 , \22243 , \22244 );
xnor \U$21869 ( \22246 , \21597 , \21602 );
not \U$21870 ( \22247 , \22246 );
not \U$21871 ( \22248 , \21594 );
and \U$21872 ( \22249 , \22247 , \22248 );
and \U$21873 ( \22250 , \22246 , \21594 );
nor \U$21874 ( \22251 , \22249 , \22250 );
not \U$21875 ( \22252 , \22251 );
and \U$21876 ( \22253 , \22245 , \22252 );
not \U$21877 ( \22254 , \22252 );
not \U$21878 ( \22255 , \22245 );
and \U$21879 ( \22256 , \22254 , \22255 );
not \U$21880 ( \22257 , \21591 );
not \U$21881 ( \22258 , \21575 );
or \U$21882 ( \22259 , \22257 , \22258 );
or \U$21883 ( \22260 , \21575 , \21591 );
nand \U$21884 ( \22261 , \22259 , \22260 );
not \U$21885 ( \22262 , \22261 );
not \U$21886 ( \22263 , \21585 );
and \U$21887 ( \22264 , \22262 , \22263 );
and \U$21888 ( \22265 , \22261 , \21585 );
nor \U$21889 ( \22266 , \22264 , \22265 );
nor \U$21890 ( \22267 , \22256 , \22266 );
nor \U$21891 ( \22268 , \22253 , \22267 );
and \U$21892 ( \22269 , \22241 , \22268 );
and \U$21893 ( \22270 , \22197 , \22240 );
nor \U$21894 ( \22271 , \22269 , \22270 );
xor \U$21895 ( \22272 , \21977 , \22271 );
xor \U$21896 ( \22273 , \21724 , \21742 );
xor \U$21897 ( \22274 , \22273 , \21768 );
xor \U$21898 ( \22275 , \21797 , \21824 );
xor \U$21899 ( \22276 , \22275 , \21850 );
xor \U$21900 ( \22277 , \22274 , \22276 );
xor \U$21901 ( \22278 , \21645 , \21668 );
xor \U$21902 ( \22279 , \22278 , \21696 );
and \U$21903 ( \22280 , \22277 , \22279 );
and \U$21904 ( \22281 , \22274 , \22276 );
or \U$21905 ( \22282 , \22280 , \22281 );
xor \U$21906 ( \22283 , \21361 , \21386 );
xor \U$21907 ( \22284 , \22283 , \21414 );
xor \U$21908 ( \22285 , \22282 , \22284 );
xor \U$21909 ( \22286 , \21443 , \21468 );
xor \U$21910 ( \22287 , \22286 , \21494 );
xor \U$21911 ( \22288 , \21882 , \21889 );
xor \U$21912 ( \22289 , \22287 , \22288 );
and \U$21913 ( \22290 , \22285 , \22289 );
and \U$21914 ( \22291 , \22282 , \22284 );
or \U$21915 ( \22292 , \22290 , \22291 );
and \U$21916 ( \22293 , \22272 , \22292 );
and \U$21917 ( \22294 , \21977 , \22271 );
or \U$21918 ( \22295 , \22293 , \22294 );
xor \U$21919 ( \22296 , \21876 , \21878 );
xor \U$21920 ( \22297 , \21620 , \21856 );
xor \U$21921 ( \22298 , \22297 , \21871 );
and \U$21922 ( \22299 , \22296 , \22298 );
xor \U$21923 ( \22300 , \21523 , \21525 );
xor \U$21924 ( \22301 , \22300 , \21528 );
xor \U$21925 ( \22302 , \21894 , \21901 );
xor \U$21926 ( \22303 , \22301 , \22302 );
xor \U$21927 ( \22304 , \21620 , \21856 );
xor \U$21928 ( \22305 , \22304 , \21871 );
and \U$21929 ( \22306 , \22303 , \22305 );
and \U$21930 ( \22307 , \22296 , \22303 );
or \U$21931 ( \22308 , \22299 , \22306 , \22307 );
xor \U$21932 ( \22309 , \22295 , \22308 );
xor \U$21933 ( \22310 , \21213 , \21217 );
xor \U$21934 ( \22311 , \22310 , \21220 );
xor \U$21935 ( \22312 , \21914 , \21919 );
xor \U$21936 ( \22313 , \22311 , \22312 );
and \U$21937 ( \22314 , \22309 , \22313 );
and \U$21938 ( \22315 , \22295 , \22308 );
or \U$21939 ( \22316 , \22314 , \22315 );
xor \U$21940 ( \22317 , \21909 , \21911 );
xor \U$21941 ( \22318 , \22317 , \21924 );
xnor \U$21942 ( \22319 , \22316 , \22318 );
not \U$21943 ( \22320 , \22319 );
not \U$21944 ( \22321 , \21571 );
not \U$21945 ( \22322 , \21568 );
or \U$21946 ( \22323 , \22321 , \22322 );
or \U$21947 ( \22324 , \21568 , \21571 );
nand \U$21948 ( \22325 , \22323 , \22324 );
not \U$21949 ( \22326 , \22325 );
and \U$21950 ( \22327 , \22320 , \22326 );
and \U$21951 ( \22328 , \22319 , \22325 );
nor \U$21952 ( \22329 , \22327 , \22328 );
xor \U$21953 ( \22330 , \22140 , \22165 );
xor \U$21954 ( \22331 , \22330 , \22191 );
xor \U$21955 ( \22332 , \22004 , \22029 );
xor \U$21956 ( \22333 , \22332 , \22032 );
xor \U$21957 ( \22334 , \22331 , \22333 );
xor \U$21958 ( \22335 , \22060 , \22085 );
xor \U$21959 ( \22336 , \22335 , \22111 );
and \U$21960 ( \22337 , \22334 , \22336 );
and \U$21961 ( \22338 , \22331 , \22333 );
or \U$21962 ( \22339 , \22337 , \22338 );
xor \U$21963 ( \22340 , \22274 , \22276 );
xor \U$21964 ( \22341 , \22340 , \22279 );
and \U$21965 ( \22342 , \22339 , \22341 );
not \U$21966 ( \22343 , \22251 );
not \U$21967 ( \22344 , \22245 );
not \U$21968 ( \22345 , \22266 );
or \U$21969 ( \22346 , \22344 , \22345 );
or \U$21970 ( \22347 , \22266 , \22245 );
nand \U$21971 ( \22348 , \22346 , \22347 );
not \U$21972 ( \22349 , \22348 );
or \U$21973 ( \22350 , \22343 , \22349 );
or \U$21974 ( \22351 , \22348 , \22251 );
nand \U$21975 ( \22352 , \22350 , \22351 );
xor \U$21976 ( \22353 , \22274 , \22276 );
xor \U$21977 ( \22354 , \22353 , \22279 );
and \U$21978 ( \22355 , \22352 , \22354 );
and \U$21979 ( \22356 , \22339 , \22352 );
or \U$21980 ( \22357 , \22342 , \22355 , \22356 );
xor \U$21981 ( \22358 , \22147 , \22154 );
xor \U$21982 ( \22359 , \22358 , \22162 );
xor \U$21983 ( \22360 , \22011 , \22018 );
xor \U$21984 ( \22361 , \22360 , \22026 );
xor \U$21985 ( \22362 , \22359 , \22361 );
xor \U$21986 ( \22363 , \21984 , \21992 );
xor \U$21987 ( \22364 , \22363 , \22001 );
and \U$21988 ( \22365 , \22362 , \22364 );
and \U$21989 ( \22366 , \22359 , \22361 );
or \U$21990 ( \22367 , \22365 , \22366 );
xor \U$21991 ( \22368 , \22042 , \22049 );
xor \U$21992 ( \22369 , \22368 , \22057 );
xor \U$21993 ( \22370 , \22067 , \22074 );
xor \U$21994 ( \22371 , \22370 , \22082 );
and \U$21995 ( \22372 , \22369 , \22371 );
xor \U$21996 ( \22373 , \22367 , \22372 );
xor \U$21997 ( \22374 , \22122 , \22129 );
xor \U$21998 ( \22375 , \22374 , \22137 );
xor \U$21999 ( \22376 , \22173 , \22180 );
xor \U$22000 ( \22377 , \22376 , \22188 );
and \U$22001 ( \22378 , \22375 , \22377 );
xor \U$22002 ( \22379 , \22093 , \22100 );
xor \U$22003 ( \22380 , \22379 , \22108 );
xor \U$22004 ( \22381 , \22173 , \22180 );
xor \U$22005 ( \22382 , \22381 , \22188 );
and \U$22006 ( \22383 , \22380 , \22382 );
and \U$22007 ( \22384 , \22375 , \22380 );
or \U$22008 ( \22385 , \22378 , \22383 , \22384 );
and \U$22009 ( \22386 , \22373 , \22385 );
and \U$22010 ( \22387 , \22367 , \22372 );
or \U$22011 ( \22388 , \22386 , \22387 );
and \U$22012 ( \22389 , \1939 , RIae773d8_75);
and \U$22013 ( \22390 , RIae77a68_89, \1937 );
nor \U$22014 ( \22391 , \22389 , \22390 );
and \U$22015 ( \22392 , \22391 , \1735 );
not \U$22016 ( \22393 , \22391 );
and \U$22017 ( \22394 , \22393 , \1734 );
nor \U$22018 ( \22395 , \22392 , \22394 );
and \U$22019 ( \22396 , \2224 , RIae77978_87);
and \U$22020 ( \22397 , RIae77798_83, \2222 );
nor \U$22021 ( \22398 , \22396 , \22397 );
and \U$22022 ( \22399 , \22398 , \2061 );
not \U$22023 ( \22400 , \22398 );
and \U$22024 ( \22401 , \22400 , \2060 );
nor \U$22025 ( \22402 , \22399 , \22401 );
xor \U$22026 ( \22403 , \22395 , \22402 );
and \U$22027 ( \22404 , \2607 , RIae77888_85);
and \U$22028 ( \22405 , RIae76f28_65, \2605 );
nor \U$22029 ( \22406 , \22404 , \22405 );
and \U$22030 ( \22407 , \22406 , \2611 );
not \U$22031 ( \22408 , \22406 );
and \U$22032 ( \22409 , \22408 , \2397 );
nor \U$22033 ( \22410 , \22407 , \22409 );
and \U$22034 ( \22411 , \22403 , \22410 );
and \U$22035 ( \22412 , \22395 , \22402 );
or \U$22036 ( \22413 , \22411 , \22412 );
and \U$22037 ( \22414 , \1376 , RIae775b8_79);
and \U$22038 ( \22415 , RIae774c8_77, \1374 );
nor \U$22039 ( \22416 , \22414 , \22415 );
and \U$22040 ( \22417 , \22416 , \1380 );
not \U$22041 ( \22418 , \22416 );
and \U$22042 ( \22419 , \22418 , \1261 );
nor \U$22043 ( \22420 , \22417 , \22419 );
xor \U$22044 ( \22421 , \22413 , \22420 );
not \U$22045 ( \22422 , \2774 );
and \U$22046 ( \22423 , \3214 , RIae76c58_59);
and \U$22047 ( \22424 , RIae77180_70, \3212 );
nor \U$22048 ( \22425 , \22423 , \22424 );
not \U$22049 ( \22426 , \22425 );
or \U$22050 ( \22427 , \22422 , \22426 );
or \U$22051 ( \22428 , \22425 , \2774 );
nand \U$22052 ( \22429 , \22427 , \22428 );
not \U$22053 ( \22430 , \2789 );
and \U$22054 ( \22431 , \2783 , RIae76e38_63);
and \U$22055 ( \22432 , RIae76d48_61, \2781 );
nor \U$22056 ( \22433 , \22431 , \22432 );
not \U$22057 ( \22434 , \22433 );
or \U$22058 ( \22435 , \22430 , \22434 );
or \U$22059 ( \22436 , \22433 , \2789 );
nand \U$22060 ( \22437 , \22435 , \22436 );
xor \U$22061 ( \22438 , \22429 , \22437 );
and \U$22062 ( \22439 , \3730 , RIae77018_67);
and \U$22063 ( \22440 , RIae771f8_71, \3728 );
nor \U$22064 ( \22441 , \22439 , \22440 );
and \U$22065 ( \22442 , \22441 , \3732 );
not \U$22066 ( \22443 , \22441 );
and \U$22067 ( \22444 , \22443 , \3422 );
nor \U$22068 ( \22445 , \22442 , \22444 );
and \U$22069 ( \22446 , \22438 , \22445 );
and \U$22070 ( \22447 , \22429 , \22437 );
or \U$22071 ( \22448 , \22446 , \22447 );
and \U$22072 ( \22449 , \22421 , \22448 );
and \U$22073 ( \22450 , \22413 , \22420 );
or \U$22074 ( \22451 , \22449 , \22450 );
and \U$22075 ( \22452 , \12180 , RIae75d58_27);
and \U$22076 ( \22453 , RIae755d8_11, \12178 );
nor \U$22077 ( \22454 , \22452 , \22453 );
and \U$22078 ( \22455 , \22454 , \12184 );
not \U$22079 ( \22456 , \22454 );
and \U$22080 ( \22457 , \22456 , \11827 );
nor \U$22081 ( \22458 , \22455 , \22457 );
and \U$22082 ( \22459 , \13059 , RIae754e8_9);
and \U$22083 ( \22460 , RIae757b8_15, \13057 );
nor \U$22084 ( \22461 , \22459 , \22460 );
and \U$22085 ( \22462 , \22461 , \13063 );
not \U$22086 ( \22463 , \22461 );
and \U$22087 ( \22464 , \22463 , \12718 );
nor \U$22088 ( \22465 , \22462 , \22464 );
xor \U$22089 ( \22466 , \22458 , \22465 );
and \U$22090 ( \22467 , \14059 , RIae756c8_13);
and \U$22091 ( \22468 , RIae75218_3, \14057 );
nor \U$22092 ( \22469 , \22467 , \22468 );
and \U$22093 ( \22470 , \22469 , \13502 );
not \U$22094 ( \22471 , \22469 );
and \U$22095 ( \22472 , \22471 , \14063 );
nor \U$22096 ( \22473 , \22470 , \22472 );
and \U$22097 ( \22474 , \22466 , \22473 );
and \U$22098 ( \22475 , \22458 , \22465 );
or \U$22099 ( \22476 , \22474 , \22475 );
and \U$22100 ( \22477 , \15726 , RIae753f8_7);
and \U$22101 ( \22478 , RIae7aab0_192, RIae763e8_41);
nor \U$22102 ( \22479 , \22477 , \22478 );
and \U$22103 ( \22480 , \22479 , \14959 );
not \U$22104 ( \22481 , \22479 );
and \U$22105 ( \22482 , \22481 , RIae7aa38_191);
nor \U$22106 ( \22483 , \22480 , \22482 );
xor \U$22107 ( \22484 , \22483 , \1261 );
and \U$22108 ( \22485 , \14964 , RIae75128_1);
and \U$22109 ( \22486 , RIae75308_5, \14962 );
nor \U$22110 ( \22487 , \22485 , \22486 );
and \U$22111 ( \22488 , \22487 , \14463 );
not \U$22112 ( \22489 , \22487 );
and \U$22113 ( \22490 , \22489 , \14462 );
nor \U$22114 ( \22491 , \22488 , \22490 );
and \U$22115 ( \22492 , \22484 , \22491 );
and \U$22116 ( \22493 , \22483 , \1261 );
or \U$22117 ( \22494 , \22492 , \22493 );
xor \U$22118 ( \22495 , \22476 , \22494 );
and \U$22119 ( \22496 , \9760 , RIae75a88_21);
and \U$22120 ( \22497 , RIae75998_19, \9758 );
nor \U$22121 ( \22498 , \22496 , \22497 );
and \U$22122 ( \22499 , \22498 , \9273 );
not \U$22123 ( \22500 , \22498 );
and \U$22124 ( \22501 , \22500 , \9764 );
nor \U$22125 ( \22502 , \22499 , \22501 );
and \U$22126 ( \22503 , \10548 , RIae758a8_17);
and \U$22127 ( \22504 , RIae75f38_31, \10546 );
nor \U$22128 ( \22505 , \22503 , \22504 );
and \U$22129 ( \22506 , \22505 , \10421 );
not \U$22130 ( \22507 , \22505 );
and \U$22131 ( \22508 , \22507 , \10118 );
nor \U$22132 ( \22509 , \22506 , \22508 );
xor \U$22133 ( \22510 , \22502 , \22509 );
and \U$22134 ( \22511 , \11470 , RIae75e48_29);
and \U$22135 ( \22512 , RIae75c68_25, \11468 );
nor \U$22136 ( \22513 , \22511 , \22512 );
and \U$22137 ( \22514 , \22513 , \10936 );
not \U$22138 ( \22515 , \22513 );
and \U$22139 ( \22516 , \22515 , \11474 );
nor \U$22140 ( \22517 , \22514 , \22516 );
and \U$22141 ( \22518 , \22510 , \22517 );
and \U$22142 ( \22519 , \22502 , \22509 );
or \U$22143 ( \22520 , \22518 , \22519 );
and \U$22144 ( \22521 , \22495 , \22520 );
and \U$22145 ( \22522 , \22476 , \22494 );
or \U$22146 ( \22523 , \22521 , \22522 );
xor \U$22147 ( \22524 , \22451 , \22523 );
and \U$22148 ( \22525 , \7633 , RIae77e28_97);
and \U$22149 ( \22526 , RIae78968_121, \7631 );
nor \U$22150 ( \22527 , \22525 , \22526 );
and \U$22151 ( \22528 , \22527 , \7206 );
not \U$22152 ( \22529 , \22527 );
and \U$22153 ( \22530 , \22529 , \7205 );
nor \U$22154 ( \22531 , \22528 , \22530 );
and \U$22155 ( \22532 , \8371 , RIae78878_119);
and \U$22156 ( \22533 , RIae78788_117, \8369 );
nor \U$22157 ( \22534 , \22532 , \22533 );
and \U$22158 ( \22535 , \22534 , \8020 );
not \U$22159 ( \22536 , \22534 );
and \U$22160 ( \22537 , \22536 , \8019 );
nor \U$22161 ( \22538 , \22535 , \22537 );
xor \U$22162 ( \22539 , \22531 , \22538 );
and \U$22163 ( \22540 , \8966 , RIae78698_115);
and \U$22164 ( \22541 , RIae75b78_23, \8964 );
nor \U$22165 ( \22542 , \22540 , \22541 );
and \U$22166 ( \22543 , \22542 , \8799 );
not \U$22167 ( \22544 , \22542 );
and \U$22168 ( \22545 , \22544 , \8789 );
nor \U$22169 ( \22546 , \22543 , \22545 );
and \U$22170 ( \22547 , \22539 , \22546 );
and \U$22171 ( \22548 , \22531 , \22538 );
or \U$22172 ( \22549 , \22547 , \22548 );
and \U$22173 ( \22550 , \4247 , RIae772e8_73);
and \U$22174 ( \22551 , RIae782d8_107, \4245 );
nor \U$22175 ( \22552 , \22550 , \22551 );
and \U$22176 ( \22553 , \22552 , \3989 );
not \U$22177 ( \22554 , \22552 );
and \U$22178 ( \22555 , \22554 , \4251 );
nor \U$22179 ( \22556 , \22553 , \22555 );
and \U$22180 ( \22557 , \4688 , RIae780f8_103);
and \U$22181 ( \22558 , RIae77f18_99, \4686 );
nor \U$22182 ( \22559 , \22557 , \22558 );
and \U$22183 ( \22560 , \22559 , \4481 );
not \U$22184 ( \22561 , \22559 );
and \U$22185 ( \22562 , \22561 , \4482 );
nor \U$22186 ( \22563 , \22560 , \22562 );
xor \U$22187 ( \22564 , \22556 , \22563 );
and \U$22188 ( \22565 , \5399 , RIae78008_101);
and \U$22189 ( \22566 , RIae781e8_105, \5397 );
nor \U$22190 ( \22567 , \22565 , \22566 );
and \U$22191 ( \22568 , \22567 , \5016 );
not \U$22192 ( \22569 , \22567 );
and \U$22193 ( \22570 , \22569 , \5403 );
nor \U$22194 ( \22571 , \22568 , \22570 );
and \U$22195 ( \22572 , \22564 , \22571 );
and \U$22196 ( \22573 , \22556 , \22563 );
or \U$22197 ( \22574 , \22572 , \22573 );
xor \U$22198 ( \22575 , \22549 , \22574 );
and \U$22199 ( \22576 , \6172 , RIae78530_112);
and \U$22200 ( \22577 , RIae77c48_93, \6170 );
nor \U$22201 ( \22578 , \22576 , \22577 );
and \U$22202 ( \22579 , \22578 , \6176 );
not \U$22203 ( \22580 , \22578 );
and \U$22204 ( \22581 , \22580 , \6175 );
nor \U$22205 ( \22582 , \22579 , \22581 );
and \U$22206 ( \22583 , \5896 , RIae785a8_113);
and \U$22207 ( \22584 , RIae783c8_109, \5894 );
nor \U$22208 ( \22585 , \22583 , \22584 );
and \U$22209 ( \22586 , \22585 , \5590 );
not \U$22210 ( \22587 , \22585 );
and \U$22211 ( \22588 , \22587 , \5589 );
nor \U$22212 ( \22589 , \22586 , \22588 );
xor \U$22213 ( \22590 , \22582 , \22589 );
and \U$22214 ( \22591 , \6941 , RIae77b58_91);
and \U$22215 ( \22592 , RIae77d38_95, \6939 );
nor \U$22216 ( \22593 , \22591 , \22592 );
and \U$22217 ( \22594 , \22593 , \6314 );
not \U$22218 ( \22595 , \22593 );
and \U$22219 ( \22596 , \22595 , \6945 );
nor \U$22220 ( \22597 , \22594 , \22596 );
and \U$22221 ( \22598 , \22590 , \22597 );
and \U$22222 ( \22599 , \22582 , \22589 );
or \U$22223 ( \22600 , \22598 , \22599 );
and \U$22224 ( \22601 , \22575 , \22600 );
and \U$22225 ( \22602 , \22549 , \22574 );
or \U$22226 ( \22603 , \22601 , \22602 );
and \U$22227 ( \22604 , \22524 , \22603 );
and \U$22228 ( \22605 , \22451 , \22523 );
or \U$22229 ( \22606 , \22604 , \22605 );
xor \U$22230 ( \22607 , \22388 , \22606 );
not \U$22231 ( \22608 , \22219 );
xor \U$22232 ( \22609 , \22235 , \22230 );
not \U$22233 ( \22610 , \22609 );
or \U$22234 ( \22611 , \22608 , \22610 );
or \U$22235 ( \22612 , \22609 , \22219 );
nand \U$22236 ( \22613 , \22611 , \22612 );
not \U$22237 ( \22614 , \22212 );
not \U$22238 ( \22615 , \22215 );
or \U$22239 ( \22616 , \22614 , \22615 );
or \U$22240 ( \22617 , \22215 , \22212 );
nand \U$22241 ( \22618 , \22616 , \22617 );
xor \U$22242 ( \22619 , \22613 , \22618 );
xor \U$22243 ( \22620 , \21832 , \21839 );
xor \U$22244 ( \22621 , \22620 , \21847 );
xor \U$22245 ( \22622 , \22199 , \22204 );
xor \U$22246 ( \22623 , \22621 , \22622 );
and \U$22247 ( \22624 , \22619 , \22623 );
and \U$22248 ( \22625 , \22613 , \22618 );
or \U$22249 ( \22626 , \22624 , \22625 );
and \U$22250 ( \22627 , \22607 , \22626 );
and \U$22251 ( \22628 , \22388 , \22606 );
or \U$22252 ( \22629 , \22627 , \22628 );
xor \U$22253 ( \22630 , \22357 , \22629 );
xor \U$22254 ( \22631 , \21593 , \21604 );
xor \U$22255 ( \22632 , \22631 , \21617 );
xor \U$22256 ( \22633 , \21965 , \21972 );
xor \U$22257 ( \22634 , \22632 , \22633 );
and \U$22258 ( \22635 , \22630 , \22634 );
and \U$22259 ( \22636 , \22357 , \22629 );
or \U$22260 ( \22637 , \22635 , \22636 );
xor \U$22261 ( \22638 , \21977 , \22271 );
xor \U$22262 ( \22639 , \22638 , \22292 );
and \U$22263 ( \22640 , \22637 , \22639 );
xor \U$22264 ( \22641 , \21620 , \21856 );
xor \U$22265 ( \22642 , \22641 , \21871 );
xor \U$22266 ( \22643 , \22296 , \22303 );
xor \U$22267 ( \22644 , \22642 , \22643 );
xor \U$22268 ( \22645 , \21977 , \22271 );
xor \U$22269 ( \22646 , \22645 , \22292 );
and \U$22270 ( \22647 , \22644 , \22646 );
and \U$22271 ( \22648 , \22637 , \22644 );
or \U$22272 ( \22649 , \22640 , \22647 , \22648 );
xor \U$22273 ( \22650 , \21874 , \21879 );
xor \U$22274 ( \22651 , \22650 , \21906 );
and \U$22275 ( \22652 , \22649 , \22651 );
xor \U$22276 ( \22653 , \22295 , \22308 );
xor \U$22277 ( \22654 , \22653 , \22313 );
xor \U$22278 ( \22655 , \21874 , \21879 );
xor \U$22279 ( \22656 , \22655 , \21906 );
and \U$22280 ( \22657 , \22654 , \22656 );
and \U$22281 ( \22658 , \22649 , \22654 );
or \U$22282 ( \22659 , \22652 , \22657 , \22658 );
not \U$22283 ( \22660 , \22659 );
or \U$22284 ( \22661 , \22329 , \22660 );
xnor \U$22285 ( \22662 , \22660 , \22329 );
xor \U$22286 ( \22663 , \21874 , \21879 );
xor \U$22287 ( \22664 , \22663 , \21906 );
xor \U$22288 ( \22665 , \22649 , \22654 );
xor \U$22289 ( \22666 , \22664 , \22665 );
xor \U$22290 ( \22667 , \21977 , \22271 );
xor \U$22291 ( \22668 , \22667 , \22292 );
xor \U$22292 ( \22669 , \22637 , \22644 );
xor \U$22293 ( \22670 , \22668 , \22669 );
not \U$22294 ( \22671 , \22670 );
xor \U$22295 ( \22672 , \22197 , \22240 );
xor \U$22296 ( \22673 , \22672 , \22268 );
not \U$22297 ( \22674 , \22673 );
xor \U$22298 ( \22675 , \22357 , \22629 );
xor \U$22299 ( \22676 , \22675 , \22634 );
nand \U$22300 ( \22677 , \22674 , \22676 );
or \U$22301 ( \22678 , \22671 , \22677 );
not \U$22302 ( \22679 , \22677 );
not \U$22303 ( \22680 , \22671 );
or \U$22304 ( \22681 , \22679 , \22680 );
xor \U$22305 ( \22682 , \22502 , \22509 );
xor \U$22306 ( \22683 , \22682 , \22517 );
xor \U$22307 ( \22684 , \22483 , \1261 );
xor \U$22308 ( \22685 , \22684 , \22491 );
and \U$22309 ( \22686 , \22683 , \22685 );
xor \U$22310 ( \22687 , \22458 , \22465 );
xor \U$22311 ( \22688 , \22687 , \22473 );
xor \U$22312 ( \22689 , \22483 , \1261 );
xor \U$22313 ( \22690 , \22689 , \22491 );
and \U$22314 ( \22691 , \22688 , \22690 );
and \U$22315 ( \22692 , \22683 , \22688 );
or \U$22316 ( \22693 , \22686 , \22691 , \22692 );
xor \U$22317 ( \22694 , \22395 , \22402 );
xor \U$22318 ( \22695 , \22694 , \22410 );
nand \U$22319 ( \22696 , RIae775b8_79, \1374 );
and \U$22320 ( \22697 , \22696 , \1380 );
not \U$22321 ( \22698 , \22696 );
and \U$22322 ( \22699 , \22698 , \1261 );
nor \U$22323 ( \22700 , \22697 , \22699 );
xor \U$22324 ( \22701 , \22695 , \22700 );
xor \U$22325 ( \22702 , \22429 , \22437 );
xor \U$22326 ( \22703 , \22702 , \22445 );
and \U$22327 ( \22704 , \22701 , \22703 );
and \U$22328 ( \22705 , \22695 , \22700 );
or \U$22329 ( \22706 , \22704 , \22705 );
xor \U$22330 ( \22707 , \22693 , \22706 );
xor \U$22331 ( \22708 , \22582 , \22589 );
xor \U$22332 ( \22709 , \22708 , \22597 );
xor \U$22333 ( \22710 , \22556 , \22563 );
xor \U$22334 ( \22711 , \22710 , \22571 );
and \U$22335 ( \22712 , \22709 , \22711 );
xor \U$22336 ( \22713 , \22531 , \22538 );
xor \U$22337 ( \22714 , \22713 , \22546 );
xor \U$22338 ( \22715 , \22556 , \22563 );
xor \U$22339 ( \22716 , \22715 , \22571 );
and \U$22340 ( \22717 , \22714 , \22716 );
and \U$22341 ( \22718 , \22709 , \22714 );
or \U$22342 ( \22719 , \22712 , \22717 , \22718 );
and \U$22343 ( \22720 , \22707 , \22719 );
and \U$22344 ( \22721 , \22693 , \22706 );
or \U$22345 ( \22722 , \22720 , \22721 );
and \U$22346 ( \22723 , \13059 , RIae755d8_11);
and \U$22347 ( \22724 , RIae754e8_9, \13057 );
nor \U$22348 ( \22725 , \22723 , \22724 );
and \U$22349 ( \22726 , \22725 , \13063 );
not \U$22350 ( \22727 , \22725 );
and \U$22351 ( \22728 , \22727 , \12718 );
nor \U$22352 ( \22729 , \22726 , \22728 );
and \U$22353 ( \22730 , \11470 , RIae75f38_31);
and \U$22354 ( \22731 , RIae75e48_29, \11468 );
nor \U$22355 ( \22732 , \22730 , \22731 );
and \U$22356 ( \22733 , \22732 , \10936 );
not \U$22357 ( \22734 , \22732 );
and \U$22358 ( \22735 , \22734 , \11474 );
nor \U$22359 ( \22736 , \22733 , \22735 );
xor \U$22360 ( \22737 , \22729 , \22736 );
and \U$22361 ( \22738 , \12180 , RIae75c68_25);
and \U$22362 ( \22739 , RIae75d58_27, \12178 );
nor \U$22363 ( \22740 , \22738 , \22739 );
and \U$22364 ( \22741 , \22740 , \12184 );
not \U$22365 ( \22742 , \22740 );
and \U$22366 ( \22743 , \22742 , \11827 );
nor \U$22367 ( \22744 , \22741 , \22743 );
and \U$22368 ( \22745 , \22737 , \22744 );
and \U$22369 ( \22746 , \22729 , \22736 );
or \U$22370 ( \22747 , \22745 , \22746 );
and \U$22371 ( \22748 , \14059 , RIae757b8_15);
and \U$22372 ( \22749 , RIae756c8_13, \14057 );
nor \U$22373 ( \22750 , \22748 , \22749 );
and \U$22374 ( \22751 , \22750 , \13502 );
not \U$22375 ( \22752 , \22750 );
and \U$22376 ( \22753 , \22752 , \14063 );
nor \U$22377 ( \22754 , \22751 , \22753 );
and \U$22378 ( \22755 , \15726 , RIae75308_5);
and \U$22379 ( \22756 , RIae7aab0_192, RIae753f8_7);
nor \U$22380 ( \22757 , \22755 , \22756 );
and \U$22381 ( \22758 , \22757 , \14959 );
not \U$22382 ( \22759 , \22757 );
and \U$22383 ( \22760 , \22759 , RIae7aa38_191);
nor \U$22384 ( \22761 , \22758 , \22760 );
xor \U$22385 ( \22762 , \22754 , \22761 );
and \U$22386 ( \22763 , \14964 , RIae75218_3);
and \U$22387 ( \22764 , RIae75128_1, \14962 );
nor \U$22388 ( \22765 , \22763 , \22764 );
and \U$22389 ( \22766 , \22765 , \14463 );
not \U$22390 ( \22767 , \22765 );
and \U$22391 ( \22768 , \22767 , \14462 );
nor \U$22392 ( \22769 , \22766 , \22768 );
and \U$22393 ( \22770 , \22762 , \22769 );
and \U$22394 ( \22771 , \22754 , \22761 );
or \U$22395 ( \22772 , \22770 , \22771 );
xor \U$22396 ( \22773 , \22747 , \22772 );
and \U$22397 ( \22774 , \8966 , RIae78788_117);
and \U$22398 ( \22775 , RIae78698_115, \8964 );
nor \U$22399 ( \22776 , \22774 , \22775 );
and \U$22400 ( \22777 , \22776 , \8799 );
not \U$22401 ( \22778 , \22776 );
and \U$22402 ( \22779 , \22778 , \8789 );
nor \U$22403 ( \22780 , \22777 , \22779 );
and \U$22404 ( \22781 , \9760 , RIae75b78_23);
and \U$22405 ( \22782 , RIae75a88_21, \9758 );
nor \U$22406 ( \22783 , \22781 , \22782 );
and \U$22407 ( \22784 , \22783 , \9273 );
not \U$22408 ( \22785 , \22783 );
and \U$22409 ( \22786 , \22785 , \9272 );
nor \U$22410 ( \22787 , \22784 , \22786 );
xor \U$22411 ( \22788 , \22780 , \22787 );
and \U$22412 ( \22789 , \10548 , RIae75998_19);
and \U$22413 ( \22790 , RIae758a8_17, \10546 );
nor \U$22414 ( \22791 , \22789 , \22790 );
and \U$22415 ( \22792 , \22791 , \10421 );
not \U$22416 ( \22793 , \22791 );
and \U$22417 ( \22794 , \22793 , \10118 );
nor \U$22418 ( \22795 , \22792 , \22794 );
and \U$22419 ( \22796 , \22788 , \22795 );
and \U$22420 ( \22797 , \22780 , \22787 );
or \U$22421 ( \22798 , \22796 , \22797 );
and \U$22422 ( \22799 , \22773 , \22798 );
and \U$22423 ( \22800 , \22747 , \22772 );
or \U$22424 ( \22801 , \22799 , \22800 );
and \U$22425 ( \22802 , \2607 , RIae77798_83);
and \U$22426 ( \22803 , RIae77888_85, \2605 );
nor \U$22427 ( \22804 , \22802 , \22803 );
and \U$22428 ( \22805 , \22804 , \2611 );
not \U$22429 ( \22806 , \22804 );
and \U$22430 ( \22807 , \22806 , \2397 );
nor \U$22431 ( \22808 , \22805 , \22807 );
not \U$22432 ( \22809 , \2789 );
and \U$22433 ( \22810 , \2783 , RIae76f28_65);
and \U$22434 ( \22811 , RIae76e38_63, \2781 );
nor \U$22435 ( \22812 , \22810 , \22811 );
not \U$22436 ( \22813 , \22812 );
or \U$22437 ( \22814 , \22809 , \22813 );
or \U$22438 ( \22815 , \22812 , \3089 );
nand \U$22439 ( \22816 , \22814 , \22815 );
xor \U$22440 ( \22817 , \22808 , \22816 );
not \U$22441 ( \22818 , \3218 );
and \U$22442 ( \22819 , \3214 , RIae76d48_61);
and \U$22443 ( \22820 , RIae76c58_59, \3212 );
nor \U$22444 ( \22821 , \22819 , \22820 );
not \U$22445 ( \22822 , \22821 );
or \U$22446 ( \22823 , \22818 , \22822 );
or \U$22447 ( \22824 , \22821 , \2774 );
nand \U$22448 ( \22825 , \22823 , \22824 );
and \U$22449 ( \22826 , \22817 , \22825 );
and \U$22450 ( \22827 , \22808 , \22816 );
or \U$22451 ( \22828 , \22826 , \22827 );
and \U$22452 ( \22829 , \1593 , RIae774c8_77);
and \U$22453 ( \22830 , RIae77720_82, \1591 );
nor \U$22454 ( \22831 , \22829 , \22830 );
and \U$22455 ( \22832 , \22831 , \1498 );
not \U$22456 ( \22833 , \22831 );
and \U$22457 ( \22834 , \22833 , \1488 );
nor \U$22458 ( \22835 , \22832 , \22834 );
xor \U$22459 ( \22836 , \22828 , \22835 );
and \U$22460 ( \22837 , \2224 , RIae77a68_89);
and \U$22461 ( \22838 , RIae77978_87, \2222 );
nor \U$22462 ( \22839 , \22837 , \22838 );
and \U$22463 ( \22840 , \22839 , \2061 );
not \U$22464 ( \22841 , \22839 );
and \U$22465 ( \22842 , \22841 , \2060 );
nor \U$22466 ( \22843 , \22840 , \22842 );
and \U$22467 ( \22844 , \1593 , RIae775b8_79);
and \U$22468 ( \22845 , RIae774c8_77, \1591 );
nor \U$22469 ( \22846 , \22844 , \22845 );
and \U$22470 ( \22847 , \22846 , \1498 );
not \U$22471 ( \22848 , \22846 );
and \U$22472 ( \22849 , \22848 , \1488 );
nor \U$22473 ( \22850 , \22847 , \22849 );
xor \U$22474 ( \22851 , \22843 , \22850 );
and \U$22475 ( \22852 , \1939 , RIae77720_82);
and \U$22476 ( \22853 , RIae773d8_75, \1937 );
nor \U$22477 ( \22854 , \22852 , \22853 );
and \U$22478 ( \22855 , \22854 , \1735 );
not \U$22479 ( \22856 , \22854 );
and \U$22480 ( \22857 , \22856 , \1734 );
nor \U$22481 ( \22858 , \22855 , \22857 );
and \U$22482 ( \22859 , \22851 , \22858 );
and \U$22483 ( \22860 , \22843 , \22850 );
or \U$22484 ( \22861 , \22859 , \22860 );
and \U$22485 ( \22862 , \22836 , \22861 );
and \U$22486 ( \22863 , \22828 , \22835 );
or \U$22487 ( \22864 , \22862 , \22863 );
xor \U$22488 ( \22865 , \22801 , \22864 );
and \U$22489 ( \22866 , \6941 , RIae77c48_93);
and \U$22490 ( \22867 , RIae77b58_91, \6939 );
nor \U$22491 ( \22868 , \22866 , \22867 );
and \U$22492 ( \22869 , \22868 , \6314 );
not \U$22493 ( \22870 , \22868 );
and \U$22494 ( \22871 , \22870 , \6945 );
nor \U$22495 ( \22872 , \22869 , \22871 );
and \U$22496 ( \22873 , \7633 , RIae77d38_95);
and \U$22497 ( \22874 , RIae77e28_97, \7631 );
nor \U$22498 ( \22875 , \22873 , \22874 );
and \U$22499 ( \22876 , \22875 , \7206 );
not \U$22500 ( \22877 , \22875 );
and \U$22501 ( \22878 , \22877 , \7205 );
nor \U$22502 ( \22879 , \22876 , \22878 );
xor \U$22503 ( \22880 , \22872 , \22879 );
and \U$22504 ( \22881 , \8371 , RIae78968_121);
and \U$22505 ( \22882 , RIae78878_119, \8369 );
nor \U$22506 ( \22883 , \22881 , \22882 );
and \U$22507 ( \22884 , \22883 , \8020 );
not \U$22508 ( \22885 , \22883 );
and \U$22509 ( \22886 , \22885 , \8019 );
nor \U$22510 ( \22887 , \22884 , \22886 );
and \U$22511 ( \22888 , \22880 , \22887 );
and \U$22512 ( \22889 , \22872 , \22879 );
or \U$22513 ( \22890 , \22888 , \22889 );
and \U$22514 ( \22891 , \3730 , RIae77180_70);
and \U$22515 ( \22892 , RIae77018_67, \3728 );
nor \U$22516 ( \22893 , \22891 , \22892 );
and \U$22517 ( \22894 , \22893 , \3732 );
not \U$22518 ( \22895 , \22893 );
and \U$22519 ( \22896 , \22895 , \3422 );
nor \U$22520 ( \22897 , \22894 , \22896 );
and \U$22521 ( \22898 , \4247 , RIae771f8_71);
and \U$22522 ( \22899 , RIae772e8_73, \4245 );
nor \U$22523 ( \22900 , \22898 , \22899 );
and \U$22524 ( \22901 , \22900 , \3989 );
not \U$22525 ( \22902 , \22900 );
and \U$22526 ( \22903 , \22902 , \4251 );
nor \U$22527 ( \22904 , \22901 , \22903 );
xor \U$22528 ( \22905 , \22897 , \22904 );
and \U$22529 ( \22906 , \4688 , RIae782d8_107);
and \U$22530 ( \22907 , RIae780f8_103, \4686 );
nor \U$22531 ( \22908 , \22906 , \22907 );
and \U$22532 ( \22909 , \22908 , \4481 );
not \U$22533 ( \22910 , \22908 );
and \U$22534 ( \22911 , \22910 , \4482 );
nor \U$22535 ( \22912 , \22909 , \22911 );
and \U$22536 ( \22913 , \22905 , \22912 );
and \U$22537 ( \22914 , \22897 , \22904 );
or \U$22538 ( \22915 , \22913 , \22914 );
xor \U$22539 ( \22916 , \22890 , \22915 );
and \U$22540 ( \22917 , \5896 , RIae781e8_105);
and \U$22541 ( \22918 , RIae785a8_113, \5894 );
nor \U$22542 ( \22919 , \22917 , \22918 );
and \U$22543 ( \22920 , \22919 , \5590 );
not \U$22544 ( \22921 , \22919 );
and \U$22545 ( \22922 , \22921 , \5589 );
nor \U$22546 ( \22923 , \22920 , \22922 );
and \U$22547 ( \22924 , \5399 , RIae77f18_99);
and \U$22548 ( \22925 , RIae78008_101, \5397 );
nor \U$22549 ( \22926 , \22924 , \22925 );
and \U$22550 ( \22927 , \22926 , \5016 );
not \U$22551 ( \22928 , \22926 );
and \U$22552 ( \22929 , \22928 , \5403 );
nor \U$22553 ( \22930 , \22927 , \22929 );
xor \U$22554 ( \22931 , \22923 , \22930 );
and \U$22555 ( \22932 , \6172 , RIae783c8_109);
and \U$22556 ( \22933 , RIae78530_112, \6170 );
nor \U$22557 ( \22934 , \22932 , \22933 );
and \U$22558 ( \22935 , \22934 , \6176 );
not \U$22559 ( \22936 , \22934 );
and \U$22560 ( \22937 , \22936 , \6175 );
nor \U$22561 ( \22938 , \22935 , \22937 );
and \U$22562 ( \22939 , \22931 , \22938 );
and \U$22563 ( \22940 , \22923 , \22930 );
or \U$22564 ( \22941 , \22939 , \22940 );
and \U$22565 ( \22942 , \22916 , \22941 );
and \U$22566 ( \22943 , \22890 , \22915 );
or \U$22567 ( \22944 , \22942 , \22943 );
and \U$22568 ( \22945 , \22865 , \22944 );
and \U$22569 ( \22946 , \22801 , \22864 );
or \U$22570 ( \22947 , \22945 , \22946 );
xor \U$22571 ( \22948 , \22722 , \22947 );
xor \U$22572 ( \22949 , \22369 , \22371 );
xor \U$22573 ( \22950 , \22359 , \22361 );
xor \U$22574 ( \22951 , \22950 , \22364 );
and \U$22575 ( \22952 , \22949 , \22951 );
xor \U$22576 ( \22953 , \22173 , \22180 );
xor \U$22577 ( \22954 , \22953 , \22188 );
xor \U$22578 ( \22955 , \22375 , \22380 );
xor \U$22579 ( \22956 , \22954 , \22955 );
xor \U$22580 ( \22957 , \22359 , \22361 );
xor \U$22581 ( \22958 , \22957 , \22364 );
and \U$22582 ( \22959 , \22956 , \22958 );
and \U$22583 ( \22960 , \22949 , \22956 );
or \U$22584 ( \22961 , \22952 , \22959 , \22960 );
and \U$22585 ( \22962 , \22948 , \22961 );
and \U$22586 ( \22963 , \22722 , \22947 );
nor \U$22587 ( \22964 , \22962 , \22963 );
xor \U$22588 ( \22965 , \22210 , \22216 );
xor \U$22589 ( \22966 , \22965 , \22237 );
or \U$22590 ( \22967 , \22964 , \22966 );
not \U$22591 ( \22968 , \22966 );
not \U$22592 ( \22969 , \22964 );
or \U$22593 ( \22970 , \22968 , \22969 );
xor \U$22594 ( \22971 , \22413 , \22420 );
xor \U$22595 ( \22972 , \22971 , \22448 );
xor \U$22596 ( \22973 , \22549 , \22574 );
xor \U$22597 ( \22974 , \22973 , \22600 );
and \U$22598 ( \22975 , \22972 , \22974 );
xor \U$22599 ( \22976 , \22476 , \22494 );
xor \U$22600 ( \22977 , \22976 , \22520 );
xor \U$22601 ( \22978 , \22549 , \22574 );
xor \U$22602 ( \22979 , \22978 , \22600 );
and \U$22603 ( \22980 , \22977 , \22979 );
and \U$22604 ( \22981 , \22972 , \22977 );
or \U$22605 ( \22982 , \22975 , \22980 , \22981 );
xor \U$22606 ( \22983 , \22331 , \22333 );
xor \U$22607 ( \22984 , \22983 , \22336 );
and \U$22608 ( \22985 , \22982 , \22984 );
xor \U$22609 ( \22986 , \22613 , \22618 );
xor \U$22610 ( \22987 , \22986 , \22623 );
xor \U$22611 ( \22988 , \22331 , \22333 );
xor \U$22612 ( \22989 , \22988 , \22336 );
and \U$22613 ( \22990 , \22987 , \22989 );
and \U$22614 ( \22991 , \22982 , \22987 );
or \U$22615 ( \22992 , \22985 , \22990 , \22991 );
nand \U$22616 ( \22993 , \22970 , \22992 );
nand \U$22617 ( \22994 , \22967 , \22993 );
xor \U$22618 ( \22995 , \22282 , \22284 );
xor \U$22619 ( \22996 , \22995 , \22289 );
xor \U$22620 ( \22997 , \22994 , \22996 );
xor \U$22621 ( \22998 , \22035 , \22114 );
xor \U$22622 ( \22999 , \22998 , \22194 );
xor \U$22623 ( \23000 , \22388 , \22606 );
xor \U$22624 ( \23001 , \23000 , \22626 );
and \U$22625 ( \23002 , \22999 , \23001 );
xor \U$22626 ( \23003 , \22274 , \22276 );
xor \U$22627 ( \23004 , \23003 , \22279 );
xor \U$22628 ( \23005 , \22339 , \22352 );
xor \U$22629 ( \23006 , \23004 , \23005 );
xor \U$22630 ( \23007 , \22388 , \22606 );
xor \U$22631 ( \23008 , \23007 , \22626 );
and \U$22632 ( \23009 , \23006 , \23008 );
and \U$22633 ( \23010 , \22999 , \23006 );
or \U$22634 ( \23011 , \23002 , \23009 , \23010 );
and \U$22635 ( \23012 , \22997 , \23011 );
and \U$22636 ( \23013 , \22994 , \22996 );
or \U$22637 ( \23014 , \23012 , \23013 );
nand \U$22638 ( \23015 , \22681 , \23014 );
nand \U$22639 ( \23016 , \22678 , \23015 );
and \U$22640 ( \23017 , \22666 , \23016 );
xor \U$22641 ( \23018 , \23016 , \22666 );
not \U$22642 ( \23019 , \23014 );
not \U$22643 ( \23020 , \22677 );
and \U$22644 ( \23021 , \23019 , \23020 );
and \U$22645 ( \23022 , \23014 , \22677 );
nor \U$22646 ( \23023 , \23021 , \23022 );
not \U$22647 ( \23024 , \23023 );
not \U$22648 ( \23025 , \22670 );
and \U$22649 ( \23026 , \23024 , \23025 );
and \U$22650 ( \23027 , \23023 , \22670 );
nor \U$22651 ( \23028 , \23026 , \23027 );
not \U$22652 ( \23029 , \22673 );
not \U$22653 ( \23030 , \22676 );
or \U$22654 ( \23031 , \23029 , \23030 );
or \U$22655 ( \23032 , \22676 , \22673 );
nand \U$22656 ( \23033 , \23031 , \23032 );
xor \U$22657 ( \23034 , \22994 , \22996 );
xor \U$22658 ( \23035 , \23034 , \23011 );
xor \U$22659 ( \23036 , \23033 , \23035 );
xor \U$22660 ( \23037 , \22722 , \22947 );
xor \U$22661 ( \23038 , \23037 , \22961 );
xor \U$22662 ( \23039 , \22451 , \22523 );
xor \U$22663 ( \23040 , \23039 , \22603 );
xor \U$22664 ( \23041 , \23038 , \23040 );
xor \U$22665 ( \23042 , \22331 , \22333 );
xor \U$22666 ( \23043 , \23042 , \22336 );
xor \U$22667 ( \23044 , \22982 , \22987 );
xor \U$22668 ( \23045 , \23043 , \23044 );
and \U$22669 ( \23046 , \23041 , \23045 );
and \U$22670 ( \23047 , \23038 , \23040 );
or \U$22671 ( \23048 , \23046 , \23047 );
not \U$22672 ( \23049 , \23048 );
xor \U$22673 ( \23050 , \22388 , \22606 );
xor \U$22674 ( \23051 , \23050 , \22626 );
xor \U$22675 ( \23052 , \22999 , \23006 );
xor \U$22676 ( \23053 , \23051 , \23052 );
not \U$22677 ( \23054 , \23053 );
or \U$22678 ( \23055 , \23049 , \23054 );
or \U$22679 ( \23056 , \23053 , \23048 );
xor \U$22680 ( \23057 , \22897 , \22904 );
xor \U$22681 ( \23058 , \23057 , \22912 );
xor \U$22682 ( \23059 , \22808 , \22816 );
xor \U$22683 ( \23060 , \23059 , \22825 );
and \U$22684 ( \23061 , \23058 , \23060 );
xor \U$22685 ( \23062 , \22923 , \22930 );
xor \U$22686 ( \23063 , \23062 , \22938 );
xor \U$22687 ( \23064 , \22808 , \22816 );
xor \U$22688 ( \23065 , \23064 , \22825 );
and \U$22689 ( \23066 , \23063 , \23065 );
and \U$22690 ( \23067 , \23058 , \23063 );
or \U$22691 ( \23068 , \23061 , \23066 , \23067 );
xor \U$22692 ( \23069 , \22780 , \22787 );
xor \U$22693 ( \23070 , \23069 , \22795 );
xor \U$22694 ( \23071 , \22872 , \22879 );
xor \U$22695 ( \23072 , \23071 , \22887 );
xor \U$22696 ( \23073 , \23070 , \23072 );
xor \U$22697 ( \23074 , \22729 , \22736 );
xor \U$22698 ( \23075 , \23074 , \22744 );
and \U$22699 ( \23076 , \23073 , \23075 );
and \U$22700 ( \23077 , \23070 , \23072 );
or \U$22701 ( \23078 , \23076 , \23077 );
xor \U$22702 ( \23079 , \23068 , \23078 );
xor \U$22703 ( \23080 , \22483 , \1261 );
xor \U$22704 ( \23081 , \23080 , \22491 );
xor \U$22705 ( \23082 , \22683 , \22688 );
xor \U$22706 ( \23083 , \23081 , \23082 );
and \U$22707 ( \23084 , \23079 , \23083 );
and \U$22708 ( \23085 , \23068 , \23078 );
or \U$22709 ( \23086 , \23084 , \23085 );
not \U$22710 ( \23087 , \3089 );
and \U$22711 ( \23088 , \2783 , RIae77888_85);
and \U$22712 ( \23089 , RIae76f28_65, \2781 );
nor \U$22713 ( \23090 , \23088 , \23089 );
not \U$22714 ( \23091 , \23090 );
or \U$22715 ( \23092 , \23087 , \23091 );
or \U$22716 ( \23093 , \23090 , \2789 );
nand \U$22717 ( \23094 , \23092 , \23093 );
not \U$22718 ( \23095 , \3218 );
and \U$22719 ( \23096 , \3214 , RIae76e38_63);
and \U$22720 ( \23097 , RIae76d48_61, \3212 );
nor \U$22721 ( \23098 , \23096 , \23097 );
not \U$22722 ( \23099 , \23098 );
or \U$22723 ( \23100 , \23095 , \23099 );
or \U$22724 ( \23101 , \23098 , \3218 );
nand \U$22725 ( \23102 , \23100 , \23101 );
xor \U$22726 ( \23103 , \23094 , \23102 );
and \U$22727 ( \23104 , \3730 , RIae76c58_59);
and \U$22728 ( \23105 , RIae77180_70, \3728 );
nor \U$22729 ( \23106 , \23104 , \23105 );
and \U$22730 ( \23107 , \23106 , \3732 );
not \U$22731 ( \23108 , \23106 );
and \U$22732 ( \23109 , \23108 , \3422 );
nor \U$22733 ( \23110 , \23107 , \23109 );
and \U$22734 ( \23111 , \23103 , \23110 );
and \U$22735 ( \23112 , \23094 , \23102 );
or \U$22736 ( \23113 , \23111 , \23112 );
and \U$22737 ( \23114 , \1939 , RIae774c8_77);
and \U$22738 ( \23115 , RIae77720_82, \1937 );
nor \U$22739 ( \23116 , \23114 , \23115 );
and \U$22740 ( \23117 , \23116 , \1735 );
not \U$22741 ( \23118 , \23116 );
and \U$22742 ( \23119 , \23118 , \1734 );
nor \U$22743 ( \23120 , \23117 , \23119 );
and \U$22744 ( \23121 , \2224 , RIae773d8_75);
and \U$22745 ( \23122 , RIae77a68_89, \2222 );
nor \U$22746 ( \23123 , \23121 , \23122 );
and \U$22747 ( \23124 , \23123 , \2061 );
not \U$22748 ( \23125 , \23123 );
and \U$22749 ( \23126 , \23125 , \2060 );
nor \U$22750 ( \23127 , \23124 , \23126 );
xor \U$22751 ( \23128 , \23120 , \23127 );
and \U$22752 ( \23129 , \2607 , RIae77978_87);
and \U$22753 ( \23130 , RIae77798_83, \2605 );
nor \U$22754 ( \23131 , \23129 , \23130 );
and \U$22755 ( \23132 , \23131 , \2611 );
not \U$22756 ( \23133 , \23131 );
and \U$22757 ( \23134 , \23133 , \2397 );
nor \U$22758 ( \23135 , \23132 , \23134 );
and \U$22759 ( \23136 , \23128 , \23135 );
and \U$22760 ( \23137 , \23120 , \23127 );
or \U$22761 ( \23138 , \23136 , \23137 );
xor \U$22762 ( \23139 , \23113 , \23138 );
xor \U$22763 ( \23140 , \22843 , \22850 );
xor \U$22764 ( \23141 , \23140 , \22858 );
and \U$22765 ( \23142 , \23139 , \23141 );
and \U$22766 ( \23143 , \23113 , \23138 );
nor \U$22767 ( \23144 , \23142 , \23143 );
and \U$22768 ( \23145 , \4247 , RIae77018_67);
and \U$22769 ( \23146 , RIae771f8_71, \4245 );
nor \U$22770 ( \23147 , \23145 , \23146 );
and \U$22771 ( \23148 , \23147 , \4251 );
not \U$22772 ( \23149 , \23147 );
and \U$22773 ( \23150 , \23149 , \3989 );
nor \U$22774 ( \23151 , \23148 , \23150 );
not \U$22775 ( \23152 , \23151 );
and \U$22776 ( \23153 , \4688 , RIae772e8_73);
and \U$22777 ( \23154 , RIae782d8_107, \4686 );
nor \U$22778 ( \23155 , \23153 , \23154 );
and \U$22779 ( \23156 , \23155 , \4482 );
not \U$22780 ( \23157 , \23155 );
and \U$22781 ( \23158 , \23157 , \4481 );
nor \U$22782 ( \23159 , \23156 , \23158 );
not \U$22783 ( \23160 , \23159 );
and \U$22784 ( \23161 , \23152 , \23160 );
and \U$22785 ( \23162 , \23159 , \23151 );
and \U$22786 ( \23163 , \5399 , RIae780f8_103);
and \U$22787 ( \23164 , RIae77f18_99, \5397 );
nor \U$22788 ( \23165 , \23163 , \23164 );
and \U$22789 ( \23166 , \23165 , \5403 );
not \U$22790 ( \23167 , \23165 );
and \U$22791 ( \23168 , \23167 , \5016 );
nor \U$22792 ( \23169 , \23166 , \23168 );
nor \U$22793 ( \23170 , \23162 , \23169 );
nor \U$22794 ( \23171 , \23161 , \23170 );
not \U$22795 ( \23172 , \23171 );
and \U$22796 ( \23173 , \7633 , RIae77b58_91);
and \U$22797 ( \23174 , RIae77d38_95, \7631 );
nor \U$22798 ( \23175 , \23173 , \23174 );
and \U$22799 ( \23176 , \23175 , \7205 );
not \U$22800 ( \23177 , \23175 );
and \U$22801 ( \23178 , \23177 , \7206 );
nor \U$22802 ( \23179 , \23176 , \23178 );
not \U$22803 ( \23180 , \23179 );
and \U$22804 ( \23181 , \8966 , RIae78878_119);
and \U$22805 ( \23182 , RIae78788_117, \8964 );
nor \U$22806 ( \23183 , \23181 , \23182 );
and \U$22807 ( \23184 , \23183 , \8789 );
not \U$22808 ( \23185 , \23183 );
and \U$22809 ( \23186 , \23185 , \8799 );
nor \U$22810 ( \23187 , \23184 , \23186 );
not \U$22811 ( \23188 , \23187 );
and \U$22812 ( \23189 , \23180 , \23188 );
and \U$22813 ( \23190 , \23187 , \23179 );
and \U$22814 ( \23191 , \8371 , RIae77e28_97);
and \U$22815 ( \23192 , RIae78968_121, \8369 );
nor \U$22816 ( \23193 , \23191 , \23192 );
and \U$22817 ( \23194 , \23193 , \8019 );
not \U$22818 ( \23195 , \23193 );
and \U$22819 ( \23196 , \23195 , \8020 );
nor \U$22820 ( \23197 , \23194 , \23196 );
nor \U$22821 ( \23198 , \23190 , \23197 );
nor \U$22822 ( \23199 , \23189 , \23198 );
not \U$22823 ( \23200 , \23199 );
and \U$22824 ( \23201 , \23172 , \23200 );
and \U$22825 ( \23202 , \23171 , \23199 );
and \U$22826 ( \23203 , \5896 , RIae78008_101);
and \U$22827 ( \23204 , RIae781e8_105, \5894 );
nor \U$22828 ( \23205 , \23203 , \23204 );
and \U$22829 ( \23206 , \23205 , \5590 );
not \U$22830 ( \23207 , \23205 );
and \U$22831 ( \23208 , \23207 , \5589 );
nor \U$22832 ( \23209 , \23206 , \23208 );
and \U$22833 ( \23210 , \6172 , RIae785a8_113);
and \U$22834 ( \23211 , RIae783c8_109, \6170 );
nor \U$22835 ( \23212 , \23210 , \23211 );
and \U$22836 ( \23213 , \23212 , \6176 );
not \U$22837 ( \23214 , \23212 );
and \U$22838 ( \23215 , \23214 , \6175 );
nor \U$22839 ( \23216 , \23213 , \23215 );
xor \U$22840 ( \23217 , \23209 , \23216 );
and \U$22841 ( \23218 , \6941 , RIae78530_112);
and \U$22842 ( \23219 , RIae77c48_93, \6939 );
nor \U$22843 ( \23220 , \23218 , \23219 );
and \U$22844 ( \23221 , \23220 , \6314 );
not \U$22845 ( \23222 , \23220 );
and \U$22846 ( \23223 , \23222 , \6945 );
nor \U$22847 ( \23224 , \23221 , \23223 );
and \U$22848 ( \23225 , \23217 , \23224 );
and \U$22849 ( \23226 , \23209 , \23216 );
or \U$22850 ( \23227 , \23225 , \23226 );
not \U$22851 ( \23228 , \23227 );
nor \U$22852 ( \23229 , \23202 , \23228 );
nor \U$22853 ( \23230 , \23201 , \23229 );
or \U$22854 ( \23231 , \23144 , \23230 );
not \U$22855 ( \23232 , \23230 );
not \U$22856 ( \23233 , \23144 );
or \U$22857 ( \23234 , \23232 , \23233 );
and \U$22858 ( \23235 , \12180 , RIae75e48_29);
and \U$22859 ( \23236 , RIae75c68_25, \12178 );
nor \U$22860 ( \23237 , \23235 , \23236 );
and \U$22861 ( \23238 , \23237 , \12184 );
not \U$22862 ( \23239 , \23237 );
and \U$22863 ( \23240 , \23239 , \11827 );
nor \U$22864 ( \23241 , \23238 , \23240 );
and \U$22865 ( \23242 , \13059 , RIae75d58_27);
and \U$22866 ( \23243 , RIae755d8_11, \13057 );
nor \U$22867 ( \23244 , \23242 , \23243 );
and \U$22868 ( \23245 , \23244 , \13063 );
not \U$22869 ( \23246 , \23244 );
and \U$22870 ( \23247 , \23246 , \12718 );
nor \U$22871 ( \23248 , \23245 , \23247 );
xor \U$22872 ( \23249 , \23241 , \23248 );
and \U$22873 ( \23250 , \14059 , RIae754e8_9);
and \U$22874 ( \23251 , RIae757b8_15, \14057 );
nor \U$22875 ( \23252 , \23250 , \23251 );
and \U$22876 ( \23253 , \23252 , \13502 );
not \U$22877 ( \23254 , \23252 );
and \U$22878 ( \23255 , \23254 , \14063 );
nor \U$22879 ( \23256 , \23253 , \23255 );
and \U$22880 ( \23257 , \23249 , \23256 );
and \U$22881 ( \23258 , \23241 , \23248 );
or \U$22882 ( \23259 , \23257 , \23258 );
and \U$22883 ( \23260 , \15726 , RIae75128_1);
and \U$22884 ( \23261 , RIae7aab0_192, RIae75308_5);
nor \U$22885 ( \23262 , \23260 , \23261 );
and \U$22886 ( \23263 , \23262 , \14959 );
not \U$22887 ( \23264 , \23262 );
and \U$22888 ( \23265 , \23264 , RIae7aa38_191);
nor \U$22889 ( \23266 , \23263 , \23265 );
xor \U$22890 ( \23267 , \23266 , \1488 );
and \U$22891 ( \23268 , \14964 , RIae756c8_13);
and \U$22892 ( \23269 , RIae75218_3, \14962 );
nor \U$22893 ( \23270 , \23268 , \23269 );
and \U$22894 ( \23271 , \23270 , \14463 );
not \U$22895 ( \23272 , \23270 );
and \U$22896 ( \23273 , \23272 , \14462 );
nor \U$22897 ( \23274 , \23271 , \23273 );
and \U$22898 ( \23275 , \23267 , \23274 );
and \U$22899 ( \23276 , \23266 , \1488 );
or \U$22900 ( \23277 , \23275 , \23276 );
xor \U$22901 ( \23278 , \23259 , \23277 );
and \U$22902 ( \23279 , \9760 , RIae78698_115);
and \U$22903 ( \23280 , RIae75b78_23, \9758 );
nor \U$22904 ( \23281 , \23279 , \23280 );
and \U$22905 ( \23282 , \23281 , \9273 );
not \U$22906 ( \23283 , \23281 );
and \U$22907 ( \23284 , \23283 , \9764 );
nor \U$22908 ( \23285 , \23282 , \23284 );
and \U$22909 ( \23286 , \10548 , RIae75a88_21);
and \U$22910 ( \23287 , RIae75998_19, \10546 );
nor \U$22911 ( \23288 , \23286 , \23287 );
and \U$22912 ( \23289 , \23288 , \10421 );
not \U$22913 ( \23290 , \23288 );
and \U$22914 ( \23291 , \23290 , \10118 );
nor \U$22915 ( \23292 , \23289 , \23291 );
xor \U$22916 ( \23293 , \23285 , \23292 );
and \U$22917 ( \23294 , \11470 , RIae758a8_17);
and \U$22918 ( \23295 , RIae75f38_31, \11468 );
nor \U$22919 ( \23296 , \23294 , \23295 );
and \U$22920 ( \23297 , \23296 , \10936 );
not \U$22921 ( \23298 , \23296 );
and \U$22922 ( \23299 , \23298 , \11474 );
nor \U$22923 ( \23300 , \23297 , \23299 );
and \U$22924 ( \23301 , \23293 , \23300 );
and \U$22925 ( \23302 , \23285 , \23292 );
or \U$22926 ( \23303 , \23301 , \23302 );
and \U$22927 ( \23304 , \23278 , \23303 );
and \U$22928 ( \23305 , \23259 , \23277 );
or \U$22929 ( \23306 , \23304 , \23305 );
nand \U$22930 ( \23307 , \23234 , \23306 );
nand \U$22931 ( \23308 , \23231 , \23307 );
xor \U$22932 ( \23309 , \23086 , \23308 );
xor \U$22933 ( \23310 , \22828 , \22835 );
xor \U$22934 ( \23311 , \23310 , \22861 );
xor \U$22935 ( \23312 , \22695 , \22700 );
xor \U$22936 ( \23313 , \23312 , \22703 );
and \U$22937 ( \23314 , \23311 , \23313 );
xor \U$22938 ( \23315 , \22556 , \22563 );
xor \U$22939 ( \23316 , \23315 , \22571 );
xor \U$22940 ( \23317 , \22709 , \22714 );
xor \U$22941 ( \23318 , \23316 , \23317 );
xor \U$22942 ( \23319 , \22695 , \22700 );
xor \U$22943 ( \23320 , \23319 , \22703 );
and \U$22944 ( \23321 , \23318 , \23320 );
and \U$22945 ( \23322 , \23311 , \23318 );
or \U$22946 ( \23323 , \23314 , \23321 , \23322 );
and \U$22947 ( \23324 , \23309 , \23323 );
and \U$22948 ( \23325 , \23086 , \23308 );
or \U$22949 ( \23326 , \23324 , \23325 );
xor \U$22950 ( \23327 , \22367 , \22372 );
xor \U$22951 ( \23328 , \23327 , \22385 );
xor \U$22952 ( \23329 , \23326 , \23328 );
xor \U$22953 ( \23330 , \22549 , \22574 );
xor \U$22954 ( \23331 , \23330 , \22600 );
xor \U$22955 ( \23332 , \22972 , \22977 );
xor \U$22956 ( \23333 , \23331 , \23332 );
xor \U$22957 ( \23334 , \22693 , \22706 );
xor \U$22958 ( \23335 , \23334 , \22719 );
and \U$22959 ( \23336 , \23333 , \23335 );
xor \U$22960 ( \23337 , \22359 , \22361 );
xor \U$22961 ( \23338 , \23337 , \22364 );
xor \U$22962 ( \23339 , \22949 , \22956 );
xor \U$22963 ( \23340 , \23338 , \23339 );
xor \U$22964 ( \23341 , \22693 , \22706 );
xor \U$22965 ( \23342 , \23341 , \22719 );
and \U$22966 ( \23343 , \23340 , \23342 );
and \U$22967 ( \23344 , \23333 , \23340 );
or \U$22968 ( \23345 , \23336 , \23343 , \23344 );
and \U$22969 ( \23346 , \23329 , \23345 );
and \U$22970 ( \23347 , \23326 , \23328 );
or \U$22971 ( \23348 , \23346 , \23347 );
nand \U$22972 ( \23349 , \23056 , \23348 );
nand \U$22973 ( \23350 , \23055 , \23349 );
and \U$22974 ( \23351 , \23036 , \23350 );
and \U$22975 ( \23352 , \23033 , \23035 );
nor \U$22976 ( \23353 , \23351 , \23352 );
or \U$22977 ( \23354 , \23028 , \23353 );
xnor \U$22978 ( \23355 , \23028 , \23353 );
not \U$22979 ( \23356 , \22964 );
not \U$22980 ( \23357 , \22992 );
or \U$22981 ( \23358 , \23356 , \23357 );
or \U$22982 ( \23359 , \22992 , \22964 );
nand \U$22983 ( \23360 , \23358 , \23359 );
not \U$22984 ( \23361 , \23360 );
not \U$22985 ( \23362 , \22966 );
and \U$22986 ( \23363 , \23361 , \23362 );
and \U$22987 ( \23364 , \23360 , \22966 );
nor \U$22988 ( \23365 , \23363 , \23364 );
not \U$22989 ( \23366 , \23365 );
xor \U$22990 ( \23367 , \22801 , \22864 );
xor \U$22991 ( \23368 , \23367 , \22944 );
xor \U$22992 ( \23369 , \23086 , \23308 );
xor \U$22993 ( \23370 , \23369 , \23323 );
and \U$22994 ( \23371 , \23368 , \23370 );
xor \U$22995 ( \23372 , \22693 , \22706 );
xor \U$22996 ( \23373 , \23372 , \22719 );
xor \U$22997 ( \23374 , \23333 , \23340 );
xor \U$22998 ( \23375 , \23373 , \23374 );
xor \U$22999 ( \23376 , \23086 , \23308 );
xor \U$23000 ( \23377 , \23376 , \23323 );
and \U$23001 ( \23378 , \23375 , \23377 );
and \U$23002 ( \23379 , \23368 , \23375 );
or \U$23003 ( \23380 , \23371 , \23378 , \23379 );
xor \U$23004 ( \23381 , \22890 , \22915 );
xor \U$23005 ( \23382 , \23381 , \22941 );
xor \U$23006 ( \23383 , \22747 , \22772 );
xor \U$23007 ( \23384 , \23383 , \22798 );
xor \U$23008 ( \23385 , \23382 , \23384 );
xor \U$23009 ( \23386 , \22695 , \22700 );
xor \U$23010 ( \23387 , \23386 , \22703 );
xor \U$23011 ( \23388 , \23311 , \23318 );
xor \U$23012 ( \23389 , \23387 , \23388 );
and \U$23013 ( \23390 , \23385 , \23389 );
and \U$23014 ( \23391 , \23382 , \23384 );
or \U$23015 ( \23392 , \23390 , \23391 );
not \U$23016 ( \23393 , \23392 );
not \U$23017 ( \23394 , \23306 );
not \U$23018 ( \23395 , \23230 );
or \U$23019 ( \23396 , \23394 , \23395 );
or \U$23020 ( \23397 , \23230 , \23306 );
nand \U$23021 ( \23398 , \23396 , \23397 );
not \U$23022 ( \23399 , \23398 );
not \U$23023 ( \23400 , \23144 );
and \U$23024 ( \23401 , \23399 , \23400 );
and \U$23025 ( \23402 , \23398 , \23144 );
nor \U$23026 ( \23403 , \23401 , \23402 );
not \U$23027 ( \23404 , \23403 );
xor \U$23028 ( \23405 , \23068 , \23078 );
xor \U$23029 ( \23406 , \23405 , \23083 );
nand \U$23030 ( \23407 , \23404 , \23406 );
or \U$23031 ( \23408 , \23393 , \23407 );
not \U$23032 ( \23409 , \23407 );
not \U$23033 ( \23410 , \23393 );
or \U$23034 ( \23411 , \23409 , \23410 );
not \U$23035 ( \23412 , \23151 );
xor \U$23036 ( \23413 , \23159 , \23169 );
not \U$23037 ( \23414 , \23413 );
or \U$23038 ( \23415 , \23412 , \23414 );
or \U$23039 ( \23416 , \23413 , \23151 );
nand \U$23040 ( \23417 , \23415 , \23416 );
xor \U$23041 ( \23418 , \23094 , \23102 );
xor \U$23042 ( \23419 , \23418 , \23110 );
xor \U$23043 ( \23420 , \23417 , \23419 );
xor \U$23044 ( \23421 , \23209 , \23216 );
xor \U$23045 ( \23422 , \23421 , \23224 );
and \U$23046 ( \23423 , \23420 , \23422 );
and \U$23047 ( \23424 , \23417 , \23419 );
or \U$23048 ( \23425 , \23423 , \23424 );
xor \U$23049 ( \23426 , \22754 , \22761 );
xor \U$23050 ( \23427 , \23426 , \22769 );
xor \U$23051 ( \23428 , \23425 , \23427 );
not \U$23052 ( \23429 , \23179 );
xor \U$23053 ( \23430 , \23197 , \23187 );
not \U$23054 ( \23431 , \23430 );
or \U$23055 ( \23432 , \23429 , \23431 );
or \U$23056 ( \23433 , \23430 , \23179 );
nand \U$23057 ( \23434 , \23432 , \23433 );
xor \U$23058 ( \23435 , \23285 , \23292 );
xor \U$23059 ( \23436 , \23435 , \23300 );
xor \U$23060 ( \23437 , \23434 , \23436 );
xor \U$23061 ( \23438 , \23241 , \23248 );
xor \U$23062 ( \23439 , \23438 , \23256 );
and \U$23063 ( \23440 , \23437 , \23439 );
and \U$23064 ( \23441 , \23434 , \23436 );
or \U$23065 ( \23442 , \23440 , \23441 );
and \U$23066 ( \23443 , \23428 , \23442 );
and \U$23067 ( \23444 , \23425 , \23427 );
or \U$23068 ( \23445 , \23443 , \23444 );
and \U$23069 ( \23446 , \8371 , RIae77d38_95);
and \U$23070 ( \23447 , RIae77e28_97, \8369 );
nor \U$23071 ( \23448 , \23446 , \23447 );
and \U$23072 ( \23449 , \23448 , \8020 );
not \U$23073 ( \23450 , \23448 );
and \U$23074 ( \23451 , \23450 , \8019 );
nor \U$23075 ( \23452 , \23449 , \23451 );
and \U$23076 ( \23453 , \6941 , RIae783c8_109);
and \U$23077 ( \23454 , RIae78530_112, \6939 );
nor \U$23078 ( \23455 , \23453 , \23454 );
and \U$23079 ( \23456 , \23455 , \6314 );
not \U$23080 ( \23457 , \23455 );
and \U$23081 ( \23458 , \23457 , \6945 );
nor \U$23082 ( \23459 , \23456 , \23458 );
xor \U$23083 ( \23460 , \23452 , \23459 );
and \U$23084 ( \23461 , \7633 , RIae77c48_93);
and \U$23085 ( \23462 , RIae77b58_91, \7631 );
nor \U$23086 ( \23463 , \23461 , \23462 );
and \U$23087 ( \23464 , \23463 , \7206 );
not \U$23088 ( \23465 , \23463 );
and \U$23089 ( \23466 , \23465 , \7205 );
nor \U$23090 ( \23467 , \23464 , \23466 );
and \U$23091 ( \23468 , \23460 , \23467 );
and \U$23092 ( \23469 , \23452 , \23459 );
or \U$23093 ( \23470 , \23468 , \23469 );
and \U$23094 ( \23471 , \5399 , RIae782d8_107);
and \U$23095 ( \23472 , RIae780f8_103, \5397 );
nor \U$23096 ( \23473 , \23471 , \23472 );
and \U$23097 ( \23474 , \23473 , \5016 );
not \U$23098 ( \23475 , \23473 );
and \U$23099 ( \23476 , \23475 , \5403 );
nor \U$23100 ( \23477 , \23474 , \23476 );
and \U$23101 ( \23478 , \5896 , RIae77f18_99);
and \U$23102 ( \23479 , RIae78008_101, \5894 );
nor \U$23103 ( \23480 , \23478 , \23479 );
and \U$23104 ( \23481 , \23480 , \5590 );
not \U$23105 ( \23482 , \23480 );
and \U$23106 ( \23483 , \23482 , \5589 );
nor \U$23107 ( \23484 , \23481 , \23483 );
xor \U$23108 ( \23485 , \23477 , \23484 );
and \U$23109 ( \23486 , \6172 , RIae781e8_105);
and \U$23110 ( \23487 , RIae785a8_113, \6170 );
nor \U$23111 ( \23488 , \23486 , \23487 );
and \U$23112 ( \23489 , \23488 , \6176 );
not \U$23113 ( \23490 , \23488 );
and \U$23114 ( \23491 , \23490 , \6175 );
nor \U$23115 ( \23492 , \23489 , \23491 );
and \U$23116 ( \23493 , \23485 , \23492 );
and \U$23117 ( \23494 , \23477 , \23484 );
or \U$23118 ( \23495 , \23493 , \23494 );
xor \U$23119 ( \23496 , \23470 , \23495 );
and \U$23120 ( \23497 , \4688 , RIae771f8_71);
and \U$23121 ( \23498 , RIae772e8_73, \4686 );
nor \U$23122 ( \23499 , \23497 , \23498 );
and \U$23123 ( \23500 , \23499 , \4481 );
not \U$23124 ( \23501 , \23499 );
and \U$23125 ( \23502 , \23501 , \4482 );
nor \U$23126 ( \23503 , \23500 , \23502 );
and \U$23127 ( \23504 , \3730 , RIae76d48_61);
and \U$23128 ( \23505 , RIae76c58_59, \3728 );
nor \U$23129 ( \23506 , \23504 , \23505 );
and \U$23130 ( \23507 , \23506 , \3732 );
not \U$23131 ( \23508 , \23506 );
and \U$23132 ( \23509 , \23508 , \3421 );
nor \U$23133 ( \23510 , \23507 , \23509 );
xor \U$23134 ( \23511 , \23503 , \23510 );
and \U$23135 ( \23512 , \4247 , RIae77180_70);
and \U$23136 ( \23513 , RIae77018_67, \4245 );
nor \U$23137 ( \23514 , \23512 , \23513 );
and \U$23138 ( \23515 , \23514 , \3989 );
not \U$23139 ( \23516 , \23514 );
and \U$23140 ( \23517 , \23516 , \4251 );
nor \U$23141 ( \23518 , \23515 , \23517 );
and \U$23142 ( \23519 , \23511 , \23518 );
and \U$23143 ( \23520 , \23503 , \23510 );
or \U$23144 ( \23521 , \23519 , \23520 );
and \U$23145 ( \23522 , \23496 , \23521 );
and \U$23146 ( \23523 , \23470 , \23495 );
or \U$23147 ( \23524 , \23522 , \23523 );
and \U$23148 ( \23525 , \12180 , RIae75f38_31);
and \U$23149 ( \23526 , RIae75e48_29, \12178 );
nor \U$23150 ( \23527 , \23525 , \23526 );
and \U$23151 ( \23528 , \23527 , \12184 );
not \U$23152 ( \23529 , \23527 );
and \U$23153 ( \23530 , \23529 , \11827 );
nor \U$23154 ( \23531 , \23528 , \23530 );
and \U$23155 ( \23532 , \11470 , RIae75998_19);
and \U$23156 ( \23533 , RIae758a8_17, \11468 );
nor \U$23157 ( \23534 , \23532 , \23533 );
and \U$23158 ( \23535 , \23534 , \10936 );
not \U$23159 ( \23536 , \23534 );
and \U$23160 ( \23537 , \23536 , \11474 );
nor \U$23161 ( \23538 , \23535 , \23537 );
xor \U$23162 ( \23539 , \23531 , \23538 );
and \U$23163 ( \23540 , \13059 , RIae75c68_25);
and \U$23164 ( \23541 , RIae75d58_27, \13057 );
nor \U$23165 ( \23542 , \23540 , \23541 );
and \U$23166 ( \23543 , \23542 , \13063 );
not \U$23167 ( \23544 , \23542 );
and \U$23168 ( \23545 , \23544 , \12718 );
nor \U$23169 ( \23546 , \23543 , \23545 );
and \U$23170 ( \23547 , \23539 , \23546 );
and \U$23171 ( \23548 , \23531 , \23538 );
or \U$23172 ( \23549 , \23547 , \23548 );
and \U$23173 ( \23550 , \14059 , RIae755d8_11);
and \U$23174 ( \23551 , RIae754e8_9, \14057 );
nor \U$23175 ( \23552 , \23550 , \23551 );
and \U$23176 ( \23553 , \23552 , \13502 );
not \U$23177 ( \23554 , \23552 );
and \U$23178 ( \23555 , \23554 , \14063 );
nor \U$23179 ( \23556 , \23553 , \23555 );
and \U$23180 ( \23557 , \15726 , RIae75218_3);
and \U$23181 ( \23558 , RIae7aab0_192, RIae75128_1);
nor \U$23182 ( \23559 , \23557 , \23558 );
and \U$23183 ( \23560 , \23559 , \14959 );
not \U$23184 ( \23561 , \23559 );
and \U$23185 ( \23562 , \23561 , RIae7aa38_191);
nor \U$23186 ( \23563 , \23560 , \23562 );
xor \U$23187 ( \23564 , \23556 , \23563 );
and \U$23188 ( \23565 , \14964 , RIae757b8_15);
and \U$23189 ( \23566 , RIae756c8_13, \14962 );
nor \U$23190 ( \23567 , \23565 , \23566 );
and \U$23191 ( \23568 , \23567 , \14463 );
not \U$23192 ( \23569 , \23567 );
and \U$23193 ( \23570 , \23569 , \14462 );
nor \U$23194 ( \23571 , \23568 , \23570 );
and \U$23195 ( \23572 , \23564 , \23571 );
and \U$23196 ( \23573 , \23556 , \23563 );
or \U$23197 ( \23574 , \23572 , \23573 );
xor \U$23198 ( \23575 , \23549 , \23574 );
and \U$23199 ( \23576 , \8966 , RIae78968_121);
and \U$23200 ( \23577 , RIae78878_119, \8964 );
nor \U$23201 ( \23578 , \23576 , \23577 );
and \U$23202 ( \23579 , \23578 , \8799 );
not \U$23203 ( \23580 , \23578 );
and \U$23204 ( \23581 , \23580 , \8789 );
nor \U$23205 ( \23582 , \23579 , \23581 );
and \U$23206 ( \23583 , \9760 , RIae78788_117);
and \U$23207 ( \23584 , RIae78698_115, \9758 );
nor \U$23208 ( \23585 , \23583 , \23584 );
and \U$23209 ( \23586 , \23585 , \9273 );
not \U$23210 ( \23587 , \23585 );
and \U$23211 ( \23588 , \23587 , \9272 );
nor \U$23212 ( \23589 , \23586 , \23588 );
xor \U$23213 ( \23590 , \23582 , \23589 );
and \U$23214 ( \23591 , \10548 , RIae75b78_23);
and \U$23215 ( \23592 , RIae75a88_21, \10546 );
nor \U$23216 ( \23593 , \23591 , \23592 );
and \U$23217 ( \23594 , \23593 , \10421 );
not \U$23218 ( \23595 , \23593 );
and \U$23219 ( \23596 , \23595 , \10118 );
nor \U$23220 ( \23597 , \23594 , \23596 );
and \U$23221 ( \23598 , \23590 , \23597 );
and \U$23222 ( \23599 , \23582 , \23589 );
or \U$23223 ( \23600 , \23598 , \23599 );
and \U$23224 ( \23601 , \23575 , \23600 );
and \U$23225 ( \23602 , \23549 , \23574 );
or \U$23226 ( \23603 , \23601 , \23602 );
xor \U$23227 ( \23604 , \23524 , \23603 );
and \U$23228 ( \23605 , \2607 , RIae77a68_89);
and \U$23229 ( \23606 , RIae77978_87, \2605 );
nor \U$23230 ( \23607 , \23605 , \23606 );
and \U$23231 ( \23608 , \23607 , \2611 );
not \U$23232 ( \23609 , \23607 );
and \U$23233 ( \23610 , \23609 , \2396 );
nor \U$23234 ( \23611 , \23608 , \23610 );
not \U$23235 ( \23612 , \2789 );
and \U$23236 ( \23613 , \2783 , RIae77798_83);
and \U$23237 ( \23614 , RIae77888_85, \2781 );
nor \U$23238 ( \23615 , \23613 , \23614 );
not \U$23239 ( \23616 , \23615 );
or \U$23240 ( \23617 , \23612 , \23616 );
or \U$23241 ( \23618 , \23615 , \3089 );
nand \U$23242 ( \23619 , \23617 , \23618 );
xor \U$23243 ( \23620 , \23611 , \23619 );
not \U$23244 ( \23621 , \2774 );
and \U$23245 ( \23622 , \3214 , RIae76f28_65);
and \U$23246 ( \23623 , RIae76e38_63, \3212 );
nor \U$23247 ( \23624 , \23622 , \23623 );
not \U$23248 ( \23625 , \23624 );
or \U$23249 ( \23626 , \23621 , \23625 );
or \U$23250 ( \23627 , \23624 , \3218 );
nand \U$23251 ( \23628 , \23626 , \23627 );
and \U$23252 ( \23629 , \23620 , \23628 );
and \U$23253 ( \23630 , \23611 , \23619 );
or \U$23254 ( \23631 , \23629 , \23630 );
nand \U$23255 ( \23632 , RIae775b8_79, \1591 );
and \U$23256 ( \23633 , \23632 , \1498 );
not \U$23257 ( \23634 , \23632 );
and \U$23258 ( \23635 , \23634 , \1488 );
nor \U$23259 ( \23636 , \23633 , \23635 );
xor \U$23260 ( \23637 , \23631 , \23636 );
xor \U$23261 ( \23638 , \23120 , \23127 );
xor \U$23262 ( \23639 , \23638 , \23135 );
and \U$23263 ( \23640 , \23637 , \23639 );
and \U$23264 ( \23641 , \23631 , \23636 );
or \U$23265 ( \23642 , \23640 , \23641 );
and \U$23266 ( \23643 , \23604 , \23642 );
and \U$23267 ( \23644 , \23524 , \23603 );
or \U$23268 ( \23645 , \23643 , \23644 );
xor \U$23269 ( \23646 , \23445 , \23645 );
xor \U$23270 ( \23647 , \23113 , \23138 );
xor \U$23271 ( \23648 , \23647 , \23141 );
xor \U$23272 ( \23649 , \23070 , \23072 );
xor \U$23273 ( \23650 , \23649 , \23075 );
and \U$23274 ( \23651 , \23648 , \23650 );
xor \U$23275 ( \23652 , \22808 , \22816 );
xor \U$23276 ( \23653 , \23652 , \22825 );
xor \U$23277 ( \23654 , \23058 , \23063 );
xor \U$23278 ( \23655 , \23653 , \23654 );
xor \U$23279 ( \23656 , \23070 , \23072 );
xor \U$23280 ( \23657 , \23656 , \23075 );
and \U$23281 ( \23658 , \23655 , \23657 );
and \U$23282 ( \23659 , \23648 , \23655 );
or \U$23283 ( \23660 , \23651 , \23658 , \23659 );
and \U$23284 ( \23661 , \23646 , \23660 );
and \U$23285 ( \23662 , \23445 , \23645 );
or \U$23286 ( \23663 , \23661 , \23662 );
nand \U$23287 ( \23664 , \23411 , \23663 );
nand \U$23288 ( \23665 , \23408 , \23664 );
xor \U$23289 ( \23666 , \23380 , \23665 );
xor \U$23290 ( \23667 , \23038 , \23040 );
xor \U$23291 ( \23668 , \23667 , \23045 );
and \U$23292 ( \23669 , \23666 , \23668 );
and \U$23293 ( \23670 , \23380 , \23665 );
or \U$23294 ( \23671 , \23669 , \23670 );
not \U$23295 ( \23672 , \23671 );
or \U$23296 ( \23673 , \23366 , \23672 );
or \U$23297 ( \23674 , \23671 , \23365 );
nand \U$23298 ( \23675 , \23673 , \23674 );
not \U$23299 ( \23676 , \23675 );
xnor \U$23300 ( \23677 , \23048 , \23348 );
not \U$23301 ( \23678 , \23677 );
not \U$23302 ( \23679 , \23053 );
and \U$23303 ( \23680 , \23678 , \23679 );
and \U$23304 ( \23681 , \23677 , \23053 );
nor \U$23305 ( \23682 , \23680 , \23681 );
not \U$23306 ( \23683 , \23682 );
and \U$23307 ( \23684 , \23676 , \23683 );
and \U$23308 ( \23685 , \23675 , \23682 );
nor \U$23309 ( \23686 , \23684 , \23685 );
xor \U$23310 ( \23687 , \23380 , \23665 );
xor \U$23311 ( \23688 , \23687 , \23668 );
xor \U$23312 ( \23689 , \23326 , \23328 );
xor \U$23313 ( \23690 , \23689 , \23345 );
xor \U$23314 ( \23691 , \23688 , \23690 );
not \U$23315 ( \23692 , \23403 );
not \U$23316 ( \23693 , \23406 );
or \U$23317 ( \23694 , \23692 , \23693 );
or \U$23318 ( \23695 , \23406 , \23403 );
nand \U$23319 ( \23696 , \23694 , \23695 );
xor \U$23320 ( \23697 , \23382 , \23384 );
xor \U$23321 ( \23698 , \23697 , \23389 );
and \U$23322 ( \23699 , \23696 , \23698 );
xor \U$23323 ( \23700 , \23445 , \23645 );
xor \U$23324 ( \23701 , \23700 , \23660 );
xor \U$23325 ( \23702 , \23382 , \23384 );
xor \U$23326 ( \23703 , \23702 , \23389 );
and \U$23327 ( \23704 , \23701 , \23703 );
and \U$23328 ( \23705 , \23696 , \23701 );
or \U$23329 ( \23706 , \23699 , \23704 , \23705 );
not \U$23330 ( \23707 , \23706 );
xor \U$23331 ( \23708 , \23086 , \23308 );
xor \U$23332 ( \23709 , \23708 , \23323 );
xor \U$23333 ( \23710 , \23368 , \23375 );
xor \U$23334 ( \23711 , \23709 , \23710 );
not \U$23335 ( \23712 , \23711 );
or \U$23336 ( \23713 , \23707 , \23712 );
or \U$23337 ( \23714 , \23711 , \23706 );
xor \U$23338 ( \23715 , \23503 , \23510 );
xor \U$23339 ( \23716 , \23715 , \23518 );
and \U$23340 ( \23717 , \1939 , RIae775b8_79);
and \U$23341 ( \23718 , RIae774c8_77, \1937 );
nor \U$23342 ( \23719 , \23717 , \23718 );
and \U$23343 ( \23720 , \23719 , \1735 );
not \U$23344 ( \23721 , \23719 );
and \U$23345 ( \23722 , \23721 , \1734 );
nor \U$23346 ( \23723 , \23720 , \23722 );
xor \U$23347 ( \23724 , \23716 , \23723 );
xor \U$23348 ( \23725 , \23611 , \23619 );
xor \U$23349 ( \23726 , \23725 , \23628 );
and \U$23350 ( \23727 , \23724 , \23726 );
and \U$23351 ( \23728 , \23716 , \23723 );
or \U$23352 ( \23729 , \23727 , \23728 );
xor \U$23353 ( \23730 , \23266 , \1488 );
xor \U$23354 ( \23731 , \23730 , \23274 );
xor \U$23355 ( \23732 , \23729 , \23731 );
xor \U$23356 ( \23733 , \23477 , \23484 );
xor \U$23357 ( \23734 , \23733 , \23492 );
xor \U$23358 ( \23735 , \23452 , \23459 );
xor \U$23359 ( \23736 , \23735 , \23467 );
and \U$23360 ( \23737 , \23734 , \23736 );
xor \U$23361 ( \23738 , \23582 , \23589 );
xor \U$23362 ( \23739 , \23738 , \23597 );
xor \U$23363 ( \23740 , \23452 , \23459 );
xor \U$23364 ( \23741 , \23740 , \23467 );
and \U$23365 ( \23742 , \23739 , \23741 );
and \U$23366 ( \23743 , \23734 , \23739 );
or \U$23367 ( \23744 , \23737 , \23742 , \23743 );
and \U$23368 ( \23745 , \23732 , \23744 );
and \U$23369 ( \23746 , \23729 , \23731 );
or \U$23370 ( \23747 , \23745 , \23746 );
and \U$23371 ( \23748 , \11470 , RIae75a88_21);
and \U$23372 ( \23749 , RIae75998_19, \11468 );
nor \U$23373 ( \23750 , \23748 , \23749 );
and \U$23374 ( \23751 , \23750 , \10936 );
not \U$23375 ( \23752 , \23750 );
and \U$23376 ( \23753 , \23752 , \11474 );
nor \U$23377 ( \23754 , \23751 , \23753 );
and \U$23378 ( \23755 , \9760 , RIae78878_119);
and \U$23379 ( \23756 , RIae78788_117, \9758 );
nor \U$23380 ( \23757 , \23755 , \23756 );
and \U$23381 ( \23758 , \23757 , \9273 );
not \U$23382 ( \23759 , \23757 );
and \U$23383 ( \23760 , \23759 , \9764 );
nor \U$23384 ( \23761 , \23758 , \23760 );
xor \U$23385 ( \23762 , \23754 , \23761 );
and \U$23386 ( \23763 , \10548 , RIae78698_115);
and \U$23387 ( \23764 , RIae75b78_23, \10546 );
nor \U$23388 ( \23765 , \23763 , \23764 );
and \U$23389 ( \23766 , \23765 , \10421 );
not \U$23390 ( \23767 , \23765 );
and \U$23391 ( \23768 , \23767 , \10118 );
nor \U$23392 ( \23769 , \23766 , \23768 );
and \U$23393 ( \23770 , \23762 , \23769 );
and \U$23394 ( \23771 , \23754 , \23761 );
or \U$23395 ( \23772 , \23770 , \23771 );
and \U$23396 ( \23773 , \15726 , RIae756c8_13);
and \U$23397 ( \23774 , RIae7aab0_192, RIae75218_3);
nor \U$23398 ( \23775 , \23773 , \23774 );
and \U$23399 ( \23776 , \23775 , \14959 );
not \U$23400 ( \23777 , \23775 );
and \U$23401 ( \23778 , \23777 , RIae7aa38_191);
nor \U$23402 ( \23779 , \23776 , \23778 );
xor \U$23403 ( \23780 , \23779 , \1734 );
and \U$23404 ( \23781 , \14964 , RIae754e8_9);
and \U$23405 ( \23782 , RIae757b8_15, \14962 );
nor \U$23406 ( \23783 , \23781 , \23782 );
and \U$23407 ( \23784 , \23783 , \14463 );
not \U$23408 ( \23785 , \23783 );
and \U$23409 ( \23786 , \23785 , \14462 );
nor \U$23410 ( \23787 , \23784 , \23786 );
and \U$23411 ( \23788 , \23780 , \23787 );
and \U$23412 ( \23789 , \23779 , \1734 );
or \U$23413 ( \23790 , \23788 , \23789 );
xor \U$23414 ( \23791 , \23772 , \23790 );
and \U$23415 ( \23792 , \12180 , RIae758a8_17);
and \U$23416 ( \23793 , RIae75f38_31, \12178 );
nor \U$23417 ( \23794 , \23792 , \23793 );
and \U$23418 ( \23795 , \23794 , \12184 );
not \U$23419 ( \23796 , \23794 );
and \U$23420 ( \23797 , \23796 , \11827 );
nor \U$23421 ( \23798 , \23795 , \23797 );
and \U$23422 ( \23799 , \13059 , RIae75e48_29);
and \U$23423 ( \23800 , RIae75c68_25, \13057 );
nor \U$23424 ( \23801 , \23799 , \23800 );
and \U$23425 ( \23802 , \23801 , \13063 );
not \U$23426 ( \23803 , \23801 );
and \U$23427 ( \23804 , \23803 , \12718 );
nor \U$23428 ( \23805 , \23802 , \23804 );
xor \U$23429 ( \23806 , \23798 , \23805 );
and \U$23430 ( \23807 , \14059 , RIae75d58_27);
and \U$23431 ( \23808 , RIae755d8_11, \14057 );
nor \U$23432 ( \23809 , \23807 , \23808 );
and \U$23433 ( \23810 , \23809 , \13502 );
not \U$23434 ( \23811 , \23809 );
and \U$23435 ( \23812 , \23811 , \14063 );
nor \U$23436 ( \23813 , \23810 , \23812 );
and \U$23437 ( \23814 , \23806 , \23813 );
and \U$23438 ( \23815 , \23798 , \23805 );
or \U$23439 ( \23816 , \23814 , \23815 );
and \U$23440 ( \23817 , \23791 , \23816 );
and \U$23441 ( \23818 , \23772 , \23790 );
or \U$23442 ( \23819 , \23817 , \23818 );
and \U$23443 ( \23820 , \2607 , RIae773d8_75);
and \U$23444 ( \23821 , RIae77a68_89, \2605 );
nor \U$23445 ( \23822 , \23820 , \23821 );
and \U$23446 ( \23823 , \23822 , \2611 );
not \U$23447 ( \23824 , \23822 );
and \U$23448 ( \23825 , \23824 , \2397 );
nor \U$23449 ( \23826 , \23823 , \23825 );
nand \U$23450 ( \23827 , RIae775b8_79, \1937 );
and \U$23451 ( \23828 , \23827 , \1735 );
not \U$23452 ( \23829 , \23827 );
and \U$23453 ( \23830 , \23829 , \1734 );
nor \U$23454 ( \23831 , \23828 , \23830 );
xor \U$23455 ( \23832 , \23826 , \23831 );
and \U$23456 ( \23833 , \2224 , RIae774c8_77);
and \U$23457 ( \23834 , RIae77720_82, \2222 );
nor \U$23458 ( \23835 , \23833 , \23834 );
and \U$23459 ( \23836 , \23835 , \2061 );
not \U$23460 ( \23837 , \23835 );
and \U$23461 ( \23838 , \23837 , \2060 );
nor \U$23462 ( \23839 , \23836 , \23838 );
and \U$23463 ( \23840 , \23832 , \23839 );
and \U$23464 ( \23841 , \23826 , \23831 );
or \U$23465 ( \23842 , \23840 , \23841 );
and \U$23466 ( \23843 , \2224 , RIae77720_82);
and \U$23467 ( \23844 , RIae773d8_75, \2222 );
nor \U$23468 ( \23845 , \23843 , \23844 );
and \U$23469 ( \23846 , \23845 , \2061 );
not \U$23470 ( \23847 , \23845 );
and \U$23471 ( \23848 , \23847 , \2060 );
nor \U$23472 ( \23849 , \23846 , \23848 );
xor \U$23473 ( \23850 , \23842 , \23849 );
not \U$23474 ( \23851 , \3089 );
and \U$23475 ( \23852 , \2783 , RIae77978_87);
and \U$23476 ( \23853 , RIae77798_83, \2781 );
nor \U$23477 ( \23854 , \23852 , \23853 );
not \U$23478 ( \23855 , \23854 );
or \U$23479 ( \23856 , \23851 , \23855 );
or \U$23480 ( \23857 , \23854 , \2789 );
nand \U$23481 ( \23858 , \23856 , \23857 );
not \U$23482 ( \23859 , \3218 );
and \U$23483 ( \23860 , \3214 , RIae77888_85);
and \U$23484 ( \23861 , RIae76f28_65, \3212 );
nor \U$23485 ( \23862 , \23860 , \23861 );
not \U$23486 ( \23863 , \23862 );
or \U$23487 ( \23864 , \23859 , \23863 );
or \U$23488 ( \23865 , \23862 , \2774 );
nand \U$23489 ( \23866 , \23864 , \23865 );
xor \U$23490 ( \23867 , \23858 , \23866 );
and \U$23491 ( \23868 , \3730 , RIae76e38_63);
and \U$23492 ( \23869 , RIae76d48_61, \3728 );
nor \U$23493 ( \23870 , \23868 , \23869 );
and \U$23494 ( \23871 , \23870 , \3732 );
not \U$23495 ( \23872 , \23870 );
and \U$23496 ( \23873 , \23872 , \3422 );
nor \U$23497 ( \23874 , \23871 , \23873 );
and \U$23498 ( \23875 , \23867 , \23874 );
and \U$23499 ( \23876 , \23858 , \23866 );
or \U$23500 ( \23877 , \23875 , \23876 );
and \U$23501 ( \23878 , \23850 , \23877 );
and \U$23502 ( \23879 , \23842 , \23849 );
or \U$23503 ( \23880 , \23878 , \23879 );
xor \U$23504 ( \23881 , \23819 , \23880 );
and \U$23505 ( \23882 , \7633 , RIae78530_112);
and \U$23506 ( \23883 , RIae77c48_93, \7631 );
nor \U$23507 ( \23884 , \23882 , \23883 );
and \U$23508 ( \23885 , \23884 , \7206 );
not \U$23509 ( \23886 , \23884 );
and \U$23510 ( \23887 , \23886 , \7205 );
nor \U$23511 ( \23888 , \23885 , \23887 );
and \U$23512 ( \23889 , \8371 , RIae77b58_91);
and \U$23513 ( \23890 , RIae77d38_95, \8369 );
nor \U$23514 ( \23891 , \23889 , \23890 );
and \U$23515 ( \23892 , \23891 , \8020 );
not \U$23516 ( \23893 , \23891 );
and \U$23517 ( \23894 , \23893 , \8019 );
nor \U$23518 ( \23895 , \23892 , \23894 );
xor \U$23519 ( \23896 , \23888 , \23895 );
and \U$23520 ( \23897 , \8966 , RIae77e28_97);
and \U$23521 ( \23898 , RIae78968_121, \8964 );
nor \U$23522 ( \23899 , \23897 , \23898 );
and \U$23523 ( \23900 , \23899 , \8799 );
not \U$23524 ( \23901 , \23899 );
and \U$23525 ( \23902 , \23901 , \8789 );
nor \U$23526 ( \23903 , \23900 , \23902 );
and \U$23527 ( \23904 , \23896 , \23903 );
and \U$23528 ( \23905 , \23888 , \23895 );
or \U$23529 ( \23906 , \23904 , \23905 );
and \U$23530 ( \23907 , \4247 , RIae76c58_59);
and \U$23531 ( \23908 , RIae77180_70, \4245 );
nor \U$23532 ( \23909 , \23907 , \23908 );
and \U$23533 ( \23910 , \23909 , \3989 );
not \U$23534 ( \23911 , \23909 );
and \U$23535 ( \23912 , \23911 , \4251 );
nor \U$23536 ( \23913 , \23910 , \23912 );
and \U$23537 ( \23914 , \4688 , RIae77018_67);
and \U$23538 ( \23915 , RIae771f8_71, \4686 );
nor \U$23539 ( \23916 , \23914 , \23915 );
and \U$23540 ( \23917 , \23916 , \4481 );
not \U$23541 ( \23918 , \23916 );
and \U$23542 ( \23919 , \23918 , \4482 );
nor \U$23543 ( \23920 , \23917 , \23919 );
xor \U$23544 ( \23921 , \23913 , \23920 );
and \U$23545 ( \23922 , \5399 , RIae772e8_73);
and \U$23546 ( \23923 , RIae782d8_107, \5397 );
nor \U$23547 ( \23924 , \23922 , \23923 );
and \U$23548 ( \23925 , \23924 , \5016 );
not \U$23549 ( \23926 , \23924 );
and \U$23550 ( \23927 , \23926 , \5403 );
nor \U$23551 ( \23928 , \23925 , \23927 );
and \U$23552 ( \23929 , \23921 , \23928 );
and \U$23553 ( \23930 , \23913 , \23920 );
or \U$23554 ( \23931 , \23929 , \23930 );
xor \U$23555 ( \23932 , \23906 , \23931 );
and \U$23556 ( \23933 , \5896 , RIae780f8_103);
and \U$23557 ( \23934 , RIae77f18_99, \5894 );
nor \U$23558 ( \23935 , \23933 , \23934 );
and \U$23559 ( \23936 , \23935 , \5590 );
not \U$23560 ( \23937 , \23935 );
and \U$23561 ( \23938 , \23937 , \5589 );
nor \U$23562 ( \23939 , \23936 , \23938 );
and \U$23563 ( \23940 , \6172 , RIae78008_101);
and \U$23564 ( \23941 , RIae781e8_105, \6170 );
nor \U$23565 ( \23942 , \23940 , \23941 );
and \U$23566 ( \23943 , \23942 , \6176 );
not \U$23567 ( \23944 , \23942 );
and \U$23568 ( \23945 , \23944 , \6175 );
nor \U$23569 ( \23946 , \23943 , \23945 );
xor \U$23570 ( \23947 , \23939 , \23946 );
and \U$23571 ( \23948 , \6941 , RIae785a8_113);
and \U$23572 ( \23949 , RIae783c8_109, \6939 );
nor \U$23573 ( \23950 , \23948 , \23949 );
and \U$23574 ( \23951 , \23950 , \6314 );
not \U$23575 ( \23952 , \23950 );
and \U$23576 ( \23953 , \23952 , \6945 );
nor \U$23577 ( \23954 , \23951 , \23953 );
and \U$23578 ( \23955 , \23947 , \23954 );
and \U$23579 ( \23956 , \23939 , \23946 );
or \U$23580 ( \23957 , \23955 , \23956 );
and \U$23581 ( \23958 , \23932 , \23957 );
and \U$23582 ( \23959 , \23906 , \23931 );
or \U$23583 ( \23960 , \23958 , \23959 );
and \U$23584 ( \23961 , \23881 , \23960 );
and \U$23585 ( \23962 , \23819 , \23880 );
or \U$23586 ( \23963 , \23961 , \23962 );
xor \U$23587 ( \23964 , \23747 , \23963 );
xor \U$23588 ( \23965 , \23631 , \23636 );
xor \U$23589 ( \23966 , \23965 , \23639 );
xor \U$23590 ( \23967 , \23417 , \23419 );
xor \U$23591 ( \23968 , \23967 , \23422 );
and \U$23592 ( \23969 , \23966 , \23968 );
xor \U$23593 ( \23970 , \23434 , \23436 );
xor \U$23594 ( \23971 , \23970 , \23439 );
xor \U$23595 ( \23972 , \23417 , \23419 );
xor \U$23596 ( \23973 , \23972 , \23422 );
and \U$23597 ( \23974 , \23971 , \23973 );
and \U$23598 ( \23975 , \23966 , \23971 );
or \U$23599 ( \23976 , \23969 , \23974 , \23975 );
and \U$23600 ( \23977 , \23964 , \23976 );
and \U$23601 ( \23978 , \23747 , \23963 );
or \U$23602 ( \23979 , \23977 , \23978 );
xor \U$23603 ( \23980 , \23524 , \23603 );
xor \U$23604 ( \23981 , \23980 , \23642 );
xor \U$23605 ( \23982 , \23425 , \23427 );
xor \U$23606 ( \23983 , \23982 , \23442 );
and \U$23607 ( \23984 , \23981 , \23983 );
xor \U$23608 ( \23985 , \23979 , \23984 );
not \U$23609 ( \23986 , \23199 );
not \U$23610 ( \23987 , \23227 );
not \U$23611 ( \23988 , \23171 );
or \U$23612 ( \23989 , \23987 , \23988 );
or \U$23613 ( \23990 , \23171 , \23227 );
nand \U$23614 ( \23991 , \23989 , \23990 );
not \U$23615 ( \23992 , \23991 );
or \U$23616 ( \23993 , \23986 , \23992 );
or \U$23617 ( \23994 , \23991 , \23199 );
nand \U$23618 ( \23995 , \23993 , \23994 );
xor \U$23619 ( \23996 , \23259 , \23277 );
xor \U$23620 ( \23997 , \23996 , \23303 );
xor \U$23621 ( \23998 , \23995 , \23997 );
xor \U$23622 ( \23999 , \23070 , \23072 );
xor \U$23623 ( \24000 , \23999 , \23075 );
xor \U$23624 ( \24001 , \23648 , \23655 );
xor \U$23625 ( \24002 , \24000 , \24001 );
and \U$23626 ( \24003 , \23998 , \24002 );
and \U$23627 ( \24004 , \23995 , \23997 );
or \U$23628 ( \24005 , \24003 , \24004 );
and \U$23629 ( \24006 , \23985 , \24005 );
and \U$23630 ( \24007 , \23979 , \23984 );
or \U$23631 ( \24008 , \24006 , \24007 );
nand \U$23632 ( \24009 , \23714 , \24008 );
nand \U$23633 ( \24010 , \23713 , \24009 );
and \U$23634 ( \24011 , \23691 , \24010 );
and \U$23635 ( \24012 , \23688 , \23690 );
nor \U$23636 ( \24013 , \24011 , \24012 );
or \U$23637 ( \24014 , \23686 , \24013 );
xnor \U$23638 ( \24015 , \24013 , \23686 );
not \U$23639 ( \24016 , \23663 );
not \U$23640 ( \24017 , \23393 );
or \U$23641 ( \24018 , \24016 , \24017 );
or \U$23642 ( \24019 , \23393 , \23663 );
nand \U$23643 ( \24020 , \24018 , \24019 );
not \U$23644 ( \24021 , \24020 );
not \U$23645 ( \24022 , \23407 );
and \U$23646 ( \24023 , \24021 , \24022 );
and \U$23647 ( \24024 , \24020 , \23407 );
nor \U$23648 ( \24025 , \24023 , \24024 );
not \U$23649 ( \24026 , \24025 );
xor \U$23650 ( \24027 , \23754 , \23761 );
xor \U$23651 ( \24028 , \24027 , \23769 );
xor \U$23652 ( \24029 , \23779 , \1734 );
xor \U$23653 ( \24030 , \24029 , \23787 );
and \U$23654 ( \24031 , \24028 , \24030 );
xor \U$23655 ( \24032 , \23798 , \23805 );
xor \U$23656 ( \24033 , \24032 , \23813 );
xor \U$23657 ( \24034 , \23779 , \1734 );
xor \U$23658 ( \24035 , \24034 , \23787 );
and \U$23659 ( \24036 , \24033 , \24035 );
and \U$23660 ( \24037 , \24028 , \24033 );
or \U$23661 ( \24038 , \24031 , \24036 , \24037 );
xor \U$23662 ( \24039 , \23531 , \23538 );
xor \U$23663 ( \24040 , \24039 , \23546 );
xor \U$23664 ( \24041 , \24038 , \24040 );
xor \U$23665 ( \24042 , \23913 , \23920 );
xor \U$23666 ( \24043 , \24042 , \23928 );
xor \U$23667 ( \24044 , \23939 , \23946 );
xor \U$23668 ( \24045 , \24044 , \23954 );
xor \U$23669 ( \24046 , \24043 , \24045 );
xor \U$23670 ( \24047 , \23888 , \23895 );
xor \U$23671 ( \24048 , \24047 , \23903 );
and \U$23672 ( \24049 , \24046 , \24048 );
and \U$23673 ( \24050 , \24043 , \24045 );
or \U$23674 ( \24051 , \24049 , \24050 );
and \U$23675 ( \24052 , \24041 , \24051 );
and \U$23676 ( \24053 , \24038 , \24040 );
or \U$23677 ( \24054 , \24052 , \24053 );
and \U$23678 ( \24055 , \5896 , RIae782d8_107);
and \U$23679 ( \24056 , RIae780f8_103, \5894 );
nor \U$23680 ( \24057 , \24055 , \24056 );
and \U$23681 ( \24058 , \24057 , \5590 );
not \U$23682 ( \24059 , \24057 );
and \U$23683 ( \24060 , \24059 , \5589 );
nor \U$23684 ( \24061 , \24058 , \24060 );
and \U$23685 ( \24062 , \5399 , RIae771f8_71);
and \U$23686 ( \24063 , RIae772e8_73, \5397 );
nor \U$23687 ( \24064 , \24062 , \24063 );
and \U$23688 ( \24065 , \24064 , \5016 );
not \U$23689 ( \24066 , \24064 );
and \U$23690 ( \24067 , \24066 , \5403 );
nor \U$23691 ( \24068 , \24065 , \24067 );
xor \U$23692 ( \24069 , \24061 , \24068 );
and \U$23693 ( \24070 , \6172 , RIae77f18_99);
and \U$23694 ( \24071 , RIae78008_101, \6170 );
nor \U$23695 ( \24072 , \24070 , \24071 );
and \U$23696 ( \24073 , \24072 , \6176 );
not \U$23697 ( \24074 , \24072 );
and \U$23698 ( \24075 , \24074 , \6175 );
nor \U$23699 ( \24076 , \24073 , \24075 );
and \U$23700 ( \24077 , \24069 , \24076 );
and \U$23701 ( \24078 , \24061 , \24068 );
or \U$23702 ( \24079 , \24077 , \24078 );
and \U$23703 ( \24080 , \3730 , RIae76f28_65);
and \U$23704 ( \24081 , RIae76e38_63, \3728 );
nor \U$23705 ( \24082 , \24080 , \24081 );
and \U$23706 ( \24083 , \24082 , \3732 );
not \U$23707 ( \24084 , \24082 );
and \U$23708 ( \24085 , \24084 , \3422 );
nor \U$23709 ( \24086 , \24083 , \24085 );
and \U$23710 ( \24087 , \4247 , RIae76d48_61);
and \U$23711 ( \24088 , RIae76c58_59, \4245 );
nor \U$23712 ( \24089 , \24087 , \24088 );
and \U$23713 ( \24090 , \24089 , \3989 );
not \U$23714 ( \24091 , \24089 );
and \U$23715 ( \24092 , \24091 , \4251 );
nor \U$23716 ( \24093 , \24090 , \24092 );
xor \U$23717 ( \24094 , \24086 , \24093 );
and \U$23718 ( \24095 , \4688 , RIae77180_70);
and \U$23719 ( \24096 , RIae77018_67, \4686 );
nor \U$23720 ( \24097 , \24095 , \24096 );
and \U$23721 ( \24098 , \24097 , \4481 );
not \U$23722 ( \24099 , \24097 );
and \U$23723 ( \24100 , \24099 , \4482 );
nor \U$23724 ( \24101 , \24098 , \24100 );
and \U$23725 ( \24102 , \24094 , \24101 );
and \U$23726 ( \24103 , \24086 , \24093 );
or \U$23727 ( \24104 , \24102 , \24103 );
xor \U$23728 ( \24105 , \24079 , \24104 );
and \U$23729 ( \24106 , \8371 , RIae77c48_93);
and \U$23730 ( \24107 , RIae77b58_91, \8369 );
nor \U$23731 ( \24108 , \24106 , \24107 );
and \U$23732 ( \24109 , \24108 , \8020 );
not \U$23733 ( \24110 , \24108 );
and \U$23734 ( \24111 , \24110 , \8019 );
nor \U$23735 ( \24112 , \24109 , \24111 );
and \U$23736 ( \24113 , \6941 , RIae781e8_105);
and \U$23737 ( \24114 , RIae785a8_113, \6939 );
nor \U$23738 ( \24115 , \24113 , \24114 );
and \U$23739 ( \24116 , \24115 , \6314 );
not \U$23740 ( \24117 , \24115 );
and \U$23741 ( \24118 , \24117 , \6945 );
nor \U$23742 ( \24119 , \24116 , \24118 );
xor \U$23743 ( \24120 , \24112 , \24119 );
and \U$23744 ( \24121 , \7633 , RIae783c8_109);
and \U$23745 ( \24122 , RIae78530_112, \7631 );
nor \U$23746 ( \24123 , \24121 , \24122 );
and \U$23747 ( \24124 , \24123 , \7206 );
not \U$23748 ( \24125 , \24123 );
and \U$23749 ( \24126 , \24125 , \7205 );
nor \U$23750 ( \24127 , \24124 , \24126 );
and \U$23751 ( \24128 , \24120 , \24127 );
and \U$23752 ( \24129 , \24112 , \24119 );
or \U$23753 ( \24130 , \24128 , \24129 );
and \U$23754 ( \24131 , \24105 , \24130 );
and \U$23755 ( \24132 , \24079 , \24104 );
or \U$23756 ( \24133 , \24131 , \24132 );
and \U$23757 ( \24134 , \11470 , RIae75b78_23);
and \U$23758 ( \24135 , RIae75a88_21, \11468 );
nor \U$23759 ( \24136 , \24134 , \24135 );
and \U$23760 ( \24137 , \24136 , \10936 );
not \U$23761 ( \24138 , \24136 );
and \U$23762 ( \24139 , \24138 , \11474 );
nor \U$23763 ( \24140 , \24137 , \24139 );
and \U$23764 ( \24141 , \12180 , RIae75998_19);
and \U$23765 ( \24142 , RIae758a8_17, \12178 );
nor \U$23766 ( \24143 , \24141 , \24142 );
and \U$23767 ( \24144 , \24143 , \12184 );
not \U$23768 ( \24145 , \24143 );
and \U$23769 ( \24146 , \24145 , \11827 );
nor \U$23770 ( \24147 , \24144 , \24146 );
xor \U$23771 ( \24148 , \24140 , \24147 );
and \U$23772 ( \24149 , \13059 , RIae75f38_31);
and \U$23773 ( \24150 , RIae75e48_29, \13057 );
nor \U$23774 ( \24151 , \24149 , \24150 );
and \U$23775 ( \24152 , \24151 , \13063 );
not \U$23776 ( \24153 , \24151 );
and \U$23777 ( \24154 , \24153 , \12718 );
nor \U$23778 ( \24155 , \24152 , \24154 );
and \U$23779 ( \24156 , \24148 , \24155 );
and \U$23780 ( \24157 , \24140 , \24147 );
or \U$23781 ( \24158 , \24156 , \24157 );
and \U$23782 ( \24159 , \14059 , RIae75c68_25);
and \U$23783 ( \24160 , RIae75d58_27, \14057 );
nor \U$23784 ( \24161 , \24159 , \24160 );
and \U$23785 ( \24162 , \24161 , \13502 );
not \U$23786 ( \24163 , \24161 );
and \U$23787 ( \24164 , \24163 , \14063 );
nor \U$23788 ( \24165 , \24162 , \24164 );
and \U$23789 ( \24166 , \15726 , RIae757b8_15);
and \U$23790 ( \24167 , RIae7aab0_192, RIae756c8_13);
nor \U$23791 ( \24168 , \24166 , \24167 );
and \U$23792 ( \24169 , \24168 , \14959 );
not \U$23793 ( \24170 , \24168 );
and \U$23794 ( \24171 , \24170 , RIae7aa38_191);
nor \U$23795 ( \24172 , \24169 , \24171 );
xor \U$23796 ( \24173 , \24165 , \24172 );
and \U$23797 ( \24174 , \14964 , RIae755d8_11);
and \U$23798 ( \24175 , RIae754e8_9, \14962 );
nor \U$23799 ( \24176 , \24174 , \24175 );
and \U$23800 ( \24177 , \24176 , \14463 );
not \U$23801 ( \24178 , \24176 );
and \U$23802 ( \24179 , \24178 , \14462 );
nor \U$23803 ( \24180 , \24177 , \24179 );
and \U$23804 ( \24181 , \24173 , \24180 );
and \U$23805 ( \24182 , \24165 , \24172 );
or \U$23806 ( \24183 , \24181 , \24182 );
xor \U$23807 ( \24184 , \24158 , \24183 );
and \U$23808 ( \24185 , \10548 , RIae78788_117);
and \U$23809 ( \24186 , RIae78698_115, \10546 );
nor \U$23810 ( \24187 , \24185 , \24186 );
and \U$23811 ( \24188 , \24187 , \10421 );
not \U$23812 ( \24189 , \24187 );
and \U$23813 ( \24190 , \24189 , \10118 );
nor \U$23814 ( \24191 , \24188 , \24190 );
and \U$23815 ( \24192 , \8966 , RIae77d38_95);
and \U$23816 ( \24193 , RIae77e28_97, \8964 );
nor \U$23817 ( \24194 , \24192 , \24193 );
and \U$23818 ( \24195 , \24194 , \8799 );
not \U$23819 ( \24196 , \24194 );
and \U$23820 ( \24197 , \24196 , \8789 );
nor \U$23821 ( \24198 , \24195 , \24197 );
xor \U$23822 ( \24199 , \24191 , \24198 );
and \U$23823 ( \24200 , \9760 , RIae78968_121);
and \U$23824 ( \24201 , RIae78878_119, \9758 );
nor \U$23825 ( \24202 , \24200 , \24201 );
and \U$23826 ( \24203 , \24202 , \9273 );
not \U$23827 ( \24204 , \24202 );
and \U$23828 ( \24205 , \24204 , \9764 );
nor \U$23829 ( \24206 , \24203 , \24205 );
and \U$23830 ( \24207 , \24199 , \24206 );
and \U$23831 ( \24208 , \24191 , \24198 );
or \U$23832 ( \24209 , \24207 , \24208 );
and \U$23833 ( \24210 , \24184 , \24209 );
and \U$23834 ( \24211 , \24158 , \24183 );
or \U$23835 ( \24212 , \24210 , \24211 );
xor \U$23836 ( \24213 , \24133 , \24212 );
and \U$23837 ( \24214 , \2607 , RIae77720_82);
and \U$23838 ( \24215 , RIae773d8_75, \2605 );
nor \U$23839 ( \24216 , \24214 , \24215 );
and \U$23840 ( \24217 , \24216 , \2611 );
not \U$23841 ( \24218 , \24216 );
and \U$23842 ( \24219 , \24218 , \2397 );
nor \U$23843 ( \24220 , \24217 , \24219 );
not \U$23844 ( \24221 , \3089 );
and \U$23845 ( \24222 , \2783 , RIae77a68_89);
and \U$23846 ( \24223 , RIae77978_87, \2781 );
nor \U$23847 ( \24224 , \24222 , \24223 );
not \U$23848 ( \24225 , \24224 );
or \U$23849 ( \24226 , \24221 , \24225 );
or \U$23850 ( \24227 , \24224 , \2789 );
nand \U$23851 ( \24228 , \24226 , \24227 );
xor \U$23852 ( \24229 , \24220 , \24228 );
not \U$23853 ( \24230 , \3218 );
and \U$23854 ( \24231 , \3214 , RIae77798_83);
and \U$23855 ( \24232 , RIae77888_85, \3212 );
nor \U$23856 ( \24233 , \24231 , \24232 );
not \U$23857 ( \24234 , \24233 );
or \U$23858 ( \24235 , \24230 , \24234 );
or \U$23859 ( \24236 , \24233 , \2774 );
nand \U$23860 ( \24237 , \24235 , \24236 );
and \U$23861 ( \24238 , \24229 , \24237 );
and \U$23862 ( \24239 , \24220 , \24228 );
or \U$23863 ( \24240 , \24238 , \24239 );
xor \U$23864 ( \24241 , \23858 , \23866 );
xor \U$23865 ( \24242 , \24241 , \23874 );
and \U$23866 ( \24243 , \24240 , \24242 );
xor \U$23867 ( \24244 , \23826 , \23831 );
xor \U$23868 ( \24245 , \24244 , \23839 );
xor \U$23869 ( \24246 , \23858 , \23866 );
xor \U$23870 ( \24247 , \24246 , \23874 );
and \U$23871 ( \24248 , \24245 , \24247 );
and \U$23872 ( \24249 , \24240 , \24245 );
or \U$23873 ( \24250 , \24243 , \24248 , \24249 );
and \U$23874 ( \24251 , \24213 , \24250 );
and \U$23875 ( \24252 , \24133 , \24212 );
or \U$23876 ( \24253 , \24251 , \24252 );
xor \U$23877 ( \24254 , \24054 , \24253 );
xor \U$23878 ( \24255 , \23556 , \23563 );
xor \U$23879 ( \24256 , \24255 , \23571 );
xor \U$23880 ( \24257 , \23716 , \23723 );
xor \U$23881 ( \24258 , \24257 , \23726 );
and \U$23882 ( \24259 , \24256 , \24258 );
xor \U$23883 ( \24260 , \23452 , \23459 );
xor \U$23884 ( \24261 , \24260 , \23467 );
xor \U$23885 ( \24262 , \23734 , \23739 );
xor \U$23886 ( \24263 , \24261 , \24262 );
xor \U$23887 ( \24264 , \23716 , \23723 );
xor \U$23888 ( \24265 , \24264 , \23726 );
and \U$23889 ( \24266 , \24263 , \24265 );
and \U$23890 ( \24267 , \24256 , \24263 );
or \U$23891 ( \24268 , \24259 , \24266 , \24267 );
and \U$23892 ( \24269 , \24254 , \24268 );
and \U$23893 ( \24270 , \24054 , \24253 );
or \U$23894 ( \24271 , \24269 , \24270 );
xor \U$23895 ( \24272 , \23549 , \23574 );
xor \U$23896 ( \24273 , \24272 , \23600 );
xor \U$23897 ( \24274 , \23470 , \23495 );
xor \U$23898 ( \24275 , \24274 , \23521 );
and \U$23899 ( \24276 , \24273 , \24275 );
xor \U$23900 ( \24277 , \23842 , \23849 );
xor \U$23901 ( \24278 , \24277 , \23877 );
xor \U$23902 ( \24279 , \23772 , \23790 );
xor \U$23903 ( \24280 , \24279 , \23816 );
xor \U$23904 ( \24281 , \24278 , \24280 );
xor \U$23905 ( \24282 , \23906 , \23931 );
xor \U$23906 ( \24283 , \24282 , \23957 );
and \U$23907 ( \24284 , \24281 , \24283 );
and \U$23908 ( \24285 , \24278 , \24280 );
or \U$23909 ( \24286 , \24284 , \24285 );
xor \U$23910 ( \24287 , \23470 , \23495 );
xor \U$23911 ( \24288 , \24287 , \23521 );
and \U$23912 ( \24289 , \24286 , \24288 );
and \U$23913 ( \24290 , \24273 , \24286 );
or \U$23914 ( \24291 , \24276 , \24289 , \24290 );
xor \U$23915 ( \24292 , \24271 , \24291 );
xor \U$23916 ( \24293 , \23819 , \23880 );
xor \U$23917 ( \24294 , \24293 , \23960 );
xor \U$23918 ( \24295 , \23729 , \23731 );
xor \U$23919 ( \24296 , \24295 , \23744 );
and \U$23920 ( \24297 , \24294 , \24296 );
xor \U$23921 ( \24298 , \23417 , \23419 );
xor \U$23922 ( \24299 , \24298 , \23422 );
xor \U$23923 ( \24300 , \23966 , \23971 );
xor \U$23924 ( \24301 , \24299 , \24300 );
xor \U$23925 ( \24302 , \23729 , \23731 );
xor \U$23926 ( \24303 , \24302 , \23744 );
and \U$23927 ( \24304 , \24301 , \24303 );
and \U$23928 ( \24305 , \24294 , \24301 );
or \U$23929 ( \24306 , \24297 , \24304 , \24305 );
and \U$23930 ( \24307 , \24292 , \24306 );
and \U$23931 ( \24308 , \24271 , \24291 );
or \U$23932 ( \24309 , \24307 , \24308 );
xor \U$23933 ( \24310 , \23981 , \23983 );
xor \U$23934 ( \24311 , \23995 , \23997 );
xor \U$23935 ( \24312 , \24311 , \24002 );
and \U$23936 ( \24313 , \24310 , \24312 );
xor \U$23937 ( \24314 , \23747 , \23963 );
xor \U$23938 ( \24315 , \24314 , \23976 );
xor \U$23939 ( \24316 , \23995 , \23997 );
xor \U$23940 ( \24317 , \24316 , \24002 );
and \U$23941 ( \24318 , \24315 , \24317 );
and \U$23942 ( \24319 , \24310 , \24315 );
or \U$23943 ( \24320 , \24313 , \24318 , \24319 );
xor \U$23944 ( \24321 , \24309 , \24320 );
xor \U$23945 ( \24322 , \23382 , \23384 );
xor \U$23946 ( \24323 , \24322 , \23389 );
xor \U$23947 ( \24324 , \23696 , \23701 );
xor \U$23948 ( \24325 , \24323 , \24324 );
and \U$23949 ( \24326 , \24321 , \24325 );
and \U$23950 ( \24327 , \24309 , \24320 );
or \U$23951 ( \24328 , \24326 , \24327 );
not \U$23952 ( \24329 , \24328 );
or \U$23953 ( \24330 , \24026 , \24329 );
or \U$23954 ( \24331 , \24328 , \24025 );
nand \U$23955 ( \24332 , \24330 , \24331 );
not \U$23956 ( \24333 , \24332 );
xnor \U$23957 ( \24334 , \24008 , \23706 );
not \U$23958 ( \24335 , \24334 );
not \U$23959 ( \24336 , \23711 );
and \U$23960 ( \24337 , \24335 , \24336 );
and \U$23961 ( \24338 , \24334 , \23711 );
nor \U$23962 ( \24339 , \24337 , \24338 );
not \U$23963 ( \24340 , \24339 );
and \U$23964 ( \24341 , \24333 , \24340 );
and \U$23965 ( \24342 , \24332 , \24339 );
nor \U$23966 ( \24343 , \24341 , \24342 );
xor \U$23967 ( \24344 , \24309 , \24320 );
xor \U$23968 ( \24345 , \24344 , \24325 );
xor \U$23969 ( \24346 , \24038 , \24040 );
xor \U$23970 ( \24347 , \24346 , \24051 );
xor \U$23971 ( \24348 , \24278 , \24280 );
xor \U$23972 ( \24349 , \24348 , \24283 );
and \U$23973 ( \24350 , \24347 , \24349 );
xor \U$23974 ( \24351 , \23716 , \23723 );
xor \U$23975 ( \24352 , \24351 , \23726 );
xor \U$23976 ( \24353 , \24256 , \24263 );
xor \U$23977 ( \24354 , \24352 , \24353 );
xor \U$23978 ( \24355 , \24278 , \24280 );
xor \U$23979 ( \24356 , \24355 , \24283 );
and \U$23980 ( \24357 , \24354 , \24356 );
and \U$23981 ( \24358 , \24347 , \24354 );
or \U$23982 ( \24359 , \24350 , \24357 , \24358 );
xor \U$23983 ( \24360 , \24112 , \24119 );
xor \U$23984 ( \24361 , \24360 , \24127 );
xor \U$23985 ( \24362 , \24191 , \24198 );
xor \U$23986 ( \24363 , \24362 , \24206 );
and \U$23987 ( \24364 , \24361 , \24363 );
xor \U$23988 ( \24365 , \24140 , \24147 );
xor \U$23989 ( \24366 , \24365 , \24155 );
xor \U$23990 ( \24367 , \24191 , \24198 );
xor \U$23991 ( \24368 , \24367 , \24206 );
and \U$23992 ( \24369 , \24366 , \24368 );
and \U$23993 ( \24370 , \24361 , \24366 );
or \U$23994 ( \24371 , \24364 , \24369 , \24370 );
xor \U$23995 ( \24372 , \24061 , \24068 );
xor \U$23996 ( \24373 , \24372 , \24076 );
xor \U$23997 ( \24374 , \24220 , \24228 );
xor \U$23998 ( \24375 , \24374 , \24237 );
xor \U$23999 ( \24376 , \24373 , \24375 );
xor \U$24000 ( \24377 , \24086 , \24093 );
xor \U$24001 ( \24378 , \24377 , \24101 );
and \U$24002 ( \24379 , \24376 , \24378 );
and \U$24003 ( \24380 , \24373 , \24375 );
or \U$24004 ( \24381 , \24379 , \24380 );
xor \U$24005 ( \24382 , \24371 , \24381 );
xor \U$24006 ( \24383 , \23779 , \1734 );
xor \U$24007 ( \24384 , \24383 , \23787 );
xor \U$24008 ( \24385 , \24028 , \24033 );
xor \U$24009 ( \24386 , \24384 , \24385 );
and \U$24010 ( \24387 , \24382 , \24386 );
and \U$24011 ( \24388 , \24371 , \24381 );
or \U$24012 ( \24389 , \24387 , \24388 );
and \U$24013 ( \24390 , \14059 , RIae75e48_29);
and \U$24014 ( \24391 , RIae75c68_25, \14057 );
nor \U$24015 ( \24392 , \24390 , \24391 );
and \U$24016 ( \24393 , \24392 , \13502 );
not \U$24017 ( \24394 , \24392 );
and \U$24018 ( \24395 , \24394 , \14063 );
nor \U$24019 ( \24396 , \24393 , \24395 );
and \U$24020 ( \24397 , \12180 , RIae75a88_21);
and \U$24021 ( \24398 , RIae75998_19, \12178 );
nor \U$24022 ( \24399 , \24397 , \24398 );
and \U$24023 ( \24400 , \24399 , \12184 );
not \U$24024 ( \24401 , \24399 );
and \U$24025 ( \24402 , \24401 , \11827 );
nor \U$24026 ( \24403 , \24400 , \24402 );
xor \U$24027 ( \24404 , \24396 , \24403 );
and \U$24028 ( \24405 , \13059 , RIae758a8_17);
and \U$24029 ( \24406 , RIae75f38_31, \13057 );
nor \U$24030 ( \24407 , \24405 , \24406 );
and \U$24031 ( \24408 , \24407 , \13063 );
not \U$24032 ( \24409 , \24407 );
and \U$24033 ( \24410 , \24409 , \12718 );
nor \U$24034 ( \24411 , \24408 , \24410 );
and \U$24035 ( \24412 , \24404 , \24411 );
and \U$24036 ( \24413 , \24396 , \24403 );
or \U$24037 ( \24414 , \24412 , \24413 );
and \U$24038 ( \24415 , \15726 , RIae754e8_9);
and \U$24039 ( \24416 , RIae7aab0_192, RIae757b8_15);
nor \U$24040 ( \24417 , \24415 , \24416 );
and \U$24041 ( \24418 , \24417 , \14959 );
not \U$24042 ( \24419 , \24417 );
and \U$24043 ( \24420 , \24419 , RIae7aa38_191);
nor \U$24044 ( \24421 , \24418 , \24420 );
xor \U$24045 ( \24422 , \24421 , \2060 );
and \U$24046 ( \24423 , \14964 , RIae75d58_27);
and \U$24047 ( \24424 , RIae755d8_11, \14962 );
nor \U$24048 ( \24425 , \24423 , \24424 );
and \U$24049 ( \24426 , \24425 , \14463 );
not \U$24050 ( \24427 , \24425 );
and \U$24051 ( \24428 , \24427 , \14462 );
nor \U$24052 ( \24429 , \24426 , \24428 );
and \U$24053 ( \24430 , \24422 , \24429 );
and \U$24054 ( \24431 , \24421 , \2060 );
or \U$24055 ( \24432 , \24430 , \24431 );
xor \U$24056 ( \24433 , \24414 , \24432 );
and \U$24057 ( \24434 , \9760 , RIae77e28_97);
and \U$24058 ( \24435 , RIae78968_121, \9758 );
nor \U$24059 ( \24436 , \24434 , \24435 );
and \U$24060 ( \24437 , \24436 , \9273 );
not \U$24061 ( \24438 , \24436 );
and \U$24062 ( \24439 , \24438 , \9272 );
nor \U$24063 ( \24440 , \24437 , \24439 );
and \U$24064 ( \24441 , \10548 , RIae78878_119);
and \U$24065 ( \24442 , RIae78788_117, \10546 );
nor \U$24066 ( \24443 , \24441 , \24442 );
and \U$24067 ( \24444 , \24443 , \10421 );
not \U$24068 ( \24445 , \24443 );
and \U$24069 ( \24446 , \24445 , \10118 );
nor \U$24070 ( \24447 , \24444 , \24446 );
xor \U$24071 ( \24448 , \24440 , \24447 );
and \U$24072 ( \24449 , \11470 , RIae78698_115);
and \U$24073 ( \24450 , RIae75b78_23, \11468 );
nor \U$24074 ( \24451 , \24449 , \24450 );
and \U$24075 ( \24452 , \24451 , \10936 );
not \U$24076 ( \24453 , \24451 );
and \U$24077 ( \24454 , \24453 , \11474 );
nor \U$24078 ( \24455 , \24452 , \24454 );
and \U$24079 ( \24456 , \24448 , \24455 );
and \U$24080 ( \24457 , \24440 , \24447 );
or \U$24081 ( \24458 , \24456 , \24457 );
and \U$24082 ( \24459 , \24433 , \24458 );
and \U$24083 ( \24460 , \24414 , \24432 );
or \U$24084 ( \24461 , \24459 , \24460 );
nand \U$24085 ( \24462 , RIae775b8_79, \2222 );
and \U$24086 ( \24463 , \24462 , \2061 );
not \U$24087 ( \24464 , \24462 );
and \U$24088 ( \24465 , \24464 , \2060 );
nor \U$24089 ( \24466 , \24463 , \24465 );
and \U$24090 ( \24467 , \2607 , RIae774c8_77);
and \U$24091 ( \24468 , RIae77720_82, \2605 );
nor \U$24092 ( \24469 , \24467 , \24468 );
and \U$24093 ( \24470 , \24469 , \2611 );
not \U$24094 ( \24471 , \24469 );
and \U$24095 ( \24472 , \24471 , \2397 );
nor \U$24096 ( \24473 , \24470 , \24472 );
and \U$24097 ( \24474 , \24466 , \24473 );
and \U$24098 ( \24475 , \2224 , RIae775b8_79);
and \U$24099 ( \24476 , RIae774c8_77, \2222 );
nor \U$24100 ( \24477 , \24475 , \24476 );
and \U$24101 ( \24478 , \24477 , \2061 );
not \U$24102 ( \24479 , \24477 );
and \U$24103 ( \24480 , \24479 , \2060 );
nor \U$24104 ( \24481 , \24478 , \24480 );
xor \U$24105 ( \24482 , \24474 , \24481 );
not \U$24106 ( \24483 , \3089 );
and \U$24107 ( \24484 , \2783 , RIae773d8_75);
and \U$24108 ( \24485 , RIae77a68_89, \2781 );
nor \U$24109 ( \24486 , \24484 , \24485 );
not \U$24110 ( \24487 , \24486 );
or \U$24111 ( \24488 , \24483 , \24487 );
or \U$24112 ( \24489 , \24486 , \2789 );
nand \U$24113 ( \24490 , \24488 , \24489 );
not \U$24114 ( \24491 , \3218 );
and \U$24115 ( \24492 , \3214 , RIae77978_87);
and \U$24116 ( \24493 , RIae77798_83, \3212 );
nor \U$24117 ( \24494 , \24492 , \24493 );
not \U$24118 ( \24495 , \24494 );
or \U$24119 ( \24496 , \24491 , \24495 );
or \U$24120 ( \24497 , \24494 , \3218 );
nand \U$24121 ( \24498 , \24496 , \24497 );
xor \U$24122 ( \24499 , \24490 , \24498 );
and \U$24123 ( \24500 , \3730 , RIae77888_85);
and \U$24124 ( \24501 , RIae76f28_65, \3728 );
nor \U$24125 ( \24502 , \24500 , \24501 );
and \U$24126 ( \24503 , \24502 , \3732 );
not \U$24127 ( \24504 , \24502 );
and \U$24128 ( \24505 , \24504 , \3422 );
nor \U$24129 ( \24506 , \24503 , \24505 );
and \U$24130 ( \24507 , \24499 , \24506 );
and \U$24131 ( \24508 , \24490 , \24498 );
or \U$24132 ( \24509 , \24507 , \24508 );
and \U$24133 ( \24510 , \24482 , \24509 );
and \U$24134 ( \24511 , \24474 , \24481 );
or \U$24135 ( \24512 , \24510 , \24511 );
xor \U$24136 ( \24513 , \24461 , \24512 );
and \U$24137 ( \24514 , \7633 , RIae785a8_113);
and \U$24138 ( \24515 , RIae783c8_109, \7631 );
nor \U$24139 ( \24516 , \24514 , \24515 );
and \U$24140 ( \24517 , \24516 , \7206 );
not \U$24141 ( \24518 , \24516 );
and \U$24142 ( \24519 , \24518 , \7205 );
nor \U$24143 ( \24520 , \24517 , \24519 );
and \U$24144 ( \24521 , \8371 , RIae78530_112);
and \U$24145 ( \24522 , RIae77c48_93, \8369 );
nor \U$24146 ( \24523 , \24521 , \24522 );
and \U$24147 ( \24524 , \24523 , \8020 );
not \U$24148 ( \24525 , \24523 );
and \U$24149 ( \24526 , \24525 , \8019 );
nor \U$24150 ( \24527 , \24524 , \24526 );
xor \U$24151 ( \24528 , \24520 , \24527 );
and \U$24152 ( \24529 , \8966 , RIae77b58_91);
and \U$24153 ( \24530 , RIae77d38_95, \8964 );
nor \U$24154 ( \24531 , \24529 , \24530 );
and \U$24155 ( \24532 , \24531 , \8799 );
not \U$24156 ( \24533 , \24531 );
and \U$24157 ( \24534 , \24533 , \8789 );
nor \U$24158 ( \24535 , \24532 , \24534 );
and \U$24159 ( \24536 , \24528 , \24535 );
and \U$24160 ( \24537 , \24520 , \24527 );
or \U$24161 ( \24538 , \24536 , \24537 );
and \U$24162 ( \24539 , \4247 , RIae76e38_63);
and \U$24163 ( \24540 , RIae76d48_61, \4245 );
nor \U$24164 ( \24541 , \24539 , \24540 );
and \U$24165 ( \24542 , \24541 , \3989 );
not \U$24166 ( \24543 , \24541 );
and \U$24167 ( \24544 , \24543 , \4251 );
nor \U$24168 ( \24545 , \24542 , \24544 );
and \U$24169 ( \24546 , \4688 , RIae76c58_59);
and \U$24170 ( \24547 , RIae77180_70, \4686 );
nor \U$24171 ( \24548 , \24546 , \24547 );
and \U$24172 ( \24549 , \24548 , \4481 );
not \U$24173 ( \24550 , \24548 );
and \U$24174 ( \24551 , \24550 , \4482 );
nor \U$24175 ( \24552 , \24549 , \24551 );
xor \U$24176 ( \24553 , \24545 , \24552 );
and \U$24177 ( \24554 , \5399 , RIae77018_67);
and \U$24178 ( \24555 , RIae771f8_71, \5397 );
nor \U$24179 ( \24556 , \24554 , \24555 );
and \U$24180 ( \24557 , \24556 , \5016 );
not \U$24181 ( \24558 , \24556 );
and \U$24182 ( \24559 , \24558 , \5403 );
nor \U$24183 ( \24560 , \24557 , \24559 );
and \U$24184 ( \24561 , \24553 , \24560 );
and \U$24185 ( \24562 , \24545 , \24552 );
or \U$24186 ( \24563 , \24561 , \24562 );
xor \U$24187 ( \24564 , \24538 , \24563 );
and \U$24188 ( \24565 , \6172 , RIae780f8_103);
and \U$24189 ( \24566 , RIae77f18_99, \6170 );
nor \U$24190 ( \24567 , \24565 , \24566 );
and \U$24191 ( \24568 , \24567 , \6176 );
not \U$24192 ( \24569 , \24567 );
and \U$24193 ( \24570 , \24569 , \6175 );
nor \U$24194 ( \24571 , \24568 , \24570 );
and \U$24195 ( \24572 , \5896 , RIae772e8_73);
and \U$24196 ( \24573 , RIae782d8_107, \5894 );
nor \U$24197 ( \24574 , \24572 , \24573 );
and \U$24198 ( \24575 , \24574 , \5590 );
not \U$24199 ( \24576 , \24574 );
and \U$24200 ( \24577 , \24576 , \5589 );
nor \U$24201 ( \24578 , \24575 , \24577 );
xor \U$24202 ( \24579 , \24571 , \24578 );
and \U$24203 ( \24580 , \6941 , RIae78008_101);
and \U$24204 ( \24581 , RIae781e8_105, \6939 );
nor \U$24205 ( \24582 , \24580 , \24581 );
and \U$24206 ( \24583 , \24582 , \6314 );
not \U$24207 ( \24584 , \24582 );
and \U$24208 ( \24585 , \24584 , \6945 );
nor \U$24209 ( \24586 , \24583 , \24585 );
and \U$24210 ( \24587 , \24579 , \24586 );
and \U$24211 ( \24588 , \24571 , \24578 );
or \U$24212 ( \24589 , \24587 , \24588 );
and \U$24213 ( \24590 , \24564 , \24589 );
and \U$24214 ( \24591 , \24538 , \24563 );
or \U$24215 ( \24592 , \24590 , \24591 );
and \U$24216 ( \24593 , \24513 , \24592 );
and \U$24217 ( \24594 , \24461 , \24512 );
or \U$24218 ( \24595 , \24593 , \24594 );
xor \U$24219 ( \24596 , \24389 , \24595 );
xor \U$24220 ( \24597 , \24079 , \24104 );
xor \U$24221 ( \24598 , \24597 , \24130 );
xor \U$24222 ( \24599 , \24043 , \24045 );
xor \U$24223 ( \24600 , \24599 , \24048 );
and \U$24224 ( \24601 , \24598 , \24600 );
xor \U$24225 ( \24602 , \23858 , \23866 );
xor \U$24226 ( \24603 , \24602 , \23874 );
xor \U$24227 ( \24604 , \24240 , \24245 );
xor \U$24228 ( \24605 , \24603 , \24604 );
xor \U$24229 ( \24606 , \24043 , \24045 );
xor \U$24230 ( \24607 , \24606 , \24048 );
and \U$24231 ( \24608 , \24605 , \24607 );
and \U$24232 ( \24609 , \24598 , \24605 );
or \U$24233 ( \24610 , \24601 , \24608 , \24609 );
and \U$24234 ( \24611 , \24596 , \24610 );
and \U$24235 ( \24612 , \24389 , \24595 );
or \U$24236 ( \24613 , \24611 , \24612 );
xor \U$24237 ( \24614 , \24359 , \24613 );
xor \U$24238 ( \24615 , \23729 , \23731 );
xor \U$24239 ( \24616 , \24615 , \23744 );
xor \U$24240 ( \24617 , \24294 , \24301 );
xor \U$24241 ( \24618 , \24616 , \24617 );
and \U$24242 ( \24619 , \24614 , \24618 );
and \U$24243 ( \24620 , \24359 , \24613 );
or \U$24244 ( \24621 , \24619 , \24620 );
xor \U$24245 ( \24622 , \24271 , \24291 );
xor \U$24246 ( \24623 , \24622 , \24306 );
xor \U$24247 ( \24624 , \24621 , \24623 );
xor \U$24248 ( \24625 , \23995 , \23997 );
xor \U$24249 ( \24626 , \24625 , \24002 );
xor \U$24250 ( \24627 , \24310 , \24315 );
xor \U$24251 ( \24628 , \24626 , \24627 );
and \U$24252 ( \24629 , \24624 , \24628 );
and \U$24253 ( \24630 , \24621 , \24623 );
or \U$24254 ( \24631 , \24629 , \24630 );
xor \U$24255 ( \24632 , \24345 , \24631 );
xor \U$24256 ( \24633 , \23979 , \23984 );
xor \U$24257 ( \24634 , \24633 , \24005 );
and \U$24258 ( \24635 , \24632 , \24634 );
and \U$24259 ( \24636 , \24345 , \24631 );
nor \U$24260 ( \24637 , \24635 , \24636 );
or \U$24261 ( \24638 , \24343 , \24637 );
xnor \U$24262 ( \24639 , \24343 , \24637 );
xor \U$24263 ( \24640 , \24054 , \24253 );
xor \U$24264 ( \24641 , \24640 , \24268 );
xor \U$24265 ( \24642 , \24359 , \24613 );
xor \U$24266 ( \24643 , \24642 , \24618 );
xor \U$24267 ( \24644 , \24641 , \24643 );
xor \U$24268 ( \24645 , \24389 , \24595 );
xor \U$24269 ( \24646 , \24645 , \24610 );
xor \U$24270 ( \24647 , \24278 , \24280 );
xor \U$24271 ( \24648 , \24647 , \24283 );
xor \U$24272 ( \24649 , \24347 , \24354 );
xor \U$24273 ( \24650 , \24648 , \24649 );
xor \U$24274 ( \24651 , \24646 , \24650 );
xor \U$24275 ( \24652 , \24538 , \24563 );
xor \U$24276 ( \24653 , \24652 , \24589 );
xor \U$24277 ( \24654 , \24414 , \24432 );
xor \U$24278 ( \24655 , \24654 , \24458 );
xor \U$24279 ( \24656 , \24653 , \24655 );
xor \U$24280 ( \24657 , \24373 , \24375 );
xor \U$24281 ( \24658 , \24657 , \24378 );
xor \U$24282 ( \24659 , \24474 , \24481 );
xor \U$24283 ( \24660 , \24659 , \24509 );
xor \U$24284 ( \24661 , \24191 , \24198 );
xor \U$24285 ( \24662 , \24661 , \24206 );
xor \U$24286 ( \24663 , \24361 , \24366 );
xor \U$24287 ( \24664 , \24662 , \24663 );
xor \U$24288 ( \24665 , \24660 , \24664 );
xor \U$24289 ( \24666 , \24658 , \24665 );
and \U$24290 ( \24667 , \24656 , \24666 );
and \U$24291 ( \24668 , \24653 , \24655 );
or \U$24292 ( \24669 , \24667 , \24668 );
xor \U$24293 ( \24670 , \24461 , \24512 );
xor \U$24294 ( \24671 , \24670 , \24592 );
xor \U$24295 ( \24672 , \24669 , \24671 );
and \U$24296 ( \24673 , \5896 , RIae771f8_71);
and \U$24297 ( \24674 , RIae772e8_73, \5894 );
nor \U$24298 ( \24675 , \24673 , \24674 );
and \U$24299 ( \24676 , \24675 , \5590 );
not \U$24300 ( \24677 , \24675 );
and \U$24301 ( \24678 , \24677 , \5589 );
nor \U$24302 ( \24679 , \24676 , \24678 );
and \U$24303 ( \24680 , \5399 , RIae77180_70);
and \U$24304 ( \24681 , RIae77018_67, \5397 );
nor \U$24305 ( \24682 , \24680 , \24681 );
and \U$24306 ( \24683 , \24682 , \5016 );
not \U$24307 ( \24684 , \24682 );
and \U$24308 ( \24685 , \24684 , \5403 );
nor \U$24309 ( \24686 , \24683 , \24685 );
xor \U$24310 ( \24687 , \24679 , \24686 );
and \U$24311 ( \24688 , \6172 , RIae782d8_107);
and \U$24312 ( \24689 , RIae780f8_103, \6170 );
nor \U$24313 ( \24690 , \24688 , \24689 );
and \U$24314 ( \24691 , \24690 , \6176 );
not \U$24315 ( \24692 , \24690 );
and \U$24316 ( \24693 , \24692 , \6175 );
nor \U$24317 ( \24694 , \24691 , \24693 );
and \U$24318 ( \24695 , \24687 , \24694 );
and \U$24319 ( \24696 , \24679 , \24686 );
or \U$24320 ( \24697 , \24695 , \24696 );
and \U$24321 ( \24698 , \4247 , RIae76f28_65);
and \U$24322 ( \24699 , RIae76e38_63, \4245 );
nor \U$24323 ( \24700 , \24698 , \24699 );
and \U$24324 ( \24701 , \24700 , \3989 );
not \U$24325 ( \24702 , \24700 );
and \U$24326 ( \24703 , \24702 , \4251 );
nor \U$24327 ( \24704 , \24701 , \24703 );
and \U$24328 ( \24705 , \3730 , RIae77798_83);
and \U$24329 ( \24706 , RIae77888_85, \3728 );
nor \U$24330 ( \24707 , \24705 , \24706 );
and \U$24331 ( \24708 , \24707 , \3732 );
not \U$24332 ( \24709 , \24707 );
and \U$24333 ( \24710 , \24709 , \3422 );
nor \U$24334 ( \24711 , \24708 , \24710 );
xor \U$24335 ( \24712 , \24704 , \24711 );
and \U$24336 ( \24713 , \4688 , RIae76d48_61);
and \U$24337 ( \24714 , RIae76c58_59, \4686 );
nor \U$24338 ( \24715 , \24713 , \24714 );
and \U$24339 ( \24716 , \24715 , \4481 );
not \U$24340 ( \24717 , \24715 );
and \U$24341 ( \24718 , \24717 , \4482 );
nor \U$24342 ( \24719 , \24716 , \24718 );
and \U$24343 ( \24720 , \24712 , \24719 );
and \U$24344 ( \24721 , \24704 , \24711 );
or \U$24345 ( \24722 , \24720 , \24721 );
xor \U$24346 ( \24723 , \24697 , \24722 );
and \U$24347 ( \24724 , \6941 , RIae77f18_99);
and \U$24348 ( \24725 , RIae78008_101, \6939 );
nor \U$24349 ( \24726 , \24724 , \24725 );
and \U$24350 ( \24727 , \24726 , \6314 );
not \U$24351 ( \24728 , \24726 );
and \U$24352 ( \24729 , \24728 , \6945 );
nor \U$24353 ( \24730 , \24727 , \24729 );
and \U$24354 ( \24731 , \7633 , RIae781e8_105);
and \U$24355 ( \24732 , RIae785a8_113, \7631 );
nor \U$24356 ( \24733 , \24731 , \24732 );
and \U$24357 ( \24734 , \24733 , \7206 );
not \U$24358 ( \24735 , \24733 );
and \U$24359 ( \24736 , \24735 , \7205 );
nor \U$24360 ( \24737 , \24734 , \24736 );
xor \U$24361 ( \24738 , \24730 , \24737 );
and \U$24362 ( \24739 , \8371 , RIae783c8_109);
and \U$24363 ( \24740 , RIae78530_112, \8369 );
nor \U$24364 ( \24741 , \24739 , \24740 );
and \U$24365 ( \24742 , \24741 , \8020 );
not \U$24366 ( \24743 , \24741 );
and \U$24367 ( \24744 , \24743 , \8019 );
nor \U$24368 ( \24745 , \24742 , \24744 );
and \U$24369 ( \24746 , \24738 , \24745 );
and \U$24370 ( \24747 , \24730 , \24737 );
or \U$24371 ( \24748 , \24746 , \24747 );
xor \U$24372 ( \24749 , \24723 , \24748 );
xor \U$24373 ( \24750 , \24571 , \24578 );
xor \U$24374 ( \24751 , \24750 , \24586 );
xor \U$24375 ( \24752 , \24545 , \24552 );
xor \U$24376 ( \24753 , \24752 , \24560 );
xor \U$24377 ( \24754 , \24751 , \24753 );
xor \U$24378 ( \24755 , \24520 , \24527 );
xor \U$24379 ( \24756 , \24755 , \24535 );
xor \U$24380 ( \24757 , \24754 , \24756 );
and \U$24381 ( \24758 , \24749 , \24757 );
and \U$24382 ( \24759 , \2607 , RIae775b8_79);
and \U$24383 ( \24760 , RIae774c8_77, \2605 );
nor \U$24384 ( \24761 , \24759 , \24760 );
and \U$24385 ( \24762 , \24761 , \2611 );
not \U$24386 ( \24763 , \24761 );
and \U$24387 ( \24764 , \24763 , \2397 );
nor \U$24388 ( \24765 , \24762 , \24764 );
not \U$24389 ( \24766 , \2789 );
and \U$24390 ( \24767 , \2783 , RIae77720_82);
and \U$24391 ( \24768 , RIae773d8_75, \2781 );
nor \U$24392 ( \24769 , \24767 , \24768 );
not \U$24393 ( \24770 , \24769 );
or \U$24394 ( \24771 , \24766 , \24770 );
or \U$24395 ( \24772 , \24769 , \2789 );
nand \U$24396 ( \24773 , \24771 , \24772 );
xor \U$24397 ( \24774 , \24765 , \24773 );
not \U$24398 ( \24775 , \2774 );
and \U$24399 ( \24776 , \3214 , RIae77a68_89);
and \U$24400 ( \24777 , RIae77978_87, \3212 );
nor \U$24401 ( \24778 , \24776 , \24777 );
not \U$24402 ( \24779 , \24778 );
or \U$24403 ( \24780 , \24775 , \24779 );
or \U$24404 ( \24781 , \24778 , \3218 );
nand \U$24405 ( \24782 , \24780 , \24781 );
and \U$24406 ( \24783 , \24774 , \24782 );
and \U$24407 ( \24784 , \24765 , \24773 );
or \U$24408 ( \24785 , \24783 , \24784 );
xor \U$24409 ( \24786 , \24466 , \24473 );
xor \U$24410 ( \24787 , \24785 , \24786 );
xor \U$24411 ( \24788 , \24490 , \24498 );
xor \U$24412 ( \24789 , \24788 , \24506 );
xor \U$24413 ( \24790 , \24787 , \24789 );
xor \U$24414 ( \24791 , \24751 , \24753 );
xor \U$24415 ( \24792 , \24791 , \24756 );
and \U$24416 ( \24793 , \24790 , \24792 );
and \U$24417 ( \24794 , \24749 , \24790 );
or \U$24418 ( \24795 , \24758 , \24793 , \24794 );
and \U$24419 ( \24796 , \7633 , RIae78008_101);
and \U$24420 ( \24797 , RIae781e8_105, \7631 );
nor \U$24421 ( \24798 , \24796 , \24797 );
and \U$24422 ( \24799 , \24798 , \7206 );
not \U$24423 ( \24800 , \24798 );
and \U$24424 ( \24801 , \24800 , \7205 );
nor \U$24425 ( \24802 , \24799 , \24801 );
and \U$24426 ( \24803 , \8371 , RIae785a8_113);
and \U$24427 ( \24804 , RIae783c8_109, \8369 );
nor \U$24428 ( \24805 , \24803 , \24804 );
and \U$24429 ( \24806 , \24805 , \8020 );
not \U$24430 ( \24807 , \24805 );
and \U$24431 ( \24808 , \24807 , \8019 );
nor \U$24432 ( \24809 , \24806 , \24808 );
xor \U$24433 ( \24810 , \24802 , \24809 );
and \U$24434 ( \24811 , \8966 , RIae78530_112);
and \U$24435 ( \24812 , RIae77c48_93, \8964 );
nor \U$24436 ( \24813 , \24811 , \24812 );
and \U$24437 ( \24814 , \24813 , \8799 );
not \U$24438 ( \24815 , \24813 );
and \U$24439 ( \24816 , \24815 , \8789 );
nor \U$24440 ( \24817 , \24814 , \24816 );
and \U$24441 ( \24818 , \24810 , \24817 );
and \U$24442 ( \24819 , \24802 , \24809 );
or \U$24443 ( \24820 , \24818 , \24819 );
and \U$24444 ( \24821 , \4247 , RIae77888_85);
and \U$24445 ( \24822 , RIae76f28_65, \4245 );
nor \U$24446 ( \24823 , \24821 , \24822 );
and \U$24447 ( \24824 , \24823 , \3989 );
not \U$24448 ( \24825 , \24823 );
and \U$24449 ( \24826 , \24825 , \4251 );
nor \U$24450 ( \24827 , \24824 , \24826 );
and \U$24451 ( \24828 , \4688 , RIae76e38_63);
and \U$24452 ( \24829 , RIae76d48_61, \4686 );
nor \U$24453 ( \24830 , \24828 , \24829 );
and \U$24454 ( \24831 , \24830 , \4481 );
not \U$24455 ( \24832 , \24830 );
and \U$24456 ( \24833 , \24832 , \4482 );
nor \U$24457 ( \24834 , \24831 , \24833 );
xor \U$24458 ( \24835 , \24827 , \24834 );
and \U$24459 ( \24836 , \5399 , RIae76c58_59);
and \U$24460 ( \24837 , RIae77180_70, \5397 );
nor \U$24461 ( \24838 , \24836 , \24837 );
and \U$24462 ( \24839 , \24838 , \5016 );
not \U$24463 ( \24840 , \24838 );
and \U$24464 ( \24841 , \24840 , \5403 );
nor \U$24465 ( \24842 , \24839 , \24841 );
and \U$24466 ( \24843 , \24835 , \24842 );
and \U$24467 ( \24844 , \24827 , \24834 );
or \U$24468 ( \24845 , \24843 , \24844 );
xor \U$24469 ( \24846 , \24820 , \24845 );
and \U$24470 ( \24847 , \6172 , RIae772e8_73);
and \U$24471 ( \24848 , RIae782d8_107, \6170 );
nor \U$24472 ( \24849 , \24847 , \24848 );
and \U$24473 ( \24850 , \24849 , \6176 );
not \U$24474 ( \24851 , \24849 );
and \U$24475 ( \24852 , \24851 , \6175 );
nor \U$24476 ( \24853 , \24850 , \24852 );
and \U$24477 ( \24854 , \5896 , RIae77018_67);
and \U$24478 ( \24855 , RIae771f8_71, \5894 );
nor \U$24479 ( \24856 , \24854 , \24855 );
and \U$24480 ( \24857 , \24856 , \5590 );
not \U$24481 ( \24858 , \24856 );
and \U$24482 ( \24859 , \24858 , \5589 );
nor \U$24483 ( \24860 , \24857 , \24859 );
xor \U$24484 ( \24861 , \24853 , \24860 );
and \U$24485 ( \24862 , \6941 , RIae780f8_103);
and \U$24486 ( \24863 , RIae77f18_99, \6939 );
nor \U$24487 ( \24864 , \24862 , \24863 );
and \U$24488 ( \24865 , \24864 , \6314 );
not \U$24489 ( \24866 , \24864 );
and \U$24490 ( \24867 , \24866 , \6945 );
nor \U$24491 ( \24868 , \24865 , \24867 );
and \U$24492 ( \24869 , \24861 , \24868 );
and \U$24493 ( \24870 , \24853 , \24860 );
or \U$24494 ( \24871 , \24869 , \24870 );
and \U$24495 ( \24872 , \24846 , \24871 );
and \U$24496 ( \24873 , \24820 , \24845 );
or \U$24497 ( \24874 , \24872 , \24873 );
and \U$24498 ( \24875 , \10548 , RIae77e28_97);
and \U$24499 ( \24876 , RIae78968_121, \10546 );
nor \U$24500 ( \24877 , \24875 , \24876 );
and \U$24501 ( \24878 , \24877 , \10421 );
not \U$24502 ( \24879 , \24877 );
and \U$24503 ( \24880 , \24879 , \10118 );
nor \U$24504 ( \24881 , \24878 , \24880 );
and \U$24505 ( \24882 , \9760 , RIae77b58_91);
and \U$24506 ( \24883 , RIae77d38_95, \9758 );
nor \U$24507 ( \24884 , \24882 , \24883 );
and \U$24508 ( \24885 , \24884 , \9273 );
not \U$24509 ( \24886 , \24884 );
and \U$24510 ( \24887 , \24886 , \9272 );
nor \U$24511 ( \24888 , \24885 , \24887 );
xor \U$24512 ( \24889 , \24881 , \24888 );
and \U$24513 ( \24890 , \11470 , RIae78878_119);
and \U$24514 ( \24891 , RIae78788_117, \11468 );
nor \U$24515 ( \24892 , \24890 , \24891 );
and \U$24516 ( \24893 , \24892 , \10936 );
not \U$24517 ( \24894 , \24892 );
and \U$24518 ( \24895 , \24894 , \11474 );
nor \U$24519 ( \24896 , \24893 , \24895 );
and \U$24520 ( \24897 , \24889 , \24896 );
and \U$24521 ( \24898 , \24881 , \24888 );
or \U$24522 ( \24899 , \24897 , \24898 );
and \U$24523 ( \24900 , \15726 , RIae75d58_27);
and \U$24524 ( \24901 , RIae7aab0_192, RIae755d8_11);
nor \U$24525 ( \24902 , \24900 , \24901 );
and \U$24526 ( \24903 , \24902 , \14959 );
not \U$24527 ( \24904 , \24902 );
and \U$24528 ( \24905 , \24904 , RIae7aa38_191);
nor \U$24529 ( \24906 , \24903 , \24905 );
xor \U$24530 ( \24907 , \24906 , \2397 );
and \U$24531 ( \24908 , \14964 , RIae75e48_29);
and \U$24532 ( \24909 , RIae75c68_25, \14962 );
nor \U$24533 ( \24910 , \24908 , \24909 );
and \U$24534 ( \24911 , \24910 , \14463 );
not \U$24535 ( \24912 , \24910 );
and \U$24536 ( \24913 , \24912 , \14462 );
nor \U$24537 ( \24914 , \24911 , \24913 );
and \U$24538 ( \24915 , \24907 , \24914 );
and \U$24539 ( \24916 , \24906 , \2397 );
or \U$24540 ( \24917 , \24915 , \24916 );
xor \U$24541 ( \24918 , \24899 , \24917 );
and \U$24542 ( \24919 , \14059 , RIae758a8_17);
and \U$24543 ( \24920 , RIae75f38_31, \14057 );
nor \U$24544 ( \24921 , \24919 , \24920 );
and \U$24545 ( \24922 , \24921 , \13502 );
not \U$24546 ( \24923 , \24921 );
and \U$24547 ( \24924 , \24923 , \14063 );
nor \U$24548 ( \24925 , \24922 , \24924 );
and \U$24549 ( \24926 , \12180 , RIae78698_115);
and \U$24550 ( \24927 , RIae75b78_23, \12178 );
nor \U$24551 ( \24928 , \24926 , \24927 );
and \U$24552 ( \24929 , \24928 , \12184 );
not \U$24553 ( \24930 , \24928 );
and \U$24554 ( \24931 , \24930 , \11827 );
nor \U$24555 ( \24932 , \24929 , \24931 );
xor \U$24556 ( \24933 , \24925 , \24932 );
and \U$24557 ( \24934 , \13059 , RIae75a88_21);
and \U$24558 ( \24935 , RIae75998_19, \13057 );
nor \U$24559 ( \24936 , \24934 , \24935 );
and \U$24560 ( \24937 , \24936 , \13063 );
not \U$24561 ( \24938 , \24936 );
and \U$24562 ( \24939 , \24938 , \12718 );
nor \U$24563 ( \24940 , \24937 , \24939 );
and \U$24564 ( \24941 , \24933 , \24940 );
and \U$24565 ( \24942 , \24925 , \24932 );
or \U$24566 ( \24943 , \24941 , \24942 );
and \U$24567 ( \24944 , \24918 , \24943 );
and \U$24568 ( \24945 , \24899 , \24917 );
or \U$24569 ( \24946 , \24944 , \24945 );
xor \U$24570 ( \24947 , \24874 , \24946 );
and \U$24571 ( \24948 , \3730 , RIae77978_87);
and \U$24572 ( \24949 , RIae77798_83, \3728 );
nor \U$24573 ( \24950 , \24948 , \24949 );
and \U$24574 ( \24951 , \24950 , \3732 );
not \U$24575 ( \24952 , \24950 );
and \U$24576 ( \24953 , \24952 , \3422 );
nor \U$24577 ( \24954 , \24951 , \24953 );
not \U$24578 ( \24955 , \2789 );
and \U$24579 ( \24956 , \2783 , RIae774c8_77);
and \U$24580 ( \24957 , RIae77720_82, \2781 );
nor \U$24581 ( \24958 , \24956 , \24957 );
not \U$24582 ( \24959 , \24958 );
or \U$24583 ( \24960 , \24955 , \24959 );
or \U$24584 ( \24961 , \24958 , \3089 );
nand \U$24585 ( \24962 , \24960 , \24961 );
xor \U$24586 ( \24963 , \24954 , \24962 );
not \U$24587 ( \24964 , \3218 );
and \U$24588 ( \24965 , \3214 , RIae773d8_75);
and \U$24589 ( \24966 , RIae77a68_89, \3212 );
nor \U$24590 ( \24967 , \24965 , \24966 );
not \U$24591 ( \24968 , \24967 );
or \U$24592 ( \24969 , \24964 , \24968 );
or \U$24593 ( \24970 , \24967 , \2774 );
nand \U$24594 ( \24971 , \24969 , \24970 );
and \U$24595 ( \24972 , \24963 , \24971 );
and \U$24596 ( \24973 , \24954 , \24962 );
or \U$24597 ( \24974 , \24972 , \24973 );
xor \U$24598 ( \24975 , \24765 , \24773 );
xor \U$24599 ( \24976 , \24975 , \24782 );
and \U$24600 ( \24977 , \24974 , \24976 );
xor \U$24601 ( \24978 , \24704 , \24711 );
xor \U$24602 ( \24979 , \24978 , \24719 );
xor \U$24603 ( \24980 , \24765 , \24773 );
xor \U$24604 ( \24981 , \24980 , \24782 );
and \U$24605 ( \24982 , \24979 , \24981 );
and \U$24606 ( \24983 , \24974 , \24979 );
or \U$24607 ( \24984 , \24977 , \24982 , \24983 );
and \U$24608 ( \24985 , \24947 , \24984 );
and \U$24609 ( \24986 , \24874 , \24946 );
or \U$24610 ( \24987 , \24985 , \24986 );
xor \U$24611 ( \24988 , \24795 , \24987 );
xor \U$24612 ( \24989 , \24730 , \24737 );
xor \U$24613 ( \24990 , \24989 , \24745 );
xor \U$24614 ( \24991 , \24679 , \24686 );
xor \U$24615 ( \24992 , \24991 , \24694 );
and \U$24616 ( \24993 , \24990 , \24992 );
and \U$24617 ( \24994 , \8966 , RIae77c48_93);
and \U$24618 ( \24995 , RIae77b58_91, \8964 );
nor \U$24619 ( \24996 , \24994 , \24995 );
and \U$24620 ( \24997 , \24996 , \8799 );
not \U$24621 ( \24998 , \24996 );
and \U$24622 ( \24999 , \24998 , \8789 );
nor \U$24623 ( \25000 , \24997 , \24999 );
and \U$24624 ( \25001 , \9760 , RIae77d38_95);
and \U$24625 ( \25002 , RIae77e28_97, \9758 );
nor \U$24626 ( \25003 , \25001 , \25002 );
and \U$24627 ( \25004 , \25003 , \9273 );
not \U$24628 ( \25005 , \25003 );
and \U$24629 ( \25006 , \25005 , \9764 );
nor \U$24630 ( \25007 , \25004 , \25006 );
xor \U$24631 ( \25008 , \25000 , \25007 );
and \U$24632 ( \25009 , \10548 , RIae78968_121);
and \U$24633 ( \25010 , RIae78878_119, \10546 );
nor \U$24634 ( \25011 , \25009 , \25010 );
and \U$24635 ( \25012 , \25011 , \10421 );
not \U$24636 ( \25013 , \25011 );
and \U$24637 ( \25014 , \25013 , \10118 );
nor \U$24638 ( \25015 , \25012 , \25014 );
xor \U$24639 ( \25016 , \25008 , \25015 );
xor \U$24640 ( \25017 , \24679 , \24686 );
xor \U$24641 ( \25018 , \25017 , \24694 );
and \U$24642 ( \25019 , \25016 , \25018 );
and \U$24643 ( \25020 , \24990 , \25016 );
or \U$24644 ( \25021 , \24993 , \25019 , \25020 );
and \U$24645 ( \25022 , \12180 , RIae75b78_23);
and \U$24646 ( \25023 , RIae75a88_21, \12178 );
nor \U$24647 ( \25024 , \25022 , \25023 );
and \U$24648 ( \25025 , \25024 , \12184 );
not \U$24649 ( \25026 , \25024 );
and \U$24650 ( \25027 , \25026 , \11827 );
nor \U$24651 ( \25028 , \25025 , \25027 );
and \U$24652 ( \25029 , \11470 , RIae78788_117);
and \U$24653 ( \25030 , RIae78698_115, \11468 );
nor \U$24654 ( \25031 , \25029 , \25030 );
and \U$24655 ( \25032 , \25031 , \10936 );
not \U$24656 ( \25033 , \25031 );
and \U$24657 ( \25034 , \25033 , \11474 );
nor \U$24658 ( \25035 , \25032 , \25034 );
xor \U$24659 ( \25036 , \25028 , \25035 );
and \U$24660 ( \25037 , \13059 , RIae75998_19);
and \U$24661 ( \25038 , RIae758a8_17, \13057 );
nor \U$24662 ( \25039 , \25037 , \25038 );
and \U$24663 ( \25040 , \25039 , \13063 );
not \U$24664 ( \25041 , \25039 );
and \U$24665 ( \25042 , \25041 , \12718 );
nor \U$24666 ( \25043 , \25040 , \25042 );
xor \U$24667 ( \25044 , \25036 , \25043 );
and \U$24668 ( \25045 , \14059 , RIae75f38_31);
and \U$24669 ( \25046 , RIae75e48_29, \14057 );
nor \U$24670 ( \25047 , \25045 , \25046 );
and \U$24671 ( \25048 , \25047 , \13502 );
not \U$24672 ( \25049 , \25047 );
and \U$24673 ( \25050 , \25049 , \14063 );
nor \U$24674 ( \25051 , \25048 , \25050 );
and \U$24675 ( \25052 , \15726 , RIae755d8_11);
and \U$24676 ( \25053 , RIae7aab0_192, RIae754e8_9);
nor \U$24677 ( \25054 , \25052 , \25053 );
and \U$24678 ( \25055 , \25054 , \14959 );
not \U$24679 ( \25056 , \25054 );
and \U$24680 ( \25057 , \25056 , RIae7aa38_191);
nor \U$24681 ( \25058 , \25055 , \25057 );
xor \U$24682 ( \25059 , \25051 , \25058 );
and \U$24683 ( \25060 , \14964 , RIae75c68_25);
and \U$24684 ( \25061 , RIae75d58_27, \14962 );
nor \U$24685 ( \25062 , \25060 , \25061 );
and \U$24686 ( \25063 , \25062 , \14463 );
not \U$24687 ( \25064 , \25062 );
and \U$24688 ( \25065 , \25064 , \14462 );
nor \U$24689 ( \25066 , \25063 , \25065 );
xor \U$24690 ( \25067 , \25059 , \25066 );
and \U$24691 ( \25068 , \25044 , \25067 );
xor \U$24692 ( \25069 , \25021 , \25068 );
xor \U$24693 ( \25070 , \24440 , \24447 );
xor \U$24694 ( \25071 , \25070 , \24455 );
xor \U$24695 ( \25072 , \24421 , \2060 );
xor \U$24696 ( \25073 , \25072 , \24429 );
xor \U$24697 ( \25074 , \24396 , \24403 );
xor \U$24698 ( \25075 , \25074 , \24411 );
xor \U$24699 ( \25076 , \25073 , \25075 );
xor \U$24700 ( \25077 , \25071 , \25076 );
and \U$24701 ( \25078 , \25069 , \25077 );
and \U$24702 ( \25079 , \25021 , \25068 );
or \U$24703 ( \25080 , \25078 , \25079 );
and \U$24704 ( \25081 , \24988 , \25080 );
and \U$24705 ( \25082 , \24795 , \24987 );
or \U$24706 ( \25083 , \25081 , \25082 );
and \U$24707 ( \25084 , \24672 , \25083 );
and \U$24708 ( \25085 , \24669 , \24671 );
or \U$24709 ( \25086 , \25084 , \25085 );
xor \U$24710 ( \25087 , \24651 , \25086 );
xor \U$24711 ( \25088 , \24440 , \24447 );
xor \U$24712 ( \25089 , \25088 , \24455 );
and \U$24713 ( \25090 , \25073 , \25089 );
xor \U$24714 ( \25091 , \24440 , \24447 );
xor \U$24715 ( \25092 , \25091 , \24455 );
and \U$24716 ( \25093 , \25075 , \25092 );
and \U$24717 ( \25094 , \25073 , \25075 );
or \U$24718 ( \25095 , \25090 , \25093 , \25094 );
xor \U$24719 ( \25096 , \24165 , \24172 );
xor \U$24720 ( \25097 , \25096 , \24180 );
xor \U$24721 ( \25098 , \25095 , \25097 );
xor \U$24722 ( \25099 , \24751 , \24753 );
and \U$24723 ( \25100 , \25099 , \24756 );
and \U$24724 ( \25101 , \24751 , \24753 );
or \U$24725 ( \25102 , \25100 , \25101 );
and \U$24726 ( \25103 , \25098 , \25102 );
and \U$24727 ( \25104 , \25095 , \25097 );
or \U$24728 ( \25105 , \25103 , \25104 );
xor \U$24729 ( \25106 , \24697 , \24722 );
and \U$24730 ( \25107 , \25106 , \24748 );
and \U$24731 ( \25108 , \24697 , \24722 );
or \U$24732 ( \25109 , \25107 , \25108 );
xor \U$24733 ( \25110 , \25000 , \25007 );
and \U$24734 ( \25111 , \25110 , \25015 );
and \U$24735 ( \25112 , \25000 , \25007 );
or \U$24736 ( \25113 , \25111 , \25112 );
xor \U$24737 ( \25114 , \25051 , \25058 );
and \U$24738 ( \25115 , \25114 , \25066 );
and \U$24739 ( \25116 , \25051 , \25058 );
or \U$24740 ( \25117 , \25115 , \25116 );
xor \U$24741 ( \25118 , \25113 , \25117 );
xor \U$24742 ( \25119 , \25028 , \25035 );
and \U$24743 ( \25120 , \25119 , \25043 );
and \U$24744 ( \25121 , \25028 , \25035 );
or \U$24745 ( \25122 , \25120 , \25121 );
and \U$24746 ( \25123 , \25118 , \25122 );
and \U$24747 ( \25124 , \25113 , \25117 );
or \U$24748 ( \25125 , \25123 , \25124 );
xor \U$24749 ( \25126 , \25109 , \25125 );
xor \U$24750 ( \25127 , \24785 , \24786 );
and \U$24751 ( \25128 , \25127 , \24789 );
and \U$24752 ( \25129 , \24785 , \24786 );
or \U$24753 ( \25130 , \25128 , \25129 );
and \U$24754 ( \25131 , \25126 , \25130 );
and \U$24755 ( \25132 , \25109 , \25125 );
or \U$24756 ( \25133 , \25131 , \25132 );
xor \U$24757 ( \25134 , \25105 , \25133 );
xor \U$24758 ( \25135 , \24373 , \24375 );
xor \U$24759 ( \25136 , \25135 , \24378 );
and \U$24760 ( \25137 , \24660 , \25136 );
xor \U$24761 ( \25138 , \24373 , \24375 );
xor \U$24762 ( \25139 , \25138 , \24378 );
and \U$24763 ( \25140 , \24664 , \25139 );
and \U$24764 ( \25141 , \24660 , \24664 );
or \U$24765 ( \25142 , \25137 , \25140 , \25141 );
and \U$24766 ( \25143 , \25134 , \25142 );
and \U$24767 ( \25144 , \25105 , \25133 );
or \U$24768 ( \25145 , \25143 , \25144 );
xor \U$24769 ( \25146 , \24133 , \24212 );
xor \U$24770 ( \25147 , \25146 , \24250 );
xor \U$24771 ( \25148 , \25145 , \25147 );
xor \U$24772 ( \25149 , \24158 , \24183 );
xor \U$24773 ( \25150 , \25149 , \24209 );
xor \U$24774 ( \25151 , \24371 , \24381 );
xor \U$24775 ( \25152 , \25151 , \24386 );
and \U$24776 ( \25153 , \25150 , \25152 );
xor \U$24777 ( \25154 , \24043 , \24045 );
xor \U$24778 ( \25155 , \25154 , \24048 );
xor \U$24779 ( \25156 , \24598 , \24605 );
xor \U$24780 ( \25157 , \25155 , \25156 );
xor \U$24781 ( \25158 , \24371 , \24381 );
xor \U$24782 ( \25159 , \25158 , \24386 );
and \U$24783 ( \25160 , \25157 , \25159 );
and \U$24784 ( \25161 , \25150 , \25157 );
or \U$24785 ( \25162 , \25153 , \25160 , \25161 );
xor \U$24786 ( \25163 , \25148 , \25162 );
and \U$24787 ( \25164 , \25087 , \25163 );
and \U$24788 ( \25165 , \24651 , \25086 );
or \U$24789 ( \25166 , \25164 , \25165 );
xor \U$24790 ( \25167 , \24644 , \25166 );
and \U$24791 ( \25168 , \24646 , \24650 );
xor \U$24792 ( \25169 , \23470 , \23495 );
xor \U$24793 ( \25170 , \25169 , \23521 );
xor \U$24794 ( \25171 , \24273 , \24286 );
xor \U$24795 ( \25172 , \25170 , \25171 );
xor \U$24796 ( \25173 , \25168 , \25172 );
xor \U$24797 ( \25174 , \25145 , \25147 );
and \U$24798 ( \25175 , \25174 , \25162 );
and \U$24799 ( \25176 , \25145 , \25147 );
or \U$24800 ( \25177 , \25175 , \25176 );
xor \U$24801 ( \25178 , \25173 , \25177 );
xor \U$24802 ( \25179 , \25167 , \25178 );
xor \U$24803 ( \25180 , \25105 , \25133 );
xor \U$24804 ( \25181 , \25180 , \25142 );
xor \U$24805 ( \25182 , \24669 , \24671 );
xor \U$24806 ( \25183 , \25182 , \25083 );
and \U$24807 ( \25184 , \25181 , \25183 );
not \U$24808 ( \25185 , \25184 );
xor \U$24809 ( \25186 , \24651 , \25086 );
xor \U$24810 ( \25187 , \25186 , \25163 );
not \U$24811 ( \25188 , \25187 );
or \U$24812 ( \25189 , \25185 , \25188 );
or \U$24813 ( \25190 , \25187 , \25184 );
xor \U$24814 ( \25191 , \25109 , \25125 );
xor \U$24815 ( \25192 , \25191 , \25130 );
xor \U$24816 ( \25193 , \24653 , \24655 );
xor \U$24817 ( \25194 , \25193 , \24666 );
and \U$24818 ( \25195 , \25192 , \25194 );
xor \U$24819 ( \25196 , \24795 , \24987 );
xor \U$24820 ( \25197 , \25196 , \25080 );
xor \U$24821 ( \25198 , \24653 , \24655 );
xor \U$24822 ( \25199 , \25198 , \24666 );
and \U$24823 ( \25200 , \25197 , \25199 );
and \U$24824 ( \25201 , \25192 , \25197 );
or \U$24825 ( \25202 , \25195 , \25200 , \25201 );
xor \U$24826 ( \25203 , \24371 , \24381 );
xor \U$24827 ( \25204 , \25203 , \24386 );
xor \U$24828 ( \25205 , \25150 , \25157 );
xor \U$24829 ( \25206 , \25204 , \25205 );
xor \U$24830 ( \25207 , \25202 , \25206 );
xor \U$24831 ( \25208 , \24820 , \24845 );
xor \U$24832 ( \25209 , \25208 , \24871 );
xor \U$24833 ( \25210 , \24899 , \24917 );
xor \U$24834 ( \25211 , \25210 , \24943 );
xor \U$24835 ( \25212 , \25209 , \25211 );
xor \U$24836 ( \25213 , \24765 , \24773 );
xor \U$24837 ( \25214 , \25213 , \24782 );
xor \U$24838 ( \25215 , \24974 , \24979 );
xor \U$24839 ( \25216 , \25214 , \25215 );
and \U$24840 ( \25217 , \25212 , \25216 );
and \U$24841 ( \25218 , \25209 , \25211 );
or \U$24842 ( \25219 , \25217 , \25218 );
and \U$24843 ( \25220 , \8371 , RIae781e8_105);
and \U$24844 ( \25221 , RIae785a8_113, \8369 );
nor \U$24845 ( \25222 , \25220 , \25221 );
and \U$24846 ( \25223 , \25222 , \8020 );
not \U$24847 ( \25224 , \25222 );
and \U$24848 ( \25225 , \25224 , \8019 );
nor \U$24849 ( \25226 , \25223 , \25225 );
and \U$24850 ( \25227 , \6941 , RIae782d8_107);
and \U$24851 ( \25228 , RIae780f8_103, \6939 );
nor \U$24852 ( \25229 , \25227 , \25228 );
and \U$24853 ( \25230 , \25229 , \6314 );
not \U$24854 ( \25231 , \25229 );
and \U$24855 ( \25232 , \25231 , \6945 );
nor \U$24856 ( \25233 , \25230 , \25232 );
xor \U$24857 ( \25234 , \25226 , \25233 );
and \U$24858 ( \25235 , \7633 , RIae77f18_99);
and \U$24859 ( \25236 , RIae78008_101, \7631 );
nor \U$24860 ( \25237 , \25235 , \25236 );
and \U$24861 ( \25238 , \25237 , \7206 );
not \U$24862 ( \25239 , \25237 );
and \U$24863 ( \25240 , \25239 , \7205 );
nor \U$24864 ( \25241 , \25238 , \25240 );
and \U$24865 ( \25242 , \25234 , \25241 );
and \U$24866 ( \25243 , \25226 , \25233 );
or \U$24867 ( \25244 , \25242 , \25243 );
and \U$24868 ( \25245 , \6172 , RIae771f8_71);
and \U$24869 ( \25246 , RIae772e8_73, \6170 );
nor \U$24870 ( \25247 , \25245 , \25246 );
and \U$24871 ( \25248 , \25247 , \6176 );
not \U$24872 ( \25249 , \25247 );
and \U$24873 ( \25250 , \25249 , \6175 );
nor \U$24874 ( \25251 , \25248 , \25250 );
and \U$24875 ( \25252 , \5399 , RIae76d48_61);
and \U$24876 ( \25253 , RIae76c58_59, \5397 );
nor \U$24877 ( \25254 , \25252 , \25253 );
and \U$24878 ( \25255 , \25254 , \5016 );
not \U$24879 ( \25256 , \25254 );
and \U$24880 ( \25257 , \25256 , \5403 );
nor \U$24881 ( \25258 , \25255 , \25257 );
xor \U$24882 ( \25259 , \25251 , \25258 );
and \U$24883 ( \25260 , \5896 , RIae77180_70);
and \U$24884 ( \25261 , RIae77018_67, \5894 );
nor \U$24885 ( \25262 , \25260 , \25261 );
and \U$24886 ( \25263 , \25262 , \5590 );
not \U$24887 ( \25264 , \25262 );
and \U$24888 ( \25265 , \25264 , \5589 );
nor \U$24889 ( \25266 , \25263 , \25265 );
and \U$24890 ( \25267 , \25259 , \25266 );
and \U$24891 ( \25268 , \25251 , \25258 );
or \U$24892 ( \25269 , \25267 , \25268 );
xor \U$24893 ( \25270 , \25244 , \25269 );
and \U$24894 ( \25271 , \4688 , RIae76f28_65);
and \U$24895 ( \25272 , RIae76e38_63, \4686 );
nor \U$24896 ( \25273 , \25271 , \25272 );
and \U$24897 ( \25274 , \25273 , \4481 );
not \U$24898 ( \25275 , \25273 );
and \U$24899 ( \25276 , \25275 , \4482 );
nor \U$24900 ( \25277 , \25274 , \25276 );
and \U$24901 ( \25278 , \3730 , RIae77a68_89);
and \U$24902 ( \25279 , RIae77978_87, \3728 );
nor \U$24903 ( \25280 , \25278 , \25279 );
and \U$24904 ( \25281 , \25280 , \3732 );
not \U$24905 ( \25282 , \25280 );
and \U$24906 ( \25283 , \25282 , \3422 );
nor \U$24907 ( \25284 , \25281 , \25283 );
xor \U$24908 ( \25285 , \25277 , \25284 );
and \U$24909 ( \25286 , \4247 , RIae77798_83);
and \U$24910 ( \25287 , RIae77888_85, \4245 );
nor \U$24911 ( \25288 , \25286 , \25287 );
and \U$24912 ( \25289 , \25288 , \3989 );
not \U$24913 ( \25290 , \25288 );
and \U$24914 ( \25291 , \25290 , \4251 );
nor \U$24915 ( \25292 , \25289 , \25291 );
and \U$24916 ( \25293 , \25285 , \25292 );
and \U$24917 ( \25294 , \25277 , \25284 );
or \U$24918 ( \25295 , \25293 , \25294 );
and \U$24919 ( \25296 , \25270 , \25295 );
and \U$24920 ( \25297 , \25244 , \25269 );
or \U$24921 ( \25298 , \25296 , \25297 );
and \U$24922 ( \25299 , \8966 , RIae783c8_109);
and \U$24923 ( \25300 , RIae78530_112, \8964 );
nor \U$24924 ( \25301 , \25299 , \25300 );
and \U$24925 ( \25302 , \25301 , \8799 );
not \U$24926 ( \25303 , \25301 );
and \U$24927 ( \25304 , \25303 , \8789 );
nor \U$24928 ( \25305 , \25302 , \25304 );
and \U$24929 ( \25306 , \9760 , RIae77c48_93);
and \U$24930 ( \25307 , RIae77b58_91, \9758 );
nor \U$24931 ( \25308 , \25306 , \25307 );
and \U$24932 ( \25309 , \25308 , \9273 );
not \U$24933 ( \25310 , \25308 );
and \U$24934 ( \25311 , \25310 , \9764 );
nor \U$24935 ( \25312 , \25309 , \25311 );
xor \U$24936 ( \25313 , \25305 , \25312 );
and \U$24937 ( \25314 , \10548 , RIae77d38_95);
and \U$24938 ( \25315 , RIae77e28_97, \10546 );
nor \U$24939 ( \25316 , \25314 , \25315 );
and \U$24940 ( \25317 , \25316 , \10421 );
not \U$24941 ( \25318 , \25316 );
and \U$24942 ( \25319 , \25318 , \10118 );
nor \U$24943 ( \25320 , \25317 , \25319 );
and \U$24944 ( \25321 , \25313 , \25320 );
and \U$24945 ( \25322 , \25305 , \25312 );
or \U$24946 ( \25323 , \25321 , \25322 );
and \U$24947 ( \25324 , \14059 , RIae75998_19);
and \U$24948 ( \25325 , RIae758a8_17, \14057 );
nor \U$24949 ( \25326 , \25324 , \25325 );
and \U$24950 ( \25327 , \25326 , \13502 );
not \U$24951 ( \25328 , \25326 );
and \U$24952 ( \25329 , \25328 , \14063 );
nor \U$24953 ( \25330 , \25327 , \25329 );
and \U$24954 ( \25331 , \15726 , RIae75c68_25);
and \U$24955 ( \25332 , RIae7aab0_192, RIae75d58_27);
nor \U$24956 ( \25333 , \25331 , \25332 );
and \U$24957 ( \25334 , \25333 , \14959 );
not \U$24958 ( \25335 , \25333 );
and \U$24959 ( \25336 , \25335 , RIae7aa38_191);
nor \U$24960 ( \25337 , \25334 , \25336 );
xor \U$24961 ( \25338 , \25330 , \25337 );
and \U$24962 ( \25339 , \14964 , RIae75f38_31);
and \U$24963 ( \25340 , RIae75e48_29, \14962 );
nor \U$24964 ( \25341 , \25339 , \25340 );
and \U$24965 ( \25342 , \25341 , \14463 );
not \U$24966 ( \25343 , \25341 );
and \U$24967 ( \25344 , \25343 , \14462 );
nor \U$24968 ( \25345 , \25342 , \25344 );
and \U$24969 ( \25346 , \25338 , \25345 );
and \U$24970 ( \25347 , \25330 , \25337 );
or \U$24971 ( \25348 , \25346 , \25347 );
xor \U$24972 ( \25349 , \25323 , \25348 );
and \U$24973 ( \25350 , \11470 , RIae78968_121);
and \U$24974 ( \25351 , RIae78878_119, \11468 );
nor \U$24975 ( \25352 , \25350 , \25351 );
and \U$24976 ( \25353 , \25352 , \10936 );
not \U$24977 ( \25354 , \25352 );
and \U$24978 ( \25355 , \25354 , \11474 );
nor \U$24979 ( \25356 , \25353 , \25355 );
and \U$24980 ( \25357 , \12180 , RIae78788_117);
and \U$24981 ( \25358 , RIae78698_115, \12178 );
nor \U$24982 ( \25359 , \25357 , \25358 );
and \U$24983 ( \25360 , \25359 , \12184 );
not \U$24984 ( \25361 , \25359 );
and \U$24985 ( \25362 , \25361 , \11827 );
nor \U$24986 ( \25363 , \25360 , \25362 );
xor \U$24987 ( \25364 , \25356 , \25363 );
and \U$24988 ( \25365 , \13059 , RIae75b78_23);
and \U$24989 ( \25366 , RIae75a88_21, \13057 );
nor \U$24990 ( \25367 , \25365 , \25366 );
and \U$24991 ( \25368 , \25367 , \13063 );
not \U$24992 ( \25369 , \25367 );
and \U$24993 ( \25370 , \25369 , \12718 );
nor \U$24994 ( \25371 , \25368 , \25370 );
and \U$24995 ( \25372 , \25364 , \25371 );
and \U$24996 ( \25373 , \25356 , \25363 );
or \U$24997 ( \25374 , \25372 , \25373 );
and \U$24998 ( \25375 , \25349 , \25374 );
and \U$24999 ( \25376 , \25323 , \25348 );
or \U$25000 ( \25377 , \25375 , \25376 );
xor \U$25001 ( \25378 , \25298 , \25377 );
xor \U$25002 ( \25379 , \24954 , \24962 );
xor \U$25003 ( \25380 , \25379 , \24971 );
nand \U$25004 ( \25381 , RIae775b8_79, \2605 );
and \U$25005 ( \25382 , \25381 , \2611 );
not \U$25006 ( \25383 , \25381 );
and \U$25007 ( \25384 , \25383 , \2397 );
nor \U$25008 ( \25385 , \25382 , \25384 );
xor \U$25009 ( \25386 , \25380 , \25385 );
xor \U$25010 ( \25387 , \24827 , \24834 );
xor \U$25011 ( \25388 , \25387 , \24842 );
and \U$25012 ( \25389 , \25386 , \25388 );
and \U$25013 ( \25390 , \25380 , \25385 );
or \U$25014 ( \25391 , \25389 , \25390 );
and \U$25015 ( \25392 , \25378 , \25391 );
and \U$25016 ( \25393 , \25298 , \25377 );
or \U$25017 ( \25394 , \25392 , \25393 );
xor \U$25018 ( \25395 , \25219 , \25394 );
xor \U$25019 ( \25396 , \24802 , \24809 );
xor \U$25020 ( \25397 , \25396 , \24817 );
xor \U$25021 ( \25398 , \24853 , \24860 );
xor \U$25022 ( \25399 , \25398 , \24868 );
and \U$25023 ( \25400 , \25397 , \25399 );
xor \U$25024 ( \25401 , \24881 , \24888 );
xor \U$25025 ( \25402 , \25401 , \24896 );
xor \U$25026 ( \25403 , \24853 , \24860 );
xor \U$25027 ( \25404 , \25403 , \24868 );
and \U$25028 ( \25405 , \25402 , \25404 );
and \U$25029 ( \25406 , \25397 , \25402 );
or \U$25030 ( \25407 , \25400 , \25405 , \25406 );
xor \U$25031 ( \25408 , \25044 , \25067 );
xor \U$25032 ( \25409 , \25407 , \25408 );
xor \U$25033 ( \25410 , \24679 , \24686 );
xor \U$25034 ( \25411 , \25410 , \24694 );
xor \U$25035 ( \25412 , \24990 , \25016 );
xor \U$25036 ( \25413 , \25411 , \25412 );
and \U$25037 ( \25414 , \25409 , \25413 );
and \U$25038 ( \25415 , \25407 , \25408 );
or \U$25039 ( \25416 , \25414 , \25415 );
and \U$25040 ( \25417 , \25395 , \25416 );
and \U$25041 ( \25418 , \25219 , \25394 );
or \U$25042 ( \25419 , \25417 , \25418 );
xor \U$25043 ( \25420 , \25095 , \25097 );
xor \U$25044 ( \25421 , \25420 , \25102 );
xor \U$25045 ( \25422 , \25419 , \25421 );
xor \U$25046 ( \25423 , \25113 , \25117 );
xor \U$25047 ( \25424 , \25423 , \25122 );
xor \U$25048 ( \25425 , \25021 , \25068 );
xor \U$25049 ( \25426 , \25425 , \25077 );
and \U$25050 ( \25427 , \25424 , \25426 );
xor \U$25051 ( \25428 , \24751 , \24753 );
xor \U$25052 ( \25429 , \25428 , \24756 );
xor \U$25053 ( \25430 , \24749 , \24790 );
xor \U$25054 ( \25431 , \25429 , \25430 );
xor \U$25055 ( \25432 , \25021 , \25068 );
xor \U$25056 ( \25433 , \25432 , \25077 );
and \U$25057 ( \25434 , \25431 , \25433 );
and \U$25058 ( \25435 , \25424 , \25431 );
or \U$25059 ( \25436 , \25427 , \25434 , \25435 );
and \U$25060 ( \25437 , \25422 , \25436 );
and \U$25061 ( \25438 , \25419 , \25421 );
or \U$25062 ( \25439 , \25437 , \25438 );
and \U$25063 ( \25440 , \25207 , \25439 );
and \U$25064 ( \25441 , \25202 , \25206 );
or \U$25065 ( \25442 , \25440 , \25441 );
nand \U$25066 ( \25443 , \25190 , \25442 );
nand \U$25067 ( \25444 , \25189 , \25443 );
and \U$25068 ( \25445 , \25179 , \25444 );
xor \U$25069 ( \25446 , \25444 , \25179 );
xor \U$25070 ( \25447 , \25181 , \25183 );
xor \U$25071 ( \25448 , \25202 , \25206 );
xor \U$25072 ( \25449 , \25448 , \25439 );
xor \U$25073 ( \25450 , \25447 , \25449 );
xor \U$25074 ( \25451 , \25356 , \25363 );
xor \U$25075 ( \25452 , \25451 , \25371 );
xor \U$25076 ( \25453 , \25330 , \25337 );
xor \U$25077 ( \25454 , \25453 , \25345 );
xor \U$25078 ( \25455 , \25452 , \25454 );
xor \U$25079 ( \25456 , \25305 , \25312 );
xor \U$25080 ( \25457 , \25456 , \25320 );
and \U$25081 ( \25458 , \25455 , \25457 );
and \U$25082 ( \25459 , \25452 , \25454 );
or \U$25083 ( \25460 , \25458 , \25459 );
xor \U$25084 ( \25461 , \24925 , \24932 );
xor \U$25085 ( \25462 , \25461 , \24940 );
xor \U$25086 ( \25463 , \25460 , \25462 );
xor \U$25087 ( \25464 , \25251 , \25258 );
xor \U$25088 ( \25465 , \25464 , \25266 );
xor \U$25089 ( \25466 , \25277 , \25284 );
xor \U$25090 ( \25467 , \25466 , \25292 );
and \U$25091 ( \25468 , \25465 , \25467 );
xor \U$25092 ( \25469 , \25226 , \25233 );
xor \U$25093 ( \25470 , \25469 , \25241 );
xor \U$25094 ( \25471 , \25277 , \25284 );
xor \U$25095 ( \25472 , \25471 , \25292 );
and \U$25096 ( \25473 , \25470 , \25472 );
and \U$25097 ( \25474 , \25465 , \25470 );
or \U$25098 ( \25475 , \25468 , \25473 , \25474 );
and \U$25099 ( \25476 , \25463 , \25475 );
and \U$25100 ( \25477 , \25460 , \25462 );
or \U$25101 ( \25478 , \25476 , \25477 );
and \U$25102 ( \25479 , \12180 , RIae78878_119);
and \U$25103 ( \25480 , RIae78788_117, \12178 );
nor \U$25104 ( \25481 , \25479 , \25480 );
and \U$25105 ( \25482 , \25481 , \12184 );
not \U$25106 ( \25483 , \25481 );
and \U$25107 ( \25484 , \25483 , \11827 );
nor \U$25108 ( \25485 , \25482 , \25484 );
and \U$25109 ( \25486 , \13059 , RIae78698_115);
and \U$25110 ( \25487 , RIae75b78_23, \13057 );
nor \U$25111 ( \25488 , \25486 , \25487 );
and \U$25112 ( \25489 , \25488 , \13063 );
not \U$25113 ( \25490 , \25488 );
and \U$25114 ( \25491 , \25490 , \12718 );
nor \U$25115 ( \25492 , \25489 , \25491 );
xor \U$25116 ( \25493 , \25485 , \25492 );
and \U$25117 ( \25494 , \14059 , RIae75a88_21);
and \U$25118 ( \25495 , RIae75998_19, \14057 );
nor \U$25119 ( \25496 , \25494 , \25495 );
and \U$25120 ( \25497 , \25496 , \13502 );
not \U$25121 ( \25498 , \25496 );
and \U$25122 ( \25499 , \25498 , \14063 );
nor \U$25123 ( \25500 , \25497 , \25499 );
and \U$25124 ( \25501 , \25493 , \25500 );
and \U$25125 ( \25502 , \25485 , \25492 );
or \U$25126 ( \25503 , \25501 , \25502 );
and \U$25127 ( \25504 , \15726 , RIae75e48_29);
and \U$25128 ( \25505 , RIae7aab0_192, RIae75c68_25);
nor \U$25129 ( \25506 , \25504 , \25505 );
and \U$25130 ( \25507 , \25506 , \14959 );
not \U$25131 ( \25508 , \25506 );
and \U$25132 ( \25509 , \25508 , RIae7aa38_191);
nor \U$25133 ( \25510 , \25507 , \25509 );
xor \U$25134 ( \25511 , \25510 , \2789 );
and \U$25135 ( \25512 , \14964 , RIae758a8_17);
and \U$25136 ( \25513 , RIae75f38_31, \14962 );
nor \U$25137 ( \25514 , \25512 , \25513 );
and \U$25138 ( \25515 , \25514 , \14463 );
not \U$25139 ( \25516 , \25514 );
and \U$25140 ( \25517 , \25516 , \14462 );
nor \U$25141 ( \25518 , \25515 , \25517 );
and \U$25142 ( \25519 , \25511 , \25518 );
and \U$25143 ( \25520 , \25510 , \2789 );
or \U$25144 ( \25521 , \25519 , \25520 );
xor \U$25145 ( \25522 , \25503 , \25521 );
and \U$25146 ( \25523 , \10548 , RIae77b58_91);
and \U$25147 ( \25524 , RIae77d38_95, \10546 );
nor \U$25148 ( \25525 , \25523 , \25524 );
and \U$25149 ( \25526 , \25525 , \10421 );
not \U$25150 ( \25527 , \25525 );
and \U$25151 ( \25528 , \25527 , \10118 );
nor \U$25152 ( \25529 , \25526 , \25528 );
and \U$25153 ( \25530 , \9760 , RIae78530_112);
and \U$25154 ( \25531 , RIae77c48_93, \9758 );
nor \U$25155 ( \25532 , \25530 , \25531 );
and \U$25156 ( \25533 , \25532 , \9273 );
not \U$25157 ( \25534 , \25532 );
and \U$25158 ( \25535 , \25534 , \9272 );
nor \U$25159 ( \25536 , \25533 , \25535 );
xor \U$25160 ( \25537 , \25529 , \25536 );
and \U$25161 ( \25538 , \11470 , RIae77e28_97);
and \U$25162 ( \25539 , RIae78968_121, \11468 );
nor \U$25163 ( \25540 , \25538 , \25539 );
and \U$25164 ( \25541 , \25540 , \10936 );
not \U$25165 ( \25542 , \25540 );
and \U$25166 ( \25543 , \25542 , \11474 );
nor \U$25167 ( \25544 , \25541 , \25543 );
and \U$25168 ( \25545 , \25537 , \25544 );
and \U$25169 ( \25546 , \25529 , \25536 );
or \U$25170 ( \25547 , \25545 , \25546 );
and \U$25171 ( \25548 , \25522 , \25547 );
and \U$25172 ( \25549 , \25503 , \25521 );
or \U$25173 ( \25550 , \25548 , \25549 );
not \U$25174 ( \25551 , \3218 );
and \U$25175 ( \25552 , \3214 , RIae77720_82);
and \U$25176 ( \25553 , RIae773d8_75, \3212 );
nor \U$25177 ( \25554 , \25552 , \25553 );
not \U$25178 ( \25555 , \25554 );
or \U$25179 ( \25556 , \25551 , \25555 );
or \U$25180 ( \25557 , \25554 , \2774 );
nand \U$25181 ( \25558 , \25556 , \25557 );
not \U$25182 ( \25559 , \2789 );
and \U$25183 ( \25560 , \2783 , RIae775b8_79);
and \U$25184 ( \25561 , RIae774c8_77, \2781 );
nor \U$25185 ( \25562 , \25560 , \25561 );
not \U$25186 ( \25563 , \25562 );
or \U$25187 ( \25564 , \25559 , \25563 );
or \U$25188 ( \25565 , \25562 , \3089 );
nand \U$25189 ( \25566 , \25564 , \25565 );
xor \U$25190 ( \25567 , \25558 , \25566 );
not \U$25191 ( \25568 , \3218 );
and \U$25192 ( \25569 , \3214 , RIae774c8_77);
and \U$25193 ( \25570 , RIae77720_82, \3212 );
nor \U$25194 ( \25571 , \25569 , \25570 );
not \U$25195 ( \25572 , \25571 );
or \U$25196 ( \25573 , \25568 , \25572 );
or \U$25197 ( \25574 , \25571 , \3218 );
nand \U$25198 ( \25575 , \25573 , \25574 );
nand \U$25199 ( \25576 , RIae775b8_79, \2781 );
not \U$25200 ( \25577 , \25576 );
not \U$25201 ( \25578 , \3089 );
or \U$25202 ( \25579 , \25577 , \25578 );
or \U$25203 ( \25580 , \2789 , \25576 );
nand \U$25204 ( \25581 , \25579 , \25580 );
xor \U$25205 ( \25582 , \25575 , \25581 );
and \U$25206 ( \25583 , \3730 , RIae773d8_75);
and \U$25207 ( \25584 , RIae77a68_89, \3728 );
nor \U$25208 ( \25585 , \25583 , \25584 );
and \U$25209 ( \25586 , \25585 , \3732 );
not \U$25210 ( \25587 , \25585 );
and \U$25211 ( \25588 , \25587 , \3421 );
nor \U$25212 ( \25589 , \25586 , \25588 );
and \U$25213 ( \25590 , \25582 , \25589 );
and \U$25214 ( \25591 , \25575 , \25581 );
or \U$25215 ( \25592 , \25590 , \25591 );
and \U$25216 ( \25593 , \25567 , \25592 );
and \U$25217 ( \25594 , \25558 , \25566 );
or \U$25218 ( \25595 , \25593 , \25594 );
xor \U$25219 ( \25596 , \25550 , \25595 );
and \U$25220 ( \25597 , \5896 , RIae76c58_59);
and \U$25221 ( \25598 , RIae77180_70, \5894 );
nor \U$25222 ( \25599 , \25597 , \25598 );
and \U$25223 ( \25600 , \25599 , \5590 );
not \U$25224 ( \25601 , \25599 );
and \U$25225 ( \25602 , \25601 , \5589 );
nor \U$25226 ( \25603 , \25600 , \25602 );
and \U$25227 ( \25604 , \6172 , RIae77018_67);
and \U$25228 ( \25605 , RIae771f8_71, \6170 );
nor \U$25229 ( \25606 , \25604 , \25605 );
and \U$25230 ( \25607 , \25606 , \6176 );
not \U$25231 ( \25608 , \25606 );
and \U$25232 ( \25609 , \25608 , \6175 );
nor \U$25233 ( \25610 , \25607 , \25609 );
xor \U$25234 ( \25611 , \25603 , \25610 );
and \U$25235 ( \25612 , \6941 , RIae772e8_73);
and \U$25236 ( \25613 , RIae782d8_107, \6939 );
nor \U$25237 ( \25614 , \25612 , \25613 );
and \U$25238 ( \25615 , \25614 , \6314 );
not \U$25239 ( \25616 , \25614 );
and \U$25240 ( \25617 , \25616 , \6945 );
nor \U$25241 ( \25618 , \25615 , \25617 );
and \U$25242 ( \25619 , \25611 , \25618 );
and \U$25243 ( \25620 , \25603 , \25610 );
or \U$25244 ( \25621 , \25619 , \25620 );
and \U$25245 ( \25622 , \4247 , RIae77978_87);
and \U$25246 ( \25623 , RIae77798_83, \4245 );
nor \U$25247 ( \25624 , \25622 , \25623 );
and \U$25248 ( \25625 , \25624 , \3989 );
not \U$25249 ( \25626 , \25624 );
and \U$25250 ( \25627 , \25626 , \4251 );
nor \U$25251 ( \25628 , \25625 , \25627 );
and \U$25252 ( \25629 , \4688 , RIae77888_85);
and \U$25253 ( \25630 , RIae76f28_65, \4686 );
nor \U$25254 ( \25631 , \25629 , \25630 );
and \U$25255 ( \25632 , \25631 , \4481 );
not \U$25256 ( \25633 , \25631 );
and \U$25257 ( \25634 , \25633 , \4482 );
nor \U$25258 ( \25635 , \25632 , \25634 );
xor \U$25259 ( \25636 , \25628 , \25635 );
and \U$25260 ( \25637 , \5399 , RIae76e38_63);
and \U$25261 ( \25638 , RIae76d48_61, \5397 );
nor \U$25262 ( \25639 , \25637 , \25638 );
and \U$25263 ( \25640 , \25639 , \5016 );
not \U$25264 ( \25641 , \25639 );
and \U$25265 ( \25642 , \25641 , \5403 );
nor \U$25266 ( \25643 , \25640 , \25642 );
and \U$25267 ( \25644 , \25636 , \25643 );
and \U$25268 ( \25645 , \25628 , \25635 );
or \U$25269 ( \25646 , \25644 , \25645 );
xor \U$25270 ( \25647 , \25621 , \25646 );
and \U$25271 ( \25648 , \8371 , RIae78008_101);
and \U$25272 ( \25649 , RIae781e8_105, \8369 );
nor \U$25273 ( \25650 , \25648 , \25649 );
and \U$25274 ( \25651 , \25650 , \8020 );
not \U$25275 ( \25652 , \25650 );
and \U$25276 ( \25653 , \25652 , \8019 );
nor \U$25277 ( \25654 , \25651 , \25653 );
and \U$25278 ( \25655 , \7633 , RIae780f8_103);
and \U$25279 ( \25656 , RIae77f18_99, \7631 );
nor \U$25280 ( \25657 , \25655 , \25656 );
and \U$25281 ( \25658 , \25657 , \7206 );
not \U$25282 ( \25659 , \25657 );
and \U$25283 ( \25660 , \25659 , \7205 );
nor \U$25284 ( \25661 , \25658 , \25660 );
xor \U$25285 ( \25662 , \25654 , \25661 );
and \U$25286 ( \25663 , \8966 , RIae785a8_113);
and \U$25287 ( \25664 , RIae783c8_109, \8964 );
nor \U$25288 ( \25665 , \25663 , \25664 );
and \U$25289 ( \25666 , \25665 , \8799 );
not \U$25290 ( \25667 , \25665 );
and \U$25291 ( \25668 , \25667 , \8789 );
nor \U$25292 ( \25669 , \25666 , \25668 );
and \U$25293 ( \25670 , \25662 , \25669 );
and \U$25294 ( \25671 , \25654 , \25661 );
or \U$25295 ( \25672 , \25670 , \25671 );
and \U$25296 ( \25673 , \25647 , \25672 );
and \U$25297 ( \25674 , \25621 , \25646 );
or \U$25298 ( \25675 , \25673 , \25674 );
and \U$25299 ( \25676 , \25596 , \25675 );
and \U$25300 ( \25677 , \25550 , \25595 );
or \U$25301 ( \25678 , \25676 , \25677 );
xor \U$25302 ( \25679 , \25478 , \25678 );
xor \U$25303 ( \25680 , \24906 , \2397 );
xor \U$25304 ( \25681 , \25680 , \24914 );
xor \U$25305 ( \25682 , \25380 , \25385 );
xor \U$25306 ( \25683 , \25682 , \25388 );
and \U$25307 ( \25684 , \25681 , \25683 );
xor \U$25308 ( \25685 , \24853 , \24860 );
xor \U$25309 ( \25686 , \25685 , \24868 );
xor \U$25310 ( \25687 , \25397 , \25402 );
xor \U$25311 ( \25688 , \25686 , \25687 );
xor \U$25312 ( \25689 , \25380 , \25385 );
xor \U$25313 ( \25690 , \25689 , \25388 );
and \U$25314 ( \25691 , \25688 , \25690 );
and \U$25315 ( \25692 , \25681 , \25688 );
or \U$25316 ( \25693 , \25684 , \25691 , \25692 );
and \U$25317 ( \25694 , \25679 , \25693 );
and \U$25318 ( \25695 , \25478 , \25678 );
or \U$25319 ( \25696 , \25694 , \25695 );
xor \U$25320 ( \25697 , \24874 , \24946 );
xor \U$25321 ( \25698 , \25697 , \24984 );
xor \U$25322 ( \25699 , \25696 , \25698 );
xor \U$25323 ( \25700 , \25298 , \25377 );
xor \U$25324 ( \25701 , \25700 , \25391 );
xor \U$25325 ( \25702 , \25209 , \25211 );
xor \U$25326 ( \25703 , \25702 , \25216 );
and \U$25327 ( \25704 , \25701 , \25703 );
xor \U$25328 ( \25705 , \25407 , \25408 );
xor \U$25329 ( \25706 , \25705 , \25413 );
xor \U$25330 ( \25707 , \25209 , \25211 );
xor \U$25331 ( \25708 , \25707 , \25216 );
and \U$25332 ( \25709 , \25706 , \25708 );
and \U$25333 ( \25710 , \25701 , \25706 );
or \U$25334 ( \25711 , \25704 , \25709 , \25710 );
and \U$25335 ( \25712 , \25699 , \25711 );
and \U$25336 ( \25713 , \25696 , \25698 );
or \U$25337 ( \25714 , \25712 , \25713 );
xor \U$25338 ( \25715 , \25219 , \25394 );
xor \U$25339 ( \25716 , \25715 , \25416 );
xor \U$25340 ( \25717 , \25021 , \25068 );
xor \U$25341 ( \25718 , \25717 , \25077 );
xor \U$25342 ( \25719 , \25424 , \25431 );
xor \U$25343 ( \25720 , \25718 , \25719 );
and \U$25344 ( \25721 , \25716 , \25720 );
xor \U$25345 ( \25722 , \25714 , \25721 );
xor \U$25346 ( \25723 , \24653 , \24655 );
xor \U$25347 ( \25724 , \25723 , \24666 );
xor \U$25348 ( \25725 , \25192 , \25197 );
xor \U$25349 ( \25726 , \25724 , \25725 );
and \U$25350 ( \25727 , \25722 , \25726 );
and \U$25351 ( \25728 , \25714 , \25721 );
or \U$25352 ( \25729 , \25727 , \25728 );
and \U$25353 ( \25730 , \25450 , \25729 );
and \U$25354 ( \25731 , \25447 , \25449 );
nor \U$25355 ( \25732 , \25730 , \25731 );
xnor \U$25356 ( \25733 , \25184 , \25442 );
not \U$25357 ( \25734 , \25733 );
not \U$25358 ( \25735 , \25187 );
and \U$25359 ( \25736 , \25734 , \25735 );
and \U$25360 ( \25737 , \25733 , \25187 );
nor \U$25361 ( \25738 , \25736 , \25737 );
or \U$25362 ( \25739 , \25732 , \25738 );
xnor \U$25363 ( \25740 , \25738 , \25732 );
and \U$25364 ( \25741 , \8371 , RIae77f18_99);
and \U$25365 ( \25742 , RIae78008_101, \8369 );
nor \U$25366 ( \25743 , \25741 , \25742 );
and \U$25367 ( \25744 , \25743 , \8020 );
not \U$25368 ( \25745 , \25743 );
and \U$25369 ( \25746 , \25745 , \8019 );
nor \U$25370 ( \25747 , \25744 , \25746 );
and \U$25371 ( \25748 , \6941 , RIae771f8_71);
and \U$25372 ( \25749 , RIae772e8_73, \6939 );
nor \U$25373 ( \25750 , \25748 , \25749 );
and \U$25374 ( \25751 , \25750 , \6314 );
not \U$25375 ( \25752 , \25750 );
and \U$25376 ( \25753 , \25752 , \6945 );
nor \U$25377 ( \25754 , \25751 , \25753 );
xor \U$25378 ( \25755 , \25747 , \25754 );
and \U$25379 ( \25756 , \7633 , RIae782d8_107);
and \U$25380 ( \25757 , RIae780f8_103, \7631 );
nor \U$25381 ( \25758 , \25756 , \25757 );
and \U$25382 ( \25759 , \25758 , \7206 );
not \U$25383 ( \25760 , \25758 );
and \U$25384 ( \25761 , \25760 , \7205 );
nor \U$25385 ( \25762 , \25759 , \25761 );
xor \U$25386 ( \25763 , \25755 , \25762 );
and \U$25387 ( \25764 , \11470 , RIae77d38_95);
and \U$25388 ( \25765 , RIae77e28_97, \11468 );
nor \U$25389 ( \25766 , \25764 , \25765 );
and \U$25390 ( \25767 , \25766 , \10936 );
not \U$25391 ( \25768 , \25766 );
and \U$25392 ( \25769 , \25768 , \11474 );
nor \U$25393 ( \25770 , \25767 , \25769 );
and \U$25394 ( \25771 , \12180 , RIae78968_121);
and \U$25395 ( \25772 , RIae78878_119, \12178 );
nor \U$25396 ( \25773 , \25771 , \25772 );
and \U$25397 ( \25774 , \25773 , \12184 );
not \U$25398 ( \25775 , \25773 );
and \U$25399 ( \25776 , \25775 , \11827 );
nor \U$25400 ( \25777 , \25774 , \25776 );
xor \U$25401 ( \25778 , \25770 , \25777 );
and \U$25402 ( \25779 , \13059 , RIae78788_117);
and \U$25403 ( \25780 , RIae78698_115, \13057 );
nor \U$25404 ( \25781 , \25779 , \25780 );
and \U$25405 ( \25782 , \25781 , \13063 );
not \U$25406 ( \25783 , \25781 );
and \U$25407 ( \25784 , \25783 , \12718 );
nor \U$25408 ( \25785 , \25782 , \25784 );
xor \U$25409 ( \25786 , \25778 , \25785 );
and \U$25410 ( \25787 , \25763 , \25786 );
and \U$25411 ( \25788 , \10548 , RIae77c48_93);
and \U$25412 ( \25789 , RIae77b58_91, \10546 );
nor \U$25413 ( \25790 , \25788 , \25789 );
and \U$25414 ( \25791 , \25790 , \10421 );
not \U$25415 ( \25792 , \25790 );
and \U$25416 ( \25793 , \25792 , \10118 );
nor \U$25417 ( \25794 , \25791 , \25793 );
and \U$25418 ( \25795 , \8966 , RIae781e8_105);
and \U$25419 ( \25796 , RIae785a8_113, \8964 );
nor \U$25420 ( \25797 , \25795 , \25796 );
and \U$25421 ( \25798 , \25797 , \8799 );
not \U$25422 ( \25799 , \25797 );
and \U$25423 ( \25800 , \25799 , \8789 );
nor \U$25424 ( \25801 , \25798 , \25800 );
xor \U$25425 ( \25802 , \25794 , \25801 );
and \U$25426 ( \25803 , \9760 , RIae783c8_109);
and \U$25427 ( \25804 , RIae78530_112, \9758 );
nor \U$25428 ( \25805 , \25803 , \25804 );
and \U$25429 ( \25806 , \25805 , \9273 );
not \U$25430 ( \25807 , \25805 );
and \U$25431 ( \25808 , \25807 , \9272 );
nor \U$25432 ( \25809 , \25806 , \25808 );
xor \U$25433 ( \25810 , \25802 , \25809 );
xor \U$25434 ( \25811 , \25770 , \25777 );
xor \U$25435 ( \25812 , \25811 , \25785 );
and \U$25436 ( \25813 , \25810 , \25812 );
and \U$25437 ( \25814 , \25763 , \25810 );
or \U$25438 ( \25815 , \25787 , \25813 , \25814 );
xor \U$25439 ( \25816 , \25510 , \2789 );
xor \U$25440 ( \25817 , \25816 , \25518 );
xor \U$25441 ( \25818 , \25815 , \25817 );
xor \U$25442 ( \25819 , \25529 , \25536 );
xor \U$25443 ( \25820 , \25819 , \25544 );
xor \U$25444 ( \25821 , \25654 , \25661 );
xor \U$25445 ( \25822 , \25821 , \25669 );
xor \U$25446 ( \25823 , \25485 , \25492 );
xor \U$25447 ( \25824 , \25823 , \25500 );
xor \U$25448 ( \25825 , \25822 , \25824 );
xor \U$25449 ( \25826 , \25820 , \25825 );
and \U$25450 ( \25827 , \25818 , \25826 );
and \U$25451 ( \25828 , \25815 , \25817 );
or \U$25452 ( \25829 , \25827 , \25828 );
and \U$25453 ( \25830 , \8371 , RIae780f8_103);
and \U$25454 ( \25831 , RIae77f18_99, \8369 );
nor \U$25455 ( \25832 , \25830 , \25831 );
and \U$25456 ( \25833 , \25832 , \8019 );
not \U$25457 ( \25834 , \25832 );
and \U$25458 ( \25835 , \25834 , \8020 );
nor \U$25459 ( \25836 , \25833 , \25835 );
and \U$25460 ( \25837 , \8966 , RIae78008_101);
and \U$25461 ( \25838 , RIae781e8_105, \8964 );
nor \U$25462 ( \25839 , \25837 , \25838 );
and \U$25463 ( \25840 , \25839 , \8789 );
not \U$25464 ( \25841 , \25839 );
and \U$25465 ( \25842 , \25841 , \8799 );
nor \U$25466 ( \25843 , \25840 , \25842 );
xor \U$25467 ( \25844 , \25836 , \25843 );
and \U$25468 ( \25845 , \7633 , RIae772e8_73);
and \U$25469 ( \25846 , RIae782d8_107, \7631 );
nor \U$25470 ( \25847 , \25845 , \25846 );
and \U$25471 ( \25848 , \25847 , \7205 );
not \U$25472 ( \25849 , \25847 );
and \U$25473 ( \25850 , \25849 , \7206 );
nor \U$25474 ( \25851 , \25848 , \25850 );
and \U$25475 ( \25852 , \25844 , \25851 );
and \U$25476 ( \25853 , \25836 , \25843 );
nor \U$25477 ( \25854 , \25852 , \25853 );
and \U$25478 ( \25855 , \6172 , RIae76c58_59);
and \U$25479 ( \25856 , RIae77180_70, \6170 );
nor \U$25480 ( \25857 , \25855 , \25856 );
and \U$25481 ( \25858 , \25857 , \6175 );
not \U$25482 ( \25859 , \25857 );
and \U$25483 ( \25860 , \25859 , \6176 );
nor \U$25484 ( \25861 , \25858 , \25860 );
and \U$25485 ( \25862 , \6941 , RIae77018_67);
and \U$25486 ( \25863 , RIae771f8_71, \6939 );
nor \U$25487 ( \25864 , \25862 , \25863 );
and \U$25488 ( \25865 , \25864 , \6945 );
not \U$25489 ( \25866 , \25864 );
and \U$25490 ( \25867 , \25866 , \6314 );
nor \U$25491 ( \25868 , \25865 , \25867 );
xor \U$25492 ( \25869 , \25861 , \25868 );
and \U$25493 ( \25870 , \5896 , RIae76e38_63);
and \U$25494 ( \25871 , RIae76d48_61, \5894 );
nor \U$25495 ( \25872 , \25870 , \25871 );
and \U$25496 ( \25873 , \25872 , \5589 );
not \U$25497 ( \25874 , \25872 );
and \U$25498 ( \25875 , \25874 , \5590 );
nor \U$25499 ( \25876 , \25873 , \25875 );
and \U$25500 ( \25877 , \25869 , \25876 );
and \U$25501 ( \25878 , \25861 , \25868 );
nor \U$25502 ( \25879 , \25877 , \25878 );
xor \U$25503 ( \25880 , \25854 , \25879 );
and \U$25504 ( \25881 , \5399 , RIae77888_85);
and \U$25505 ( \25882 , RIae76f28_65, \5397 );
nor \U$25506 ( \25883 , \25881 , \25882 );
and \U$25507 ( \25884 , \25883 , \5016 );
not \U$25508 ( \25885 , \25883 );
and \U$25509 ( \25886 , \25885 , \5403 );
nor \U$25510 ( \25887 , \25884 , \25886 );
and \U$25511 ( \25888 , \4247 , RIae773d8_75);
and \U$25512 ( \25889 , RIae77a68_89, \4245 );
nor \U$25513 ( \25890 , \25888 , \25889 );
and \U$25514 ( \25891 , \25890 , \3989 );
not \U$25515 ( \25892 , \25890 );
and \U$25516 ( \25893 , \25892 , \4251 );
nor \U$25517 ( \25894 , \25891 , \25893 );
xor \U$25518 ( \25895 , \25887 , \25894 );
and \U$25519 ( \25896 , \4688 , RIae77978_87);
and \U$25520 ( \25897 , RIae77798_83, \4686 );
nor \U$25521 ( \25898 , \25896 , \25897 );
and \U$25522 ( \25899 , \25898 , \4481 );
not \U$25523 ( \25900 , \25898 );
and \U$25524 ( \25901 , \25900 , \4482 );
nor \U$25525 ( \25902 , \25899 , \25901 );
and \U$25526 ( \25903 , \25895 , \25902 );
and \U$25527 ( \25904 , \25887 , \25894 );
or \U$25528 ( \25905 , \25903 , \25904 );
and \U$25529 ( \25906 , \25880 , \25905 );
and \U$25530 ( \25907 , \25854 , \25879 );
or \U$25531 ( \25908 , \25906 , \25907 );
and \U$25532 ( \25909 , \15726 , RIae758a8_17);
and \U$25533 ( \25910 , RIae7aab0_192, RIae75f38_31);
nor \U$25534 ( \25911 , \25909 , \25910 );
and \U$25535 ( \25912 , \25911 , \14959 );
not \U$25536 ( \25913 , \25911 );
and \U$25537 ( \25914 , \25913 , RIae7aa38_191);
nor \U$25538 ( \25915 , \25912 , \25914 );
xor \U$25539 ( \25916 , \25915 , \3218 );
and \U$25540 ( \25917 , \14964 , RIae75a88_21);
and \U$25541 ( \25918 , RIae75998_19, \14962 );
nor \U$25542 ( \25919 , \25917 , \25918 );
and \U$25543 ( \25920 , \25919 , \14463 );
not \U$25544 ( \25921 , \25919 );
and \U$25545 ( \25922 , \25921 , \14462 );
nor \U$25546 ( \25923 , \25920 , \25922 );
and \U$25547 ( \25924 , \25916 , \25923 );
and \U$25548 ( \25925 , \25915 , \3218 );
or \U$25549 ( \25926 , \25924 , \25925 );
not \U$25550 ( \25927 , \25926 );
and \U$25551 ( \25928 , \13059 , RIae78878_119);
and \U$25552 ( \25929 , RIae78788_117, \13057 );
nor \U$25553 ( \25930 , \25928 , \25929 );
and \U$25554 ( \25931 , \25930 , \12718 );
not \U$25555 ( \25932 , \25930 );
and \U$25556 ( \25933 , \25932 , \13063 );
nor \U$25557 ( \25934 , \25931 , \25933 );
and \U$25558 ( \25935 , \14059 , RIae78698_115);
and \U$25559 ( \25936 , RIae75b78_23, \14057 );
nor \U$25560 ( \25937 , \25935 , \25936 );
and \U$25561 ( \25938 , \25937 , \14063 );
not \U$25562 ( \25939 , \25937 );
and \U$25563 ( \25940 , \25939 , \13502 );
nor \U$25564 ( \25941 , \25938 , \25940 );
xor \U$25565 ( \25942 , \25934 , \25941 );
and \U$25566 ( \25943 , \12180 , RIae77e28_97);
and \U$25567 ( \25944 , RIae78968_121, \12178 );
nor \U$25568 ( \25945 , \25943 , \25944 );
and \U$25569 ( \25946 , \25945 , \11827 );
not \U$25570 ( \25947 , \25945 );
and \U$25571 ( \25948 , \25947 , \12184 );
nor \U$25572 ( \25949 , \25946 , \25948 );
and \U$25573 ( \25950 , \25942 , \25949 );
and \U$25574 ( \25951 , \25934 , \25941 );
nor \U$25575 ( \25952 , \25950 , \25951 );
not \U$25576 ( \25953 , \25952 );
or \U$25577 ( \25954 , \25927 , \25953 );
or \U$25578 ( \25955 , \25952 , \25926 );
and \U$25579 ( \25956 , \9760 , RIae785a8_113);
and \U$25580 ( \25957 , RIae783c8_109, \9758 );
nor \U$25581 ( \25958 , \25956 , \25957 );
and \U$25582 ( \25959 , \25958 , \9272 );
not \U$25583 ( \25960 , \25958 );
and \U$25584 ( \25961 , \25960 , \9273 );
nor \U$25585 ( \25962 , \25959 , \25961 );
and \U$25586 ( \25963 , \10548 , RIae78530_112);
and \U$25587 ( \25964 , RIae77c48_93, \10546 );
nor \U$25588 ( \25965 , \25963 , \25964 );
and \U$25589 ( \25966 , \25965 , \10118 );
not \U$25590 ( \25967 , \25965 );
and \U$25591 ( \25968 , \25967 , \10421 );
nor \U$25592 ( \25969 , \25966 , \25968 );
or \U$25593 ( \25970 , \25962 , \25969 );
not \U$25594 ( \25971 , \25969 );
not \U$25595 ( \25972 , \25962 );
or \U$25596 ( \25973 , \25971 , \25972 );
and \U$25597 ( \25974 , \11470 , RIae77b58_91);
and \U$25598 ( \25975 , RIae77d38_95, \11468 );
nor \U$25599 ( \25976 , \25974 , \25975 );
and \U$25600 ( \25977 , \25976 , \10936 );
not \U$25601 ( \25978 , \25976 );
and \U$25602 ( \25979 , \25978 , \11474 );
nor \U$25603 ( \25980 , \25977 , \25979 );
nand \U$25604 ( \25981 , \25973 , \25980 );
nand \U$25605 ( \25982 , \25970 , \25981 );
nand \U$25606 ( \25983 , \25955 , \25982 );
nand \U$25607 ( \25984 , \25954 , \25983 );
xor \U$25608 ( \25985 , \25908 , \25984 );
not \U$25609 ( \25986 , \2774 );
and \U$25610 ( \25987 , \3214 , RIae775b8_79);
and \U$25611 ( \25988 , RIae774c8_77, \3212 );
nor \U$25612 ( \25989 , \25987 , \25988 );
not \U$25613 ( \25990 , \25989 );
or \U$25614 ( \25991 , \25986 , \25990 );
or \U$25615 ( \25992 , \25989 , \3218 );
nand \U$25616 ( \25993 , \25991 , \25992 );
and \U$25617 ( \25994 , \5896 , RIae76d48_61);
and \U$25618 ( \25995 , RIae76c58_59, \5894 );
nor \U$25619 ( \25996 , \25994 , \25995 );
and \U$25620 ( \25997 , \25996 , \5590 );
not \U$25621 ( \25998 , \25996 );
and \U$25622 ( \25999 , \25998 , \5589 );
nor \U$25623 ( \26000 , \25997 , \25999 );
and \U$25624 ( \26001 , \5399 , RIae76f28_65);
and \U$25625 ( \26002 , RIae76e38_63, \5397 );
nor \U$25626 ( \26003 , \26001 , \26002 );
and \U$25627 ( \26004 , \26003 , \5016 );
not \U$25628 ( \26005 , \26003 );
and \U$25629 ( \26006 , \26005 , \5403 );
nor \U$25630 ( \26007 , \26004 , \26006 );
xor \U$25631 ( \26008 , \26000 , \26007 );
and \U$25632 ( \26009 , \6172 , RIae77180_70);
and \U$25633 ( \26010 , RIae77018_67, \6170 );
nor \U$25634 ( \26011 , \26009 , \26010 );
and \U$25635 ( \26012 , \26011 , \6176 );
not \U$25636 ( \26013 , \26011 );
and \U$25637 ( \26014 , \26013 , \6175 );
nor \U$25638 ( \26015 , \26012 , \26014 );
xor \U$25639 ( \26016 , \26008 , \26015 );
and \U$25640 ( \26017 , \25993 , \26016 );
and \U$25641 ( \26018 , \3730 , RIae77720_82);
and \U$25642 ( \26019 , RIae773d8_75, \3728 );
nor \U$25643 ( \26020 , \26018 , \26019 );
and \U$25644 ( \26021 , \26020 , \3732 );
not \U$25645 ( \26022 , \26020 );
and \U$25646 ( \26023 , \26022 , \3422 );
nor \U$25647 ( \26024 , \26021 , \26023 );
and \U$25648 ( \26025 , \4247 , RIae77a68_89);
and \U$25649 ( \26026 , RIae77978_87, \4245 );
nor \U$25650 ( \26027 , \26025 , \26026 );
and \U$25651 ( \26028 , \26027 , \3989 );
not \U$25652 ( \26029 , \26027 );
and \U$25653 ( \26030 , \26029 , \4251 );
nor \U$25654 ( \26031 , \26028 , \26030 );
xor \U$25655 ( \26032 , \26024 , \26031 );
and \U$25656 ( \26033 , \4688 , RIae77798_83);
and \U$25657 ( \26034 , RIae77888_85, \4686 );
nor \U$25658 ( \26035 , \26033 , \26034 );
and \U$25659 ( \26036 , \26035 , \4481 );
not \U$25660 ( \26037 , \26035 );
and \U$25661 ( \26038 , \26037 , \4482 );
nor \U$25662 ( \26039 , \26036 , \26038 );
xor \U$25663 ( \26040 , \26032 , \26039 );
xor \U$25664 ( \26041 , \26000 , \26007 );
xor \U$25665 ( \26042 , \26041 , \26015 );
and \U$25666 ( \26043 , \26040 , \26042 );
and \U$25667 ( \26044 , \25993 , \26040 );
or \U$25668 ( \26045 , \26017 , \26043 , \26044 );
and \U$25669 ( \26046 , \25985 , \26045 );
and \U$25670 ( \26047 , \25908 , \25984 );
or \U$25671 ( \26048 , \26046 , \26047 );
xor \U$25672 ( \26049 , \25829 , \26048 );
xor \U$25673 ( \26050 , \25770 , \25777 );
and \U$25674 ( \26051 , \26050 , \25785 );
and \U$25675 ( \26052 , \25770 , \25777 );
or \U$25676 ( \26053 , \26051 , \26052 );
and \U$25677 ( \26054 , \15726 , RIae75f38_31);
and \U$25678 ( \26055 , RIae7aab0_192, RIae75e48_29);
nor \U$25679 ( \26056 , \26054 , \26055 );
and \U$25680 ( \26057 , \26056 , RIae7aa38_191);
not \U$25681 ( \26058 , \26056 );
and \U$25682 ( \26059 , \26058 , \14959 );
nor \U$25683 ( \26060 , \26057 , \26059 );
and \U$25684 ( \26061 , \14964 , RIae75998_19);
and \U$25685 ( \26062 , RIae758a8_17, \14962 );
nor \U$25686 ( \26063 , \26061 , \26062 );
and \U$25687 ( \26064 , \26063 , \14462 );
not \U$25688 ( \26065 , \26063 );
and \U$25689 ( \26066 , \26065 , \14463 );
nor \U$25690 ( \26067 , \26064 , \26066 );
xor \U$25691 ( \26068 , \26060 , \26067 );
and \U$25692 ( \26069 , \14059 , RIae75b78_23);
and \U$25693 ( \26070 , RIae75a88_21, \14057 );
nor \U$25694 ( \26071 , \26069 , \26070 );
and \U$25695 ( \26072 , \26071 , \14063 );
not \U$25696 ( \26073 , \26071 );
and \U$25697 ( \26074 , \26073 , \13502 );
nor \U$25698 ( \26075 , \26072 , \26074 );
and \U$25699 ( \26076 , \26068 , \26075 );
and \U$25700 ( \26077 , \26060 , \26067 );
nor \U$25701 ( \26078 , \26076 , \26077 );
xor \U$25702 ( \26079 , \26053 , \26078 );
xor \U$25703 ( \26080 , \25794 , \25801 );
and \U$25704 ( \26081 , \26080 , \25809 );
and \U$25705 ( \26082 , \25794 , \25801 );
or \U$25706 ( \26083 , \26081 , \26082 );
xor \U$25707 ( \26084 , \26079 , \26083 );
xor \U$25708 ( \26085 , \25747 , \25754 );
and \U$25709 ( \26086 , \26085 , \25762 );
and \U$25710 ( \26087 , \25747 , \25754 );
or \U$25711 ( \26088 , \26086 , \26087 );
xor \U$25712 ( \26089 , \26000 , \26007 );
and \U$25713 ( \26090 , \26089 , \26015 );
and \U$25714 ( \26091 , \26000 , \26007 );
or \U$25715 ( \26092 , \26090 , \26091 );
xor \U$25716 ( \26093 , \26088 , \26092 );
xor \U$25717 ( \26094 , \26024 , \26031 );
and \U$25718 ( \26095 , \26094 , \26039 );
and \U$25719 ( \26096 , \26024 , \26031 );
or \U$25720 ( \26097 , \26095 , \26096 );
xor \U$25721 ( \26098 , \26093 , \26097 );
and \U$25722 ( \26099 , \26084 , \26098 );
xor \U$25723 ( \26100 , \25628 , \25635 );
xor \U$25724 ( \26101 , \26100 , \25643 );
xor \U$25725 ( \26102 , \25575 , \25581 );
xor \U$25726 ( \26103 , \26102 , \25589 );
xor \U$25727 ( \26104 , \25603 , \25610 );
xor \U$25728 ( \26105 , \26104 , \25618 );
xor \U$25729 ( \26106 , \26103 , \26105 );
xor \U$25730 ( \26107 , \26101 , \26106 );
xor \U$25731 ( \26108 , \26088 , \26092 );
xor \U$25732 ( \26109 , \26108 , \26097 );
and \U$25733 ( \26110 , \26107 , \26109 );
and \U$25734 ( \26111 , \26084 , \26107 );
or \U$25735 ( \26112 , \26099 , \26110 , \26111 );
and \U$25736 ( \26113 , \26049 , \26112 );
and \U$25737 ( \26114 , \25829 , \26048 );
or \U$25738 ( \26115 , \26113 , \26114 );
xor \U$25739 ( \26116 , \25460 , \25462 );
xor \U$25740 ( \26117 , \26116 , \25475 );
xor \U$25741 ( \26118 , \26115 , \26117 );
xor \U$25742 ( \26119 , \25503 , \25521 );
xor \U$25743 ( \26120 , \26119 , \25547 );
xor \U$25744 ( \26121 , \25558 , \25566 );
xor \U$25745 ( \26122 , \26121 , \25592 );
xor \U$25746 ( \26123 , \25621 , \25646 );
xor \U$25747 ( \26124 , \26123 , \25672 );
xor \U$25748 ( \26125 , \26122 , \26124 );
xor \U$25749 ( \26126 , \26120 , \26125 );
xor \U$25750 ( \26127 , \26088 , \26092 );
and \U$25751 ( \26128 , \26127 , \26097 );
and \U$25752 ( \26129 , \26088 , \26092 );
or \U$25753 ( \26130 , \26128 , \26129 );
xor \U$25754 ( \26131 , \26053 , \26078 );
and \U$25755 ( \26132 , \26131 , \26083 );
and \U$25756 ( \26133 , \26053 , \26078 );
or \U$25757 ( \26134 , \26132 , \26133 );
xor \U$25758 ( \26135 , \26130 , \26134 );
xor \U$25759 ( \26136 , \25628 , \25635 );
xor \U$25760 ( \26137 , \26136 , \25643 );
and \U$25761 ( \26138 , \26103 , \26137 );
xor \U$25762 ( \26139 , \25628 , \25635 );
xor \U$25763 ( \26140 , \26139 , \25643 );
and \U$25764 ( \26141 , \26105 , \26140 );
and \U$25765 ( \26142 , \26103 , \26105 );
or \U$25766 ( \26143 , \26138 , \26141 , \26142 );
xor \U$25767 ( \26144 , \26135 , \26143 );
and \U$25768 ( \26145 , \26126 , \26144 );
xor \U$25769 ( \26146 , \25452 , \25454 );
xor \U$25770 ( \26147 , \26146 , \25457 );
xor \U$25771 ( \26148 , \25529 , \25536 );
xor \U$25772 ( \26149 , \26148 , \25544 );
and \U$25773 ( \26150 , \25822 , \26149 );
xor \U$25774 ( \26151 , \25529 , \25536 );
xor \U$25775 ( \26152 , \26151 , \25544 );
and \U$25776 ( \26153 , \25824 , \26152 );
and \U$25777 ( \26154 , \25822 , \25824 );
or \U$25778 ( \26155 , \26150 , \26153 , \26154 );
xor \U$25779 ( \26156 , \25277 , \25284 );
xor \U$25780 ( \26157 , \26156 , \25292 );
xor \U$25781 ( \26158 , \25465 , \25470 );
xor \U$25782 ( \26159 , \26157 , \26158 );
xor \U$25783 ( \26160 , \26155 , \26159 );
xor \U$25784 ( \26161 , \26147 , \26160 );
xor \U$25785 ( \26162 , \26130 , \26134 );
xor \U$25786 ( \26163 , \26162 , \26143 );
and \U$25787 ( \26164 , \26161 , \26163 );
and \U$25788 ( \26165 , \26126 , \26161 );
or \U$25789 ( \26166 , \26145 , \26164 , \26165 );
and \U$25790 ( \26167 , \26118 , \26166 );
and \U$25791 ( \26168 , \26115 , \26117 );
or \U$25792 ( \26169 , \26167 , \26168 );
xor \U$25793 ( \26170 , \25478 , \25678 );
xor \U$25794 ( \26171 , \26170 , \25693 );
xor \U$25795 ( \26172 , \26169 , \26171 );
xor \U$25796 ( \26173 , \25550 , \25595 );
xor \U$25797 ( \26174 , \26173 , \25675 );
xor \U$25798 ( \26175 , \25323 , \25348 );
xor \U$25799 ( \26176 , \26175 , \25374 );
xor \U$25800 ( \26177 , \25244 , \25269 );
xor \U$25801 ( \26178 , \26177 , \25295 );
xor \U$25802 ( \26179 , \26176 , \26178 );
xor \U$25803 ( \26180 , \25380 , \25385 );
xor \U$25804 ( \26181 , \26180 , \25388 );
xor \U$25805 ( \26182 , \25681 , \25688 );
xor \U$25806 ( \26183 , \26181 , \26182 );
xor \U$25807 ( \26184 , \26179 , \26183 );
and \U$25808 ( \26185 , \26174 , \26184 );
xor \U$25809 ( \26186 , \25503 , \25521 );
xor \U$25810 ( \26187 , \26186 , \25547 );
and \U$25811 ( \26188 , \26122 , \26187 );
xor \U$25812 ( \26189 , \25503 , \25521 );
xor \U$25813 ( \26190 , \26189 , \25547 );
and \U$25814 ( \26191 , \26124 , \26190 );
and \U$25815 ( \26192 , \26122 , \26124 );
or \U$25816 ( \26193 , \26188 , \26191 , \26192 );
xor \U$25817 ( \26194 , \26130 , \26134 );
and \U$25818 ( \26195 , \26194 , \26143 );
and \U$25819 ( \26196 , \26130 , \26134 );
or \U$25820 ( \26197 , \26195 , \26196 );
xor \U$25821 ( \26198 , \26193 , \26197 );
xor \U$25822 ( \26199 , \25452 , \25454 );
xor \U$25823 ( \26200 , \26199 , \25457 );
and \U$25824 ( \26201 , \26155 , \26200 );
xor \U$25825 ( \26202 , \25452 , \25454 );
xor \U$25826 ( \26203 , \26202 , \25457 );
and \U$25827 ( \26204 , \26159 , \26203 );
and \U$25828 ( \26205 , \26155 , \26159 );
or \U$25829 ( \26206 , \26201 , \26204 , \26205 );
xor \U$25830 ( \26207 , \26198 , \26206 );
xor \U$25831 ( \26208 , \26176 , \26178 );
xor \U$25832 ( \26209 , \26208 , \26183 );
and \U$25833 ( \26210 , \26207 , \26209 );
and \U$25834 ( \26211 , \26174 , \26207 );
or \U$25835 ( \26212 , \26185 , \26210 , \26211 );
and \U$25836 ( \26213 , \26172 , \26212 );
and \U$25837 ( \26214 , \26169 , \26171 );
or \U$25838 ( \26215 , \26213 , \26214 );
not \U$25839 ( \26216 , \26215 );
xor \U$25840 ( \26217 , \26193 , \26197 );
and \U$25841 ( \26218 , \26217 , \26206 );
and \U$25842 ( \26219 , \26193 , \26197 );
or \U$25843 ( \26220 , \26218 , \26219 );
xor \U$25844 ( \26221 , \26176 , \26178 );
and \U$25845 ( \26222 , \26221 , \26183 );
and \U$25846 ( \26223 , \26176 , \26178 );
or \U$25847 ( \26224 , \26222 , \26223 );
xor \U$25848 ( \26225 , \26220 , \26224 );
xor \U$25849 ( \26226 , \25209 , \25211 );
xor \U$25850 ( \26227 , \26226 , \25216 );
xor \U$25851 ( \26228 , \25701 , \25706 );
xor \U$25852 ( \26229 , \26227 , \26228 );
and \U$25853 ( \26230 , \26225 , \26229 );
and \U$25854 ( \26231 , \26220 , \26224 );
or \U$25855 ( \26232 , \26230 , \26231 );
xor \U$25856 ( \26233 , \25696 , \25698 );
xor \U$25857 ( \26234 , \26233 , \25711 );
xnor \U$25858 ( \26235 , \26232 , \26234 );
not \U$25859 ( \26236 , \26235 );
xor \U$25860 ( \26237 , \25716 , \25720 );
not \U$25861 ( \26238 , \26237 );
and \U$25862 ( \26239 , \26236 , \26238 );
and \U$25863 ( \26240 , \26235 , \26237 );
nor \U$25864 ( \26241 , \26239 , \26240 );
not \U$25865 ( \26242 , \26241 );
or \U$25866 ( \26243 , \26216 , \26242 );
or \U$25867 ( \26244 , \26241 , \26215 );
nand \U$25868 ( \26245 , \26243 , \26244 );
xor \U$25869 ( \26246 , \26220 , \26224 );
xor \U$25870 ( \26247 , \26246 , \26229 );
not \U$25871 ( \26248 , \26247 );
xor \U$25872 ( \26249 , \26169 , \26171 );
xor \U$25873 ( \26250 , \26249 , \26212 );
not \U$25874 ( \26251 , \26250 );
or \U$25875 ( \26252 , \26248 , \26251 );
or \U$25876 ( \26253 , \26250 , \26247 );
xor \U$25877 ( \26254 , \26115 , \26117 );
xor \U$25878 ( \26255 , \26254 , \26166 );
not \U$25879 ( \26256 , \26255 );
xor \U$25880 ( \26257 , \26176 , \26178 );
xor \U$25881 ( \26258 , \26257 , \26183 );
xor \U$25882 ( \26259 , \26174 , \26207 );
xor \U$25883 ( \26260 , \26258 , \26259 );
not \U$25884 ( \26261 , \26260 );
or \U$25885 ( \26262 , \26256 , \26261 );
or \U$25886 ( \26263 , \26260 , \26255 );
xor \U$25887 ( \26264 , \25908 , \25984 );
xor \U$25888 ( \26265 , \26264 , \26045 );
xor \U$25889 ( \26266 , \25815 , \25817 );
xor \U$25890 ( \26267 , \26266 , \25826 );
and \U$25891 ( \26268 , \26265 , \26267 );
xor \U$25892 ( \26269 , \26088 , \26092 );
xor \U$25893 ( \26270 , \26269 , \26097 );
xor \U$25894 ( \26271 , \26084 , \26107 );
xor \U$25895 ( \26272 , \26270 , \26271 );
xor \U$25896 ( \26273 , \25815 , \25817 );
xor \U$25897 ( \26274 , \26273 , \25826 );
and \U$25898 ( \26275 , \26272 , \26274 );
and \U$25899 ( \26276 , \26265 , \26272 );
or \U$25900 ( \26277 , \26268 , \26275 , \26276 );
xor \U$25901 ( \26278 , \25934 , \25941 );
xor \U$25902 ( \26279 , \26278 , \25949 );
not \U$25903 ( \26280 , \26279 );
xor \U$25904 ( \26281 , \25915 , \3218 );
xor \U$25905 ( \26282 , \26281 , \25923 );
nand \U$25906 ( \26283 , \26280 , \26282 );
xor \U$25907 ( \26284 , \26060 , \26067 );
xor \U$25908 ( \26285 , \26284 , \26075 );
xor \U$25909 ( \26286 , \26283 , \26285 );
xor \U$25910 ( \26287 , \25861 , \25868 );
xor \U$25911 ( \26288 , \26287 , \25876 );
not \U$25912 ( \26289 , \26288 );
not \U$25913 ( \26290 , \25969 );
not \U$25914 ( \26291 , \25980 );
or \U$25915 ( \26292 , \26290 , \26291 );
or \U$25916 ( \26293 , \25969 , \25980 );
nand \U$25917 ( \26294 , \26292 , \26293 );
not \U$25918 ( \26295 , \26294 );
not \U$25919 ( \26296 , \25962 );
and \U$25920 ( \26297 , \26295 , \26296 );
and \U$25921 ( \26298 , \26294 , \25962 );
nor \U$25922 ( \26299 , \26297 , \26298 );
not \U$25923 ( \26300 , \26299 );
and \U$25924 ( \26301 , \26289 , \26300 );
and \U$25925 ( \26302 , \26299 , \26288 );
xor \U$25926 ( \26303 , \25836 , \25843 );
xor \U$25927 ( \26304 , \26303 , \25851 );
nor \U$25928 ( \26305 , \26302 , \26304 );
nor \U$25929 ( \26306 , \26301 , \26305 );
and \U$25930 ( \26307 , \26286 , \26306 );
and \U$25931 ( \26308 , \26283 , \26285 );
or \U$25932 ( \26309 , \26307 , \26308 );
and \U$25933 ( \26310 , \12180 , RIae77d38_95);
and \U$25934 ( \26311 , RIae77e28_97, \12178 );
nor \U$25935 ( \26312 , \26310 , \26311 );
and \U$25936 ( \26313 , \26312 , \12184 );
not \U$25937 ( \26314 , \26312 );
and \U$25938 ( \26315 , \26314 , \11827 );
nor \U$25939 ( \26316 , \26313 , \26315 );
and \U$25940 ( \26317 , \11470 , RIae77c48_93);
and \U$25941 ( \26318 , RIae77b58_91, \11468 );
nor \U$25942 ( \26319 , \26317 , \26318 );
and \U$25943 ( \26320 , \26319 , \10936 );
not \U$25944 ( \26321 , \26319 );
and \U$25945 ( \26322 , \26321 , \11474 );
nor \U$25946 ( \26323 , \26320 , \26322 );
xor \U$25947 ( \26324 , \26316 , \26323 );
and \U$25948 ( \26325 , \13059 , RIae78968_121);
and \U$25949 ( \26326 , RIae78878_119, \13057 );
nor \U$25950 ( \26327 , \26325 , \26326 );
and \U$25951 ( \26328 , \26327 , \13063 );
not \U$25952 ( \26329 , \26327 );
and \U$25953 ( \26330 , \26329 , \12718 );
nor \U$25954 ( \26331 , \26328 , \26330 );
and \U$25955 ( \26332 , \26324 , \26331 );
and \U$25956 ( \26333 , \26316 , \26323 );
or \U$25957 ( \26334 , \26332 , \26333 );
and \U$25958 ( \26335 , \14059 , RIae78788_117);
and \U$25959 ( \26336 , RIae78698_115, \14057 );
nor \U$25960 ( \26337 , \26335 , \26336 );
and \U$25961 ( \26338 , \26337 , \13502 );
not \U$25962 ( \26339 , \26337 );
and \U$25963 ( \26340 , \26339 , \14063 );
nor \U$25964 ( \26341 , \26338 , \26340 );
and \U$25965 ( \26342 , \15726 , RIae75998_19);
and \U$25966 ( \26343 , RIae7aab0_192, RIae758a8_17);
nor \U$25967 ( \26344 , \26342 , \26343 );
and \U$25968 ( \26345 , \26344 , \14959 );
not \U$25969 ( \26346 , \26344 );
and \U$25970 ( \26347 , \26346 , RIae7aa38_191);
nor \U$25971 ( \26348 , \26345 , \26347 );
xor \U$25972 ( \26349 , \26341 , \26348 );
and \U$25973 ( \26350 , \14964 , RIae75b78_23);
and \U$25974 ( \26351 , RIae75a88_21, \14962 );
nor \U$25975 ( \26352 , \26350 , \26351 );
and \U$25976 ( \26353 , \26352 , \14463 );
not \U$25977 ( \26354 , \26352 );
and \U$25978 ( \26355 , \26354 , \14462 );
nor \U$25979 ( \26356 , \26353 , \26355 );
and \U$25980 ( \26357 , \26349 , \26356 );
and \U$25981 ( \26358 , \26341 , \26348 );
or \U$25982 ( \26359 , \26357 , \26358 );
xor \U$25983 ( \26360 , \26334 , \26359 );
and \U$25984 ( \26361 , \8966 , RIae77f18_99);
and \U$25985 ( \26362 , RIae78008_101, \8964 );
nor \U$25986 ( \26363 , \26361 , \26362 );
and \U$25987 ( \26364 , \26363 , \8799 );
not \U$25988 ( \26365 , \26363 );
and \U$25989 ( \26366 , \26365 , \8789 );
nor \U$25990 ( \26367 , \26364 , \26366 );
and \U$25991 ( \26368 , \9760 , RIae781e8_105);
and \U$25992 ( \26369 , RIae785a8_113, \9758 );
nor \U$25993 ( \26370 , \26368 , \26369 );
and \U$25994 ( \26371 , \26370 , \9273 );
not \U$25995 ( \26372 , \26370 );
and \U$25996 ( \26373 , \26372 , \9764 );
nor \U$25997 ( \26374 , \26371 , \26373 );
xor \U$25998 ( \26375 , \26367 , \26374 );
and \U$25999 ( \26376 , \10548 , RIae783c8_109);
and \U$26000 ( \26377 , RIae78530_112, \10546 );
nor \U$26001 ( \26378 , \26376 , \26377 );
and \U$26002 ( \26379 , \26378 , \10421 );
not \U$26003 ( \26380 , \26378 );
and \U$26004 ( \26381 , \26380 , \10118 );
nor \U$26005 ( \26382 , \26379 , \26381 );
and \U$26006 ( \26383 , \26375 , \26382 );
and \U$26007 ( \26384 , \26367 , \26374 );
or \U$26008 ( \26385 , \26383 , \26384 );
and \U$26009 ( \26386 , \26360 , \26385 );
and \U$26010 ( \26387 , \26334 , \26359 );
nor \U$26011 ( \26388 , \26386 , \26387 );
nand \U$26012 ( \26389 , RIae775b8_79, \3212 );
not \U$26013 ( \26390 , \26389 );
not \U$26014 ( \26391 , \2774 );
or \U$26015 ( \26392 , \26390 , \26391 );
or \U$26016 ( \26393 , \2774 , \26389 );
nand \U$26017 ( \26394 , \26392 , \26393 );
and \U$26018 ( \26395 , \3730 , RIae774c8_77);
and \U$26019 ( \26396 , RIae77720_82, \3728 );
nor \U$26020 ( \26397 , \26395 , \26396 );
and \U$26021 ( \26398 , \26397 , \3732 );
not \U$26022 ( \26399 , \26397 );
and \U$26023 ( \26400 , \26399 , \3422 );
nor \U$26024 ( \26401 , \26398 , \26400 );
xor \U$26025 ( \26402 , \26394 , \26401 );
xor \U$26026 ( \26403 , \25887 , \25894 );
xor \U$26027 ( \26404 , \26403 , \25902 );
and \U$26028 ( \26405 , \26402 , \26404 );
and \U$26029 ( \26406 , \26394 , \26401 );
nor \U$26030 ( \26407 , \26405 , \26406 );
xor \U$26031 ( \26408 , \26388 , \26407 );
and \U$26032 ( \26409 , \5399 , RIae77798_83);
and \U$26033 ( \26410 , RIae77888_85, \5397 );
nor \U$26034 ( \26411 , \26409 , \26410 );
and \U$26035 ( \26412 , \26411 , \5016 );
not \U$26036 ( \26413 , \26411 );
and \U$26037 ( \26414 , \26413 , \5403 );
nor \U$26038 ( \26415 , \26412 , \26414 );
and \U$26039 ( \26416 , \5896 , RIae76f28_65);
and \U$26040 ( \26417 , RIae76e38_63, \5894 );
nor \U$26041 ( \26418 , \26416 , \26417 );
and \U$26042 ( \26419 , \26418 , \5590 );
not \U$26043 ( \26420 , \26418 );
and \U$26044 ( \26421 , \26420 , \5589 );
nor \U$26045 ( \26422 , \26419 , \26421 );
xor \U$26046 ( \26423 , \26415 , \26422 );
and \U$26047 ( \26424 , \6172 , RIae76d48_61);
and \U$26048 ( \26425 , RIae76c58_59, \6170 );
nor \U$26049 ( \26426 , \26424 , \26425 );
and \U$26050 ( \26427 , \26426 , \6176 );
not \U$26051 ( \26428 , \26426 );
and \U$26052 ( \26429 , \26428 , \6175 );
nor \U$26053 ( \26430 , \26427 , \26429 );
and \U$26054 ( \26431 , \26423 , \26430 );
and \U$26055 ( \26432 , \26415 , \26422 );
or \U$26056 ( \26433 , \26431 , \26432 );
and \U$26057 ( \26434 , \4688 , RIae77a68_89);
and \U$26058 ( \26435 , RIae77978_87, \4686 );
nor \U$26059 ( \26436 , \26434 , \26435 );
and \U$26060 ( \26437 , \26436 , \4481 );
not \U$26061 ( \26438 , \26436 );
and \U$26062 ( \26439 , \26438 , \4482 );
nor \U$26063 ( \26440 , \26437 , \26439 );
and \U$26064 ( \26441 , \3730 , RIae775b8_79);
and \U$26065 ( \26442 , RIae774c8_77, \3728 );
nor \U$26066 ( \26443 , \26441 , \26442 );
and \U$26067 ( \26444 , \26443 , \3732 );
not \U$26068 ( \26445 , \26443 );
and \U$26069 ( \26446 , \26445 , \3422 );
nor \U$26070 ( \26447 , \26444 , \26446 );
xor \U$26071 ( \26448 , \26440 , \26447 );
and \U$26072 ( \26449 , \4247 , RIae77720_82);
and \U$26073 ( \26450 , RIae773d8_75, \4245 );
nor \U$26074 ( \26451 , \26449 , \26450 );
and \U$26075 ( \26452 , \26451 , \3989 );
not \U$26076 ( \26453 , \26451 );
and \U$26077 ( \26454 , \26453 , \4251 );
nor \U$26078 ( \26455 , \26452 , \26454 );
and \U$26079 ( \26456 , \26448 , \26455 );
and \U$26080 ( \26457 , \26440 , \26447 );
or \U$26081 ( \26458 , \26456 , \26457 );
xor \U$26082 ( \26459 , \26433 , \26458 );
and \U$26083 ( \26460 , \6941 , RIae77180_70);
and \U$26084 ( \26461 , RIae77018_67, \6939 );
nor \U$26085 ( \26462 , \26460 , \26461 );
and \U$26086 ( \26463 , \26462 , \6314 );
not \U$26087 ( \26464 , \26462 );
and \U$26088 ( \26465 , \26464 , \6945 );
nor \U$26089 ( \26466 , \26463 , \26465 );
and \U$26090 ( \26467 , \7633 , RIae771f8_71);
and \U$26091 ( \26468 , RIae772e8_73, \7631 );
nor \U$26092 ( \26469 , \26467 , \26468 );
and \U$26093 ( \26470 , \26469 , \7206 );
not \U$26094 ( \26471 , \26469 );
and \U$26095 ( \26472 , \26471 , \7205 );
nor \U$26096 ( \26473 , \26470 , \26472 );
xor \U$26097 ( \26474 , \26466 , \26473 );
and \U$26098 ( \26475 , \8371 , RIae782d8_107);
and \U$26099 ( \26476 , RIae780f8_103, \8369 );
nor \U$26100 ( \26477 , \26475 , \26476 );
and \U$26101 ( \26478 , \26477 , \8020 );
not \U$26102 ( \26479 , \26477 );
and \U$26103 ( \26480 , \26479 , \8019 );
nor \U$26104 ( \26481 , \26478 , \26480 );
and \U$26105 ( \26482 , \26474 , \26481 );
and \U$26106 ( \26483 , \26466 , \26473 );
or \U$26107 ( \26484 , \26482 , \26483 );
and \U$26108 ( \26485 , \26459 , \26484 );
and \U$26109 ( \26486 , \26433 , \26458 );
nor \U$26110 ( \26487 , \26485 , \26486 );
and \U$26111 ( \26488 , \26408 , \26487 );
and \U$26112 ( \26489 , \26388 , \26407 );
or \U$26113 ( \26490 , \26488 , \26489 );
xor \U$26114 ( \26491 , \26309 , \26490 );
xor \U$26115 ( \26492 , \25770 , \25777 );
xor \U$26116 ( \26493 , \26492 , \25785 );
xor \U$26117 ( \26494 , \25763 , \25810 );
xor \U$26118 ( \26495 , \26493 , \26494 );
xor \U$26119 ( \26496 , \25854 , \25879 );
xor \U$26120 ( \26497 , \26496 , \25905 );
xor \U$26121 ( \26498 , \26495 , \26497 );
xor \U$26122 ( \26499 , \26000 , \26007 );
xor \U$26123 ( \26500 , \26499 , \26015 );
xor \U$26124 ( \26501 , \25993 , \26040 );
xor \U$26125 ( \26502 , \26500 , \26501 );
and \U$26126 ( \26503 , \26498 , \26502 );
and \U$26127 ( \26504 , \26495 , \26497 );
nor \U$26128 ( \26505 , \26503 , \26504 );
and \U$26129 ( \26506 , \26491 , \26505 );
and \U$26130 ( \26507 , \26309 , \26490 );
nor \U$26131 ( \26508 , \26506 , \26507 );
xor \U$26132 ( \26509 , \26277 , \26508 );
xor \U$26133 ( \26510 , \26130 , \26134 );
xor \U$26134 ( \26511 , \26510 , \26143 );
xor \U$26135 ( \26512 , \26126 , \26161 );
xor \U$26136 ( \26513 , \26511 , \26512 );
and \U$26137 ( \26514 , \26509 , \26513 );
and \U$26138 ( \26515 , \26277 , \26508 );
or \U$26139 ( \26516 , \26514 , \26515 );
nand \U$26140 ( \26517 , \26263 , \26516 );
nand \U$26141 ( \26518 , \26262 , \26517 );
nand \U$26142 ( \26519 , \26253 , \26518 );
nand \U$26143 ( \26520 , \26252 , \26519 );
and \U$26144 ( \26521 , \26245 , \26520 );
xor \U$26145 ( \26522 , \26520 , \26245 );
xnor \U$26146 ( \26523 , \26518 , \26250 );
not \U$26147 ( \26524 , \26523 );
not \U$26148 ( \26525 , \26247 );
and \U$26149 ( \26526 , \26524 , \26525 );
and \U$26150 ( \26527 , \26523 , \26247 );
nor \U$26151 ( \26528 , \26526 , \26527 );
xnor \U$26152 ( \26529 , \26516 , \26255 );
not \U$26153 ( \26530 , \26529 );
not \U$26154 ( \26531 , \26260 );
and \U$26155 ( \26532 , \26530 , \26531 );
and \U$26156 ( \26533 , \26529 , \26260 );
nor \U$26157 ( \26534 , \26532 , \26533 );
not \U$26158 ( \26535 , \26534 );
xor \U$26159 ( \26536 , \26283 , \26285 );
xor \U$26160 ( \26537 , \26536 , \26306 );
xnor \U$26161 ( \26538 , \25952 , \25982 );
not \U$26162 ( \26539 , \26538 );
not \U$26163 ( \26540 , \25926 );
and \U$26164 ( \26541 , \26539 , \26540 );
and \U$26165 ( \26542 , \26538 , \25926 );
nor \U$26166 ( \26543 , \26541 , \26542 );
or \U$26167 ( \26544 , \26537 , \26543 );
not \U$26168 ( \26545 , \26543 );
not \U$26169 ( \26546 , \26537 );
or \U$26170 ( \26547 , \26545 , \26546 );
xor \U$26171 ( \26548 , \26495 , \26497 );
xor \U$26172 ( \26549 , \26548 , \26502 );
nand \U$26173 ( \26550 , \26547 , \26549 );
nand \U$26174 ( \26551 , \26544 , \26550 );
xor \U$26175 ( \26552 , \26334 , \26359 );
xor \U$26176 ( \26553 , \26552 , \26385 );
xor \U$26177 ( \26554 , \26394 , \26401 );
xor \U$26178 ( \26555 , \26554 , \26404 );
xor \U$26179 ( \26556 , \26553 , \26555 );
xor \U$26180 ( \26557 , \26433 , \26458 );
xor \U$26181 ( \26558 , \26557 , \26484 );
and \U$26182 ( \26559 , \26556 , \26558 );
and \U$26183 ( \26560 , \26553 , \26555 );
or \U$26184 ( \26561 , \26559 , \26560 );
and \U$26185 ( \26562 , \6941 , RIae76c58_59);
and \U$26186 ( \26563 , RIae77180_70, \6939 );
nor \U$26187 ( \26564 , \26562 , \26563 );
and \U$26188 ( \26565 , \26564 , \6945 );
not \U$26189 ( \26566 , \26564 );
and \U$26190 ( \26567 , \26566 , \6314 );
nor \U$26191 ( \26568 , \26565 , \26567 );
and \U$26192 ( \26569 , \5896 , RIae77888_85);
and \U$26193 ( \26570 , RIae76f28_65, \5894 );
nor \U$26194 ( \26571 , \26569 , \26570 );
and \U$26195 ( \26572 , \26571 , \5589 );
not \U$26196 ( \26573 , \26571 );
and \U$26197 ( \26574 , \26573 , \5590 );
nor \U$26198 ( \26575 , \26572 , \26574 );
xor \U$26199 ( \26576 , \26568 , \26575 );
and \U$26200 ( \26577 , \6172 , RIae76e38_63);
and \U$26201 ( \26578 , RIae76d48_61, \6170 );
nor \U$26202 ( \26579 , \26577 , \26578 );
and \U$26203 ( \26580 , \26579 , \6175 );
not \U$26204 ( \26581 , \26579 );
and \U$26205 ( \26582 , \26581 , \6176 );
nor \U$26206 ( \26583 , \26580 , \26582 );
and \U$26207 ( \26584 , \26576 , \26583 );
and \U$26208 ( \26585 , \26568 , \26575 );
or \U$26209 ( \26586 , \26584 , \26585 );
and \U$26210 ( \26587 , \7633 , RIae77018_67);
and \U$26211 ( \26588 , RIae771f8_71, \7631 );
nor \U$26212 ( \26589 , \26587 , \26588 );
and \U$26213 ( \26590 , \26589 , \7205 );
not \U$26214 ( \26591 , \26589 );
and \U$26215 ( \26592 , \26591 , \7206 );
nor \U$26216 ( \26593 , \26590 , \26592 );
not \U$26217 ( \26594 , \26593 );
and \U$26218 ( \26595 , \8966 , RIae780f8_103);
and \U$26219 ( \26596 , RIae77f18_99, \8964 );
nor \U$26220 ( \26597 , \26595 , \26596 );
and \U$26221 ( \26598 , \26597 , \8789 );
not \U$26222 ( \26599 , \26597 );
and \U$26223 ( \26600 , \26599 , \8799 );
nor \U$26224 ( \26601 , \26598 , \26600 );
not \U$26225 ( \26602 , \26601 );
and \U$26226 ( \26603 , \26594 , \26602 );
and \U$26227 ( \26604 , \26601 , \26593 );
and \U$26228 ( \26605 , \8371 , RIae772e8_73);
and \U$26229 ( \26606 , RIae782d8_107, \8369 );
nor \U$26230 ( \26607 , \26605 , \26606 );
and \U$26231 ( \26608 , \26607 , \8019 );
not \U$26232 ( \26609 , \26607 );
and \U$26233 ( \26610 , \26609 , \8020 );
nor \U$26234 ( \26611 , \26608 , \26610 );
nor \U$26235 ( \26612 , \26604 , \26611 );
nor \U$26236 ( \26613 , \26603 , \26612 );
xor \U$26237 ( \26614 , \26586 , \26613 );
and \U$26238 ( \26615 , \4247 , RIae774c8_77);
and \U$26239 ( \26616 , RIae77720_82, \4245 );
nor \U$26240 ( \26617 , \26615 , \26616 );
and \U$26241 ( \26618 , \26617 , \4251 );
not \U$26242 ( \26619 , \26617 );
and \U$26243 ( \26620 , \26619 , \3989 );
nor \U$26244 ( \26621 , \26618 , \26620 );
and \U$26245 ( \26622 , \4688 , RIae773d8_75);
and \U$26246 ( \26623 , RIae77a68_89, \4686 );
nor \U$26247 ( \26624 , \26622 , \26623 );
and \U$26248 ( \26625 , \26624 , \4482 );
not \U$26249 ( \26626 , \26624 );
and \U$26250 ( \26627 , \26626 , \4481 );
nor \U$26251 ( \26628 , \26625 , \26627 );
xor \U$26252 ( \26629 , \26621 , \26628 );
and \U$26253 ( \26630 , \5399 , RIae77978_87);
and \U$26254 ( \26631 , RIae77798_83, \5397 );
nor \U$26255 ( \26632 , \26630 , \26631 );
and \U$26256 ( \26633 , \26632 , \5403 );
not \U$26257 ( \26634 , \26632 );
and \U$26258 ( \26635 , \26634 , \5016 );
nor \U$26259 ( \26636 , \26633 , \26635 );
and \U$26260 ( \26637 , \26629 , \26636 );
and \U$26261 ( \26638 , \26621 , \26628 );
or \U$26262 ( \26639 , \26637 , \26638 );
and \U$26263 ( \26640 , \26614 , \26639 );
and \U$26264 ( \26641 , \26586 , \26613 );
nor \U$26265 ( \26642 , \26640 , \26641 );
and \U$26266 ( \26643 , \14059 , RIae78878_119);
and \U$26267 ( \26644 , RIae78788_117, \14057 );
nor \U$26268 ( \26645 , \26643 , \26644 );
and \U$26269 ( \26646 , \26645 , \13502 );
not \U$26270 ( \26647 , \26645 );
and \U$26271 ( \26648 , \26647 , \14063 );
nor \U$26272 ( \26649 , \26646 , \26648 );
and \U$26273 ( \26650 , \12180 , RIae77b58_91);
and \U$26274 ( \26651 , RIae77d38_95, \12178 );
nor \U$26275 ( \26652 , \26650 , \26651 );
and \U$26276 ( \26653 , \26652 , \12184 );
not \U$26277 ( \26654 , \26652 );
and \U$26278 ( \26655 , \26654 , \11827 );
nor \U$26279 ( \26656 , \26653 , \26655 );
xor \U$26280 ( \26657 , \26649 , \26656 );
and \U$26281 ( \26658 , \13059 , RIae77e28_97);
and \U$26282 ( \26659 , RIae78968_121, \13057 );
nor \U$26283 ( \26660 , \26658 , \26659 );
and \U$26284 ( \26661 , \26660 , \13063 );
not \U$26285 ( \26662 , \26660 );
and \U$26286 ( \26663 , \26662 , \12718 );
nor \U$26287 ( \26664 , \26661 , \26663 );
and \U$26288 ( \26665 , \26657 , \26664 );
and \U$26289 ( \26666 , \26649 , \26656 );
or \U$26290 ( \26667 , \26665 , \26666 );
and \U$26291 ( \26668 , \15726 , RIae75a88_21);
and \U$26292 ( \26669 , RIae7aab0_192, RIae75998_19);
nor \U$26293 ( \26670 , \26668 , \26669 );
and \U$26294 ( \26671 , \26670 , \14959 );
not \U$26295 ( \26672 , \26670 );
and \U$26296 ( \26673 , \26672 , RIae7aa38_191);
nor \U$26297 ( \26674 , \26671 , \26673 );
xor \U$26298 ( \26675 , \26674 , \3422 );
and \U$26299 ( \26676 , \14964 , RIae78698_115);
and \U$26300 ( \26677 , RIae75b78_23, \14962 );
nor \U$26301 ( \26678 , \26676 , \26677 );
and \U$26302 ( \26679 , \26678 , \14463 );
not \U$26303 ( \26680 , \26678 );
and \U$26304 ( \26681 , \26680 , \14462 );
nor \U$26305 ( \26682 , \26679 , \26681 );
and \U$26306 ( \26683 , \26675 , \26682 );
and \U$26307 ( \26684 , \26674 , \3422 );
or \U$26308 ( \26685 , \26683 , \26684 );
xor \U$26309 ( \26686 , \26667 , \26685 );
and \U$26310 ( \26687 , \11470 , RIae78530_112);
and \U$26311 ( \26688 , RIae77c48_93, \11468 );
nor \U$26312 ( \26689 , \26687 , \26688 );
and \U$26313 ( \26690 , \26689 , \10936 );
not \U$26314 ( \26691 , \26689 );
and \U$26315 ( \26692 , \26691 , \11474 );
nor \U$26316 ( \26693 , \26690 , \26692 );
and \U$26317 ( \26694 , \9760 , RIae78008_101);
and \U$26318 ( \26695 , RIae781e8_105, \9758 );
nor \U$26319 ( \26696 , \26694 , \26695 );
and \U$26320 ( \26697 , \26696 , \9273 );
not \U$26321 ( \26698 , \26696 );
and \U$26322 ( \26699 , \26698 , \9764 );
nor \U$26323 ( \26700 , \26697 , \26699 );
xor \U$26324 ( \26701 , \26693 , \26700 );
and \U$26325 ( \26702 , \10548 , RIae785a8_113);
and \U$26326 ( \26703 , RIae783c8_109, \10546 );
nor \U$26327 ( \26704 , \26702 , \26703 );
and \U$26328 ( \26705 , \26704 , \10421 );
not \U$26329 ( \26706 , \26704 );
and \U$26330 ( \26707 , \26706 , \10118 );
nor \U$26331 ( \26708 , \26705 , \26707 );
and \U$26332 ( \26709 , \26701 , \26708 );
and \U$26333 ( \26710 , \26693 , \26700 );
or \U$26334 ( \26711 , \26709 , \26710 );
and \U$26335 ( \26712 , \26686 , \26711 );
and \U$26336 ( \26713 , \26667 , \26685 );
or \U$26337 ( \26714 , \26712 , \26713 );
xor \U$26338 ( \26715 , \26642 , \26714 );
xor \U$26339 ( \26716 , \26415 , \26422 );
xor \U$26340 ( \26717 , \26716 , \26430 );
xor \U$26341 ( \26718 , \26440 , \26447 );
xor \U$26342 ( \26719 , \26718 , \26455 );
xor \U$26343 ( \26720 , \26717 , \26719 );
xor \U$26344 ( \26721 , \26466 , \26473 );
xor \U$26345 ( \26722 , \26721 , \26481 );
and \U$26346 ( \26723 , \26720 , \26722 );
and \U$26347 ( \26724 , \26717 , \26719 );
or \U$26348 ( \26725 , \26723 , \26724 );
and \U$26349 ( \26726 , \26715 , \26725 );
and \U$26350 ( \26727 , \26642 , \26714 );
or \U$26351 ( \26728 , \26726 , \26727 );
xor \U$26352 ( \26729 , \26561 , \26728 );
xor \U$26353 ( \26730 , \26341 , \26348 );
xor \U$26354 ( \26731 , \26730 , \26356 );
xor \U$26355 ( \26732 , \26316 , \26323 );
xor \U$26356 ( \26733 , \26732 , \26331 );
and \U$26357 ( \26734 , \26731 , \26733 );
xor \U$26358 ( \26735 , \26367 , \26374 );
xor \U$26359 ( \26736 , \26735 , \26382 );
xor \U$26360 ( \26737 , \26316 , \26323 );
xor \U$26361 ( \26738 , \26737 , \26331 );
and \U$26362 ( \26739 , \26736 , \26738 );
and \U$26363 ( \26740 , \26731 , \26736 );
or \U$26364 ( \26741 , \26734 , \26739 , \26740 );
not \U$26365 ( \26742 , \26279 );
not \U$26366 ( \26743 , \26282 );
or \U$26367 ( \26744 , \26742 , \26743 );
or \U$26368 ( \26745 , \26282 , \26279 );
nand \U$26369 ( \26746 , \26744 , \26745 );
xor \U$26370 ( \26747 , \26741 , \26746 );
not \U$26371 ( \26748 , \26288 );
xor \U$26372 ( \26749 , \26304 , \26299 );
not \U$26373 ( \26750 , \26749 );
or \U$26374 ( \26751 , \26748 , \26750 );
or \U$26375 ( \26752 , \26749 , \26288 );
nand \U$26376 ( \26753 , \26751 , \26752 );
and \U$26377 ( \26754 , \26747 , \26753 );
and \U$26378 ( \26755 , \26741 , \26746 );
or \U$26379 ( \26756 , \26754 , \26755 );
and \U$26380 ( \26757 , \26729 , \26756 );
and \U$26381 ( \26758 , \26561 , \26728 );
or \U$26382 ( \26759 , \26757 , \26758 );
xor \U$26383 ( \26760 , \26551 , \26759 );
xor \U$26384 ( \26761 , \25815 , \25817 );
xor \U$26385 ( \26762 , \26761 , \25826 );
xor \U$26386 ( \26763 , \26265 , \26272 );
xor \U$26387 ( \26764 , \26762 , \26763 );
and \U$26388 ( \26765 , \26760 , \26764 );
and \U$26389 ( \26766 , \26551 , \26759 );
or \U$26390 ( \26767 , \26765 , \26766 );
xor \U$26391 ( \26768 , \25829 , \26048 );
xor \U$26392 ( \26769 , \26768 , \26112 );
xor \U$26393 ( \26770 , \26767 , \26769 );
xor \U$26394 ( \26771 , \26277 , \26508 );
xor \U$26395 ( \26772 , \26771 , \26513 );
and \U$26396 ( \26773 , \26770 , \26772 );
and \U$26397 ( \26774 , \26767 , \26769 );
or \U$26398 ( \26775 , \26773 , \26774 );
nand \U$26399 ( \26776 , \26535 , \26775 );
or \U$26400 ( \26777 , \26528 , \26776 );
xnor \U$26401 ( \26778 , \26776 , \26528 );
xor \U$26402 ( \26779 , \26767 , \26769 );
xor \U$26403 ( \26780 , \26779 , \26772 );
not \U$26404 ( \26781 , \26780 );
xnor \U$26405 ( \26782 , \26543 , \26537 );
not \U$26406 ( \26783 , \26782 );
not \U$26407 ( \26784 , \26549 );
and \U$26408 ( \26785 , \26783 , \26784 );
and \U$26409 ( \26786 , \26782 , \26549 );
nor \U$26410 ( \26787 , \26785 , \26786 );
not \U$26411 ( \26788 , \26787 );
xor \U$26412 ( \26789 , \26561 , \26728 );
xor \U$26413 ( \26790 , \26789 , \26756 );
nand \U$26414 ( \26791 , \26788 , \26790 );
xor \U$26415 ( \26792 , \26309 , \26490 );
xor \U$26416 ( \26793 , \26792 , \26505 );
xor \U$26417 ( \26794 , \26791 , \26793 );
xor \U$26418 ( \26795 , \26642 , \26714 );
xor \U$26419 ( \26796 , \26795 , \26725 );
xor \U$26420 ( \26797 , \26553 , \26555 );
xor \U$26421 ( \26798 , \26797 , \26558 );
and \U$26422 ( \26799 , \26796 , \26798 );
xor \U$26423 ( \26800 , \26741 , \26746 );
xor \U$26424 ( \26801 , \26800 , \26753 );
xor \U$26425 ( \26802 , \26553 , \26555 );
xor \U$26426 ( \26803 , \26802 , \26558 );
and \U$26427 ( \26804 , \26801 , \26803 );
and \U$26428 ( \26805 , \26796 , \26801 );
or \U$26429 ( \26806 , \26799 , \26804 , \26805 );
not \U$26430 ( \26807 , \26806 );
not \U$26431 ( \26808 , \26807 );
xor \U$26432 ( \26809 , \26388 , \26407 );
xor \U$26433 ( \26810 , \26809 , \26487 );
not \U$26434 ( \26811 , \26810 );
and \U$26435 ( \26812 , \26808 , \26811 );
and \U$26436 ( \26813 , \26807 , \26810 );
not \U$26437 ( \26814 , \26593 );
xor \U$26438 ( \26815 , \26611 , \26601 );
not \U$26439 ( \26816 , \26815 );
or \U$26440 ( \26817 , \26814 , \26816 );
or \U$26441 ( \26818 , \26815 , \26593 );
nand \U$26442 ( \26819 , \26817 , \26818 );
xor \U$26443 ( \26820 , \26649 , \26656 );
xor \U$26444 ( \26821 , \26820 , \26664 );
and \U$26445 ( \26822 , \26819 , \26821 );
xor \U$26446 ( \26823 , \26693 , \26700 );
xor \U$26447 ( \26824 , \26823 , \26708 );
xor \U$26448 ( \26825 , \26649 , \26656 );
xor \U$26449 ( \26826 , \26825 , \26664 );
and \U$26450 ( \26827 , \26824 , \26826 );
and \U$26451 ( \26828 , \26819 , \26824 );
or \U$26452 ( \26829 , \26822 , \26827 , \26828 );
xor \U$26453 ( \26830 , \26717 , \26719 );
xor \U$26454 ( \26831 , \26830 , \26722 );
and \U$26455 ( \26832 , \26829 , \26831 );
xor \U$26456 ( \26833 , \26316 , \26323 );
xor \U$26457 ( \26834 , \26833 , \26331 );
xor \U$26458 ( \26835 , \26731 , \26736 );
xor \U$26459 ( \26836 , \26834 , \26835 );
xor \U$26460 ( \26837 , \26717 , \26719 );
xor \U$26461 ( \26838 , \26837 , \26722 );
and \U$26462 ( \26839 , \26836 , \26838 );
and \U$26463 ( \26840 , \26829 , \26836 );
or \U$26464 ( \26841 , \26832 , \26839 , \26840 );
xor \U$26465 ( \26842 , \26586 , \26613 );
xor \U$26466 ( \26843 , \26842 , \26639 );
not \U$26467 ( \26844 , \26843 );
xor \U$26468 ( \26845 , \26667 , \26685 );
xor \U$26469 ( \26846 , \26845 , \26711 );
nand \U$26470 ( \26847 , \26844 , \26846 );
not \U$26471 ( \26848 , \26847 );
and \U$26472 ( \26849 , \26841 , \26848 );
not \U$26473 ( \26850 , \26841 );
not \U$26474 ( \26851 , \26848 );
and \U$26475 ( \26852 , \26850 , \26851 );
and \U$26476 ( \26853 , \14059 , RIae78968_121);
and \U$26477 ( \26854 , RIae78878_119, \14057 );
nor \U$26478 ( \26855 , \26853 , \26854 );
and \U$26479 ( \26856 , \26855 , \14063 );
not \U$26480 ( \26857 , \26855 );
and \U$26481 ( \26858 , \26857 , \13502 );
nor \U$26482 ( \26859 , \26856 , \26858 );
not \U$26483 ( \26860 , \26859 );
and \U$26484 ( \26861 , \15726 , RIae75b78_23);
and \U$26485 ( \26862 , RIae7aab0_192, RIae75a88_21);
nor \U$26486 ( \26863 , \26861 , \26862 );
and \U$26487 ( \26864 , \26863 , RIae7aa38_191);
not \U$26488 ( \26865 , \26863 );
and \U$26489 ( \26866 , \26865 , \14959 );
nor \U$26490 ( \26867 , \26864 , \26866 );
not \U$26491 ( \26868 , \26867 );
and \U$26492 ( \26869 , \26860 , \26868 );
and \U$26493 ( \26870 , \26859 , \26867 );
and \U$26494 ( \26871 , \14964 , RIae78788_117);
and \U$26495 ( \26872 , RIae78698_115, \14962 );
nor \U$26496 ( \26873 , \26871 , \26872 );
and \U$26497 ( \26874 , \26873 , \14462 );
not \U$26498 ( \26875 , \26873 );
and \U$26499 ( \26876 , \26875 , \14463 );
nor \U$26500 ( \26877 , \26874 , \26876 );
nor \U$26501 ( \26878 , \26870 , \26877 );
nor \U$26502 ( \26879 , \26869 , \26878 );
and \U$26503 ( \26880 , \9760 , RIae77f18_99);
and \U$26504 ( \26881 , RIae78008_101, \9758 );
nor \U$26505 ( \26882 , \26880 , \26881 );
and \U$26506 ( \26883 , \26882 , \9273 );
not \U$26507 ( \26884 , \26882 );
and \U$26508 ( \26885 , \26884 , \9764 );
nor \U$26509 ( \26886 , \26883 , \26885 );
and \U$26510 ( \26887 , \10548 , RIae781e8_105);
and \U$26511 ( \26888 , RIae785a8_113, \10546 );
nor \U$26512 ( \26889 , \26887 , \26888 );
and \U$26513 ( \26890 , \26889 , \10421 );
not \U$26514 ( \26891 , \26889 );
and \U$26515 ( \26892 , \26891 , \10118 );
nor \U$26516 ( \26893 , \26890 , \26892 );
xor \U$26517 ( \26894 , \26886 , \26893 );
and \U$26518 ( \26895 , \8966 , RIae782d8_107);
and \U$26519 ( \26896 , RIae780f8_103, \8964 );
nor \U$26520 ( \26897 , \26895 , \26896 );
and \U$26521 ( \26898 , \26897 , \8799 );
not \U$26522 ( \26899 , \26897 );
and \U$26523 ( \26900 , \26899 , \8789 );
nor \U$26524 ( \26901 , \26898 , \26900 );
and \U$26525 ( \26902 , \26894 , \26901 );
and \U$26526 ( \26903 , \26886 , \26893 );
nor \U$26527 ( \26904 , \26902 , \26903 );
xor \U$26528 ( \26905 , \26879 , \26904 );
and \U$26529 ( \26906 , \11470 , RIae783c8_109);
and \U$26530 ( \26907 , RIae78530_112, \11468 );
nor \U$26531 ( \26908 , \26906 , \26907 );
and \U$26532 ( \26909 , \26908 , \11474 );
not \U$26533 ( \26910 , \26908 );
and \U$26534 ( \26911 , \26910 , \10936 );
nor \U$26535 ( \26912 , \26909 , \26911 );
not \U$26536 ( \26913 , \26912 );
and \U$26537 ( \26914 , \12180 , RIae77c48_93);
and \U$26538 ( \26915 , RIae77b58_91, \12178 );
nor \U$26539 ( \26916 , \26914 , \26915 );
and \U$26540 ( \26917 , \26916 , \11827 );
not \U$26541 ( \26918 , \26916 );
and \U$26542 ( \26919 , \26918 , \12184 );
nor \U$26543 ( \26920 , \26917 , \26919 );
not \U$26544 ( \26921 , \26920 );
and \U$26545 ( \26922 , \26913 , \26921 );
and \U$26546 ( \26923 , \26920 , \26912 );
and \U$26547 ( \26924 , \13059 , RIae77d38_95);
and \U$26548 ( \26925 , RIae77e28_97, \13057 );
nor \U$26549 ( \26926 , \26924 , \26925 );
and \U$26550 ( \26927 , \26926 , \12718 );
not \U$26551 ( \26928 , \26926 );
and \U$26552 ( \26929 , \26928 , \13063 );
nor \U$26553 ( \26930 , \26927 , \26929 );
nor \U$26554 ( \26931 , \26923 , \26930 );
nor \U$26555 ( \26932 , \26922 , \26931 );
and \U$26556 ( \26933 , \26905 , \26932 );
and \U$26557 ( \26934 , \26879 , \26904 );
nor \U$26558 ( \26935 , \26933 , \26934 );
and \U$26559 ( \26936 , \5399 , RIae77a68_89);
and \U$26560 ( \26937 , RIae77978_87, \5397 );
nor \U$26561 ( \26938 , \26936 , \26937 );
and \U$26562 ( \26939 , \26938 , \5403 );
not \U$26563 ( \26940 , \26938 );
and \U$26564 ( \26941 , \26940 , \5016 );
nor \U$26565 ( \26942 , \26939 , \26941 );
not \U$26566 ( \26943 , \26942 );
and \U$26567 ( \26944 , \5896 , RIae77798_83);
and \U$26568 ( \26945 , RIae77888_85, \5894 );
nor \U$26569 ( \26946 , \26944 , \26945 );
and \U$26570 ( \26947 , \26946 , \5589 );
not \U$26571 ( \26948 , \26946 );
and \U$26572 ( \26949 , \26948 , \5590 );
nor \U$26573 ( \26950 , \26947 , \26949 );
not \U$26574 ( \26951 , \26950 );
and \U$26575 ( \26952 , \26943 , \26951 );
and \U$26576 ( \26953 , \26950 , \26942 );
and \U$26577 ( \26954 , \6172 , RIae76f28_65);
and \U$26578 ( \26955 , RIae76e38_63, \6170 );
nor \U$26579 ( \26956 , \26954 , \26955 );
and \U$26580 ( \26957 , \26956 , \6175 );
not \U$26581 ( \26958 , \26956 );
and \U$26582 ( \26959 , \26958 , \6176 );
nor \U$26583 ( \26960 , \26957 , \26959 );
nor \U$26584 ( \26961 , \26953 , \26960 );
nor \U$26585 ( \26962 , \26952 , \26961 );
and \U$26586 ( \26963 , \4247 , RIae775b8_79);
and \U$26587 ( \26964 , RIae774c8_77, \4245 );
nor \U$26588 ( \26965 , \26963 , \26964 );
and \U$26589 ( \26966 , \26965 , \4251 );
not \U$26590 ( \26967 , \26965 );
and \U$26591 ( \26968 , \26967 , \3989 );
nor \U$26592 ( \26969 , \26966 , \26968 );
not \U$26593 ( \26970 , \26969 );
and \U$26594 ( \26971 , \4688 , RIae77720_82);
and \U$26595 ( \26972 , RIae773d8_75, \4686 );
nor \U$26596 ( \26973 , \26971 , \26972 );
and \U$26597 ( \26974 , \26973 , \4481 );
not \U$26598 ( \26975 , \26973 );
and \U$26599 ( \26976 , \26975 , \4482 );
nor \U$26600 ( \26977 , \26974 , \26976 );
nand \U$26601 ( \26978 , \26970 , \26977 );
or \U$26602 ( \26979 , \26962 , \26978 );
not \U$26603 ( \26980 , \26978 );
not \U$26604 ( \26981 , \26962 );
or \U$26605 ( \26982 , \26980 , \26981 );
and \U$26606 ( \26983 , \8371 , RIae771f8_71);
and \U$26607 ( \26984 , RIae772e8_73, \8369 );
nor \U$26608 ( \26985 , \26983 , \26984 );
and \U$26609 ( \26986 , \26985 , \8020 );
not \U$26610 ( \26987 , \26985 );
and \U$26611 ( \26988 , \26987 , \8019 );
nor \U$26612 ( \26989 , \26986 , \26988 );
and \U$26613 ( \26990 , \6941 , RIae76d48_61);
and \U$26614 ( \26991 , RIae76c58_59, \6939 );
nor \U$26615 ( \26992 , \26990 , \26991 );
and \U$26616 ( \26993 , \26992 , \6314 );
not \U$26617 ( \26994 , \26992 );
and \U$26618 ( \26995 , \26994 , \6945 );
nor \U$26619 ( \26996 , \26993 , \26995 );
xor \U$26620 ( \26997 , \26989 , \26996 );
and \U$26621 ( \26998 , \7633 , RIae77180_70);
and \U$26622 ( \26999 , RIae77018_67, \7631 );
nor \U$26623 ( \27000 , \26998 , \26999 );
and \U$26624 ( \27001 , \27000 , \7206 );
not \U$26625 ( \27002 , \27000 );
and \U$26626 ( \27003 , \27002 , \7205 );
nor \U$26627 ( \27004 , \27001 , \27003 );
and \U$26628 ( \27005 , \26997 , \27004 );
and \U$26629 ( \27006 , \26989 , \26996 );
or \U$26630 ( \27007 , \27005 , \27006 );
nand \U$26631 ( \27008 , \26982 , \27007 );
nand \U$26632 ( \27009 , \26979 , \27008 );
xor \U$26633 ( \27010 , \26935 , \27009 );
nand \U$26634 ( \27011 , RIae775b8_79, \3728 );
and \U$26635 ( \27012 , \27011 , \3422 );
not \U$26636 ( \27013 , \27011 );
and \U$26637 ( \27014 , \27013 , \3732 );
nor \U$26638 ( \27015 , \27012 , \27014 );
xor \U$26639 ( \27016 , \26568 , \26575 );
xor \U$26640 ( \27017 , \27016 , \26583 );
xor \U$26641 ( \27018 , \27015 , \27017 );
xor \U$26642 ( \27019 , \26621 , \26628 );
xor \U$26643 ( \27020 , \27019 , \26636 );
and \U$26644 ( \27021 , \27018 , \27020 );
and \U$26645 ( \27022 , \27015 , \27017 );
nor \U$26646 ( \27023 , \27021 , \27022 );
and \U$26647 ( \27024 , \27010 , \27023 );
and \U$26648 ( \27025 , \26935 , \27009 );
nor \U$26649 ( \27026 , \27024 , \27025 );
nor \U$26650 ( \27027 , \26852 , \27026 );
nor \U$26651 ( \27028 , \26849 , \27027 );
nor \U$26652 ( \27029 , \26813 , \27028 );
nor \U$26653 ( \27030 , \26812 , \27029 );
and \U$26654 ( \27031 , \26794 , \27030 );
and \U$26655 ( \27032 , \26791 , \26793 );
or \U$26656 ( \27033 , \27031 , \27032 );
not \U$26657 ( \27034 , \27033 );
and \U$26658 ( \27035 , \26781 , \27034 );
and \U$26659 ( \27036 , \26780 , \27033 );
nor \U$26660 ( \27037 , \27035 , \27036 );
xor \U$26661 ( \27038 , \26791 , \26793 );
xor \U$26662 ( \27039 , \27038 , \27030 );
not \U$26663 ( \27040 , \27039 );
xor \U$26664 ( \27041 , \26551 , \26759 );
xor \U$26665 ( \27042 , \27041 , \26764 );
nand \U$26666 ( \27043 , \27040 , \27042 );
or \U$26667 ( \27044 , \27037 , \27043 );
xnor \U$26668 ( \27045 , \27043 , \27037 );
not \U$26669 ( \27046 , \27007 );
not \U$26670 ( \27047 , \26962 );
or \U$26671 ( \27048 , \27046 , \27047 );
or \U$26672 ( \27049 , \26962 , \27007 );
nand \U$26673 ( \27050 , \27048 , \27049 );
not \U$26674 ( \27051 , \27050 );
not \U$26675 ( \27052 , \26978 );
and \U$26676 ( \27053 , \27051 , \27052 );
and \U$26677 ( \27054 , \27050 , \26978 );
nor \U$26678 ( \27055 , \27053 , \27054 );
xor \U$26679 ( \27056 , \26879 , \26904 );
xor \U$26680 ( \27057 , \27056 , \26932 );
xor \U$26681 ( \27058 , \27055 , \27057 );
xor \U$26682 ( \27059 , \27015 , \27017 );
xor \U$26683 ( \27060 , \27059 , \27020 );
and \U$26684 ( \27061 , \27058 , \27060 );
and \U$26685 ( \27062 , \27055 , \27057 );
nor \U$26686 ( \27063 , \27061 , \27062 );
and \U$26687 ( \27064 , \6172 , RIae77888_85);
and \U$26688 ( \27065 , RIae76f28_65, \6170 );
nor \U$26689 ( \27066 , \27064 , \27065 );
and \U$26690 ( \27067 , \27066 , \6176 );
not \U$26691 ( \27068 , \27066 );
and \U$26692 ( \27069 , \27068 , \6175 );
nor \U$26693 ( \27070 , \27067 , \27069 );
and \U$26694 ( \27071 , \5896 , RIae77978_87);
and \U$26695 ( \27072 , RIae77798_83, \5894 );
nor \U$26696 ( \27073 , \27071 , \27072 );
and \U$26697 ( \27074 , \27073 , \5590 );
not \U$26698 ( \27075 , \27073 );
and \U$26699 ( \27076 , \27075 , \5589 );
nor \U$26700 ( \27077 , \27074 , \27076 );
xor \U$26701 ( \27078 , \27070 , \27077 );
and \U$26702 ( \27079 , \6941 , RIae76e38_63);
and \U$26703 ( \27080 , RIae76d48_61, \6939 );
nor \U$26704 ( \27081 , \27079 , \27080 );
and \U$26705 ( \27082 , \27081 , \6314 );
not \U$26706 ( \27083 , \27081 );
and \U$26707 ( \27084 , \27083 , \6945 );
nor \U$26708 ( \27085 , \27082 , \27084 );
and \U$26709 ( \27086 , \27078 , \27085 );
and \U$26710 ( \27087 , \27070 , \27077 );
or \U$26711 ( \27088 , \27086 , \27087 );
and \U$26712 ( \27089 , \4688 , RIae774c8_77);
and \U$26713 ( \27090 , RIae77720_82, \4686 );
nor \U$26714 ( \27091 , \27089 , \27090 );
and \U$26715 ( \27092 , \27091 , \4481 );
not \U$26716 ( \27093 , \27091 );
and \U$26717 ( \27094 , \27093 , \4482 );
nor \U$26718 ( \27095 , \27092 , \27094 );
nand \U$26719 ( \27096 , RIae775b8_79, \4245 );
and \U$26720 ( \27097 , \27096 , \3989 );
not \U$26721 ( \27098 , \27096 );
and \U$26722 ( \27099 , \27098 , \4251 );
nor \U$26723 ( \27100 , \27097 , \27099 );
xor \U$26724 ( \27101 , \27095 , \27100 );
and \U$26725 ( \27102 , \5399 , RIae773d8_75);
and \U$26726 ( \27103 , RIae77a68_89, \5397 );
nor \U$26727 ( \27104 , \27102 , \27103 );
and \U$26728 ( \27105 , \27104 , \5016 );
not \U$26729 ( \27106 , \27104 );
and \U$26730 ( \27107 , \27106 , \5403 );
nor \U$26731 ( \27108 , \27105 , \27107 );
and \U$26732 ( \27109 , \27101 , \27108 );
and \U$26733 ( \27110 , \27095 , \27100 );
or \U$26734 ( \27111 , \27109 , \27110 );
xor \U$26735 ( \27112 , \27088 , \27111 );
and \U$26736 ( \27113 , \8371 , RIae77018_67);
and \U$26737 ( \27114 , RIae771f8_71, \8369 );
nor \U$26738 ( \27115 , \27113 , \27114 );
and \U$26739 ( \27116 , \27115 , \8020 );
not \U$26740 ( \27117 , \27115 );
and \U$26741 ( \27118 , \27117 , \8019 );
nor \U$26742 ( \27119 , \27116 , \27118 );
and \U$26743 ( \27120 , \7633 , RIae76c58_59);
and \U$26744 ( \27121 , RIae77180_70, \7631 );
nor \U$26745 ( \27122 , \27120 , \27121 );
and \U$26746 ( \27123 , \27122 , \7206 );
not \U$26747 ( \27124 , \27122 );
and \U$26748 ( \27125 , \27124 , \7205 );
nor \U$26749 ( \27126 , \27123 , \27125 );
xor \U$26750 ( \27127 , \27119 , \27126 );
and \U$26751 ( \27128 , \8966 , RIae772e8_73);
and \U$26752 ( \27129 , RIae782d8_107, \8964 );
nor \U$26753 ( \27130 , \27128 , \27129 );
and \U$26754 ( \27131 , \27130 , \8799 );
not \U$26755 ( \27132 , \27130 );
and \U$26756 ( \27133 , \27132 , \8789 );
nor \U$26757 ( \27134 , \27131 , \27133 );
and \U$26758 ( \27135 , \27127 , \27134 );
and \U$26759 ( \27136 , \27119 , \27126 );
or \U$26760 ( \27137 , \27135 , \27136 );
and \U$26761 ( \27138 , \27112 , \27137 );
and \U$26762 ( \27139 , \27088 , \27111 );
or \U$26763 ( \27140 , \27138 , \27139 );
and \U$26764 ( \27141 , \9760 , RIae780f8_103);
and \U$26765 ( \27142 , RIae77f18_99, \9758 );
nor \U$26766 ( \27143 , \27141 , \27142 );
and \U$26767 ( \27144 , \27143 , \9273 );
not \U$26768 ( \27145 , \27143 );
and \U$26769 ( \27146 , \27145 , \9272 );
nor \U$26770 ( \27147 , \27144 , \27146 );
and \U$26771 ( \27148 , \10548 , RIae78008_101);
and \U$26772 ( \27149 , RIae781e8_105, \10546 );
nor \U$26773 ( \27150 , \27148 , \27149 );
and \U$26774 ( \27151 , \27150 , \10421 );
not \U$26775 ( \27152 , \27150 );
and \U$26776 ( \27153 , \27152 , \10118 );
nor \U$26777 ( \27154 , \27151 , \27153 );
xor \U$26778 ( \27155 , \27147 , \27154 );
and \U$26779 ( \27156 , \11470 , RIae785a8_113);
and \U$26780 ( \27157 , RIae783c8_109, \11468 );
nor \U$26781 ( \27158 , \27156 , \27157 );
and \U$26782 ( \27159 , \27158 , \10936 );
not \U$26783 ( \27160 , \27158 );
and \U$26784 ( \27161 , \27160 , \11474 );
nor \U$26785 ( \27162 , \27159 , \27161 );
and \U$26786 ( \27163 , \27155 , \27162 );
and \U$26787 ( \27164 , \27147 , \27154 );
or \U$26788 ( \27165 , \27163 , \27164 );
and \U$26789 ( \27166 , \15726 , RIae78698_115);
and \U$26790 ( \27167 , RIae7aab0_192, RIae75b78_23);
nor \U$26791 ( \27168 , \27166 , \27167 );
and \U$26792 ( \27169 , \27168 , \14959 );
not \U$26793 ( \27170 , \27168 );
and \U$26794 ( \27171 , \27170 , RIae7aa38_191);
nor \U$26795 ( \27172 , \27169 , \27171 );
xor \U$26796 ( \27173 , \27172 , \4251 );
and \U$26797 ( \27174 , \14964 , RIae78878_119);
and \U$26798 ( \27175 , RIae78788_117, \14962 );
nor \U$26799 ( \27176 , \27174 , \27175 );
and \U$26800 ( \27177 , \27176 , \14463 );
not \U$26801 ( \27178 , \27176 );
and \U$26802 ( \27179 , \27178 , \14462 );
nor \U$26803 ( \27180 , \27177 , \27179 );
and \U$26804 ( \27181 , \27173 , \27180 );
and \U$26805 ( \27182 , \27172 , \4251 );
or \U$26806 ( \27183 , \27181 , \27182 );
xor \U$26807 ( \27184 , \27165 , \27183 );
and \U$26808 ( \27185 , \12180 , RIae78530_112);
and \U$26809 ( \27186 , RIae77c48_93, \12178 );
nor \U$26810 ( \27187 , \27185 , \27186 );
and \U$26811 ( \27188 , \27187 , \12184 );
not \U$26812 ( \27189 , \27187 );
and \U$26813 ( \27190 , \27189 , \11827 );
nor \U$26814 ( \27191 , \27188 , \27190 );
and \U$26815 ( \27192 , \13059 , RIae77b58_91);
and \U$26816 ( \27193 , RIae77d38_95, \13057 );
nor \U$26817 ( \27194 , \27192 , \27193 );
and \U$26818 ( \27195 , \27194 , \13063 );
not \U$26819 ( \27196 , \27194 );
and \U$26820 ( \27197 , \27196 , \12718 );
nor \U$26821 ( \27198 , \27195 , \27197 );
xor \U$26822 ( \27199 , \27191 , \27198 );
and \U$26823 ( \27200 , \14059 , RIae77e28_97);
and \U$26824 ( \27201 , RIae78968_121, \14057 );
nor \U$26825 ( \27202 , \27200 , \27201 );
and \U$26826 ( \27203 , \27202 , \13502 );
not \U$26827 ( \27204 , \27202 );
and \U$26828 ( \27205 , \27204 , \14063 );
nor \U$26829 ( \27206 , \27203 , \27205 );
and \U$26830 ( \27207 , \27199 , \27206 );
and \U$26831 ( \27208 , \27191 , \27198 );
or \U$26832 ( \27209 , \27207 , \27208 );
and \U$26833 ( \27210 , \27184 , \27209 );
and \U$26834 ( \27211 , \27165 , \27183 );
or \U$26835 ( \27212 , \27210 , \27211 );
xor \U$26836 ( \27213 , \27140 , \27212 );
not \U$26837 ( \27214 , \26942 );
xor \U$26838 ( \27215 , \26950 , \26960 );
not \U$26839 ( \27216 , \27215 );
or \U$26840 ( \27217 , \27214 , \27216 );
or \U$26841 ( \27218 , \27215 , \26942 );
nand \U$26842 ( \27219 , \27217 , \27218 );
not \U$26843 ( \27220 , \26969 );
not \U$26844 ( \27221 , \26977 );
or \U$26845 ( \27222 , \27220 , \27221 );
or \U$26846 ( \27223 , \26969 , \26977 );
nand \U$26847 ( \27224 , \27222 , \27223 );
xor \U$26848 ( \27225 , \27219 , \27224 );
xor \U$26849 ( \27226 , \26989 , \26996 );
xor \U$26850 ( \27227 , \27226 , \27004 );
and \U$26851 ( \27228 , \27225 , \27227 );
and \U$26852 ( \27229 , \27219 , \27224 );
or \U$26853 ( \27230 , \27228 , \27229 );
and \U$26854 ( \27231 , \27213 , \27230 );
and \U$26855 ( \27232 , \27140 , \27212 );
or \U$26856 ( \27233 , \27231 , \27232 );
xor \U$26857 ( \27234 , \27063 , \27233 );
not \U$26858 ( \27235 , \26859 );
xor \U$26859 ( \27236 , \26867 , \26877 );
not \U$26860 ( \27237 , \27236 );
or \U$26861 ( \27238 , \27235 , \27237 );
or \U$26862 ( \27239 , \27236 , \26859 );
nand \U$26863 ( \27240 , \27238 , \27239 );
xor \U$26864 ( \27241 , \26886 , \26893 );
xor \U$26865 ( \27242 , \27241 , \26901 );
xor \U$26866 ( \27243 , \27240 , \27242 );
not \U$26867 ( \27244 , \26912 );
xor \U$26868 ( \27245 , \26920 , \26930 );
not \U$26869 ( \27246 , \27245 );
or \U$26870 ( \27247 , \27244 , \27246 );
or \U$26871 ( \27248 , \27245 , \26912 );
nand \U$26872 ( \27249 , \27247 , \27248 );
and \U$26873 ( \27250 , \27243 , \27249 );
and \U$26874 ( \27251 , \27240 , \27242 );
or \U$26875 ( \27252 , \27250 , \27251 );
xor \U$26876 ( \27253 , \26674 , \3422 );
xor \U$26877 ( \27254 , \27253 , \26682 );
xor \U$26878 ( \27255 , \27252 , \27254 );
xor \U$26879 ( \27256 , \26649 , \26656 );
xor \U$26880 ( \27257 , \27256 , \26664 );
xor \U$26881 ( \27258 , \26819 , \26824 );
xor \U$26882 ( \27259 , \27257 , \27258 );
and \U$26883 ( \27260 , \27255 , \27259 );
and \U$26884 ( \27261 , \27252 , \27254 );
or \U$26885 ( \27262 , \27260 , \27261 );
and \U$26886 ( \27263 , \27234 , \27262 );
and \U$26887 ( \27264 , \27063 , \27233 );
or \U$26888 ( \27265 , \27263 , \27264 );
xor \U$26889 ( \27266 , \26935 , \27009 );
xor \U$26890 ( \27267 , \27266 , \27023 );
not \U$26891 ( \27268 , \26846 );
not \U$26892 ( \27269 , \26843 );
or \U$26893 ( \27270 , \27268 , \27269 );
or \U$26894 ( \27271 , \26843 , \26846 );
nand \U$26895 ( \27272 , \27270 , \27271 );
xor \U$26896 ( \27273 , \27267 , \27272 );
xor \U$26897 ( \27274 , \26717 , \26719 );
xor \U$26898 ( \27275 , \27274 , \26722 );
xor \U$26899 ( \27276 , \26829 , \26836 );
xor \U$26900 ( \27277 , \27275 , \27276 );
and \U$26901 ( \27278 , \27273 , \27277 );
and \U$26902 ( \27279 , \27267 , \27272 );
or \U$26903 ( \27280 , \27278 , \27279 );
xor \U$26904 ( \27281 , \27265 , \27280 );
xor \U$26905 ( \27282 , \26553 , \26555 );
xor \U$26906 ( \27283 , \27282 , \26558 );
xor \U$26907 ( \27284 , \26796 , \26801 );
xor \U$26908 ( \27285 , \27283 , \27284 );
and \U$26909 ( \27286 , \27281 , \27285 );
and \U$26910 ( \27287 , \27265 , \27280 );
or \U$26911 ( \27288 , \27286 , \27287 );
not \U$26912 ( \27289 , \26810 );
xor \U$26913 ( \27290 , \27028 , \26807 );
not \U$26914 ( \27291 , \27290 );
or \U$26915 ( \27292 , \27289 , \27291 );
or \U$26916 ( \27293 , \27290 , \26810 );
nand \U$26917 ( \27294 , \27292 , \27293 );
xnor \U$26918 ( \27295 , \27288 , \27294 );
not \U$26919 ( \27296 , \27295 );
not \U$26920 ( \27297 , \26790 );
not \U$26921 ( \27298 , \26787 );
or \U$26922 ( \27299 , \27297 , \27298 );
or \U$26923 ( \27300 , \26787 , \26790 );
nand \U$26924 ( \27301 , \27299 , \27300 );
not \U$26925 ( \27302 , \27301 );
and \U$26926 ( \27303 , \27296 , \27302 );
and \U$26927 ( \27304 , \27295 , \27301 );
nor \U$26928 ( \27305 , \27303 , \27304 );
xor \U$26929 ( \27306 , \27265 , \27280 );
xor \U$26930 ( \27307 , \27306 , \27285 );
not \U$26931 ( \27308 , \26847 );
not \U$26932 ( \27309 , \27026 );
not \U$26933 ( \27310 , \26841 );
or \U$26934 ( \27311 , \27309 , \27310 );
or \U$26935 ( \27312 , \26841 , \27026 );
nand \U$26936 ( \27313 , \27311 , \27312 );
not \U$26937 ( \27314 , \27313 );
or \U$26938 ( \27315 , \27308 , \27314 );
or \U$26939 ( \27316 , \27313 , \26847 );
nand \U$26940 ( \27317 , \27315 , \27316 );
xor \U$26941 ( \27318 , \27307 , \27317 );
xor \U$26942 ( \27319 , \27055 , \27057 );
xor \U$26943 ( \27320 , \27319 , \27060 );
xor \U$26944 ( \27321 , \27070 , \27077 );
xor \U$26945 ( \27322 , \27321 , \27085 );
xor \U$26946 ( \27323 , \27119 , \27126 );
xor \U$26947 ( \27324 , \27323 , \27134 );
and \U$26948 ( \27325 , \27322 , \27324 );
xor \U$26949 ( \27326 , \27147 , \27154 );
xor \U$26950 ( \27327 , \27326 , \27162 );
xor \U$26951 ( \27328 , \27119 , \27126 );
xor \U$26952 ( \27329 , \27328 , \27134 );
and \U$26953 ( \27330 , \27327 , \27329 );
and \U$26954 ( \27331 , \27322 , \27327 );
or \U$26955 ( \27332 , \27325 , \27330 , \27331 );
and \U$26956 ( \27333 , \11470 , RIae781e8_105);
and \U$26957 ( \27334 , RIae785a8_113, \11468 );
nor \U$26958 ( \27335 , \27333 , \27334 );
and \U$26959 ( \27336 , \27335 , \10936 );
not \U$26960 ( \27337 , \27335 );
and \U$26961 ( \27338 , \27337 , \11474 );
nor \U$26962 ( \27339 , \27336 , \27338 );
and \U$26963 ( \27340 , \12180 , RIae783c8_109);
and \U$26964 ( \27341 , RIae78530_112, \12178 );
nor \U$26965 ( \27342 , \27340 , \27341 );
and \U$26966 ( \27343 , \27342 , \12184 );
not \U$26967 ( \27344 , \27342 );
and \U$26968 ( \27345 , \27344 , \11827 );
nor \U$26969 ( \27346 , \27343 , \27345 );
xor \U$26970 ( \27347 , \27339 , \27346 );
and \U$26971 ( \27348 , \13059 , RIae77c48_93);
and \U$26972 ( \27349 , RIae77b58_91, \13057 );
nor \U$26973 ( \27350 , \27348 , \27349 );
and \U$26974 ( \27351 , \27350 , \13063 );
not \U$26975 ( \27352 , \27350 );
and \U$26976 ( \27353 , \27352 , \12718 );
nor \U$26977 ( \27354 , \27351 , \27353 );
and \U$26978 ( \27355 , \27347 , \27354 );
and \U$26979 ( \27356 , \27339 , \27346 );
or \U$26980 ( \27357 , \27355 , \27356 );
and \U$26981 ( \27358 , \14059 , RIae77d38_95);
and \U$26982 ( \27359 , RIae77e28_97, \14057 );
nor \U$26983 ( \27360 , \27358 , \27359 );
and \U$26984 ( \27361 , \27360 , \13502 );
not \U$26985 ( \27362 , \27360 );
and \U$26986 ( \27363 , \27362 , \14063 );
nor \U$26987 ( \27364 , \27361 , \27363 );
and \U$26988 ( \27365 , \15726 , RIae78788_117);
and \U$26989 ( \27366 , RIae7aab0_192, RIae78698_115);
nor \U$26990 ( \27367 , \27365 , \27366 );
and \U$26991 ( \27368 , \27367 , \14959 );
not \U$26992 ( \27369 , \27367 );
and \U$26993 ( \27370 , \27369 , RIae7aa38_191);
nor \U$26994 ( \27371 , \27368 , \27370 );
xor \U$26995 ( \27372 , \27364 , \27371 );
and \U$26996 ( \27373 , \14964 , RIae78968_121);
and \U$26997 ( \27374 , RIae78878_119, \14962 );
nor \U$26998 ( \27375 , \27373 , \27374 );
and \U$26999 ( \27376 , \27375 , \14463 );
not \U$27000 ( \27377 , \27375 );
and \U$27001 ( \27378 , \27377 , \14462 );
nor \U$27002 ( \27379 , \27376 , \27378 );
and \U$27003 ( \27380 , \27372 , \27379 );
and \U$27004 ( \27381 , \27364 , \27371 );
or \U$27005 ( \27382 , \27380 , \27381 );
xor \U$27006 ( \27383 , \27357 , \27382 );
and \U$27007 ( \27384 , \10548 , RIae77f18_99);
and \U$27008 ( \27385 , RIae78008_101, \10546 );
nor \U$27009 ( \27386 , \27384 , \27385 );
and \U$27010 ( \27387 , \27386 , \10421 );
not \U$27011 ( \27388 , \27386 );
and \U$27012 ( \27389 , \27388 , \10118 );
nor \U$27013 ( \27390 , \27387 , \27389 );
and \U$27014 ( \27391 , \8966 , RIae771f8_71);
and \U$27015 ( \27392 , RIae772e8_73, \8964 );
nor \U$27016 ( \27393 , \27391 , \27392 );
and \U$27017 ( \27394 , \27393 , \8799 );
not \U$27018 ( \27395 , \27393 );
and \U$27019 ( \27396 , \27395 , \8789 );
nor \U$27020 ( \27397 , \27394 , \27396 );
xor \U$27021 ( \27398 , \27390 , \27397 );
and \U$27022 ( \27399 , \9760 , RIae782d8_107);
and \U$27023 ( \27400 , RIae780f8_103, \9758 );
nor \U$27024 ( \27401 , \27399 , \27400 );
and \U$27025 ( \27402 , \27401 , \9273 );
not \U$27026 ( \27403 , \27401 );
and \U$27027 ( \27404 , \27403 , \9764 );
nor \U$27028 ( \27405 , \27402 , \27404 );
and \U$27029 ( \27406 , \27398 , \27405 );
and \U$27030 ( \27407 , \27390 , \27397 );
or \U$27031 ( \27408 , \27406 , \27407 );
and \U$27032 ( \27409 , \27383 , \27408 );
and \U$27033 ( \27410 , \27357 , \27382 );
or \U$27034 ( \27411 , \27409 , \27410 );
xor \U$27035 ( \27412 , \27332 , \27411 );
and \U$27036 ( \27413 , \6941 , RIae76f28_65);
and \U$27037 ( \27414 , RIae76e38_63, \6939 );
nor \U$27038 ( \27415 , \27413 , \27414 );
and \U$27039 ( \27416 , \27415 , \6314 );
not \U$27040 ( \27417 , \27415 );
and \U$27041 ( \27418 , \27417 , \6945 );
nor \U$27042 ( \27419 , \27416 , \27418 );
and \U$27043 ( \27420 , \7633 , RIae76d48_61);
and \U$27044 ( \27421 , RIae76c58_59, \7631 );
nor \U$27045 ( \27422 , \27420 , \27421 );
and \U$27046 ( \27423 , \27422 , \7206 );
not \U$27047 ( \27424 , \27422 );
and \U$27048 ( \27425 , \27424 , \7205 );
nor \U$27049 ( \27426 , \27423 , \27425 );
xor \U$27050 ( \27427 , \27419 , \27426 );
and \U$27051 ( \27428 , \8371 , RIae77180_70);
and \U$27052 ( \27429 , RIae77018_67, \8369 );
nor \U$27053 ( \27430 , \27428 , \27429 );
and \U$27054 ( \27431 , \27430 , \8020 );
not \U$27055 ( \27432 , \27430 );
and \U$27056 ( \27433 , \27432 , \8019 );
nor \U$27057 ( \27434 , \27431 , \27433 );
and \U$27058 ( \27435 , \27427 , \27434 );
and \U$27059 ( \27436 , \27419 , \27426 );
or \U$27060 ( \27437 , \27435 , \27436 );
and \U$27061 ( \27438 , \5399 , RIae77720_82);
and \U$27062 ( \27439 , RIae773d8_75, \5397 );
nor \U$27063 ( \27440 , \27438 , \27439 );
and \U$27064 ( \27441 , \27440 , \5016 );
not \U$27065 ( \27442 , \27440 );
and \U$27066 ( \27443 , \27442 , \5403 );
nor \U$27067 ( \27444 , \27441 , \27443 );
and \U$27068 ( \27445 , \5896 , RIae77a68_89);
and \U$27069 ( \27446 , RIae77978_87, \5894 );
nor \U$27070 ( \27447 , \27445 , \27446 );
and \U$27071 ( \27448 , \27447 , \5590 );
not \U$27072 ( \27449 , \27447 );
and \U$27073 ( \27450 , \27449 , \5589 );
nor \U$27074 ( \27451 , \27448 , \27450 );
xor \U$27075 ( \27452 , \27444 , \27451 );
and \U$27076 ( \27453 , \6172 , RIae77798_83);
and \U$27077 ( \27454 , RIae77888_85, \6170 );
nor \U$27078 ( \27455 , \27453 , \27454 );
and \U$27079 ( \27456 , \27455 , \6176 );
not \U$27080 ( \27457 , \27455 );
and \U$27081 ( \27458 , \27457 , \6175 );
nor \U$27082 ( \27459 , \27456 , \27458 );
and \U$27083 ( \27460 , \27452 , \27459 );
and \U$27084 ( \27461 , \27444 , \27451 );
or \U$27085 ( \27462 , \27460 , \27461 );
xor \U$27086 ( \27463 , \27437 , \27462 );
xor \U$27087 ( \27464 , \27095 , \27100 );
xor \U$27088 ( \27465 , \27464 , \27108 );
and \U$27089 ( \27466 , \27463 , \27465 );
and \U$27090 ( \27467 , \27437 , \27462 );
or \U$27091 ( \27468 , \27466 , \27467 );
and \U$27092 ( \27469 , \27412 , \27468 );
and \U$27093 ( \27470 , \27332 , \27411 );
nor \U$27094 ( \27471 , \27469 , \27470 );
or \U$27095 ( \27472 , \27320 , \27471 );
not \U$27096 ( \27473 , \27471 );
not \U$27097 ( \27474 , \27320 );
or \U$27098 ( \27475 , \27473 , \27474 );
xor \U$27099 ( \27476 , \27088 , \27111 );
xor \U$27100 ( \27477 , \27476 , \27137 );
xor \U$27101 ( \27478 , \27219 , \27224 );
xor \U$27102 ( \27479 , \27478 , \27227 );
and \U$27103 ( \27480 , \27477 , \27479 );
xor \U$27104 ( \27481 , \27240 , \27242 );
xor \U$27105 ( \27482 , \27481 , \27249 );
xor \U$27106 ( \27483 , \27219 , \27224 );
xor \U$27107 ( \27484 , \27483 , \27227 );
and \U$27108 ( \27485 , \27482 , \27484 );
and \U$27109 ( \27486 , \27477 , \27482 );
or \U$27110 ( \27487 , \27480 , \27485 , \27486 );
nand \U$27111 ( \27488 , \27475 , \27487 );
nand \U$27112 ( \27489 , \27472 , \27488 );
xor \U$27113 ( \27490 , \27063 , \27233 );
xor \U$27114 ( \27491 , \27490 , \27262 );
and \U$27115 ( \27492 , \27489 , \27491 );
xor \U$27116 ( \27493 , \27267 , \27272 );
xor \U$27117 ( \27494 , \27493 , \27277 );
xor \U$27118 ( \27495 , \27063 , \27233 );
xor \U$27119 ( \27496 , \27495 , \27262 );
and \U$27120 ( \27497 , \27494 , \27496 );
and \U$27121 ( \27498 , \27489 , \27494 );
or \U$27122 ( \27499 , \27492 , \27497 , \27498 );
and \U$27123 ( \27500 , \27318 , \27499 );
and \U$27124 ( \27501 , \27307 , \27317 );
nor \U$27125 ( \27502 , \27500 , \27501 );
or \U$27126 ( \27503 , \27305 , \27502 );
xnor \U$27127 ( \27504 , \27502 , \27305 );
xor \U$27128 ( \27505 , \27140 , \27212 );
xor \U$27129 ( \27506 , \27505 , \27230 );
not \U$27130 ( \27507 , \27506 );
not \U$27131 ( \27508 , \27471 );
not \U$27132 ( \27509 , \27487 );
or \U$27133 ( \27510 , \27508 , \27509 );
or \U$27134 ( \27511 , \27487 , \27471 );
nand \U$27135 ( \27512 , \27510 , \27511 );
not \U$27136 ( \27513 , \27512 );
not \U$27137 ( \27514 , \27320 );
and \U$27138 ( \27515 , \27513 , \27514 );
and \U$27139 ( \27516 , \27512 , \27320 );
nor \U$27140 ( \27517 , \27515 , \27516 );
not \U$27141 ( \27518 , \27517 );
or \U$27142 ( \27519 , \27507 , \27518 );
or \U$27143 ( \27520 , \27517 , \27506 );
nand \U$27144 ( \27521 , \27519 , \27520 );
and \U$27145 ( \27522 , \8966 , RIae77180_70);
and \U$27146 ( \27523 , RIae77018_67, \8964 );
nor \U$27147 ( \27524 , \27522 , \27523 );
and \U$27148 ( \27525 , \27524 , \8789 );
not \U$27149 ( \27526 , \27524 );
and \U$27150 ( \27527 , \27526 , \8799 );
nor \U$27151 ( \27528 , \27525 , \27527 );
not \U$27152 ( \27529 , \27528 );
and \U$27153 ( \27530 , \9760 , RIae771f8_71);
and \U$27154 ( \27531 , RIae772e8_73, \9758 );
nor \U$27155 ( \27532 , \27530 , \27531 );
and \U$27156 ( \27533 , \27532 , \9272 );
not \U$27157 ( \27534 , \27532 );
and \U$27158 ( \27535 , \27534 , \9273 );
nor \U$27159 ( \27536 , \27533 , \27535 );
not \U$27160 ( \27537 , \27536 );
and \U$27161 ( \27538 , \27529 , \27537 );
and \U$27162 ( \27539 , \27536 , \27528 );
and \U$27163 ( \27540 , \10548 , RIae782d8_107);
and \U$27164 ( \27541 , RIae780f8_103, \10546 );
nor \U$27165 ( \27542 , \27540 , \27541 );
and \U$27166 ( \27543 , \27542 , \10118 );
not \U$27167 ( \27544 , \27542 );
and \U$27168 ( \27545 , \27544 , \10421 );
nor \U$27169 ( \27546 , \27543 , \27545 );
nor \U$27170 ( \27547 , \27539 , \27546 );
nor \U$27171 ( \27548 , \27538 , \27547 );
and \U$27172 ( \27549 , \11470 , RIae77f18_99);
and \U$27173 ( \27550 , RIae78008_101, \11468 );
nor \U$27174 ( \27551 , \27549 , \27550 );
and \U$27175 ( \27552 , \27551 , \11474 );
not \U$27176 ( \27553 , \27551 );
and \U$27177 ( \27554 , \27553 , \10936 );
nor \U$27178 ( \27555 , \27552 , \27554 );
not \U$27179 ( \27556 , \27555 );
and \U$27180 ( \27557 , \13059 , RIae783c8_109);
and \U$27181 ( \27558 , RIae78530_112, \13057 );
nor \U$27182 ( \27559 , \27557 , \27558 );
and \U$27183 ( \27560 , \27559 , \12718 );
not \U$27184 ( \27561 , \27559 );
and \U$27185 ( \27562 , \27561 , \13063 );
nor \U$27186 ( \27563 , \27560 , \27562 );
not \U$27187 ( \27564 , \27563 );
and \U$27188 ( \27565 , \27556 , \27564 );
and \U$27189 ( \27566 , \27563 , \27555 );
and \U$27190 ( \27567 , \12180 , RIae781e8_105);
and \U$27191 ( \27568 , RIae785a8_113, \12178 );
nor \U$27192 ( \27569 , \27567 , \27568 );
and \U$27193 ( \27570 , \27569 , \11827 );
not \U$27194 ( \27571 , \27569 );
and \U$27195 ( \27572 , \27571 , \12184 );
nor \U$27196 ( \27573 , \27570 , \27572 );
nor \U$27197 ( \27574 , \27566 , \27573 );
nor \U$27198 ( \27575 , \27565 , \27574 );
xor \U$27199 ( \27576 , \27548 , \27575 );
and \U$27200 ( \27577 , \14964 , RIae77d38_95);
and \U$27201 ( \27578 , RIae77e28_97, \14962 );
nor \U$27202 ( \27579 , \27577 , \27578 );
and \U$27203 ( \27580 , \27579 , \14463 );
not \U$27204 ( \27581 , \27579 );
and \U$27205 ( \27582 , \27581 , \14462 );
nor \U$27206 ( \27583 , \27580 , \27582 );
and \U$27207 ( \27584 , \15726 , RIae78968_121);
and \U$27208 ( \27585 , RIae7aab0_192, RIae78878_119);
nor \U$27209 ( \27586 , \27584 , \27585 );
and \U$27210 ( \27587 , \27586 , \14959 );
not \U$27211 ( \27588 , \27586 );
and \U$27212 ( \27589 , \27588 , RIae7aa38_191);
nor \U$27213 ( \27590 , \27587 , \27589 );
xor \U$27214 ( \27591 , \27583 , \27590 );
and \U$27215 ( \27592 , \14059 , RIae77c48_93);
and \U$27216 ( \27593 , RIae77b58_91, \14057 );
nor \U$27217 ( \27594 , \27592 , \27593 );
and \U$27218 ( \27595 , \27594 , \13502 );
not \U$27219 ( \27596 , \27594 );
and \U$27220 ( \27597 , \27596 , \14063 );
nor \U$27221 ( \27598 , \27595 , \27597 );
and \U$27222 ( \27599 , \27591 , \27598 );
and \U$27223 ( \27600 , \27583 , \27590 );
nor \U$27224 ( \27601 , \27599 , \27600 );
and \U$27225 ( \27602 , \27576 , \27601 );
and \U$27226 ( \27603 , \27548 , \27575 );
nor \U$27227 ( \27604 , \27602 , \27603 );
and \U$27228 ( \27605 , \6941 , RIae77798_83);
and \U$27229 ( \27606 , RIae77888_85, \6939 );
nor \U$27230 ( \27607 , \27605 , \27606 );
and \U$27231 ( \27608 , \27607 , \6314 );
not \U$27232 ( \27609 , \27607 );
and \U$27233 ( \27610 , \27609 , \6945 );
nor \U$27234 ( \27611 , \27608 , \27610 );
and \U$27235 ( \27612 , \7633 , RIae76f28_65);
and \U$27236 ( \27613 , RIae76e38_63, \7631 );
nor \U$27237 ( \27614 , \27612 , \27613 );
and \U$27238 ( \27615 , \27614 , \7206 );
not \U$27239 ( \27616 , \27614 );
and \U$27240 ( \27617 , \27616 , \7205 );
nor \U$27241 ( \27618 , \27615 , \27617 );
xor \U$27242 ( \27619 , \27611 , \27618 );
and \U$27243 ( \27620 , \8371 , RIae76d48_61);
and \U$27244 ( \27621 , RIae76c58_59, \8369 );
nor \U$27245 ( \27622 , \27620 , \27621 );
and \U$27246 ( \27623 , \27622 , \8020 );
not \U$27247 ( \27624 , \27622 );
and \U$27248 ( \27625 , \27624 , \8019 );
nor \U$27249 ( \27626 , \27623 , \27625 );
and \U$27250 ( \27627 , \27619 , \27626 );
and \U$27251 ( \27628 , \27611 , \27618 );
or \U$27252 ( \27629 , \27627 , \27628 );
and \U$27253 ( \27630 , \5399 , RIae774c8_77);
and \U$27254 ( \27631 , RIae77720_82, \5397 );
nor \U$27255 ( \27632 , \27630 , \27631 );
and \U$27256 ( \27633 , \27632 , \5016 );
not \U$27257 ( \27634 , \27632 );
and \U$27258 ( \27635 , \27634 , \5403 );
nor \U$27259 ( \27636 , \27633 , \27635 );
xor \U$27260 ( \27637 , \27629 , \27636 );
and \U$27261 ( \27638 , \6172 , RIae77a68_89);
and \U$27262 ( \27639 , RIae77978_87, \6170 );
nor \U$27263 ( \27640 , \27638 , \27639 );
and \U$27264 ( \27641 , \27640 , \6176 );
not \U$27265 ( \27642 , \27640 );
and \U$27266 ( \27643 , \27642 , \6175 );
nor \U$27267 ( \27644 , \27641 , \27643 );
and \U$27268 ( \27645 , \5399 , RIae775b8_79);
and \U$27269 ( \27646 , RIae774c8_77, \5397 );
nor \U$27270 ( \27647 , \27645 , \27646 );
and \U$27271 ( \27648 , \27647 , \5016 );
not \U$27272 ( \27649 , \27647 );
and \U$27273 ( \27650 , \27649 , \5403 );
nor \U$27274 ( \27651 , \27648 , \27650 );
xor \U$27275 ( \27652 , \27644 , \27651 );
and \U$27276 ( \27653 , \5896 , RIae77720_82);
and \U$27277 ( \27654 , RIae773d8_75, \5894 );
nor \U$27278 ( \27655 , \27653 , \27654 );
and \U$27279 ( \27656 , \27655 , \5590 );
not \U$27280 ( \27657 , \27655 );
and \U$27281 ( \27658 , \27657 , \5589 );
nor \U$27282 ( \27659 , \27656 , \27658 );
and \U$27283 ( \27660 , \27652 , \27659 );
and \U$27284 ( \27661 , \27644 , \27651 );
or \U$27285 ( \27662 , \27660 , \27661 );
and \U$27286 ( \27663 , \27637 , \27662 );
and \U$27287 ( \27664 , \27629 , \27636 );
or \U$27288 ( \27665 , \27663 , \27664 );
xor \U$27289 ( \27666 , \27604 , \27665 );
and \U$27290 ( \27667 , \5896 , RIae773d8_75);
and \U$27291 ( \27668 , RIae77a68_89, \5894 );
nor \U$27292 ( \27669 , \27667 , \27668 );
and \U$27293 ( \27670 , \27669 , \5590 );
not \U$27294 ( \27671 , \27669 );
and \U$27295 ( \27672 , \27671 , \5589 );
nor \U$27296 ( \27673 , \27670 , \27672 );
and \U$27297 ( \27674 , \6172 , RIae77978_87);
and \U$27298 ( \27675 , RIae77798_83, \6170 );
nor \U$27299 ( \27676 , \27674 , \27675 );
and \U$27300 ( \27677 , \27676 , \6176 );
not \U$27301 ( \27678 , \27676 );
and \U$27302 ( \27679 , \27678 , \6175 );
nor \U$27303 ( \27680 , \27677 , \27679 );
xor \U$27304 ( \27681 , \27673 , \27680 );
and \U$27305 ( \27682 , \6941 , RIae77888_85);
and \U$27306 ( \27683 , RIae76f28_65, \6939 );
nor \U$27307 ( \27684 , \27682 , \27683 );
and \U$27308 ( \27685 , \27684 , \6314 );
not \U$27309 ( \27686 , \27684 );
and \U$27310 ( \27687 , \27686 , \6945 );
nor \U$27311 ( \27688 , \27685 , \27687 );
xor \U$27312 ( \27689 , \27681 , \27688 );
nand \U$27313 ( \27690 , RIae775b8_79, \4686 );
and \U$27314 ( \27691 , \27690 , \4481 );
not \U$27315 ( \27692 , \27690 );
and \U$27316 ( \27693 , \27692 , \4482 );
nor \U$27317 ( \27694 , \27691 , \27693 );
xor \U$27318 ( \27695 , \27689 , \27694 );
and \U$27319 ( \27696 , \8966 , RIae77018_67);
and \U$27320 ( \27697 , RIae771f8_71, \8964 );
nor \U$27321 ( \27698 , \27696 , \27697 );
and \U$27322 ( \27699 , \27698 , \8799 );
not \U$27323 ( \27700 , \27698 );
and \U$27324 ( \27701 , \27700 , \8789 );
nor \U$27325 ( \27702 , \27699 , \27701 );
and \U$27326 ( \27703 , \7633 , RIae76e38_63);
and \U$27327 ( \27704 , RIae76d48_61, \7631 );
nor \U$27328 ( \27705 , \27703 , \27704 );
and \U$27329 ( \27706 , \27705 , \7206 );
not \U$27330 ( \27707 , \27705 );
and \U$27331 ( \27708 , \27707 , \7205 );
nor \U$27332 ( \27709 , \27706 , \27708 );
xor \U$27333 ( \27710 , \27702 , \27709 );
and \U$27334 ( \27711 , \8371 , RIae76c58_59);
and \U$27335 ( \27712 , RIae77180_70, \8369 );
nor \U$27336 ( \27713 , \27711 , \27712 );
and \U$27337 ( \27714 , \27713 , \8020 );
not \U$27338 ( \27715 , \27713 );
and \U$27339 ( \27716 , \27715 , \8019 );
nor \U$27340 ( \27717 , \27714 , \27716 );
xor \U$27341 ( \27718 , \27710 , \27717 );
and \U$27342 ( \27719 , \27695 , \27718 );
and \U$27343 ( \27720 , \27689 , \27694 );
or \U$27344 ( \27721 , \27719 , \27720 );
and \U$27345 ( \27722 , \27666 , \27721 );
and \U$27346 ( \27723 , \27604 , \27665 );
or \U$27347 ( \27724 , \27722 , \27723 );
xor \U$27348 ( \27725 , \27364 , \27371 );
xor \U$27349 ( \27726 , \27725 , \27379 );
xor \U$27350 ( \27727 , \27339 , \27346 );
xor \U$27351 ( \27728 , \27727 , \27354 );
and \U$27352 ( \27729 , \27726 , \27728 );
and \U$27353 ( \27730 , \12180 , RIae785a8_113);
and \U$27354 ( \27731 , RIae783c8_109, \12178 );
nor \U$27355 ( \27732 , \27730 , \27731 );
and \U$27356 ( \27733 , \27732 , \12184 );
not \U$27357 ( \27734 , \27732 );
and \U$27358 ( \27735 , \27734 , \11827 );
nor \U$27359 ( \27736 , \27733 , \27735 );
and \U$27360 ( \27737 , \13059 , RIae78530_112);
and \U$27361 ( \27738 , RIae77c48_93, \13057 );
nor \U$27362 ( \27739 , \27737 , \27738 );
and \U$27363 ( \27740 , \27739 , \13063 );
not \U$27364 ( \27741 , \27739 );
and \U$27365 ( \27742 , \27741 , \12718 );
nor \U$27366 ( \27743 , \27740 , \27742 );
xor \U$27367 ( \27744 , \27736 , \27743 );
and \U$27368 ( \27745 , \14059 , RIae77b58_91);
and \U$27369 ( \27746 , RIae77d38_95, \14057 );
nor \U$27370 ( \27747 , \27745 , \27746 );
and \U$27371 ( \27748 , \27747 , \13502 );
not \U$27372 ( \27749 , \27747 );
and \U$27373 ( \27750 , \27749 , \14063 );
nor \U$27374 ( \27751 , \27748 , \27750 );
xor \U$27375 ( \27752 , \27744 , \27751 );
and \U$27376 ( \27753 , \9760 , RIae772e8_73);
and \U$27377 ( \27754 , RIae782d8_107, \9758 );
nor \U$27378 ( \27755 , \27753 , \27754 );
and \U$27379 ( \27756 , \27755 , \9273 );
not \U$27380 ( \27757 , \27755 );
and \U$27381 ( \27758 , \27757 , \9272 );
nor \U$27382 ( \27759 , \27756 , \27758 );
and \U$27383 ( \27760 , \10548 , RIae780f8_103);
and \U$27384 ( \27761 , RIae77f18_99, \10546 );
nor \U$27385 ( \27762 , \27760 , \27761 );
and \U$27386 ( \27763 , \27762 , \10421 );
not \U$27387 ( \27764 , \27762 );
and \U$27388 ( \27765 , \27764 , \10118 );
nor \U$27389 ( \27766 , \27763 , \27765 );
xor \U$27390 ( \27767 , \27759 , \27766 );
and \U$27391 ( \27768 , \11470 , RIae78008_101);
and \U$27392 ( \27769 , RIae781e8_105, \11468 );
nor \U$27393 ( \27770 , \27768 , \27769 );
and \U$27394 ( \27771 , \27770 , \10936 );
not \U$27395 ( \27772 , \27770 );
and \U$27396 ( \27773 , \27772 , \11474 );
nor \U$27397 ( \27774 , \27771 , \27773 );
xor \U$27398 ( \27775 , \27767 , \27774 );
and \U$27399 ( \27776 , \27752 , \27775 );
and \U$27400 ( \27777 , \15726 , RIae78878_119);
and \U$27401 ( \27778 , RIae7aab0_192, RIae78788_117);
nor \U$27402 ( \27779 , \27777 , \27778 );
and \U$27403 ( \27780 , \27779 , \14959 );
not \U$27404 ( \27781 , \27779 );
and \U$27405 ( \27782 , \27781 , RIae7aa38_191);
nor \U$27406 ( \27783 , \27780 , \27782 );
xor \U$27407 ( \27784 , \27783 , \4482 );
and \U$27408 ( \27785 , \14964 , RIae77e28_97);
and \U$27409 ( \27786 , RIae78968_121, \14962 );
nor \U$27410 ( \27787 , \27785 , \27786 );
and \U$27411 ( \27788 , \27787 , \14463 );
not \U$27412 ( \27789 , \27787 );
and \U$27413 ( \27790 , \27789 , \14462 );
nor \U$27414 ( \27791 , \27788 , \27790 );
xor \U$27415 ( \27792 , \27784 , \27791 );
xor \U$27416 ( \27793 , \27759 , \27766 );
xor \U$27417 ( \27794 , \27793 , \27774 );
and \U$27418 ( \27795 , \27792 , \27794 );
and \U$27419 ( \27796 , \27752 , \27792 );
or \U$27420 ( \27797 , \27776 , \27795 , \27796 );
xor \U$27421 ( \27798 , \27339 , \27346 );
xor \U$27422 ( \27799 , \27798 , \27354 );
and \U$27423 ( \27800 , \27797 , \27799 );
and \U$27424 ( \27801 , \27726 , \27797 );
or \U$27425 ( \27802 , \27729 , \27800 , \27801 );
xor \U$27426 ( \27803 , \27724 , \27802 );
xor \U$27427 ( \27804 , \27673 , \27680 );
and \U$27428 ( \27805 , \27804 , \27688 );
and \U$27429 ( \27806 , \27673 , \27680 );
or \U$27430 ( \27807 , \27805 , \27806 );
and \U$27431 ( \27808 , \4688 , RIae775b8_79);
and \U$27432 ( \27809 , RIae774c8_77, \4686 );
nor \U$27433 ( \27810 , \27808 , \27809 );
and \U$27434 ( \27811 , \27810 , \4481 );
not \U$27435 ( \27812 , \27810 );
and \U$27436 ( \27813 , \27812 , \4482 );
nor \U$27437 ( \27814 , \27811 , \27813 );
xor \U$27438 ( \27815 , \27807 , \27814 );
xor \U$27439 ( \27816 , \27702 , \27709 );
and \U$27440 ( \27817 , \27816 , \27717 );
and \U$27441 ( \27818 , \27702 , \27709 );
or \U$27442 ( \27819 , \27817 , \27818 );
xor \U$27443 ( \27820 , \27815 , \27819 );
xor \U$27444 ( \27821 , \27736 , \27743 );
and \U$27445 ( \27822 , \27821 , \27751 );
and \U$27446 ( \27823 , \27736 , \27743 );
or \U$27447 ( \27824 , \27822 , \27823 );
xor \U$27448 ( \27825 , \27783 , \4482 );
and \U$27449 ( \27826 , \27825 , \27791 );
and \U$27450 ( \27827 , \27783 , \4482 );
or \U$27451 ( \27828 , \27826 , \27827 );
xor \U$27452 ( \27829 , \27824 , \27828 );
xor \U$27453 ( \27830 , \27759 , \27766 );
and \U$27454 ( \27831 , \27830 , \27774 );
and \U$27455 ( \27832 , \27759 , \27766 );
or \U$27456 ( \27833 , \27831 , \27832 );
xor \U$27457 ( \27834 , \27829 , \27833 );
and \U$27458 ( \27835 , \27820 , \27834 );
xor \U$27459 ( \27836 , \27419 , \27426 );
xor \U$27460 ( \27837 , \27836 , \27434 );
xor \U$27461 ( \27838 , \27444 , \27451 );
xor \U$27462 ( \27839 , \27838 , \27459 );
xor \U$27463 ( \27840 , \27390 , \27397 );
xor \U$27464 ( \27841 , \27840 , \27405 );
xor \U$27465 ( \27842 , \27839 , \27841 );
xor \U$27466 ( \27843 , \27837 , \27842 );
xor \U$27467 ( \27844 , \27824 , \27828 );
xor \U$27468 ( \27845 , \27844 , \27833 );
and \U$27469 ( \27846 , \27843 , \27845 );
and \U$27470 ( \27847 , \27820 , \27843 );
or \U$27471 ( \27848 , \27835 , \27846 , \27847 );
and \U$27472 ( \27849 , \27803 , \27848 );
and \U$27473 ( \27850 , \27724 , \27802 );
or \U$27474 ( \27851 , \27849 , \27850 );
xor \U$27475 ( \27852 , \27437 , \27462 );
xor \U$27476 ( \27853 , \27852 , \27465 );
xor \U$27477 ( \27854 , \27357 , \27382 );
xor \U$27478 ( \27855 , \27854 , \27408 );
xor \U$27479 ( \27856 , \27853 , \27855 );
xor \U$27480 ( \27857 , \27172 , \4251 );
xor \U$27481 ( \27858 , \27857 , \27180 );
xor \U$27482 ( \27859 , \27191 , \27198 );
xor \U$27483 ( \27860 , \27859 , \27206 );
xor \U$27484 ( \27861 , \27858 , \27860 );
xor \U$27485 ( \27862 , \27119 , \27126 );
xor \U$27486 ( \27863 , \27862 , \27134 );
xor \U$27487 ( \27864 , \27322 , \27327 );
xor \U$27488 ( \27865 , \27863 , \27864 );
xor \U$27489 ( \27866 , \27861 , \27865 );
and \U$27490 ( \27867 , \27856 , \27866 );
xor \U$27491 ( \27868 , \27824 , \27828 );
and \U$27492 ( \27869 , \27868 , \27833 );
and \U$27493 ( \27870 , \27824 , \27828 );
or \U$27494 ( \27871 , \27869 , \27870 );
xor \U$27495 ( \27872 , \27807 , \27814 );
and \U$27496 ( \27873 , \27872 , \27819 );
and \U$27497 ( \27874 , \27807 , \27814 );
or \U$27498 ( \27875 , \27873 , \27874 );
xor \U$27499 ( \27876 , \27871 , \27875 );
xor \U$27500 ( \27877 , \27419 , \27426 );
xor \U$27501 ( \27878 , \27877 , \27434 );
and \U$27502 ( \27879 , \27839 , \27878 );
xor \U$27503 ( \27880 , \27419 , \27426 );
xor \U$27504 ( \27881 , \27880 , \27434 );
and \U$27505 ( \27882 , \27841 , \27881 );
and \U$27506 ( \27883 , \27839 , \27841 );
or \U$27507 ( \27884 , \27879 , \27882 , \27883 );
xor \U$27508 ( \27885 , \27876 , \27884 );
xor \U$27509 ( \27886 , \27858 , \27860 );
xor \U$27510 ( \27887 , \27886 , \27865 );
and \U$27511 ( \27888 , \27885 , \27887 );
and \U$27512 ( \27889 , \27856 , \27885 );
or \U$27513 ( \27890 , \27867 , \27888 , \27889 );
xor \U$27514 ( \27891 , \27851 , \27890 );
xor \U$27515 ( \27892 , \27332 , \27411 );
xor \U$27516 ( \27893 , \27892 , \27468 );
xor \U$27517 ( \27894 , \27165 , \27183 );
xor \U$27518 ( \27895 , \27894 , \27209 );
xor \U$27519 ( \27896 , \27893 , \27895 );
xor \U$27520 ( \27897 , \27219 , \27224 );
xor \U$27521 ( \27898 , \27897 , \27227 );
xor \U$27522 ( \27899 , \27477 , \27482 );
xor \U$27523 ( \27900 , \27898 , \27899 );
xor \U$27524 ( \27901 , \27896 , \27900 );
and \U$27525 ( \27902 , \27891 , \27901 );
and \U$27526 ( \27903 , \27851 , \27890 );
or \U$27527 ( \27904 , \27902 , \27903 );
xor \U$27528 ( \27905 , \27521 , \27904 );
xor \U$27529 ( \27906 , \27871 , \27875 );
and \U$27530 ( \27907 , \27906 , \27884 );
and \U$27531 ( \27908 , \27871 , \27875 );
or \U$27532 ( \27909 , \27907 , \27908 );
and \U$27533 ( \27910 , \27853 , \27855 );
xor \U$27534 ( \27911 , \27909 , \27910 );
xor \U$27535 ( \27912 , \27858 , \27860 );
and \U$27536 ( \27913 , \27912 , \27865 );
and \U$27537 ( \27914 , \27858 , \27860 );
or \U$27538 ( \27915 , \27913 , \27914 );
and \U$27539 ( \27916 , \27911 , \27915 );
and \U$27540 ( \27917 , \27909 , \27910 );
or \U$27541 ( \27918 , \27916 , \27917 );
xor \U$27542 ( \27919 , \27252 , \27254 );
xor \U$27543 ( \27920 , \27919 , \27259 );
xor \U$27544 ( \27921 , \27918 , \27920 );
xor \U$27545 ( \27922 , \27893 , \27895 );
and \U$27546 ( \27923 , \27922 , \27900 );
and \U$27547 ( \27924 , \27893 , \27895 );
or \U$27548 ( \27925 , \27923 , \27924 );
xor \U$27549 ( \27926 , \27921 , \27925 );
xor \U$27550 ( \27927 , \27905 , \27926 );
xor \U$27551 ( \27928 , \27909 , \27910 );
xor \U$27552 ( \27929 , \27928 , \27915 );
not \U$27553 ( \27930 , \27929 );
xor \U$27554 ( \27931 , \27851 , \27890 );
xor \U$27555 ( \27932 , \27931 , \27901 );
not \U$27556 ( \27933 , \27932 );
or \U$27557 ( \27934 , \27930 , \27933 );
or \U$27558 ( \27935 , \27932 , \27929 );
xor \U$27559 ( \27936 , \27629 , \27636 );
xor \U$27560 ( \27937 , \27936 , \27662 );
xor \U$27561 ( \27938 , \27689 , \27694 );
xor \U$27562 ( \27939 , \27938 , \27718 );
and \U$27563 ( \27940 , \27937 , \27939 );
xor \U$27564 ( \27941 , \27759 , \27766 );
xor \U$27565 ( \27942 , \27941 , \27774 );
xor \U$27566 ( \27943 , \27752 , \27792 );
xor \U$27567 ( \27944 , \27942 , \27943 );
xor \U$27568 ( \27945 , \27689 , \27694 );
xor \U$27569 ( \27946 , \27945 , \27718 );
and \U$27570 ( \27947 , \27944 , \27946 );
and \U$27571 ( \27948 , \27937 , \27944 );
or \U$27572 ( \27949 , \27940 , \27947 , \27948 );
and \U$27573 ( \27950 , \8371 , RIae76e38_63);
and \U$27574 ( \27951 , RIae76d48_61, \8369 );
nor \U$27575 ( \27952 , \27950 , \27951 );
and \U$27576 ( \27953 , \27952 , \8020 );
not \U$27577 ( \27954 , \27952 );
and \U$27578 ( \27955 , \27954 , \8019 );
nor \U$27579 ( \27956 , \27953 , \27955 );
and \U$27580 ( \27957 , \7633 , RIae77888_85);
and \U$27581 ( \27958 , RIae76f28_65, \7631 );
nor \U$27582 ( \27959 , \27957 , \27958 );
and \U$27583 ( \27960 , \27959 , \7206 );
not \U$27584 ( \27961 , \27959 );
and \U$27585 ( \27962 , \27961 , \7205 );
nor \U$27586 ( \27963 , \27960 , \27962 );
xor \U$27587 ( \27964 , \27956 , \27963 );
and \U$27588 ( \27965 , \8966 , RIae76c58_59);
and \U$27589 ( \27966 , RIae77180_70, \8964 );
nor \U$27590 ( \27967 , \27965 , \27966 );
and \U$27591 ( \27968 , \27967 , \8799 );
not \U$27592 ( \27969 , \27967 );
and \U$27593 ( \27970 , \27969 , \8789 );
nor \U$27594 ( \27971 , \27968 , \27970 );
and \U$27595 ( \27972 , \27964 , \27971 );
and \U$27596 ( \27973 , \27956 , \27963 );
or \U$27597 ( \27974 , \27972 , \27973 );
and \U$27598 ( \27975 , \6172 , RIae773d8_75);
and \U$27599 ( \27976 , RIae77a68_89, \6170 );
nor \U$27600 ( \27977 , \27975 , \27976 );
and \U$27601 ( \27978 , \27977 , \6175 );
not \U$27602 ( \27979 , \27977 );
and \U$27603 ( \27980 , \27979 , \6176 );
nor \U$27604 ( \27981 , \27978 , \27980 );
and \U$27605 ( \27982 , \6941 , RIae77978_87);
and \U$27606 ( \27983 , RIae77798_83, \6939 );
nor \U$27607 ( \27984 , \27982 , \27983 );
and \U$27608 ( \27985 , \27984 , \6945 );
not \U$27609 ( \27986 , \27984 );
and \U$27610 ( \27987 , \27986 , \6314 );
nor \U$27611 ( \27988 , \27985 , \27987 );
xor \U$27612 ( \27989 , \27981 , \27988 );
and \U$27613 ( \27990 , \5896 , RIae774c8_77);
and \U$27614 ( \27991 , RIae77720_82, \5894 );
nor \U$27615 ( \27992 , \27990 , \27991 );
and \U$27616 ( \27993 , \27992 , \5589 );
not \U$27617 ( \27994 , \27992 );
and \U$27618 ( \27995 , \27994 , \5590 );
nor \U$27619 ( \27996 , \27993 , \27995 );
and \U$27620 ( \27997 , \27989 , \27996 );
and \U$27621 ( \27998 , \27981 , \27988 );
nor \U$27622 ( \27999 , \27997 , \27998 );
xor \U$27623 ( \28000 , \27974 , \27999 );
xor \U$27624 ( \28001 , \27644 , \27651 );
xor \U$27625 ( \28002 , \28001 , \27659 );
and \U$27626 ( \28003 , \28000 , \28002 );
and \U$27627 ( \28004 , \27974 , \27999 );
or \U$27628 ( \28005 , \28003 , \28004 );
and \U$27629 ( \28006 , \11470 , RIae780f8_103);
and \U$27630 ( \28007 , RIae77f18_99, \11468 );
nor \U$27631 ( \28008 , \28006 , \28007 );
and \U$27632 ( \28009 , \28008 , \10936 );
not \U$27633 ( \28010 , \28008 );
and \U$27634 ( \28011 , \28010 , \11474 );
nor \U$27635 ( \28012 , \28009 , \28011 );
and \U$27636 ( \28013 , \9760 , RIae77018_67);
and \U$27637 ( \28014 , RIae771f8_71, \9758 );
nor \U$27638 ( \28015 , \28013 , \28014 );
and \U$27639 ( \28016 , \28015 , \9273 );
not \U$27640 ( \28017 , \28015 );
and \U$27641 ( \28018 , \28017 , \9764 );
nor \U$27642 ( \28019 , \28016 , \28018 );
xor \U$27643 ( \28020 , \28012 , \28019 );
and \U$27644 ( \28021 , \10548 , RIae772e8_73);
and \U$27645 ( \28022 , RIae782d8_107, \10546 );
nor \U$27646 ( \28023 , \28021 , \28022 );
and \U$27647 ( \28024 , \28023 , \10421 );
not \U$27648 ( \28025 , \28023 );
and \U$27649 ( \28026 , \28025 , \10118 );
nor \U$27650 ( \28027 , \28024 , \28026 );
and \U$27651 ( \28028 , \28020 , \28027 );
and \U$27652 ( \28029 , \28012 , \28019 );
or \U$27653 ( \28030 , \28028 , \28029 );
and \U$27654 ( \28031 , \15726 , RIae77e28_97);
and \U$27655 ( \28032 , RIae7aab0_192, RIae78968_121);
nor \U$27656 ( \28033 , \28031 , \28032 );
and \U$27657 ( \28034 , \28033 , \14959 );
not \U$27658 ( \28035 , \28033 );
and \U$27659 ( \28036 , \28035 , RIae7aa38_191);
nor \U$27660 ( \28037 , \28034 , \28036 );
xor \U$27661 ( \28038 , \28037 , \5403 );
and \U$27662 ( \28039 , \14964 , RIae77b58_91);
and \U$27663 ( \28040 , RIae77d38_95, \14962 );
nor \U$27664 ( \28041 , \28039 , \28040 );
or \U$27665 ( \28042 , \28041 , \14462 );
nand \U$27666 ( \28043 , \14462 , \28041 );
nand \U$27667 ( \28044 , \28042 , \28043 );
and \U$27668 ( \28045 , \28038 , \28044 );
and \U$27669 ( \28046 , \28037 , \5403 );
or \U$27670 ( \28047 , \28045 , \28046 );
xor \U$27671 ( \28048 , \28030 , \28047 );
and \U$27672 ( \28049 , \13059 , RIae785a8_113);
and \U$27673 ( \28050 , RIae783c8_109, \13057 );
nor \U$27674 ( \28051 , \28049 , \28050 );
and \U$27675 ( \28052 , \28051 , \13063 );
not \U$27676 ( \28053 , \28051 );
and \U$27677 ( \28054 , \28053 , \12718 );
nor \U$27678 ( \28055 , \28052 , \28054 );
and \U$27679 ( \28056 , \12180 , RIae78008_101);
and \U$27680 ( \28057 , RIae781e8_105, \12178 );
nor \U$27681 ( \28058 , \28056 , \28057 );
and \U$27682 ( \28059 , \28058 , \12184 );
not \U$27683 ( \28060 , \28058 );
and \U$27684 ( \28061 , \28060 , \11827 );
nor \U$27685 ( \28062 , \28059 , \28061 );
xor \U$27686 ( \28063 , \28055 , \28062 );
and \U$27687 ( \28064 , \14059 , RIae78530_112);
and \U$27688 ( \28065 , RIae77c48_93, \14057 );
nor \U$27689 ( \28066 , \28064 , \28065 );
and \U$27690 ( \28067 , \28066 , \13502 );
not \U$27691 ( \28068 , \28066 );
and \U$27692 ( \28069 , \28068 , \14063 );
nor \U$27693 ( \28070 , \28067 , \28069 );
and \U$27694 ( \28071 , \28063 , \28070 );
and \U$27695 ( \28072 , \28055 , \28062 );
or \U$27696 ( \28073 , \28071 , \28072 );
and \U$27697 ( \28074 , \28048 , \28073 );
and \U$27698 ( \28075 , \28030 , \28047 );
or \U$27699 ( \28076 , \28074 , \28075 );
xor \U$27700 ( \28077 , \28005 , \28076 );
not \U$27701 ( \28078 , \27555 );
xor \U$27702 ( \28079 , \27573 , \27563 );
not \U$27703 ( \28080 , \28079 );
or \U$27704 ( \28081 , \28078 , \28080 );
or \U$27705 ( \28082 , \28079 , \27555 );
nand \U$27706 ( \28083 , \28081 , \28082 );
xor \U$27707 ( \28084 , \27611 , \27618 );
xor \U$27708 ( \28085 , \28084 , \27626 );
xor \U$27709 ( \28086 , \28083 , \28085 );
not \U$27710 ( \28087 , \27528 );
xor \U$27711 ( \28088 , \27536 , \27546 );
not \U$27712 ( \28089 , \28088 );
or \U$27713 ( \28090 , \28087 , \28089 );
or \U$27714 ( \28091 , \28088 , \27528 );
nand \U$27715 ( \28092 , \28090 , \28091 );
and \U$27716 ( \28093 , \28086 , \28092 );
and \U$27717 ( \28094 , \28083 , \28085 );
or \U$27718 ( \28095 , \28093 , \28094 );
and \U$27719 ( \28096 , \28077 , \28095 );
and \U$27720 ( \28097 , \28005 , \28076 );
or \U$27721 ( \28098 , \28096 , \28097 );
xor \U$27722 ( \28099 , \27949 , \28098 );
xor \U$27723 ( \28100 , \27824 , \27828 );
xor \U$27724 ( \28101 , \28100 , \27833 );
xor \U$27725 ( \28102 , \27820 , \27843 );
xor \U$27726 ( \28103 , \28101 , \28102 );
and \U$27727 ( \28104 , \28099 , \28103 );
and \U$27728 ( \28105 , \27949 , \28098 );
or \U$27729 ( \28106 , \28104 , \28105 );
xor \U$27730 ( \28107 , \27604 , \27665 );
xor \U$27731 ( \28108 , \28107 , \27721 );
xor \U$27732 ( \28109 , \27339 , \27346 );
xor \U$27733 ( \28110 , \28109 , \27354 );
xor \U$27734 ( \28111 , \27726 , \27797 );
xor \U$27735 ( \28112 , \28110 , \28111 );
and \U$27736 ( \28113 , \28108 , \28112 );
xor \U$27737 ( \28114 , \28106 , \28113 );
xor \U$27738 ( \28115 , \27858 , \27860 );
xor \U$27739 ( \28116 , \28115 , \27865 );
xor \U$27740 ( \28117 , \27856 , \27885 );
xor \U$27741 ( \28118 , \28116 , \28117 );
and \U$27742 ( \28119 , \28114 , \28118 );
and \U$27743 ( \28120 , \28106 , \28113 );
or \U$27744 ( \28121 , \28119 , \28120 );
nand \U$27745 ( \28122 , \27935 , \28121 );
nand \U$27746 ( \28123 , \27934 , \28122 );
and \U$27747 ( \28124 , \27927 , \28123 );
xor \U$27748 ( \28125 , \28123 , \27927 );
xnor \U$27749 ( \28126 , \27929 , \28121 );
not \U$27750 ( \28127 , \28126 );
not \U$27751 ( \28128 , \27932 );
and \U$27752 ( \28129 , \28127 , \28128 );
and \U$27753 ( \28130 , \28126 , \27932 );
nor \U$27754 ( \28131 , \28129 , \28130 );
xor \U$27755 ( \28132 , \28106 , \28113 );
xor \U$27756 ( \28133 , \28132 , \28118 );
xor \U$27757 ( \28134 , \27724 , \27802 );
xor \U$27758 ( \28135 , \28134 , \27848 );
xor \U$27759 ( \28136 , \28133 , \28135 );
xor \U$27760 ( \28137 , \27583 , \27590 );
xor \U$27761 ( \28138 , \28137 , \27598 );
xor \U$27762 ( \28139 , \27974 , \27999 );
xor \U$27763 ( \28140 , \28139 , \28002 );
and \U$27764 ( \28141 , \28138 , \28140 );
xor \U$27765 ( \28142 , \28083 , \28085 );
xor \U$27766 ( \28143 , \28142 , \28092 );
xor \U$27767 ( \28144 , \27974 , \27999 );
xor \U$27768 ( \28145 , \28144 , \28002 );
and \U$27769 ( \28146 , \28143 , \28145 );
and \U$27770 ( \28147 , \28138 , \28143 );
or \U$27771 ( \28148 , \28141 , \28146 , \28147 );
not \U$27772 ( \28149 , \28148 );
xor \U$27773 ( \28150 , \27548 , \27575 );
xor \U$27774 ( \28151 , \28150 , \27601 );
or \U$27775 ( \28152 , \28149 , \28151 );
not \U$27776 ( \28153 , \28151 );
not \U$27777 ( \28154 , \28149 );
or \U$27778 ( \28155 , \28153 , \28154 );
and \U$27779 ( \28156 , \8966 , RIae76d48_61);
and \U$27780 ( \28157 , RIae76c58_59, \8964 );
nor \U$27781 ( \28158 , \28156 , \28157 );
and \U$27782 ( \28159 , \28158 , \8799 );
not \U$27783 ( \28160 , \28158 );
and \U$27784 ( \28161 , \28160 , \8789 );
nor \U$27785 ( \28162 , \28159 , \28161 );
and \U$27786 ( \28163 , \9760 , RIae77180_70);
and \U$27787 ( \28164 , RIae77018_67, \9758 );
nor \U$27788 ( \28165 , \28163 , \28164 );
and \U$27789 ( \28166 , \28165 , \9273 );
not \U$27790 ( \28167 , \28165 );
and \U$27791 ( \28168 , \28167 , \9764 );
nor \U$27792 ( \28169 , \28166 , \28168 );
xor \U$27793 ( \28170 , \28162 , \28169 );
and \U$27794 ( \28171 , \10548 , RIae771f8_71);
and \U$27795 ( \28172 , RIae772e8_73, \10546 );
nor \U$27796 ( \28173 , \28171 , \28172 );
and \U$27797 ( \28174 , \28173 , \10421 );
not \U$27798 ( \28175 , \28173 );
and \U$27799 ( \28176 , \28175 , \10118 );
nor \U$27800 ( \28177 , \28174 , \28176 );
and \U$27801 ( \28178 , \28170 , \28177 );
and \U$27802 ( \28179 , \28162 , \28169 );
or \U$27803 ( \28180 , \28178 , \28179 );
and \U$27804 ( \28181 , \14059 , RIae783c8_109);
and \U$27805 ( \28182 , RIae78530_112, \14057 );
nor \U$27806 ( \28183 , \28181 , \28182 );
and \U$27807 ( \28184 , \28183 , \13502 );
not \U$27808 ( \28185 , \28183 );
and \U$27809 ( \28186 , \28185 , \14063 );
nor \U$27810 ( \28187 , \28184 , \28186 );
and \U$27811 ( \28188 , \15726 , RIae77d38_95);
and \U$27812 ( \28189 , RIae7aab0_192, RIae77e28_97);
nor \U$27813 ( \28190 , \28188 , \28189 );
and \U$27814 ( \28191 , \28190 , \14959 );
not \U$27815 ( \28192 , \28190 );
and \U$27816 ( \28193 , \28192 , RIae7aa38_191);
nor \U$27817 ( \28194 , \28191 , \28193 );
xor \U$27818 ( \28195 , \28187 , \28194 );
and \U$27819 ( \28196 , \14964 , RIae77c48_93);
and \U$27820 ( \28197 , RIae77b58_91, \14962 );
nor \U$27821 ( \28198 , \28196 , \28197 );
and \U$27822 ( \28199 , \28198 , \14463 );
not \U$27823 ( \28200 , \28198 );
and \U$27824 ( \28201 , \28200 , \14462 );
nor \U$27825 ( \28202 , \28199 , \28201 );
and \U$27826 ( \28203 , \28195 , \28202 );
and \U$27827 ( \28204 , \28187 , \28194 );
or \U$27828 ( \28205 , \28203 , \28204 );
xor \U$27829 ( \28206 , \28180 , \28205 );
and \U$27830 ( \28207 , \11470 , RIae782d8_107);
and \U$27831 ( \28208 , RIae780f8_103, \11468 );
nor \U$27832 ( \28209 , \28207 , \28208 );
and \U$27833 ( \28210 , \28209 , \10936 );
not \U$27834 ( \28211 , \28209 );
and \U$27835 ( \28212 , \28211 , \11474 );
nor \U$27836 ( \28213 , \28210 , \28212 );
and \U$27837 ( \28214 , \12180 , RIae77f18_99);
and \U$27838 ( \28215 , RIae78008_101, \12178 );
nor \U$27839 ( \28216 , \28214 , \28215 );
and \U$27840 ( \28217 , \28216 , \12184 );
not \U$27841 ( \28218 , \28216 );
and \U$27842 ( \28219 , \28218 , \11827 );
nor \U$27843 ( \28220 , \28217 , \28219 );
xor \U$27844 ( \28221 , \28213 , \28220 );
and \U$27845 ( \28222 , \13059 , RIae781e8_105);
and \U$27846 ( \28223 , RIae785a8_113, \13057 );
nor \U$27847 ( \28224 , \28222 , \28223 );
and \U$27848 ( \28225 , \28224 , \13063 );
not \U$27849 ( \28226 , \28224 );
and \U$27850 ( \28227 , \28226 , \12718 );
nor \U$27851 ( \28228 , \28225 , \28227 );
and \U$27852 ( \28229 , \28221 , \28228 );
and \U$27853 ( \28230 , \28213 , \28220 );
or \U$27854 ( \28231 , \28229 , \28230 );
and \U$27855 ( \28232 , \28206 , \28231 );
and \U$27856 ( \28233 , \28180 , \28205 );
nor \U$27857 ( \28234 , \28232 , \28233 );
xor \U$27858 ( \28235 , \28055 , \28062 );
xor \U$27859 ( \28236 , \28235 , \28070 );
xor \U$27860 ( \28237 , \28012 , \28019 );
xor \U$27861 ( \28238 , \28237 , \28027 );
and \U$27862 ( \28239 , \28236 , \28238 );
xor \U$27863 ( \28240 , \27956 , \27963 );
xor \U$27864 ( \28241 , \28240 , \27971 );
xor \U$27865 ( \28242 , \28012 , \28019 );
xor \U$27866 ( \28243 , \28242 , \28027 );
and \U$27867 ( \28244 , \28241 , \28243 );
and \U$27868 ( \28245 , \28236 , \28241 );
or \U$27869 ( \28246 , \28239 , \28244 , \28245 );
not \U$27870 ( \28247 , \28246 );
xor \U$27871 ( \28248 , \28234 , \28247 );
xor \U$27872 ( \28249 , \27981 , \27988 );
xor \U$27873 ( \28250 , \28249 , \27996 );
not \U$27874 ( \28251 , \28250 );
nand \U$27875 ( \28252 , RIae775b8_79, \5397 );
and \U$27876 ( \28253 , \28252 , \5403 );
not \U$27877 ( \28254 , \28252 );
and \U$27878 ( \28255 , \28254 , \5016 );
nor \U$27879 ( \28256 , \28253 , \28255 );
not \U$27880 ( \28257 , \28256 );
and \U$27881 ( \28258 , \28251 , \28257 );
and \U$27882 ( \28259 , \28250 , \28256 );
and \U$27883 ( \28260 , \7633 , RIae77798_83);
and \U$27884 ( \28261 , RIae77888_85, \7631 );
nor \U$27885 ( \28262 , \28260 , \28261 );
and \U$27886 ( \28263 , \28262 , \7206 );
not \U$27887 ( \28264 , \28262 );
and \U$27888 ( \28265 , \28264 , \7205 );
nor \U$27889 ( \28266 , \28263 , \28265 );
and \U$27890 ( \28267 , \8371 , RIae76f28_65);
and \U$27891 ( \28268 , RIae76e38_63, \8369 );
nor \U$27892 ( \28269 , \28267 , \28268 );
and \U$27893 ( \28270 , \28269 , \8020 );
not \U$27894 ( \28271 , \28269 );
and \U$27895 ( \28272 , \28271 , \8019 );
nor \U$27896 ( \28273 , \28270 , \28272 );
xor \U$27897 ( \28274 , \28266 , \28273 );
and \U$27898 ( \28275 , \6941 , RIae77a68_89);
and \U$27899 ( \28276 , RIae77978_87, \6939 );
nor \U$27900 ( \28277 , \28275 , \28276 );
and \U$27901 ( \28278 , \28277 , \6314 );
not \U$27902 ( \28279 , \28277 );
and \U$27903 ( \28280 , \28279 , \6945 );
nor \U$27904 ( \28281 , \28278 , \28280 );
and \U$27905 ( \28282 , \28274 , \28281 );
and \U$27906 ( \28283 , \28266 , \28273 );
nor \U$27907 ( \28284 , \28282 , \28283 );
nor \U$27908 ( \28285 , \28259 , \28284 );
nor \U$27909 ( \28286 , \28258 , \28285 );
and \U$27910 ( \28287 , \28248 , \28286 );
and \U$27911 ( \28288 , \28234 , \28247 );
nor \U$27912 ( \28289 , \28287 , \28288 );
nand \U$27913 ( \28290 , \28155 , \28289 );
nand \U$27914 ( \28291 , \28152 , \28290 );
xor \U$27915 ( \28292 , \28108 , \28112 );
xor \U$27916 ( \28293 , \28291 , \28292 );
xor \U$27917 ( \28294 , \27949 , \28098 );
xor \U$27918 ( \28295 , \28294 , \28103 );
and \U$27919 ( \28296 , \28293 , \28295 );
and \U$27920 ( \28297 , \28291 , \28292 );
or \U$27921 ( \28298 , \28296 , \28297 );
and \U$27922 ( \28299 , \28136 , \28298 );
and \U$27923 ( \28300 , \28133 , \28135 );
nor \U$27924 ( \28301 , \28299 , \28300 );
or \U$27925 ( \28302 , \28131 , \28301 );
xnor \U$27926 ( \28303 , \28301 , \28131 );
xor \U$27927 ( \28304 , \28133 , \28135 );
xor \U$27928 ( \28305 , \28304 , \28298 );
xor \U$27929 ( \28306 , \28234 , \28247 );
xor \U$27930 ( \28307 , \28306 , \28286 );
not \U$27931 ( \28308 , \28307 );
xor \U$27932 ( \28309 , \27974 , \27999 );
xor \U$27933 ( \28310 , \28309 , \28002 );
xor \U$27934 ( \28311 , \28138 , \28143 );
xor \U$27935 ( \28312 , \28310 , \28311 );
nand \U$27936 ( \28313 , \28308 , \28312 );
not \U$27937 ( \28314 , \28313 );
xor \U$27938 ( \28315 , \27689 , \27694 );
xor \U$27939 ( \28316 , \28315 , \27718 );
xor \U$27940 ( \28317 , \27937 , \27944 );
xor \U$27941 ( \28318 , \28316 , \28317 );
and \U$27942 ( \28319 , \28314 , \28318 );
and \U$27943 ( \28320 , \9760 , RIae76c58_59);
and \U$27944 ( \28321 , RIae77180_70, \9758 );
nor \U$27945 ( \28322 , \28320 , \28321 );
and \U$27946 ( \28323 , \28322 , \9273 );
not \U$27947 ( \28324 , \28322 );
and \U$27948 ( \28325 , \28324 , \9764 );
nor \U$27949 ( \28326 , \28323 , \28325 );
and \U$27950 ( \28327 , \10548 , RIae77018_67);
and \U$27951 ( \28328 , RIae771f8_71, \10546 );
nor \U$27952 ( \28329 , \28327 , \28328 );
and \U$27953 ( \28330 , \28329 , \10421 );
not \U$27954 ( \28331 , \28329 );
and \U$27955 ( \28332 , \28331 , \10118 );
nor \U$27956 ( \28333 , \28330 , \28332 );
xor \U$27957 ( \28334 , \28326 , \28333 );
and \U$27958 ( \28335 , \11470 , RIae772e8_73);
and \U$27959 ( \28336 , RIae782d8_107, \11468 );
nor \U$27960 ( \28337 , \28335 , \28336 );
and \U$27961 ( \28338 , \28337 , \10936 );
not \U$27962 ( \28339 , \28337 );
and \U$27963 ( \28340 , \28339 , \11474 );
nor \U$27964 ( \28341 , \28338 , \28340 );
and \U$27965 ( \28342 , \28334 , \28341 );
and \U$27966 ( \28343 , \28326 , \28333 );
or \U$27967 ( \28344 , \28342 , \28343 );
and \U$27968 ( \28345 , \15726 , RIae77b58_91);
and \U$27969 ( \28346 , RIae7aab0_192, RIae77d38_95);
nor \U$27970 ( \28347 , \28345 , \28346 );
and \U$27971 ( \28348 , \28347 , \14959 );
not \U$27972 ( \28349 , \28347 );
and \U$27973 ( \28350 , \28349 , RIae7aa38_191);
nor \U$27974 ( \28351 , \28348 , \28350 );
xor \U$27975 ( \28352 , \28351 , \5589 );
and \U$27976 ( \28353 , \14964 , RIae78530_112);
and \U$27977 ( \28354 , RIae77c48_93, \14962 );
nor \U$27978 ( \28355 , \28353 , \28354 );
and \U$27979 ( \28356 , \28355 , \14463 );
not \U$27980 ( \28357 , \28355 );
and \U$27981 ( \28358 , \28357 , \14462 );
nor \U$27982 ( \28359 , \28356 , \28358 );
and \U$27983 ( \28360 , \28352 , \28359 );
and \U$27984 ( \28361 , \28351 , \5589 );
or \U$27985 ( \28362 , \28360 , \28361 );
xor \U$27986 ( \28363 , \28344 , \28362 );
and \U$27987 ( \28364 , \14059 , RIae785a8_113);
and \U$27988 ( \28365 , RIae783c8_109, \14057 );
nor \U$27989 ( \28366 , \28364 , \28365 );
and \U$27990 ( \28367 , \28366 , \13502 );
not \U$27991 ( \28368 , \28366 );
and \U$27992 ( \28369 , \28368 , \14063 );
nor \U$27993 ( \28370 , \28367 , \28369 );
and \U$27994 ( \28371 , \12180 , RIae780f8_103);
and \U$27995 ( \28372 , RIae77f18_99, \12178 );
nor \U$27996 ( \28373 , \28371 , \28372 );
and \U$27997 ( \28374 , \28373 , \12184 );
not \U$27998 ( \28375 , \28373 );
and \U$27999 ( \28376 , \28375 , \11827 );
nor \U$28000 ( \28377 , \28374 , \28376 );
xor \U$28001 ( \28378 , \28370 , \28377 );
and \U$28002 ( \28379 , \13059 , RIae78008_101);
and \U$28003 ( \28380 , RIae781e8_105, \13057 );
nor \U$28004 ( \28381 , \28379 , \28380 );
and \U$28005 ( \28382 , \28381 , \13063 );
not \U$28006 ( \28383 , \28381 );
and \U$28007 ( \28384 , \28383 , \12718 );
nor \U$28008 ( \28385 , \28382 , \28384 );
and \U$28009 ( \28386 , \28378 , \28385 );
and \U$28010 ( \28387 , \28370 , \28377 );
or \U$28011 ( \28388 , \28386 , \28387 );
and \U$28012 ( \28389 , \28363 , \28388 );
and \U$28013 ( \28390 , \28344 , \28362 );
or \U$28014 ( \28391 , \28389 , \28390 );
and \U$28015 ( \28392 , \6941 , RIae773d8_75);
and \U$28016 ( \28393 , RIae77a68_89, \6939 );
nor \U$28017 ( \28394 , \28392 , \28393 );
and \U$28018 ( \28395 , \28394 , \6314 );
not \U$28019 ( \28396 , \28394 );
and \U$28020 ( \28397 , \28396 , \6945 );
nor \U$28021 ( \28398 , \28395 , \28397 );
nand \U$28022 ( \28399 , RIae775b8_79, \5894 );
and \U$28023 ( \28400 , \28399 , \5590 );
not \U$28024 ( \28401 , \28399 );
and \U$28025 ( \28402 , \28401 , \5589 );
nor \U$28026 ( \28403 , \28400 , \28402 );
xor \U$28027 ( \28404 , \28398 , \28403 );
and \U$28028 ( \28405 , \6172 , RIae774c8_77);
and \U$28029 ( \28406 , RIae77720_82, \6170 );
nor \U$28030 ( \28407 , \28405 , \28406 );
and \U$28031 ( \28408 , \28407 , \6176 );
not \U$28032 ( \28409 , \28407 );
and \U$28033 ( \28410 , \28409 , \6175 );
nor \U$28034 ( \28411 , \28408 , \28410 );
and \U$28035 ( \28412 , \28404 , \28411 );
and \U$28036 ( \28413 , \28398 , \28403 );
or \U$28037 ( \28414 , \28412 , \28413 );
and \U$28038 ( \28415 , \6172 , RIae77720_82);
and \U$28039 ( \28416 , RIae773d8_75, \6170 );
nor \U$28040 ( \28417 , \28415 , \28416 );
and \U$28041 ( \28418 , \28417 , \6176 );
not \U$28042 ( \28419 , \28417 );
and \U$28043 ( \28420 , \28419 , \6175 );
nor \U$28044 ( \28421 , \28418 , \28420 );
xor \U$28045 ( \28422 , \28414 , \28421 );
and \U$28046 ( \28423 , \8966 , RIae76e38_63);
and \U$28047 ( \28424 , RIae76d48_61, \8964 );
nor \U$28048 ( \28425 , \28423 , \28424 );
and \U$28049 ( \28426 , \28425 , \8799 );
not \U$28050 ( \28427 , \28425 );
and \U$28051 ( \28428 , \28427 , \8789 );
nor \U$28052 ( \28429 , \28426 , \28428 );
and \U$28053 ( \28430 , \7633 , RIae77978_87);
and \U$28054 ( \28431 , RIae77798_83, \7631 );
nor \U$28055 ( \28432 , \28430 , \28431 );
and \U$28056 ( \28433 , \28432 , \7206 );
not \U$28057 ( \28434 , \28432 );
and \U$28058 ( \28435 , \28434 , \7205 );
nor \U$28059 ( \28436 , \28433 , \28435 );
xor \U$28060 ( \28437 , \28429 , \28436 );
and \U$28061 ( \28438 , \8371 , RIae77888_85);
and \U$28062 ( \28439 , RIae76f28_65, \8369 );
nor \U$28063 ( \28440 , \28438 , \28439 );
and \U$28064 ( \28441 , \28440 , \8020 );
not \U$28065 ( \28442 , \28440 );
and \U$28066 ( \28443 , \28442 , \8019 );
nor \U$28067 ( \28444 , \28441 , \28443 );
and \U$28068 ( \28445 , \28437 , \28444 );
and \U$28069 ( \28446 , \28429 , \28436 );
or \U$28070 ( \28447 , \28445 , \28446 );
and \U$28071 ( \28448 , \28422 , \28447 );
and \U$28072 ( \28449 , \28414 , \28421 );
or \U$28073 ( \28450 , \28448 , \28449 );
xor \U$28074 ( \28451 , \28391 , \28450 );
and \U$28075 ( \28452 , \5896 , RIae775b8_79);
and \U$28076 ( \28453 , RIae774c8_77, \5894 );
nor \U$28077 ( \28454 , \28452 , \28453 );
and \U$28078 ( \28455 , \28454 , \5590 );
not \U$28079 ( \28456 , \28454 );
and \U$28080 ( \28457 , \28456 , \5589 );
nor \U$28081 ( \28458 , \28455 , \28457 );
xor \U$28082 ( \28459 , \28162 , \28169 );
xor \U$28083 ( \28460 , \28459 , \28177 );
and \U$28084 ( \28461 , \28458 , \28460 );
xor \U$28085 ( \28462 , \28266 , \28273 );
xor \U$28086 ( \28463 , \28462 , \28281 );
xor \U$28087 ( \28464 , \28162 , \28169 );
xor \U$28088 ( \28465 , \28464 , \28177 );
and \U$28089 ( \28466 , \28463 , \28465 );
and \U$28090 ( \28467 , \28458 , \28463 );
or \U$28091 ( \28468 , \28461 , \28466 , \28467 );
and \U$28092 ( \28469 , \28451 , \28468 );
and \U$28093 ( \28470 , \28391 , \28450 );
or \U$28094 ( \28471 , \28469 , \28470 );
xor \U$28095 ( \28472 , \28030 , \28047 );
xor \U$28096 ( \28473 , \28472 , \28073 );
xor \U$28097 ( \28474 , \28471 , \28473 );
not \U$28098 ( \28475 , \28250 );
xor \U$28099 ( \28476 , \28256 , \28284 );
not \U$28100 ( \28477 , \28476 );
or \U$28101 ( \28478 , \28475 , \28477 );
or \U$28102 ( \28479 , \28476 , \28250 );
nand \U$28103 ( \28480 , \28478 , \28479 );
xor \U$28104 ( \28481 , \28037 , \5403 );
xor \U$28105 ( \28482 , \28481 , \28044 );
xor \U$28106 ( \28483 , \28480 , \28482 );
xor \U$28107 ( \28484 , \28012 , \28019 );
xor \U$28108 ( \28485 , \28484 , \28027 );
xor \U$28109 ( \28486 , \28236 , \28241 );
xor \U$28110 ( \28487 , \28485 , \28486 );
and \U$28111 ( \28488 , \28483 , \28487 );
and \U$28112 ( \28489 , \28480 , \28482 );
or \U$28113 ( \28490 , \28488 , \28489 );
and \U$28114 ( \28491 , \28474 , \28490 );
and \U$28115 ( \28492 , \28471 , \28473 );
or \U$28116 ( \28493 , \28491 , \28492 );
not \U$28117 ( \28494 , \28318 );
nand \U$28118 ( \28495 , \28494 , \28313 );
and \U$28119 ( \28496 , \28493 , \28495 );
nor \U$28120 ( \28497 , \28319 , \28496 );
not \U$28121 ( \28498 , \28289 );
not \U$28122 ( \28499 , \28149 );
or \U$28123 ( \28500 , \28498 , \28499 );
or \U$28124 ( \28501 , \28149 , \28289 );
nand \U$28125 ( \28502 , \28500 , \28501 );
not \U$28126 ( \28503 , \28502 );
not \U$28127 ( \28504 , \28151 );
and \U$28128 ( \28505 , \28503 , \28504 );
and \U$28129 ( \28506 , \28502 , \28151 );
nor \U$28130 ( \28507 , \28505 , \28506 );
not \U$28131 ( \28508 , \28507 );
xor \U$28132 ( \28509 , \28005 , \28076 );
xor \U$28133 ( \28510 , \28509 , \28095 );
nand \U$28134 ( \28511 , \28508 , \28510 );
or \U$28135 ( \28512 , \28497 , \28511 );
not \U$28136 ( \28513 , \28511 );
not \U$28137 ( \28514 , \28497 );
or \U$28138 ( \28515 , \28513 , \28514 );
xor \U$28139 ( \28516 , \28291 , \28292 );
xor \U$28140 ( \28517 , \28516 , \28295 );
nand \U$28141 ( \28518 , \28515 , \28517 );
nand \U$28142 ( \28519 , \28512 , \28518 );
and \U$28143 ( \28520 , \28305 , \28519 );
xor \U$28144 ( \28521 , \28519 , \28305 );
not \U$28145 ( \28522 , \28517 );
xnor \U$28146 ( \28523 , \28511 , \28497 );
not \U$28147 ( \28524 , \28523 );
and \U$28148 ( \28525 , \28522 , \28524 );
and \U$28149 ( \28526 , \28523 , \28517 );
nor \U$28150 ( \28527 , \28525 , \28526 );
not \U$28151 ( \28528 , \28510 );
not \U$28152 ( \28529 , \28507 );
or \U$28153 ( \28530 , \28528 , \28529 );
or \U$28154 ( \28531 , \28507 , \28510 );
nand \U$28155 ( \28532 , \28530 , \28531 );
not \U$28156 ( \28533 , \28307 );
not \U$28157 ( \28534 , \28312 );
or \U$28158 ( \28535 , \28533 , \28534 );
or \U$28159 ( \28536 , \28312 , \28307 );
nand \U$28160 ( \28537 , \28535 , \28536 );
xor \U$28161 ( \28538 , \28213 , \28220 );
xor \U$28162 ( \28539 , \28538 , \28228 );
xor \U$28163 ( \28540 , \28187 , \28194 );
xor \U$28164 ( \28541 , \28540 , \28202 );
xor \U$28165 ( \28542 , \28539 , \28541 );
xor \U$28166 ( \28543 , \28162 , \28169 );
xor \U$28167 ( \28544 , \28543 , \28177 );
xor \U$28168 ( \28545 , \28458 , \28463 );
xor \U$28169 ( \28546 , \28544 , \28545 );
and \U$28170 ( \28547 , \28542 , \28546 );
and \U$28171 ( \28548 , \28539 , \28541 );
or \U$28172 ( \28549 , \28547 , \28548 );
xor \U$28173 ( \28550 , \28180 , \28205 );
xor \U$28174 ( \28551 , \28550 , \28231 );
xor \U$28175 ( \28552 , \28549 , \28551 );
xor \U$28176 ( \28553 , \28398 , \28403 );
xor \U$28177 ( \28554 , \28553 , \28411 );
and \U$28178 ( \28555 , \6941 , RIae77720_82);
and \U$28179 ( \28556 , RIae773d8_75, \6939 );
nor \U$28180 ( \28557 , \28555 , \28556 );
and \U$28181 ( \28558 , \28557 , \6945 );
not \U$28182 ( \28559 , \28557 );
and \U$28183 ( \28560 , \28559 , \6314 );
nor \U$28184 ( \28561 , \28558 , \28560 );
and \U$28185 ( \28562 , \8371 , RIae77798_83);
and \U$28186 ( \28563 , RIae77888_85, \8369 );
nor \U$28187 ( \28564 , \28562 , \28563 );
and \U$28188 ( \28565 , \28564 , \8019 );
not \U$28189 ( \28566 , \28564 );
and \U$28190 ( \28567 , \28566 , \8020 );
nor \U$28191 ( \28568 , \28565 , \28567 );
or \U$28192 ( \28569 , \28561 , \28568 );
not \U$28193 ( \28570 , \28568 );
not \U$28194 ( \28571 , \28561 );
or \U$28195 ( \28572 , \28570 , \28571 );
and \U$28196 ( \28573 , \7633 , RIae77a68_89);
and \U$28197 ( \28574 , RIae77978_87, \7631 );
nor \U$28198 ( \28575 , \28573 , \28574 );
and \U$28199 ( \28576 , \28575 , \7206 );
not \U$28200 ( \28577 , \28575 );
and \U$28201 ( \28578 , \28577 , \7205 );
nor \U$28202 ( \28579 , \28576 , \28578 );
nand \U$28203 ( \28580 , \28572 , \28579 );
nand \U$28204 ( \28581 , \28569 , \28580 );
xor \U$28205 ( \28582 , \28554 , \28581 );
xor \U$28206 ( \28583 , \28429 , \28436 );
xor \U$28207 ( \28584 , \28583 , \28444 );
and \U$28208 ( \28585 , \28582 , \28584 );
and \U$28209 ( \28586 , \28554 , \28581 );
or \U$28210 ( \28587 , \28585 , \28586 );
and \U$28211 ( \28588 , \12180 , RIae782d8_107);
and \U$28212 ( \28589 , RIae780f8_103, \12178 );
nor \U$28213 ( \28590 , \28588 , \28589 );
and \U$28214 ( \28591 , \28590 , \11827 );
not \U$28215 ( \28592 , \28590 );
and \U$28216 ( \28593 , \28592 , \12184 );
nor \U$28217 ( \28594 , \28591 , \28593 );
and \U$28218 ( \28595 , \13059 , RIae77f18_99);
and \U$28219 ( \28596 , RIae78008_101, \13057 );
nor \U$28220 ( \28597 , \28595 , \28596 );
and \U$28221 ( \28598 , \28597 , \12718 );
not \U$28222 ( \28599 , \28597 );
and \U$28223 ( \28600 , \28599 , \13063 );
nor \U$28224 ( \28601 , \28598 , \28600 );
xor \U$28225 ( \28602 , \28594 , \28601 );
and \U$28226 ( \28603 , \11470 , RIae771f8_71);
and \U$28227 ( \28604 , RIae772e8_73, \11468 );
nor \U$28228 ( \28605 , \28603 , \28604 );
and \U$28229 ( \28606 , \28605 , \11474 );
not \U$28230 ( \28607 , \28605 );
and \U$28231 ( \28608 , \28607 , \10936 );
nor \U$28232 ( \28609 , \28606 , \28608 );
and \U$28233 ( \28610 , \28602 , \28609 );
and \U$28234 ( \28611 , \28594 , \28601 );
nor \U$28235 ( \28612 , \28610 , \28611 );
and \U$28236 ( \28613 , \15726 , RIae77c48_93);
and \U$28237 ( \28614 , RIae7aab0_192, RIae77b58_91);
nor \U$28238 ( \28615 , \28613 , \28614 );
and \U$28239 ( \28616 , \28615 , RIae7aa38_191);
not \U$28240 ( \28617 , \28615 );
and \U$28241 ( \28618 , \28617 , \14959 );
nor \U$28242 ( \28619 , \28616 , \28618 );
and \U$28243 ( \28620 , \14964 , RIae783c8_109);
and \U$28244 ( \28621 , RIae78530_112, \14962 );
nor \U$28245 ( \28622 , \28620 , \28621 );
and \U$28246 ( \28623 , \28622 , \14462 );
not \U$28247 ( \28624 , \28622 );
and \U$28248 ( \28625 , \28624 , \14463 );
nor \U$28249 ( \28626 , \28623 , \28625 );
xor \U$28250 ( \28627 , \28619 , \28626 );
and \U$28251 ( \28628 , \14059 , RIae781e8_105);
and \U$28252 ( \28629 , RIae785a8_113, \14057 );
nor \U$28253 ( \28630 , \28628 , \28629 );
and \U$28254 ( \28631 , \28630 , \14063 );
not \U$28255 ( \28632 , \28630 );
and \U$28256 ( \28633 , \28632 , \13502 );
nor \U$28257 ( \28634 , \28631 , \28633 );
and \U$28258 ( \28635 , \28627 , \28634 );
and \U$28259 ( \28636 , \28619 , \28626 );
nor \U$28260 ( \28637 , \28635 , \28636 );
xor \U$28261 ( \28638 , \28612 , \28637 );
and \U$28262 ( \28639 , \8966 , RIae76f28_65);
and \U$28263 ( \28640 , RIae76e38_63, \8964 );
nor \U$28264 ( \28641 , \28639 , \28640 );
and \U$28265 ( \28642 , \28641 , \8789 );
not \U$28266 ( \28643 , \28641 );
and \U$28267 ( \28644 , \28643 , \8799 );
nor \U$28268 ( \28645 , \28642 , \28644 );
and \U$28269 ( \28646 , \9760 , RIae76d48_61);
and \U$28270 ( \28647 , RIae76c58_59, \9758 );
nor \U$28271 ( \28648 , \28646 , \28647 );
and \U$28272 ( \28649 , \28648 , \9272 );
not \U$28273 ( \28650 , \28648 );
and \U$28274 ( \28651 , \28650 , \9273 );
nor \U$28275 ( \28652 , \28649 , \28651 );
or \U$28276 ( \28653 , \28645 , \28652 );
not \U$28277 ( \28654 , \28652 );
not \U$28278 ( \28655 , \28645 );
or \U$28279 ( \28656 , \28654 , \28655 );
and \U$28280 ( \28657 , \10548 , RIae77180_70);
and \U$28281 ( \28658 , RIae77018_67, \10546 );
nor \U$28282 ( \28659 , \28657 , \28658 );
and \U$28283 ( \28660 , \28659 , \10421 );
not \U$28284 ( \28661 , \28659 );
and \U$28285 ( \28662 , \28661 , \10118 );
nor \U$28286 ( \28663 , \28660 , \28662 );
nand \U$28287 ( \28664 , \28656 , \28663 );
nand \U$28288 ( \28665 , \28653 , \28664 );
and \U$28289 ( \28666 , \28638 , \28665 );
and \U$28290 ( \28667 , \28612 , \28637 );
or \U$28291 ( \28668 , \28666 , \28667 );
xor \U$28292 ( \28669 , \28587 , \28668 );
xor \U$28293 ( \28670 , \28326 , \28333 );
xor \U$28294 ( \28671 , \28670 , \28341 );
xor \U$28295 ( \28672 , \28370 , \28377 );
xor \U$28296 ( \28673 , \28672 , \28385 );
and \U$28297 ( \28674 , \28671 , \28673 );
xor \U$28298 ( \28675 , \28351 , \5589 );
xor \U$28299 ( \28676 , \28675 , \28359 );
xor \U$28300 ( \28677 , \28370 , \28377 );
xor \U$28301 ( \28678 , \28677 , \28385 );
and \U$28302 ( \28679 , \28676 , \28678 );
and \U$28303 ( \28680 , \28671 , \28676 );
or \U$28304 ( \28681 , \28674 , \28679 , \28680 );
and \U$28305 ( \28682 , \28669 , \28681 );
and \U$28306 ( \28683 , \28587 , \28668 );
or \U$28307 ( \28684 , \28682 , \28683 );
and \U$28308 ( \28685 , \28552 , \28684 );
and \U$28309 ( \28686 , \28549 , \28551 );
or \U$28310 ( \28687 , \28685 , \28686 );
xor \U$28311 ( \28688 , \28537 , \28687 );
xor \U$28312 ( \28689 , \28471 , \28473 );
xor \U$28313 ( \28690 , \28689 , \28490 );
and \U$28314 ( \28691 , \28688 , \28690 );
and \U$28315 ( \28692 , \28537 , \28687 );
or \U$28316 ( \28693 , \28691 , \28692 );
xor \U$28317 ( \28694 , \28532 , \28693 );
not \U$28318 ( \28695 , \28318 );
not \U$28319 ( \28696 , \28493 );
not \U$28320 ( \28697 , \28313 );
and \U$28321 ( \28698 , \28696 , \28697 );
and \U$28322 ( \28699 , \28493 , \28313 );
nor \U$28323 ( \28700 , \28698 , \28699 );
not \U$28324 ( \28701 , \28700 );
or \U$28325 ( \28702 , \28695 , \28701 );
or \U$28326 ( \28703 , \28700 , \28318 );
nand \U$28327 ( \28704 , \28702 , \28703 );
and \U$28328 ( \28705 , \28694 , \28704 );
and \U$28329 ( \28706 , \28532 , \28693 );
nor \U$28330 ( \28707 , \28705 , \28706 );
or \U$28331 ( \28708 , \28527 , \28707 );
xnor \U$28332 ( \28709 , \28527 , \28707 );
xor \U$28333 ( \28710 , \28391 , \28450 );
xor \U$28334 ( \28711 , \28710 , \28468 );
xor \U$28335 ( \28712 , \28549 , \28551 );
xor \U$28336 ( \28713 , \28712 , \28684 );
xor \U$28337 ( \28714 , \28711 , \28713 );
and \U$28338 ( \28715 , \7633 , RIae773d8_75);
and \U$28339 ( \28716 , RIae77a68_89, \7631 );
nor \U$28340 ( \28717 , \28715 , \28716 );
and \U$28341 ( \28718 , \28717 , \7206 );
not \U$28342 ( \28719 , \28717 );
and \U$28343 ( \28720 , \28719 , \7205 );
nor \U$28344 ( \28721 , \28718 , \28720 );
and \U$28345 ( \28722 , \8371 , RIae77978_87);
and \U$28346 ( \28723 , RIae77798_83, \8369 );
nor \U$28347 ( \28724 , \28722 , \28723 );
and \U$28348 ( \28725 , \28724 , \8020 );
not \U$28349 ( \28726 , \28724 );
and \U$28350 ( \28727 , \28726 , \8019 );
nor \U$28351 ( \28728 , \28725 , \28727 );
xor \U$28352 ( \28729 , \28721 , \28728 );
and \U$28353 ( \28730 , \8966 , RIae77888_85);
and \U$28354 ( \28731 , RIae76f28_65, \8964 );
nor \U$28355 ( \28732 , \28730 , \28731 );
and \U$28356 ( \28733 , \28732 , \8799 );
not \U$28357 ( \28734 , \28732 );
and \U$28358 ( \28735 , \28734 , \8789 );
nor \U$28359 ( \28736 , \28733 , \28735 );
and \U$28360 ( \28737 , \28729 , \28736 );
and \U$28361 ( \28738 , \28721 , \28728 );
or \U$28362 ( \28739 , \28737 , \28738 );
nand \U$28363 ( \28740 , RIae775b8_79, \6170 );
and \U$28364 ( \28741 , \28740 , \6176 );
not \U$28365 ( \28742 , \28740 );
and \U$28366 ( \28743 , \28742 , \6175 );
nor \U$28367 ( \28744 , \28741 , \28743 );
and \U$28368 ( \28745 , \6941 , RIae774c8_77);
and \U$28369 ( \28746 , RIae77720_82, \6939 );
nor \U$28370 ( \28747 , \28745 , \28746 );
and \U$28371 ( \28748 , \28747 , \6314 );
not \U$28372 ( \28749 , \28747 );
and \U$28373 ( \28750 , \28749 , \6945 );
nor \U$28374 ( \28751 , \28748 , \28750 );
and \U$28375 ( \28752 , \28744 , \28751 );
xnor \U$28376 ( \28753 , \28739 , \28752 );
not \U$28377 ( \28754 , \28753 );
and \U$28378 ( \28755 , \6172 , RIae775b8_79);
and \U$28379 ( \28756 , RIae774c8_77, \6170 );
nor \U$28380 ( \28757 , \28755 , \28756 );
and \U$28381 ( \28758 , \28757 , \6176 );
not \U$28382 ( \28759 , \28757 );
and \U$28383 ( \28760 , \28759 , \6175 );
nor \U$28384 ( \28761 , \28758 , \28760 );
not \U$28385 ( \28762 , \28761 );
and \U$28386 ( \28763 , \28754 , \28762 );
and \U$28387 ( \28764 , \28753 , \28761 );
nor \U$28388 ( \28765 , \28763 , \28764 );
xor \U$28389 ( \28766 , \28619 , \28626 );
xor \U$28390 ( \28767 , \28766 , \28634 );
xor \U$28391 ( \28768 , \28765 , \28767 );
not \U$28392 ( \28769 , \28568 );
not \U$28393 ( \28770 , \28579 );
or \U$28394 ( \28771 , \28769 , \28770 );
or \U$28395 ( \28772 , \28568 , \28579 );
nand \U$28396 ( \28773 , \28771 , \28772 );
not \U$28397 ( \28774 , \28773 );
not \U$28398 ( \28775 , \28561 );
and \U$28399 ( \28776 , \28774 , \28775 );
and \U$28400 ( \28777 , \28773 , \28561 );
nor \U$28401 ( \28778 , \28776 , \28777 );
xor \U$28402 ( \28779 , \28594 , \28601 );
xor \U$28403 ( \28780 , \28779 , \28609 );
xor \U$28404 ( \28781 , \28778 , \28780 );
not \U$28405 ( \28782 , \28652 );
not \U$28406 ( \28783 , \28663 );
or \U$28407 ( \28784 , \28782 , \28783 );
or \U$28408 ( \28785 , \28652 , \28663 );
nand \U$28409 ( \28786 , \28784 , \28785 );
not \U$28410 ( \28787 , \28786 );
not \U$28411 ( \28788 , \28645 );
and \U$28412 ( \28789 , \28787 , \28788 );
and \U$28413 ( \28790 , \28786 , \28645 );
nor \U$28414 ( \28791 , \28789 , \28790 );
xor \U$28415 ( \28792 , \28781 , \28791 );
and \U$28416 ( \28793 , \28768 , \28792 );
and \U$28417 ( \28794 , \28765 , \28767 );
or \U$28418 ( \28795 , \28793 , \28794 );
and \U$28419 ( \28796 , \9760 , RIae76e38_63);
and \U$28420 ( \28797 , RIae76d48_61, \9758 );
nor \U$28421 ( \28798 , \28796 , \28797 );
and \U$28422 ( \28799 , \28798 , \9273 );
not \U$28423 ( \28800 , \28798 );
and \U$28424 ( \28801 , \28800 , \9764 );
nor \U$28425 ( \28802 , \28799 , \28801 );
and \U$28426 ( \28803 , \10548 , RIae76c58_59);
and \U$28427 ( \28804 , RIae77180_70, \10546 );
nor \U$28428 ( \28805 , \28803 , \28804 );
and \U$28429 ( \28806 , \28805 , \10421 );
not \U$28430 ( \28807 , \28805 );
and \U$28431 ( \28808 , \28807 , \10118 );
nor \U$28432 ( \28809 , \28806 , \28808 );
xor \U$28433 ( \28810 , \28802 , \28809 );
and \U$28434 ( \28811 , \11470 , RIae77018_67);
and \U$28435 ( \28812 , RIae771f8_71, \11468 );
nor \U$28436 ( \28813 , \28811 , \28812 );
and \U$28437 ( \28814 , \28813 , \10936 );
not \U$28438 ( \28815 , \28813 );
and \U$28439 ( \28816 , \28815 , \11474 );
nor \U$28440 ( \28817 , \28814 , \28816 );
xor \U$28441 ( \28818 , \28810 , \28817 );
and \U$28442 ( \28819 , \12180 , RIae772e8_73);
and \U$28443 ( \28820 , RIae782d8_107, \12178 );
nor \U$28444 ( \28821 , \28819 , \28820 );
and \U$28445 ( \28822 , \28821 , \12184 );
not \U$28446 ( \28823 , \28821 );
and \U$28447 ( \28824 , \28823 , \11827 );
nor \U$28448 ( \28825 , \28822 , \28824 );
and \U$28449 ( \28826 , \13059 , RIae780f8_103);
and \U$28450 ( \28827 , RIae77f18_99, \13057 );
nor \U$28451 ( \28828 , \28826 , \28827 );
and \U$28452 ( \28829 , \28828 , \13063 );
not \U$28453 ( \28830 , \28828 );
and \U$28454 ( \28831 , \28830 , \12718 );
nor \U$28455 ( \28832 , \28829 , \28831 );
xor \U$28456 ( \28833 , \28825 , \28832 );
and \U$28457 ( \28834 , \14059 , RIae78008_101);
and \U$28458 ( \28835 , RIae781e8_105, \14057 );
nor \U$28459 ( \28836 , \28834 , \28835 );
and \U$28460 ( \28837 , \28836 , \13502 );
not \U$28461 ( \28838 , \28836 );
and \U$28462 ( \28839 , \28838 , \14063 );
nor \U$28463 ( \28840 , \28837 , \28839 );
xor \U$28464 ( \28841 , \28833 , \28840 );
and \U$28465 ( \28842 , \28818 , \28841 );
and \U$28466 ( \28843 , \15726 , RIae78530_112);
and \U$28467 ( \28844 , RIae7aab0_192, RIae77c48_93);
nor \U$28468 ( \28845 , \28843 , \28844 );
and \U$28469 ( \28846 , \28845 , \14959 );
not \U$28470 ( \28847 , \28845 );
and \U$28471 ( \28848 , \28847 , RIae7aa38_191);
nor \U$28472 ( \28849 , \28846 , \28848 );
xor \U$28473 ( \28850 , \28849 , \6175 );
and \U$28474 ( \28851 , \14964 , RIae785a8_113);
and \U$28475 ( \28852 , RIae783c8_109, \14962 );
nor \U$28476 ( \28853 , \28851 , \28852 );
and \U$28477 ( \28854 , \28853 , \14463 );
not \U$28478 ( \28855 , \28853 );
and \U$28479 ( \28856 , \28855 , \14462 );
nor \U$28480 ( \28857 , \28854 , \28856 );
xor \U$28481 ( \28858 , \28850 , \28857 );
xor \U$28482 ( \28859 , \28825 , \28832 );
xor \U$28483 ( \28860 , \28859 , \28840 );
and \U$28484 ( \28861 , \28858 , \28860 );
and \U$28485 ( \28862 , \28818 , \28858 );
or \U$28486 ( \28863 , \28842 , \28861 , \28862 );
and \U$28487 ( \28864 , \9760 , RIae76f28_65);
and \U$28488 ( \28865 , RIae76e38_63, \9758 );
nor \U$28489 ( \28866 , \28864 , \28865 );
and \U$28490 ( \28867 , \28866 , \9273 );
not \U$28491 ( \28868 , \28866 );
and \U$28492 ( \28869 , \28868 , \9764 );
nor \U$28493 ( \28870 , \28867 , \28869 );
and \U$28494 ( \28871 , \8966 , RIae77798_83);
and \U$28495 ( \28872 , RIae77888_85, \8964 );
nor \U$28496 ( \28873 , \28871 , \28872 );
and \U$28497 ( \28874 , \28873 , \8799 );
not \U$28498 ( \28875 , \28873 );
and \U$28499 ( \28876 , \28875 , \8789 );
nor \U$28500 ( \28877 , \28874 , \28876 );
xor \U$28501 ( \28878 , \28870 , \28877 );
and \U$28502 ( \28879 , \10548 , RIae76d48_61);
and \U$28503 ( \28880 , RIae76c58_59, \10546 );
nor \U$28504 ( \28881 , \28879 , \28880 );
and \U$28505 ( \28882 , \28881 , \10421 );
not \U$28506 ( \28883 , \28881 );
and \U$28507 ( \28884 , \28883 , \10118 );
nor \U$28508 ( \28885 , \28882 , \28884 );
and \U$28509 ( \28886 , \28878 , \28885 );
and \U$28510 ( \28887 , \28870 , \28877 );
or \U$28511 ( \28888 , \28886 , \28887 );
and \U$28512 ( \28889 , \14059 , RIae77f18_99);
and \U$28513 ( \28890 , RIae78008_101, \14057 );
nor \U$28514 ( \28891 , \28889 , \28890 );
and \U$28515 ( \28892 , \28891 , \14063 );
not \U$28516 ( \28893 , \28891 );
and \U$28517 ( \28894 , \28893 , \13502 );
nor \U$28518 ( \28895 , \28892 , \28894 );
and \U$28519 ( \28896 , \15726 , RIae783c8_109);
and \U$28520 ( \28897 , RIae7aab0_192, RIae78530_112);
nor \U$28521 ( \28898 , \28896 , \28897 );
and \U$28522 ( \28899 , \28898 , RIae7aa38_191);
not \U$28523 ( \28900 , \28898 );
and \U$28524 ( \28901 , \28900 , \14959 );
nor \U$28525 ( \28902 , \28899 , \28901 );
or \U$28526 ( \28903 , \28895 , \28902 );
not \U$28527 ( \28904 , \28902 );
not \U$28528 ( \28905 , \28895 );
or \U$28529 ( \28906 , \28904 , \28905 );
and \U$28530 ( \28907 , \14964 , RIae781e8_105);
and \U$28531 ( \28908 , RIae785a8_113, \14962 );
nor \U$28532 ( \28909 , \28907 , \28908 );
and \U$28533 ( \28910 , \28909 , \14463 );
not \U$28534 ( \28911 , \28909 );
and \U$28535 ( \28912 , \28911 , \14462 );
nor \U$28536 ( \28913 , \28910 , \28912 );
nand \U$28537 ( \28914 , \28906 , \28913 );
nand \U$28538 ( \28915 , \28903 , \28914 );
xor \U$28539 ( \28916 , \28888 , \28915 );
and \U$28540 ( \28917 , \11470 , RIae77180_70);
and \U$28541 ( \28918 , RIae77018_67, \11468 );
nor \U$28542 ( \28919 , \28917 , \28918 );
and \U$28543 ( \28920 , \28919 , \10936 );
not \U$28544 ( \28921 , \28919 );
and \U$28545 ( \28922 , \28921 , \11474 );
nor \U$28546 ( \28923 , \28920 , \28922 );
and \U$28547 ( \28924 , \12180 , RIae771f8_71);
and \U$28548 ( \28925 , RIae772e8_73, \12178 );
nor \U$28549 ( \28926 , \28924 , \28925 );
and \U$28550 ( \28927 , \28926 , \12184 );
not \U$28551 ( \28928 , \28926 );
and \U$28552 ( \28929 , \28928 , \11827 );
nor \U$28553 ( \28930 , \28927 , \28929 );
xor \U$28554 ( \28931 , \28923 , \28930 );
and \U$28555 ( \28932 , \13059 , RIae782d8_107);
and \U$28556 ( \28933 , RIae780f8_103, \13057 );
nor \U$28557 ( \28934 , \28932 , \28933 );
and \U$28558 ( \28935 , \28934 , \13063 );
not \U$28559 ( \28936 , \28934 );
and \U$28560 ( \28937 , \28936 , \12718 );
nor \U$28561 ( \28938 , \28935 , \28937 );
and \U$28562 ( \28939 , \28931 , \28938 );
and \U$28563 ( \28940 , \28923 , \28930 );
or \U$28564 ( \28941 , \28939 , \28940 );
and \U$28565 ( \28942 , \28916 , \28941 );
and \U$28566 ( \28943 , \28888 , \28915 );
or \U$28567 ( \28944 , \28942 , \28943 );
xor \U$28568 ( \28945 , \28863 , \28944 );
and \U$28569 ( \28946 , \7633 , RIae77720_82);
and \U$28570 ( \28947 , RIae773d8_75, \7631 );
nor \U$28571 ( \28948 , \28946 , \28947 );
and \U$28572 ( \28949 , \28948 , \7206 );
not \U$28573 ( \28950 , \28948 );
and \U$28574 ( \28951 , \28950 , \7205 );
nor \U$28575 ( \28952 , \28949 , \28951 );
and \U$28576 ( \28953 , \6941 , RIae775b8_79);
and \U$28577 ( \28954 , RIae774c8_77, \6939 );
nor \U$28578 ( \28955 , \28953 , \28954 );
and \U$28579 ( \28956 , \28955 , \6314 );
not \U$28580 ( \28957 , \28955 );
and \U$28581 ( \28958 , \28957 , \6945 );
nor \U$28582 ( \28959 , \28956 , \28958 );
xor \U$28583 ( \28960 , \28952 , \28959 );
and \U$28584 ( \28961 , \8371 , RIae77a68_89);
and \U$28585 ( \28962 , RIae77978_87, \8369 );
nor \U$28586 ( \28963 , \28961 , \28962 );
and \U$28587 ( \28964 , \28963 , \8020 );
not \U$28588 ( \28965 , \28963 );
and \U$28589 ( \28966 , \28965 , \8019 );
nor \U$28590 ( \28967 , \28964 , \28966 );
and \U$28591 ( \28968 , \28960 , \28967 );
and \U$28592 ( \28969 , \28952 , \28959 );
or \U$28593 ( \28970 , \28968 , \28969 );
xor \U$28594 ( \28971 , \28744 , \28751 );
xor \U$28595 ( \28972 , \28970 , \28971 );
xor \U$28596 ( \28973 , \28721 , \28728 );
xor \U$28597 ( \28974 , \28973 , \28736 );
and \U$28598 ( \28975 , \28972 , \28974 );
and \U$28599 ( \28976 , \28970 , \28971 );
or \U$28600 ( \28977 , \28975 , \28976 );
and \U$28601 ( \28978 , \28945 , \28977 );
and \U$28602 ( \28979 , \28863 , \28944 );
nor \U$28603 ( \28980 , \28978 , \28979 );
or \U$28604 ( \28981 , \28795 , \28980 );
not \U$28605 ( \28982 , \28980 );
not \U$28606 ( \28983 , \28795 );
or \U$28607 ( \28984 , \28982 , \28983 );
xor \U$28608 ( \28985 , \28554 , \28581 );
xor \U$28609 ( \28986 , \28985 , \28584 );
xor \U$28610 ( \28987 , \28612 , \28637 );
xor \U$28611 ( \28988 , \28987 , \28665 );
xor \U$28612 ( \28989 , \28370 , \28377 );
xor \U$28613 ( \28990 , \28989 , \28385 );
xor \U$28614 ( \28991 , \28671 , \28676 );
xor \U$28615 ( \28992 , \28990 , \28991 );
xor \U$28616 ( \28993 , \28988 , \28992 );
xor \U$28617 ( \28994 , \28986 , \28993 );
nand \U$28618 ( \28995 , \28984 , \28994 );
nand \U$28619 ( \28996 , \28981 , \28995 );
xor \U$28620 ( \28997 , \28802 , \28809 );
and \U$28621 ( \28998 , \28997 , \28817 );
and \U$28622 ( \28999 , \28802 , \28809 );
or \U$28623 ( \29000 , \28998 , \28999 );
xor \U$28624 ( \29001 , \28849 , \6175 );
and \U$28625 ( \29002 , \29001 , \28857 );
and \U$28626 ( \29003 , \28849 , \6175 );
or \U$28627 ( \29004 , \29002 , \29003 );
xor \U$28628 ( \29005 , \29000 , \29004 );
xor \U$28629 ( \29006 , \28825 , \28832 );
and \U$28630 ( \29007 , \29006 , \28840 );
and \U$28631 ( \29008 , \28825 , \28832 );
or \U$28632 ( \29009 , \29007 , \29008 );
and \U$28633 ( \29010 , \29005 , \29009 );
and \U$28634 ( \29011 , \29000 , \29004 );
or \U$28635 ( \29012 , \29010 , \29011 );
not \U$28636 ( \29013 , \28761 );
not \U$28637 ( \29014 , \28752 );
or \U$28638 ( \29015 , \29013 , \29014 );
or \U$28639 ( \29016 , \28752 , \28761 );
nand \U$28640 ( \29017 , \29016 , \28739 );
nand \U$28641 ( \29018 , \29015 , \29017 );
xor \U$28642 ( \29019 , \29012 , \29018 );
xor \U$28643 ( \29020 , \28778 , \28780 );
and \U$28644 ( \29021 , \29020 , \28791 );
and \U$28645 ( \29022 , \28778 , \28780 );
nor \U$28646 ( \29023 , \29021 , \29022 );
and \U$28647 ( \29024 , \29019 , \29023 );
and \U$28648 ( \29025 , \29012 , \29018 );
or \U$28649 ( \29026 , \29024 , \29025 );
xor \U$28650 ( \29027 , \28414 , \28421 );
xor \U$28651 ( \29028 , \29027 , \28447 );
xor \U$28652 ( \29029 , \29026 , \29028 );
xor \U$28653 ( \29030 , \28554 , \28581 );
xor \U$28654 ( \29031 , \29030 , \28584 );
and \U$28655 ( \29032 , \28988 , \29031 );
xor \U$28656 ( \29033 , \28554 , \28581 );
xor \U$28657 ( \29034 , \29033 , \28584 );
and \U$28658 ( \29035 , \28992 , \29034 );
and \U$28659 ( \29036 , \28988 , \28992 );
or \U$28660 ( \29037 , \29032 , \29035 , \29036 );
xor \U$28661 ( \29038 , \29029 , \29037 );
and \U$28662 ( \29039 , \28996 , \29038 );
xor \U$28663 ( \29040 , \28539 , \28541 );
xor \U$28664 ( \29041 , \29040 , \28546 );
xor \U$28665 ( \29042 , \28344 , \28362 );
xor \U$28666 ( \29043 , \29042 , \28388 );
xor \U$28667 ( \29044 , \28587 , \28668 );
xor \U$28668 ( \29045 , \29044 , \28681 );
xor \U$28669 ( \29046 , \29043 , \29045 );
xor \U$28670 ( \29047 , \29041 , \29046 );
xor \U$28671 ( \29048 , \29026 , \29028 );
xor \U$28672 ( \29049 , \29048 , \29037 );
and \U$28673 ( \29050 , \29047 , \29049 );
and \U$28674 ( \29051 , \28996 , \29047 );
or \U$28675 ( \29052 , \29039 , \29050 , \29051 );
xor \U$28676 ( \29053 , \28714 , \29052 );
xor \U$28677 ( \29054 , \28539 , \28541 );
xor \U$28678 ( \29055 , \29054 , \28546 );
and \U$28679 ( \29056 , \29043 , \29055 );
xor \U$28680 ( \29057 , \28539 , \28541 );
xor \U$28681 ( \29058 , \29057 , \28546 );
and \U$28682 ( \29059 , \29045 , \29058 );
and \U$28683 ( \29060 , \29043 , \29045 );
or \U$28684 ( \29061 , \29056 , \29059 , \29060 );
xor \U$28685 ( \29062 , \28480 , \28482 );
xor \U$28686 ( \29063 , \29062 , \28487 );
xor \U$28687 ( \29064 , \29061 , \29063 );
xor \U$28688 ( \29065 , \29026 , \29028 );
and \U$28689 ( \29066 , \29065 , \29037 );
and \U$28690 ( \29067 , \29026 , \29028 );
or \U$28691 ( \29068 , \29066 , \29067 );
xor \U$28692 ( \29069 , \29064 , \29068 );
and \U$28693 ( \29070 , \29053 , \29069 );
and \U$28694 ( \29071 , \28714 , \29052 );
nor \U$28695 ( \29072 , \29070 , \29071 );
and \U$28696 ( \29073 , \28711 , \28713 );
xor \U$28697 ( \29074 , \29061 , \29063 );
and \U$28698 ( \29075 , \29074 , \29068 );
and \U$28699 ( \29076 , \29061 , \29063 );
or \U$28700 ( \29077 , \29075 , \29076 );
xnor \U$28701 ( \29078 , \29073 , \29077 );
not \U$28702 ( \29079 , \29078 );
xor \U$28703 ( \29080 , \28537 , \28687 );
xor \U$28704 ( \29081 , \29080 , \28690 );
not \U$28705 ( \29082 , \29081 );
and \U$28706 ( \29083 , \29079 , \29082 );
and \U$28707 ( \29084 , \29078 , \29081 );
nor \U$28708 ( \29085 , \29083 , \29084 );
or \U$28709 ( \29086 , \29072 , \29085 );
xnor \U$28710 ( \29087 , \29085 , \29072 );
xor \U$28711 ( \29088 , \29026 , \29028 );
xor \U$28712 ( \29089 , \29088 , \29037 );
xor \U$28713 ( \29090 , \28996 , \29047 );
xor \U$28714 ( \29091 , \29089 , \29090 );
not \U$28715 ( \29092 , \29091 );
xor \U$28716 ( \29093 , \29012 , \29018 );
xor \U$28717 ( \29094 , \29093 , \29023 );
not \U$28718 ( \29095 , \29094 );
xor \U$28719 ( \29096 , \28765 , \28767 );
xor \U$28720 ( \29097 , \29096 , \28792 );
not \U$28721 ( \29098 , \29097 );
xor \U$28722 ( \29099 , \28863 , \28944 );
xor \U$28723 ( \29100 , \29099 , \28977 );
nand \U$28724 ( \29101 , \29098 , \29100 );
nand \U$28725 ( \29102 , \29095 , \29101 );
and \U$28726 ( \29103 , \15726 , RIae785a8_113);
and \U$28727 ( \29104 , RIae7aab0_192, RIae783c8_109);
nor \U$28728 ( \29105 , \29103 , \29104 );
and \U$28729 ( \29106 , \29105 , \14959 );
not \U$28730 ( \29107 , \29105 );
and \U$28731 ( \29108 , \29107 , RIae7aa38_191);
nor \U$28732 ( \29109 , \29106 , \29108 );
xor \U$28733 ( \29110 , \29109 , \6945 );
and \U$28734 ( \29111 , \14964 , RIae78008_101);
and \U$28735 ( \29112 , RIae781e8_105, \14962 );
nor \U$28736 ( \29113 , \29111 , \29112 );
and \U$28737 ( \29114 , \29113 , \14463 );
not \U$28738 ( \29115 , \29113 );
and \U$28739 ( \29116 , \29115 , \14462 );
nor \U$28740 ( \29117 , \29114 , \29116 );
and \U$28741 ( \29118 , \29110 , \29117 );
and \U$28742 ( \29119 , \29109 , \6945 );
or \U$28743 ( \29120 , \29118 , \29119 );
and \U$28744 ( \29121 , \12180 , RIae77018_67);
and \U$28745 ( \29122 , RIae771f8_71, \12178 );
nor \U$28746 ( \29123 , \29121 , \29122 );
and \U$28747 ( \29124 , \29123 , \12184 );
not \U$28748 ( \29125 , \29123 );
and \U$28749 ( \29126 , \29125 , \11827 );
nor \U$28750 ( \29127 , \29124 , \29126 );
and \U$28751 ( \29128 , \13059 , RIae772e8_73);
and \U$28752 ( \29129 , RIae782d8_107, \13057 );
nor \U$28753 ( \29130 , \29128 , \29129 );
and \U$28754 ( \29131 , \29130 , \13063 );
not \U$28755 ( \29132 , \29130 );
and \U$28756 ( \29133 , \29132 , \12718 );
nor \U$28757 ( \29134 , \29131 , \29133 );
xor \U$28758 ( \29135 , \29127 , \29134 );
and \U$28759 ( \29136 , \14059 , RIae780f8_103);
and \U$28760 ( \29137 , RIae77f18_99, \14057 );
nor \U$28761 ( \29138 , \29136 , \29137 );
and \U$28762 ( \29139 , \29138 , \13502 );
not \U$28763 ( \29140 , \29138 );
and \U$28764 ( \29141 , \29140 , \14063 );
nor \U$28765 ( \29142 , \29139 , \29141 );
and \U$28766 ( \29143 , \29135 , \29142 );
and \U$28767 ( \29144 , \29127 , \29134 );
or \U$28768 ( \29145 , \29143 , \29144 );
xor \U$28769 ( \29146 , \29120 , \29145 );
and \U$28770 ( \29147 , \9760 , RIae77888_85);
and \U$28771 ( \29148 , RIae76f28_65, \9758 );
nor \U$28772 ( \29149 , \29147 , \29148 );
and \U$28773 ( \29150 , \29149 , \9273 );
not \U$28774 ( \29151 , \29149 );
and \U$28775 ( \29152 , \29151 , \9764 );
nor \U$28776 ( \29153 , \29150 , \29152 );
and \U$28777 ( \29154 , \10548 , RIae76e38_63);
and \U$28778 ( \29155 , RIae76d48_61, \10546 );
nor \U$28779 ( \29156 , \29154 , \29155 );
and \U$28780 ( \29157 , \29156 , \10421 );
not \U$28781 ( \29158 , \29156 );
and \U$28782 ( \29159 , \29158 , \10118 );
nor \U$28783 ( \29160 , \29157 , \29159 );
xor \U$28784 ( \29161 , \29153 , \29160 );
and \U$28785 ( \29162 , \11470 , RIae76c58_59);
and \U$28786 ( \29163 , RIae77180_70, \11468 );
nor \U$28787 ( \29164 , \29162 , \29163 );
and \U$28788 ( \29165 , \29164 , \10936 );
not \U$28789 ( \29166 , \29164 );
and \U$28790 ( \29167 , \29166 , \11474 );
nor \U$28791 ( \29168 , \29165 , \29167 );
and \U$28792 ( \29169 , \29161 , \29168 );
and \U$28793 ( \29170 , \29153 , \29160 );
or \U$28794 ( \29171 , \29169 , \29170 );
and \U$28795 ( \29172 , \29146 , \29171 );
and \U$28796 ( \29173 , \29120 , \29145 );
nor \U$28797 ( \29174 , \29172 , \29173 );
not \U$28798 ( \29175 , \29174 );
not \U$28799 ( \29176 , \28902 );
not \U$28800 ( \29177 , \28913 );
or \U$28801 ( \29178 , \29176 , \29177 );
or \U$28802 ( \29179 , \28913 , \28902 );
nand \U$28803 ( \29180 , \29178 , \29179 );
not \U$28804 ( \29181 , \29180 );
not \U$28805 ( \29182 , \28895 );
and \U$28806 ( \29183 , \29181 , \29182 );
and \U$28807 ( \29184 , \29180 , \28895 );
nor \U$28808 ( \29185 , \29183 , \29184 );
not \U$28809 ( \29186 , \29185 );
xor \U$28810 ( \29187 , \28923 , \28930 );
xor \U$28811 ( \29188 , \29187 , \28938 );
nand \U$28812 ( \29189 , \29186 , \29188 );
not \U$28813 ( \29190 , \29189 );
and \U$28814 ( \29191 , \29175 , \29190 );
and \U$28815 ( \29192 , \29174 , \29189 );
xor \U$28816 ( \29193 , \28870 , \28877 );
xor \U$28817 ( \29194 , \29193 , \28885 );
xor \U$28818 ( \29195 , \28952 , \28959 );
xor \U$28819 ( \29196 , \29195 , \28967 );
and \U$28820 ( \29197 , \29194 , \29196 );
not \U$28821 ( \29198 , \29196 );
not \U$28822 ( \29199 , \29194 );
and \U$28823 ( \29200 , \29198 , \29199 );
and \U$28824 ( \29201 , \8371 , RIae773d8_75);
and \U$28825 ( \29202 , RIae77a68_89, \8369 );
nor \U$28826 ( \29203 , \29201 , \29202 );
and \U$28827 ( \29204 , \29203 , \8020 );
not \U$28828 ( \29205 , \29203 );
and \U$28829 ( \29206 , \29205 , \8019 );
nor \U$28830 ( \29207 , \29204 , \29206 );
and \U$28831 ( \29208 , \8966 , RIae77978_87);
and \U$28832 ( \29209 , RIae77798_83, \8964 );
nor \U$28833 ( \29210 , \29208 , \29209 );
and \U$28834 ( \29211 , \29210 , \8799 );
not \U$28835 ( \29212 , \29210 );
and \U$28836 ( \29213 , \29212 , \8789 );
nor \U$28837 ( \29214 , \29211 , \29213 );
xor \U$28838 ( \29215 , \29207 , \29214 );
and \U$28839 ( \29216 , \7633 , RIae774c8_77);
and \U$28840 ( \29217 , RIae77720_82, \7631 );
nor \U$28841 ( \29218 , \29216 , \29217 );
and \U$28842 ( \29219 , \29218 , \7206 );
not \U$28843 ( \29220 , \29218 );
and \U$28844 ( \29221 , \29220 , \7205 );
nor \U$28845 ( \29222 , \29219 , \29221 );
and \U$28846 ( \29223 , \29215 , \29222 );
and \U$28847 ( \29224 , \29207 , \29214 );
nor \U$28848 ( \29225 , \29223 , \29224 );
nor \U$28849 ( \29226 , \29200 , \29225 );
nor \U$28850 ( \29227 , \29197 , \29226 );
nor \U$28851 ( \29228 , \29192 , \29227 );
nor \U$28852 ( \29229 , \29191 , \29228 );
xor \U$28853 ( \29230 , \29000 , \29004 );
xor \U$28854 ( \29231 , \29230 , \29009 );
not \U$28855 ( \29232 , \29231 );
or \U$28856 ( \29233 , \29229 , \29232 );
not \U$28857 ( \29234 , \29232 );
not \U$28858 ( \29235 , \29229 );
or \U$28859 ( \29236 , \29234 , \29235 );
xor \U$28860 ( \29237 , \28888 , \28915 );
xor \U$28861 ( \29238 , \29237 , \28941 );
xor \U$28862 ( \29239 , \28970 , \28971 );
xor \U$28863 ( \29240 , \29239 , \28974 );
and \U$28864 ( \29241 , \29238 , \29240 );
xor \U$28865 ( \29242 , \28825 , \28832 );
xor \U$28866 ( \29243 , \29242 , \28840 );
xor \U$28867 ( \29244 , \28818 , \28858 );
xor \U$28868 ( \29245 , \29243 , \29244 );
xor \U$28869 ( \29246 , \28970 , \28971 );
xor \U$28870 ( \29247 , \29246 , \28974 );
and \U$28871 ( \29248 , \29245 , \29247 );
and \U$28872 ( \29249 , \29238 , \29245 );
or \U$28873 ( \29250 , \29241 , \29248 , \29249 );
nand \U$28874 ( \29251 , \29236 , \29250 );
nand \U$28875 ( \29252 , \29233 , \29251 );
and \U$28876 ( \29253 , \29102 , \29252 );
not \U$28877 ( \29254 , \29101 );
and \U$28878 ( \29255 , \29094 , \29254 );
nor \U$28879 ( \29256 , \29253 , \29255 );
not \U$28880 ( \29257 , \29256 );
and \U$28881 ( \29258 , \29092 , \29257 );
and \U$28882 ( \29259 , \29091 , \29256 );
nor \U$28883 ( \29260 , \29258 , \29259 );
xnor \U$28884 ( \29261 , \28980 , \28795 );
not \U$28885 ( \29262 , \29261 );
not \U$28886 ( \29263 , \28994 );
and \U$28887 ( \29264 , \29262 , \29263 );
and \U$28888 ( \29265 , \29261 , \28994 );
nor \U$28889 ( \29266 , \29264 , \29265 );
not \U$28890 ( \29267 , \29266 );
not \U$28891 ( \29268 , \29094 );
not \U$28892 ( \29269 , \29252 );
not \U$28893 ( \29270 , \29101 );
and \U$28894 ( \29271 , \29269 , \29270 );
and \U$28895 ( \29272 , \29252 , \29101 );
nor \U$28896 ( \29273 , \29271 , \29272 );
not \U$28897 ( \29274 , \29273 );
or \U$28898 ( \29275 , \29268 , \29274 );
or \U$28899 ( \29276 , \29273 , \29094 );
nand \U$28900 ( \29277 , \29275 , \29276 );
nand \U$28901 ( \29278 , \29267 , \29277 );
or \U$28902 ( \29279 , \29260 , \29278 );
xnor \U$28903 ( \29280 , \29278 , \29260 );
not \U$28904 ( \29281 , \29266 );
not \U$28905 ( \29282 , \29277 );
or \U$28906 ( \29283 , \29281 , \29282 );
or \U$28907 ( \29284 , \29277 , \29266 );
nand \U$28908 ( \29285 , \29283 , \29284 );
not \U$28909 ( \29286 , \29250 );
not \U$28910 ( \29287 , \29229 );
and \U$28911 ( \29288 , \29286 , \29287 );
and \U$28912 ( \29289 , \29250 , \29229 );
nor \U$28913 ( \29290 , \29288 , \29289 );
not \U$28914 ( \29291 , \29290 );
not \U$28915 ( \29292 , \29231 );
and \U$28916 ( \29293 , \29291 , \29292 );
and \U$28917 ( \29294 , \29290 , \29231 );
nor \U$28918 ( \29295 , \29293 , \29294 );
not \U$28919 ( \29296 , \29100 );
not \U$28920 ( \29297 , \29097 );
and \U$28921 ( \29298 , \29296 , \29297 );
and \U$28922 ( \29299 , \29100 , \29097 );
nor \U$28923 ( \29300 , \29298 , \29299 );
or \U$28924 ( \29301 , \29295 , \29300 );
not \U$28925 ( \29302 , \29300 );
not \U$28926 ( \29303 , \29295 );
or \U$28927 ( \29304 , \29302 , \29303 );
xor \U$28928 ( \29305 , \29120 , \29145 );
xor \U$28929 ( \29306 , \29305 , \29171 );
not \U$28930 ( \29307 , \29188 );
not \U$28931 ( \29308 , \29185 );
or \U$28932 ( \29309 , \29307 , \29308 );
or \U$28933 ( \29310 , \29185 , \29188 );
nand \U$28934 ( \29311 , \29309 , \29310 );
xor \U$28935 ( \29312 , \29306 , \29311 );
not \U$28936 ( \29313 , \29225 );
not \U$28937 ( \29314 , \29194 );
or \U$28938 ( \29315 , \29313 , \29314 );
or \U$28939 ( \29316 , \29194 , \29225 );
nand \U$28940 ( \29317 , \29315 , \29316 );
xor \U$28941 ( \29318 , \29196 , \29317 );
and \U$28942 ( \29319 , \29312 , \29318 );
and \U$28943 ( \29320 , \29306 , \29311 );
or \U$28944 ( \29321 , \29319 , \29320 );
and \U$28945 ( \29322 , \10548 , RIae76f28_65);
and \U$28946 ( \29323 , RIae76e38_63, \10546 );
nor \U$28947 ( \29324 , \29322 , \29323 );
and \U$28948 ( \29325 , \29324 , \10421 );
not \U$28949 ( \29326 , \29324 );
and \U$28950 ( \29327 , \29326 , \10118 );
nor \U$28951 ( \29328 , \29325 , \29327 );
and \U$28952 ( \29329 , \8966 , RIae77a68_89);
and \U$28953 ( \29330 , RIae77978_87, \8964 );
nor \U$28954 ( \29331 , \29329 , \29330 );
and \U$28955 ( \29332 , \29331 , \8799 );
not \U$28956 ( \29333 , \29331 );
and \U$28957 ( \29334 , \29333 , \8789 );
nor \U$28958 ( \29335 , \29332 , \29334 );
xor \U$28959 ( \29336 , \29328 , \29335 );
and \U$28960 ( \29337 , \9760 , RIae77798_83);
and \U$28961 ( \29338 , RIae77888_85, \9758 );
nor \U$28962 ( \29339 , \29337 , \29338 );
and \U$28963 ( \29340 , \29339 , \9273 );
not \U$28964 ( \29341 , \29339 );
and \U$28965 ( \29342 , \29341 , \9272 );
nor \U$28966 ( \29343 , \29340 , \29342 );
and \U$28967 ( \29344 , \29336 , \29343 );
and \U$28968 ( \29345 , \29328 , \29335 );
or \U$28969 ( \29346 , \29344 , \29345 );
and \U$28970 ( \29347 , \14059 , RIae782d8_107);
and \U$28971 ( \29348 , RIae780f8_103, \14057 );
nor \U$28972 ( \29349 , \29347 , \29348 );
and \U$28973 ( \29350 , \29349 , \13502 );
not \U$28974 ( \29351 , \29349 );
and \U$28975 ( \29352 , \29351 , \14063 );
nor \U$28976 ( \29353 , \29350 , \29352 );
and \U$28977 ( \29354 , \15726 , RIae781e8_105);
and \U$28978 ( \29355 , RIae7aab0_192, RIae785a8_113);
nor \U$28979 ( \29356 , \29354 , \29355 );
and \U$28980 ( \29357 , \29356 , \14959 );
not \U$28981 ( \29358 , \29356 );
and \U$28982 ( \29359 , \29358 , RIae7aa38_191);
nor \U$28983 ( \29360 , \29357 , \29359 );
xor \U$28984 ( \29361 , \29353 , \29360 );
and \U$28985 ( \29362 , \14964 , RIae77f18_99);
and \U$28986 ( \29363 , RIae78008_101, \14962 );
nor \U$28987 ( \29364 , \29362 , \29363 );
and \U$28988 ( \29365 , \29364 , \14463 );
not \U$28989 ( \29366 , \29364 );
and \U$28990 ( \29367 , \29366 , \14462 );
nor \U$28991 ( \29368 , \29365 , \29367 );
and \U$28992 ( \29369 , \29361 , \29368 );
and \U$28993 ( \29370 , \29353 , \29360 );
or \U$28994 ( \29371 , \29369 , \29370 );
xor \U$28995 ( \29372 , \29346 , \29371 );
and \U$28996 ( \29373 , \11470 , RIae76d48_61);
and \U$28997 ( \29374 , RIae76c58_59, \11468 );
nor \U$28998 ( \29375 , \29373 , \29374 );
and \U$28999 ( \29376 , \29375 , \10936 );
not \U$29000 ( \29377 , \29375 );
and \U$29001 ( \29378 , \29377 , \11474 );
nor \U$29002 ( \29379 , \29376 , \29378 );
and \U$29003 ( \29380 , \12180 , RIae77180_70);
and \U$29004 ( \29381 , RIae77018_67, \12178 );
nor \U$29005 ( \29382 , \29380 , \29381 );
and \U$29006 ( \29383 , \29382 , \12184 );
not \U$29007 ( \29384 , \29382 );
and \U$29008 ( \29385 , \29384 , \11827 );
nor \U$29009 ( \29386 , \29383 , \29385 );
xor \U$29010 ( \29387 , \29379 , \29386 );
and \U$29011 ( \29388 , \13059 , RIae771f8_71);
and \U$29012 ( \29389 , RIae772e8_73, \13057 );
nor \U$29013 ( \29390 , \29388 , \29389 );
and \U$29014 ( \29391 , \29390 , \13063 );
not \U$29015 ( \29392 , \29390 );
and \U$29016 ( \29393 , \29392 , \12718 );
nor \U$29017 ( \29394 , \29391 , \29393 );
and \U$29018 ( \29395 , \29387 , \29394 );
and \U$29019 ( \29396 , \29379 , \29386 );
or \U$29020 ( \29397 , \29395 , \29396 );
and \U$29021 ( \29398 , \29372 , \29397 );
and \U$29022 ( \29399 , \29346 , \29371 );
or \U$29023 ( \29400 , \29398 , \29399 );
xor \U$29024 ( \29401 , \29127 , \29134 );
xor \U$29025 ( \29402 , \29401 , \29142 );
xor \U$29026 ( \29403 , \29109 , \6945 );
xor \U$29027 ( \29404 , \29403 , \29117 );
and \U$29028 ( \29405 , \29402 , \29404 );
xor \U$29029 ( \29406 , \29400 , \29405 );
nand \U$29030 ( \29407 , RIae775b8_79, \6939 );
and \U$29031 ( \29408 , \29407 , \6314 );
not \U$29032 ( \29409 , \29407 );
and \U$29033 ( \29410 , \29409 , \6945 );
nor \U$29034 ( \29411 , \29408 , \29410 );
xor \U$29035 ( \29412 , \29153 , \29160 );
xor \U$29036 ( \29413 , \29412 , \29168 );
and \U$29037 ( \29414 , \29411 , \29413 );
xor \U$29038 ( \29415 , \29207 , \29214 );
xor \U$29039 ( \29416 , \29415 , \29222 );
xor \U$29040 ( \29417 , \29153 , \29160 );
xor \U$29041 ( \29418 , \29417 , \29168 );
and \U$29042 ( \29419 , \29416 , \29418 );
and \U$29043 ( \29420 , \29411 , \29416 );
or \U$29044 ( \29421 , \29414 , \29419 , \29420 );
and \U$29045 ( \29422 , \29406 , \29421 );
and \U$29046 ( \29423 , \29400 , \29405 );
or \U$29047 ( \29424 , \29422 , \29423 );
xor \U$29048 ( \29425 , \29321 , \29424 );
xor \U$29049 ( \29426 , \28970 , \28971 );
xor \U$29050 ( \29427 , \29426 , \28974 );
xor \U$29051 ( \29428 , \29238 , \29245 );
xor \U$29052 ( \29429 , \29427 , \29428 );
and \U$29053 ( \29430 , \29425 , \29429 );
and \U$29054 ( \29431 , \29321 , \29424 );
or \U$29055 ( \29432 , \29430 , \29431 );
nand \U$29056 ( \29433 , \29304 , \29432 );
nand \U$29057 ( \29434 , \29301 , \29433 );
and \U$29058 ( \29435 , \29285 , \29434 );
xor \U$29059 ( \29436 , \29434 , \29285 );
not \U$29060 ( \29437 , \29432 );
not \U$29061 ( \29438 , \29295 );
or \U$29062 ( \29439 , \29437 , \29438 );
or \U$29063 ( \29440 , \29295 , \29432 );
nand \U$29064 ( \29441 , \29439 , \29440 );
not \U$29065 ( \29442 , \29441 );
not \U$29066 ( \29443 , \29300 );
and \U$29067 ( \29444 , \29442 , \29443 );
and \U$29068 ( \29445 , \29441 , \29300 );
nor \U$29069 ( \29446 , \29444 , \29445 );
xor \U$29070 ( \29447 , \29321 , \29424 );
xor \U$29071 ( \29448 , \29447 , \29429 );
xor \U$29072 ( \29449 , \29402 , \29404 );
xor \U$29073 ( \29450 , \29346 , \29371 );
xor \U$29074 ( \29451 , \29450 , \29397 );
and \U$29075 ( \29452 , \29449 , \29451 );
xor \U$29076 ( \29453 , \29153 , \29160 );
xor \U$29077 ( \29454 , \29453 , \29168 );
xor \U$29078 ( \29455 , \29411 , \29416 );
xor \U$29079 ( \29456 , \29454 , \29455 );
xor \U$29080 ( \29457 , \29346 , \29371 );
xor \U$29081 ( \29458 , \29457 , \29397 );
and \U$29082 ( \29459 , \29456 , \29458 );
and \U$29083 ( \29460 , \29449 , \29456 );
or \U$29084 ( \29461 , \29452 , \29459 , \29460 );
and \U$29085 ( \29462 , \12180 , RIae76c58_59);
and \U$29086 ( \29463 , RIae77180_70, \12178 );
nor \U$29087 ( \29464 , \29462 , \29463 );
and \U$29088 ( \29465 , \29464 , \12184 );
not \U$29089 ( \29466 , \29464 );
and \U$29090 ( \29467 , \29466 , \11827 );
nor \U$29091 ( \29468 , \29465 , \29467 );
and \U$29092 ( \29469 , \13059 , RIae77018_67);
and \U$29093 ( \29470 , RIae771f8_71, \13057 );
nor \U$29094 ( \29471 , \29469 , \29470 );
and \U$29095 ( \29472 , \29471 , \13063 );
not \U$29096 ( \29473 , \29471 );
and \U$29097 ( \29474 , \29473 , \12718 );
nor \U$29098 ( \29475 , \29472 , \29474 );
xor \U$29099 ( \29476 , \29468 , \29475 );
and \U$29100 ( \29477 , \14059 , RIae772e8_73);
and \U$29101 ( \29478 , RIae782d8_107, \14057 );
nor \U$29102 ( \29479 , \29477 , \29478 );
and \U$29103 ( \29480 , \29479 , \13502 );
not \U$29104 ( \29481 , \29479 );
and \U$29105 ( \29482 , \29481 , \14063 );
nor \U$29106 ( \29483 , \29480 , \29482 );
and \U$29107 ( \29484 , \29476 , \29483 );
and \U$29108 ( \29485 , \29468 , \29475 );
or \U$29109 ( \29486 , \29484 , \29485 );
and \U$29110 ( \29487 , \15726 , RIae78008_101);
and \U$29111 ( \29488 , RIae7aab0_192, RIae781e8_105);
nor \U$29112 ( \29489 , \29487 , \29488 );
and \U$29113 ( \29490 , \29489 , \14959 );
not \U$29114 ( \29491 , \29489 );
and \U$29115 ( \29492 , \29491 , RIae7aa38_191);
nor \U$29116 ( \29493 , \29490 , \29492 );
xor \U$29117 ( \29494 , \29493 , \7205 );
and \U$29118 ( \29495 , \14964 , RIae780f8_103);
and \U$29119 ( \29496 , RIae77f18_99, \14962 );
nor \U$29120 ( \29497 , \29495 , \29496 );
and \U$29121 ( \29498 , \29497 , \14463 );
not \U$29122 ( \29499 , \29497 );
and \U$29123 ( \29500 , \29499 , \14462 );
nor \U$29124 ( \29501 , \29498 , \29500 );
and \U$29125 ( \29502 , \29494 , \29501 );
and \U$29126 ( \29503 , \29493 , \7205 );
or \U$29127 ( \29504 , \29502 , \29503 );
xor \U$29128 ( \29505 , \29486 , \29504 );
and \U$29129 ( \29506 , \11470 , RIae76e38_63);
and \U$29130 ( \29507 , RIae76d48_61, \11468 );
nor \U$29131 ( \29508 , \29506 , \29507 );
and \U$29132 ( \29509 , \29508 , \10936 );
not \U$29133 ( \29510 , \29508 );
and \U$29134 ( \29511 , \29510 , \11474 );
nor \U$29135 ( \29512 , \29509 , \29511 );
and \U$29136 ( \29513 , \9760 , RIae77978_87);
and \U$29137 ( \29514 , RIae77798_83, \9758 );
nor \U$29138 ( \29515 , \29513 , \29514 );
and \U$29139 ( \29516 , \29515 , \9273 );
not \U$29140 ( \29517 , \29515 );
and \U$29141 ( \29518 , \29517 , \9764 );
nor \U$29142 ( \29519 , \29516 , \29518 );
xor \U$29143 ( \29520 , \29512 , \29519 );
and \U$29144 ( \29521 , \10548 , RIae77888_85);
and \U$29145 ( \29522 , RIae76f28_65, \10546 );
nor \U$29146 ( \29523 , \29521 , \29522 );
and \U$29147 ( \29524 , \29523 , \10421 );
not \U$29148 ( \29525 , \29523 );
and \U$29149 ( \29526 , \29525 , \10118 );
nor \U$29150 ( \29527 , \29524 , \29526 );
and \U$29151 ( \29528 , \29520 , \29527 );
and \U$29152 ( \29529 , \29512 , \29519 );
or \U$29153 ( \29530 , \29528 , \29529 );
and \U$29154 ( \29531 , \29505 , \29530 );
and \U$29155 ( \29532 , \29486 , \29504 );
or \U$29156 ( \29533 , \29531 , \29532 );
and \U$29157 ( \29534 , \8371 , RIae77720_82);
and \U$29158 ( \29535 , RIae773d8_75, \8369 );
nor \U$29159 ( \29536 , \29534 , \29535 );
and \U$29160 ( \29537 , \29536 , \8020 );
not \U$29161 ( \29538 , \29536 );
and \U$29162 ( \29539 , \29538 , \8019 );
nor \U$29163 ( \29540 , \29537 , \29539 );
and \U$29164 ( \29541 , \7633 , RIae775b8_79);
and \U$29165 ( \29542 , RIae774c8_77, \7631 );
nor \U$29166 ( \29543 , \29541 , \29542 );
and \U$29167 ( \29544 , \29543 , \7206 );
not \U$29168 ( \29545 , \29543 );
and \U$29169 ( \29546 , \29545 , \7205 );
nor \U$29170 ( \29547 , \29544 , \29546 );
xor \U$29171 ( \29548 , \29540 , \29547 );
and \U$29172 ( \29549 , \8371 , RIae774c8_77);
and \U$29173 ( \29550 , RIae77720_82, \8369 );
nor \U$29174 ( \29551 , \29549 , \29550 );
and \U$29175 ( \29552 , \29551 , \8020 );
not \U$29176 ( \29553 , \29551 );
and \U$29177 ( \29554 , \29553 , \8019 );
nor \U$29178 ( \29555 , \29552 , \29554 );
nand \U$29179 ( \29556 , RIae775b8_79, \7631 );
and \U$29180 ( \29557 , \29556 , \7206 );
not \U$29181 ( \29558 , \29556 );
and \U$29182 ( \29559 , \29558 , \7205 );
nor \U$29183 ( \29560 , \29557 , \29559 );
xor \U$29184 ( \29561 , \29555 , \29560 );
and \U$29185 ( \29562 , \8966 , RIae773d8_75);
and \U$29186 ( \29563 , RIae77a68_89, \8964 );
nor \U$29187 ( \29564 , \29562 , \29563 );
and \U$29188 ( \29565 , \29564 , \8799 );
not \U$29189 ( \29566 , \29564 );
and \U$29190 ( \29567 , \29566 , \8789 );
nor \U$29191 ( \29568 , \29565 , \29567 );
and \U$29192 ( \29569 , \29561 , \29568 );
and \U$29193 ( \29570 , \29555 , \29560 );
or \U$29194 ( \29571 , \29569 , \29570 );
and \U$29195 ( \29572 , \29548 , \29571 );
and \U$29196 ( \29573 , \29540 , \29547 );
or \U$29197 ( \29574 , \29572 , \29573 );
xor \U$29198 ( \29575 , \29533 , \29574 );
xor \U$29199 ( \29576 , \29353 , \29360 );
xor \U$29200 ( \29577 , \29576 , \29368 );
xor \U$29201 ( \29578 , \29379 , \29386 );
xor \U$29202 ( \29579 , \29578 , \29394 );
and \U$29203 ( \29580 , \29577 , \29579 );
xor \U$29204 ( \29581 , \29328 , \29335 );
xor \U$29205 ( \29582 , \29581 , \29343 );
xor \U$29206 ( \29583 , \29379 , \29386 );
xor \U$29207 ( \29584 , \29583 , \29394 );
and \U$29208 ( \29585 , \29582 , \29584 );
and \U$29209 ( \29586 , \29577 , \29582 );
or \U$29210 ( \29587 , \29580 , \29585 , \29586 );
and \U$29211 ( \29588 , \29575 , \29587 );
and \U$29212 ( \29589 , \29533 , \29574 );
or \U$29213 ( \29590 , \29588 , \29589 );
xor \U$29214 ( \29591 , \29461 , \29590 );
xor \U$29215 ( \29592 , \29306 , \29311 );
xor \U$29216 ( \29593 , \29592 , \29318 );
and \U$29217 ( \29594 , \29591 , \29593 );
and \U$29218 ( \29595 , \29461 , \29590 );
or \U$29219 ( \29596 , \29594 , \29595 );
xor \U$29220 ( \29597 , \29448 , \29596 );
not \U$29221 ( \29598 , \29189 );
xor \U$29222 ( \29599 , \29174 , \29227 );
not \U$29223 ( \29600 , \29599 );
or \U$29224 ( \29601 , \29598 , \29600 );
or \U$29225 ( \29602 , \29599 , \29189 );
nand \U$29226 ( \29603 , \29601 , \29602 );
and \U$29227 ( \29604 , \29597 , \29603 );
and \U$29228 ( \29605 , \29448 , \29596 );
nor \U$29229 ( \29606 , \29604 , \29605 );
or \U$29230 ( \29607 , \29446 , \29606 );
xnor \U$29231 ( \29608 , \29606 , \29446 );
xor \U$29232 ( \29609 , \29448 , \29596 );
xor \U$29233 ( \29610 , \29609 , \29603 );
xor \U$29234 ( \29611 , \29400 , \29405 );
xor \U$29235 ( \29612 , \29611 , \29421 );
not \U$29236 ( \29613 , \29612 );
xor \U$29237 ( \29614 , \29461 , \29590 );
xor \U$29238 ( \29615 , \29614 , \29593 );
not \U$29239 ( \29616 , \29615 );
or \U$29240 ( \29617 , \29613 , \29616 );
or \U$29241 ( \29618 , \29615 , \29612 );
xor \U$29242 ( \29619 , \29555 , \29560 );
xor \U$29243 ( \29620 , \29619 , \29568 );
xor \U$29244 ( \29621 , \29512 , \29519 );
xor \U$29245 ( \29622 , \29621 , \29527 );
and \U$29246 ( \29623 , \29620 , \29622 );
xor \U$29247 ( \29624 , \29468 , \29475 );
xor \U$29248 ( \29625 , \29624 , \29483 );
xor \U$29249 ( \29626 , \29512 , \29519 );
xor \U$29250 ( \29627 , \29626 , \29527 );
and \U$29251 ( \29628 , \29625 , \29627 );
and \U$29252 ( \29629 , \29620 , \29625 );
or \U$29253 ( \29630 , \29623 , \29628 , \29629 );
and \U$29254 ( \29631 , \8966 , RIae77720_82);
and \U$29255 ( \29632 , RIae773d8_75, \8964 );
nor \U$29256 ( \29633 , \29631 , \29632 );
and \U$29257 ( \29634 , \29633 , \8799 );
not \U$29258 ( \29635 , \29633 );
and \U$29259 ( \29636 , \29635 , \8789 );
nor \U$29260 ( \29637 , \29634 , \29636 );
and \U$29261 ( \29638 , \9760 , RIae77a68_89);
and \U$29262 ( \29639 , RIae77978_87, \9758 );
nor \U$29263 ( \29640 , \29638 , \29639 );
and \U$29264 ( \29641 , \29640 , \9273 );
not \U$29265 ( \29642 , \29640 );
and \U$29266 ( \29643 , \29642 , \9764 );
nor \U$29267 ( \29644 , \29641 , \29643 );
xor \U$29268 ( \29645 , \29637 , \29644 );
and \U$29269 ( \29646 , \10548 , RIae77798_83);
and \U$29270 ( \29647 , RIae77888_85, \10546 );
nor \U$29271 ( \29648 , \29646 , \29647 );
and \U$29272 ( \29649 , \29648 , \10421 );
not \U$29273 ( \29650 , \29648 );
and \U$29274 ( \29651 , \29650 , \10118 );
nor \U$29275 ( \29652 , \29649 , \29651 );
and \U$29276 ( \29653 , \29645 , \29652 );
and \U$29277 ( \29654 , \29637 , \29644 );
or \U$29278 ( \29655 , \29653 , \29654 );
and \U$29279 ( \29656 , \14964 , RIae782d8_107);
and \U$29280 ( \29657 , RIae780f8_103, \14962 );
nor \U$29281 ( \29658 , \29656 , \29657 );
and \U$29282 ( \29659 , \29658 , \14463 );
not \U$29283 ( \29660 , \29658 );
and \U$29284 ( \29661 , \29660 , \14462 );
nor \U$29285 ( \29662 , \29659 , \29661 );
and \U$29286 ( \29663 , \15726 , RIae77f18_99);
and \U$29287 ( \29664 , RIae7aab0_192, RIae78008_101);
nor \U$29288 ( \29665 , \29663 , \29664 );
and \U$29289 ( \29666 , \29665 , \14959 );
not \U$29290 ( \29667 , \29665 );
and \U$29291 ( \29668 , \29667 , RIae7aa38_191);
nor \U$29292 ( \29669 , \29666 , \29668 );
xor \U$29293 ( \29670 , \29662 , \29669 );
and \U$29294 ( \29671 , \14059 , RIae771f8_71);
and \U$29295 ( \29672 , RIae772e8_73, \14057 );
nor \U$29296 ( \29673 , \29671 , \29672 );
and \U$29297 ( \29674 , \29673 , \13502 );
not \U$29298 ( \29675 , \29673 );
and \U$29299 ( \29676 , \29675 , \14063 );
nor \U$29300 ( \29677 , \29674 , \29676 );
and \U$29301 ( \29678 , \29670 , \29677 );
and \U$29302 ( \29679 , \29662 , \29669 );
or \U$29303 ( \29680 , \29678 , \29679 );
xor \U$29304 ( \29681 , \29655 , \29680 );
and \U$29305 ( \29682 , \13059 , RIae77180_70);
and \U$29306 ( \29683 , RIae77018_67, \13057 );
nor \U$29307 ( \29684 , \29682 , \29683 );
and \U$29308 ( \29685 , \29684 , \13063 );
not \U$29309 ( \29686 , \29684 );
and \U$29310 ( \29687 , \29686 , \12718 );
nor \U$29311 ( \29688 , \29685 , \29687 );
and \U$29312 ( \29689 , \11470 , RIae76f28_65);
and \U$29313 ( \29690 , RIae76e38_63, \11468 );
nor \U$29314 ( \29691 , \29689 , \29690 );
and \U$29315 ( \29692 , \29691 , \10936 );
not \U$29316 ( \29693 , \29691 );
and \U$29317 ( \29694 , \29693 , \11474 );
nor \U$29318 ( \29695 , \29692 , \29694 );
xor \U$29319 ( \29696 , \29688 , \29695 );
and \U$29320 ( \29697 , \12180 , RIae76d48_61);
and \U$29321 ( \29698 , RIae76c58_59, \12178 );
nor \U$29322 ( \29699 , \29697 , \29698 );
and \U$29323 ( \29700 , \29699 , \12184 );
not \U$29324 ( \29701 , \29699 );
and \U$29325 ( \29702 , \29701 , \11827 );
nor \U$29326 ( \29703 , \29700 , \29702 );
and \U$29327 ( \29704 , \29696 , \29703 );
and \U$29328 ( \29705 , \29688 , \29695 );
or \U$29329 ( \29706 , \29704 , \29705 );
and \U$29330 ( \29707 , \29681 , \29706 );
and \U$29331 ( \29708 , \29655 , \29680 );
or \U$29332 ( \29709 , \29707 , \29708 );
xor \U$29333 ( \29710 , \29630 , \29709 );
xor \U$29334 ( \29711 , \29379 , \29386 );
xor \U$29335 ( \29712 , \29711 , \29394 );
xor \U$29336 ( \29713 , \29577 , \29582 );
xor \U$29337 ( \29714 , \29712 , \29713 );
and \U$29338 ( \29715 , \29710 , \29714 );
and \U$29339 ( \29716 , \29630 , \29709 );
or \U$29340 ( \29717 , \29715 , \29716 );
xor \U$29341 ( \29718 , \29533 , \29574 );
xor \U$29342 ( \29719 , \29718 , \29587 );
and \U$29343 ( \29720 , \29717 , \29719 );
xor \U$29344 ( \29721 , \29346 , \29371 );
xor \U$29345 ( \29722 , \29721 , \29397 );
xor \U$29346 ( \29723 , \29449 , \29456 );
xor \U$29347 ( \29724 , \29722 , \29723 );
xor \U$29348 ( \29725 , \29533 , \29574 );
xor \U$29349 ( \29726 , \29725 , \29587 );
and \U$29350 ( \29727 , \29724 , \29726 );
and \U$29351 ( \29728 , \29717 , \29724 );
or \U$29352 ( \29729 , \29720 , \29727 , \29728 );
nand \U$29353 ( \29730 , \29618 , \29729 );
nand \U$29354 ( \29731 , \29617 , \29730 );
and \U$29355 ( \29732 , \29610 , \29731 );
xor \U$29356 ( \29733 , \29731 , \29610 );
xnor \U$29357 ( \29734 , \29612 , \29729 );
not \U$29358 ( \29735 , \29734 );
not \U$29359 ( \29736 , \29615 );
and \U$29360 ( \29737 , \29735 , \29736 );
and \U$29361 ( \29738 , \29734 , \29615 );
nor \U$29362 ( \29739 , \29737 , \29738 );
xor \U$29363 ( \29740 , \29533 , \29574 );
xor \U$29364 ( \29741 , \29740 , \29587 );
xor \U$29365 ( \29742 , \29717 , \29724 );
xor \U$29366 ( \29743 , \29741 , \29742 );
xor \U$29367 ( \29744 , \29486 , \29504 );
xor \U$29368 ( \29745 , \29744 , \29530 );
xor \U$29369 ( \29746 , \29630 , \29709 );
xor \U$29370 ( \29747 , \29746 , \29714 );
and \U$29371 ( \29748 , \29745 , \29747 );
xor \U$29372 ( \29749 , \29743 , \29748 );
xor \U$29373 ( \29750 , \29655 , \29680 );
xor \U$29374 ( \29751 , \29750 , \29706 );
xor \U$29375 ( \29752 , \29512 , \29519 );
xor \U$29376 ( \29753 , \29752 , \29527 );
xor \U$29377 ( \29754 , \29620 , \29625 );
xor \U$29378 ( \29755 , \29753 , \29754 );
and \U$29379 ( \29756 , \29751 , \29755 );
xor \U$29380 ( \29757 , \29540 , \29547 );
xor \U$29381 ( \29758 , \29757 , \29571 );
xor \U$29382 ( \29759 , \29756 , \29758 );
and \U$29383 ( \29760 , \9760 , RIae773d8_75);
and \U$29384 ( \29761 , RIae77a68_89, \9758 );
nor \U$29385 ( \29762 , \29760 , \29761 );
and \U$29386 ( \29763 , \29762 , \9273 );
not \U$29387 ( \29764 , \29762 );
and \U$29388 ( \29765 , \29764 , \9764 );
nor \U$29389 ( \29766 , \29763 , \29765 );
and \U$29390 ( \29767 , \10548 , RIae77978_87);
and \U$29391 ( \29768 , RIae77798_83, \10546 );
nor \U$29392 ( \29769 , \29767 , \29768 );
and \U$29393 ( \29770 , \29769 , \10421 );
not \U$29394 ( \29771 , \29769 );
and \U$29395 ( \29772 , \29771 , \10118 );
nor \U$29396 ( \29773 , \29770 , \29772 );
xor \U$29397 ( \29774 , \29766 , \29773 );
and \U$29398 ( \29775 , \11470 , RIae77888_85);
and \U$29399 ( \29776 , RIae76f28_65, \11468 );
nor \U$29400 ( \29777 , \29775 , \29776 );
and \U$29401 ( \29778 , \29777 , \10936 );
not \U$29402 ( \29779 , \29777 );
and \U$29403 ( \29780 , \29779 , \11474 );
nor \U$29404 ( \29781 , \29778 , \29780 );
and \U$29405 ( \29782 , \29774 , \29781 );
and \U$29406 ( \29783 , \29766 , \29773 );
or \U$29407 ( \29784 , \29782 , \29783 );
and \U$29408 ( \29785 , \15726 , RIae780f8_103);
and \U$29409 ( \29786 , RIae7aab0_192, RIae77f18_99);
nor \U$29410 ( \29787 , \29785 , \29786 );
and \U$29411 ( \29788 , \29787 , \14959 );
not \U$29412 ( \29789 , \29787 );
and \U$29413 ( \29790 , \29789 , RIae7aa38_191);
nor \U$29414 ( \29791 , \29788 , \29790 );
xor \U$29415 ( \29792 , \29791 , \8019 );
and \U$29416 ( \29793 , \14964 , RIae772e8_73);
and \U$29417 ( \29794 , RIae782d8_107, \14962 );
nor \U$29418 ( \29795 , \29793 , \29794 );
and \U$29419 ( \29796 , \29795 , \14463 );
not \U$29420 ( \29797 , \29795 );
and \U$29421 ( \29798 , \29797 , \14462 );
nor \U$29422 ( \29799 , \29796 , \29798 );
and \U$29423 ( \29800 , \29792 , \29799 );
and \U$29424 ( \29801 , \29791 , \8019 );
or \U$29425 ( \29802 , \29800 , \29801 );
xor \U$29426 ( \29803 , \29784 , \29802 );
and \U$29427 ( \29804 , \12180 , RIae76e38_63);
and \U$29428 ( \29805 , RIae76d48_61, \12178 );
nor \U$29429 ( \29806 , \29804 , \29805 );
and \U$29430 ( \29807 , \29806 , \12184 );
not \U$29431 ( \29808 , \29806 );
and \U$29432 ( \29809 , \29808 , \11827 );
nor \U$29433 ( \29810 , \29807 , \29809 );
and \U$29434 ( \29811 , \13059 , RIae76c58_59);
and \U$29435 ( \29812 , RIae77180_70, \13057 );
nor \U$29436 ( \29813 , \29811 , \29812 );
and \U$29437 ( \29814 , \29813 , \13063 );
not \U$29438 ( \29815 , \29813 );
and \U$29439 ( \29816 , \29815 , \12718 );
nor \U$29440 ( \29817 , \29814 , \29816 );
xor \U$29441 ( \29818 , \29810 , \29817 );
and \U$29442 ( \29819 , \14059 , RIae77018_67);
and \U$29443 ( \29820 , RIae771f8_71, \14057 );
nor \U$29444 ( \29821 , \29819 , \29820 );
and \U$29445 ( \29822 , \29821 , \13502 );
not \U$29446 ( \29823 , \29821 );
and \U$29447 ( \29824 , \29823 , \14063 );
nor \U$29448 ( \29825 , \29822 , \29824 );
and \U$29449 ( \29826 , \29818 , \29825 );
and \U$29450 ( \29827 , \29810 , \29817 );
or \U$29451 ( \29828 , \29826 , \29827 );
and \U$29452 ( \29829 , \29803 , \29828 );
and \U$29453 ( \29830 , \29784 , \29802 );
or \U$29454 ( \29831 , \29829 , \29830 );
xor \U$29455 ( \29832 , \29493 , \7205 );
xor \U$29456 ( \29833 , \29832 , \29501 );
xor \U$29457 ( \29834 , \29831 , \29833 );
and \U$29458 ( \29835 , \8371 , RIae775b8_79);
and \U$29459 ( \29836 , RIae774c8_77, \8369 );
nor \U$29460 ( \29837 , \29835 , \29836 );
and \U$29461 ( \29838 , \29837 , \8020 );
not \U$29462 ( \29839 , \29837 );
and \U$29463 ( \29840 , \29839 , \8019 );
nor \U$29464 ( \29841 , \29838 , \29840 );
xor \U$29465 ( \29842 , \29637 , \29644 );
xor \U$29466 ( \29843 , \29842 , \29652 );
and \U$29467 ( \29844 , \29841 , \29843 );
xor \U$29468 ( \29845 , \29688 , \29695 );
xor \U$29469 ( \29846 , \29845 , \29703 );
xor \U$29470 ( \29847 , \29637 , \29644 );
xor \U$29471 ( \29848 , \29847 , \29652 );
and \U$29472 ( \29849 , \29846 , \29848 );
and \U$29473 ( \29850 , \29841 , \29846 );
or \U$29474 ( \29851 , \29844 , \29849 , \29850 );
and \U$29475 ( \29852 , \29834 , \29851 );
and \U$29476 ( \29853 , \29831 , \29833 );
or \U$29477 ( \29854 , \29852 , \29853 );
and \U$29478 ( \29855 , \29759 , \29854 );
and \U$29479 ( \29856 , \29756 , \29758 );
or \U$29480 ( \29857 , \29855 , \29856 );
and \U$29481 ( \29858 , \29749 , \29857 );
and \U$29482 ( \29859 , \29743 , \29748 );
nor \U$29483 ( \29860 , \29858 , \29859 );
or \U$29484 ( \29861 , \29739 , \29860 );
xnor \U$29485 ( \29862 , \29860 , \29739 );
xor \U$29486 ( \29863 , \29791 , \8019 );
xor \U$29487 ( \29864 , \29863 , \29799 );
and \U$29488 ( \29865 , \8966 , RIae774c8_77);
and \U$29489 ( \29866 , RIae77720_82, \8964 );
nor \U$29490 ( \29867 , \29865 , \29866 );
and \U$29491 ( \29868 , \29867 , \8799 );
not \U$29492 ( \29869 , \29867 );
and \U$29493 ( \29870 , \29869 , \8789 );
nor \U$29494 ( \29871 , \29868 , \29870 );
nand \U$29495 ( \29872 , RIae775b8_79, \8369 );
and \U$29496 ( \29873 , \29872 , \8020 );
not \U$29497 ( \29874 , \29872 );
and \U$29498 ( \29875 , \29874 , \8019 );
nor \U$29499 ( \29876 , \29873 , \29875 );
xor \U$29500 ( \29877 , \29871 , \29876 );
xor \U$29501 ( \29878 , \29766 , \29773 );
xor \U$29502 ( \29879 , \29878 , \29781 );
xor \U$29503 ( \29880 , \29877 , \29879 );
and \U$29504 ( \29881 , \29864 , \29880 );
and \U$29505 ( \29882 , \12180 , RIae76f28_65);
and \U$29506 ( \29883 , RIae76e38_63, \12178 );
nor \U$29507 ( \29884 , \29882 , \29883 );
and \U$29508 ( \29885 , \29884 , \12184 );
not \U$29509 ( \29886 , \29884 );
and \U$29510 ( \29887 , \29886 , \11827 );
nor \U$29511 ( \29888 , \29885 , \29887 );
and \U$29512 ( \29889 , \11470 , RIae77798_83);
and \U$29513 ( \29890 , RIae77888_85, \11468 );
nor \U$29514 ( \29891 , \29889 , \29890 );
and \U$29515 ( \29892 , \29891 , \10936 );
not \U$29516 ( \29893 , \29891 );
and \U$29517 ( \29894 , \29893 , \11474 );
nor \U$29518 ( \29895 , \29892 , \29894 );
xor \U$29519 ( \29896 , \29888 , \29895 );
and \U$29520 ( \29897 , \13059 , RIae76d48_61);
and \U$29521 ( \29898 , RIae76c58_59, \13057 );
nor \U$29522 ( \29899 , \29897 , \29898 );
and \U$29523 ( \29900 , \29899 , \13063 );
not \U$29524 ( \29901 , \29899 );
and \U$29525 ( \29902 , \29901 , \12718 );
nor \U$29526 ( \29903 , \29900 , \29902 );
and \U$29527 ( \29904 , \29896 , \29903 );
and \U$29528 ( \29905 , \29888 , \29895 );
or \U$29529 ( \29906 , \29904 , \29905 );
and \U$29530 ( \29907 , \14059 , RIae77180_70);
and \U$29531 ( \29908 , RIae77018_67, \14057 );
nor \U$29532 ( \29909 , \29907 , \29908 );
and \U$29533 ( \29910 , \29909 , \14063 );
not \U$29534 ( \29911 , \29909 );
and \U$29535 ( \29912 , \29911 , \13502 );
nor \U$29536 ( \29913 , \29910 , \29912 );
and \U$29537 ( \29914 , \15726 , RIae782d8_107);
and \U$29538 ( \29915 , RIae7aab0_192, RIae780f8_103);
nor \U$29539 ( \29916 , \29914 , \29915 );
and \U$29540 ( \29917 , \29916 , RIae7aa38_191);
not \U$29541 ( \29918 , \29916 );
and \U$29542 ( \29919 , \29918 , \14959 );
nor \U$29543 ( \29920 , \29917 , \29919 );
or \U$29544 ( \29921 , \29913 , \29920 );
not \U$29545 ( \29922 , \29920 );
not \U$29546 ( \29923 , \29913 );
or \U$29547 ( \29924 , \29922 , \29923 );
and \U$29548 ( \29925 , \14964 , RIae771f8_71);
and \U$29549 ( \29926 , RIae772e8_73, \14962 );
nor \U$29550 ( \29927 , \29925 , \29926 );
and \U$29551 ( \29928 , \29927 , \14463 );
not \U$29552 ( \29929 , \29927 );
and \U$29553 ( \29930 , \29929 , \14462 );
nor \U$29554 ( \29931 , \29928 , \29930 );
nand \U$29555 ( \29932 , \29924 , \29931 );
nand \U$29556 ( \29933 , \29921 , \29932 );
xor \U$29557 ( \29934 , \29906 , \29933 );
and \U$29558 ( \29935 , \8966 , RIae775b8_79);
and \U$29559 ( \29936 , RIae774c8_77, \8964 );
nor \U$29560 ( \29937 , \29935 , \29936 );
and \U$29561 ( \29938 , \29937 , \8789 );
not \U$29562 ( \29939 , \29937 );
and \U$29563 ( \29940 , \29939 , \8799 );
nor \U$29564 ( \29941 , \29938 , \29940 );
and \U$29565 ( \29942 , \9760 , RIae77720_82);
and \U$29566 ( \29943 , RIae773d8_75, \9758 );
nor \U$29567 ( \29944 , \29942 , \29943 );
and \U$29568 ( \29945 , \29944 , \9272 );
not \U$29569 ( \29946 , \29944 );
and \U$29570 ( \29947 , \29946 , \9273 );
nor \U$29571 ( \29948 , \29945 , \29947 );
or \U$29572 ( \29949 , \29941 , \29948 );
not \U$29573 ( \29950 , \29948 );
not \U$29574 ( \29951 , \29941 );
or \U$29575 ( \29952 , \29950 , \29951 );
and \U$29576 ( \29953 , \10548 , RIae77a68_89);
and \U$29577 ( \29954 , RIae77978_87, \10546 );
nor \U$29578 ( \29955 , \29953 , \29954 );
and \U$29579 ( \29956 , \29955 , \10421 );
not \U$29580 ( \29957 , \29955 );
and \U$29581 ( \29958 , \29957 , \10118 );
nor \U$29582 ( \29959 , \29956 , \29958 );
nand \U$29583 ( \29960 , \29952 , \29959 );
nand \U$29584 ( \29961 , \29949 , \29960 );
xor \U$29585 ( \29962 , \29934 , \29961 );
xor \U$29586 ( \29963 , \29871 , \29876 );
xor \U$29587 ( \29964 , \29963 , \29879 );
and \U$29588 ( \29965 , \29962 , \29964 );
and \U$29589 ( \29966 , \29864 , \29962 );
or \U$29590 ( \29967 , \29881 , \29965 , \29966 );
xor \U$29591 ( \29968 , \29637 , \29644 );
xor \U$29592 ( \29969 , \29968 , \29652 );
xor \U$29593 ( \29970 , \29841 , \29846 );
xor \U$29594 ( \29971 , \29969 , \29970 );
xor \U$29595 ( \29972 , \29967 , \29971 );
and \U$29596 ( \29973 , \13059 , RIae76e38_63);
and \U$29597 ( \29974 , RIae76d48_61, \13057 );
nor \U$29598 ( \29975 , \29973 , \29974 );
and \U$29599 ( \29976 , \29975 , \13063 );
not \U$29600 ( \29977 , \29975 );
and \U$29601 ( \29978 , \29977 , \12718 );
nor \U$29602 ( \29979 , \29976 , \29978 );
and \U$29603 ( \29980 , \12180 , RIae77888_85);
and \U$29604 ( \29981 , RIae76f28_65, \12178 );
nor \U$29605 ( \29982 , \29980 , \29981 );
and \U$29606 ( \29983 , \29982 , \12184 );
not \U$29607 ( \29984 , \29982 );
and \U$29608 ( \29985 , \29984 , \11827 );
nor \U$29609 ( \29986 , \29983 , \29985 );
xor \U$29610 ( \29987 , \29979 , \29986 );
and \U$29611 ( \29988 , \14059 , RIae76c58_59);
and \U$29612 ( \29989 , RIae77180_70, \14057 );
nor \U$29613 ( \29990 , \29988 , \29989 );
and \U$29614 ( \29991 , \29990 , \13502 );
not \U$29615 ( \29992 , \29990 );
and \U$29616 ( \29993 , \29992 , \14063 );
nor \U$29617 ( \29994 , \29991 , \29993 );
and \U$29618 ( \29995 , \29987 , \29994 );
and \U$29619 ( \29996 , \29979 , \29986 );
or \U$29620 ( \29997 , \29995 , \29996 );
and \U$29621 ( \29998 , \15726 , RIae772e8_73);
and \U$29622 ( \29999 , RIae7aab0_192, RIae782d8_107);
nor \U$29623 ( \30000 , \29998 , \29999 );
and \U$29624 ( \30001 , \30000 , \14959 );
not \U$29625 ( \30002 , \30000 );
and \U$29626 ( \30003 , \30002 , RIae7aa38_191);
nor \U$29627 ( \30004 , \30001 , \30003 );
xor \U$29628 ( \30005 , \30004 , \8789 );
and \U$29629 ( \30006 , \14964 , RIae77018_67);
and \U$29630 ( \30007 , RIae771f8_71, \14962 );
nor \U$29631 ( \30008 , \30006 , \30007 );
and \U$29632 ( \30009 , \30008 , \14463 );
not \U$29633 ( \30010 , \30008 );
and \U$29634 ( \30011 , \30010 , \14462 );
nor \U$29635 ( \30012 , \30009 , \30011 );
and \U$29636 ( \30013 , \30005 , \30012 );
and \U$29637 ( \30014 , \30004 , \8789 );
or \U$29638 ( \30015 , \30013 , \30014 );
xor \U$29639 ( \30016 , \29997 , \30015 );
and \U$29640 ( \30017 , \9760 , RIae774c8_77);
and \U$29641 ( \30018 , RIae77720_82, \9758 );
nor \U$29642 ( \30019 , \30017 , \30018 );
and \U$29643 ( \30020 , \30019 , \9273 );
not \U$29644 ( \30021 , \30019 );
and \U$29645 ( \30022 , \30021 , \9272 );
nor \U$29646 ( \30023 , \30020 , \30022 );
and \U$29647 ( \30024 , \10548 , RIae773d8_75);
and \U$29648 ( \30025 , RIae77a68_89, \10546 );
nor \U$29649 ( \30026 , \30024 , \30025 );
and \U$29650 ( \30027 , \30026 , \10421 );
not \U$29651 ( \30028 , \30026 );
and \U$29652 ( \30029 , \30028 , \10118 );
nor \U$29653 ( \30030 , \30027 , \30029 );
xor \U$29654 ( \30031 , \30023 , \30030 );
and \U$29655 ( \30032 , \11470 , RIae77978_87);
and \U$29656 ( \30033 , RIae77798_83, \11468 );
nor \U$29657 ( \30034 , \30032 , \30033 );
and \U$29658 ( \30035 , \30034 , \10936 );
not \U$29659 ( \30036 , \30034 );
and \U$29660 ( \30037 , \30036 , \11474 );
nor \U$29661 ( \30038 , \30035 , \30037 );
and \U$29662 ( \30039 , \30031 , \30038 );
and \U$29663 ( \30040 , \30023 , \30030 );
or \U$29664 ( \30041 , \30039 , \30040 );
and \U$29665 ( \30042 , \30016 , \30041 );
and \U$29666 ( \30043 , \29997 , \30015 );
or \U$29667 ( \30044 , \30042 , \30043 );
xor \U$29668 ( \30045 , \29810 , \29817 );
xor \U$29669 ( \30046 , \30045 , \29825 );
xor \U$29670 ( \30047 , \30044 , \30046 );
not \U$29671 ( \30048 , \29920 );
not \U$29672 ( \30049 , \29931 );
or \U$29673 ( \30050 , \30048 , \30049 );
or \U$29674 ( \30051 , \29931 , \29920 );
nand \U$29675 ( \30052 , \30050 , \30051 );
not \U$29676 ( \30053 , \30052 );
not \U$29677 ( \30054 , \29913 );
and \U$29678 ( \30055 , \30053 , \30054 );
and \U$29679 ( \30056 , \30052 , \29913 );
nor \U$29680 ( \30057 , \30055 , \30056 );
not \U$29681 ( \30058 , \29948 );
not \U$29682 ( \30059 , \29959 );
or \U$29683 ( \30060 , \30058 , \30059 );
or \U$29684 ( \30061 , \29948 , \29959 );
nand \U$29685 ( \30062 , \30060 , \30061 );
not \U$29686 ( \30063 , \30062 );
not \U$29687 ( \30064 , \29941 );
and \U$29688 ( \30065 , \30063 , \30064 );
and \U$29689 ( \30066 , \30062 , \29941 );
nor \U$29690 ( \30067 , \30065 , \30066 );
or \U$29691 ( \30068 , \30057 , \30067 );
not \U$29692 ( \30069 , \30067 );
not \U$29693 ( \30070 , \30057 );
or \U$29694 ( \30071 , \30069 , \30070 );
xor \U$29695 ( \30072 , \29888 , \29895 );
xor \U$29696 ( \30073 , \30072 , \29903 );
nand \U$29697 ( \30074 , \30071 , \30073 );
nand \U$29698 ( \30075 , \30068 , \30074 );
and \U$29699 ( \30076 , \30047 , \30075 );
and \U$29700 ( \30077 , \30044 , \30046 );
or \U$29701 ( \30078 , \30076 , \30077 );
xor \U$29702 ( \30079 , \29972 , \30078 );
xor \U$29703 ( \30080 , \30044 , \30046 );
xor \U$29704 ( \30081 , \30080 , \30075 );
not \U$29705 ( \30082 , \30081 );
xor \U$29706 ( \30083 , \29871 , \29876 );
xor \U$29707 ( \30084 , \30083 , \29879 );
xor \U$29708 ( \30085 , \29864 , \29962 );
xor \U$29709 ( \30086 , \30084 , \30085 );
not \U$29710 ( \30087 , \30086 );
or \U$29711 ( \30088 , \30082 , \30087 );
or \U$29712 ( \30089 , \30086 , \30081 );
not \U$29713 ( \30090 , \30073 );
not \U$29714 ( \30091 , \30057 );
or \U$29715 ( \30092 , \30090 , \30091 );
or \U$29716 ( \30093 , \30057 , \30073 );
nand \U$29717 ( \30094 , \30092 , \30093 );
not \U$29718 ( \30095 , \30094 );
not \U$29719 ( \30096 , \30067 );
and \U$29720 ( \30097 , \30095 , \30096 );
and \U$29721 ( \30098 , \30094 , \30067 );
nor \U$29722 ( \30099 , \30097 , \30098 );
and \U$29723 ( \30100 , \14964 , RIae77180_70);
and \U$29724 ( \30101 , RIae77018_67, \14962 );
nor \U$29725 ( \30102 , \30100 , \30101 );
and \U$29726 ( \30103 , \30102 , \14463 );
not \U$29727 ( \30104 , \30102 );
and \U$29728 ( \30105 , \30104 , \14462 );
nor \U$29729 ( \30106 , \30103 , \30105 );
and \U$29730 ( \30107 , \15726 , RIae771f8_71);
and \U$29731 ( \30108 , RIae7aab0_192, RIae772e8_73);
nor \U$29732 ( \30109 , \30107 , \30108 );
and \U$29733 ( \30110 , \30109 , \14959 );
not \U$29734 ( \30111 , \30109 );
and \U$29735 ( \30112 , \30111 , RIae7aa38_191);
nor \U$29736 ( \30113 , \30110 , \30112 );
xor \U$29737 ( \30114 , \30106 , \30113 );
and \U$29738 ( \30115 , \14059 , RIae76d48_61);
and \U$29739 ( \30116 , RIae76c58_59, \14057 );
nor \U$29740 ( \30117 , \30115 , \30116 );
and \U$29741 ( \30118 , \30117 , \13502 );
not \U$29742 ( \30119 , \30117 );
and \U$29743 ( \30120 , \30119 , \14063 );
nor \U$29744 ( \30121 , \30118 , \30120 );
and \U$29745 ( \30122 , \30114 , \30121 );
and \U$29746 ( \30123 , \30106 , \30113 );
nor \U$29747 ( \30124 , \30122 , \30123 );
not \U$29748 ( \30125 , \30124 );
and \U$29749 ( \30126 , \9760 , RIae775b8_79);
and \U$29750 ( \30127 , RIae774c8_77, \9758 );
nor \U$29751 ( \30128 , \30126 , \30127 );
and \U$29752 ( \30129 , \30128 , \9272 );
not \U$29753 ( \30130 , \30128 );
and \U$29754 ( \30131 , \30130 , \9273 );
nor \U$29755 ( \30132 , \30129 , \30131 );
not \U$29756 ( \30133 , \30132 );
and \U$29757 ( \30134 , \10548 , RIae77720_82);
and \U$29758 ( \30135 , RIae773d8_75, \10546 );
nor \U$29759 ( \30136 , \30134 , \30135 );
and \U$29760 ( \30137 , \30136 , \10421 );
not \U$29761 ( \30138 , \30136 );
and \U$29762 ( \30139 , \30138 , \10118 );
nor \U$29763 ( \30140 , \30137 , \30139 );
nand \U$29764 ( \30141 , \30133 , \30140 );
not \U$29765 ( \30142 , \30141 );
and \U$29766 ( \30143 , \30125 , \30142 );
and \U$29767 ( \30144 , \30124 , \30141 );
and \U$29768 ( \30145 , \12180 , RIae77798_83);
and \U$29769 ( \30146 , RIae77888_85, \12178 );
nor \U$29770 ( \30147 , \30145 , \30146 );
and \U$29771 ( \30148 , \30147 , \12184 );
not \U$29772 ( \30149 , \30147 );
and \U$29773 ( \30150 , \30149 , \11827 );
nor \U$29774 ( \30151 , \30148 , \30150 );
and \U$29775 ( \30152 , \13059 , RIae76f28_65);
and \U$29776 ( \30153 , RIae76e38_63, \13057 );
nor \U$29777 ( \30154 , \30152 , \30153 );
and \U$29778 ( \30155 , \30154 , \13063 );
not \U$29779 ( \30156 , \30154 );
and \U$29780 ( \30157 , \30156 , \12718 );
nor \U$29781 ( \30158 , \30155 , \30157 );
xor \U$29782 ( \30159 , \30151 , \30158 );
and \U$29783 ( \30160 , \11470 , RIae77a68_89);
and \U$29784 ( \30161 , RIae77978_87, \11468 );
nor \U$29785 ( \30162 , \30160 , \30161 );
and \U$29786 ( \30163 , \30162 , \10936 );
not \U$29787 ( \30164 , \30162 );
and \U$29788 ( \30165 , \30164 , \11474 );
nor \U$29789 ( \30166 , \30163 , \30165 );
and \U$29790 ( \30167 , \30159 , \30166 );
and \U$29791 ( \30168 , \30151 , \30158 );
nor \U$29792 ( \30169 , \30167 , \30168 );
nor \U$29793 ( \30170 , \30144 , \30169 );
nor \U$29794 ( \30171 , \30143 , \30170 );
or \U$29795 ( \30172 , \30099 , \30171 );
not \U$29796 ( \30173 , \30171 );
not \U$29797 ( \30174 , \30099 );
or \U$29798 ( \30175 , \30173 , \30174 );
nand \U$29799 ( \30176 , RIae775b8_79, \8964 );
and \U$29800 ( \30177 , \30176 , \8799 );
not \U$29801 ( \30178 , \30176 );
and \U$29802 ( \30179 , \30178 , \8789 );
nor \U$29803 ( \30180 , \30177 , \30179 );
xor \U$29804 ( \30181 , \29979 , \29986 );
xor \U$29805 ( \30182 , \30181 , \29994 );
and \U$29806 ( \30183 , \30180 , \30182 );
xor \U$29807 ( \30184 , \30023 , \30030 );
xor \U$29808 ( \30185 , \30184 , \30038 );
xor \U$29809 ( \30186 , \29979 , \29986 );
xor \U$29810 ( \30187 , \30186 , \29994 );
and \U$29811 ( \30188 , \30185 , \30187 );
and \U$29812 ( \30189 , \30180 , \30185 );
or \U$29813 ( \30190 , \30183 , \30188 , \30189 );
nand \U$29814 ( \30191 , \30175 , \30190 );
nand \U$29815 ( \30192 , \30172 , \30191 );
nand \U$29816 ( \30193 , \30089 , \30192 );
nand \U$29817 ( \30194 , \30088 , \30193 );
xnor \U$29818 ( \30195 , \30079 , \30194 );
not \U$29819 ( \30196 , \30195 );
xor \U$29820 ( \30197 , \29784 , \29802 );
xor \U$29821 ( \30198 , \30197 , \29828 );
xor \U$29822 ( \30199 , \29871 , \29876 );
and \U$29823 ( \30200 , \30199 , \29879 );
and \U$29824 ( \30201 , \29871 , \29876 );
or \U$29825 ( \30202 , \30200 , \30201 );
xor \U$29826 ( \30203 , \29662 , \29669 );
xor \U$29827 ( \30204 , \30203 , \29677 );
xor \U$29828 ( \30205 , \30202 , \30204 );
xor \U$29829 ( \30206 , \29906 , \29933 );
and \U$29830 ( \30207 , \30206 , \29961 );
and \U$29831 ( \30208 , \29906 , \29933 );
or \U$29832 ( \30209 , \30207 , \30208 );
xor \U$29833 ( \30210 , \30205 , \30209 );
xor \U$29834 ( \30211 , \30198 , \30210 );
not \U$29835 ( \30212 , \30211 );
and \U$29836 ( \30213 , \30196 , \30212 );
and \U$29837 ( \30214 , \30195 , \30211 );
nor \U$29838 ( \30215 , \30213 , \30214 );
xnor \U$29839 ( \30216 , \30192 , \30081 );
not \U$29840 ( \30217 , \30216 );
not \U$29841 ( \30218 , \30086 );
and \U$29842 ( \30219 , \30217 , \30218 );
and \U$29843 ( \30220 , \30216 , \30086 );
nor \U$29844 ( \30221 , \30219 , \30220 );
not \U$29845 ( \30222 , \30221 );
not \U$29846 ( \30223 , \30141 );
xor \U$29847 ( \30224 , \30124 , \30169 );
not \U$29848 ( \30225 , \30224 );
or \U$29849 ( \30226 , \30223 , \30225 );
or \U$29850 ( \30227 , \30224 , \30141 );
nand \U$29851 ( \30228 , \30226 , \30227 );
xor \U$29852 ( \30229 , \29979 , \29986 );
xor \U$29853 ( \30230 , \30229 , \29994 );
xor \U$29854 ( \30231 , \30180 , \30185 );
xor \U$29855 ( \30232 , \30230 , \30231 );
and \U$29856 ( \30233 , \30228 , \30232 );
xor \U$29857 ( \30234 , \29997 , \30015 );
xor \U$29858 ( \30235 , \30234 , \30041 );
xor \U$29859 ( \30236 , \30233 , \30235 );
and \U$29860 ( \30237 , \12180 , RIae77978_87);
and \U$29861 ( \30238 , RIae77798_83, \12178 );
nor \U$29862 ( \30239 , \30237 , \30238 );
and \U$29863 ( \30240 , \30239 , \11827 );
not \U$29864 ( \30241 , \30239 );
and \U$29865 ( \30242 , \30241 , \12184 );
nor \U$29866 ( \30243 , \30240 , \30242 );
and \U$29867 ( \30244 , \13059 , RIae77888_85);
and \U$29868 ( \30245 , RIae76f28_65, \13057 );
nor \U$29869 ( \30246 , \30244 , \30245 );
and \U$29870 ( \30247 , \30246 , \12718 );
not \U$29871 ( \30248 , \30246 );
and \U$29872 ( \30249 , \30248 , \13063 );
nor \U$29873 ( \30250 , \30247 , \30249 );
xor \U$29874 ( \30251 , \30243 , \30250 );
and \U$29875 ( \30252 , \14059 , RIae76e38_63);
and \U$29876 ( \30253 , RIae76d48_61, \14057 );
nor \U$29877 ( \30254 , \30252 , \30253 );
and \U$29878 ( \30255 , \30254 , \14063 );
not \U$29879 ( \30256 , \30254 );
and \U$29880 ( \30257 , \30256 , \13502 );
nor \U$29881 ( \30258 , \30255 , \30257 );
and \U$29882 ( \30259 , \30251 , \30258 );
and \U$29883 ( \30260 , \30243 , \30250 );
or \U$29884 ( \30261 , \30259 , \30260 );
and \U$29885 ( \30262 , \15726 , RIae77018_67);
and \U$29886 ( \30263 , RIae7aab0_192, RIae771f8_71);
nor \U$29887 ( \30264 , \30262 , \30263 );
and \U$29888 ( \30265 , \30264 , \14959 );
not \U$29889 ( \30266 , \30264 );
and \U$29890 ( \30267 , \30266 , RIae7aa38_191);
nor \U$29891 ( \30268 , \30265 , \30267 );
and \U$29892 ( \30269 , \30268 , \9764 );
not \U$29893 ( \30270 , \30268 );
not \U$29894 ( \30271 , \9272 );
and \U$29895 ( \30272 , \30270 , \30271 );
and \U$29896 ( \30273 , \14964 , RIae76c58_59);
and \U$29897 ( \30274 , RIae77180_70, \14962 );
nor \U$29898 ( \30275 , \30273 , \30274 );
and \U$29899 ( \30276 , \30275 , \14462 );
not \U$29900 ( \30277 , \30275 );
and \U$29901 ( \30278 , \30277 , \14463 );
nor \U$29902 ( \30279 , \30276 , \30278 );
nor \U$29903 ( \30280 , \30272 , \30279 );
nor \U$29904 ( \30281 , \30269 , \30280 );
or \U$29905 ( \30282 , \30261 , \30281 );
not \U$29906 ( \30283 , \30281 );
not \U$29907 ( \30284 , \30261 );
or \U$29908 ( \30285 , \30283 , \30284 );
nand \U$29909 ( \30286 , RIae775b8_79, \9758 );
and \U$29910 ( \30287 , \30286 , \9273 );
not \U$29911 ( \30288 , \30286 );
and \U$29912 ( \30289 , \30288 , \9764 );
nor \U$29913 ( \30290 , \30287 , \30289 );
not \U$29914 ( \30291 , \30290 );
and \U$29915 ( \30292 , \10548 , RIae774c8_77);
and \U$29916 ( \30293 , RIae77720_82, \10546 );
nor \U$29917 ( \30294 , \30292 , \30293 );
and \U$29918 ( \30295 , \30294 , \10421 );
not \U$29919 ( \30296 , \30294 );
and \U$29920 ( \30297 , \30296 , \10118 );
nor \U$29921 ( \30298 , \30295 , \30297 );
not \U$29922 ( \30299 , \30298 );
or \U$29923 ( \30300 , \30291 , \30299 );
or \U$29924 ( \30301 , \30298 , \30290 );
and \U$29925 ( \30302 , \11470 , RIae773d8_75);
and \U$29926 ( \30303 , RIae77a68_89, \11468 );
nor \U$29927 ( \30304 , \30302 , \30303 );
and \U$29928 ( \30305 , \30304 , \10936 );
not \U$29929 ( \30306 , \30304 );
and \U$29930 ( \30307 , \30306 , \11474 );
nor \U$29931 ( \30308 , \30305 , \30307 );
nand \U$29932 ( \30309 , \30301 , \30308 );
nand \U$29933 ( \30310 , \30300 , \30309 );
nand \U$29934 ( \30311 , \30285 , \30310 );
nand \U$29935 ( \30312 , \30282 , \30311 );
xor \U$29936 ( \30313 , \30004 , \8789 );
xor \U$29937 ( \30314 , \30313 , \30012 );
xor \U$29938 ( \30315 , \30312 , \30314 );
not \U$29939 ( \30316 , \30132 );
not \U$29940 ( \30317 , \30140 );
or \U$29941 ( \30318 , \30316 , \30317 );
or \U$29942 ( \30319 , \30132 , \30140 );
nand \U$29943 ( \30320 , \30318 , \30319 );
not \U$29944 ( \30321 , \30320 );
xor \U$29945 ( \30322 , \30106 , \30113 );
xor \U$29946 ( \30323 , \30322 , \30121 );
not \U$29947 ( \30324 , \30323 );
or \U$29948 ( \30325 , \30321 , \30324 );
or \U$29949 ( \30326 , \30323 , \30320 );
xor \U$29950 ( \30327 , \30151 , \30158 );
xor \U$29951 ( \30328 , \30327 , \30166 );
nand \U$29952 ( \30329 , \30326 , \30328 );
nand \U$29953 ( \30330 , \30325 , \30329 );
and \U$29954 ( \30331 , \30315 , \30330 );
and \U$29955 ( \30332 , \30312 , \30314 );
or \U$29956 ( \30333 , \30331 , \30332 );
and \U$29957 ( \30334 , \30236 , \30333 );
and \U$29958 ( \30335 , \30233 , \30235 );
or \U$29959 ( \30336 , \30334 , \30335 );
nand \U$29960 ( \30337 , \30222 , \30336 );
or \U$29961 ( \30338 , \30215 , \30337 );
xnor \U$29962 ( \30339 , \30337 , \30215 );
not \U$29963 ( \30340 , \30336 );
not \U$29964 ( \30341 , \30221 );
or \U$29965 ( \30342 , \30340 , \30341 );
or \U$29966 ( \30343 , \30221 , \30336 );
nand \U$29967 ( \30344 , \30342 , \30343 );
xor \U$29968 ( \30345 , \30233 , \30235 );
xor \U$29969 ( \30346 , \30345 , \30333 );
not \U$29970 ( \30347 , \30346 );
not \U$29971 ( \30348 , \30171 );
not \U$29972 ( \30349 , \30190 );
or \U$29973 ( \30350 , \30348 , \30349 );
or \U$29974 ( \30351 , \30190 , \30171 );
nand \U$29975 ( \30352 , \30350 , \30351 );
not \U$29976 ( \30353 , \30352 );
not \U$29977 ( \30354 , \30099 );
and \U$29978 ( \30355 , \30353 , \30354 );
and \U$29979 ( \30356 , \30352 , \30099 );
nor \U$29980 ( \30357 , \30355 , \30356 );
nor \U$29981 ( \30358 , \30347 , \30357 );
and \U$29982 ( \30359 , \30344 , \30358 );
xor \U$29983 ( \30360 , \30358 , \30344 );
not \U$29984 ( \30361 , \30346 );
not \U$29985 ( \30362 , \30357 );
and \U$29986 ( \30363 , \30361 , \30362 );
and \U$29987 ( \30364 , \30346 , \30357 );
nor \U$29988 ( \30365 , \30363 , \30364 );
xor \U$29989 ( \30366 , \30312 , \30314 );
xor \U$29990 ( \30367 , \30366 , \30330 );
xor \U$29991 ( \30368 , \30228 , \30232 );
and \U$29992 ( \30369 , \30367 , \30368 );
not \U$29993 ( \30370 , \30367 );
not \U$29994 ( \30371 , \30368 );
and \U$29995 ( \30372 , \30370 , \30371 );
xnor \U$29996 ( \30373 , \30308 , \30298 );
not \U$29997 ( \30374 , \30373 );
not \U$29998 ( \30375 , \30290 );
and \U$29999 ( \30376 , \30374 , \30375 );
and \U$30000 ( \30377 , \30373 , \30290 );
nor \U$30001 ( \30378 , \30376 , \30377 );
not \U$30002 ( \30379 , \30378 );
and \U$30003 ( \30380 , \14059 , RIae76f28_65);
and \U$30004 ( \30381 , RIae76e38_63, \14057 );
nor \U$30005 ( \30382 , \30380 , \30381 );
and \U$30006 ( \30383 , \30382 , \14063 );
not \U$30007 ( \30384 , \30382 );
and \U$30008 ( \30385 , \30384 , \13502 );
nor \U$30009 ( \30386 , \30383 , \30385 );
not \U$30010 ( \30387 , \30386 );
and \U$30011 ( \30388 , \15726 , RIae77180_70);
and \U$30012 ( \30389 , RIae7aab0_192, RIae77018_67);
nor \U$30013 ( \30390 , \30388 , \30389 );
and \U$30014 ( \30391 , \30390 , RIae7aa38_191);
not \U$30015 ( \30392 , \30390 );
and \U$30016 ( \30393 , \30392 , \14959 );
nor \U$30017 ( \30394 , \30391 , \30393 );
not \U$30018 ( \30395 , \30394 );
and \U$30019 ( \30396 , \30387 , \30395 );
and \U$30020 ( \30397 , \30386 , \30394 );
and \U$30021 ( \30398 , \14964 , RIae76d48_61);
and \U$30022 ( \30399 , RIae76c58_59, \14962 );
nor \U$30023 ( \30400 , \30398 , \30399 );
and \U$30024 ( \30401 , \30400 , \14462 );
not \U$30025 ( \30402 , \30400 );
and \U$30026 ( \30403 , \30402 , \14463 );
nor \U$30027 ( \30404 , \30401 , \30403 );
nor \U$30028 ( \30405 , \30397 , \30404 );
nor \U$30029 ( \30406 , \30396 , \30405 );
not \U$30030 ( \30407 , \30406 );
and \U$30031 ( \30408 , \30379 , \30407 );
and \U$30032 ( \30409 , \30378 , \30406 );
and \U$30033 ( \30410 , \12180 , RIae77a68_89);
and \U$30034 ( \30411 , RIae77978_87, \12178 );
nor \U$30035 ( \30412 , \30410 , \30411 );
and \U$30036 ( \30413 , \30412 , \11827 );
not \U$30037 ( \30414 , \30412 );
and \U$30038 ( \30415 , \30414 , \12184 );
nor \U$30039 ( \30416 , \30413 , \30415 );
and \U$30040 ( \30417 , \13059 , RIae77798_83);
and \U$30041 ( \30418 , RIae77888_85, \13057 );
nor \U$30042 ( \30419 , \30417 , \30418 );
and \U$30043 ( \30420 , \30419 , \12718 );
not \U$30044 ( \30421 , \30419 );
and \U$30045 ( \30422 , \30421 , \13063 );
nor \U$30046 ( \30423 , \30420 , \30422 );
or \U$30047 ( \30424 , \30416 , \30423 );
and \U$30048 ( \30425 , \30423 , \30416 );
and \U$30049 ( \30426 , \11470 , RIae77720_82);
and \U$30050 ( \30427 , RIae773d8_75, \11468 );
nor \U$30051 ( \30428 , \30426 , \30427 );
and \U$30052 ( \30429 , \30428 , \11474 );
not \U$30053 ( \30430 , \30428 );
and \U$30054 ( \30431 , \30430 , \10936 );
nor \U$30055 ( \30432 , \30429 , \30431 );
nor \U$30056 ( \30433 , \30425 , \30432 );
not \U$30057 ( \30434 , \30433 );
nand \U$30058 ( \30435 , \30424 , \30434 );
not \U$30059 ( \30436 , \30435 );
nor \U$30060 ( \30437 , \30409 , \30436 );
nor \U$30061 ( \30438 , \30408 , \30437 );
xor \U$30062 ( \30439 , \30243 , \30250 );
xor \U$30063 ( \30440 , \30439 , \30258 );
not \U$30064 ( \30441 , \30440 );
not \U$30065 ( \30442 , \9273 );
not \U$30066 ( \30443 , \30268 );
not \U$30067 ( \30444 , \30279 );
or \U$30068 ( \30445 , \30443 , \30444 );
or \U$30069 ( \30446 , \30279 , \30268 );
nand \U$30070 ( \30447 , \30445 , \30446 );
not \U$30071 ( \30448 , \30447 );
or \U$30072 ( \30449 , \30442 , \30448 );
or \U$30073 ( \30450 , \30447 , \9273 );
nand \U$30074 ( \30451 , \30449 , \30450 );
nand \U$30075 ( \30452 , \30441 , \30451 );
xor \U$30076 ( \30453 , \30438 , \30452 );
xnor \U$30077 ( \30454 , \30328 , \30323 );
not \U$30078 ( \30455 , \30454 );
not \U$30079 ( \30456 , \30320 );
and \U$30080 ( \30457 , \30455 , \30456 );
and \U$30081 ( \30458 , \30454 , \30320 );
nor \U$30082 ( \30459 , \30457 , \30458 );
and \U$30083 ( \30460 , \30453 , \30459 );
and \U$30084 ( \30461 , \30438 , \30452 );
or \U$30085 ( \30462 , \30460 , \30461 );
nor \U$30086 ( \30463 , \30372 , \30462 );
nor \U$30087 ( \30464 , \30369 , \30463 );
or \U$30088 ( \30465 , \30365 , \30464 );
xnor \U$30089 ( \30466 , \30464 , \30365 );
and \U$30090 ( \30467 , \14964 , RIae76f28_65);
and \U$30091 ( \30468 , RIae76e38_63, \14962 );
nor \U$30092 ( \30469 , \30467 , \30468 );
and \U$30093 ( \30470 , \30469 , \14462 );
not \U$30094 ( \30471 , \30469 );
and \U$30095 ( \30472 , \30471 , \14463 );
nor \U$30096 ( \30473 , \30470 , \30472 );
and \U$30097 ( \30474 , \15726 , RIae76d48_61);
and \U$30098 ( \30475 , RIae7aab0_192, RIae76c58_59);
nor \U$30099 ( \30476 , \30474 , \30475 );
and \U$30100 ( \30477 , \30476 , RIae7aa38_191);
not \U$30101 ( \30478 , \30476 );
and \U$30102 ( \30479 , \30478 , \14959 );
nor \U$30103 ( \30480 , \30477 , \30479 );
xor \U$30104 ( \30481 , \30473 , \30480 );
and \U$30105 ( \30482 , \14059 , RIae77798_83);
and \U$30106 ( \30483 , RIae77888_85, \14057 );
nor \U$30107 ( \30484 , \30482 , \30483 );
and \U$30108 ( \30485 , \30484 , \14063 );
not \U$30109 ( \30486 , \30484 );
and \U$30110 ( \30487 , \30486 , \13502 );
nor \U$30111 ( \30488 , \30485 , \30487 );
and \U$30112 ( \30489 , \30481 , \30488 );
and \U$30113 ( \30490 , \30473 , \30480 );
or \U$30114 ( \30491 , \30489 , \30490 );
not \U$30115 ( \30492 , \30491 );
and \U$30116 ( \30493 , \11470 , RIae774c8_77);
and \U$30117 ( \30494 , RIae77720_82, \11468 );
nor \U$30118 ( \30495 , \30493 , \30494 );
and \U$30119 ( \30496 , \30495 , \11474 );
not \U$30120 ( \30497 , \30495 );
and \U$30121 ( \30498 , \30497 , \10936 );
nor \U$30122 ( \30499 , \30496 , \30498 );
not \U$30123 ( \30500 , \30499 );
and \U$30124 ( \30501 , \30492 , \30500 );
and \U$30125 ( \30502 , \30491 , \30499 );
and \U$30126 ( \30503 , \12180 , RIae77720_82);
and \U$30127 ( \30504 , RIae773d8_75, \12178 );
nor \U$30128 ( \30505 , \30503 , \30504 );
and \U$30129 ( \30506 , \30505 , \11827 );
not \U$30130 ( \30507 , \30505 );
and \U$30131 ( \30508 , \30507 , \12184 );
nor \U$30132 ( \30509 , \30506 , \30508 );
and \U$30133 ( \30510 , \13059 , RIae77a68_89);
and \U$30134 ( \30511 , RIae77978_87, \13057 );
nor \U$30135 ( \30512 , \30510 , \30511 );
and \U$30136 ( \30513 , \30512 , \12718 );
not \U$30137 ( \30514 , \30512 );
and \U$30138 ( \30515 , \30514 , \13063 );
nor \U$30139 ( \30516 , \30513 , \30515 );
or \U$30140 ( \30517 , \30509 , \30516 );
and \U$30141 ( \30518 , \30516 , \30509 );
and \U$30142 ( \30519 , \11470 , RIae775b8_79);
and \U$30143 ( \30520 , RIae774c8_77, \11468 );
nor \U$30144 ( \30521 , \30519 , \30520 );
and \U$30145 ( \30522 , \30521 , \11474 );
not \U$30146 ( \30523 , \30521 );
and \U$30147 ( \30524 , \30523 , \10936 );
nor \U$30148 ( \30525 , \30522 , \30524 );
nor \U$30149 ( \30526 , \30518 , \30525 );
not \U$30150 ( \30527 , \30526 );
nand \U$30151 ( \30528 , \30517 , \30527 );
not \U$30152 ( \30529 , \30528 );
nor \U$30153 ( \30530 , \30502 , \30529 );
nor \U$30154 ( \30531 , \30501 , \30530 );
not \U$30155 ( \30532 , \30531 );
nand \U$30156 ( \30533 , RIae775b8_79, \10546 );
and \U$30157 ( \30534 , \30533 , \10421 );
not \U$30158 ( \30535 , \30533 );
and \U$30159 ( \30536 , \30535 , \10118 );
nor \U$30160 ( \30537 , \30534 , \30536 );
and \U$30161 ( \30538 , \13059 , RIae77978_87);
and \U$30162 ( \30539 , RIae77798_83, \13057 );
nor \U$30163 ( \30540 , \30538 , \30539 );
and \U$30164 ( \30541 , \30540 , \13063 );
not \U$30165 ( \30542 , \30540 );
and \U$30166 ( \30543 , \30542 , \12718 );
nor \U$30167 ( \30544 , \30541 , \30543 );
and \U$30168 ( \30545 , \12180 , RIae773d8_75);
and \U$30169 ( \30546 , RIae77a68_89, \12178 );
nor \U$30170 ( \30547 , \30545 , \30546 );
and \U$30171 ( \30548 , \30547 , \12184 );
not \U$30172 ( \30549 , \30547 );
and \U$30173 ( \30550 , \30549 , \11827 );
nor \U$30174 ( \30551 , \30548 , \30550 );
xor \U$30175 ( \30552 , \30544 , \30551 );
and \U$30176 ( \30553 , \14059 , RIae77888_85);
and \U$30177 ( \30554 , RIae76f28_65, \14057 );
nor \U$30178 ( \30555 , \30553 , \30554 );
and \U$30179 ( \30556 , \30555 , \13502 );
not \U$30180 ( \30557 , \30555 );
and \U$30181 ( \30558 , \30557 , \14063 );
nor \U$30182 ( \30559 , \30556 , \30558 );
xor \U$30183 ( \30560 , \30552 , \30559 );
and \U$30184 ( \30561 , \30537 , \30560 );
and \U$30185 ( \30562 , \15726 , RIae76c58_59);
and \U$30186 ( \30563 , RIae7aab0_192, RIae77180_70);
nor \U$30187 ( \30564 , \30562 , \30563 );
and \U$30188 ( \30565 , \30564 , \14959 );
not \U$30189 ( \30566 , \30564 );
and \U$30190 ( \30567 , \30566 , RIae7aa38_191);
nor \U$30191 ( \30568 , \30565 , \30567 );
xor \U$30192 ( \30569 , \30568 , \10118 );
and \U$30193 ( \30570 , \14964 , RIae76e38_63);
and \U$30194 ( \30571 , RIae76d48_61, \14962 );
nor \U$30195 ( \30572 , \30570 , \30571 );
and \U$30196 ( \30573 , \30572 , \14463 );
not \U$30197 ( \30574 , \30572 );
and \U$30198 ( \30575 , \30574 , \14462 );
nor \U$30199 ( \30576 , \30573 , \30575 );
xor \U$30200 ( \30577 , \30569 , \30576 );
xor \U$30201 ( \30578 , \30544 , \30551 );
xor \U$30202 ( \30579 , \30578 , \30559 );
and \U$30203 ( \30580 , \30577 , \30579 );
and \U$30204 ( \30581 , \30537 , \30577 );
or \U$30205 ( \30582 , \30561 , \30580 , \30581 );
not \U$30206 ( \30583 , \30582 );
or \U$30207 ( \30584 , \30532 , \30583 );
or \U$30208 ( \30585 , \30582 , \30531 );
nand \U$30209 ( \30586 , \30584 , \30585 );
not \U$30210 ( \30587 , \30586 );
xor \U$30211 ( \30588 , \30416 , \30423 );
not \U$30212 ( \30589 , \30588 );
not \U$30213 ( \30590 , \30432 );
and \U$30214 ( \30591 , \30589 , \30590 );
and \U$30215 ( \30592 , \30588 , \30432 );
nor \U$30216 ( \30593 , \30591 , \30592 );
not \U$30217 ( \30594 , \30593 );
and \U$30218 ( \30595 , \30587 , \30594 );
and \U$30219 ( \30596 , \30586 , \30593 );
nor \U$30220 ( \30597 , \30595 , \30596 );
not \U$30221 ( \30598 , \30386 );
xor \U$30222 ( \30599 , \30394 , \30404 );
not \U$30223 ( \30600 , \30599 );
or \U$30224 ( \30601 , \30598 , \30600 );
or \U$30225 ( \30602 , \30599 , \30386 );
nand \U$30226 ( \30603 , \30601 , \30602 );
xor \U$30227 ( \30604 , \30568 , \10118 );
and \U$30228 ( \30605 , \30604 , \30576 );
and \U$30229 ( \30606 , \30568 , \10118 );
or \U$30230 ( \30607 , \30605 , \30606 );
and \U$30231 ( \30608 , \10548 , RIae775b8_79);
and \U$30232 ( \30609 , RIae774c8_77, \10546 );
nor \U$30233 ( \30610 , \30608 , \30609 );
and \U$30234 ( \30611 , \30610 , \10421 );
not \U$30235 ( \30612 , \30610 );
and \U$30236 ( \30613 , \30612 , \10118 );
nor \U$30237 ( \30614 , \30611 , \30613 );
xor \U$30238 ( \30615 , \30607 , \30614 );
xor \U$30239 ( \30616 , \30544 , \30551 );
and \U$30240 ( \30617 , \30616 , \30559 );
and \U$30241 ( \30618 , \30544 , \30551 );
or \U$30242 ( \30619 , \30617 , \30618 );
xor \U$30243 ( \30620 , \30615 , \30619 );
xor \U$30244 ( \30621 , \30603 , \30620 );
not \U$30245 ( \30622 , \30621 );
or \U$30246 ( \30623 , \30597 , \30622 );
not \U$30247 ( \30624 , \30622 );
not \U$30248 ( \30625 , \30597 );
or \U$30249 ( \30626 , \30624 , \30625 );
not \U$30250 ( \30627 , \30499 );
not \U$30251 ( \30628 , \30528 );
not \U$30252 ( \30629 , \30491 );
or \U$30253 ( \30630 , \30628 , \30629 );
or \U$30254 ( \30631 , \30491 , \30528 );
nand \U$30255 ( \30632 , \30630 , \30631 );
not \U$30256 ( \30633 , \30632 );
or \U$30257 ( \30634 , \30627 , \30633 );
or \U$30258 ( \30635 , \30632 , \30499 );
nand \U$30259 ( \30636 , \30634 , \30635 );
xor \U$30260 ( \30637 , \30509 , \30516 );
not \U$30261 ( \30638 , \30637 );
not \U$30262 ( \30639 , \30525 );
and \U$30263 ( \30640 , \30638 , \30639 );
and \U$30264 ( \30641 , \30637 , \30525 );
nor \U$30265 ( \30642 , \30640 , \30641 );
and \U$30266 ( \30643 , \15726 , RIae76e38_63);
and \U$30267 ( \30644 , RIae7aab0_192, RIae76d48_61);
nor \U$30268 ( \30645 , \30643 , \30644 );
and \U$30269 ( \30646 , \30645 , \14959 );
not \U$30270 ( \30647 , \30645 );
and \U$30271 ( \30648 , \30647 , RIae7aa38_191);
nor \U$30272 ( \30649 , \30646 , \30648 );
and \U$30273 ( \30650 , \30649 , \11474 );
not \U$30274 ( \30651 , \30649 );
not \U$30275 ( \30652 , \11474 );
and \U$30276 ( \30653 , \30651 , \30652 );
and \U$30277 ( \30654 , \14964 , RIae77888_85);
and \U$30278 ( \30655 , RIae76f28_65, \14962 );
nor \U$30279 ( \30656 , \30654 , \30655 );
and \U$30280 ( \30657 , \30656 , \14462 );
not \U$30281 ( \30658 , \30656 );
and \U$30282 ( \30659 , \30658 , \14463 );
nor \U$30283 ( \30660 , \30657 , \30659 );
nor \U$30284 ( \30661 , \30653 , \30660 );
nor \U$30285 ( \30662 , \30650 , \30661 );
or \U$30286 ( \30663 , \30642 , \30662 );
not \U$30287 ( \30664 , \30662 );
not \U$30288 ( \30665 , \30642 );
or \U$30289 ( \30666 , \30664 , \30665 );
and \U$30290 ( \30667 , \13059 , RIae773d8_75);
and \U$30291 ( \30668 , RIae77a68_89, \13057 );
nor \U$30292 ( \30669 , \30667 , \30668 );
and \U$30293 ( \30670 , \30669 , \12718 );
not \U$30294 ( \30671 , \30669 );
and \U$30295 ( \30672 , \30671 , \13063 );
nor \U$30296 ( \30673 , \30670 , \30672 );
and \U$30297 ( \30674 , \14059 , RIae77978_87);
and \U$30298 ( \30675 , RIae77798_83, \14057 );
nor \U$30299 ( \30676 , \30674 , \30675 );
and \U$30300 ( \30677 , \30676 , \14063 );
not \U$30301 ( \30678 , \30676 );
and \U$30302 ( \30679 , \30678 , \13502 );
nor \U$30303 ( \30680 , \30677 , \30679 );
xor \U$30304 ( \30681 , \30673 , \30680 );
and \U$30305 ( \30682 , \12180 , RIae774c8_77);
and \U$30306 ( \30683 , RIae77720_82, \12178 );
nor \U$30307 ( \30684 , \30682 , \30683 );
and \U$30308 ( \30685 , \30684 , \11827 );
not \U$30309 ( \30686 , \30684 );
and \U$30310 ( \30687 , \30686 , \12184 );
nor \U$30311 ( \30688 , \30685 , \30687 );
and \U$30312 ( \30689 , \30681 , \30688 );
and \U$30313 ( \30690 , \30673 , \30680 );
nor \U$30314 ( \30691 , \30689 , \30690 );
nand \U$30315 ( \30692 , \30666 , \30691 );
nand \U$30316 ( \30693 , \30663 , \30692 );
xor \U$30317 ( \30694 , \30636 , \30693 );
xor \U$30318 ( \30695 , \30544 , \30551 );
xor \U$30319 ( \30696 , \30695 , \30559 );
xor \U$30320 ( \30697 , \30537 , \30577 );
xor \U$30321 ( \30698 , \30696 , \30697 );
and \U$30322 ( \30699 , \30694 , \30698 );
and \U$30323 ( \30700 , \30636 , \30693 );
or \U$30324 ( \30701 , \30699 , \30700 );
nand \U$30325 ( \30702 , \30626 , \30701 );
nand \U$30326 ( \30703 , \30623 , \30702 );
not \U$30327 ( \30704 , \30440 );
not \U$30328 ( \30705 , \30451 );
or \U$30329 ( \30706 , \30704 , \30705 );
or \U$30330 ( \30707 , \30451 , \30440 );
nand \U$30331 ( \30708 , \30706 , \30707 );
xor \U$30332 ( \30709 , \30607 , \30614 );
and \U$30333 ( \30710 , \30709 , \30619 );
and \U$30334 ( \30711 , \30607 , \30614 );
or \U$30335 ( \30712 , \30710 , \30711 );
xor \U$30336 ( \30713 , \30708 , \30712 );
not \U$30337 ( \30714 , \30378 );
not \U$30338 ( \30715 , \30435 );
not \U$30339 ( \30716 , \30406 );
or \U$30340 ( \30717 , \30715 , \30716 );
or \U$30341 ( \30718 , \30406 , \30435 );
nand \U$30342 ( \30719 , \30717 , \30718 );
not \U$30343 ( \30720 , \30719 );
or \U$30344 ( \30721 , \30714 , \30720 );
or \U$30345 ( \30722 , \30719 , \30378 );
nand \U$30346 ( \30723 , \30721 , \30722 );
xor \U$30347 ( \30724 , \30713 , \30723 );
and \U$30348 ( \30725 , \30603 , \30620 );
xor \U$30349 ( \30726 , \30724 , \30725 );
or \U$30350 ( \30727 , \30531 , \30593 );
not \U$30351 ( \30728 , \30593 );
not \U$30352 ( \30729 , \30531 );
or \U$30353 ( \30730 , \30728 , \30729 );
nand \U$30354 ( \30731 , \30730 , \30582 );
nand \U$30355 ( \30732 , \30727 , \30731 );
xor \U$30356 ( \30733 , \30726 , \30732 );
and \U$30357 ( \30734 , \30703 , \30733 );
xor \U$30358 ( \30735 , \30733 , \30703 );
and \U$30359 ( \30736 , \14964 , RIae77798_83);
and \U$30360 ( \30737 , RIae77888_85, \14962 );
nor \U$30361 ( \30738 , \30736 , \30737 );
and \U$30362 ( \30739 , \30738 , \14463 );
not \U$30363 ( \30740 , \30738 );
and \U$30364 ( \30741 , \30740 , \14462 );
nor \U$30365 ( \30742 , \30739 , \30741 );
and \U$30366 ( \30743 , \15726 , RIae76f28_65);
and \U$30367 ( \30744 , RIae7aab0_192, RIae76e38_63);
nor \U$30368 ( \30745 , \30743 , \30744 );
and \U$30369 ( \30746 , \30745 , \14959 );
not \U$30370 ( \30747 , \30745 );
and \U$30371 ( \30748 , \30747 , RIae7aa38_191);
nor \U$30372 ( \30749 , \30746 , \30748 );
xor \U$30373 ( \30750 , \30742 , \30749 );
and \U$30374 ( \30751 , \14059 , RIae77a68_89);
and \U$30375 ( \30752 , RIae77978_87, \14057 );
nor \U$30376 ( \30753 , \30751 , \30752 );
and \U$30377 ( \30754 , \30753 , \13502 );
not \U$30378 ( \30755 , \30753 );
and \U$30379 ( \30756 , \30755 , \14063 );
nor \U$30380 ( \30757 , \30754 , \30756 );
and \U$30381 ( \30758 , \30750 , \30757 );
and \U$30382 ( \30759 , \30742 , \30749 );
nor \U$30383 ( \30760 , \30758 , \30759 );
nand \U$30384 ( \30761 , RIae775b8_79, \11468 );
and \U$30385 ( \30762 , \30761 , \11474 );
not \U$30386 ( \30763 , \30761 );
and \U$30387 ( \30764 , \30763 , \10936 );
nor \U$30388 ( \30765 , \30762 , \30764 );
xor \U$30389 ( \30766 , \30760 , \30765 );
xor \U$30390 ( \30767 , \30673 , \30680 );
xor \U$30391 ( \30768 , \30767 , \30688 );
and \U$30392 ( \30769 , \30766 , \30768 );
and \U$30393 ( \30770 , \30760 , \30765 );
or \U$30394 ( \30771 , \30769 , \30770 );
xor \U$30395 ( \30772 , \30473 , \30480 );
xor \U$30396 ( \30773 , \30772 , \30488 );
xor \U$30397 ( \30774 , \30771 , \30773 );
not \U$30398 ( \30775 , \30662 );
not \U$30399 ( \30776 , \30691 );
or \U$30400 ( \30777 , \30775 , \30776 );
or \U$30401 ( \30778 , \30691 , \30662 );
nand \U$30402 ( \30779 , \30777 , \30778 );
not \U$30403 ( \30780 , \30779 );
not \U$30404 ( \30781 , \30642 );
and \U$30405 ( \30782 , \30780 , \30781 );
and \U$30406 ( \30783 , \30779 , \30642 );
nor \U$30407 ( \30784 , \30782 , \30783 );
xor \U$30408 ( \30785 , \30774 , \30784 );
not \U$30409 ( \30786 , \30785 );
and \U$30410 ( \30787 , \15726 , RIae77888_85);
and \U$30411 ( \30788 , RIae7aab0_192, RIae76f28_65);
nor \U$30412 ( \30789 , \30787 , \30788 );
and \U$30413 ( \30790 , \30789 , \14959 );
not \U$30414 ( \30791 , \30789 );
and \U$30415 ( \30792 , \30791 , RIae7aa38_191);
nor \U$30416 ( \30793 , \30790 , \30792 );
xor \U$30417 ( \30794 , \30793 , \11827 );
and \U$30418 ( \30795 , \14964 , RIae77978_87);
and \U$30419 ( \30796 , RIae77798_83, \14962 );
nor \U$30420 ( \30797 , \30795 , \30796 );
and \U$30421 ( \30798 , \30797 , \14463 );
not \U$30422 ( \30799 , \30797 );
and \U$30423 ( \30800 , \30799 , \14462 );
nor \U$30424 ( \30801 , \30798 , \30800 );
and \U$30425 ( \30802 , \30794 , \30801 );
and \U$30426 ( \30803 , \30793 , \11827 );
or \U$30427 ( \30804 , \30802 , \30803 );
and \U$30428 ( \30805 , \13059 , RIae77720_82);
and \U$30429 ( \30806 , RIae773d8_75, \13057 );
nor \U$30430 ( \30807 , \30805 , \30806 );
and \U$30431 ( \30808 , \30807 , \13063 );
not \U$30432 ( \30809 , \30807 );
and \U$30433 ( \30810 , \30809 , \12718 );
nor \U$30434 ( \30811 , \30808 , \30810 );
xor \U$30435 ( \30812 , \30804 , \30811 );
and \U$30436 ( \30813 , \14059 , RIae773d8_75);
and \U$30437 ( \30814 , RIae77a68_89, \14057 );
nor \U$30438 ( \30815 , \30813 , \30814 );
and \U$30439 ( \30816 , \30815 , \13502 );
not \U$30440 ( \30817 , \30815 );
and \U$30441 ( \30818 , \30817 , \14063 );
nor \U$30442 ( \30819 , \30816 , \30818 );
nand \U$30443 ( \30820 , RIae775b8_79, \12178 );
and \U$30444 ( \30821 , \30820 , \12184 );
not \U$30445 ( \30822 , \30820 );
and \U$30446 ( \30823 , \30822 , \11827 );
nor \U$30447 ( \30824 , \30821 , \30823 );
xor \U$30448 ( \30825 , \30819 , \30824 );
and \U$30449 ( \30826 , \13059 , RIae774c8_77);
and \U$30450 ( \30827 , RIae77720_82, \13057 );
nor \U$30451 ( \30828 , \30826 , \30827 );
and \U$30452 ( \30829 , \30828 , \13063 );
not \U$30453 ( \30830 , \30828 );
and \U$30454 ( \30831 , \30830 , \12718 );
nor \U$30455 ( \30832 , \30829 , \30831 );
and \U$30456 ( \30833 , \30825 , \30832 );
and \U$30457 ( \30834 , \30819 , \30824 );
or \U$30458 ( \30835 , \30833 , \30834 );
and \U$30459 ( \30836 , \30812 , \30835 );
and \U$30460 ( \30837 , \30804 , \30811 );
or \U$30461 ( \30838 , \30836 , \30837 );
not \U$30462 ( \30839 , \10936 );
not \U$30463 ( \30840 , \30649 );
not \U$30464 ( \30841 , \30660 );
or \U$30465 ( \30842 , \30840 , \30841 );
or \U$30466 ( \30843 , \30660 , \30649 );
nand \U$30467 ( \30844 , \30842 , \30843 );
not \U$30468 ( \30845 , \30844 );
or \U$30469 ( \30846 , \30839 , \30845 );
or \U$30470 ( \30847 , \30844 , \10936 );
nand \U$30471 ( \30848 , \30846 , \30847 );
xor \U$30472 ( \30849 , \30838 , \30848 );
and \U$30473 ( \30850 , \12180 , RIae775b8_79);
and \U$30474 ( \30851 , RIae774c8_77, \12178 );
nor \U$30475 ( \30852 , \30850 , \30851 );
and \U$30476 ( \30853 , \30852 , \12184 );
not \U$30477 ( \30854 , \30852 );
and \U$30478 ( \30855 , \30854 , \11827 );
nor \U$30479 ( \30856 , \30853 , \30855 );
xor \U$30480 ( \30857 , \30742 , \30749 );
xor \U$30481 ( \30858 , \30857 , \30757 );
and \U$30482 ( \30859 , \30856 , \30858 );
and \U$30483 ( \30860 , \30849 , \30859 );
and \U$30484 ( \30861 , \30838 , \30848 );
or \U$30485 ( \30862 , \30860 , \30861 );
not \U$30486 ( \30863 , \30862 );
and \U$30487 ( \30864 , \30786 , \30863 );
and \U$30488 ( \30865 , \30785 , \30862 );
nor \U$30489 ( \30866 , \30864 , \30865 );
xor \U$30490 ( \30867 , \30760 , \30765 );
xor \U$30491 ( \30868 , \30867 , \30768 );
not \U$30492 ( \30869 , \30868 );
xor \U$30493 ( \30870 , \30838 , \30848 );
xor \U$30494 ( \30871 , \30870 , \30859 );
nand \U$30495 ( \30872 , \30869 , \30871 );
or \U$30496 ( \30873 , \30866 , \30872 );
xnor \U$30497 ( \30874 , \30872 , \30866 );
and \U$30498 ( \30875 , \15726 , RIae77978_87);
and \U$30499 ( \30876 , RIae7aab0_192, RIae77798_83);
nor \U$30500 ( \30877 , \30875 , \30876 );
and \U$30501 ( \30878 , \30877 , \14959 );
not \U$30502 ( \30879 , \30877 );
and \U$30503 ( \30880 , \30879 , RIae7aa38_191);
nor \U$30504 ( \30881 , \30878 , \30880 );
xor \U$30505 ( \30882 , \30881 , \12718 );
and \U$30506 ( \30883 , \14964 , RIae773d8_75);
and \U$30507 ( \30884 , RIae77a68_89, \14962 );
nor \U$30508 ( \30885 , \30883 , \30884 );
and \U$30509 ( \30886 , \30885 , \14463 );
not \U$30510 ( \30887 , \30885 );
and \U$30511 ( \30888 , \30887 , \14462 );
nor \U$30512 ( \30889 , \30886 , \30888 );
xor \U$30513 ( \30890 , \30882 , \30889 );
nand \U$30514 ( \30891 , RIae775b8_79, \13057 );
and \U$30515 ( \30892 , \30891 , \13063 );
not \U$30516 ( \30893 , \30891 );
and \U$30517 ( \30894 , \30893 , \12718 );
nor \U$30518 ( \30895 , \30892 , \30894 );
not \U$30519 ( \30896 , \30895 );
and \U$30520 ( \30897 , \14059 , RIae774c8_77);
and \U$30521 ( \30898 , RIae77720_82, \14057 );
nor \U$30522 ( \30899 , \30897 , \30898 );
and \U$30523 ( \30900 , \30899 , \14063 );
not \U$30524 ( \30901 , \30899 );
and \U$30525 ( \30902 , \30901 , \13502 );
nor \U$30526 ( \30903 , \30900 , \30902 );
not \U$30527 ( \30904 , \30903 );
or \U$30528 ( \30905 , \30896 , \30904 );
or \U$30529 ( \30906 , \30903 , \30895 );
nand \U$30530 ( \30907 , \30905 , \30906 );
and \U$30531 ( \30908 , \30890 , \30907 );
not \U$30532 ( \30909 , \30890 );
not \U$30533 ( \30910 , \30907 );
and \U$30534 ( \30911 , \30909 , \30910 );
and \U$30535 ( \30912 , \14059 , RIae775b8_79);
and \U$30536 ( \30913 , RIae774c8_77, \14057 );
nor \U$30537 ( \30914 , \30912 , \30913 );
and \U$30538 ( \30915 , \30914 , \14063 );
not \U$30539 ( \30916 , \30914 );
and \U$30540 ( \30917 , \30916 , \13502 );
nor \U$30541 ( \30918 , \30915 , \30917 );
and \U$30542 ( \30919 , \15726 , RIae77a68_89);
and \U$30543 ( \30920 , RIae7aab0_192, RIae77978_87);
nor \U$30544 ( \30921 , \30919 , \30920 );
and \U$30545 ( \30922 , \30921 , RIae7aa38_191);
not \U$30546 ( \30923 , \30921 );
and \U$30547 ( \30924 , \30923 , \14959 );
nor \U$30548 ( \30925 , \30922 , \30924 );
xor \U$30549 ( \30926 , \30918 , \30925 );
and \U$30550 ( \30927 , \14964 , RIae77720_82);
and \U$30551 ( \30928 , RIae773d8_75, \14962 );
nor \U$30552 ( \30929 , \30927 , \30928 );
and \U$30553 ( \30930 , \30929 , \14462 );
not \U$30554 ( \30931 , \30929 );
and \U$30555 ( \30932 , \30931 , \14463 );
nor \U$30556 ( \30933 , \30930 , \30932 );
and \U$30557 ( \30934 , \30926 , \30933 );
and \U$30558 ( \30935 , \30918 , \30925 );
or \U$30559 ( \30936 , \30934 , \30935 );
nor \U$30560 ( \30937 , \30911 , \30936 );
nor \U$30561 ( \30938 , \30908 , \30937 );
and \U$30562 ( \30939 , \13059 , RIae775b8_79);
and \U$30563 ( \30940 , RIae774c8_77, \13057 );
nor \U$30564 ( \30941 , \30939 , \30940 );
and \U$30565 ( \30942 , \30941 , \12718 );
not \U$30566 ( \30943 , \30941 );
and \U$30567 ( \30944 , \30943 , \13063 );
nor \U$30568 ( \30945 , \30942 , \30944 );
not \U$30569 ( \30946 , \30945 );
not \U$30570 ( \30947 , \30903 );
nand \U$30571 ( \30948 , \30947 , \30895 );
not \U$30572 ( \30949 , \30948 );
xor \U$30573 ( \30950 , \30881 , \12718 );
and \U$30574 ( \30951 , \30950 , \30889 );
and \U$30575 ( \30952 , \30881 , \12718 );
or \U$30576 ( \30953 , \30951 , \30952 );
not \U$30577 ( \30954 , \30953 );
or \U$30578 ( \30955 , \30949 , \30954 );
or \U$30579 ( \30956 , \30953 , \30948 );
nand \U$30580 ( \30957 , \30955 , \30956 );
not \U$30581 ( \30958 , \30957 );
or \U$30582 ( \30959 , \30946 , \30958 );
or \U$30583 ( \30960 , \30957 , \30945 );
nand \U$30584 ( \30961 , \30959 , \30960 );
not \U$30585 ( \30962 , \30961 );
and \U$30586 ( \30963 , \15726 , RIae77798_83);
and \U$30587 ( \30964 , RIae7aab0_192, RIae77888_85);
nor \U$30588 ( \30965 , \30963 , \30964 );
and \U$30589 ( \30966 , \30965 , RIae7aa38_191);
not \U$30590 ( \30967 , \30965 );
and \U$30591 ( \30968 , \30967 , \14959 );
nor \U$30592 ( \30969 , \30966 , \30968 );
not \U$30593 ( \30970 , \30969 );
and \U$30594 ( \30971 , \14964 , RIae77a68_89);
and \U$30595 ( \30972 , RIae77978_87, \14962 );
nor \U$30596 ( \30973 , \30971 , \30972 );
and \U$30597 ( \30974 , \30973 , \14463 );
not \U$30598 ( \30975 , \30973 );
and \U$30599 ( \30976 , \30975 , \14462 );
nor \U$30600 ( \30977 , \30974 , \30976 );
not \U$30601 ( \30978 , \30977 );
or \U$30602 ( \30979 , \30970 , \30978 );
or \U$30603 ( \30980 , \30977 , \30969 );
nand \U$30604 ( \30981 , \30979 , \30980 );
not \U$30605 ( \30982 , \30981 );
and \U$30606 ( \30983 , \14059 , RIae77720_82);
and \U$30607 ( \30984 , RIae773d8_75, \14057 );
nor \U$30608 ( \30985 , \30983 , \30984 );
and \U$30609 ( \30986 , \30985 , \14063 );
not \U$30610 ( \30987 , \30985 );
and \U$30611 ( \30988 , \30987 , \13502 );
nor \U$30612 ( \30989 , \30986 , \30988 );
not \U$30613 ( \30990 , \30989 );
and \U$30614 ( \30991 , \30982 , \30990 );
and \U$30615 ( \30992 , \30981 , \30989 );
nor \U$30616 ( \30993 , \30991 , \30992 );
not \U$30617 ( \30994 , \30993 );
and \U$30618 ( \30995 , \30962 , \30994 );
and \U$30619 ( \30996 , \30961 , \30993 );
nor \U$30620 ( \30997 , \30995 , \30996 );
xor \U$30621 ( \30998 , \30938 , \30997 );
and \U$30622 ( \30999 , \14964 , RIae775b8_79);
and \U$30623 ( \31000 , RIae774c8_77, \14962 );
nor \U$30624 ( \31001 , \30999 , \31000 );
and \U$30625 ( \31002 , \31001 , \14463 );
not \U$30626 ( \31003 , \31001 );
and \U$30627 ( \31004 , \31003 , \14462 );
nor \U$30628 ( \31005 , \31002 , \31004 );
not \U$30629 ( \31006 , \31005 );
and \U$30630 ( \31007 , \15726 , RIae77720_82);
and \U$30631 ( \31008 , RIae7aab0_192, RIae773d8_75);
nor \U$30632 ( \31009 , \31007 , \31008 );
and \U$30633 ( \31010 , \31009 , RIae7aa38_191);
not \U$30634 ( \31011 , \31009 );
and \U$30635 ( \31012 , \31011 , \14959 );
nor \U$30636 ( \31013 , \31010 , \31012 );
nor \U$30637 ( \31014 , \31006 , \31013 );
nand \U$30638 ( \31015 , RIae775b8_79, \14057 );
and \U$30639 ( \31016 , \31015 , \14063 );
not \U$30640 ( \31017 , \31015 );
and \U$30641 ( \31018 , \31017 , \13502 );
nor \U$30642 ( \31019 , \31016 , \31018 );
not \U$30643 ( \31020 , \31019 );
and \U$30644 ( \31021 , \15726 , RIae773d8_75);
and \U$30645 ( \31022 , RIae7aab0_192, RIae77a68_89);
nor \U$30646 ( \31023 , \31021 , \31022 );
and \U$30647 ( \31024 , \31023 , \14959 );
not \U$30648 ( \31025 , \31023 );
and \U$30649 ( \31026 , \31025 , RIae7aa38_191);
nor \U$30650 ( \31027 , \31024 , \31026 );
xor \U$30651 ( \31028 , \31027 , \14063 );
and \U$30652 ( \31029 , \14964 , RIae774c8_77);
and \U$30653 ( \31030 , RIae77720_82, \14962 );
nor \U$30654 ( \31031 , \31029 , \31030 );
and \U$30655 ( \31032 , \31031 , \14463 );
not \U$30656 ( \31033 , \31031 );
and \U$30657 ( \31034 , \31033 , \14462 );
nor \U$30658 ( \31035 , \31032 , \31034 );
xor \U$30659 ( \31036 , \31028 , \31035 );
not \U$30660 ( \31037 , \31036 );
or \U$30661 ( \31038 , \31020 , \31037 );
or \U$30662 ( \31039 , \31036 , \31019 );
nand \U$30663 ( \31040 , \31038 , \31039 );
xor \U$30664 ( \31041 , \31014 , \31040 );
and \U$30665 ( \31042 , \15726 , RIae774c8_77);
and \U$30666 ( \31043 , RIae7aab0_192, RIae77720_82);
nor \U$30667 ( \31044 , \31042 , \31043 );
and \U$30668 ( \31045 , \31044 , \14959 );
not \U$30669 ( \31046 , \31044 );
and \U$30670 ( \31047 , \31046 , RIae7aa38_191);
nor \U$30671 ( \31048 , \31045 , \31047 );
nand \U$30672 ( \31049 , \14462 , \31048 );
not \U$30673 ( \31050 , \31005 );
not \U$30674 ( \31051 , \31013 );
and \U$30675 ( \31052 , \31050 , \31051 );
and \U$30676 ( \31053 , \31005 , \31013 );
nor \U$30677 ( \31054 , \31052 , \31053 );
xnor \U$30678 ( \31055 , \31049 , \31054 );
nand \U$30679 ( \31056 , RIae775b8_79, \14962 );
and \U$30680 ( \31057 , \31056 , \14463 );
not \U$30681 ( \31058 , \31056 );
and \U$30682 ( \31059 , \31058 , \14462 );
nor \U$30683 ( \31060 , \31057 , \31059 );
and \U$30684 ( \31061 , \31048 , \14462 );
not \U$30685 ( \31062 , \31048 );
and \U$30686 ( \31063 , \31062 , \14463 );
nor \U$30687 ( \31064 , \31061 , \31063 );
xor \U$30688 ( \31065 , \31060 , \31064 );
nand \U$30689 ( \31066 , RIae775b8_79, RIae7aab0_192);
and \U$30690 ( \31067 , \31066 , RIae7aa38_191);
and \U$30691 ( \31068 , \15726 , RIae775b8_79);
and \U$30692 ( \31069 , RIae7aab0_192, RIae774c8_77);
nor \U$30693 ( \31070 , \31068 , \31069 );
and \U$30694 ( \31071 , \31070 , \14959 );
not \U$30695 ( \31072 , \31070 );
and \U$30696 ( \31073 , \31072 , RIae7aa38_191);
nor \U$30697 ( \31074 , \31071 , \31073 );
and \U$30698 ( \31075 , \31067 , \31074 );
and \U$30699 ( \31076 , \31065 , \31075 );
and \U$30700 ( \31077 , \31060 , \31064 );
nor \U$30701 ( \31078 , \31076 , \31077 );
or \U$30702 ( \31079 , \31055 , \31078 );
or \U$30703 ( \31080 , \31049 , \31054 );
nand \U$30704 ( \31081 , \31079 , \31080 );
and \U$30705 ( \31082 , \31041 , \31081 );
and \U$30706 ( \31083 , \31014 , \31040 );
nor \U$30707 ( \31084 , \31082 , \31083 );
not \U$30708 ( \31085 , \31019 );
nand \U$30709 ( \31086 , \31085 , \31036 );
xor \U$30710 ( \31087 , \30918 , \30925 );
xor \U$30711 ( \31088 , \31087 , \30933 );
not \U$30712 ( \31089 , \31088 );
xor \U$30713 ( \31090 , \31027 , \14063 );
and \U$30714 ( \31091 , \31090 , \31035 );
and \U$30715 ( \31092 , \31027 , \14063 );
or \U$30716 ( \31093 , \31091 , \31092 );
not \U$30717 ( \31094 , \31093 );
and \U$30718 ( \31095 , \31089 , \31094 );
and \U$30719 ( \31096 , \31088 , \31093 );
nor \U$30720 ( \31097 , \31095 , \31096 );
xnor \U$30721 ( \31098 , \31086 , \31097 );
or \U$30722 ( \31099 , \31084 , \31098 );
or \U$30723 ( \31100 , \31086 , \31097 );
nand \U$30724 ( \31101 , \31099 , \31100 );
not \U$30725 ( \31102 , \31093 );
nor \U$30726 ( \31103 , \31102 , \31088 );
not \U$30727 ( \31104 , \30907 );
not \U$30728 ( \31105 , \30890 );
not \U$30729 ( \31106 , \30936 );
and \U$30730 ( \31107 , \31105 , \31106 );
and \U$30731 ( \31108 , \30890 , \30936 );
nor \U$30732 ( \31109 , \31107 , \31108 );
not \U$30733 ( \31110 , \31109 );
or \U$30734 ( \31111 , \31104 , \31110 );
or \U$30735 ( \31112 , \31109 , \30907 );
nand \U$30736 ( \31113 , \31111 , \31112 );
xor \U$30737 ( \31114 , \31103 , \31113 );
and \U$30738 ( \31115 , \31101 , \31114 );
and \U$30739 ( \31116 , \31103 , \31113 );
nor \U$30740 ( \31117 , \31115 , \31116 );
and \U$30741 ( \31118 , \30998 , \31117 );
and \U$30742 ( \31119 , \30938 , \30997 );
nor \U$30743 ( \31120 , \31118 , \31119 );
not \U$30744 ( \31121 , \30961 );
nor \U$30745 ( \31122 , \31121 , \30993 );
not \U$30746 ( \31123 , \30948 );
not \U$30747 ( \31124 , \30945 );
and \U$30748 ( \31125 , \31123 , \31124 );
and \U$30749 ( \31126 , \30948 , \30945 );
not \U$30750 ( \31127 , \30953 );
nor \U$30751 ( \31128 , \31126 , \31127 );
nor \U$30752 ( \31129 , \31125 , \31128 );
not \U$30753 ( \31130 , \31129 );
xor \U$30754 ( \31131 , \30819 , \30824 );
xor \U$30755 ( \31132 , \31131 , \30832 );
or \U$30756 ( \31133 , \30989 , \30969 );
not \U$30757 ( \31134 , \30969 );
not \U$30758 ( \31135 , \30989 );
or \U$30759 ( \31136 , \31134 , \31135 );
nand \U$30760 ( \31137 , \31136 , \30977 );
nand \U$30761 ( \31138 , \31133 , \31137 );
xor \U$30762 ( \31139 , \30793 , \11827 );
xor \U$30763 ( \31140 , \31139 , \30801 );
xor \U$30764 ( \31141 , \31138 , \31140 );
xor \U$30765 ( \31142 , \31132 , \31141 );
not \U$30766 ( \31143 , \31142 );
or \U$30767 ( \31144 , \31130 , \31143 );
or \U$30768 ( \31145 , \31142 , \31129 );
nand \U$30769 ( \31146 , \31144 , \31145 );
xor \U$30770 ( \31147 , \31122 , \31146 );
and \U$30771 ( \31148 , \31120 , \31147 );
and \U$30772 ( \31149 , \31122 , \31146 );
nor \U$30773 ( \31150 , \31148 , \31149 );
not \U$30774 ( \31151 , \31129 );
nand \U$30775 ( \31152 , \31151 , \31142 );
xor \U$30776 ( \31153 , \30804 , \30811 );
xor \U$30777 ( \31154 , \31153 , \30835 );
xor \U$30778 ( \31155 , \30819 , \30824 );
xor \U$30779 ( \31156 , \31155 , \30832 );
and \U$30780 ( \31157 , \31138 , \31156 );
xor \U$30781 ( \31158 , \30819 , \30824 );
xor \U$30782 ( \31159 , \31158 , \30832 );
and \U$30783 ( \31160 , \31140 , \31159 );
and \U$30784 ( \31161 , \31138 , \31140 );
or \U$30785 ( \31162 , \31157 , \31160 , \31161 );
xnor \U$30786 ( \31163 , \31154 , \31162 );
not \U$30787 ( \31164 , \31163 );
xor \U$30788 ( \31165 , \30856 , \30858 );
not \U$30789 ( \31166 , \31165 );
and \U$30790 ( \31167 , \31164 , \31166 );
and \U$30791 ( \31168 , \31163 , \31165 );
nor \U$30792 ( \31169 , \31167 , \31168 );
xnor \U$30793 ( \31170 , \31152 , \31169 );
or \U$30794 ( \31171 , \31150 , \31170 );
or \U$30795 ( \31172 , \31152 , \31169 );
nand \U$30796 ( \31173 , \31171 , \31172 );
not \U$30797 ( \31174 , \31165 );
not \U$30798 ( \31175 , \31154 );
or \U$30799 ( \31176 , \31174 , \31175 );
or \U$30800 ( \31177 , \31154 , \31165 );
nand \U$30801 ( \31178 , \31177 , \31162 );
nand \U$30802 ( \31179 , \31176 , \31178 );
not \U$30803 ( \31180 , \30868 );
not \U$30804 ( \31181 , \30871 );
or \U$30805 ( \31182 , \31180 , \31181 );
or \U$30806 ( \31183 , \30871 , \30868 );
nand \U$30807 ( \31184 , \31182 , \31183 );
xor \U$30808 ( \31185 , \31179 , \31184 );
and \U$30809 ( \31186 , \31173 , \31185 );
and \U$30810 ( \31187 , \31179 , \31184 );
nor \U$30811 ( \31188 , \31186 , \31187 );
or \U$30812 ( \31189 , \30874 , \31188 );
nand \U$30813 ( \31190 , \30873 , \31189 );
not \U$30814 ( \31191 , \30862 );
nor \U$30815 ( \31192 , \31191 , \30785 );
xor \U$30816 ( \31193 , \30771 , \30773 );
and \U$30817 ( \31194 , \31193 , \30784 );
and \U$30818 ( \31195 , \30771 , \30773 );
or \U$30819 ( \31196 , \31194 , \31195 );
not \U$30820 ( \31197 , \31196 );
xor \U$30821 ( \31198 , \30636 , \30693 );
xor \U$30822 ( \31199 , \31198 , \30698 );
not \U$30823 ( \31200 , \31199 );
or \U$30824 ( \31201 , \31197 , \31200 );
or \U$30825 ( \31202 , \31199 , \31196 );
nand \U$30826 ( \31203 , \31201 , \31202 );
xor \U$30827 ( \31204 , \31192 , \31203 );
and \U$30828 ( \31205 , \31190 , \31204 );
and \U$30829 ( \31206 , \31192 , \31203 );
nor \U$30830 ( \31207 , \31205 , \31206 );
not \U$30831 ( \31208 , \31196 );
nand \U$30832 ( \31209 , \31208 , \31199 );
not \U$30833 ( \31210 , \30597 );
not \U$30834 ( \31211 , \30701 );
and \U$30835 ( \31212 , \31210 , \31211 );
and \U$30836 ( \31213 , \30597 , \30701 );
nor \U$30837 ( \31214 , \31212 , \31213 );
not \U$30838 ( \31215 , \31214 );
not \U$30839 ( \31216 , \30621 );
and \U$30840 ( \31217 , \31215 , \31216 );
and \U$30841 ( \31218 , \31214 , \30621 );
nor \U$30842 ( \31219 , \31217 , \31218 );
xnor \U$30843 ( \31220 , \31209 , \31219 );
or \U$30844 ( \31221 , \31207 , \31220 );
or \U$30845 ( \31222 , \31209 , \31219 );
nand \U$30846 ( \31223 , \31221 , \31222 );
and \U$30847 ( \31224 , \30735 , \31223 );
nor \U$30848 ( \31225 , \30734 , \31224 );
not \U$30849 ( \31226 , \30281 );
not \U$30850 ( \31227 , \30310 );
or \U$30851 ( \31228 , \31226 , \31227 );
or \U$30852 ( \31229 , \30310 , \30281 );
nand \U$30853 ( \31230 , \31228 , \31229 );
not \U$30854 ( \31231 , \31230 );
not \U$30855 ( \31232 , \30261 );
and \U$30856 ( \31233 , \31231 , \31232 );
and \U$30857 ( \31234 , \31230 , \30261 );
nor \U$30858 ( \31235 , \31233 , \31234 );
not \U$30859 ( \31236 , \31235 );
xor \U$30860 ( \31237 , \30708 , \30712 );
and \U$30861 ( \31238 , \31237 , \30723 );
and \U$30862 ( \31239 , \30708 , \30712 );
or \U$30863 ( \31240 , \31238 , \31239 );
not \U$30864 ( \31241 , \31240 );
or \U$30865 ( \31242 , \31236 , \31241 );
or \U$30866 ( \31243 , \31240 , \31235 );
nand \U$30867 ( \31244 , \31242 , \31243 );
not \U$30868 ( \31245 , \31244 );
xor \U$30869 ( \31246 , \30438 , \30452 );
xor \U$30870 ( \31247 , \31246 , \30459 );
not \U$30871 ( \31248 , \31247 );
and \U$30872 ( \31249 , \31245 , \31248 );
and \U$30873 ( \31250 , \31244 , \31247 );
nor \U$30874 ( \31251 , \31249 , \31250 );
xor \U$30875 ( \31252 , \30724 , \30725 );
and \U$30876 ( \31253 , \31252 , \30732 );
and \U$30877 ( \31254 , \30724 , \30725 );
nor \U$30878 ( \31255 , \31253 , \31254 );
xnor \U$30879 ( \31256 , \31251 , \31255 );
or \U$30880 ( \31257 , \31225 , \31256 );
or \U$30881 ( \31258 , \31255 , \31251 );
nand \U$30882 ( \31259 , \31257 , \31258 );
or \U$30883 ( \31260 , \31247 , \31235 );
not \U$30884 ( \31261 , \31235 );
not \U$30885 ( \31262 , \31247 );
or \U$30886 ( \31263 , \31261 , \31262 );
nand \U$30887 ( \31264 , \31263 , \31240 );
nand \U$30888 ( \31265 , \31260 , \31264 );
not \U$30889 ( \31266 , \30368 );
not \U$30890 ( \31267 , \30367 );
not \U$30891 ( \31268 , \30462 );
and \U$30892 ( \31269 , \31267 , \31268 );
and \U$30893 ( \31270 , \30462 , \30367 );
nor \U$30894 ( \31271 , \31269 , \31270 );
not \U$30895 ( \31272 , \31271 );
or \U$30896 ( \31273 , \31266 , \31272 );
or \U$30897 ( \31274 , \31271 , \30368 );
nand \U$30898 ( \31275 , \31273 , \31274 );
xor \U$30899 ( \31276 , \31265 , \31275 );
and \U$30900 ( \31277 , \31259 , \31276 );
and \U$30901 ( \31278 , \31265 , \31275 );
nor \U$30902 ( \31279 , \31277 , \31278 );
or \U$30903 ( \31280 , \30466 , \31279 );
nand \U$30904 ( \31281 , \30465 , \31280 );
and \U$30905 ( \31282 , \30360 , \31281 );
nor \U$30906 ( \31283 , \30359 , \31282 );
or \U$30907 ( \31284 , \30339 , \31283 );
nand \U$30908 ( \31285 , \30338 , \31284 );
not \U$30909 ( \31286 , \30211 );
not \U$30910 ( \31287 , \30079 );
or \U$30911 ( \31288 , \31286 , \31287 );
or \U$30912 ( \31289 , \30079 , \30211 );
nand \U$30913 ( \31290 , \31289 , \30194 );
nand \U$30914 ( \31291 , \31288 , \31290 );
xor \U$30915 ( \31292 , \29751 , \29755 );
xor \U$30916 ( \31293 , \30202 , \30204 );
and \U$30917 ( \31294 , \31293 , \30209 );
and \U$30918 ( \31295 , \30202 , \30204 );
or \U$30919 ( \31296 , \31294 , \31295 );
xor \U$30920 ( \31297 , \31292 , \31296 );
xor \U$30921 ( \31298 , \29831 , \29833 );
xor \U$30922 ( \31299 , \31298 , \29851 );
xor \U$30923 ( \31300 , \31297 , \31299 );
and \U$30924 ( \31301 , \30198 , \30210 );
xor \U$30925 ( \31302 , \31300 , \31301 );
xor \U$30926 ( \31303 , \29967 , \29971 );
and \U$30927 ( \31304 , \31303 , \30078 );
and \U$30928 ( \31305 , \29967 , \29971 );
or \U$30929 ( \31306 , \31304 , \31305 );
xor \U$30930 ( \31307 , \31302 , \31306 );
xor \U$30931 ( \31308 , \31291 , \31307 );
and \U$30932 ( \31309 , \31285 , \31308 );
and \U$30933 ( \31310 , \31291 , \31307 );
nor \U$30934 ( \31311 , \31309 , \31310 );
xor \U$30935 ( \31312 , \31292 , \31296 );
and \U$30936 ( \31313 , \31312 , \31299 );
and \U$30937 ( \31314 , \31292 , \31296 );
or \U$30938 ( \31315 , \31313 , \31314 );
xor \U$30939 ( \31316 , \29756 , \29758 );
xor \U$30940 ( \31317 , \31316 , \29854 );
xnor \U$30941 ( \31318 , \31315 , \31317 );
not \U$30942 ( \31319 , \31318 );
xor \U$30943 ( \31320 , \29745 , \29747 );
not \U$30944 ( \31321 , \31320 );
and \U$30945 ( \31322 , \31319 , \31321 );
and \U$30946 ( \31323 , \31318 , \31320 );
nor \U$30947 ( \31324 , \31322 , \31323 );
xor \U$30948 ( \31325 , \31300 , \31301 );
and \U$30949 ( \31326 , \31325 , \31306 );
and \U$30950 ( \31327 , \31300 , \31301 );
nor \U$30951 ( \31328 , \31326 , \31327 );
xnor \U$30952 ( \31329 , \31324 , \31328 );
or \U$30953 ( \31330 , \31311 , \31329 );
or \U$30954 ( \31331 , \31324 , \31328 );
nand \U$30955 ( \31332 , \31330 , \31331 );
not \U$30956 ( \31333 , \31320 );
not \U$30957 ( \31334 , \31317 );
or \U$30958 ( \31335 , \31333 , \31334 );
or \U$30959 ( \31336 , \31317 , \31320 );
nand \U$30960 ( \31337 , \31336 , \31315 );
nand \U$30961 ( \31338 , \31335 , \31337 );
xor \U$30962 ( \31339 , \29743 , \29748 );
xor \U$30963 ( \31340 , \31339 , \29857 );
xor \U$30964 ( \31341 , \31338 , \31340 );
and \U$30965 ( \31342 , \31332 , \31341 );
and \U$30966 ( \31343 , \31338 , \31340 );
nor \U$30967 ( \31344 , \31342 , \31343 );
or \U$30968 ( \31345 , \29862 , \31344 );
nand \U$30969 ( \31346 , \29861 , \31345 );
and \U$30970 ( \31347 , \29733 , \31346 );
nor \U$30971 ( \31348 , \29732 , \31347 );
or \U$30972 ( \31349 , \29608 , \31348 );
nand \U$30973 ( \31350 , \29607 , \31349 );
and \U$30974 ( \31351 , \29436 , \31350 );
nor \U$30975 ( \31352 , \29435 , \31351 );
or \U$30976 ( \31353 , \29280 , \31352 );
nand \U$30977 ( \31354 , \29279 , \31353 );
not \U$30978 ( \31355 , \29091 );
nor \U$30979 ( \31356 , \31355 , \29256 );
xor \U$30980 ( \31357 , \28714 , \29052 );
xor \U$30981 ( \31358 , \31357 , \29069 );
xor \U$30982 ( \31359 , \31356 , \31358 );
and \U$30983 ( \31360 , \31354 , \31359 );
and \U$30984 ( \31361 , \31356 , \31358 );
nor \U$30985 ( \31362 , \31360 , \31361 );
or \U$30986 ( \31363 , \29087 , \31362 );
nand \U$30987 ( \31364 , \29086 , \31363 );
not \U$30988 ( \31365 , \29073 );
not \U$30989 ( \31366 , \29081 );
or \U$30990 ( \31367 , \31365 , \31366 );
or \U$30991 ( \31368 , \29081 , \29073 );
nand \U$30992 ( \31369 , \31368 , \29077 );
nand \U$30993 ( \31370 , \31367 , \31369 );
xor \U$30994 ( \31371 , \28532 , \28693 );
xor \U$30995 ( \31372 , \31371 , \28704 );
xor \U$30996 ( \31373 , \31370 , \31372 );
and \U$30997 ( \31374 , \31364 , \31373 );
and \U$30998 ( \31375 , \31370 , \31372 );
nor \U$30999 ( \31376 , \31374 , \31375 );
or \U$31000 ( \31377 , \28709 , \31376 );
nand \U$31001 ( \31378 , \28708 , \31377 );
and \U$31002 ( \31379 , \28521 , \31378 );
nor \U$31003 ( \31380 , \28520 , \31379 );
or \U$31004 ( \31381 , \28303 , \31380 );
nand \U$31005 ( \31382 , \28302 , \31381 );
and \U$31006 ( \31383 , \28125 , \31382 );
nor \U$31007 ( \31384 , \28124 , \31383 );
xor \U$31008 ( \31385 , \27918 , \27920 );
and \U$31009 ( \31386 , \31385 , \27925 );
and \U$31010 ( \31387 , \27918 , \27920 );
or \U$31011 ( \31388 , \31386 , \31387 );
not \U$31012 ( \31389 , \31388 );
not \U$31013 ( \31390 , \27517 );
nand \U$31014 ( \31391 , \31390 , \27506 );
not \U$31015 ( \31392 , \31391 );
and \U$31016 ( \31393 , \31389 , \31392 );
and \U$31017 ( \31394 , \31388 , \31391 );
nor \U$31018 ( \31395 , \31393 , \31394 );
not \U$31019 ( \31396 , \31395 );
xor \U$31020 ( \31397 , \27063 , \27233 );
xor \U$31021 ( \31398 , \31397 , \27262 );
xor \U$31022 ( \31399 , \27489 , \27494 );
xor \U$31023 ( \31400 , \31398 , \31399 );
not \U$31024 ( \31401 , \31400 );
and \U$31025 ( \31402 , \31396 , \31401 );
and \U$31026 ( \31403 , \31395 , \31400 );
nor \U$31027 ( \31404 , \31402 , \31403 );
xor \U$31028 ( \31405 , \27521 , \27904 );
and \U$31029 ( \31406 , \31405 , \27926 );
and \U$31030 ( \31407 , \27521 , \27904 );
nor \U$31031 ( \31408 , \31406 , \31407 );
xnor \U$31032 ( \31409 , \31404 , \31408 );
or \U$31033 ( \31410 , \31384 , \31409 );
or \U$31034 ( \31411 , \31404 , \31408 );
nand \U$31035 ( \31412 , \31410 , \31411 );
not \U$31036 ( \31413 , \31400 );
or \U$31037 ( \31414 , \31413 , \31391 );
not \U$31038 ( \31415 , \31391 );
not \U$31039 ( \31416 , \31413 );
or \U$31040 ( \31417 , \31415 , \31416 );
nand \U$31041 ( \31418 , \31417 , \31388 );
nand \U$31042 ( \31419 , \31414 , \31418 );
xor \U$31043 ( \31420 , \27307 , \27317 );
xor \U$31044 ( \31421 , \31420 , \27499 );
xor \U$31045 ( \31422 , \31419 , \31421 );
and \U$31046 ( \31423 , \31412 , \31422 );
and \U$31047 ( \31424 , \31419 , \31421 );
nor \U$31048 ( \31425 , \31423 , \31424 );
or \U$31049 ( \31426 , \27504 , \31425 );
nand \U$31050 ( \31427 , \27503 , \31426 );
not \U$31051 ( \31428 , \27301 );
not \U$31052 ( \31429 , \27294 );
or \U$31053 ( \31430 , \31428 , \31429 );
or \U$31054 ( \31431 , \27294 , \27301 );
nand \U$31055 ( \31432 , \31431 , \27288 );
nand \U$31056 ( \31433 , \31430 , \31432 );
not \U$31057 ( \31434 , \27042 );
not \U$31058 ( \31435 , \27039 );
or \U$31059 ( \31436 , \31434 , \31435 );
or \U$31060 ( \31437 , \27039 , \27042 );
nand \U$31061 ( \31438 , \31436 , \31437 );
xor \U$31062 ( \31439 , \31433 , \31438 );
and \U$31063 ( \31440 , \31427 , \31439 );
and \U$31064 ( \31441 , \31433 , \31438 );
nor \U$31065 ( \31442 , \31440 , \31441 );
or \U$31066 ( \31443 , \27045 , \31442 );
nand \U$31067 ( \31444 , \27044 , \31443 );
not \U$31068 ( \31445 , \26780 );
nor \U$31069 ( \31446 , \31445 , \27033 );
not \U$31070 ( \31447 , \26775 );
not \U$31071 ( \31448 , \26534 );
or \U$31072 ( \31449 , \31447 , \31448 );
or \U$31073 ( \31450 , \26534 , \26775 );
nand \U$31074 ( \31451 , \31449 , \31450 );
xor \U$31075 ( \31452 , \31446 , \31451 );
and \U$31076 ( \31453 , \31444 , \31452 );
and \U$31077 ( \31454 , \31446 , \31451 );
nor \U$31078 ( \31455 , \31453 , \31454 );
or \U$31079 ( \31456 , \26778 , \31455 );
nand \U$31080 ( \31457 , \26777 , \31456 );
and \U$31081 ( \31458 , \26522 , \31457 );
nor \U$31082 ( \31459 , \26521 , \31458 );
not \U$31083 ( \31460 , \26241 );
nand \U$31084 ( \31461 , \31460 , \26215 );
xor \U$31085 ( \31462 , \25419 , \25421 );
xor \U$31086 ( \31463 , \31462 , \25436 );
not \U$31087 ( \31464 , \26237 );
not \U$31088 ( \31465 , \26234 );
or \U$31089 ( \31466 , \31464 , \31465 );
or \U$31090 ( \31467 , \26234 , \26237 );
nand \U$31091 ( \31468 , \31467 , \26232 );
nand \U$31092 ( \31469 , \31466 , \31468 );
xnor \U$31093 ( \31470 , \31463 , \31469 );
not \U$31094 ( \31471 , \31470 );
xor \U$31095 ( \31472 , \25714 , \25721 );
xor \U$31096 ( \31473 , \31472 , \25726 );
not \U$31097 ( \31474 , \31473 );
and \U$31098 ( \31475 , \31471 , \31474 );
and \U$31099 ( \31476 , \31470 , \31473 );
nor \U$31100 ( \31477 , \31475 , \31476 );
xnor \U$31101 ( \31478 , \31461 , \31477 );
or \U$31102 ( \31479 , \31459 , \31478 );
or \U$31103 ( \31480 , \31461 , \31477 );
nand \U$31104 ( \31481 , \31479 , \31480 );
not \U$31105 ( \31482 , \31463 );
not \U$31106 ( \31483 , \31473 );
or \U$31107 ( \31484 , \31482 , \31483 );
or \U$31108 ( \31485 , \31473 , \31463 );
nand \U$31109 ( \31486 , \31485 , \31469 );
nand \U$31110 ( \31487 , \31484 , \31486 );
xor \U$31111 ( \31488 , \25447 , \25449 );
xor \U$31112 ( \31489 , \31488 , \25729 );
xor \U$31113 ( \31490 , \31487 , \31489 );
and \U$31114 ( \31491 , \31481 , \31490 );
and \U$31115 ( \31492 , \31487 , \31489 );
nor \U$31116 ( \31493 , \31491 , \31492 );
or \U$31117 ( \31494 , \25740 , \31493 );
nand \U$31118 ( \31495 , \25739 , \31494 );
and \U$31119 ( \31496 , \25446 , \31495 );
nor \U$31120 ( \31497 , \25445 , \31496 );
xor \U$31121 ( \31498 , \25168 , \25172 );
and \U$31122 ( \31499 , \31498 , \25177 );
and \U$31123 ( \31500 , \25168 , \25172 );
or \U$31124 ( \31501 , \31499 , \31500 );
and \U$31125 ( \31502 , \24641 , \24643 );
xnor \U$31126 ( \31503 , \31501 , \31502 );
not \U$31127 ( \31504 , \31503 );
xor \U$31128 ( \31505 , \24621 , \24623 );
xor \U$31129 ( \31506 , \31505 , \24628 );
not \U$31130 ( \31507 , \31506 );
and \U$31131 ( \31508 , \31504 , \31507 );
and \U$31132 ( \31509 , \31503 , \31506 );
nor \U$31133 ( \31510 , \31508 , \31509 );
xor \U$31134 ( \31511 , \24644 , \25166 );
and \U$31135 ( \31512 , \31511 , \25178 );
and \U$31136 ( \31513 , \24644 , \25166 );
nor \U$31137 ( \31514 , \31512 , \31513 );
xnor \U$31138 ( \31515 , \31510 , \31514 );
or \U$31139 ( \31516 , \31497 , \31515 );
or \U$31140 ( \31517 , \31510 , \31514 );
nand \U$31141 ( \31518 , \31516 , \31517 );
xor \U$31142 ( \31519 , \24345 , \24631 );
xor \U$31143 ( \31520 , \31519 , \24634 );
not \U$31144 ( \31521 , \31502 );
not \U$31145 ( \31522 , \31506 );
or \U$31146 ( \31523 , \31521 , \31522 );
or \U$31147 ( \31524 , \31506 , \31502 );
nand \U$31148 ( \31525 , \31524 , \31501 );
nand \U$31149 ( \31526 , \31523 , \31525 );
xor \U$31150 ( \31527 , \31520 , \31526 );
and \U$31151 ( \31528 , \31518 , \31527 );
and \U$31152 ( \31529 , \31520 , \31526 );
nor \U$31153 ( \31530 , \31528 , \31529 );
or \U$31154 ( \31531 , \24639 , \31530 );
nand \U$31155 ( \31532 , \24638 , \31531 );
or \U$31156 ( \31533 , \24339 , \24025 );
not \U$31157 ( \31534 , \24025 );
not \U$31158 ( \31535 , \24339 );
or \U$31159 ( \31536 , \31534 , \31535 );
nand \U$31160 ( \31537 , \31536 , \24328 );
nand \U$31161 ( \31538 , \31533 , \31537 );
xor \U$31162 ( \31539 , \23688 , \23690 );
xor \U$31163 ( \31540 , \31539 , \24010 );
xor \U$31164 ( \31541 , \31538 , \31540 );
and \U$31165 ( \31542 , \31532 , \31541 );
and \U$31166 ( \31543 , \31538 , \31540 );
nor \U$31167 ( \31544 , \31542 , \31543 );
or \U$31168 ( \31545 , \24015 , \31544 );
nand \U$31169 ( \31546 , \24014 , \31545 );
or \U$31170 ( \31547 , \23682 , \23365 );
not \U$31171 ( \31548 , \23365 );
not \U$31172 ( \31549 , \23682 );
or \U$31173 ( \31550 , \31548 , \31549 );
nand \U$31174 ( \31551 , \31550 , \23671 );
nand \U$31175 ( \31552 , \31547 , \31551 );
xor \U$31176 ( \31553 , \23033 , \23035 );
xor \U$31177 ( \31554 , \31553 , \23350 );
xor \U$31178 ( \31555 , \31552 , \31554 );
and \U$31179 ( \31556 , \31546 , \31555 );
and \U$31180 ( \31557 , \31552 , \31554 );
nor \U$31181 ( \31558 , \31556 , \31557 );
or \U$31182 ( \31559 , \23355 , \31558 );
nand \U$31183 ( \31560 , \23354 , \31559 );
and \U$31184 ( \31561 , \23018 , \31560 );
nor \U$31185 ( \31562 , \23017 , \31561 );
or \U$31186 ( \31563 , \22662 , \31562 );
nand \U$31187 ( \31564 , \22661 , \31563 );
not \U$31188 ( \31565 , \22325 );
not \U$31189 ( \31566 , \22318 );
or \U$31190 ( \31567 , \31565 , \31566 );
or \U$31191 ( \31568 , \22318 , \22325 );
nand \U$31192 ( \31569 , \31568 , \22316 );
nand \U$31193 ( \31570 , \31567 , \31569 );
not \U$31194 ( \31571 , \21949 );
not \U$31195 ( \31572 , \21960 );
or \U$31196 ( \31573 , \31571 , \31572 );
or \U$31197 ( \31574 , \21960 , \21949 );
nand \U$31198 ( \31575 , \31573 , \31574 );
xor \U$31199 ( \31576 , \31570 , \31575 );
and \U$31200 ( \31577 , \31564 , \31576 );
and \U$31201 ( \31578 , \31570 , \31575 );
nor \U$31202 ( \31579 , \31577 , \31578 );
or \U$31203 ( \31580 , \21963 , \31579 );
nand \U$31204 ( \31581 , \21962 , \31580 );
and \U$31205 ( \31582 , \21934 , \31581 );
nor \U$31206 ( \31583 , \21933 , \31582 );
not \U$31207 ( \31584 , \21554 );
nand \U$31208 ( \31585 , \31584 , \21186 );
not \U$31209 ( \31586 , \20373 );
not \U$31210 ( \31587 , \20399 );
or \U$31211 ( \31588 , \31586 , \31587 );
or \U$31212 ( \31589 , \20399 , \20373 );
nand \U$31213 ( \31590 , \31588 , \31589 );
not \U$31214 ( \31591 , \31590 );
not \U$31215 ( \31592 , \20383 );
and \U$31216 ( \31593 , \31591 , \31592 );
and \U$31217 ( \31594 , \31590 , \20383 );
nor \U$31218 ( \31595 , \31593 , \31594 );
not \U$31219 ( \31596 , \31595 );
xor \U$31220 ( \31597 , \21157 , \21179 );
and \U$31221 ( \31598 , \31597 , \21184 );
and \U$31222 ( \31599 , \21157 , \21179 );
or \U$31223 ( \31600 , \31598 , \31599 );
not \U$31224 ( \31601 , \31600 );
and \U$31225 ( \31602 , \31596 , \31601 );
and \U$31226 ( \31603 , \31595 , \31600 );
nor \U$31227 ( \31604 , \31602 , \31603 );
not \U$31228 ( \31605 , \31604 );
xor \U$31229 ( \31606 , \19956 , \19958 );
xor \U$31230 ( \31607 , \31606 , \19963 );
xor \U$31231 ( \31608 , \20004 , \20009 );
xor \U$31232 ( \31609 , \31607 , \31608 );
not \U$31233 ( \31610 , \31609 );
and \U$31234 ( \31611 , \31605 , \31610 );
and \U$31235 ( \31612 , \31604 , \31609 );
nor \U$31236 ( \31613 , \31611 , \31612 );
not \U$31237 ( \31614 , \31613 );
xor \U$31238 ( \31615 , \21146 , \21152 );
and \U$31239 ( \31616 , \31615 , \21185 );
and \U$31240 ( \31617 , \21146 , \21152 );
or \U$31241 ( \31618 , \31616 , \31617 );
not \U$31242 ( \31619 , \31618 );
and \U$31243 ( \31620 , \31614 , \31619 );
and \U$31244 ( \31621 , \31613 , \31618 );
nor \U$31245 ( \31622 , \31620 , \31621 );
xnor \U$31246 ( \31623 , \31585 , \31622 );
or \U$31247 ( \31624 , \31583 , \31623 );
or \U$31248 ( \31625 , \31585 , \31622 );
nand \U$31249 ( \31626 , \31624 , \31625 );
not \U$31250 ( \31627 , \31618 );
nor \U$31251 ( \31628 , \31627 , \31613 );
xor \U$31252 ( \31629 , \19954 , \19966 );
xor \U$31253 ( \31630 , \31629 , \19971 );
xor \U$31254 ( \31631 , \20002 , \20014 );
xor \U$31255 ( \31632 , \31631 , \20401 );
xor \U$31256 ( \31633 , \31630 , \31632 );
not \U$31257 ( \31634 , \31609 );
or \U$31258 ( \31635 , \31595 , \31634 );
not \U$31259 ( \31636 , \31634 );
not \U$31260 ( \31637 , \31595 );
or \U$31261 ( \31638 , \31636 , \31637 );
nand \U$31262 ( \31639 , \31638 , \31600 );
nand \U$31263 ( \31640 , \31635 , \31639 );
xor \U$31264 ( \31641 , \31633 , \31640 );
xor \U$31265 ( \31642 , \31628 , \31641 );
and \U$31266 ( \31643 , \31626 , \31642 );
and \U$31267 ( \31644 , \31628 , \31641 );
nor \U$31268 ( \31645 , \31643 , \31644 );
not \U$31269 ( \31646 , \19999 );
not \U$31270 ( \31647 , \20404 );
and \U$31271 ( \31648 , \31646 , \31647 );
and \U$31272 ( \31649 , \19999 , \20404 );
nor \U$31273 ( \31650 , \31648 , \31649 );
xor \U$31274 ( \31651 , \31630 , \31632 );
and \U$31275 ( \31652 , \31651 , \31640 );
and \U$31276 ( \31653 , \31630 , \31632 );
nor \U$31277 ( \31654 , \31652 , \31653 );
xnor \U$31278 ( \31655 , \31650 , \31654 );
or \U$31279 ( \31656 , \31645 , \31655 );
or \U$31280 ( \31657 , \31650 , \31654 );
nand \U$31281 ( \31658 , \31656 , \31657 );
and \U$31282 ( \31659 , \20407 , \31658 );
nor \U$31283 ( \31660 , \20406 , \31659 );
not \U$31284 ( \31661 , \19980 );
nand \U$31285 ( \31662 , \31661 , \19993 );
xor \U$31286 ( \31663 , \18773 , \18785 );
xor \U$31287 ( \31664 , \31663 , \19162 );
xor \U$31288 ( \31665 , \19142 , \19144 );
xor \U$31289 ( \31666 , \31665 , \19159 );
and \U$31290 ( \31667 , \19987 , \31666 );
xor \U$31291 ( \31668 , \19142 , \19144 );
xor \U$31292 ( \31669 , \31668 , \19159 );
and \U$31293 ( \31670 , \19991 , \31669 );
and \U$31294 ( \31671 , \19987 , \19991 );
or \U$31295 ( \31672 , \31667 , \31670 , \31671 );
xnor \U$31296 ( \31673 , \31664 , \31672 );
not \U$31297 ( \31674 , \31673 );
xor \U$31298 ( \31675 , \18725 , \18737 );
xor \U$31299 ( \31676 , \31675 , \18742 );
not \U$31300 ( \31677 , \31676 );
and \U$31301 ( \31678 , \31674 , \31677 );
and \U$31302 ( \31679 , \31673 , \31676 );
nor \U$31303 ( \31680 , \31678 , \31679 );
xnor \U$31304 ( \31681 , \31662 , \31680 );
or \U$31305 ( \31682 , \31660 , \31681 );
or \U$31306 ( \31683 , \31662 , \31680 );
nand \U$31307 ( \31684 , \31682 , \31683 );
not \U$31308 ( \31685 , \31676 );
not \U$31309 ( \31686 , \31664 );
or \U$31310 ( \31687 , \31685 , \31686 );
or \U$31311 ( \31688 , \31664 , \31676 );
nand \U$31312 ( \31689 , \31688 , \31672 );
nand \U$31313 ( \31690 , \31687 , \31689 );
not \U$31314 ( \31691 , \19165 );
not \U$31315 ( \31692 , \19170 );
or \U$31316 ( \31693 , \31691 , \31692 );
or \U$31317 ( \31694 , \19170 , \19165 );
nand \U$31318 ( \31695 , \31693 , \31694 );
xor \U$31319 ( \31696 , \31690 , \31695 );
and \U$31320 ( \31697 , \31684 , \31696 );
and \U$31321 ( \31698 , \31690 , \31695 );
nor \U$31322 ( \31699 , \31697 , \31698 );
or \U$31323 ( \31700 , \19176 , \31699 );
nand \U$31324 ( \31701 , \19172 , \31700 );
and \U$31325 ( \31702 , \18768 , \31701 );
nor \U$31326 ( \31703 , \18767 , \31702 );
not \U$31327 ( \31704 , \17922 );
not \U$31328 ( \31705 , \17933 );
and \U$31329 ( \31706 , \31704 , \31705 );
and \U$31330 ( \31707 , \17922 , \17933 );
not \U$31331 ( \31708 , \18353 );
nor \U$31332 ( \31709 , \31707 , \31708 );
nor \U$31333 ( \31710 , \31706 , \31709 );
or \U$31334 ( \31711 , \17918 , \17820 );
not \U$31335 ( \31712 , \17820 );
not \U$31336 ( \31713 , \17918 );
or \U$31337 ( \31714 , \31712 , \31713 );
nand \U$31338 ( \31715 , \31714 , \17899 );
nand \U$31339 ( \31716 , \31711 , \31715 );
xor \U$31340 ( \31717 , \15588 , \15598 );
xor \U$31341 ( \31718 , \31717 , \15603 );
xor \U$31342 ( \31719 , \16502 , \16509 );
xor \U$31343 ( \31720 , \31718 , \31719 );
not \U$31344 ( \31721 , \31720 );
or \U$31345 ( \31722 , \17908 , \17906 );
not \U$31346 ( \31723 , \17906 );
not \U$31347 ( \31724 , \17908 );
or \U$31348 ( \31725 , \31723 , \31724 );
nand \U$31349 ( \31726 , \31725 , \17914 );
nand \U$31350 ( \31727 , \31722 , \31726 );
not \U$31351 ( \31728 , \31727 );
not \U$31352 ( \31729 , \17876 );
not \U$31353 ( \31730 , \17831 );
and \U$31354 ( \31731 , \31729 , \31730 );
and \U$31355 ( \31732 , \17876 , \17831 );
nor \U$31356 ( \31733 , \31732 , \17894 );
nor \U$31357 ( \31734 , \31731 , \31733 );
not \U$31358 ( \31735 , \31734 );
and \U$31359 ( \31736 , \31728 , \31735 );
and \U$31360 ( \31737 , \31727 , \31734 );
nor \U$31361 ( \31738 , \31736 , \31737 );
not \U$31362 ( \31739 , \31738 );
or \U$31363 ( \31740 , \31721 , \31739 );
or \U$31364 ( \31741 , \31738 , \31720 );
nand \U$31365 ( \31742 , \31740 , \31741 );
xnor \U$31366 ( \31743 , \31716 , \31742 );
not \U$31367 ( \31744 , \31743 );
xor \U$31368 ( \31745 , \16099 , \16479 );
xor \U$31369 ( \31746 , \31745 , \16494 );
xor \U$31370 ( \31747 , \16609 , \16611 );
xor \U$31371 ( \31748 , \31747 , \17057 );
xor \U$31372 ( \31749 , \31746 , \31748 );
not \U$31373 ( \31750 , \31749 );
and \U$31374 ( \31751 , \31744 , \31750 );
and \U$31375 ( \31752 , \31743 , \31749 );
nor \U$31376 ( \31753 , \31751 , \31752 );
xnor \U$31377 ( \31754 , \31710 , \31753 );
or \U$31378 ( \31755 , \31703 , \31754 );
or \U$31379 ( \31756 , \31710 , \31753 );
nand \U$31380 ( \31757 , \31755 , \31756 );
not \U$31381 ( \31758 , \31749 );
not \U$31382 ( \31759 , \31742 );
or \U$31383 ( \31760 , \31758 , \31759 );
or \U$31384 ( \31761 , \31742 , \31749 );
nand \U$31385 ( \31762 , \31761 , \31716 );
nand \U$31386 ( \31763 , \31760 , \31762 );
xor \U$31387 ( \31764 , \16595 , \17060 );
xor \U$31388 ( \31765 , \31764 , \17063 );
not \U$31389 ( \31766 , \31765 );
and \U$31390 ( \31767 , \31727 , \31720 );
not \U$31391 ( \31768 , \31727 );
not \U$31392 ( \31769 , \31720 );
and \U$31393 ( \31770 , \31768 , \31769 );
nor \U$31394 ( \31771 , \31770 , \31734 );
nor \U$31395 ( \31772 , \31767 , \31771 );
not \U$31396 ( \31773 , \31772 );
and \U$31397 ( \31774 , \31746 , \31748 );
not \U$31398 ( \31775 , \31774 );
and \U$31399 ( \31776 , \31773 , \31775 );
and \U$31400 ( \31777 , \31772 , \31774 );
nor \U$31401 ( \31778 , \31776 , \31777 );
not \U$31402 ( \31779 , \31778 );
or \U$31403 ( \31780 , \31766 , \31779 );
or \U$31404 ( \31781 , \31778 , \31765 );
nand \U$31405 ( \31782 , \31780 , \31781 );
xor \U$31406 ( \31783 , \31763 , \31782 );
and \U$31407 ( \31784 , \31757 , \31783 );
and \U$31408 ( \31785 , \31763 , \31782 );
nor \U$31409 ( \31786 , \31784 , \31785 );
and \U$31410 ( \31787 , \31765 , \31774 );
not \U$31411 ( \31788 , \31765 );
not \U$31412 ( \31789 , \31774 );
and \U$31413 ( \31790 , \31788 , \31789 );
nor \U$31414 ( \31791 , \31790 , \31772 );
nor \U$31415 ( \31792 , \31787 , \31791 );
xnor \U$31416 ( \31793 , \16591 , \17066 );
not \U$31417 ( \31794 , \31793 );
not \U$31418 ( \31795 , \16588 );
and \U$31419 ( \31796 , \31794 , \31795 );
and \U$31420 ( \31797 , \31793 , \16588 );
nor \U$31421 ( \31798 , \31796 , \31797 );
xnor \U$31422 ( \31799 , \31792 , \31798 );
or \U$31423 ( \31800 , \31786 , \31799 );
or \U$31424 ( \31801 , \31792 , \31798 );
nand \U$31425 ( \31802 , \31800 , \31801 );
and \U$31426 ( \31803 , \17070 , \31802 );
nor \U$31427 ( \31804 , \17069 , \31803 );
xnor \U$31428 ( \31805 , \16554 , \16583 );
or \U$31429 ( \31806 , \31804 , \31805 );
nand \U$31430 ( \31807 , \16585 , \31806 );
xor \U$31431 ( \31808 , \16563 , \16565 );
and \U$31432 ( \31809 , \31808 , \16582 );
and \U$31433 ( \31810 , \16563 , \16565 );
or \U$31434 ( \31811 , \31809 , \31810 );
xor \U$31435 ( \31812 , \16570 , \16576 );
and \U$31436 ( \31813 , \31812 , \16581 );
and \U$31437 ( \31814 , \16570 , \16576 );
or \U$31438 ( \31815 , \31813 , \31814 );
not \U$31439 ( \31816 , \31815 );
not \U$31440 ( \31817 , \15160 );
not \U$31441 ( \31818 , \14725 );
or \U$31442 ( \31819 , \31817 , \31818 );
or \U$31443 ( \31820 , \14725 , \15160 );
nand \U$31444 ( \31821 , \31819 , \31820 );
not \U$31445 ( \31822 , \31821 );
not \U$31446 ( \31823 , \14729 );
and \U$31447 ( \31824 , \31822 , \31823 );
and \U$31448 ( \31825 , \31821 , \14729 );
nor \U$31449 ( \31826 , \31824 , \31825 );
not \U$31450 ( \31827 , \31826 );
or \U$31451 ( \31828 , \31816 , \31827 );
or \U$31452 ( \31829 , \31826 , \31815 );
nand \U$31453 ( \31830 , \31828 , \31829 );
xor \U$31454 ( \31831 , \31811 , \31830 );
and \U$31455 ( \31832 , \31807 , \31831 );
and \U$31456 ( \31833 , \31830 , \31811 );
nor \U$31457 ( \31834 , \31832 , \31833 );
not \U$31458 ( \31835 , \31826 );
nand \U$31459 ( \31836 , \31835 , \31815 );
not \U$31460 ( \31837 , \15162 );
not \U$31461 ( \31838 , \14717 );
or \U$31462 ( \31839 , \31837 , \31838 );
or \U$31463 ( \31840 , \14717 , \15162 );
nand \U$31464 ( \31841 , \31839 , \31840 );
not \U$31465 ( \31842 , \31841 );
not \U$31466 ( \31843 , \14719 );
and \U$31467 ( \31844 , \31842 , \31843 );
and \U$31468 ( \31845 , \31841 , \14719 );
nor \U$31469 ( \31846 , \31844 , \31845 );
xnor \U$31470 ( \31847 , \31836 , \31846 );
or \U$31471 ( \31848 , \31834 , \31847 );
or \U$31472 ( \31849 , \31836 , \31846 );
nand \U$31473 ( \31850 , \31848 , \31849 );
and \U$31474 ( \31851 , \15171 , \31850 );
nor \U$31475 ( \31852 , \15170 , \31851 );
or \U$31476 ( \31853 , \14715 , \31852 );
nand \U$31477 ( \31854 , \14714 , \31853 );
not \U$31478 ( \31855 , \13804 );
nor \U$31479 ( \31856 , \31855 , \14260 );
xor \U$31480 ( \31857 , \13751 , \13770 );
and \U$31481 ( \31858 , \31857 , \13803 );
and \U$31482 ( \31859 , \13751 , \13770 );
or \U$31483 ( \31860 , \31858 , \31859 );
xor \U$31484 ( \31861 , \12481 , \12875 );
xor \U$31485 ( \31862 , \31861 , \12880 );
xor \U$31486 ( \31863 , \31860 , \31862 );
xor \U$31487 ( \31864 , \12060 , \12425 );
xor \U$31488 ( \31865 , \31864 , \12442 );
not \U$31489 ( \31866 , \31865 );
xor \U$31490 ( \31867 , \13795 , \13797 );
and \U$31491 ( \31868 , \31867 , \13802 );
and \U$31492 ( \31869 , \13795 , \13797 );
or \U$31493 ( \31870 , \31868 , \31869 );
not \U$31494 ( \31871 , \31870 );
not \U$31495 ( \31872 , \13761 );
nand \U$31496 ( \31873 , \31872 , \13766 );
not \U$31497 ( \31874 , \31873 );
and \U$31498 ( \31875 , \31871 , \31874 );
and \U$31499 ( \31876 , \31870 , \31873 );
nor \U$31500 ( \31877 , \31875 , \31876 );
not \U$31501 ( \31878 , \31877 );
or \U$31502 ( \31879 , \31866 , \31878 );
or \U$31503 ( \31880 , \31877 , \31865 );
nand \U$31504 ( \31881 , \31879 , \31880 );
xor \U$31505 ( \31882 , \31863 , \31881 );
xor \U$31506 ( \31883 , \31856 , \31882 );
and \U$31507 ( \31884 , \31854 , \31883 );
and \U$31508 ( \31885 , \31856 , \31882 );
nor \U$31509 ( \31886 , \31884 , \31885 );
not \U$31510 ( \31887 , \31886 );
xor \U$31511 ( \31888 , \31860 , \31862 );
and \U$31512 ( \31889 , \31888 , \31881 );
and \U$31513 ( \31890 , \31860 , \31862 );
or \U$31514 ( \31891 , \31889 , \31890 );
and \U$31515 ( \31892 , \31870 , \31865 );
not \U$31516 ( \31893 , \31870 );
not \U$31517 ( \31894 , \31865 );
and \U$31518 ( \31895 , \31893 , \31894 );
nor \U$31519 ( \31896 , \31895 , \31873 );
nor \U$31520 ( \31897 , \31892 , \31896 );
not \U$31521 ( \31898 , \31897 );
xor \U$31522 ( \31899 , \12030 , \12445 );
xor \U$31523 ( \31900 , \31899 , \12448 );
xor \U$31524 ( \31901 , \12464 , \12883 );
xor \U$31525 ( \31902 , \31900 , \31901 );
not \U$31526 ( \31903 , \31902 );
or \U$31527 ( \31904 , \31898 , \31903 );
or \U$31528 ( \31905 , \31902 , \31897 );
nand \U$31529 ( \31906 , \31904 , \31905 );
xor \U$31530 ( \31907 , \31891 , \31906 );
and \U$31531 ( \31908 , \31887 , \31907 );
and \U$31532 ( \31909 , \31906 , \31891 );
nor \U$31533 ( \31910 , \31908 , \31909 );
not \U$31534 ( \31911 , \31897 );
nand \U$31535 ( \31912 , \31911 , \31902 );
not \U$31536 ( \31913 , \12895 );
not \U$31537 ( \31914 , \12888 );
and \U$31538 ( \31915 , \31913 , \31914 );
and \U$31539 ( \31916 , \12895 , \12888 );
nor \U$31540 ( \31917 , \31915 , \31916 );
xnor \U$31541 ( \31918 , \31912 , \31917 );
or \U$31542 ( \31919 , \31910 , \31918 );
or \U$31543 ( \31920 , \31912 , \31917 );
nand \U$31544 ( \31921 , \31919 , \31920 );
and \U$31545 ( \31922 , \12898 , \31921 );
nor \U$31546 ( \31923 , \12897 , \31922 );
not \U$31547 ( \31924 , \12458 );
nand \U$31548 ( \31925 , \31924 , \12453 );
not \U$31549 ( \31926 , \12001 );
not \U$31550 ( \31927 , \11612 );
and \U$31551 ( \31928 , \31926 , \31927 );
and \U$31552 ( \31929 , \12001 , \11612 );
nor \U$31553 ( \31930 , \31928 , \31929 );
xnor \U$31554 ( \31931 , \31925 , \31930 );
or \U$31555 ( \31932 , \31923 , \31931 );
or \U$31556 ( \31933 , \31925 , \31930 );
nand \U$31557 ( \31934 , \31932 , \31933 );
and \U$31558 ( \31935 , \12004 , \31934 );
nor \U$31559 ( \31936 , \12003 , \31935 );
xor \U$31560 ( \31937 , \11199 , \11201 );
not \U$31561 ( \31938 , \31937 );
not \U$31562 ( \31939 , \11598 );
nand \U$31563 ( \31940 , \31939 , \11206 );
not \U$31564 ( \31941 , \31940 );
and \U$31565 ( \31942 , \31938 , \31941 );
and \U$31566 ( \31943 , \31937 , \31940 );
nor \U$31567 ( \31944 , \31942 , \31943 );
or \U$31568 ( \31945 , \31936 , \31944 );
not \U$31569 ( \31946 , \31937 );
or \U$31570 ( \31947 , \31940 , \31946 );
nand \U$31571 ( \31948 , \31945 , \31947 );
and \U$31572 ( \31949 , \11204 , \31948 );
nor \U$31573 ( \31950 , \11203 , \31949 );
not \U$31574 ( \31951 , \31950 );
and \U$31575 ( \31952 , \10818 , \31951 );
nor \U$31576 ( \31953 , \10817 , \31952 );
not \U$31577 ( \31954 , \10414 );
nand \U$31578 ( \31955 , \31954 , \10411 );
not \U$31579 ( \31956 , \9670 );
not \U$31580 ( \31957 , \10041 );
and \U$31581 ( \31958 , \31956 , \31957 );
and \U$31582 ( \31959 , \9670 , \10041 );
nor \U$31583 ( \31960 , \31958 , \31959 );
xnor \U$31584 ( \31961 , \31955 , \31960 );
or \U$31585 ( \31962 , \31953 , \31961 );
or \U$31586 ( \31963 , \31955 , \31960 );
nand \U$31587 ( \31964 , \31962 , \31963 );
and \U$31588 ( \31965 , \10044 , \31964 );
nor \U$31589 ( \31966 , \10043 , \31965 );
not \U$31590 ( \31967 , \31966 );
and \U$31591 ( \31968 , \9641 , \9667 );
xor \U$31592 ( \31969 , \9645 , \9647 );
and \U$31593 ( \31970 , \31969 , \9666 );
and \U$31594 ( \31971 , \9645 , \9647 );
nor \U$31595 ( \31972 , \31970 , \31971 );
not \U$31596 ( \31973 , \31972 );
xor \U$31597 ( \31974 , \8170 , \8172 );
xor \U$31598 ( \31975 , \31974 , \8193 );
xor \U$31599 ( \31976 , \9652 , \9660 );
and \U$31600 ( \31977 , \31976 , \9665 );
and \U$31601 ( \31978 , \9652 , \9660 );
or \U$31602 ( \31979 , \31977 , \31978 );
xor \U$31603 ( \31980 , \8548 , \8560 );
xor \U$31604 ( \31981 , \31980 , \8563 );
xor \U$31605 ( \31982 , \31979 , \31981 );
xor \U$31606 ( \31983 , \31975 , \31982 );
not \U$31607 ( \31984 , \31983 );
or \U$31608 ( \31985 , \31973 , \31984 );
or \U$31609 ( \31986 , \31983 , \31972 );
nand \U$31610 ( \31987 , \31985 , \31986 );
xor \U$31611 ( \31988 , \31968 , \31987 );
and \U$31612 ( \31989 , \31967 , \31988 );
and \U$31613 ( \31990 , \31968 , \31987 );
nor \U$31614 ( \31991 , \31989 , \31990 );
not \U$31615 ( \31992 , \31972 );
nand \U$31616 ( \31993 , \31992 , \31983 );
xor \U$31617 ( \31994 , \8566 , \8571 );
xor \U$31618 ( \31995 , \31994 , \8574 );
not \U$31619 ( \31996 , \31995 );
xor \U$31620 ( \31997 , \8170 , \8172 );
xor \U$31621 ( \31998 , \31997 , \8193 );
and \U$31622 ( \31999 , \31979 , \31998 );
xor \U$31623 ( \32000 , \8170 , \8172 );
xor \U$31624 ( \32001 , \32000 , \8193 );
and \U$31625 ( \32002 , \31981 , \32001 );
and \U$31626 ( \32003 , \31979 , \31981 );
or \U$31627 ( \32004 , \31999 , \32002 , \32003 );
not \U$31628 ( \32005 , \32004 );
not \U$31629 ( \32006 , \32005 );
and \U$31630 ( \32007 , \31996 , \32006 );
and \U$31631 ( \32008 , \31995 , \32005 );
nor \U$31632 ( \32009 , \32007 , \32008 );
xnor \U$31633 ( \32010 , \31993 , \32009 );
or \U$31634 ( \32011 , \31991 , \32010 );
or \U$31635 ( \32012 , \31993 , \32009 );
nand \U$31636 ( \32013 , \32011 , \32012 );
not \U$31637 ( \32014 , \31995 );
nor \U$31638 ( \32015 , \32014 , \32005 );
not \U$31639 ( \32016 , \8577 );
not \U$31640 ( \32017 , \8230 );
or \U$31641 ( \32018 , \32016 , \32017 );
or \U$31642 ( \32019 , \8230 , \8577 );
nand \U$31643 ( \32020 , \32018 , \32019 );
xor \U$31644 ( \32021 , \32015 , \32020 );
and \U$31645 ( \32022 , \32013 , \32021 );
and \U$31646 ( \32023 , \32020 , \32015 );
nor \U$31647 ( \32024 , \32022 , \32023 );
or \U$31648 ( \32025 , \8580 , \32024 );
nand \U$31649 ( \32026 , \8579 , \32025 );
and \U$31650 ( \32027 , \8215 , \32026 );
nor \U$31651 ( \32028 , \8214 , \32027 );
not \U$31652 ( \32029 , \32028 );
and \U$31653 ( \32030 , \7865 , \32029 );
nor \U$31654 ( \32031 , \7864 , \32030 );
not \U$31655 ( \32032 , \32031 );
xor \U$31656 ( \32033 , \7857 , \7859 );
and \U$31657 ( \32034 , \32033 , \7862 );
and \U$31658 ( \32035 , \7857 , \7859 );
or \U$31659 ( \32036 , \32034 , \32035 );
xor \U$31660 ( \32037 , \6857 , \6871 );
xor \U$31661 ( \32038 , \32037 , \6902 );
xor \U$31662 ( \32039 , \32036 , \32038 );
and \U$31663 ( \32040 , \32032 , \32039 );
and \U$31664 ( \32041 , \32036 , \32038 );
nor \U$31665 ( \32042 , \32040 , \32041 );
not \U$31666 ( \32043 , \32042 );
and \U$31667 ( \32044 , \6926 , \32043 );
nor \U$31668 ( \32045 , \6925 , \32044 );
xor \U$31669 ( \32046 , \6914 , \6916 );
and \U$31670 ( \32047 , \32046 , \6919 );
and \U$31671 ( \32048 , \6914 , \6916 );
or \U$31672 ( \32049 , \32047 , \32048 );
xor \U$31673 ( \32050 , \6049 , \6051 );
xor \U$31674 ( \32051 , \32050 , \6054 );
xor \U$31675 ( \32052 , \32049 , \32051 );
not \U$31676 ( \32053 , \32052 );
not \U$31677 ( \32054 , \6909 );
nand \U$31678 ( \32055 , \32054 , \6920 );
not \U$31679 ( \32056 , \32055 );
and \U$31680 ( \32057 , \32053 , \32056 );
and \U$31681 ( \32058 , \32052 , \32055 );
nor \U$31682 ( \32059 , \32057 , \32058 );
or \U$31683 ( \32060 , \32045 , \32059 );
not \U$31684 ( \32061 , \32052 );
or \U$31685 ( \32062 , \32055 , \32061 );
nand \U$31686 ( \32063 , \32060 , \32062 );
and \U$31687 ( \32064 , \32049 , \32051 );
not \U$31688 ( \32065 , \6057 );
not \U$31689 ( \32066 , \5784 );
or \U$31690 ( \32067 , \32065 , \32066 );
or \U$31691 ( \32068 , \5784 , \6057 );
nand \U$31692 ( \32069 , \32067 , \32068 );
xor \U$31693 ( \32070 , \32064 , \32069 );
and \U$31694 ( \32071 , \32063 , \32070 );
and \U$31695 ( \32072 , \32064 , \32069 );
nor \U$31696 ( \32073 , \32071 , \32072 );
or \U$31697 ( \32074 , \6060 , \32073 );
nand \U$31698 ( \32075 , \6059 , \32074 );
and \U$31699 ( \32076 , \5769 , \32075 );
nor \U$31700 ( \32077 , \5768 , \32076 );
or \U$31701 ( \32078 , \5500 , \32077 );
nand \U$31702 ( \32079 , \5499 , \32078 );
and \U$31703 ( \32080 , \5217 , \32079 );
nor \U$31704 ( \32081 , \5216 , \32080 );
not \U$31705 ( \32082 , \32081 );
and \U$31706 ( \32083 , \4926 , \4944 );
xor \U$31707 ( \32084 , \4928 , \4938 );
and \U$31708 ( \32085 , \32084 , \4943 );
and \U$31709 ( \32086 , \4928 , \4938 );
or \U$31710 ( \32087 , \32085 , \32086 );
not \U$31711 ( \32088 , \32087 );
xor \U$31712 ( \32089 , \4428 , \4430 );
xor \U$31713 ( \32090 , \32089 , \4433 );
not \U$31714 ( \32091 , \32090 );
or \U$31715 ( \32092 , \32088 , \32091 );
or \U$31716 ( \32093 , \32090 , \32087 );
nand \U$31717 ( \32094 , \32092 , \32093 );
xor \U$31718 ( \32095 , \32083 , \32094 );
and \U$31719 ( \32096 , \32082 , \32095 );
and \U$31720 ( \32097 , \32094 , \32083 );
nor \U$31721 ( \32098 , \32096 , \32097 );
not \U$31722 ( \32099 , \32090 );
nand \U$31723 ( \32100 , \32099 , \32087 );
not \U$31724 ( \32101 , \4199 );
not \U$31725 ( \32102 , \4436 );
and \U$31726 ( \32103 , \32101 , \32102 );
and \U$31727 ( \32104 , \4199 , \4436 );
nor \U$31728 ( \32105 , \32103 , \32104 );
xnor \U$31729 ( \32106 , \32100 , \32105 );
or \U$31730 ( \32107 , \32098 , \32106 );
or \U$31731 ( \32108 , \32100 , \32105 );
nand \U$31732 ( \32109 , \32107 , \32108 );
and \U$31733 ( \32110 , \4439 , \32109 );
nor \U$31734 ( \32111 , \4438 , \32110 );
or \U$31735 ( \32112 , \4184 , \32111 );
nand \U$31736 ( \32113 , \4183 , \32112 );
not \U$31737 ( \32114 , \3639 );
nor \U$31738 ( \32115 , \32114 , \3912 );
xor \U$31739 ( \32116 , \2937 , \3065 );
and \U$31740 ( \32117 , \32116 , \3120 );
and \U$31741 ( \32118 , \2937 , \3065 );
or \U$31742 ( \32119 , \32117 , \32118 );
and \U$31743 ( \32120 , \2408 , \2611 );
not \U$31744 ( \32121 , \2408 );
and \U$31745 ( \32122 , \32121 , \2397 );
nor \U$31746 ( \32123 , \32120 , \32122 );
not \U$31747 ( \32124 , \32123 );
not \U$31748 ( \32125 , \2394 );
and \U$31749 ( \32126 , \32124 , \32125 );
and \U$31750 ( \32127 , \32123 , \2394 );
nor \U$31751 ( \32128 , \32126 , \32127 );
xor \U$31752 ( \32129 , \2520 , \2521 );
xor \U$31753 ( \32130 , \32129 , \2552 );
xor \U$31754 ( \32131 , \32128 , \32130 );
xor \U$31755 ( \32132 , \2649 , \2651 );
xor \U$31756 ( \32133 , \32132 , \2662 );
xor \U$31757 ( \32134 , \32131 , \32133 );
not \U$31758 ( \32135 , \32134 );
xor \U$31759 ( \32136 , \3086 , \3094 );
and \U$31760 ( \32137 , \32136 , \3101 );
and \U$31761 ( \32138 , \3086 , \3094 );
or \U$31762 ( \32139 , \32137 , \32138 );
xor \U$31763 ( \32140 , \3072 , \2520 );
and \U$31764 ( \32141 , \32140 , \3079 );
and \U$31765 ( \32142 , \3072 , \2520 );
or \U$31766 ( \32143 , \32141 , \32142 );
xor \U$31767 ( \32144 , \32139 , \32143 );
xor \U$31768 ( \32145 , \3109 , \3115 );
and \U$31769 ( \32146 , \32145 , \3118 );
and \U$31770 ( \32147 , \3109 , \3115 );
or \U$31771 ( \32148 , \32146 , \32147 );
xor \U$31772 ( \32149 , \32144 , \32148 );
not \U$31773 ( \32150 , \32149 );
or \U$31774 ( \32151 , \32135 , \32150 );
or \U$31775 ( \32152 , \32134 , \32149 );
nand \U$31776 ( \32153 , \32151 , \32152 );
xor \U$31777 ( \32154 , \32119 , \32153 );
xor \U$31778 ( \32155 , \2581 , \2615 );
xor \U$31779 ( \32156 , \32155 , \2643 );
not \U$31780 ( \32157 , \32156 );
and \U$31781 ( \32158 , \3618 , \3612 );
not \U$31782 ( \32159 , \3618 );
not \U$31783 ( \32160 , \3612 );
and \U$31784 ( \32161 , \32159 , \32160 );
nor \U$31785 ( \32162 , \32161 , \3607 );
nor \U$31786 ( \32163 , \32158 , \32162 );
xor \U$31787 ( \32164 , \3080 , \3102 );
and \U$31788 ( \32165 , \32164 , \3119 );
and \U$31789 ( \32166 , \3080 , \3102 );
nor \U$31790 ( \32167 , \32165 , \32166 );
xor \U$31791 ( \32168 , \32163 , \32167 );
not \U$31792 ( \32169 , \32168 );
or \U$31793 ( \32170 , \32157 , \32169 );
or \U$31794 ( \32171 , \32168 , \32156 );
nand \U$31795 ( \32172 , \32170 , \32171 );
xor \U$31796 ( \32173 , \32154 , \32172 );
not \U$31797 ( \32174 , \32173 );
and \U$31798 ( \32175 , \3631 , \3121 );
not \U$31799 ( \32176 , \3631 );
not \U$31800 ( \32177 , \3121 );
and \U$31801 ( \32178 , \32176 , \32177 );
nor \U$31802 ( \32179 , \32178 , \3596 );
nor \U$31803 ( \32180 , \32175 , \32179 );
not \U$31804 ( \32181 , \32180 );
xor \U$31805 ( \32182 , \3603 , \3623 );
and \U$31806 ( \32183 , \32182 , \3630 );
and \U$31807 ( \32184 , \3603 , \3623 );
or \U$31808 ( \32185 , \32183 , \32184 );
not \U$31809 ( \32186 , \32185 );
and \U$31810 ( \32187 , \32181 , \32186 );
and \U$31811 ( \32188 , \32180 , \32185 );
nor \U$31812 ( \32189 , \32187 , \32188 );
not \U$31813 ( \32190 , \32189 );
or \U$31814 ( \32191 , \32174 , \32190 );
or \U$31815 ( \32192 , \32189 , \32173 );
nand \U$31816 ( \32193 , \32191 , \32192 );
xor \U$31817 ( \32194 , \32115 , \32193 );
and \U$31818 ( \32195 , \32113 , \32194 );
and \U$31819 ( \32196 , \32115 , \32193 );
nor \U$31820 ( \32197 , \32195 , \32196 );
xor \U$31821 ( \32198 , \32119 , \32153 );
and \U$31822 ( \32199 , \32198 , \32172 );
and \U$31823 ( \32200 , \32119 , \32153 );
or \U$31824 ( \32201 , \32199 , \32200 );
not \U$31825 ( \32202 , \32201 );
not \U$31826 ( \32203 , \32134 );
nand \U$31827 ( \32204 , \32203 , \32149 );
xor \U$31828 ( \32205 , \2555 , \2646 );
xor \U$31829 ( \32206 , \32205 , \2665 );
xor \U$31830 ( \32207 , \32204 , \32206 );
not \U$31831 ( \32208 , \32163 );
not \U$31832 ( \32209 , \32156 );
and \U$31833 ( \32210 , \32208 , \32209 );
and \U$31834 ( \32211 , \32163 , \32156 );
nor \U$31835 ( \32212 , \32211 , \32167 );
nor \U$31836 ( \32213 , \32210 , \32212 );
xor \U$31837 ( \32214 , \32207 , \32213 );
not \U$31838 ( \32215 , \32214 );
and \U$31839 ( \32216 , \32202 , \32215 );
and \U$31840 ( \32217 , \32201 , \32214 );
nor \U$31841 ( \32218 , \32216 , \32217 );
not \U$31842 ( \32219 , \32218 );
xor \U$31843 ( \32220 , \32128 , \32130 );
and \U$31844 ( \32221 , \32220 , \32133 );
and \U$31845 ( \32222 , \32128 , \32130 );
nor \U$31846 ( \32223 , \32221 , \32222 );
xor \U$31847 ( \32224 , \32139 , \32143 );
and \U$31848 ( \32225 , \32224 , \32148 );
and \U$31849 ( \32226 , \32139 , \32143 );
or \U$31850 ( \32227 , \32225 , \32226 );
xor \U$31851 ( \32228 , \32223 , \32227 );
xor \U$31852 ( \32229 , \2387 , \2410 );
xor \U$31853 ( \32230 , \32229 , \2438 );
xor \U$31854 ( \32231 , \2507 , \2514 );
xor \U$31855 ( \32232 , \32230 , \32231 );
xor \U$31856 ( \32233 , \32228 , \32232 );
not \U$31857 ( \32234 , \32233 );
and \U$31858 ( \32235 , \32219 , \32234 );
and \U$31859 ( \32236 , \32218 , \32233 );
nor \U$31860 ( \32237 , \32235 , \32236 );
and \U$31861 ( \32238 , \32173 , \32185 );
not \U$31862 ( \32239 , \32173 );
not \U$31863 ( \32240 , \32185 );
and \U$31864 ( \32241 , \32239 , \32240 );
nor \U$31865 ( \32242 , \32241 , \32180 );
nor \U$31866 ( \32243 , \32238 , \32242 );
xnor \U$31867 ( \32244 , \32237 , \32243 );
or \U$31868 ( \32245 , \32197 , \32244 );
or \U$31869 ( \32246 , \32237 , \32243 );
nand \U$31870 ( \32247 , \32245 , \32246 );
not \U$31871 ( \32248 , \32233 );
or \U$31872 ( \32249 , \32214 , \32248 );
not \U$31873 ( \32250 , \32248 );
not \U$31874 ( \32251 , \32214 );
or \U$31875 ( \32252 , \32250 , \32251 );
nand \U$31876 ( \32253 , \32252 , \32201 );
nand \U$31877 ( \32254 , \32249 , \32253 );
xor \U$31878 ( \32255 , \32204 , \32206 );
and \U$31879 ( \32256 , \32255 , \32213 );
and \U$31880 ( \32257 , \32204 , \32206 );
or \U$31881 ( \32258 , \32256 , \32257 );
not \U$31882 ( \32259 , \32258 );
xor \U$31883 ( \32260 , \32223 , \32227 );
and \U$31884 ( \32261 , \32260 , \32232 );
and \U$31885 ( \32262 , \32223 , \32227 );
or \U$31886 ( \32263 , \32261 , \32262 );
xor \U$31887 ( \32264 , \2441 , \2480 );
xor \U$31888 ( \32265 , \32264 , \2493 );
xor \U$31889 ( \32266 , \32263 , \32265 );
xor \U$31890 ( \32267 , \2519 , \2668 );
xor \U$31891 ( \32268 , \32267 , \2673 );
xor \U$31892 ( \32269 , \32266 , \32268 );
not \U$31893 ( \32270 , \32269 );
or \U$31894 ( \32271 , \32259 , \32270 );
or \U$31895 ( \32272 , \32269 , \32258 );
nand \U$31896 ( \32273 , \32271 , \32272 );
xor \U$31897 ( \32274 , \32254 , \32273 );
and \U$31898 ( \32275 , \32247 , \32274 );
and \U$31899 ( \32276 , \32254 , \32273 );
nor \U$31900 ( \32277 , \32275 , \32276 );
not \U$31901 ( \32278 , \32258 );
nand \U$31902 ( \32279 , \32278 , \32269 );
xor \U$31903 ( \32280 , \2676 , \2682 );
xor \U$31904 ( \32281 , \32280 , \2689 );
not \U$31905 ( \32282 , \32281 );
xor \U$31906 ( \32283 , \32263 , \32265 );
and \U$31907 ( \32284 , \32283 , \32268 );
and \U$31908 ( \32285 , \32263 , \32265 );
or \U$31909 ( \32286 , \32284 , \32285 );
not \U$31910 ( \32287 , \32286 );
and \U$31911 ( \32288 , \32282 , \32287 );
and \U$31912 ( \32289 , \32281 , \32286 );
nor \U$31913 ( \32290 , \32288 , \32289 );
xnor \U$31914 ( \32291 , \32279 , \32290 );
or \U$31915 ( \32292 , \32277 , \32291 );
or \U$31916 ( \32293 , \32279 , \32290 );
nand \U$31917 ( \32294 , \32292 , \32293 );
not \U$31918 ( \32295 , \32286 );
nor \U$31919 ( \32296 , \32295 , \32281 );
not \U$31920 ( \32297 , \2692 );
not \U$31921 ( \32298 , \2695 );
or \U$31922 ( \32299 , \32297 , \32298 );
or \U$31923 ( \32300 , \2695 , \2692 );
nand \U$31924 ( \32301 , \32299 , \32300 );
xor \U$31925 ( \32302 , \32296 , \32301 );
and \U$31926 ( \32303 , \32294 , \32302 );
and \U$31927 ( \32304 , \32296 , \32301 );
nor \U$31928 ( \32305 , \32303 , \32304 );
or \U$31929 ( \32306 , \2698 , \32305 );
nand \U$31930 ( \32307 , \2697 , \32306 );
not \U$31931 ( \32308 , \2334 );
nor \U$31932 ( \32309 , \32308 , \2501 );
and \U$31933 ( \32310 , \2172 , \2326 );
not \U$31934 ( \32311 , \2172 );
not \U$31935 ( \32312 , \2326 );
and \U$31936 ( \32313 , \32311 , \32312 );
nor \U$31937 ( \32314 , \32313 , \2323 );
nor \U$31938 ( \32315 , \32310 , \32314 );
not \U$31939 ( \32316 , \32315 );
xor \U$31940 ( \32317 , \2147 , \2149 );
xor \U$31941 ( \32318 , \32317 , \2152 );
not \U$31942 ( \32319 , \32318 );
or \U$31943 ( \32320 , \32316 , \32319 );
or \U$31944 ( \32321 , \32318 , \32315 );
nand \U$31945 ( \32322 , \32320 , \32321 );
xor \U$31946 ( \32323 , \32309 , \32322 );
and \U$31947 ( \32324 , \32307 , \32323 );
and \U$31948 ( \32325 , \32309 , \32322 );
nor \U$31949 ( \32326 , \32324 , \32325 );
not \U$31950 ( \32327 , \32315 );
nand \U$31951 ( \32328 , \32327 , \32318 );
not \U$31952 ( \32329 , \2162 );
not \U$31953 ( \32330 , \2155 );
and \U$31954 ( \32331 , \32329 , \32330 );
and \U$31955 ( \32332 , \2162 , \2155 );
nor \U$31956 ( \32333 , \32331 , \32332 );
xnor \U$31957 ( \32334 , \32328 , \32333 );
or \U$31958 ( \32335 , \32326 , \32334 );
or \U$31959 ( \32336 , \32328 , \32333 );
nand \U$31960 ( \32337 , \32335 , \32336 );
and \U$31961 ( \32338 , \2170 , \32337 );
nor \U$31962 ( \32339 , \2169 , \32338 );
or \U$31963 ( \32340 , \2011 , \32339 );
nand \U$31964 ( \32341 , \2010 , \32340 );
and \U$31965 ( \32342 , \1830 , \32341 );
nor \U$31966 ( \32343 , \1829 , \32342 );
not \U$31967 ( \32344 , \1824 );
nand \U$31968 ( \32345 , \32344 , \1819 );
not \U$31969 ( \32346 , \1328 );
not \U$31970 ( \32347 , \1447 );
and \U$31971 ( \32348 , \32346 , \32347 );
and \U$31972 ( \32349 , \1328 , \1447 );
nor \U$31973 ( \32350 , \32348 , \32349 );
xnor \U$31974 ( \32351 , \32345 , \32350 );
or \U$31975 ( \32352 , \32343 , \32351 );
or \U$31976 ( \32353 , \32345 , \32350 );
nand \U$31977 ( \32354 , \32352 , \32353 );
and \U$31978 ( \32355 , \1450 , \32354 );
nor \U$31979 ( \32356 , \1449 , \32355 );
or \U$31980 ( \32357 , \1321 , \32356 );
nand \U$31981 ( \32358 , \1320 , \32357 );
xor \U$31982 ( \32359 , \974 , \1078 );
not \U$31983 ( \32360 , \1195 );
nor \U$31984 ( \32361 , \32360 , \1091 );
xor \U$31985 ( \32362 , \32359 , \32361 );
and \U$31986 ( \32363 , \32358 , \32362 );
and \U$31987 ( \32364 , \32359 , \32361 );
nor \U$31988 ( \32365 , \32363 , \32364 );
not \U$31989 ( \32366 , \32365 );
and \U$31990 ( \32367 , \1081 , \32366 );
nor \U$31991 ( \32368 , \1080 , \32367 );
or \U$31992 ( \32369 , \954 , \32368 );
nand \U$31993 ( \32370 , \953 , \32369 );
and \U$31994 ( \32371 , \768 , \32370 );
nor \U$31995 ( \32372 , \767 , \32371 );
not \U$31996 ( \32373 , \762 );
nand \U$31997 ( \32374 , \32373 , \755 );
xor \U$31998 ( \32375 , \467 , \471 );
xor \U$31999 ( \32376 , \32375 , \480 );
not \U$32000 ( \32377 , \32376 );
xor \U$32001 ( \32378 , \727 , \728 );
and \U$32002 ( \32379 , \32378 , \753 );
and \U$32003 ( \32380 , \727 , \728 );
or \U$32004 ( \32381 , \32379 , \32380 );
not \U$32005 ( \32382 , \32381 );
or \U$32006 ( \32383 , \32377 , \32382 );
or \U$32007 ( \32384 , \32381 , \32376 );
nand \U$32008 ( \32385 , \32383 , \32384 );
not \U$32009 ( \32386 , \32385 );
not \U$32010 ( \32387 , \728 );
xor \U$32011 ( \32388 , \737 , \743 );
and \U$32012 ( \32389 , \32388 , \752 );
and \U$32013 ( \32390 , \737 , \743 );
or \U$32014 ( \32391 , \32389 , \32390 );
not \U$32015 ( \32392 , \32391 );
or \U$32016 ( \32393 , \32387 , \32392 );
or \U$32017 ( \32394 , \32391 , \728 );
nand \U$32018 ( \32395 , \32393 , \32394 );
not \U$32019 ( \32396 , \32395 );
nand \U$32020 ( \32397 , RIae76898_51, RIae78b48_125);
not \U$32021 ( \32398 , \32397 );
and \U$32022 ( \32399 , \32396 , \32398 );
and \U$32023 ( \32400 , \32395 , \32397 );
nor \U$32024 ( \32401 , \32399 , \32400 );
not \U$32025 ( \32402 , \32401 );
and \U$32026 ( \32403 , \32386 , \32402 );
and \U$32027 ( \32404 , \32385 , \32401 );
nor \U$32028 ( \32405 , \32403 , \32404 );
not \U$32029 ( \32406 , \32405 );
xor \U$32030 ( \32407 , \718 , \722 );
and \U$32031 ( \32408 , \32407 , \754 );
and \U$32032 ( \32409 , \718 , \722 );
or \U$32033 ( \32410 , \32408 , \32409 );
not \U$32034 ( \32411 , \32410 );
and \U$32035 ( \32412 , \32406 , \32411 );
and \U$32036 ( \32413 , \32405 , \32410 );
nor \U$32037 ( \32414 , \32412 , \32413 );
xnor \U$32038 ( \32415 , \32374 , \32414 );
or \U$32039 ( \32416 , \32372 , \32415 );
or \U$32040 ( \32417 , \32374 , \32414 );
nand \U$32041 ( \32418 , \32416 , \32417 );
not \U$32042 ( \32419 , \32410 );
nor \U$32043 ( \32420 , \32419 , \32405 );
or \U$32044 ( \32421 , \485 , \483 );
nand \U$32045 ( \32422 , \32421 , \486 );
or \U$32046 ( \32423 , \32401 , \32376 );
not \U$32047 ( \32424 , \32376 );
not \U$32048 ( \32425 , \32401 );
or \U$32049 ( \32426 , \32424 , \32425 );
nand \U$32050 ( \32427 , \32426 , \32381 );
nand \U$32051 ( \32428 , \32423 , \32427 );
xor \U$32052 ( \32429 , \32422 , \32428 );
or \U$32053 ( \32430 , \728 , \32397 );
not \U$32054 ( \32431 , \32397 );
not \U$32055 ( \32432 , \728 );
or \U$32056 ( \32433 , \32431 , \32432 );
nand \U$32057 ( \32434 , \32433 , \32391 );
nand \U$32058 ( \32435 , \32430 , \32434 );
xor \U$32059 ( \32436 , \32429 , \32435 );
xor \U$32060 ( \32437 , \32420 , \32436 );
and \U$32061 ( \32438 , \32418 , \32437 );
and \U$32062 ( \32439 , \32420 , \32436 );
nor \U$32063 ( \32440 , \32438 , \32439 );
not \U$32064 ( \32441 , \455 );
not \U$32065 ( \32442 , \486 );
or \U$32066 ( \32443 , \32441 , \32442 );
or \U$32067 ( \32444 , \486 , \455 );
nand \U$32068 ( \32445 , \32443 , \32444 );
not \U$32069 ( \32446 , \32445 );
not \U$32070 ( \32447 , \428 );
and \U$32071 ( \32448 , \32446 , \32447 );
and \U$32072 ( \32449 , \32445 , \428 );
nor \U$32073 ( \32450 , \32448 , \32449 );
xor \U$32074 ( \32451 , \32422 , \32428 );
and \U$32075 ( \32452 , \32451 , \32435 );
and \U$32076 ( \32453 , \32422 , \32428 );
nor \U$32077 ( \32454 , \32452 , \32453 );
xnor \U$32078 ( \32455 , \32450 , \32454 );
or \U$32079 ( \32456 , \32440 , \32455 );
or \U$32080 ( \32457 , \32450 , \32454 );
nand \U$32081 ( \32458 , \32456 , \32457 );
and \U$32082 ( \32459 , \489 , \32458 );
and \U$32083 ( \32460 , \488 , \418 );
and \U$32084 ( \32461 , \398 , \417 );
nor \U$32085 ( \32462 , \32459 , \32460 , \32461 );
not \U$32086 ( \32463 , \32462 );
nand \U$32087 ( \32464 , RIae78e18_131, RIae78b48_125);
not \U$32088 ( \32465 , \32464 );
nand \U$32089 ( \32466 , RIae78d28_129, RIae78b48_125);
nand \U$32090 ( \32467 , RIae78e18_131, \384 );
not \U$32091 ( \32468 , \32467 );
not \U$32092 ( \32469 , \388 );
and \U$32093 ( \32470 , \32468 , \32469 );
and \U$32094 ( \32471 , \32467 , \392 );
nor \U$32095 ( \32472 , \32470 , \32471 );
nand \U$32096 ( \32473 , \32466 , \32472 );
not \U$32097 ( \32474 , \32473 );
or \U$32098 ( \32475 , \32465 , \32474 );
or \U$32099 ( \32476 , \32473 , \32464 );
nand \U$32100 ( \32477 , \32475 , \32476 );
not \U$32101 ( \32478 , \32477 );
and \U$32102 ( \32479 , \32463 , \32478 );
and \U$32103 ( \32480 , \32462 , \32477 );
nor \U$32104 ( \32481 , \32479 , \32480 );
not \U$32105 ( \32482 , \32481 );
or \U$32106 ( \32483 , \32472 , \32466 );
nand \U$32107 ( \32484 , \32483 , \32473 );
nand \U$32108 ( \32485 , RIae78ad0_124, RIae78b48_125);
or \U$32109 ( \32486 , \400 , \32485 );
not \U$32110 ( \32487 , \32485 );
not \U$32111 ( \32488 , \402 );
or \U$32112 ( \32489 , \32487 , \32488 );
not \U$32113 ( \32490 , \388 );
and \U$32114 ( \32491 , \384 , RIae78d28_129);
and \U$32115 ( \32492 , RIae78e18_131, \382 );
nor \U$32116 ( \32493 , \32491 , \32492 );
not \U$32117 ( \32494 , \32493 );
or \U$32118 ( \32495 , \32490 , \32494 );
or \U$32119 ( \32496 , \32493 , \388 );
nand \U$32120 ( \32497 , \32495 , \32496 );
nand \U$32121 ( \32498 , \32489 , \32497 );
nand \U$32122 ( \32499 , \32486 , \32498 );
xor \U$32123 ( \32500 , \32484 , \32499 );
not \U$32124 ( \32501 , \402 );
not \U$32125 ( \32502 , \32497 );
or \U$32126 ( \32503 , \32501 , \32502 );
or \U$32127 ( \32504 , \32497 , \400 );
nand \U$32128 ( \32505 , \32503 , \32504 );
not \U$32129 ( \32506 , \32505 );
not \U$32130 ( \32507 , \32485 );
and \U$32131 ( \32508 , \32506 , \32507 );
and \U$32132 ( \32509 , \32505 , \32485 );
nor \U$32133 ( \32510 , \32508 , \32509 );
nand \U$32134 ( \32511 , RIae78e18_131, \436 );
not \U$32135 ( \32512 , \32511 );
not \U$32136 ( \32513 , \400 );
and \U$32137 ( \32514 , \32512 , \32513 );
and \U$32138 ( \32515 , \32511 , \400 );
nor \U$32139 ( \32516 , \32514 , \32515 );
nand \U$32140 ( \32517 , RIae76be0_58, RIae78b48_125);
xor \U$32141 ( \32518 , \32516 , \32517 );
and \U$32142 ( \32519 , \384 , RIae78ad0_124);
and \U$32143 ( \32520 , RIae78d28_129, \382 );
nor \U$32144 ( \32521 , \32519 , \32520 );
not \U$32145 ( \32522 , \32521 );
not \U$32146 ( \32523 , \392 );
and \U$32147 ( \32524 , \32522 , \32523 );
and \U$32148 ( \32525 , \32521 , \388 );
nor \U$32149 ( \32526 , \32524 , \32525 );
and \U$32150 ( \32527 , \32518 , \32526 );
and \U$32151 ( \32528 , \32516 , \32517 );
or \U$32152 ( \32529 , \32527 , \32528 );
or \U$32153 ( \32530 , \32510 , \32529 );
not \U$32154 ( \32531 , \32529 );
not \U$32155 ( \32532 , \32510 );
or \U$32156 ( \32533 , \32531 , \32532 );
and \U$32157 ( \32534 , \384 , RIae76be0_58);
and \U$32158 ( \32535 , RIae78ad0_124, \382 );
nor \U$32159 ( \32536 , \32534 , \32535 );
not \U$32160 ( \32537 , \32536 );
not \U$32161 ( \32538 , \392 );
and \U$32162 ( \32539 , \32537 , \32538 );
and \U$32163 ( \32540 , \32536 , \388 );
nor \U$32164 ( \32541 , \32539 , \32540 );
xor \U$32165 ( \32542 , \32541 , \471 );
and \U$32166 ( \32543 , \436 , RIae78d28_129);
and \U$32167 ( \32544 , RIae78e18_131, \434 );
nor \U$32168 ( \32545 , \32543 , \32544 );
not \U$32169 ( \32546 , \32545 );
not \U$32170 ( \32547 , \402 );
and \U$32171 ( \32548 , \32546 , \32547 );
and \U$32172 ( \32549 , \32545 , \402 );
nor \U$32173 ( \32550 , \32548 , \32549 );
and \U$32174 ( \32551 , \32542 , \32550 );
and \U$32175 ( \32552 , \32541 , \471 );
or \U$32176 ( \32553 , \32551 , \32552 );
xor \U$32177 ( \32554 , \32516 , \32517 );
xor \U$32178 ( \32555 , \32554 , \32526 );
nand \U$32179 ( \32556 , \32553 , \32555 );
nand \U$32180 ( \32557 , \32533 , \32556 );
nand \U$32181 ( \32558 , \32530 , \32557 );
xor \U$32182 ( \32559 , \32500 , \32558 );
xor \U$32183 ( \32560 , \32541 , \471 );
xor \U$32184 ( \32561 , \32560 , \32550 );
not \U$32185 ( \32562 , \32561 );
not \U$32186 ( \32563 , \402 );
and \U$32187 ( \32564 , \436 , RIae76be0_58);
and \U$32188 ( \32565 , RIae78ad0_124, \434 );
nor \U$32189 ( \32566 , \32564 , \32565 );
not \U$32190 ( \32567 , \32566 );
or \U$32191 ( \32568 , \32563 , \32567 );
or \U$32192 ( \32569 , \32566 , \402 );
nand \U$32193 ( \32570 , \32568 , \32569 );
xor \U$32194 ( \32571 , \32570 , \504 );
not \U$32195 ( \32572 , \471 );
and \U$32196 ( \32573 , \514 , RIae78d28_129);
and \U$32197 ( \32574 , RIae78e18_131, \512 );
nor \U$32198 ( \32575 , \32573 , \32574 );
not \U$32199 ( \32576 , \32575 );
or \U$32200 ( \32577 , \32572 , \32576 );
or \U$32201 ( \32578 , \32575 , \469 );
nand \U$32202 ( \32579 , \32577 , \32578 );
and \U$32203 ( \32580 , \32571 , \32579 );
and \U$32204 ( \32581 , \32570 , \504 );
or \U$32205 ( \32582 , \32580 , \32581 );
nand \U$32206 ( \32583 , RIae76820_50, RIae78b48_125);
xor \U$32207 ( \32584 , \32582 , \32583 );
not \U$32208 ( \32585 , \392 );
and \U$32209 ( \32586 , \384 , RIae76910_52);
and \U$32210 ( \32587 , RIae76be0_58, \382 );
nor \U$32211 ( \32588 , \32586 , \32587 );
not \U$32212 ( \32589 , \32588 );
or \U$32213 ( \32590 , \32585 , \32589 );
or \U$32214 ( \32591 , \32588 , \388 );
nand \U$32215 ( \32592 , \32590 , \32591 );
not \U$32216 ( \32593 , \471 );
nand \U$32217 ( \32594 , RIae78e18_131, \514 );
not \U$32218 ( \32595 , \32594 );
or \U$32219 ( \32596 , \32593 , \32595 );
or \U$32220 ( \32597 , \32594 , \469 );
nand \U$32221 ( \32598 , \32596 , \32597 );
xor \U$32222 ( \32599 , \32592 , \32598 );
not \U$32223 ( \32600 , \400 );
and \U$32224 ( \32601 , \436 , RIae78ad0_124);
and \U$32225 ( \32602 , RIae78d28_129, \434 );
nor \U$32226 ( \32603 , \32601 , \32602 );
not \U$32227 ( \32604 , \32603 );
or \U$32228 ( \32605 , \32600 , \32604 );
or \U$32229 ( \32606 , \32603 , \400 );
nand \U$32230 ( \32607 , \32605 , \32606 );
xor \U$32231 ( \32608 , \32599 , \32607 );
and \U$32232 ( \32609 , \32584 , \32608 );
and \U$32233 ( \32610 , \32582 , \32583 );
or \U$32234 ( \32611 , \32609 , \32610 );
not \U$32235 ( \32612 , \32611 );
or \U$32236 ( \32613 , \32562 , \32612 );
or \U$32237 ( \32614 , \32611 , \32561 );
nand \U$32238 ( \32615 , \32613 , \32614 );
not \U$32239 ( \32616 , \32615 );
not \U$32240 ( \32617 , \32583 );
xor \U$32241 ( \32618 , \32592 , \32598 );
and \U$32242 ( \32619 , \32618 , \32607 );
and \U$32243 ( \32620 , \32592 , \32598 );
or \U$32244 ( \32621 , \32619 , \32620 );
not \U$32245 ( \32622 , \32621 );
or \U$32246 ( \32623 , \32617 , \32622 );
or \U$32247 ( \32624 , \32621 , \32583 );
nand \U$32248 ( \32625 , \32623 , \32624 );
not \U$32249 ( \32626 , \32625 );
nand \U$32250 ( \32627 , RIae76910_52, RIae78b48_125);
not \U$32251 ( \32628 , \32627 );
and \U$32252 ( \32629 , \32626 , \32628 );
and \U$32253 ( \32630 , \32625 , \32627 );
nor \U$32254 ( \32631 , \32629 , \32630 );
not \U$32255 ( \32632 , \32631 );
and \U$32256 ( \32633 , \32616 , \32632 );
and \U$32257 ( \32634 , \32615 , \32631 );
nor \U$32258 ( \32635 , \32633 , \32634 );
not \U$32259 ( \32636 , \32635 );
not \U$32260 ( \32637 , RIae76a00_54);
nor \U$32261 ( \32638 , \32637 , \491 );
xor \U$32262 ( \32639 , \32570 , \504 );
xor \U$32263 ( \32640 , \32639 , \32579 );
and \U$32264 ( \32641 , \32638 , \32640 );
nand \U$32265 ( \32642 , RIae76af0_56, RIae78b48_125);
and \U$32266 ( \32643 , \384 , RIae76a00_54);
and \U$32267 ( \32644 , RIae76820_50, \382 );
nor \U$32268 ( \32645 , \32643 , \32644 );
not \U$32269 ( \32646 , \32645 );
not \U$32270 ( \32647 , \388 );
and \U$32271 ( \32648 , \32646 , \32647 );
and \U$32272 ( \32649 , \32645 , \388 );
nor \U$32273 ( \32650 , \32648 , \32649 );
nand \U$32274 ( \32651 , \32642 , \32650 );
not \U$32275 ( \32652 , \388 );
and \U$32276 ( \32653 , \384 , RIae76820_50);
and \U$32277 ( \32654 , RIae76910_52, \382 );
nor \U$32278 ( \32655 , \32653 , \32654 );
not \U$32279 ( \32656 , \32655 );
or \U$32280 ( \32657 , \32652 , \32656 );
or \U$32281 ( \32658 , \32655 , \388 );
nand \U$32282 ( \32659 , \32657 , \32658 );
xor \U$32283 ( \32660 , \32651 , \32659 );
not \U$32284 ( \32661 , \400 );
and \U$32285 ( \32662 , \436 , RIae76910_52);
and \U$32286 ( \32663 , RIae76be0_58, \434 );
nor \U$32287 ( \32664 , \32662 , \32663 );
not \U$32288 ( \32665 , \32664 );
or \U$32289 ( \32666 , \32661 , \32665 );
or \U$32290 ( \32667 , \32664 , \400 );
nand \U$32291 ( \32668 , \32666 , \32667 );
nand \U$32292 ( \32669 , RIae78e18_131, \558 );
and \U$32293 ( \32670 , \32669 , \504 );
not \U$32294 ( \32671 , \32669 );
and \U$32295 ( \32672 , \32671 , \562 );
nor \U$32296 ( \32673 , \32670 , \32672 );
xor \U$32297 ( \32674 , \32668 , \32673 );
not \U$32298 ( \32675 , \471 );
and \U$32299 ( \32676 , \514 , RIae78ad0_124);
and \U$32300 ( \32677 , RIae78d28_129, \512 );
nor \U$32301 ( \32678 , \32676 , \32677 );
not \U$32302 ( \32679 , \32678 );
or \U$32303 ( \32680 , \32675 , \32679 );
or \U$32304 ( \32681 , \32678 , \471 );
nand \U$32305 ( \32682 , \32680 , \32681 );
and \U$32306 ( \32683 , \32674 , \32682 );
and \U$32307 ( \32684 , \32668 , \32673 );
or \U$32308 ( \32685 , \32683 , \32684 );
and \U$32309 ( \32686 , \32660 , \32685 );
and \U$32310 ( \32687 , \32651 , \32659 );
or \U$32311 ( \32688 , \32686 , \32687 );
xor \U$32312 ( \32689 , \32641 , \32688 );
xor \U$32313 ( \32690 , \32582 , \32583 );
xor \U$32314 ( \32691 , \32690 , \32608 );
and \U$32315 ( \32692 , \32689 , \32691 );
and \U$32316 ( \32693 , \32641 , \32688 );
or \U$32317 ( \32694 , \32692 , \32693 );
not \U$32318 ( \32695 , \32694 );
and \U$32319 ( \32696 , \32636 , \32695 );
and \U$32320 ( \32697 , \32635 , \32694 );
nor \U$32321 ( \32698 , \32696 , \32697 );
xor \U$32322 ( \32699 , \32651 , \32659 );
xor \U$32323 ( \32700 , \32699 , \32685 );
xor \U$32324 ( \32701 , \32638 , \32640 );
and \U$32325 ( \32702 , \32700 , \32701 );
not \U$32326 ( \32703 , \32700 );
not \U$32327 ( \32704 , \32701 );
and \U$32328 ( \32705 , \32703 , \32704 );
and \U$32329 ( \32706 , \558 , RIae78d28_129);
and \U$32330 ( \32707 , RIae78e18_131, \556 );
nor \U$32331 ( \32708 , \32706 , \32707 );
and \U$32332 ( \32709 , \32708 , \504 );
not \U$32333 ( \32710 , \32708 );
and \U$32334 ( \32711 , \32710 , \562 );
nor \U$32335 ( \32712 , \32709 , \32711 );
xor \U$32336 ( \32713 , \32712 , \588 );
not \U$32337 ( \32714 , \471 );
and \U$32338 ( \32715 , \514 , RIae76be0_58);
and \U$32339 ( \32716 , RIae78ad0_124, \512 );
nor \U$32340 ( \32717 , \32715 , \32716 );
not \U$32341 ( \32718 , \32717 );
or \U$32342 ( \32719 , \32714 , \32718 );
or \U$32343 ( \32720 , \32717 , \471 );
nand \U$32344 ( \32721 , \32719 , \32720 );
and \U$32345 ( \32722 , \32713 , \32721 );
and \U$32346 ( \32723 , \32712 , \588 );
or \U$32347 ( \32724 , \32722 , \32723 );
and \U$32348 ( \32725 , \384 , RIae76af0_56);
and \U$32349 ( \32726 , RIae76a00_54, \382 );
nor \U$32350 ( \32727 , \32725 , \32726 );
not \U$32351 ( \32728 , \32727 );
not \U$32352 ( \32729 , \392 );
and \U$32353 ( \32730 , \32728 , \32729 );
and \U$32354 ( \32731 , \32727 , \392 );
nor \U$32355 ( \32732 , \32730 , \32731 );
nand \U$32356 ( \32733 , RIae76280_38, RIae78b48_125);
or \U$32357 ( \32734 , \32732 , \32733 );
not \U$32358 ( \32735 , \32733 );
not \U$32359 ( \32736 , \32732 );
or \U$32360 ( \32737 , \32735 , \32736 );
not \U$32361 ( \32738 , \402 );
and \U$32362 ( \32739 , \436 , RIae76820_50);
and \U$32363 ( \32740 , RIae76910_52, \434 );
nor \U$32364 ( \32741 , \32739 , \32740 );
not \U$32365 ( \32742 , \32741 );
or \U$32366 ( \32743 , \32738 , \32742 );
or \U$32367 ( \32744 , \32741 , \402 );
nand \U$32368 ( \32745 , \32743 , \32744 );
nand \U$32369 ( \32746 , \32737 , \32745 );
nand \U$32370 ( \32747 , \32734 , \32746 );
xor \U$32371 ( \32748 , \32724 , \32747 );
or \U$32372 ( \32749 , \32650 , \32642 );
nand \U$32373 ( \32750 , \32749 , \32651 );
and \U$32374 ( \32751 , \32748 , \32750 );
and \U$32375 ( \32752 , \32724 , \32747 );
nor \U$32376 ( \32753 , \32751 , \32752 );
nor \U$32377 ( \32754 , \32705 , \32753 );
nor \U$32378 ( \32755 , \32702 , \32754 );
not \U$32379 ( \32756 , \32755 );
xor \U$32380 ( \32757 , \32641 , \32688 );
xor \U$32381 ( \32758 , \32757 , \32691 );
nand \U$32382 ( \32759 , \32756 , \32758 );
or \U$32383 ( \32760 , \32698 , \32759 );
xnor \U$32384 ( \32761 , \32759 , \32698 );
not \U$32385 ( \32762 , \32701 );
not \U$32386 ( \32763 , \32700 );
not \U$32387 ( \32764 , \32753 );
and \U$32388 ( \32765 , \32763 , \32764 );
and \U$32389 ( \32766 , \32700 , \32753 );
nor \U$32390 ( \32767 , \32765 , \32766 );
not \U$32391 ( \32768 , \32767 );
or \U$32392 ( \32769 , \32762 , \32768 );
or \U$32393 ( \32770 , \32767 , \32701 );
nand \U$32394 ( \32771 , \32769 , \32770 );
not \U$32395 ( \32772 , \32771 );
xor \U$32396 ( \32773 , \32724 , \32747 );
xor \U$32397 ( \32774 , \32773 , \32750 );
xor \U$32398 ( \32775 , \32668 , \32673 );
xor \U$32399 ( \32776 , \32775 , \32682 );
and \U$32400 ( \32777 , \32774 , \32776 );
not \U$32401 ( \32778 , \32774 );
not \U$32402 ( \32779 , \32776 );
and \U$32403 ( \32780 , \32778 , \32779 );
and \U$32404 ( \32781 , \514 , RIae76910_52);
and \U$32405 ( \32782 , RIae76be0_58, \512 );
nor \U$32406 ( \32783 , \32781 , \32782 );
not \U$32407 ( \32784 , \32783 );
not \U$32408 ( \32785 , \471 );
and \U$32409 ( \32786 , \32784 , \32785 );
and \U$32410 ( \32787 , \32783 , \471 );
nor \U$32411 ( \32788 , \32786 , \32787 );
and \U$32412 ( \32789 , \558 , RIae78ad0_124);
and \U$32413 ( \32790 , RIae78d28_129, \556 );
nor \U$32414 ( \32791 , \32789 , \32790 );
and \U$32415 ( \32792 , \32791 , \562 );
not \U$32416 ( \32793 , \32791 );
and \U$32417 ( \32794 , \32793 , \504 );
nor \U$32418 ( \32795 , \32792 , \32794 );
or \U$32419 ( \32796 , \32788 , \32795 );
not \U$32420 ( \32797 , \32795 );
not \U$32421 ( \32798 , \32788 );
or \U$32422 ( \32799 , \32797 , \32798 );
nand \U$32423 ( \32800 , RIae78e18_131, \672 );
and \U$32424 ( \32801 , \32800 , \588 );
not \U$32425 ( \32802 , \32800 );
and \U$32426 ( \32803 , \32802 , \587 );
nor \U$32427 ( \32804 , \32801 , \32803 );
nand \U$32428 ( \32805 , \32799 , \32804 );
nand \U$32429 ( \32806 , \32796 , \32805 );
and \U$32430 ( \32807 , \436 , RIae76a00_54);
and \U$32431 ( \32808 , RIae76820_50, \434 );
nor \U$32432 ( \32809 , \32807 , \32808 );
not \U$32433 ( \32810 , \32809 );
not \U$32434 ( \32811 , \402 );
and \U$32435 ( \32812 , \32810 , \32811 );
and \U$32436 ( \32813 , \32809 , \402 );
nor \U$32437 ( \32814 , \32812 , \32813 );
nand \U$32438 ( \32815 , RIae76370_40, RIae78b48_125);
or \U$32439 ( \32816 , \32814 , \32815 );
not \U$32440 ( \32817 , \32815 );
not \U$32441 ( \32818 , \32814 );
or \U$32442 ( \32819 , \32817 , \32818 );
not \U$32443 ( \32820 , \392 );
and \U$32444 ( \32821 , \384 , RIae76280_38);
and \U$32445 ( \32822 , RIae76af0_56, \382 );
nor \U$32446 ( \32823 , \32821 , \32822 );
not \U$32447 ( \32824 , \32823 );
or \U$32448 ( \32825 , \32820 , \32824 );
or \U$32449 ( \32826 , \32823 , \392 );
nand \U$32450 ( \32827 , \32825 , \32826 );
nand \U$32451 ( \32828 , \32819 , \32827 );
nand \U$32452 ( \32829 , \32816 , \32828 );
and \U$32453 ( \32830 , \32806 , \32829 );
not \U$32454 ( \32831 , \32806 );
not \U$32455 ( \32832 , \32829 );
and \U$32456 ( \32833 , \32831 , \32832 );
not \U$32457 ( \32834 , \32732 );
not \U$32458 ( \32835 , \32745 );
or \U$32459 ( \32836 , \32834 , \32835 );
or \U$32460 ( \32837 , \32732 , \32745 );
nand \U$32461 ( \32838 , \32836 , \32837 );
not \U$32462 ( \32839 , \32838 );
not \U$32463 ( \32840 , \32733 );
and \U$32464 ( \32841 , \32839 , \32840 );
and \U$32465 ( \32842 , \32838 , \32733 );
nor \U$32466 ( \32843 , \32841 , \32842 );
nor \U$32467 ( \32844 , \32833 , \32843 );
nor \U$32468 ( \32845 , \32830 , \32844 );
nor \U$32469 ( \32846 , \32780 , \32845 );
nor \U$32470 ( \32847 , \32777 , \32846 );
nor \U$32471 ( \32848 , \32772 , \32847 );
not \U$32472 ( \32849 , \32758 );
not \U$32473 ( \32850 , \32755 );
or \U$32474 ( \32851 , \32849 , \32850 );
or \U$32475 ( \32852 , \32755 , \32758 );
nand \U$32476 ( \32853 , \32851 , \32852 );
and \U$32477 ( \32854 , \32848 , \32853 );
xor \U$32478 ( \32855 , \32848 , \32853 );
not \U$32479 ( \32856 , \32774 );
not \U$32480 ( \32857 , \32845 );
not \U$32481 ( \32858 , \32776 );
and \U$32482 ( \32859 , \32857 , \32858 );
and \U$32483 ( \32860 , \32845 , \32776 );
nor \U$32484 ( \32861 , \32859 , \32860 );
not \U$32485 ( \32862 , \32861 );
or \U$32486 ( \32863 , \32856 , \32862 );
or \U$32487 ( \32864 , \32861 , \32774 );
nand \U$32488 ( \32865 , \32863 , \32864 );
and \U$32489 ( \32866 , \672 , RIae78d28_129);
and \U$32490 ( \32867 , RIae78e18_131, \670 );
nor \U$32491 ( \32868 , \32866 , \32867 );
and \U$32492 ( \32869 , \32868 , \587 );
not \U$32493 ( \32870 , \32868 );
and \U$32494 ( \32871 , \32870 , \588 );
nor \U$32495 ( \32872 , \32869 , \32871 );
xor \U$32496 ( \32873 , \32872 , \787 );
and \U$32497 ( \32874 , \558 , RIae76be0_58);
and \U$32498 ( \32875 , RIae78ad0_124, \556 );
nor \U$32499 ( \32876 , \32874 , \32875 );
and \U$32500 ( \32877 , \32876 , \562 );
not \U$32501 ( \32878 , \32876 );
and \U$32502 ( \32879 , \32878 , \504 );
nor \U$32503 ( \32880 , \32877 , \32879 );
and \U$32504 ( \32881 , \32873 , \32880 );
and \U$32505 ( \32882 , \32872 , \787 );
or \U$32506 ( \32883 , \32881 , \32882 );
and \U$32507 ( \32884 , \436 , RIae76af0_56);
and \U$32508 ( \32885 , RIae76a00_54, \434 );
nor \U$32509 ( \32886 , \32884 , \32885 );
not \U$32510 ( \32887 , \32886 );
not \U$32511 ( \32888 , \400 );
and \U$32512 ( \32889 , \32887 , \32888 );
and \U$32513 ( \32890 , \32886 , \400 );
nor \U$32514 ( \32891 , \32889 , \32890 );
and \U$32515 ( \32892 , \384 , RIae76370_40);
and \U$32516 ( \32893 , RIae76280_38, \382 );
nor \U$32517 ( \32894 , \32892 , \32893 );
not \U$32518 ( \32895 , \32894 );
not \U$32519 ( \32896 , \392 );
and \U$32520 ( \32897 , \32895 , \32896 );
and \U$32521 ( \32898 , \32894 , \392 );
nor \U$32522 ( \32899 , \32897 , \32898 );
xor \U$32523 ( \32900 , \32891 , \32899 );
and \U$32524 ( \32901 , \514 , RIae76820_50);
and \U$32525 ( \32902 , RIae76910_52, \512 );
nor \U$32526 ( \32903 , \32901 , \32902 );
not \U$32527 ( \32904 , \32903 );
not \U$32528 ( \32905 , \469 );
and \U$32529 ( \32906 , \32904 , \32905 );
and \U$32530 ( \32907 , \32903 , \471 );
nor \U$32531 ( \32908 , \32906 , \32907 );
and \U$32532 ( \32909 , \32900 , \32908 );
and \U$32533 ( \32910 , \32891 , \32899 );
or \U$32534 ( \32911 , \32909 , \32910 );
nand \U$32535 ( \32912 , \32883 , \32911 );
xor \U$32536 ( \32913 , \32712 , \588 );
xor \U$32537 ( \32914 , \32913 , \32721 );
xor \U$32538 ( \32915 , \32912 , \32914 );
not \U$32539 ( \32916 , \32843 );
xor \U$32540 ( \32917 , \32806 , \32829 );
not \U$32541 ( \32918 , \32917 );
or \U$32542 ( \32919 , \32916 , \32918 );
or \U$32543 ( \32920 , \32917 , \32843 );
nand \U$32544 ( \32921 , \32919 , \32920 );
and \U$32545 ( \32922 , \32915 , \32921 );
and \U$32546 ( \32923 , \32912 , \32914 );
or \U$32547 ( \32924 , \32922 , \32923 );
and \U$32548 ( \32925 , \32865 , \32924 );
not \U$32549 ( \32926 , \32865 );
not \U$32550 ( \32927 , \32924 );
and \U$32551 ( \32928 , \32926 , \32927 );
xor \U$32552 ( \32929 , \32912 , \32914 );
xor \U$32553 ( \32930 , \32929 , \32921 );
or \U$32554 ( \32931 , \32911 , \32883 );
nand \U$32555 ( \32932 , \32931 , \32912 );
not \U$32556 ( \32933 , \32932 );
not \U$32557 ( \32934 , \32804 );
not \U$32558 ( \32935 , \32795 );
or \U$32559 ( \32936 , \32934 , \32935 );
or \U$32560 ( \32937 , \32795 , \32804 );
nand \U$32561 ( \32938 , \32936 , \32937 );
not \U$32562 ( \32939 , \32938 );
not \U$32563 ( \32940 , \32788 );
and \U$32564 ( \32941 , \32939 , \32940 );
and \U$32565 ( \32942 , \32938 , \32788 );
nor \U$32566 ( \32943 , \32941 , \32942 );
nor \U$32567 ( \32944 , \32933 , \32943 );
and \U$32568 ( \32945 , \32930 , \32944 );
not \U$32569 ( \32946 , \32930 );
not \U$32570 ( \32947 , \32944 );
and \U$32571 ( \32948 , \32946 , \32947 );
not \U$32572 ( \32949 , \469 );
and \U$32573 ( \32950 , \514 , RIae76a00_54);
and \U$32574 ( \32951 , RIae76820_50, \512 );
nor \U$32575 ( \32952 , \32950 , \32951 );
not \U$32576 ( \32953 , \32952 );
or \U$32577 ( \32954 , \32949 , \32953 );
or \U$32578 ( \32955 , \32952 , \469 );
nand \U$32579 ( \32956 , \32954 , \32955 );
not \U$32580 ( \32957 , \392 );
and \U$32581 ( \32958 , \384 , RIae760a0_34);
and \U$32582 ( \32959 , RIae76370_40, \382 );
nor \U$32583 ( \32960 , \32958 , \32959 );
not \U$32584 ( \32961 , \32960 );
or \U$32585 ( \32962 , \32957 , \32961 );
or \U$32586 ( \32963 , \32960 , \392 );
nand \U$32587 ( \32964 , \32962 , \32963 );
xor \U$32588 ( \32965 , \32956 , \32964 );
not \U$32589 ( \32966 , \402 );
and \U$32590 ( \32967 , \436 , RIae76280_38);
and \U$32591 ( \32968 , RIae76af0_56, \434 );
nor \U$32592 ( \32969 , \32967 , \32968 );
not \U$32593 ( \32970 , \32969 );
or \U$32594 ( \32971 , \32966 , \32970 );
or \U$32595 ( \32972 , \32969 , \400 );
nand \U$32596 ( \32973 , \32971 , \32972 );
and \U$32597 ( \32974 , \32965 , \32973 );
and \U$32598 ( \32975 , \32956 , \32964 );
or \U$32599 ( \32976 , \32974 , \32975 );
and \U$32600 ( \32977 , \558 , RIae76910_52);
and \U$32601 ( \32978 , RIae76be0_58, \556 );
nor \U$32602 ( \32979 , \32977 , \32978 );
and \U$32603 ( \32980 , \32979 , \504 );
not \U$32604 ( \32981 , \32979 );
and \U$32605 ( \32982 , \32981 , \562 );
nor \U$32606 ( \32983 , \32980 , \32982 );
not \U$32607 ( \32984 , \787 );
nand \U$32608 ( \32985 , RIae78e18_131, \883 );
not \U$32609 ( \32986 , \32985 );
or \U$32610 ( \32987 , \32984 , \32986 );
or \U$32611 ( \32988 , \32985 , \789 );
nand \U$32612 ( \32989 , \32987 , \32988 );
xor \U$32613 ( \32990 , \32983 , \32989 );
and \U$32614 ( \32991 , \672 , RIae78ad0_124);
and \U$32615 ( \32992 , RIae78d28_129, \670 );
nor \U$32616 ( \32993 , \32991 , \32992 );
and \U$32617 ( \32994 , \32993 , \588 );
not \U$32618 ( \32995 , \32993 );
and \U$32619 ( \32996 , \32995 , \587 );
nor \U$32620 ( \32997 , \32994 , \32996 );
and \U$32621 ( \32998 , \32990 , \32997 );
and \U$32622 ( \32999 , \32983 , \32989 );
or \U$32623 ( \33000 , \32998 , \32999 );
xor \U$32624 ( \33001 , \32976 , \33000 );
nand \U$32625 ( \33002 , RIae76190_36, RIae78b48_125);
not \U$32626 ( \33003 , \33002 );
and \U$32627 ( \33004 , \33001 , \33003 );
and \U$32628 ( \33005 , \32976 , \33000 );
or \U$32629 ( \33006 , \33004 , \33005 );
not \U$32630 ( \33007 , \33006 );
not \U$32631 ( \33008 , \32814 );
not \U$32632 ( \33009 , \32827 );
or \U$32633 ( \33010 , \33008 , \33009 );
or \U$32634 ( \33011 , \32814 , \32827 );
nand \U$32635 ( \33012 , \33010 , \33011 );
not \U$32636 ( \33013 , \33012 );
not \U$32637 ( \33014 , \32815 );
and \U$32638 ( \33015 , \33013 , \33014 );
and \U$32639 ( \33016 , \33012 , \32815 );
nor \U$32640 ( \33017 , \33015 , \33016 );
xor \U$32641 ( \33018 , \33007 , \33017 );
nand \U$32642 ( \33019 , RIae760a0_34, RIae78b48_125);
xor \U$32643 ( \33020 , \32891 , \32899 );
xor \U$32644 ( \33021 , \33020 , \32908 );
and \U$32645 ( \33022 , \33019 , \33021 );
xor \U$32646 ( \33023 , \32872 , \787 );
xor \U$32647 ( \33024 , \33023 , \32880 );
xor \U$32648 ( \33025 , \32891 , \32899 );
xor \U$32649 ( \33026 , \33025 , \32908 );
and \U$32650 ( \33027 , \33024 , \33026 );
and \U$32651 ( \33028 , \33019 , \33024 );
or \U$32652 ( \33029 , \33022 , \33027 , \33028 );
and \U$32653 ( \33030 , \33018 , \33029 );
and \U$32654 ( \33031 , \33007 , \33017 );
or \U$32655 ( \33032 , \33030 , \33031 );
nor \U$32656 ( \33033 , \32948 , \33032 );
nor \U$32657 ( \33034 , \32945 , \33033 );
nor \U$32658 ( \33035 , \32928 , \33034 );
nor \U$32659 ( \33036 , \32925 , \33035 );
not \U$32660 ( \33037 , \32771 );
not \U$32661 ( \33038 , \32847 );
and \U$32662 ( \33039 , \33037 , \33038 );
and \U$32663 ( \33040 , \32771 , \32847 );
nor \U$32664 ( \33041 , \33039 , \33040 );
or \U$32665 ( \33042 , \33036 , \33041 );
xnor \U$32666 ( \33043 , \33041 , \33036 );
not \U$32667 ( \33044 , \32865 );
not \U$32668 ( \33045 , \33034 );
not \U$32669 ( \33046 , \32924 );
and \U$32670 ( \33047 , \33045 , \33046 );
and \U$32671 ( \33048 , \33034 , \32924 );
nor \U$32672 ( \33049 , \33047 , \33048 );
not \U$32673 ( \33050 , \33049 );
or \U$32674 ( \33051 , \33044 , \33050 );
or \U$32675 ( \33052 , \33049 , \32865 );
nand \U$32676 ( \33053 , \33051 , \33052 );
not \U$32677 ( \33054 , \32930 );
not \U$32678 ( \33055 , \33032 );
not \U$32679 ( \33056 , \32944 );
and \U$32680 ( \33057 , \33055 , \33056 );
and \U$32681 ( \33058 , \33032 , \32944 );
nor \U$32682 ( \33059 , \33057 , \33058 );
not \U$32683 ( \33060 , \33059 );
or \U$32684 ( \33061 , \33054 , \33060 );
or \U$32685 ( \33062 , \33059 , \32930 );
nand \U$32686 ( \33063 , \33061 , \33062 );
not \U$32687 ( \33064 , \33063 );
xor \U$32688 ( \33065 , \32956 , \32964 );
xor \U$32689 ( \33066 , \33065 , \32973 );
and \U$32690 ( \33067 , \33002 , \33066 );
xor \U$32691 ( \33068 , \32983 , \32989 );
xor \U$32692 ( \33069 , \33068 , \32997 );
xor \U$32693 ( \33070 , \32956 , \32964 );
xor \U$32694 ( \33071 , \33070 , \32973 );
and \U$32695 ( \33072 , \33069 , \33071 );
and \U$32696 ( \33073 , \33002 , \33069 );
or \U$32697 ( \33074 , \33067 , \33072 , \33073 );
and \U$32698 ( \33075 , \672 , RIae76be0_58);
and \U$32699 ( \33076 , RIae78ad0_124, \670 );
nor \U$32700 ( \33077 , \33075 , \33076 );
and \U$32701 ( \33078 , \33077 , \588 );
not \U$32702 ( \33079 , \33077 );
and \U$32703 ( \33080 , \33079 , \587 );
nor \U$32704 ( \33081 , \33078 , \33080 );
xor \U$32705 ( \33082 , \33081 , \1012 );
not \U$32706 ( \33083 , \787 );
and \U$32707 ( \33084 , \883 , RIae78d28_129);
and \U$32708 ( \33085 , RIae78e18_131, \881 );
nor \U$32709 ( \33086 , \33084 , \33085 );
not \U$32710 ( \33087 , \33086 );
or \U$32711 ( \33088 , \33083 , \33087 );
or \U$32712 ( \33089 , \33086 , \789 );
nand \U$32713 ( \33090 , \33088 , \33089 );
and \U$32714 ( \33091 , \33082 , \33090 );
and \U$32715 ( \33092 , \33081 , \1012 );
or \U$32716 ( \33093 , \33091 , \33092 );
not \U$32717 ( \33094 , RIae76640_46);
nor \U$32718 ( \33095 , \33094 , \491 );
not \U$32719 ( \33096 , \392 );
and \U$32720 ( \33097 , \384 , RIae76190_36);
and \U$32721 ( \33098 , RIae760a0_34, \382 );
nor \U$32722 ( \33099 , \33097 , \33098 );
not \U$32723 ( \33100 , \33099 );
or \U$32724 ( \33101 , \33096 , \33100 );
or \U$32725 ( \33102 , \33099 , \388 );
nand \U$32726 ( \33103 , \33101 , \33102 );
and \U$32727 ( \33104 , \33095 , \33103 );
xor \U$32728 ( \33105 , \33093 , \33104 );
not \U$32729 ( \33106 , \402 );
and \U$32730 ( \33107 , \436 , RIae76370_40);
and \U$32731 ( \33108 , RIae76280_38, \434 );
nor \U$32732 ( \33109 , \33107 , \33108 );
not \U$32733 ( \33110 , \33109 );
or \U$32734 ( \33111 , \33106 , \33110 );
or \U$32735 ( \33112 , \33109 , \400 );
nand \U$32736 ( \33113 , \33111 , \33112 );
not \U$32737 ( \33114 , \471 );
and \U$32738 ( \33115 , \514 , RIae76af0_56);
and \U$32739 ( \33116 , RIae76a00_54, \512 );
nor \U$32740 ( \33117 , \33115 , \33116 );
not \U$32741 ( \33118 , \33117 );
or \U$32742 ( \33119 , \33114 , \33118 );
or \U$32743 ( \33120 , \33117 , \469 );
nand \U$32744 ( \33121 , \33119 , \33120 );
xor \U$32745 ( \33122 , \33113 , \33121 );
and \U$32746 ( \33123 , \558 , RIae76820_50);
and \U$32747 ( \33124 , RIae76910_52, \556 );
nor \U$32748 ( \33125 , \33123 , \33124 );
and \U$32749 ( \33126 , \33125 , \504 );
not \U$32750 ( \33127 , \33125 );
and \U$32751 ( \33128 , \33127 , \562 );
nor \U$32752 ( \33129 , \33126 , \33128 );
and \U$32753 ( \33130 , \33122 , \33129 );
and \U$32754 ( \33131 , \33113 , \33121 );
or \U$32755 ( \33132 , \33130 , \33131 );
and \U$32756 ( \33133 , \33105 , \33132 );
and \U$32757 ( \33134 , \33093 , \33104 );
or \U$32758 ( \33135 , \33133 , \33134 );
and \U$32759 ( \33136 , \33074 , \33135 );
not \U$32760 ( \33137 , \33074 );
not \U$32761 ( \33138 , \33135 );
and \U$32762 ( \33139 , \33137 , \33138 );
xor \U$32763 ( \33140 , \32891 , \32899 );
xor \U$32764 ( \33141 , \33140 , \32908 );
xor \U$32765 ( \33142 , \33019 , \33024 );
xor \U$32766 ( \33143 , \33141 , \33142 );
nor \U$32767 ( \33144 , \33139 , \33143 );
nor \U$32768 ( \33145 , \33136 , \33144 );
not \U$32769 ( \33146 , \32932 );
not \U$32770 ( \33147 , \32943 );
and \U$32771 ( \33148 , \33146 , \33147 );
and \U$32772 ( \33149 , \32932 , \32943 );
nor \U$32773 ( \33150 , \33148 , \33149 );
xor \U$32774 ( \33151 , \33145 , \33150 );
xor \U$32775 ( \33152 , \33007 , \33017 );
xor \U$32776 ( \33153 , \33152 , \33029 );
and \U$32777 ( \33154 , \33151 , \33153 );
and \U$32778 ( \33155 , \33145 , \33150 );
or \U$32779 ( \33156 , \33154 , \33155 );
nor \U$32780 ( \33157 , \33064 , \33156 );
and \U$32781 ( \33158 , \33053 , \33157 );
xor \U$32782 ( \33159 , \33157 , \33053 );
and \U$32783 ( \33160 , \558 , RIae76370_40);
and \U$32784 ( \33161 , RIae76280_38, \556 );
nor \U$32785 ( \33162 , \33160 , \33161 );
and \U$32786 ( \33163 , \33162 , \562 );
not \U$32787 ( \33164 , \33162 );
and \U$32788 ( \33165 , \33164 , \504 );
nor \U$32789 ( \33166 , \33163 , \33165 );
and \U$32790 ( \33167 , \672 , RIae76af0_56);
and \U$32791 ( \33168 , RIae76a00_54, \670 );
nor \U$32792 ( \33169 , \33167 , \33168 );
and \U$32793 ( \33170 , \33169 , \587 );
not \U$32794 ( \33171 , \33169 );
and \U$32795 ( \33172 , \33171 , \588 );
nor \U$32796 ( \33173 , \33170 , \33172 );
xor \U$32797 ( \33174 , \33166 , \33173 );
and \U$32798 ( \33175 , \883 , RIae76820_50);
and \U$32799 ( \33176 , RIae76910_52, \881 );
nor \U$32800 ( \33177 , \33175 , \33176 );
not \U$32801 ( \33178 , \33177 );
not \U$32802 ( \33179 , \787 );
and \U$32803 ( \33180 , \33178 , \33179 );
and \U$32804 ( \33181 , \33177 , \787 );
nor \U$32805 ( \33182 , \33180 , \33181 );
and \U$32806 ( \33183 , \33174 , \33182 );
and \U$32807 ( \33184 , \33166 , \33173 );
or \U$32808 ( \33185 , \33183 , \33184 );
and \U$32809 ( \33186 , \1138 , RIae76be0_58);
and \U$32810 ( \33187 , RIae78ad0_124, \1136 );
nor \U$32811 ( \33188 , \33186 , \33187 );
and \U$32812 ( \33189 , \33188 , \1142 );
not \U$32813 ( \33190 , \33188 );
and \U$32814 ( \33191 , \33190 , \1012 );
nor \U$32815 ( \33192 , \33189 , \33191 );
not \U$32816 ( \33193 , \33192 );
not \U$32817 ( \33194 , \1488 );
and \U$32818 ( \33195 , \33193 , \33194 );
and \U$32819 ( \33196 , \33192 , \1488 );
and \U$32820 ( \33197 , \1376 , RIae78d28_129);
and \U$32821 ( \33198 , RIae78e18_131, \1374 );
nor \U$32822 ( \33199 , \33197 , \33198 );
and \U$32823 ( \33200 , \33199 , \1261 );
not \U$32824 ( \33201 , \33199 );
and \U$32825 ( \33202 , \33201 , \1380 );
nor \U$32826 ( \33203 , \33200 , \33202 );
nor \U$32827 ( \33204 , \33196 , \33203 );
nor \U$32828 ( \33205 , \33195 , \33204 );
xor \U$32829 ( \33206 , \33185 , \33205 );
and \U$32830 ( \33207 , \514 , RIae76190_36);
and \U$32831 ( \33208 , RIae760a0_34, \512 );
nor \U$32832 ( \33209 , \33207 , \33208 );
not \U$32833 ( \33210 , \33209 );
not \U$32834 ( \33211 , \471 );
and \U$32835 ( \33212 , \33210 , \33211 );
and \U$32836 ( \33213 , \33209 , \469 );
nor \U$32837 ( \33214 , \33212 , \33213 );
and \U$32838 ( \33215 , \384 , RIae76460_42);
and \U$32839 ( \33216 , RIae76550_44, \382 );
nor \U$32840 ( \33217 , \33215 , \33216 );
not \U$32841 ( \33218 , \33217 );
not \U$32842 ( \33219 , \392 );
and \U$32843 ( \33220 , \33218 , \33219 );
and \U$32844 ( \33221 , \33217 , \388 );
nor \U$32845 ( \33222 , \33220 , \33221 );
xor \U$32846 ( \33223 , \33214 , \33222 );
and \U$32847 ( \33224 , \436 , RIae76730_48);
and \U$32848 ( \33225 , RIae76640_46, \434 );
nor \U$32849 ( \33226 , \33224 , \33225 );
not \U$32850 ( \33227 , \33226 );
not \U$32851 ( \33228 , \402 );
and \U$32852 ( \33229 , \33227 , \33228 );
and \U$32853 ( \33230 , \33226 , \402 );
nor \U$32854 ( \33231 , \33229 , \33230 );
and \U$32855 ( \33232 , \33223 , \33231 );
and \U$32856 ( \33233 , \33214 , \33222 );
or \U$32857 ( \33234 , \33232 , \33233 );
and \U$32858 ( \33235 , \33206 , \33234 );
and \U$32859 ( \33236 , \33185 , \33205 );
or \U$32860 ( \33237 , \33235 , \33236 );
and \U$32861 ( \33238 , \384 , RIae76550_44);
and \U$32862 ( \33239 , RIae76730_48, \382 );
nor \U$32863 ( \33240 , \33238 , \33239 );
not \U$32864 ( \33241 , \33240 );
not \U$32865 ( \33242 , \388 );
and \U$32866 ( \33243 , \33241 , \33242 );
and \U$32867 ( \33244 , \33240 , \388 );
nor \U$32868 ( \33245 , \33243 , \33244 );
nand \U$32869 ( \33246 , RIae76460_42, RIae78b48_125);
xor \U$32870 ( \33247 , \33245 , \33246 );
and \U$32871 ( \33248 , \436 , RIae76640_46);
and \U$32872 ( \33249 , RIae76190_36, \434 );
nor \U$32873 ( \33250 , \33248 , \33249 );
not \U$32874 ( \33251 , \33250 );
not \U$32875 ( \33252 , \402 );
and \U$32876 ( \33253 , \33251 , \33252 );
and \U$32877 ( \33254 , \33250 , \400 );
nor \U$32878 ( \33255 , \33253 , \33254 );
xor \U$32879 ( \33256 , \33247 , \33255 );
and \U$32880 ( \33257 , \672 , RIae76a00_54);
and \U$32881 ( \33258 , RIae76820_50, \670 );
nor \U$32882 ( \33259 , \33257 , \33258 );
and \U$32883 ( \33260 , \33259 , \587 );
not \U$32884 ( \33261 , \33259 );
and \U$32885 ( \33262 , \33261 , \588 );
nor \U$32886 ( \33263 , \33260 , \33262 );
and \U$32887 ( \33264 , \514 , RIae760a0_34);
and \U$32888 ( \33265 , RIae76370_40, \512 );
nor \U$32889 ( \33266 , \33264 , \33265 );
not \U$32890 ( \33267 , \33266 );
not \U$32891 ( \33268 , \471 );
and \U$32892 ( \33269 , \33267 , \33268 );
and \U$32893 ( \33270 , \33266 , \471 );
nor \U$32894 ( \33271 , \33269 , \33270 );
xor \U$32895 ( \33272 , \33263 , \33271 );
and \U$32896 ( \33273 , \558 , RIae76280_38);
and \U$32897 ( \33274 , RIae76af0_56, \556 );
nor \U$32898 ( \33275 , \33273 , \33274 );
and \U$32899 ( \33276 , \33275 , \562 );
not \U$32900 ( \33277 , \33275 );
and \U$32901 ( \33278 , \33277 , \504 );
nor \U$32902 ( \33279 , \33276 , \33278 );
xor \U$32903 ( \33280 , \33272 , \33279 );
nand \U$32904 ( \33281 , \33256 , \33280 );
not \U$32905 ( \33282 , \33281 );
xor \U$32906 ( \33283 , \33237 , \33282 );
and \U$32907 ( \33284 , \384 , RIae76730_48);
and \U$32908 ( \33285 , RIae76640_46, \382 );
nor \U$32909 ( \33286 , \33284 , \33285 );
not \U$32910 ( \33287 , \33286 );
not \U$32911 ( \33288 , \392 );
and \U$32912 ( \33289 , \33287 , \33288 );
and \U$32913 ( \33290 , \33286 , \388 );
nor \U$32914 ( \33291 , \33289 , \33290 );
nand \U$32915 ( \33292 , RIae76550_44, RIae78b48_125);
xor \U$32916 ( \33293 , \33291 , \33292 );
and \U$32917 ( \33294 , \436 , RIae76190_36);
and \U$32918 ( \33295 , RIae760a0_34, \434 );
nor \U$32919 ( \33296 , \33294 , \33295 );
not \U$32920 ( \33297 , \33296 );
not \U$32921 ( \33298 , \402 );
and \U$32922 ( \33299 , \33297 , \33298 );
and \U$32923 ( \33300 , \33296 , \402 );
nor \U$32924 ( \33301 , \33299 , \33300 );
xor \U$32925 ( \33302 , \33293 , \33301 );
and \U$32926 ( \33303 , \1138 , RIae78d28_129);
and \U$32927 ( \33304 , RIae78e18_131, \1136 );
nor \U$32928 ( \33305 , \33303 , \33304 );
and \U$32929 ( \33306 , \33305 , \1142 );
not \U$32930 ( \33307 , \33305 );
and \U$32931 ( \33308 , \33307 , \1012 );
nor \U$32932 ( \33309 , \33306 , \33308 );
and \U$32933 ( \33310 , \33309 , \1261 );
not \U$32934 ( \33311 , \33309 );
and \U$32935 ( \33312 , \33311 , \1380 );
nor \U$32936 ( \33313 , \33310 , \33312 );
not \U$32937 ( \33314 , \33313 );
and \U$32938 ( \33315 , \883 , RIae76be0_58);
and \U$32939 ( \33316 , RIae78ad0_124, \881 );
nor \U$32940 ( \33317 , \33315 , \33316 );
not \U$32941 ( \33318 , \33317 );
not \U$32942 ( \33319 , \787 );
and \U$32943 ( \33320 , \33318 , \33319 );
and \U$32944 ( \33321 , \33317 , \789 );
nor \U$32945 ( \33322 , \33320 , \33321 );
not \U$32946 ( \33323 , \33322 );
and \U$32947 ( \33324 , \33314 , \33323 );
and \U$32948 ( \33325 , \33313 , \33322 );
nor \U$32949 ( \33326 , \33324 , \33325 );
and \U$32950 ( \33327 , \672 , RIae76820_50);
and \U$32951 ( \33328 , RIae76910_52, \670 );
nor \U$32952 ( \33329 , \33327 , \33328 );
and \U$32953 ( \33330 , \33329 , \587 );
not \U$32954 ( \33331 , \33329 );
and \U$32955 ( \33332 , \33331 , \588 );
nor \U$32956 ( \33333 , \33330 , \33332 );
and \U$32957 ( \33334 , \514 , RIae76370_40);
and \U$32958 ( \33335 , RIae76280_38, \512 );
nor \U$32959 ( \33336 , \33334 , \33335 );
not \U$32960 ( \33337 , \33336 );
not \U$32961 ( \33338 , \471 );
and \U$32962 ( \33339 , \33337 , \33338 );
and \U$32963 ( \33340 , \33336 , \471 );
nor \U$32964 ( \33341 , \33339 , \33340 );
xor \U$32965 ( \33342 , \33333 , \33341 );
and \U$32966 ( \33343 , \558 , RIae76af0_56);
and \U$32967 ( \33344 , RIae76a00_54, \556 );
nor \U$32968 ( \33345 , \33343 , \33344 );
and \U$32969 ( \33346 , \33345 , \562 );
not \U$32970 ( \33347 , \33345 );
and \U$32971 ( \33348 , \33347 , \504 );
nor \U$32972 ( \33349 , \33346 , \33348 );
xor \U$32973 ( \33350 , \33342 , \33349 );
xor \U$32974 ( \33351 , \33326 , \33350 );
xor \U$32975 ( \33352 , \33302 , \33351 );
and \U$32976 ( \33353 , \33283 , \33352 );
and \U$32977 ( \33354 , \33237 , \33282 );
or \U$32978 ( \33355 , \33353 , \33354 );
or \U$32979 ( \33356 , \33309 , \1261 );
and \U$32980 ( \33357 , \33309 , \1261 );
nor \U$32981 ( \33358 , \33357 , \33322 );
not \U$32982 ( \33359 , \33358 );
nand \U$32983 ( \33360 , \33356 , \33359 );
not \U$32984 ( \33361 , \33360 );
xor \U$32985 ( \33362 , \33291 , \33292 );
and \U$32986 ( \33363 , \33362 , \33301 );
and \U$32987 ( \33364 , \33291 , \33292 );
or \U$32988 ( \33365 , \33363 , \33364 );
not \U$32989 ( \33366 , \33365 );
or \U$32990 ( \33367 , \33361 , \33366 );
or \U$32991 ( \33368 , \33365 , \33360 );
nand \U$32992 ( \33369 , \33367 , \33368 );
not \U$32993 ( \33370 , \33369 );
xor \U$32994 ( \33371 , \33333 , \33341 );
and \U$32995 ( \33372 , \33371 , \33349 );
and \U$32996 ( \33373 , \33333 , \33341 );
or \U$32997 ( \33374 , \33372 , \33373 );
not \U$32998 ( \33375 , \33374 );
and \U$32999 ( \33376 , \33370 , \33375 );
and \U$33000 ( \33377 , \33369 , \33374 );
nor \U$33001 ( \33378 , \33376 , \33377 );
xor \U$33002 ( \33379 , \33355 , \33378 );
xor \U$33003 ( \33380 , \33291 , \33292 );
xor \U$33004 ( \33381 , \33380 , \33301 );
and \U$33005 ( \33382 , \33326 , \33381 );
xor \U$33006 ( \33383 , \33291 , \33292 );
xor \U$33007 ( \33384 , \33383 , \33301 );
and \U$33008 ( \33385 , \33350 , \33384 );
and \U$33009 ( \33386 , \33326 , \33350 );
or \U$33010 ( \33387 , \33382 , \33385 , \33386 );
and \U$33011 ( \33388 , \883 , RIae76910_52);
and \U$33012 ( \33389 , RIae76be0_58, \881 );
nor \U$33013 ( \33390 , \33388 , \33389 );
not \U$33014 ( \33391 , \33390 );
not \U$33015 ( \33392 , \787 );
and \U$33016 ( \33393 , \33391 , \33392 );
and \U$33017 ( \33394 , \33390 , \787 );
nor \U$33018 ( \33395 , \33393 , \33394 );
nand \U$33019 ( \33396 , RIae78e18_131, \1376 );
and \U$33020 ( \33397 , \33396 , \1261 );
not \U$33021 ( \33398 , \33396 );
and \U$33022 ( \33399 , \33398 , \1380 );
nor \U$33023 ( \33400 , \33397 , \33399 );
xor \U$33024 ( \33401 , \33395 , \33400 );
and \U$33025 ( \33402 , \1138 , RIae78ad0_124);
and \U$33026 ( \33403 , RIae78d28_129, \1136 );
nor \U$33027 ( \33404 , \33402 , \33403 );
and \U$33028 ( \33405 , \33404 , \1142 );
not \U$33029 ( \33406 , \33404 );
and \U$33030 ( \33407 , \33406 , \1012 );
nor \U$33031 ( \33408 , \33405 , \33407 );
and \U$33032 ( \33409 , \33401 , \33408 );
and \U$33033 ( \33410 , \33395 , \33400 );
or \U$33034 ( \33411 , \33409 , \33410 );
xor \U$33035 ( \33412 , \33245 , \33246 );
and \U$33036 ( \33413 , \33412 , \33255 );
and \U$33037 ( \33414 , \33245 , \33246 );
or \U$33038 ( \33415 , \33413 , \33414 );
xor \U$33039 ( \33416 , \33411 , \33415 );
xor \U$33040 ( \33417 , \33263 , \33271 );
and \U$33041 ( \33418 , \33417 , \33279 );
and \U$33042 ( \33419 , \33263 , \33271 );
or \U$33043 ( \33420 , \33418 , \33419 );
and \U$33044 ( \33421 , \33416 , \33420 );
and \U$33045 ( \33422 , \33411 , \33415 );
or \U$33046 ( \33423 , \33421 , \33422 );
xor \U$33047 ( \33424 , \33387 , \33423 );
nand \U$33048 ( \33425 , RIae78e18_131, \1138 );
and \U$33049 ( \33426 , \33425 , \1012 );
not \U$33050 ( \33427 , \33425 );
and \U$33051 ( \33428 , \33427 , \1142 );
nor \U$33052 ( \33429 , \33426 , \33428 );
not \U$33053 ( \33430 , \33429 );
and \U$33054 ( \33431 , \883 , RIae78ad0_124);
and \U$33055 ( \33432 , RIae78d28_129, \881 );
nor \U$33056 ( \33433 , \33431 , \33432 );
not \U$33057 ( \33434 , \33433 );
not \U$33058 ( \33435 , \789 );
and \U$33059 ( \33436 , \33434 , \33435 );
and \U$33060 ( \33437 , \33433 , \789 );
nor \U$33061 ( \33438 , \33436 , \33437 );
not \U$33062 ( \33439 , \33438 );
or \U$33063 ( \33440 , \33430 , \33439 );
or \U$33064 ( \33441 , \33438 , \33429 );
nand \U$33065 ( \33442 , \33440 , \33441 );
not \U$33066 ( \33443 , \33442 );
and \U$33067 ( \33444 , \672 , RIae76910_52);
and \U$33068 ( \33445 , RIae76be0_58, \670 );
nor \U$33069 ( \33446 , \33444 , \33445 );
and \U$33070 ( \33447 , \33446 , \587 );
not \U$33071 ( \33448 , \33446 );
and \U$33072 ( \33449 , \33448 , \588 );
nor \U$33073 ( \33450 , \33447 , \33449 );
not \U$33074 ( \33451 , \33450 );
and \U$33075 ( \33452 , \33443 , \33451 );
and \U$33076 ( \33453 , \33442 , \33450 );
nor \U$33077 ( \33454 , \33452 , \33453 );
and \U$33078 ( \33455 , \514 , RIae76280_38);
and \U$33079 ( \33456 , RIae76af0_56, \512 );
nor \U$33080 ( \33457 , \33455 , \33456 );
not \U$33081 ( \33458 , \33457 );
not \U$33082 ( \33459 , \469 );
and \U$33083 ( \33460 , \33458 , \33459 );
and \U$33084 ( \33461 , \33457 , \471 );
nor \U$33085 ( \33462 , \33460 , \33461 );
and \U$33086 ( \33463 , \558 , RIae76a00_54);
and \U$33087 ( \33464 , RIae76820_50, \556 );
nor \U$33088 ( \33465 , \33463 , \33464 );
and \U$33089 ( \33466 , \33465 , \562 );
not \U$33090 ( \33467 , \33465 );
and \U$33091 ( \33468 , \33467 , \504 );
nor \U$33092 ( \33469 , \33466 , \33468 );
xor \U$33093 ( \33470 , \33462 , \33469 );
and \U$33094 ( \33471 , \436 , RIae760a0_34);
and \U$33095 ( \33472 , RIae76370_40, \434 );
nor \U$33096 ( \33473 , \33471 , \33472 );
not \U$33097 ( \33474 , \33473 );
not \U$33098 ( \33475 , \402 );
and \U$33099 ( \33476 , \33474 , \33475 );
and \U$33100 ( \33477 , \33473 , \400 );
nor \U$33101 ( \33478 , \33476 , \33477 );
xor \U$33102 ( \33479 , \33470 , \33478 );
xnor \U$33103 ( \33480 , \33454 , \33479 );
not \U$33104 ( \33481 , \33480 );
and \U$33105 ( \33482 , \384 , RIae76640_46);
and \U$33106 ( \33483 , RIae76190_36, \382 );
nor \U$33107 ( \33484 , \33482 , \33483 );
not \U$33108 ( \33485 , \33484 );
not \U$33109 ( \33486 , \388 );
and \U$33110 ( \33487 , \33485 , \33486 );
and \U$33111 ( \33488 , \33484 , \388 );
nor \U$33112 ( \33489 , \33487 , \33488 );
nand \U$33113 ( \33490 , RIae76730_48, RIae78b48_125);
or \U$33114 ( \33491 , \33489 , \33490 );
nand \U$33115 ( \33492 , \33490 , \33489 );
nand \U$33116 ( \33493 , \33491 , \33492 );
not \U$33117 ( \33494 , \33493 );
and \U$33118 ( \33495 , \33481 , \33494 );
and \U$33119 ( \33496 , \33480 , \33493 );
nor \U$33120 ( \33497 , \33495 , \33496 );
xor \U$33121 ( \33498 , \33424 , \33497 );
xor \U$33122 ( \33499 , \33379 , \33498 );
not \U$33123 ( \33500 , \33499 );
and \U$33124 ( \33501 , \1138 , RIae76910_52);
and \U$33125 ( \33502 , RIae76be0_58, \1136 );
nor \U$33126 ( \33503 , \33501 , \33502 );
and \U$33127 ( \33504 , \33503 , \1142 );
not \U$33128 ( \33505 , \33503 );
and \U$33129 ( \33506 , \33505 , \1012 );
nor \U$33130 ( \33507 , \33504 , \33506 );
not \U$33131 ( \33508 , \33507 );
and \U$33132 ( \33509 , \1376 , RIae78ad0_124);
and \U$33133 ( \33510 , RIae78d28_129, \1374 );
nor \U$33134 ( \33511 , \33509 , \33510 );
and \U$33135 ( \33512 , \33511 , \1261 );
not \U$33136 ( \33513 , \33511 );
and \U$33137 ( \33514 , \33513 , \1380 );
nor \U$33138 ( \33515 , \33512 , \33514 );
not \U$33139 ( \33516 , \33515 );
and \U$33140 ( \33517 , \33508 , \33516 );
and \U$33141 ( \33518 , \33515 , \33507 );
nand \U$33142 ( \33519 , RIae78e18_131, \1593 );
and \U$33143 ( \33520 , \33519 , \1488 );
not \U$33144 ( \33521 , \33519 );
and \U$33145 ( \33522 , \33521 , \1498 );
nor \U$33146 ( \33523 , \33520 , \33522 );
nor \U$33147 ( \33524 , \33518 , \33523 );
nor \U$33148 ( \33525 , \33517 , \33524 );
not \U$33149 ( \33526 , \33525 );
and \U$33150 ( \33527 , \384 , RIae75470_8);
and \U$33151 ( \33528 , RIae76460_42, \382 );
nor \U$33152 ( \33529 , \33527 , \33528 );
not \U$33153 ( \33530 , \33529 );
not \U$33154 ( \33531 , \388 );
and \U$33155 ( \33532 , \33530 , \33531 );
and \U$33156 ( \33533 , \33529 , \388 );
nor \U$33157 ( \33534 , \33532 , \33533 );
and \U$33158 ( \33535 , \436 , RIae76550_44);
and \U$33159 ( \33536 , RIae76730_48, \434 );
nor \U$33160 ( \33537 , \33535 , \33536 );
not \U$33161 ( \33538 , \33537 );
not \U$33162 ( \33539 , \402 );
and \U$33163 ( \33540 , \33538 , \33539 );
and \U$33164 ( \33541 , \33537 , \402 );
nor \U$33165 ( \33542 , \33540 , \33541 );
xor \U$33166 ( \33543 , \33534 , \33542 );
and \U$33167 ( \33544 , \514 , RIae76640_46);
and \U$33168 ( \33545 , RIae76190_36, \512 );
nor \U$33169 ( \33546 , \33544 , \33545 );
not \U$33170 ( \33547 , \33546 );
not \U$33171 ( \33548 , \469 );
and \U$33172 ( \33549 , \33547 , \33548 );
and \U$33173 ( \33550 , \33546 , \471 );
nor \U$33174 ( \33551 , \33549 , \33550 );
and \U$33175 ( \33552 , \33543 , \33551 );
and \U$33176 ( \33553 , \33534 , \33542 );
or \U$33177 ( \33554 , \33552 , \33553 );
not \U$33178 ( \33555 , \33554 );
and \U$33179 ( \33556 , \33526 , \33555 );
and \U$33180 ( \33557 , \33525 , \33554 );
and \U$33181 ( \33558 , \672 , RIae76280_38);
and \U$33182 ( \33559 , RIae76af0_56, \670 );
nor \U$33183 ( \33560 , \33558 , \33559 );
and \U$33184 ( \33561 , \33560 , \588 );
not \U$33185 ( \33562 , \33560 );
and \U$33186 ( \33563 , \33562 , \587 );
nor \U$33187 ( \33564 , \33561 , \33563 );
not \U$33188 ( \33565 , \789 );
and \U$33189 ( \33566 , \883 , RIae76a00_54);
and \U$33190 ( \33567 , RIae76820_50, \881 );
nor \U$33191 ( \33568 , \33566 , \33567 );
not \U$33192 ( \33569 , \33568 );
or \U$33193 ( \33570 , \33565 , \33569 );
or \U$33194 ( \33571 , \33568 , \787 );
nand \U$33195 ( \33572 , \33570 , \33571 );
xor \U$33196 ( \33573 , \33564 , \33572 );
and \U$33197 ( \33574 , \558 , RIae760a0_34);
and \U$33198 ( \33575 , RIae76370_40, \556 );
nor \U$33199 ( \33576 , \33574 , \33575 );
and \U$33200 ( \33577 , \33576 , \504 );
not \U$33201 ( \33578 , \33576 );
and \U$33202 ( \33579 , \33578 , \562 );
nor \U$33203 ( \33580 , \33577 , \33579 );
and \U$33204 ( \33581 , \33573 , \33580 );
and \U$33205 ( \33582 , \33564 , \33572 );
nor \U$33206 ( \33583 , \33581 , \33582 );
nor \U$33207 ( \33584 , \33557 , \33583 );
nor \U$33208 ( \33585 , \33556 , \33584 );
not \U$33209 ( \33586 , \33585 );
xor \U$33210 ( \33587 , \33395 , \33400 );
xor \U$33211 ( \33588 , \33587 , \33408 );
not \U$33212 ( \33589 , \33588 );
and \U$33213 ( \33590 , \33586 , \33589 );
and \U$33214 ( \33591 , \33585 , \33588 );
xor \U$33215 ( \33592 , \33214 , \33222 );
xor \U$33216 ( \33593 , \33592 , \33231 );
not \U$33217 ( \33594 , \33593 );
nand \U$33218 ( \33595 , RIae75470_8, RIae78b48_125);
not \U$33219 ( \33596 , \33595 );
and \U$33220 ( \33597 , \33594 , \33596 );
and \U$33221 ( \33598 , \33593 , \33595 );
xor \U$33222 ( \33599 , \33166 , \33173 );
xor \U$33223 ( \33600 , \33599 , \33182 );
nor \U$33224 ( \33601 , \33598 , \33600 );
nor \U$33225 ( \33602 , \33597 , \33601 );
nor \U$33226 ( \33603 , \33591 , \33602 );
nor \U$33227 ( \33604 , \33590 , \33603 );
xor \U$33228 ( \33605 , \33411 , \33415 );
xor \U$33229 ( \33606 , \33605 , \33420 );
xor \U$33230 ( \33607 , \33604 , \33606 );
xor \U$33231 ( \33608 , \33237 , \33282 );
xor \U$33232 ( \33609 , \33608 , \33352 );
and \U$33233 ( \33610 , \33607 , \33609 );
and \U$33234 ( \33611 , \33604 , \33606 );
or \U$33235 ( \33612 , \33610 , \33611 );
not \U$33236 ( \33613 , \33612 );
xor \U$33237 ( \33614 , \33604 , \33606 );
xor \U$33238 ( \33615 , \33614 , \33609 );
xor \U$33239 ( \33616 , \33185 , \33205 );
xor \U$33240 ( \33617 , \33616 , \33234 );
not \U$33241 ( \33618 , \33617 );
not \U$33242 ( \33619 , \33588 );
xor \U$33243 ( \33620 , \33585 , \33602 );
not \U$33244 ( \33621 , \33620 );
or \U$33245 ( \33622 , \33619 , \33621 );
or \U$33246 ( \33623 , \33620 , \33588 );
nand \U$33247 ( \33624 , \33622 , \33623 );
nand \U$33248 ( \33625 , \33618 , \33624 );
or \U$33249 ( \33626 , \33615 , \33625 );
not \U$33250 ( \33627 , \33625 );
not \U$33251 ( \33628 , \33615 );
or \U$33252 ( \33629 , \33627 , \33628 );
xor \U$33253 ( \33630 , \33564 , \33572 );
xor \U$33254 ( \33631 , \33630 , \33580 );
not \U$33255 ( \33632 , \33507 );
xor \U$33256 ( \33633 , \33523 , \33515 );
not \U$33257 ( \33634 , \33633 );
or \U$33258 ( \33635 , \33632 , \33634 );
or \U$33259 ( \33636 , \33633 , \33507 );
nand \U$33260 ( \33637 , \33635 , \33636 );
and \U$33261 ( \33638 , \33631 , \33637 );
nand \U$33262 ( \33639 , RIae75380_6, RIae78b48_125);
xor \U$33263 ( \33640 , \33534 , \33542 );
xor \U$33264 ( \33641 , \33640 , \33551 );
nand \U$33265 ( \33642 , \33639 , \33641 );
xor \U$33266 ( \33643 , \33638 , \33642 );
and \U$33267 ( \33644 , \514 , RIae76730_48);
and \U$33268 ( \33645 , RIae76640_46, \512 );
nor \U$33269 ( \33646 , \33644 , \33645 );
not \U$33270 ( \33647 , \33646 );
not \U$33271 ( \33648 , \469 );
and \U$33272 ( \33649 , \33647 , \33648 );
and \U$33273 ( \33650 , \33646 , \469 );
nor \U$33274 ( \33651 , \33649 , \33650 );
and \U$33275 ( \33652 , \558 , RIae76190_36);
and \U$33276 ( \33653 , RIae760a0_34, \556 );
nor \U$33277 ( \33654 , \33652 , \33653 );
and \U$33278 ( \33655 , \33654 , \562 );
not \U$33279 ( \33656 , \33654 );
and \U$33280 ( \33657 , \33656 , \504 );
nor \U$33281 ( \33658 , \33655 , \33657 );
xor \U$33282 ( \33659 , \33651 , \33658 );
and \U$33283 ( \33660 , \436 , RIae76460_42);
and \U$33284 ( \33661 , RIae76550_44, \434 );
nor \U$33285 ( \33662 , \33660 , \33661 );
not \U$33286 ( \33663 , \33662 );
not \U$33287 ( \33664 , \400 );
and \U$33288 ( \33665 , \33663 , \33664 );
and \U$33289 ( \33666 , \33662 , \400 );
nor \U$33290 ( \33667 , \33665 , \33666 );
and \U$33291 ( \33668 , \33659 , \33667 );
and \U$33292 ( \33669 , \33651 , \33658 );
nor \U$33293 ( \33670 , \33668 , \33669 );
and \U$33294 ( \33671 , \1376 , RIae76be0_58);
and \U$33295 ( \33672 , RIae78ad0_124, \1374 );
nor \U$33296 ( \33673 , \33671 , \33672 );
and \U$33297 ( \33674 , \33673 , \1380 );
not \U$33298 ( \33675 , \33673 );
and \U$33299 ( \33676 , \33675 , \1261 );
nor \U$33300 ( \33677 , \33674 , \33676 );
xor \U$33301 ( \33678 , \33677 , \1735 );
and \U$33302 ( \33679 , \1593 , RIae78d28_129);
and \U$33303 ( \33680 , RIae78e18_131, \1591 );
nor \U$33304 ( \33681 , \33679 , \33680 );
and \U$33305 ( \33682 , \33681 , \1498 );
not \U$33306 ( \33683 , \33681 );
and \U$33307 ( \33684 , \33683 , \1488 );
nor \U$33308 ( \33685 , \33682 , \33684 );
and \U$33309 ( \33686 , \33678 , \33685 );
and \U$33310 ( \33687 , \33677 , \1735 );
or \U$33311 ( \33688 , \33686 , \33687 );
xor \U$33312 ( \33689 , \33670 , \33688 );
and \U$33313 ( \33690 , \672 , RIae76370_40);
and \U$33314 ( \33691 , RIae76280_38, \670 );
nor \U$33315 ( \33692 , \33690 , \33691 );
and \U$33316 ( \33693 , \33692 , \587 );
not \U$33317 ( \33694 , \33692 );
and \U$33318 ( \33695 , \33694 , \588 );
nor \U$33319 ( \33696 , \33693 , \33695 );
and \U$33320 ( \33697 , \883 , RIae76af0_56);
and \U$33321 ( \33698 , RIae76a00_54, \881 );
nor \U$33322 ( \33699 , \33697 , \33698 );
not \U$33323 ( \33700 , \33699 );
not \U$33324 ( \33701 , \787 );
and \U$33325 ( \33702 , \33700 , \33701 );
and \U$33326 ( \33703 , \33699 , \789 );
nor \U$33327 ( \33704 , \33702 , \33703 );
or \U$33328 ( \33705 , \33696 , \33704 );
not \U$33329 ( \33706 , \33704 );
not \U$33330 ( \33707 , \33696 );
or \U$33331 ( \33708 , \33706 , \33707 );
and \U$33332 ( \33709 , \1138 , RIae76820_50);
and \U$33333 ( \33710 , RIae76910_52, \1136 );
nor \U$33334 ( \33711 , \33709 , \33710 );
and \U$33335 ( \33712 , \33711 , \1012 );
not \U$33336 ( \33713 , \33711 );
and \U$33337 ( \33714 , \33713 , \1142 );
nor \U$33338 ( \33715 , \33712 , \33714 );
nand \U$33339 ( \33716 , \33708 , \33715 );
nand \U$33340 ( \33717 , \33705 , \33716 );
and \U$33341 ( \33718 , \33689 , \33717 );
and \U$33342 ( \33719 , \33670 , \33688 );
or \U$33343 ( \33720 , \33718 , \33719 );
and \U$33344 ( \33721 , \33643 , \33720 );
and \U$33345 ( \33722 , \33638 , \33642 );
or \U$33346 ( \33723 , \33721 , \33722 );
or \U$33347 ( \33724 , \33256 , \33280 );
nand \U$33348 ( \33725 , \33724 , \33281 );
xor \U$33349 ( \33726 , \33723 , \33725 );
not \U$33350 ( \33727 , \33554 );
xor \U$33351 ( \33728 , \33525 , \33583 );
not \U$33352 ( \33729 , \33728 );
or \U$33353 ( \33730 , \33727 , \33729 );
or \U$33354 ( \33731 , \33728 , \33554 );
nand \U$33355 ( \33732 , \33730 , \33731 );
not \U$33356 ( \33733 , \33192 );
and \U$33357 ( \33734 , \33203 , \1488 );
not \U$33358 ( \33735 , \33203 );
and \U$33359 ( \33736 , \33735 , \1498 );
nor \U$33360 ( \33737 , \33734 , \33736 );
not \U$33361 ( \33738 , \33737 );
or \U$33362 ( \33739 , \33733 , \33738 );
or \U$33363 ( \33740 , \33737 , \33192 );
nand \U$33364 ( \33741 , \33739 , \33740 );
xor \U$33365 ( \33742 , \33732 , \33741 );
not \U$33366 ( \33743 , \33593 );
xor \U$33367 ( \33744 , \33595 , \33600 );
not \U$33368 ( \33745 , \33744 );
or \U$33369 ( \33746 , \33743 , \33745 );
or \U$33370 ( \33747 , \33744 , \33593 );
nand \U$33371 ( \33748 , \33746 , \33747 );
and \U$33372 ( \33749 , \33742 , \33748 );
and \U$33373 ( \33750 , \33732 , \33741 );
or \U$33374 ( \33751 , \33749 , \33750 );
and \U$33375 ( \33752 , \33726 , \33751 );
and \U$33376 ( \33753 , \33723 , \33725 );
or \U$33377 ( \33754 , \33752 , \33753 );
nand \U$33378 ( \33755 , \33629 , \33754 );
nand \U$33379 ( \33756 , \33626 , \33755 );
not \U$33380 ( \33757 , \33756 );
or \U$33381 ( \33758 , \33613 , \33757 );
or \U$33382 ( \33759 , \33756 , \33612 );
nand \U$33383 ( \33760 , \33758 , \33759 );
not \U$33384 ( \33761 , \33760 );
or \U$33385 ( \33762 , \33500 , \33761 );
or \U$33386 ( \33763 , \33760 , \33499 );
nand \U$33387 ( \33764 , \33762 , \33763 );
not \U$33388 ( \33765 , \33617 );
not \U$33389 ( \33766 , \33624 );
or \U$33390 ( \33767 , \33765 , \33766 );
or \U$33391 ( \33768 , \33624 , \33617 );
nand \U$33392 ( \33769 , \33767 , \33768 );
not \U$33393 ( \33770 , \33769 );
xor \U$33394 ( \33771 , \33723 , \33725 );
xor \U$33395 ( \33772 , \33771 , \33751 );
not \U$33396 ( \33773 , \33772 );
or \U$33397 ( \33774 , \33770 , \33773 );
or \U$33398 ( \33775 , \33772 , \33769 );
or \U$33399 ( \33776 , \33641 , \33639 );
nand \U$33400 ( \33777 , \33776 , \33642 );
xor \U$33401 ( \33778 , \33631 , \33637 );
xor \U$33402 ( \33779 , \33777 , \33778 );
xor \U$33403 ( \33780 , \33670 , \33688 );
xor \U$33404 ( \33781 , \33780 , \33717 );
and \U$33405 ( \33782 , \33779 , \33781 );
and \U$33406 ( \33783 , \33777 , \33778 );
or \U$33407 ( \33784 , \33782 , \33783 );
and \U$33408 ( \33785 , \436 , RIae75470_8);
and \U$33409 ( \33786 , RIae76460_42, \434 );
nor \U$33410 ( \33787 , \33785 , \33786 );
not \U$33411 ( \33788 , \33787 );
not \U$33412 ( \33789 , \400 );
and \U$33413 ( \33790 , \33788 , \33789 );
and \U$33414 ( \33791 , \33787 , \400 );
nor \U$33415 ( \33792 , \33790 , \33791 );
not \U$33416 ( \33793 , \33792 );
and \U$33417 ( \33794 , \558 , RIae76640_46);
and \U$33418 ( \33795 , RIae76190_36, \556 );
nor \U$33419 ( \33796 , \33794 , \33795 );
and \U$33420 ( \33797 , \33796 , \562 );
not \U$33421 ( \33798 , \33796 );
and \U$33422 ( \33799 , \33798 , \504 );
nor \U$33423 ( \33800 , \33797 , \33799 );
not \U$33424 ( \33801 , \33800 );
and \U$33425 ( \33802 , \33793 , \33801 );
and \U$33426 ( \33803 , \33800 , \33792 );
and \U$33427 ( \33804 , \514 , RIae76550_44);
and \U$33428 ( \33805 , RIae76730_48, \512 );
nor \U$33429 ( \33806 , \33804 , \33805 );
not \U$33430 ( \33807 , \33806 );
not \U$33431 ( \33808 , \471 );
and \U$33432 ( \33809 , \33807 , \33808 );
and \U$33433 ( \33810 , \33806 , \469 );
nor \U$33434 ( \33811 , \33809 , \33810 );
nor \U$33435 ( \33812 , \33803 , \33811 );
nor \U$33436 ( \33813 , \33802 , \33812 );
and \U$33437 ( \33814 , \672 , RIae760a0_34);
and \U$33438 ( \33815 , RIae76370_40, \670 );
nor \U$33439 ( \33816 , \33814 , \33815 );
and \U$33440 ( \33817 , \33816 , \587 );
not \U$33441 ( \33818 , \33816 );
and \U$33442 ( \33819 , \33818 , \588 );
nor \U$33443 ( \33820 , \33817 , \33819 );
not \U$33444 ( \33821 , \33820 );
and \U$33445 ( \33822 , \1138 , RIae76a00_54);
and \U$33446 ( \33823 , RIae76820_50, \1136 );
nor \U$33447 ( \33824 , \33822 , \33823 );
and \U$33448 ( \33825 , \33824 , \1142 );
not \U$33449 ( \33826 , \33824 );
and \U$33450 ( \33827 , \33826 , \1012 );
nor \U$33451 ( \33828 , \33825 , \33827 );
not \U$33452 ( \33829 , \33828 );
and \U$33453 ( \33830 , \33821 , \33829 );
and \U$33454 ( \33831 , \33828 , \33820 );
and \U$33455 ( \33832 , \883 , RIae76280_38);
and \U$33456 ( \33833 , RIae76af0_56, \881 );
nor \U$33457 ( \33834 , \33832 , \33833 );
not \U$33458 ( \33835 , \33834 );
not \U$33459 ( \33836 , \789 );
and \U$33460 ( \33837 , \33835 , \33836 );
and \U$33461 ( \33838 , \33834 , \787 );
nor \U$33462 ( \33839 , \33837 , \33838 );
nor \U$33463 ( \33840 , \33831 , \33839 );
nor \U$33464 ( \33841 , \33830 , \33840 );
xor \U$33465 ( \33842 , \33813 , \33841 );
and \U$33466 ( \33843 , \1376 , RIae76910_52);
and \U$33467 ( \33844 , RIae76be0_58, \1374 );
nor \U$33468 ( \33845 , \33843 , \33844 );
and \U$33469 ( \33846 , \33845 , \1261 );
not \U$33470 ( \33847 , \33845 );
and \U$33471 ( \33848 , \33847 , \1380 );
nor \U$33472 ( \33849 , \33846 , \33848 );
not \U$33473 ( \33850 , \33849 );
and \U$33474 ( \33851 , \1593 , RIae78ad0_124);
and \U$33475 ( \33852 , RIae78d28_129, \1591 );
nor \U$33476 ( \33853 , \33851 , \33852 );
and \U$33477 ( \33854 , \33853 , \1488 );
not \U$33478 ( \33855 , \33853 );
and \U$33479 ( \33856 , \33855 , \1498 );
nor \U$33480 ( \33857 , \33854 , \33856 );
not \U$33481 ( \33858 , \33857 );
and \U$33482 ( \33859 , \33850 , \33858 );
and \U$33483 ( \33860 , \33857 , \33849 );
nand \U$33484 ( \33861 , RIae78e18_131, \1939 );
and \U$33485 ( \33862 , \33861 , \1734 );
not \U$33486 ( \33863 , \33861 );
and \U$33487 ( \33864 , \33863 , \1735 );
nor \U$33488 ( \33865 , \33862 , \33864 );
nor \U$33489 ( \33866 , \33860 , \33865 );
nor \U$33490 ( \33867 , \33859 , \33866 );
and \U$33491 ( \33868 , \33842 , \33867 );
and \U$33492 ( \33869 , \33813 , \33841 );
nor \U$33493 ( \33870 , \33868 , \33869 );
and \U$33494 ( \33871 , \384 , RIae75380_6);
and \U$33495 ( \33872 , RIae75470_8, \382 );
nor \U$33496 ( \33873 , \33871 , \33872 );
not \U$33497 ( \33874 , \33873 );
not \U$33498 ( \33875 , \388 );
and \U$33499 ( \33876 , \33874 , \33875 );
and \U$33500 ( \33877 , \33873 , \388 );
nor \U$33501 ( \33878 , \33876 , \33877 );
nand \U$33502 ( \33879 , RIae751a0_2, RIae78b48_125);
or \U$33503 ( \33880 , \33878 , \33879 );
not \U$33504 ( \33881 , \33879 );
not \U$33505 ( \33882 , \33878 );
or \U$33506 ( \33883 , \33881 , \33882 );
nand \U$33507 ( \33884 , RIae75290_4, RIae78b48_125);
and \U$33508 ( \33885 , \384 , RIae751a0_2);
and \U$33509 ( \33886 , RIae75380_6, \382 );
nor \U$33510 ( \33887 , \33885 , \33886 );
not \U$33511 ( \33888 , \33887 );
not \U$33512 ( \33889 , \388 );
and \U$33513 ( \33890 , \33888 , \33889 );
and \U$33514 ( \33891 , \33887 , \392 );
nor \U$33515 ( \33892 , \33890 , \33891 );
nand \U$33516 ( \33893 , \33884 , \33892 );
nand \U$33517 ( \33894 , \33883 , \33893 );
nand \U$33518 ( \33895 , \33880 , \33894 );
xor \U$33519 ( \33896 , \33870 , \33895 );
xor \U$33520 ( \33897 , \33651 , \33658 );
xor \U$33521 ( \33898 , \33897 , \33667 );
not \U$33522 ( \33899 , \33704 );
not \U$33523 ( \33900 , \33715 );
or \U$33524 ( \33901 , \33899 , \33900 );
or \U$33525 ( \33902 , \33704 , \33715 );
nand \U$33526 ( \33903 , \33901 , \33902 );
not \U$33527 ( \33904 , \33903 );
not \U$33528 ( \33905 , \33696 );
and \U$33529 ( \33906 , \33904 , \33905 );
and \U$33530 ( \33907 , \33903 , \33696 );
nor \U$33531 ( \33908 , \33906 , \33907 );
or \U$33532 ( \33909 , \33898 , \33908 );
not \U$33533 ( \33910 , \33908 );
not \U$33534 ( \33911 , \33898 );
or \U$33535 ( \33912 , \33910 , \33911 );
xor \U$33536 ( \33913 , \33677 , \1735 );
xor \U$33537 ( \33914 , \33913 , \33685 );
nand \U$33538 ( \33915 , \33912 , \33914 );
nand \U$33539 ( \33916 , \33909 , \33915 );
and \U$33540 ( \33917 , \33896 , \33916 );
and \U$33541 ( \33918 , \33870 , \33895 );
or \U$33542 ( \33919 , \33917 , \33918 );
xor \U$33543 ( \33920 , \33784 , \33919 );
xor \U$33544 ( \33921 , \33732 , \33741 );
xor \U$33545 ( \33922 , \33921 , \33748 );
and \U$33546 ( \33923 , \33920 , \33922 );
and \U$33547 ( \33924 , \33784 , \33919 );
or \U$33548 ( \33925 , \33923 , \33924 );
nand \U$33549 ( \33926 , \33775 , \33925 );
nand \U$33550 ( \33927 , \33774 , \33926 );
not \U$33551 ( \33928 , \33927 );
not \U$33552 ( \33929 , \33625 );
not \U$33553 ( \33930 , \33754 );
or \U$33554 ( \33931 , \33929 , \33930 );
or \U$33555 ( \33932 , \33754 , \33625 );
nand \U$33556 ( \33933 , \33931 , \33932 );
not \U$33557 ( \33934 , \33933 );
not \U$33558 ( \33935 , \33615 );
and \U$33559 ( \33936 , \33934 , \33935 );
and \U$33560 ( \33937 , \33933 , \33615 );
nor \U$33561 ( \33938 , \33936 , \33937 );
nor \U$33562 ( \33939 , \33928 , \33938 );
and \U$33563 ( \33940 , \33764 , \33939 );
xor \U$33564 ( \33941 , \33939 , \33764 );
not \U$33565 ( \33942 , \33927 );
not \U$33566 ( \33943 , \33938 );
and \U$33567 ( \33944 , \33942 , \33943 );
and \U$33568 ( \33945 , \33927 , \33938 );
nor \U$33569 ( \33946 , \33944 , \33945 );
xnor \U$33570 ( \33947 , \33925 , \33772 );
not \U$33571 ( \33948 , \33947 );
not \U$33572 ( \33949 , \33769 );
and \U$33573 ( \33950 , \33948 , \33949 );
and \U$33574 ( \33951 , \33947 , \33769 );
nor \U$33575 ( \33952 , \33950 , \33951 );
not \U$33576 ( \33953 , \33952 );
not \U$33577 ( \33954 , \33878 );
not \U$33578 ( \33955 , \33893 );
or \U$33579 ( \33956 , \33954 , \33955 );
or \U$33580 ( \33957 , \33893 , \33878 );
nand \U$33581 ( \33958 , \33956 , \33957 );
not \U$33582 ( \33959 , \33958 );
not \U$33583 ( \33960 , \33879 );
and \U$33584 ( \33961 , \33959 , \33960 );
and \U$33585 ( \33962 , \33958 , \33879 );
nor \U$33586 ( \33963 , \33961 , \33962 );
xor \U$33587 ( \33964 , \33813 , \33841 );
xor \U$33588 ( \33965 , \33964 , \33867 );
xor \U$33589 ( \33966 , \33963 , \33965 );
not \U$33590 ( \33967 , \33908 );
not \U$33591 ( \33968 , \33914 );
or \U$33592 ( \33969 , \33967 , \33968 );
or \U$33593 ( \33970 , \33914 , \33908 );
nand \U$33594 ( \33971 , \33969 , \33970 );
not \U$33595 ( \33972 , \33971 );
not \U$33596 ( \33973 , \33898 );
and \U$33597 ( \33974 , \33972 , \33973 );
and \U$33598 ( \33975 , \33971 , \33898 );
nor \U$33599 ( \33976 , \33974 , \33975 );
and \U$33600 ( \33977 , \33966 , \33976 );
and \U$33601 ( \33978 , \33963 , \33965 );
nor \U$33602 ( \33979 , \33977 , \33978 );
not \U$33603 ( \33980 , \33820 );
xor \U$33604 ( \33981 , \33839 , \33828 );
not \U$33605 ( \33982 , \33981 );
or \U$33606 ( \33983 , \33980 , \33982 );
or \U$33607 ( \33984 , \33981 , \33820 );
nand \U$33608 ( \33985 , \33983 , \33984 );
not \U$33609 ( \33986 , \33849 );
xor \U$33610 ( \33987 , \33865 , \33857 );
not \U$33611 ( \33988 , \33987 );
or \U$33612 ( \33989 , \33986 , \33988 );
or \U$33613 ( \33990 , \33987 , \33849 );
nand \U$33614 ( \33991 , \33989 , \33990 );
and \U$33615 ( \33992 , \33985 , \33991 );
not \U$33616 ( \33993 , \33992 );
and \U$33617 ( \33994 , \558 , RIae76730_48);
and \U$33618 ( \33995 , RIae76640_46, \556 );
nor \U$33619 ( \33996 , \33994 , \33995 );
and \U$33620 ( \33997 , \33996 , \562 );
not \U$33621 ( \33998 , \33996 );
and \U$33622 ( \33999 , \33998 , \504 );
nor \U$33623 ( \34000 , \33997 , \33999 );
and \U$33624 ( \34001 , \672 , RIae76190_36);
and \U$33625 ( \34002 , RIae760a0_34, \670 );
nor \U$33626 ( \34003 , \34001 , \34002 );
and \U$33627 ( \34004 , \34003 , \587 );
not \U$33628 ( \34005 , \34003 );
and \U$33629 ( \34006 , \34005 , \588 );
nor \U$33630 ( \34007 , \34004 , \34006 );
xor \U$33631 ( \34008 , \34000 , \34007 );
and \U$33632 ( \34009 , \514 , RIae76460_42);
and \U$33633 ( \34010 , RIae76550_44, \512 );
nor \U$33634 ( \34011 , \34009 , \34010 );
not \U$33635 ( \34012 , \34011 );
not \U$33636 ( \34013 , \471 );
and \U$33637 ( \34014 , \34012 , \34013 );
and \U$33638 ( \34015 , \34011 , \469 );
nor \U$33639 ( \34016 , \34014 , \34015 );
and \U$33640 ( \34017 , \34008 , \34016 );
and \U$33641 ( \34018 , \34000 , \34007 );
nor \U$33642 ( \34019 , \34017 , \34018 );
and \U$33643 ( \34020 , \1939 , RIae78d28_129);
and \U$33644 ( \34021 , RIae78e18_131, \1937 );
nor \U$33645 ( \34022 , \34020 , \34021 );
and \U$33646 ( \34023 , \34022 , \1734 );
not \U$33647 ( \34024 , \34022 );
and \U$33648 ( \34025 , \34024 , \1735 );
nor \U$33649 ( \34026 , \34023 , \34025 );
or \U$33650 ( \34027 , \34026 , \2060 );
and \U$33651 ( \34028 , \34026 , \2060 );
and \U$33652 ( \34029 , \1593 , RIae76be0_58);
and \U$33653 ( \34030 , RIae78ad0_124, \1591 );
nor \U$33654 ( \34031 , \34029 , \34030 );
and \U$33655 ( \34032 , \34031 , \1488 );
not \U$33656 ( \34033 , \34031 );
and \U$33657 ( \34034 , \34033 , \1498 );
nor \U$33658 ( \34035 , \34032 , \34034 );
nor \U$33659 ( \34036 , \34028 , \34035 );
not \U$33660 ( \34037 , \34036 );
nand \U$33661 ( \34038 , \34027 , \34037 );
xor \U$33662 ( \34039 , \34019 , \34038 );
not \U$33663 ( \34040 , \787 );
and \U$33664 ( \34041 , \883 , RIae76370_40);
and \U$33665 ( \34042 , RIae76280_38, \881 );
nor \U$33666 ( \34043 , \34041 , \34042 );
not \U$33667 ( \34044 , \34043 );
or \U$33668 ( \34045 , \34040 , \34044 );
or \U$33669 ( \34046 , \34043 , \789 );
nand \U$33670 ( \34047 , \34045 , \34046 );
and \U$33671 ( \34048 , \1138 , RIae76af0_56);
and \U$33672 ( \34049 , RIae76a00_54, \1136 );
nor \U$33673 ( \34050 , \34048 , \34049 );
and \U$33674 ( \34051 , \34050 , \1012 );
not \U$33675 ( \34052 , \34050 );
and \U$33676 ( \34053 , \34052 , \1142 );
nor \U$33677 ( \34054 , \34051 , \34053 );
xor \U$33678 ( \34055 , \34047 , \34054 );
and \U$33679 ( \34056 , \1376 , RIae76820_50);
and \U$33680 ( \34057 , RIae76910_52, \1374 );
nor \U$33681 ( \34058 , \34056 , \34057 );
and \U$33682 ( \34059 , \34058 , \1380 );
not \U$33683 ( \34060 , \34058 );
and \U$33684 ( \34061 , \34060 , \1261 );
nor \U$33685 ( \34062 , \34059 , \34061 );
and \U$33686 ( \34063 , \34055 , \34062 );
and \U$33687 ( \34064 , \34047 , \34054 );
or \U$33688 ( \34065 , \34063 , \34064 );
and \U$33689 ( \34066 , \34039 , \34065 );
and \U$33690 ( \34067 , \34019 , \34038 );
or \U$33691 ( \34068 , \34066 , \34067 );
not \U$33692 ( \34069 , \34068 );
or \U$33693 ( \34070 , \33993 , \34069 );
or \U$33694 ( \34071 , \34068 , \33992 );
and \U$33695 ( \34072 , \436 , RIae75380_6);
and \U$33696 ( \34073 , RIae75470_8, \434 );
nor \U$33697 ( \34074 , \34072 , \34073 );
not \U$33698 ( \34075 , \34074 );
not \U$33699 ( \34076 , \400 );
and \U$33700 ( \34077 , \34075 , \34076 );
and \U$33701 ( \34078 , \34074 , \402 );
nor \U$33702 ( \34079 , \34077 , \34078 );
nand \U$33703 ( \34080 , RIae75740_14, RIae78b48_125);
or \U$33704 ( \34081 , \34079 , \34080 );
not \U$33705 ( \34082 , \34080 );
not \U$33706 ( \34083 , \34079 );
or \U$33707 ( \34084 , \34082 , \34083 );
not \U$33708 ( \34085 , \388 );
and \U$33709 ( \34086 , \384 , RIae75290_4);
and \U$33710 ( \34087 , RIae751a0_2, \382 );
nor \U$33711 ( \34088 , \34086 , \34087 );
not \U$33712 ( \34089 , \34088 );
or \U$33713 ( \34090 , \34085 , \34089 );
or \U$33714 ( \34091 , \34088 , \392 );
nand \U$33715 ( \34092 , \34090 , \34091 );
nand \U$33716 ( \34093 , \34084 , \34092 );
nand \U$33717 ( \34094 , \34081 , \34093 );
or \U$33718 ( \34095 , \33892 , \33884 );
nand \U$33719 ( \34096 , \34095 , \33893 );
xor \U$33720 ( \34097 , \34094 , \34096 );
not \U$33721 ( \34098 , \33792 );
xor \U$33722 ( \34099 , \33811 , \33800 );
not \U$33723 ( \34100 , \34099 );
or \U$33724 ( \34101 , \34098 , \34100 );
or \U$33725 ( \34102 , \34099 , \33792 );
nand \U$33726 ( \34103 , \34101 , \34102 );
and \U$33727 ( \34104 , \34097 , \34103 );
and \U$33728 ( \34105 , \34094 , \34096 );
or \U$33729 ( \34106 , \34104 , \34105 );
nand \U$33730 ( \34107 , \34071 , \34106 );
nand \U$33731 ( \34108 , \34070 , \34107 );
xor \U$33732 ( \34109 , \33979 , \34108 );
xor \U$33733 ( \34110 , \33777 , \33778 );
xor \U$33734 ( \34111 , \34110 , \33781 );
and \U$33735 ( \34112 , \34109 , \34111 );
and \U$33736 ( \34113 , \33979 , \34108 );
or \U$33737 ( \34114 , \34112 , \34113 );
xor \U$33738 ( \34115 , \33638 , \33642 );
xor \U$33739 ( \34116 , \34115 , \33720 );
xor \U$33740 ( \34117 , \34114 , \34116 );
xor \U$33741 ( \34118 , \33784 , \33919 );
xor \U$33742 ( \34119 , \34118 , \33922 );
and \U$33743 ( \34120 , \34117 , \34119 );
and \U$33744 ( \34121 , \34114 , \34116 );
or \U$33745 ( \34122 , \34120 , \34121 );
nand \U$33746 ( \34123 , \33953 , \34122 );
or \U$33747 ( \34124 , \33946 , \34123 );
xnor \U$33748 ( \34125 , \33946 , \34123 );
not \U$33749 ( \34126 , \34122 );
not \U$33750 ( \34127 , \33952 );
or \U$33751 ( \34128 , \34126 , \34127 );
or \U$33752 ( \34129 , \33952 , \34122 );
nand \U$33753 ( \34130 , \34128 , \34129 );
xor \U$33754 ( \34131 , \34114 , \34116 );
xor \U$33755 ( \34132 , \34131 , \34119 );
not \U$33756 ( \34133 , \34132 );
xor \U$33757 ( \34134 , \33963 , \33965 );
xor \U$33758 ( \34135 , \34134 , \33976 );
and \U$33759 ( \34136 , \558 , RIae76550_44);
and \U$33760 ( \34137 , RIae76730_48, \556 );
nor \U$33761 ( \34138 , \34136 , \34137 );
and \U$33762 ( \34139 , \34138 , \504 );
not \U$33763 ( \34140 , \34138 );
and \U$33764 ( \34141 , \34140 , \562 );
nor \U$33765 ( \34142 , \34139 , \34141 );
and \U$33766 ( \34143 , \672 , RIae76640_46);
and \U$33767 ( \34144 , RIae76190_36, \670 );
nor \U$33768 ( \34145 , \34143 , \34144 );
and \U$33769 ( \34146 , \34145 , \588 );
not \U$33770 ( \34147 , \34145 );
and \U$33771 ( \34148 , \34147 , \587 );
nor \U$33772 ( \34149 , \34146 , \34148 );
xor \U$33773 ( \34150 , \34142 , \34149 );
not \U$33774 ( \34151 , \469 );
and \U$33775 ( \34152 , \514 , RIae75470_8);
and \U$33776 ( \34153 , RIae76460_42, \512 );
nor \U$33777 ( \34154 , \34152 , \34153 );
not \U$33778 ( \34155 , \34154 );
or \U$33779 ( \34156 , \34151 , \34155 );
or \U$33780 ( \34157 , \34154 , \469 );
nand \U$33781 ( \34158 , \34156 , \34157 );
and \U$33782 ( \34159 , \34150 , \34158 );
and \U$33783 ( \34160 , \34142 , \34149 );
nor \U$33784 ( \34161 , \34159 , \34160 );
and \U$33785 ( \34162 , \1593 , RIae76910_52);
and \U$33786 ( \34163 , RIae76be0_58, \1591 );
nor \U$33787 ( \34164 , \34162 , \34163 );
and \U$33788 ( \34165 , \34164 , \1488 );
not \U$33789 ( \34166 , \34164 );
and \U$33790 ( \34167 , \34166 , \1498 );
nor \U$33791 ( \34168 , \34165 , \34167 );
not \U$33792 ( \34169 , \34168 );
and \U$33793 ( \34170 , \1939 , RIae78ad0_124);
and \U$33794 ( \34171 , RIae78d28_129, \1937 );
nor \U$33795 ( \34172 , \34170 , \34171 );
and \U$33796 ( \34173 , \34172 , \1734 );
not \U$33797 ( \34174 , \34172 );
and \U$33798 ( \34175 , \34174 , \1735 );
nor \U$33799 ( \34176 , \34173 , \34175 );
not \U$33800 ( \34177 , \34176 );
and \U$33801 ( \34178 , \34169 , \34177 );
and \U$33802 ( \34179 , \34176 , \34168 );
nand \U$33803 ( \34180 , RIae78e18_131, \2224 );
and \U$33804 ( \34181 , \34180 , \2060 );
not \U$33805 ( \34182 , \34180 );
and \U$33806 ( \34183 , \34182 , \2061 );
nor \U$33807 ( \34184 , \34181 , \34183 );
nor \U$33808 ( \34185 , \34179 , \34184 );
nor \U$33809 ( \34186 , \34178 , \34185 );
xor \U$33810 ( \34187 , \34161 , \34186 );
and \U$33811 ( \34188 , \883 , RIae760a0_34);
and \U$33812 ( \34189 , RIae76370_40, \881 );
nor \U$33813 ( \34190 , \34188 , \34189 );
not \U$33814 ( \34191 , \34190 );
not \U$33815 ( \34192 , \789 );
and \U$33816 ( \34193 , \34191 , \34192 );
and \U$33817 ( \34194 , \34190 , \789 );
nor \U$33818 ( \34195 , \34193 , \34194 );
not \U$33819 ( \34196 , \34195 );
and \U$33820 ( \34197 , \1138 , RIae76280_38);
and \U$33821 ( \34198 , RIae76af0_56, \1136 );
nor \U$33822 ( \34199 , \34197 , \34198 );
and \U$33823 ( \34200 , \34199 , \1142 );
not \U$33824 ( \34201 , \34199 );
and \U$33825 ( \34202 , \34201 , \1012 );
nor \U$33826 ( \34203 , \34200 , \34202 );
not \U$33827 ( \34204 , \34203 );
and \U$33828 ( \34205 , \34196 , \34204 );
and \U$33829 ( \34206 , \34203 , \34195 );
and \U$33830 ( \34207 , \1376 , RIae76a00_54);
and \U$33831 ( \34208 , RIae76820_50, \1374 );
nor \U$33832 ( \34209 , \34207 , \34208 );
and \U$33833 ( \34210 , \34209 , \1261 );
not \U$33834 ( \34211 , \34209 );
and \U$33835 ( \34212 , \34211 , \1380 );
nor \U$33836 ( \34213 , \34210 , \34212 );
nor \U$33837 ( \34214 , \34206 , \34213 );
nor \U$33838 ( \34215 , \34205 , \34214 );
and \U$33839 ( \34216 , \34187 , \34215 );
and \U$33840 ( \34217 , \34161 , \34186 );
or \U$33841 ( \34218 , \34216 , \34217 );
and \U$33842 ( \34219 , \34026 , \2060 );
not \U$33843 ( \34220 , \34026 );
and \U$33844 ( \34221 , \34220 , \2061 );
nor \U$33845 ( \34222 , \34219 , \34221 );
not \U$33846 ( \34223 , \34222 );
not \U$33847 ( \34224 , \34035 );
and \U$33848 ( \34225 , \34223 , \34224 );
and \U$33849 ( \34226 , \34222 , \34035 );
nor \U$33850 ( \34227 , \34225 , \34226 );
not \U$33851 ( \34228 , \34227 );
xor \U$33852 ( \34229 , \34047 , \34054 );
xor \U$33853 ( \34230 , \34229 , \34062 );
nand \U$33854 ( \34231 , \34228 , \34230 );
xor \U$33855 ( \34232 , \34218 , \34231 );
not \U$33856 ( \34233 , \34079 );
not \U$33857 ( \34234 , \34092 );
or \U$33858 ( \34235 , \34233 , \34234 );
or \U$33859 ( \34236 , \34079 , \34092 );
nand \U$33860 ( \34237 , \34235 , \34236 );
not \U$33861 ( \34238 , \34237 );
not \U$33862 ( \34239 , \34080 );
and \U$33863 ( \34240 , \34238 , \34239 );
and \U$33864 ( \34241 , \34237 , \34080 );
nor \U$33865 ( \34242 , \34240 , \34241 );
and \U$33866 ( \34243 , \384 , RIae75740_14);
and \U$33867 ( \34244 , RIae75290_4, \382 );
nor \U$33868 ( \34245 , \34243 , \34244 );
not \U$33869 ( \34246 , \34245 );
not \U$33870 ( \34247 , \388 );
and \U$33871 ( \34248 , \34246 , \34247 );
and \U$33872 ( \34249 , \34245 , \392 );
nor \U$33873 ( \34250 , \34248 , \34249 );
nand \U$33874 ( \34251 , RIae75830_16, RIae78b48_125);
xor \U$33875 ( \34252 , \34250 , \34251 );
and \U$33876 ( \34253 , \436 , RIae751a0_2);
and \U$33877 ( \34254 , RIae75380_6, \434 );
nor \U$33878 ( \34255 , \34253 , \34254 );
not \U$33879 ( \34256 , \34255 );
not \U$33880 ( \34257 , \402 );
and \U$33881 ( \34258 , \34256 , \34257 );
and \U$33882 ( \34259 , \34255 , \400 );
nor \U$33883 ( \34260 , \34258 , \34259 );
and \U$33884 ( \34261 , \34252 , \34260 );
and \U$33885 ( \34262 , \34250 , \34251 );
or \U$33886 ( \34263 , \34261 , \34262 );
xor \U$33887 ( \34264 , \34242 , \34263 );
xor \U$33888 ( \34265 , \34000 , \34007 );
xor \U$33889 ( \34266 , \34265 , \34016 );
and \U$33890 ( \34267 , \34264 , \34266 );
and \U$33891 ( \34268 , \34242 , \34263 );
or \U$33892 ( \34269 , \34267 , \34268 );
and \U$33893 ( \34270 , \34232 , \34269 );
and \U$33894 ( \34271 , \34218 , \34231 );
or \U$33895 ( \34272 , \34270 , \34271 );
or \U$33896 ( \34273 , \34135 , \34272 );
not \U$33897 ( \34274 , \34272 );
not \U$33898 ( \34275 , \34135 );
or \U$33899 ( \34276 , \34274 , \34275 );
xor \U$33900 ( \34277 , \33985 , \33991 );
not \U$33901 ( \34278 , \34277 );
xor \U$33902 ( \34279 , \34019 , \34038 );
xor \U$33903 ( \34280 , \34279 , \34065 );
not \U$33904 ( \34281 , \34280 );
or \U$33905 ( \34282 , \34278 , \34281 );
or \U$33906 ( \34283 , \34280 , \34277 );
xor \U$33907 ( \34284 , \34094 , \34096 );
xor \U$33908 ( \34285 , \34284 , \34103 );
nand \U$33909 ( \34286 , \34283 , \34285 );
nand \U$33910 ( \34287 , \34282 , \34286 );
nand \U$33911 ( \34288 , \34276 , \34287 );
nand \U$33912 ( \34289 , \34273 , \34288 );
xor \U$33913 ( \34290 , \33870 , \33895 );
xor \U$33914 ( \34291 , \34290 , \33916 );
and \U$33915 ( \34292 , \34289 , \34291 );
xor \U$33916 ( \34293 , \33979 , \34108 );
xor \U$33917 ( \34294 , \34293 , \34111 );
or \U$33918 ( \34295 , \34289 , \34291 );
and \U$33919 ( \34296 , \34294 , \34295 );
nor \U$33920 ( \34297 , \34292 , \34296 );
nor \U$33921 ( \34298 , \34133 , \34297 );
and \U$33922 ( \34299 , \34130 , \34298 );
xor \U$33923 ( \34300 , \34298 , \34130 );
not \U$33924 ( \34301 , \34132 );
not \U$33925 ( \34302 , \34297 );
and \U$33926 ( \34303 , \34301 , \34302 );
and \U$33927 ( \34304 , \34132 , \34297 );
nor \U$33928 ( \34305 , \34303 , \34304 );
not \U$33929 ( \34306 , \34272 );
not \U$33930 ( \34307 , \34287 );
or \U$33931 ( \34308 , \34306 , \34307 );
or \U$33932 ( \34309 , \34287 , \34272 );
nand \U$33933 ( \34310 , \34308 , \34309 );
not \U$33934 ( \34311 , \34310 );
not \U$33935 ( \34312 , \34135 );
and \U$33936 ( \34313 , \34311 , \34312 );
and \U$33937 ( \34314 , \34310 , \34135 );
nor \U$33938 ( \34315 , \34313 , \34314 );
not \U$33939 ( \34316 , \34315 );
xnor \U$33940 ( \34317 , \34068 , \34106 );
not \U$33941 ( \34318 , \34317 );
not \U$33942 ( \34319 , \33992 );
and \U$33943 ( \34320 , \34318 , \34319 );
and \U$33944 ( \34321 , \34317 , \33992 );
nor \U$33945 ( \34322 , \34320 , \34321 );
not \U$33946 ( \34323 , \34322 );
and \U$33947 ( \34324 , \34316 , \34323 );
and \U$33948 ( \34325 , \34315 , \34322 );
not \U$33949 ( \34326 , \34227 );
not \U$33950 ( \34327 , \34230 );
and \U$33951 ( \34328 , \34326 , \34327 );
and \U$33952 ( \34329 , \34227 , \34230 );
nor \U$33953 ( \34330 , \34328 , \34329 );
xor \U$33954 ( \34331 , \34161 , \34186 );
xor \U$33955 ( \34332 , \34331 , \34215 );
and \U$33956 ( \34333 , \34330 , \34332 );
xor \U$33957 ( \34334 , \34242 , \34263 );
xor \U$33958 ( \34335 , \34334 , \34266 );
xor \U$33959 ( \34336 , \34161 , \34186 );
xor \U$33960 ( \34337 , \34336 , \34215 );
and \U$33961 ( \34338 , \34335 , \34337 );
and \U$33962 ( \34339 , \34330 , \34335 );
or \U$33963 ( \34340 , \34333 , \34338 , \34339 );
xor \U$33964 ( \34341 , \34142 , \34149 );
xor \U$33965 ( \34342 , \34341 , \34158 );
not \U$33966 ( \34343 , \34168 );
xor \U$33967 ( \34344 , \34184 , \34176 );
not \U$33968 ( \34345 , \34344 );
or \U$33969 ( \34346 , \34343 , \34345 );
or \U$33970 ( \34347 , \34344 , \34168 );
nand \U$33971 ( \34348 , \34346 , \34347 );
xor \U$33972 ( \34349 , \34342 , \34348 );
not \U$33973 ( \34350 , \34195 );
xor \U$33974 ( \34351 , \34203 , \34213 );
not \U$33975 ( \34352 , \34351 );
or \U$33976 ( \34353 , \34350 , \34352 );
or \U$33977 ( \34354 , \34351 , \34195 );
nand \U$33978 ( \34355 , \34353 , \34354 );
and \U$33979 ( \34356 , \34349 , \34355 );
and \U$33980 ( \34357 , \34342 , \34348 );
or \U$33981 ( \34358 , \34356 , \34357 );
and \U$33982 ( \34359 , \384 , RIae75830_16);
and \U$33983 ( \34360 , RIae75740_14, \382 );
nor \U$33984 ( \34361 , \34359 , \34360 );
not \U$33985 ( \34362 , \34361 );
not \U$33986 ( \34363 , \388 );
and \U$33987 ( \34364 , \34362 , \34363 );
and \U$33988 ( \34365 , \34361 , \392 );
nor \U$33989 ( \34366 , \34364 , \34365 );
not \U$33990 ( \34367 , \34366 );
and \U$33991 ( \34368 , \436 , RIae75290_4);
and \U$33992 ( \34369 , RIae751a0_2, \434 );
nor \U$33993 ( \34370 , \34368 , \34369 );
not \U$33994 ( \34371 , \34370 );
not \U$33995 ( \34372 , \402 );
and \U$33996 ( \34373 , \34371 , \34372 );
and \U$33997 ( \34374 , \34370 , \400 );
nor \U$33998 ( \34375 , \34373 , \34374 );
not \U$33999 ( \34376 , \34375 );
and \U$34000 ( \34377 , \34367 , \34376 );
and \U$34001 ( \34378 , \34375 , \34366 );
and \U$34002 ( \34379 , \514 , RIae75380_6);
and \U$34003 ( \34380 , RIae75470_8, \512 );
nor \U$34004 ( \34381 , \34379 , \34380 );
not \U$34005 ( \34382 , \34381 );
not \U$34006 ( \34383 , \469 );
and \U$34007 ( \34384 , \34382 , \34383 );
and \U$34008 ( \34385 , \34381 , \469 );
nor \U$34009 ( \34386 , \34384 , \34385 );
nor \U$34010 ( \34387 , \34378 , \34386 );
nor \U$34011 ( \34388 , \34377 , \34387 );
xor \U$34012 ( \34389 , \34250 , \34251 );
xor \U$34013 ( \34390 , \34389 , \34260 );
nand \U$34014 ( \34391 , \34388 , \34390 );
and \U$34015 ( \34392 , \34358 , \34391 );
not \U$34016 ( \34393 , \34358 );
not \U$34017 ( \34394 , \34391 );
and \U$34018 ( \34395 , \34393 , \34394 );
and \U$34019 ( \34396 , \1138 , RIae76370_40);
and \U$34020 ( \34397 , RIae76280_38, \1136 );
nor \U$34021 ( \34398 , \34396 , \34397 );
and \U$34022 ( \34399 , \34398 , \1012 );
not \U$34023 ( \34400 , \34398 );
and \U$34024 ( \34401 , \34400 , \1142 );
nor \U$34025 ( \34402 , \34399 , \34401 );
and \U$34026 ( \34403 , \1376 , RIae76af0_56);
and \U$34027 ( \34404 , RIae76a00_54, \1374 );
nor \U$34028 ( \34405 , \34403 , \34404 );
and \U$34029 ( \34406 , \34405 , \1380 );
not \U$34030 ( \34407 , \34405 );
and \U$34031 ( \34408 , \34407 , \1261 );
nor \U$34032 ( \34409 , \34406 , \34408 );
xor \U$34033 ( \34410 , \34402 , \34409 );
and \U$34034 ( \34411 , \1593 , RIae76820_50);
and \U$34035 ( \34412 , RIae76910_52, \1591 );
nor \U$34036 ( \34413 , \34411 , \34412 );
and \U$34037 ( \34414 , \34413 , \1498 );
not \U$34038 ( \34415 , \34413 );
and \U$34039 ( \34416 , \34415 , \1488 );
nor \U$34040 ( \34417 , \34414 , \34416 );
and \U$34041 ( \34418 , \34410 , \34417 );
and \U$34042 ( \34419 , \34402 , \34409 );
or \U$34043 ( \34420 , \34418 , \34419 );
and \U$34044 ( \34421 , \2224 , RIae78d28_129);
and \U$34045 ( \34422 , RIae78e18_131, \2222 );
nor \U$34046 ( \34423 , \34421 , \34422 );
and \U$34047 ( \34424 , \34423 , \2061 );
not \U$34048 ( \34425 , \34423 );
and \U$34049 ( \34426 , \34425 , \2060 );
nor \U$34050 ( \34427 , \34424 , \34426 );
xor \U$34051 ( \34428 , \34427 , \2611 );
and \U$34052 ( \34429 , \1939 , RIae76be0_58);
and \U$34053 ( \34430 , RIae78ad0_124, \1937 );
nor \U$34054 ( \34431 , \34429 , \34430 );
and \U$34055 ( \34432 , \34431 , \1735 );
not \U$34056 ( \34433 , \34431 );
and \U$34057 ( \34434 , \34433 , \1734 );
nor \U$34058 ( \34435 , \34432 , \34434 );
and \U$34059 ( \34436 , \34428 , \34435 );
and \U$34060 ( \34437 , \34427 , \2611 );
or \U$34061 ( \34438 , \34436 , \34437 );
xor \U$34062 ( \34439 , \34420 , \34438 );
not \U$34063 ( \34440 , \789 );
and \U$34064 ( \34441 , \883 , RIae76190_36);
and \U$34065 ( \34442 , RIae760a0_34, \881 );
nor \U$34066 ( \34443 , \34441 , \34442 );
not \U$34067 ( \34444 , \34443 );
or \U$34068 ( \34445 , \34440 , \34444 );
or \U$34069 ( \34446 , \34443 , \787 );
nand \U$34070 ( \34447 , \34445 , \34446 );
and \U$34071 ( \34448 , \558 , RIae76460_42);
and \U$34072 ( \34449 , RIae76550_44, \556 );
nor \U$34073 ( \34450 , \34448 , \34449 );
and \U$34074 ( \34451 , \34450 , \504 );
not \U$34075 ( \34452 , \34450 );
and \U$34076 ( \34453 , \34452 , \562 );
nor \U$34077 ( \34454 , \34451 , \34453 );
xor \U$34078 ( \34455 , \34447 , \34454 );
and \U$34079 ( \34456 , \672 , RIae76730_48);
and \U$34080 ( \34457 , RIae76640_46, \670 );
nor \U$34081 ( \34458 , \34456 , \34457 );
and \U$34082 ( \34459 , \34458 , \588 );
not \U$34083 ( \34460 , \34458 );
and \U$34084 ( \34461 , \34460 , \587 );
nor \U$34085 ( \34462 , \34459 , \34461 );
and \U$34086 ( \34463 , \34455 , \34462 );
and \U$34087 ( \34464 , \34447 , \34454 );
or \U$34088 ( \34465 , \34463 , \34464 );
and \U$34089 ( \34466 , \34439 , \34465 );
and \U$34090 ( \34467 , \34420 , \34438 );
nor \U$34091 ( \34468 , \34466 , \34467 );
nor \U$34092 ( \34469 , \34395 , \34468 );
nor \U$34093 ( \34470 , \34392 , \34469 );
xor \U$34094 ( \34471 , \34340 , \34470 );
xnor \U$34095 ( \34472 , \34280 , \34285 );
not \U$34096 ( \34473 , \34472 );
not \U$34097 ( \34474 , \34277 );
and \U$34098 ( \34475 , \34473 , \34474 );
and \U$34099 ( \34476 , \34472 , \34277 );
nor \U$34100 ( \34477 , \34475 , \34476 );
and \U$34101 ( \34478 , \34471 , \34477 );
and \U$34102 ( \34479 , \34340 , \34470 );
or \U$34103 ( \34480 , \34478 , \34479 );
nor \U$34104 ( \34481 , \34325 , \34480 );
nor \U$34105 ( \34482 , \34324 , \34481 );
not \U$34106 ( \34483 , \34482 );
not \U$34107 ( \34484 , \34294 );
xnor \U$34108 ( \34485 , \34291 , \34289 );
not \U$34109 ( \34486 , \34485 );
or \U$34110 ( \34487 , \34484 , \34486 );
or \U$34111 ( \34488 , \34485 , \34294 );
nand \U$34112 ( \34489 , \34487 , \34488 );
nand \U$34113 ( \34490 , \34483 , \34489 );
or \U$34114 ( \34491 , \34305 , \34490 );
xnor \U$34115 ( \34492 , \34490 , \34305 );
not \U$34116 ( \34493 , \34482 );
not \U$34117 ( \34494 , \34489 );
or \U$34118 ( \34495 , \34493 , \34494 );
or \U$34119 ( \34496 , \34489 , \34482 );
nand \U$34120 ( \34497 , \34495 , \34496 );
not \U$34121 ( \34498 , \34315 );
xor \U$34122 ( \34499 , \34322 , \34480 );
not \U$34123 ( \34500 , \34499 );
or \U$34124 ( \34501 , \34498 , \34500 );
or \U$34125 ( \34502 , \34499 , \34315 );
nand \U$34126 ( \34503 , \34501 , \34502 );
not \U$34127 ( \34504 , \34503 );
xor \U$34128 ( \34505 , \34161 , \34186 );
xor \U$34129 ( \34506 , \34505 , \34215 );
xor \U$34130 ( \34507 , \34330 , \34335 );
xor \U$34131 ( \34508 , \34506 , \34507 );
not \U$34132 ( \34509 , \34508 );
and \U$34133 ( \34510 , \1138 , RIae760a0_34);
and \U$34134 ( \34511 , RIae76370_40, \1136 );
nor \U$34135 ( \34512 , \34510 , \34511 );
and \U$34136 ( \34513 , \34512 , \1142 );
not \U$34137 ( \34514 , \34512 );
and \U$34138 ( \34515 , \34514 , \1012 );
nor \U$34139 ( \34516 , \34513 , \34515 );
not \U$34140 ( \34517 , \34516 );
and \U$34141 ( \34518 , \1593 , RIae76a00_54);
and \U$34142 ( \34519 , RIae76820_50, \1591 );
nor \U$34143 ( \34520 , \34518 , \34519 );
and \U$34144 ( \34521 , \34520 , \1488 );
not \U$34145 ( \34522 , \34520 );
and \U$34146 ( \34523 , \34522 , \1498 );
nor \U$34147 ( \34524 , \34521 , \34523 );
not \U$34148 ( \34525 , \34524 );
and \U$34149 ( \34526 , \34517 , \34525 );
and \U$34150 ( \34527 , \34524 , \34516 );
and \U$34151 ( \34528 , \1376 , RIae76280_38);
and \U$34152 ( \34529 , RIae76af0_56, \1374 );
nor \U$34153 ( \34530 , \34528 , \34529 );
and \U$34154 ( \34531 , \34530 , \1261 );
not \U$34155 ( \34532 , \34530 );
and \U$34156 ( \34533 , \34532 , \1380 );
nor \U$34157 ( \34534 , \34531 , \34533 );
nor \U$34158 ( \34535 , \34527 , \34534 );
nor \U$34159 ( \34536 , \34526 , \34535 );
and \U$34160 ( \34537 , \1939 , RIae76910_52);
and \U$34161 ( \34538 , RIae76be0_58, \1937 );
nor \U$34162 ( \34539 , \34537 , \34538 );
and \U$34163 ( \34540 , \34539 , \1734 );
not \U$34164 ( \34541 , \34539 );
and \U$34165 ( \34542 , \34541 , \1735 );
nor \U$34166 ( \34543 , \34540 , \34542 );
not \U$34167 ( \34544 , \34543 );
and \U$34168 ( \34545 , \2224 , RIae78ad0_124);
and \U$34169 ( \34546 , RIae78d28_129, \2222 );
nor \U$34170 ( \34547 , \34545 , \34546 );
and \U$34171 ( \34548 , \34547 , \2060 );
not \U$34172 ( \34549 , \34547 );
and \U$34173 ( \34550 , \34549 , \2061 );
nor \U$34174 ( \34551 , \34548 , \34550 );
not \U$34175 ( \34552 , \34551 );
and \U$34176 ( \34553 , \34544 , \34552 );
and \U$34177 ( \34554 , \34551 , \34543 );
nand \U$34178 ( \34555 , RIae78e18_131, \2607 );
and \U$34179 ( \34556 , \34555 , \2397 );
not \U$34180 ( \34557 , \34555 );
and \U$34181 ( \34558 , \34557 , \2611 );
nor \U$34182 ( \34559 , \34556 , \34558 );
nor \U$34183 ( \34560 , \34554 , \34559 );
nor \U$34184 ( \34561 , \34553 , \34560 );
xor \U$34185 ( \34562 , \34536 , \34561 );
and \U$34186 ( \34563 , \558 , RIae75470_8);
and \U$34187 ( \34564 , RIae76460_42, \556 );
nor \U$34188 ( \34565 , \34563 , \34564 );
and \U$34189 ( \34566 , \34565 , \562 );
not \U$34190 ( \34567 , \34565 );
and \U$34191 ( \34568 , \34567 , \504 );
nor \U$34192 ( \34569 , \34566 , \34568 );
not \U$34193 ( \34570 , \34569 );
and \U$34194 ( \34571 , \672 , RIae76550_44);
and \U$34195 ( \34572 , RIae76730_48, \670 );
nor \U$34196 ( \34573 , \34571 , \34572 );
and \U$34197 ( \34574 , \34573 , \587 );
not \U$34198 ( \34575 , \34573 );
and \U$34199 ( \34576 , \34575 , \588 );
nor \U$34200 ( \34577 , \34574 , \34576 );
not \U$34201 ( \34578 , \34577 );
and \U$34202 ( \34579 , \34570 , \34578 );
and \U$34203 ( \34580 , \34577 , \34569 );
and \U$34204 ( \34581 , \883 , RIae76640_46);
and \U$34205 ( \34582 , RIae76190_36, \881 );
nor \U$34206 ( \34583 , \34581 , \34582 );
not \U$34207 ( \34584 , \34583 );
not \U$34208 ( \34585 , \789 );
and \U$34209 ( \34586 , \34584 , \34585 );
and \U$34210 ( \34587 , \34583 , \789 );
nor \U$34211 ( \34588 , \34586 , \34587 );
nor \U$34212 ( \34589 , \34580 , \34588 );
nor \U$34213 ( \34590 , \34579 , \34589 );
and \U$34214 ( \34591 , \34562 , \34590 );
and \U$34215 ( \34592 , \34536 , \34561 );
or \U$34216 ( \34593 , \34591 , \34592 );
nand \U$34217 ( \34594 , RIae75650_12, RIae78b48_125);
not \U$34218 ( \34595 , \34594 );
nand \U$34219 ( \34596 , RIae75560_10, RIae78b48_125);
not \U$34220 ( \34597 , \34596 );
and \U$34221 ( \34598 , \34595 , \34597 );
and \U$34222 ( \34599 , \34594 , \34596 );
not \U$34223 ( \34600 , \400 );
and \U$34224 ( \34601 , \436 , RIae75740_14);
and \U$34225 ( \34602 , RIae75290_4, \434 );
nor \U$34226 ( \34603 , \34601 , \34602 );
not \U$34227 ( \34604 , \34603 );
or \U$34228 ( \34605 , \34600 , \34604 );
or \U$34229 ( \34606 , \34603 , \402 );
nand \U$34230 ( \34607 , \34605 , \34606 );
not \U$34231 ( \34608 , \388 );
and \U$34232 ( \34609 , \384 , RIae75560_10);
and \U$34233 ( \34610 , RIae75830_16, \382 );
nor \U$34234 ( \34611 , \34609 , \34610 );
not \U$34235 ( \34612 , \34611 );
or \U$34236 ( \34613 , \34608 , \34612 );
or \U$34237 ( \34614 , \34611 , \388 );
nand \U$34238 ( \34615 , \34613 , \34614 );
xor \U$34239 ( \34616 , \34607 , \34615 );
not \U$34240 ( \34617 , \469 );
and \U$34241 ( \34618 , \514 , RIae751a0_2);
and \U$34242 ( \34619 , RIae75380_6, \512 );
nor \U$34243 ( \34620 , \34618 , \34619 );
not \U$34244 ( \34621 , \34620 );
or \U$34245 ( \34622 , \34617 , \34621 );
or \U$34246 ( \34623 , \34620 , \469 );
nand \U$34247 ( \34624 , \34622 , \34623 );
and \U$34248 ( \34625 , \34616 , \34624 );
and \U$34249 ( \34626 , \34607 , \34615 );
or \U$34250 ( \34627 , \34625 , \34626 );
not \U$34251 ( \34628 , \34627 );
nor \U$34252 ( \34629 , \34599 , \34628 );
nor \U$34253 ( \34630 , \34598 , \34629 );
xor \U$34254 ( \34631 , \34593 , \34630 );
not \U$34255 ( \34632 , \34366 );
xor \U$34256 ( \34633 , \34375 , \34386 );
not \U$34257 ( \34634 , \34633 );
or \U$34258 ( \34635 , \34632 , \34634 );
or \U$34259 ( \34636 , \34633 , \34366 );
nand \U$34260 ( \34637 , \34635 , \34636 );
xor \U$34261 ( \34638 , \34402 , \34409 );
xor \U$34262 ( \34639 , \34638 , \34417 );
xor \U$34263 ( \34640 , \34637 , \34639 );
xor \U$34264 ( \34641 , \34447 , \34454 );
xor \U$34265 ( \34642 , \34641 , \34462 );
and \U$34266 ( \34643 , \34640 , \34642 );
and \U$34267 ( \34644 , \34637 , \34639 );
nor \U$34268 ( \34645 , \34643 , \34644 );
and \U$34269 ( \34646 , \34631 , \34645 );
and \U$34270 ( \34647 , \34593 , \34630 );
or \U$34271 ( \34648 , \34646 , \34647 );
not \U$34272 ( \34649 , \34648 );
and \U$34273 ( \34650 , \34509 , \34649 );
and \U$34274 ( \34651 , \34508 , \34648 );
xor \U$34275 ( \34652 , \34420 , \34438 );
xor \U$34276 ( \34653 , \34652 , \34465 );
or \U$34277 ( \34654 , \34390 , \34388 );
nand \U$34278 ( \34655 , \34654 , \34391 );
xor \U$34279 ( \34656 , \34653 , \34655 );
xor \U$34280 ( \34657 , \34342 , \34348 );
xor \U$34281 ( \34658 , \34657 , \34355 );
and \U$34282 ( \34659 , \34656 , \34658 );
and \U$34283 ( \34660 , \34653 , \34655 );
or \U$34284 ( \34661 , \34659 , \34660 );
not \U$34285 ( \34662 , \34661 );
nor \U$34286 ( \34663 , \34651 , \34662 );
nor \U$34287 ( \34664 , \34650 , \34663 );
xor \U$34288 ( \34665 , \34218 , \34231 );
xor \U$34289 ( \34666 , \34665 , \34269 );
xor \U$34290 ( \34667 , \34664 , \34666 );
xor \U$34291 ( \34668 , \34340 , \34470 );
xor \U$34292 ( \34669 , \34668 , \34477 );
and \U$34293 ( \34670 , \34667 , \34669 );
and \U$34294 ( \34671 , \34664 , \34666 );
or \U$34295 ( \34672 , \34670 , \34671 );
nor \U$34296 ( \34673 , \34504 , \34672 );
and \U$34297 ( \34674 , \34497 , \34673 );
xor \U$34298 ( \34675 , \34673 , \34497 );
and \U$34299 ( \34676 , \514 , RIae75290_4);
and \U$34300 ( \34677 , RIae751a0_2, \512 );
nor \U$34301 ( \34678 , \34676 , \34677 );
not \U$34302 ( \34679 , \34678 );
not \U$34303 ( \34680 , \469 );
and \U$34304 ( \34681 , \34679 , \34680 );
and \U$34305 ( \34682 , \34678 , \471 );
nor \U$34306 ( \34683 , \34681 , \34682 );
and \U$34307 ( \34684 , \558 , RIae75380_6);
and \U$34308 ( \34685 , RIae75470_8, \556 );
nor \U$34309 ( \34686 , \34684 , \34685 );
and \U$34310 ( \34687 , \34686 , \562 );
not \U$34311 ( \34688 , \34686 );
and \U$34312 ( \34689 , \34688 , \504 );
nor \U$34313 ( \34690 , \34687 , \34689 );
xor \U$34314 ( \34691 , \34683 , \34690 );
and \U$34315 ( \34692 , \436 , RIae75830_16);
and \U$34316 ( \34693 , RIae75740_14, \434 );
nor \U$34317 ( \34694 , \34692 , \34693 );
not \U$34318 ( \34695 , \34694 );
not \U$34319 ( \34696 , \400 );
and \U$34320 ( \34697 , \34695 , \34696 );
and \U$34321 ( \34698 , \34694 , \400 );
nor \U$34322 ( \34699 , \34697 , \34698 );
and \U$34323 ( \34700 , \34691 , \34699 );
and \U$34324 ( \34701 , \34683 , \34690 );
nor \U$34325 ( \34702 , \34700 , \34701 );
xor \U$34326 ( \34703 , \34702 , \34594 );
xor \U$34327 ( \34704 , \34607 , \34615 );
xor \U$34328 ( \34705 , \34704 , \34624 );
and \U$34329 ( \34706 , \34703 , \34705 );
and \U$34330 ( \34707 , \34702 , \34594 );
or \U$34331 ( \34708 , \34706 , \34707 );
and \U$34332 ( \34709 , \883 , RIae76730_48);
and \U$34333 ( \34710 , RIae76640_46, \881 );
nor \U$34334 ( \34711 , \34709 , \34710 );
not \U$34335 ( \34712 , \34711 );
not \U$34336 ( \34713 , \787 );
and \U$34337 ( \34714 , \34712 , \34713 );
and \U$34338 ( \34715 , \34711 , \787 );
nor \U$34339 ( \34716 , \34714 , \34715 );
and \U$34340 ( \34717 , \1138 , RIae76190_36);
and \U$34341 ( \34718 , RIae760a0_34, \1136 );
nor \U$34342 ( \34719 , \34717 , \34718 );
and \U$34343 ( \34720 , \34719 , \1142 );
not \U$34344 ( \34721 , \34719 );
and \U$34345 ( \34722 , \34721 , \1012 );
nor \U$34346 ( \34723 , \34720 , \34722 );
xor \U$34347 ( \34724 , \34716 , \34723 );
and \U$34348 ( \34725 , \672 , RIae76460_42);
and \U$34349 ( \34726 , RIae76550_44, \670 );
nor \U$34350 ( \34727 , \34725 , \34726 );
and \U$34351 ( \34728 , \34727 , \587 );
not \U$34352 ( \34729 , \34727 );
and \U$34353 ( \34730 , \34729 , \588 );
nor \U$34354 ( \34731 , \34728 , \34730 );
and \U$34355 ( \34732 , \34724 , \34731 );
and \U$34356 ( \34733 , \34716 , \34723 );
nor \U$34357 ( \34734 , \34732 , \34733 );
and \U$34358 ( \34735 , \2224 , RIae76be0_58);
and \U$34359 ( \34736 , RIae78ad0_124, \2222 );
nor \U$34360 ( \34737 , \34735 , \34736 );
and \U$34361 ( \34738 , \34737 , \2060 );
not \U$34362 ( \34739 , \34737 );
and \U$34363 ( \34740 , \34739 , \2061 );
nor \U$34364 ( \34741 , \34738 , \34740 );
or \U$34365 ( \34742 , \34741 , \3089 );
not \U$34366 ( \34743 , \2789 );
not \U$34367 ( \34744 , \34741 );
or \U$34368 ( \34745 , \34743 , \34744 );
and \U$34369 ( \34746 , \2607 , RIae78d28_129);
and \U$34370 ( \34747 , RIae78e18_131, \2605 );
nor \U$34371 ( \34748 , \34746 , \34747 );
and \U$34372 ( \34749 , \34748 , \2611 );
not \U$34373 ( \34750 , \34748 );
and \U$34374 ( \34751 , \34750 , \2397 );
nor \U$34375 ( \34752 , \34749 , \34751 );
nand \U$34376 ( \34753 , \34745 , \34752 );
nand \U$34377 ( \34754 , \34742 , \34753 );
xor \U$34378 ( \34755 , \34734 , \34754 );
and \U$34379 ( \34756 , \1593 , RIae76af0_56);
and \U$34380 ( \34757 , RIae76a00_54, \1591 );
nor \U$34381 ( \34758 , \34756 , \34757 );
and \U$34382 ( \34759 , \34758 , \1488 );
not \U$34383 ( \34760 , \34758 );
and \U$34384 ( \34761 , \34760 , \1498 );
nor \U$34385 ( \34762 , \34759 , \34761 );
and \U$34386 ( \34763 , \1939 , RIae76820_50);
and \U$34387 ( \34764 , RIae76910_52, \1937 );
nor \U$34388 ( \34765 , \34763 , \34764 );
and \U$34389 ( \34766 , \34765 , \1734 );
not \U$34390 ( \34767 , \34765 );
and \U$34391 ( \34768 , \34767 , \1735 );
nor \U$34392 ( \34769 , \34766 , \34768 );
xor \U$34393 ( \34770 , \34762 , \34769 );
and \U$34394 ( \34771 , \1376 , RIae76370_40);
and \U$34395 ( \34772 , RIae76280_38, \1374 );
nor \U$34396 ( \34773 , \34771 , \34772 );
and \U$34397 ( \34774 , \34773 , \1261 );
not \U$34398 ( \34775 , \34773 );
and \U$34399 ( \34776 , \34775 , \1380 );
nor \U$34400 ( \34777 , \34774 , \34776 );
and \U$34401 ( \34778 , \34770 , \34777 );
and \U$34402 ( \34779 , \34762 , \34769 );
nor \U$34403 ( \34780 , \34778 , \34779 );
and \U$34404 ( \34781 , \34755 , \34780 );
and \U$34405 ( \34782 , \34734 , \34754 );
or \U$34406 ( \34783 , \34781 , \34782 );
xor \U$34407 ( \34784 , \34708 , \34783 );
not \U$34408 ( \34785 , \34516 );
xor \U$34409 ( \34786 , \34534 , \34524 );
not \U$34410 ( \34787 , \34786 );
or \U$34411 ( \34788 , \34785 , \34787 );
or \U$34412 ( \34789 , \34786 , \34516 );
nand \U$34413 ( \34790 , \34788 , \34789 );
not \U$34414 ( \34791 , \34543 );
xor \U$34415 ( \34792 , \34559 , \34551 );
not \U$34416 ( \34793 , \34792 );
or \U$34417 ( \34794 , \34791 , \34793 );
or \U$34418 ( \34795 , \34792 , \34543 );
nand \U$34419 ( \34796 , \34794 , \34795 );
xor \U$34420 ( \34797 , \34790 , \34796 );
not \U$34421 ( \34798 , \34569 );
xor \U$34422 ( \34799 , \34577 , \34588 );
not \U$34423 ( \34800 , \34799 );
or \U$34424 ( \34801 , \34798 , \34800 );
or \U$34425 ( \34802 , \34799 , \34569 );
nand \U$34426 ( \34803 , \34801 , \34802 );
and \U$34427 ( \34804 , \34797 , \34803 );
and \U$34428 ( \34805 , \34790 , \34796 );
or \U$34429 ( \34806 , \34804 , \34805 );
and \U$34430 ( \34807 , \34784 , \34806 );
and \U$34431 ( \34808 , \34708 , \34783 );
or \U$34432 ( \34809 , \34807 , \34808 );
not \U$34433 ( \34810 , \34596 );
not \U$34434 ( \34811 , \34594 );
not \U$34435 ( \34812 , \34627 );
or \U$34436 ( \34813 , \34811 , \34812 );
or \U$34437 ( \34814 , \34627 , \34594 );
nand \U$34438 ( \34815 , \34813 , \34814 );
not \U$34439 ( \34816 , \34815 );
or \U$34440 ( \34817 , \34810 , \34816 );
or \U$34441 ( \34818 , \34815 , \34596 );
nand \U$34442 ( \34819 , \34817 , \34818 );
xor \U$34443 ( \34820 , \34427 , \2611 );
xor \U$34444 ( \34821 , \34820 , \34435 );
xor \U$34445 ( \34822 , \34819 , \34821 );
xor \U$34446 ( \34823 , \34637 , \34639 );
xor \U$34447 ( \34824 , \34823 , \34642 );
and \U$34448 ( \34825 , \34822 , \34824 );
and \U$34449 ( \34826 , \34819 , \34821 );
or \U$34450 ( \34827 , \34825 , \34826 );
xor \U$34451 ( \34828 , \34809 , \34827 );
xor \U$34452 ( \34829 , \34653 , \34655 );
xor \U$34453 ( \34830 , \34829 , \34658 );
xor \U$34454 ( \34831 , \34828 , \34830 );
xor \U$34455 ( \34832 , \34593 , \34630 );
xor \U$34456 ( \34833 , \34832 , \34645 );
not \U$34457 ( \34834 , \34833 );
xor \U$34458 ( \34835 , \34819 , \34821 );
xor \U$34459 ( \34836 , \34835 , \34824 );
xor \U$34460 ( \34837 , \34708 , \34783 );
xor \U$34461 ( \34838 , \34837 , \34806 );
and \U$34462 ( \34839 , \34836 , \34838 );
not \U$34463 ( \34840 , \34839 );
and \U$34464 ( \34841 , \2224 , RIae76910_52);
and \U$34465 ( \34842 , RIae76be0_58, \2222 );
nor \U$34466 ( \34843 , \34841 , \34842 );
and \U$34467 ( \34844 , \34843 , \2060 );
not \U$34468 ( \34845 , \34843 );
and \U$34469 ( \34846 , \34845 , \2061 );
nor \U$34470 ( \34847 , \34844 , \34846 );
not \U$34471 ( \34848 , \34847 );
and \U$34472 ( \34849 , \2607 , RIae78ad0_124);
and \U$34473 ( \34850 , RIae78d28_129, \2605 );
nor \U$34474 ( \34851 , \34849 , \34850 );
and \U$34475 ( \34852 , \34851 , \2397 );
not \U$34476 ( \34853 , \34851 );
and \U$34477 ( \34854 , \34853 , \2611 );
nor \U$34478 ( \34855 , \34852 , \34854 );
not \U$34479 ( \34856 , \34855 );
and \U$34480 ( \34857 , \34848 , \34856 );
and \U$34481 ( \34858 , \34855 , \34847 );
nand \U$34482 ( \34859 , RIae78e18_131, \2783 );
not \U$34483 ( \34860 , \34859 );
not \U$34484 ( \34861 , \3089 );
and \U$34485 ( \34862 , \34860 , \34861 );
and \U$34486 ( \34863 , \34859 , \2789 );
nor \U$34487 ( \34864 , \34862 , \34863 );
nor \U$34488 ( \34865 , \34858 , \34864 );
nor \U$34489 ( \34866 , \34857 , \34865 );
and \U$34490 ( \34867 , \672 , RIae75470_8);
and \U$34491 ( \34868 , RIae76460_42, \670 );
nor \U$34492 ( \34869 , \34867 , \34868 );
and \U$34493 ( \34870 , \34869 , \587 );
not \U$34494 ( \34871 , \34869 );
and \U$34495 ( \34872 , \34871 , \588 );
nor \U$34496 ( \34873 , \34870 , \34872 );
not \U$34497 ( \34874 , \34873 );
and \U$34498 ( \34875 , \1138 , RIae76640_46);
and \U$34499 ( \34876 , RIae76190_36, \1136 );
nor \U$34500 ( \34877 , \34875 , \34876 );
and \U$34501 ( \34878 , \34877 , \1142 );
not \U$34502 ( \34879 , \34877 );
and \U$34503 ( \34880 , \34879 , \1012 );
nor \U$34504 ( \34881 , \34878 , \34880 );
not \U$34505 ( \34882 , \34881 );
and \U$34506 ( \34883 , \34874 , \34882 );
and \U$34507 ( \34884 , \34881 , \34873 );
and \U$34508 ( \34885 , \883 , RIae76550_44);
and \U$34509 ( \34886 , RIae76730_48, \881 );
nor \U$34510 ( \34887 , \34885 , \34886 );
not \U$34511 ( \34888 , \34887 );
not \U$34512 ( \34889 , \787 );
and \U$34513 ( \34890 , \34888 , \34889 );
and \U$34514 ( \34891 , \34887 , \789 );
nor \U$34515 ( \34892 , \34890 , \34891 );
nor \U$34516 ( \34893 , \34884 , \34892 );
nor \U$34517 ( \34894 , \34883 , \34893 );
or \U$34518 ( \34895 , \34866 , \34894 );
not \U$34519 ( \34896 , \34866 );
not \U$34520 ( \34897 , \34894 );
or \U$34521 ( \34898 , \34896 , \34897 );
and \U$34522 ( \34899 , \1939 , RIae76a00_54);
and \U$34523 ( \34900 , RIae76820_50, \1937 );
nor \U$34524 ( \34901 , \34899 , \34900 );
and \U$34525 ( \34902 , \34901 , \1735 );
not \U$34526 ( \34903 , \34901 );
and \U$34527 ( \34904 , \34903 , \1734 );
nor \U$34528 ( \34905 , \34902 , \34904 );
and \U$34529 ( \34906 , \1376 , RIae760a0_34);
and \U$34530 ( \34907 , RIae76370_40, \1374 );
nor \U$34531 ( \34908 , \34906 , \34907 );
and \U$34532 ( \34909 , \34908 , \1380 );
not \U$34533 ( \34910 , \34908 );
and \U$34534 ( \34911 , \34910 , \1261 );
nor \U$34535 ( \34912 , \34909 , \34911 );
xor \U$34536 ( \34913 , \34905 , \34912 );
and \U$34537 ( \34914 , \1593 , RIae76280_38);
and \U$34538 ( \34915 , RIae76af0_56, \1591 );
nor \U$34539 ( \34916 , \34914 , \34915 );
and \U$34540 ( \34917 , \34916 , \1498 );
not \U$34541 ( \34918 , \34916 );
and \U$34542 ( \34919 , \34918 , \1488 );
nor \U$34543 ( \34920 , \34917 , \34919 );
and \U$34544 ( \34921 , \34913 , \34920 );
and \U$34545 ( \34922 , \34905 , \34912 );
or \U$34546 ( \34923 , \34921 , \34922 );
nand \U$34547 ( \34924 , \34898 , \34923 );
nand \U$34548 ( \34925 , \34895 , \34924 );
nand \U$34549 ( \34926 , RIae75ce0_26, RIae78b48_125);
and \U$34550 ( \34927 , \384 , RIae75dd0_28);
and \U$34551 ( \34928 , RIae75650_12, \382 );
nor \U$34552 ( \34929 , \34927 , \34928 );
not \U$34553 ( \34930 , \34929 );
not \U$34554 ( \34931 , \388 );
and \U$34555 ( \34932 , \34930 , \34931 );
and \U$34556 ( \34933 , \34929 , \388 );
nor \U$34557 ( \34934 , \34932 , \34933 );
nand \U$34558 ( \34935 , \34926 , \34934 );
not \U$34559 ( \34936 , \392 );
and \U$34560 ( \34937 , \384 , RIae75650_12);
and \U$34561 ( \34938 , RIae75560_10, \382 );
nor \U$34562 ( \34939 , \34937 , \34938 );
not \U$34563 ( \34940 , \34939 );
or \U$34564 ( \34941 , \34936 , \34940 );
or \U$34565 ( \34942 , \34939 , \392 );
nand \U$34566 ( \34943 , \34941 , \34942 );
xor \U$34567 ( \34944 , \34935 , \34943 );
not \U$34568 ( \34945 , \402 );
and \U$34569 ( \34946 , \436 , RIae75560_10);
and \U$34570 ( \34947 , RIae75830_16, \434 );
nor \U$34571 ( \34948 , \34946 , \34947 );
not \U$34572 ( \34949 , \34948 );
or \U$34573 ( \34950 , \34945 , \34949 );
or \U$34574 ( \34951 , \34948 , \402 );
nand \U$34575 ( \34952 , \34950 , \34951 );
not \U$34576 ( \34953 , \469 );
and \U$34577 ( \34954 , \514 , RIae75740_14);
and \U$34578 ( \34955 , RIae75290_4, \512 );
nor \U$34579 ( \34956 , \34954 , \34955 );
not \U$34580 ( \34957 , \34956 );
or \U$34581 ( \34958 , \34953 , \34957 );
or \U$34582 ( \34959 , \34956 , \469 );
nand \U$34583 ( \34960 , \34958 , \34959 );
xor \U$34584 ( \34961 , \34952 , \34960 );
and \U$34585 ( \34962 , \558 , RIae751a0_2);
and \U$34586 ( \34963 , RIae75380_6, \556 );
nor \U$34587 ( \34964 , \34962 , \34963 );
and \U$34588 ( \34965 , \34964 , \504 );
not \U$34589 ( \34966 , \34964 );
and \U$34590 ( \34967 , \34966 , \562 );
nor \U$34591 ( \34968 , \34965 , \34967 );
and \U$34592 ( \34969 , \34961 , \34968 );
and \U$34593 ( \34970 , \34952 , \34960 );
or \U$34594 ( \34971 , \34969 , \34970 );
and \U$34595 ( \34972 , \34944 , \34971 );
and \U$34596 ( \34973 , \34935 , \34943 );
or \U$34597 ( \34974 , \34972 , \34973 );
and \U$34598 ( \34975 , \34925 , \34974 );
not \U$34599 ( \34976 , \34925 );
not \U$34600 ( \34977 , \34974 );
and \U$34601 ( \34978 , \34976 , \34977 );
xor \U$34602 ( \34979 , \34716 , \34723 );
xor \U$34603 ( \34980 , \34979 , \34731 );
nand \U$34604 ( \34981 , RIae75dd0_28, RIae78b48_125);
xor \U$34605 ( \34982 , \34980 , \34981 );
xor \U$34606 ( \34983 , \34683 , \34690 );
xor \U$34607 ( \34984 , \34983 , \34699 );
and \U$34608 ( \34985 , \34982 , \34984 );
and \U$34609 ( \34986 , \34980 , \34981 );
or \U$34610 ( \34987 , \34985 , \34986 );
nor \U$34611 ( \34988 , \34978 , \34987 );
nor \U$34612 ( \34989 , \34975 , \34988 );
not \U$34613 ( \34990 , \34989 );
xor \U$34614 ( \34991 , \34536 , \34561 );
xor \U$34615 ( \34992 , \34991 , \34590 );
not \U$34616 ( \34993 , \34992 );
and \U$34617 ( \34994 , \34990 , \34993 );
and \U$34618 ( \34995 , \34989 , \34992 );
xor \U$34619 ( \34996 , \34702 , \34594 );
xor \U$34620 ( \34997 , \34996 , \34705 );
xor \U$34621 ( \34998 , \34734 , \34754 );
xor \U$34622 ( \34999 , \34998 , \34780 );
xor \U$34623 ( \35000 , \34997 , \34999 );
xor \U$34624 ( \35001 , \34790 , \34796 );
xor \U$34625 ( \35002 , \35001 , \34803 );
and \U$34626 ( \35003 , \35000 , \35002 );
and \U$34627 ( \35004 , \34997 , \34999 );
nor \U$34628 ( \35005 , \35003 , \35004 );
nor \U$34629 ( \35006 , \34995 , \35005 );
nor \U$34630 ( \35007 , \34994 , \35006 );
not \U$34631 ( \35008 , \35007 );
or \U$34632 ( \35009 , \34840 , \35008 );
or \U$34633 ( \35010 , \35007 , \34839 );
nand \U$34634 ( \35011 , \35009 , \35010 );
not \U$34635 ( \35012 , \35011 );
or \U$34636 ( \35013 , \34834 , \35012 );
or \U$34637 ( \35014 , \35011 , \34833 );
nand \U$34638 ( \35015 , \35013 , \35014 );
xor \U$34639 ( \35016 , \34831 , \35015 );
and \U$34640 ( \35017 , \436 , RIae75650_12);
and \U$34641 ( \35018 , RIae75560_10, \434 );
nor \U$34642 ( \35019 , \35017 , \35018 );
not \U$34643 ( \35020 , \35019 );
not \U$34644 ( \35021 , \402 );
and \U$34645 ( \35022 , \35020 , \35021 );
and \U$34646 ( \35023 , \35019 , \402 );
nor \U$34647 ( \35024 , \35022 , \35023 );
nand \U$34648 ( \35025 , RIae75ec0_30, RIae78b48_125);
or \U$34649 ( \35026 , \35024 , \35025 );
not \U$34650 ( \35027 , \35025 );
not \U$34651 ( \35028 , \35024 );
or \U$34652 ( \35029 , \35027 , \35028 );
not \U$34653 ( \35030 , \388 );
and \U$34654 ( \35031 , \384 , RIae75ce0_26);
and \U$34655 ( \35032 , RIae75dd0_28, \382 );
nor \U$34656 ( \35033 , \35031 , \35032 );
not \U$34657 ( \35034 , \35033 );
or \U$34658 ( \35035 , \35030 , \35034 );
or \U$34659 ( \35036 , \35033 , \392 );
nand \U$34660 ( \35037 , \35035 , \35036 );
nand \U$34661 ( \35038 , \35029 , \35037 );
nand \U$34662 ( \35039 , \35026 , \35038 );
or \U$34663 ( \35040 , \34934 , \34926 );
nand \U$34664 ( \35041 , \35040 , \34935 );
xor \U$34665 ( \35042 , \35039 , \35041 );
and \U$34666 ( \35043 , \558 , RIae75290_4);
and \U$34667 ( \35044 , RIae751a0_2, \556 );
nor \U$34668 ( \35045 , \35043 , \35044 );
and \U$34669 ( \35046 , \35045 , \562 );
not \U$34670 ( \35047 , \35045 );
and \U$34671 ( \35048 , \35047 , \504 );
nor \U$34672 ( \35049 , \35046 , \35048 );
and \U$34673 ( \35050 , \672 , RIae75380_6);
and \U$34674 ( \35051 , RIae75470_8, \670 );
nor \U$34675 ( \35052 , \35050 , \35051 );
and \U$34676 ( \35053 , \35052 , \587 );
not \U$34677 ( \35054 , \35052 );
and \U$34678 ( \35055 , \35054 , \588 );
nor \U$34679 ( \35056 , \35053 , \35055 );
xor \U$34680 ( \35057 , \35049 , \35056 );
and \U$34681 ( \35058 , \514 , RIae75830_16);
and \U$34682 ( \35059 , RIae75740_14, \512 );
nor \U$34683 ( \35060 , \35058 , \35059 );
not \U$34684 ( \35061 , \35060 );
not \U$34685 ( \35062 , \469 );
and \U$34686 ( \35063 , \35061 , \35062 );
and \U$34687 ( \35064 , \35060 , \469 );
nor \U$34688 ( \35065 , \35063 , \35064 );
and \U$34689 ( \35066 , \35057 , \35065 );
and \U$34690 ( \35067 , \35049 , \35056 );
nor \U$34691 ( \35068 , \35066 , \35067 );
and \U$34692 ( \35069 , \35042 , \35068 );
and \U$34693 ( \35070 , \35039 , \35041 );
or \U$34694 ( \35071 , \35069 , \35070 );
and \U$34695 ( \35072 , \2783 , RIae78d28_129);
and \U$34696 ( \35073 , RIae78e18_131, \2781 );
nor \U$34697 ( \35074 , \35072 , \35073 );
not \U$34698 ( \35075 , \35074 );
not \U$34699 ( \35076 , \3089 );
and \U$34700 ( \35077 , \35075 , \35076 );
and \U$34701 ( \35078 , \35074 , \2789 );
nor \U$34702 ( \35079 , \35077 , \35078 );
xor \U$34703 ( \35080 , \35079 , \3218 );
and \U$34704 ( \35081 , \2607 , RIae76be0_58);
and \U$34705 ( \35082 , RIae78ad0_124, \2605 );
nor \U$34706 ( \35083 , \35081 , \35082 );
and \U$34707 ( \35084 , \35083 , \2397 );
not \U$34708 ( \35085 , \35083 );
and \U$34709 ( \35086 , \35085 , \2611 );
nor \U$34710 ( \35087 , \35084 , \35086 );
and \U$34711 ( \35088 , \35080 , \35087 );
and \U$34712 ( \35089 , \35079 , \3218 );
or \U$34713 ( \35090 , \35088 , \35089 );
and \U$34714 ( \35091 , \1939 , RIae76af0_56);
and \U$34715 ( \35092 , RIae76a00_54, \1937 );
nor \U$34716 ( \35093 , \35091 , \35092 );
and \U$34717 ( \35094 , \35093 , \1734 );
not \U$34718 ( \35095 , \35093 );
and \U$34719 ( \35096 , \35095 , \1735 );
nor \U$34720 ( \35097 , \35094 , \35096 );
and \U$34721 ( \35098 , \1593 , RIae76370_40);
and \U$34722 ( \35099 , RIae76280_38, \1591 );
nor \U$34723 ( \35100 , \35098 , \35099 );
and \U$34724 ( \35101 , \35100 , \1488 );
not \U$34725 ( \35102 , \35100 );
and \U$34726 ( \35103 , \35102 , \1498 );
nor \U$34727 ( \35104 , \35101 , \35103 );
xor \U$34728 ( \35105 , \35097 , \35104 );
and \U$34729 ( \35106 , \2224 , RIae76820_50);
and \U$34730 ( \35107 , RIae76910_52, \2222 );
nor \U$34731 ( \35108 , \35106 , \35107 );
and \U$34732 ( \35109 , \35108 , \2060 );
not \U$34733 ( \35110 , \35108 );
and \U$34734 ( \35111 , \35110 , \2061 );
nor \U$34735 ( \35112 , \35109 , \35111 );
and \U$34736 ( \35113 , \35105 , \35112 );
and \U$34737 ( \35114 , \35097 , \35104 );
or \U$34738 ( \35115 , \35113 , \35114 );
xor \U$34739 ( \35116 , \35090 , \35115 );
and \U$34740 ( \35117 , \1138 , RIae76730_48);
and \U$34741 ( \35118 , RIae76640_46, \1136 );
nor \U$34742 ( \35119 , \35117 , \35118 );
and \U$34743 ( \35120 , \35119 , \1142 );
not \U$34744 ( \35121 , \35119 );
and \U$34745 ( \35122 , \35121 , \1012 );
nor \U$34746 ( \35123 , \35120 , \35122 );
and \U$34747 ( \35124 , \883 , RIae76460_42);
and \U$34748 ( \35125 , RIae76550_44, \881 );
nor \U$34749 ( \35126 , \35124 , \35125 );
not \U$34750 ( \35127 , \35126 );
not \U$34751 ( \35128 , \789 );
and \U$34752 ( \35129 , \35127 , \35128 );
and \U$34753 ( \35130 , \35126 , \787 );
nor \U$34754 ( \35131 , \35129 , \35130 );
xor \U$34755 ( \35132 , \35123 , \35131 );
and \U$34756 ( \35133 , \1376 , RIae76190_36);
and \U$34757 ( \35134 , RIae760a0_34, \1374 );
nor \U$34758 ( \35135 , \35133 , \35134 );
and \U$34759 ( \35136 , \35135 , \1261 );
not \U$34760 ( \35137 , \35135 );
and \U$34761 ( \35138 , \35137 , \1380 );
nor \U$34762 ( \35139 , \35136 , \35138 );
and \U$34763 ( \35140 , \35132 , \35139 );
and \U$34764 ( \35141 , \35123 , \35131 );
or \U$34765 ( \35142 , \35140 , \35141 );
and \U$34766 ( \35143 , \35116 , \35142 );
and \U$34767 ( \35144 , \35090 , \35115 );
nor \U$34768 ( \35145 , \35143 , \35144 );
xor \U$34769 ( \35146 , \35071 , \35145 );
not \U$34770 ( \35147 , \34873 );
xor \U$34771 ( \35148 , \34892 , \34881 );
not \U$34772 ( \35149 , \35148 );
or \U$34773 ( \35150 , \35147 , \35149 );
or \U$34774 ( \35151 , \35148 , \34873 );
nand \U$34775 ( \35152 , \35150 , \35151 );
xor \U$34776 ( \35153 , \34952 , \34960 );
xor \U$34777 ( \35154 , \35153 , \34968 );
and \U$34778 ( \35155 , \35152 , \35154 );
xor \U$34779 ( \35156 , \34905 , \34912 );
xor \U$34780 ( \35157 , \35156 , \34920 );
xor \U$34781 ( \35158 , \34952 , \34960 );
xor \U$34782 ( \35159 , \35158 , \34968 );
and \U$34783 ( \35160 , \35157 , \35159 );
and \U$34784 ( \35161 , \35152 , \35157 );
or \U$34785 ( \35162 , \35155 , \35160 , \35161 );
and \U$34786 ( \35163 , \35146 , \35162 );
and \U$34787 ( \35164 , \35071 , \35145 );
or \U$34788 ( \35165 , \35163 , \35164 );
not \U$34789 ( \35166 , \2789 );
not \U$34790 ( \35167 , \34752 );
or \U$34791 ( \35168 , \35166 , \35167 );
or \U$34792 ( \35169 , \34752 , \2789 );
nand \U$34793 ( \35170 , \35168 , \35169 );
not \U$34794 ( \35171 , \35170 );
not \U$34795 ( \35172 , \34741 );
and \U$34796 ( \35173 , \35171 , \35172 );
and \U$34797 ( \35174 , \35170 , \34741 );
nor \U$34798 ( \35175 , \35173 , \35174 );
xor \U$34799 ( \35176 , \34762 , \34769 );
xor \U$34800 ( \35177 , \35176 , \34777 );
or \U$34801 ( \35178 , \35175 , \35177 );
and \U$34802 ( \35179 , \35175 , \35177 );
xor \U$34803 ( \35180 , \34980 , \34981 );
xor \U$34804 ( \35181 , \35180 , \34984 );
nor \U$34805 ( \35182 , \35179 , \35181 );
not \U$34806 ( \35183 , \35182 );
nand \U$34807 ( \35184 , \35178 , \35183 );
xor \U$34808 ( \35185 , \35165 , \35184 );
xor \U$34809 ( \35186 , \34997 , \34999 );
xor \U$34810 ( \35187 , \35186 , \35002 );
and \U$34811 ( \35188 , \35185 , \35187 );
and \U$34812 ( \35189 , \35165 , \35184 );
or \U$34813 ( \35190 , \35188 , \35189 );
xor \U$34814 ( \35191 , \34836 , \34838 );
xor \U$34815 ( \35192 , \35190 , \35191 );
not \U$34816 ( \35193 , \34992 );
xor \U$34817 ( \35194 , \34989 , \35005 );
not \U$34818 ( \35195 , \35194 );
or \U$34819 ( \35196 , \35193 , \35195 );
or \U$34820 ( \35197 , \35194 , \34992 );
nand \U$34821 ( \35198 , \35196 , \35197 );
and \U$34822 ( \35199 , \35192 , \35198 );
and \U$34823 ( \35200 , \35190 , \35191 );
or \U$34824 ( \35201 , \35199 , \35200 );
and \U$34825 ( \35202 , \35016 , \35201 );
and \U$34826 ( \35203 , \34831 , \35015 );
nor \U$34827 ( \35204 , \35202 , \35203 );
xor \U$34828 ( \35205 , \34809 , \34827 );
and \U$34829 ( \35206 , \35205 , \34830 );
and \U$34830 ( \35207 , \34809 , \34827 );
or \U$34831 ( \35208 , \35206 , \35207 );
not \U$34832 ( \35209 , \34391 );
not \U$34833 ( \35210 , \34358 );
not \U$34834 ( \35211 , \34468 );
and \U$34835 ( \35212 , \35210 , \35211 );
and \U$34836 ( \35213 , \34358 , \34468 );
nor \U$34837 ( \35214 , \35212 , \35213 );
not \U$34838 ( \35215 , \35214 );
or \U$34839 ( \35216 , \35209 , \35215 );
or \U$34840 ( \35217 , \35214 , \34391 );
nand \U$34841 ( \35218 , \35216 , \35217 );
xor \U$34842 ( \35219 , \35208 , \35218 );
not \U$34843 ( \35220 , \34508 );
not \U$34844 ( \35221 , \34648 );
not \U$34845 ( \35222 , \34661 );
or \U$34846 ( \35223 , \35221 , \35222 );
or \U$34847 ( \35224 , \34661 , \34648 );
nand \U$34848 ( \35225 , \35223 , \35224 );
not \U$34849 ( \35226 , \35225 );
or \U$34850 ( \35227 , \35220 , \35226 );
or \U$34851 ( \35228 , \35225 , \34508 );
nand \U$34852 ( \35229 , \35227 , \35228 );
xor \U$34853 ( \35230 , \35219 , \35229 );
not \U$34854 ( \35231 , \35230 );
not \U$34855 ( \35232 , \34833 );
and \U$34856 ( \35233 , \34839 , \35232 );
not \U$34857 ( \35234 , \34839 );
not \U$34858 ( \35235 , \35232 );
and \U$34859 ( \35236 , \35234 , \35235 );
nor \U$34860 ( \35237 , \35236 , \35007 );
nor \U$34861 ( \35238 , \35233 , \35237 );
not \U$34862 ( \35239 , \35238 );
and \U$34863 ( \35240 , \35231 , \35239 );
and \U$34864 ( \35241 , \35230 , \35238 );
nor \U$34865 ( \35242 , \35240 , \35241 );
or \U$34866 ( \35243 , \35204 , \35242 );
xnor \U$34867 ( \35244 , \35242 , \35204 );
xor \U$34868 ( \35245 , \34935 , \34943 );
xor \U$34869 ( \35246 , \35245 , \34971 );
not \U$34870 ( \35247 , \35246 );
and \U$34871 ( \35248 , \1593 , RIae760a0_34);
and \U$34872 ( \35249 , RIae76370_40, \1591 );
nor \U$34873 ( \35250 , \35248 , \35249 );
and \U$34874 ( \35251 , \35250 , \1488 );
not \U$34875 ( \35252 , \35250 );
and \U$34876 ( \35253 , \35252 , \1498 );
nor \U$34877 ( \35254 , \35251 , \35253 );
and \U$34878 ( \35255 , \1939 , RIae76280_38);
and \U$34879 ( \35256 , RIae76af0_56, \1937 );
nor \U$34880 ( \35257 , \35255 , \35256 );
and \U$34881 ( \35258 , \35257 , \1734 );
not \U$34882 ( \35259 , \35257 );
and \U$34883 ( \35260 , \35259 , \1735 );
nor \U$34884 ( \35261 , \35258 , \35260 );
xor \U$34885 ( \35262 , \35254 , \35261 );
and \U$34886 ( \35263 , \2224 , RIae76a00_54);
and \U$34887 ( \35264 , RIae76820_50, \2222 );
nor \U$34888 ( \35265 , \35263 , \35264 );
and \U$34889 ( \35266 , \35265 , \2060 );
not \U$34890 ( \35267 , \35265 );
and \U$34891 ( \35268 , \35267 , \2061 );
nor \U$34892 ( \35269 , \35266 , \35268 );
and \U$34893 ( \35270 , \35262 , \35269 );
and \U$34894 ( \35271 , \35254 , \35261 );
or \U$34895 ( \35272 , \35270 , \35271 );
and \U$34896 ( \35273 , \2607 , RIae76910_52);
and \U$34897 ( \35274 , RIae76be0_58, \2605 );
nor \U$34898 ( \35275 , \35273 , \35274 );
and \U$34899 ( \35276 , \35275 , \2397 );
not \U$34900 ( \35277 , \35275 );
and \U$34901 ( \35278 , \35277 , \2611 );
nor \U$34902 ( \35279 , \35276 , \35278 );
nand \U$34903 ( \35280 , RIae78e18_131, \3214 );
not \U$34904 ( \35281 , \35280 );
not \U$34905 ( \35282 , \3218 );
and \U$34906 ( \35283 , \35281 , \35282 );
and \U$34907 ( \35284 , \35280 , \3218 );
nor \U$34908 ( \35285 , \35283 , \35284 );
xor \U$34909 ( \35286 , \35279 , \35285 );
and \U$34910 ( \35287 , \2783 , RIae78ad0_124);
and \U$34911 ( \35288 , RIae78d28_129, \2781 );
nor \U$34912 ( \35289 , \35287 , \35288 );
not \U$34913 ( \35290 , \35289 );
not \U$34914 ( \35291 , \3089 );
and \U$34915 ( \35292 , \35290 , \35291 );
and \U$34916 ( \35293 , \35289 , \3089 );
nor \U$34917 ( \35294 , \35292 , \35293 );
and \U$34918 ( \35295 , \35286 , \35294 );
and \U$34919 ( \35296 , \35279 , \35285 );
or \U$34920 ( \35297 , \35295 , \35296 );
xor \U$34921 ( \35298 , \35272 , \35297 );
and \U$34922 ( \35299 , \1376 , RIae76640_46);
and \U$34923 ( \35300 , RIae76190_36, \1374 );
nor \U$34924 ( \35301 , \35299 , \35300 );
and \U$34925 ( \35302 , \35301 , \1261 );
not \U$34926 ( \35303 , \35301 );
and \U$34927 ( \35304 , \35303 , \1380 );
nor \U$34928 ( \35305 , \35302 , \35304 );
and \U$34929 ( \35306 , \883 , RIae75470_8);
and \U$34930 ( \35307 , RIae76460_42, \881 );
nor \U$34931 ( \35308 , \35306 , \35307 );
not \U$34932 ( \35309 , \35308 );
not \U$34933 ( \35310 , \787 );
and \U$34934 ( \35311 , \35309 , \35310 );
and \U$34935 ( \35312 , \35308 , \787 );
nor \U$34936 ( \35313 , \35311 , \35312 );
xor \U$34937 ( \35314 , \35305 , \35313 );
and \U$34938 ( \35315 , \1138 , RIae76550_44);
and \U$34939 ( \35316 , RIae76730_48, \1136 );
nor \U$34940 ( \35317 , \35315 , \35316 );
and \U$34941 ( \35318 , \35317 , \1142 );
not \U$34942 ( \35319 , \35317 );
and \U$34943 ( \35320 , \35319 , \1012 );
nor \U$34944 ( \35321 , \35318 , \35320 );
and \U$34945 ( \35322 , \35314 , \35321 );
and \U$34946 ( \35323 , \35305 , \35313 );
or \U$34947 ( \35324 , \35322 , \35323 );
and \U$34948 ( \35325 , \35298 , \35324 );
and \U$34949 ( \35326 , \35272 , \35297 );
or \U$34950 ( \35327 , \35325 , \35326 );
and \U$34951 ( \35328 , \558 , RIae75740_14);
and \U$34952 ( \35329 , RIae75290_4, \556 );
nor \U$34953 ( \35330 , \35328 , \35329 );
and \U$34954 ( \35331 , \35330 , \562 );
not \U$34955 ( \35332 , \35330 );
and \U$34956 ( \35333 , \35332 , \504 );
nor \U$34957 ( \35334 , \35331 , \35333 );
and \U$34958 ( \35335 , \514 , RIae75560_10);
and \U$34959 ( \35336 , RIae75830_16, \512 );
nor \U$34960 ( \35337 , \35335 , \35336 );
not \U$34961 ( \35338 , \35337 );
not \U$34962 ( \35339 , \469 );
and \U$34963 ( \35340 , \35338 , \35339 );
and \U$34964 ( \35341 , \35337 , \469 );
nor \U$34965 ( \35342 , \35340 , \35341 );
xor \U$34966 ( \35343 , \35334 , \35342 );
and \U$34967 ( \35344 , \672 , RIae751a0_2);
and \U$34968 ( \35345 , RIae75380_6, \670 );
nor \U$34969 ( \35346 , \35344 , \35345 );
and \U$34970 ( \35347 , \35346 , \587 );
not \U$34971 ( \35348 , \35346 );
and \U$34972 ( \35349 , \35348 , \588 );
nor \U$34973 ( \35350 , \35347 , \35349 );
and \U$34974 ( \35351 , \35343 , \35350 );
and \U$34975 ( \35352 , \35334 , \35342 );
or \U$34976 ( \35353 , \35351 , \35352 );
and \U$34977 ( \35354 , \436 , RIae75dd0_28);
and \U$34978 ( \35355 , RIae75650_12, \434 );
nor \U$34979 ( \35356 , \35354 , \35355 );
not \U$34980 ( \35357 , \35356 );
not \U$34981 ( \35358 , \400 );
and \U$34982 ( \35359 , \35357 , \35358 );
and \U$34983 ( \35360 , \35356 , \400 );
nor \U$34984 ( \35361 , \35359 , \35360 );
nand \U$34985 ( \35362 , RIae75fb0_32, RIae78b48_125);
xor \U$34986 ( \35363 , \35361 , \35362 );
and \U$34987 ( \35364 , \384 , RIae75ec0_30);
and \U$34988 ( \35365 , RIae75ce0_26, \382 );
nor \U$34989 ( \35366 , \35364 , \35365 );
not \U$34990 ( \35367 , \35366 );
not \U$34991 ( \35368 , \392 );
and \U$34992 ( \35369 , \35367 , \35368 );
and \U$34993 ( \35370 , \35366 , \392 );
nor \U$34994 ( \35371 , \35369 , \35370 );
and \U$34995 ( \35372 , \35363 , \35371 );
and \U$34996 ( \35373 , \35361 , \35362 );
or \U$34997 ( \35374 , \35372 , \35373 );
xor \U$34998 ( \35375 , \35353 , \35374 );
not \U$34999 ( \35376 , \35024 );
not \U$35000 ( \35377 , \35037 );
or \U$35001 ( \35378 , \35376 , \35377 );
or \U$35002 ( \35379 , \35024 , \35037 );
nand \U$35003 ( \35380 , \35378 , \35379 );
not \U$35004 ( \35381 , \35380 );
not \U$35005 ( \35382 , \35025 );
and \U$35006 ( \35383 , \35381 , \35382 );
and \U$35007 ( \35384 , \35380 , \35025 );
nor \U$35008 ( \35385 , \35383 , \35384 );
and \U$35009 ( \35386 , \35375 , \35385 );
and \U$35010 ( \35387 , \35353 , \35374 );
or \U$35011 ( \35388 , \35386 , \35387 );
xor \U$35012 ( \35389 , \35327 , \35388 );
xor \U$35013 ( \35390 , \35049 , \35056 );
xor \U$35014 ( \35391 , \35390 , \35065 );
xor \U$35015 ( \35392 , \35123 , \35131 );
xor \U$35016 ( \35393 , \35392 , \35139 );
and \U$35017 ( \35394 , \35391 , \35393 );
xor \U$35018 ( \35395 , \35097 , \35104 );
xor \U$35019 ( \35396 , \35395 , \35112 );
xor \U$35020 ( \35397 , \35123 , \35131 );
xor \U$35021 ( \35398 , \35397 , \35139 );
and \U$35022 ( \35399 , \35396 , \35398 );
and \U$35023 ( \35400 , \35391 , \35396 );
or \U$35024 ( \35401 , \35394 , \35399 , \35400 );
and \U$35025 ( \35402 , \35389 , \35401 );
and \U$35026 ( \35403 , \35327 , \35388 );
nor \U$35027 ( \35404 , \35402 , \35403 );
not \U$35028 ( \35405 , \35404 );
or \U$35029 ( \35406 , \35247 , \35405 );
or \U$35030 ( \35407 , \35404 , \35246 );
not \U$35031 ( \35408 , \34847 );
xor \U$35032 ( \35409 , \34864 , \34855 );
not \U$35033 ( \35410 , \35409 );
or \U$35034 ( \35411 , \35408 , \35410 );
or \U$35035 ( \35412 , \35409 , \34847 );
nand \U$35036 ( \35413 , \35411 , \35412 );
xor \U$35037 ( \35414 , \35039 , \35041 );
xor \U$35038 ( \35415 , \35414 , \35068 );
and \U$35039 ( \35416 , \35413 , \35415 );
xor \U$35040 ( \35417 , \34952 , \34960 );
xor \U$35041 ( \35418 , \35417 , \34968 );
xor \U$35042 ( \35419 , \35152 , \35157 );
xor \U$35043 ( \35420 , \35418 , \35419 );
xor \U$35044 ( \35421 , \35039 , \35041 );
xor \U$35045 ( \35422 , \35421 , \35068 );
and \U$35046 ( \35423 , \35420 , \35422 );
and \U$35047 ( \35424 , \35413 , \35420 );
or \U$35048 ( \35425 , \35416 , \35423 , \35424 );
nand \U$35049 ( \35426 , \35407 , \35425 );
nand \U$35050 ( \35427 , \35406 , \35426 );
not \U$35051 ( \35428 , \34987 );
xor \U$35052 ( \35429 , \34974 , \34925 );
not \U$35053 ( \35430 , \35429 );
or \U$35054 ( \35431 , \35428 , \35430 );
or \U$35055 ( \35432 , \35429 , \34987 );
nand \U$35056 ( \35433 , \35431 , \35432 );
xor \U$35057 ( \35434 , \35427 , \35433 );
not \U$35058 ( \35435 , \35181 );
xor \U$35059 ( \35436 , \35175 , \35177 );
not \U$35060 ( \35437 , \35436 );
and \U$35061 ( \35438 , \35435 , \35437 );
and \U$35062 ( \35439 , \35181 , \35436 );
nor \U$35063 ( \35440 , \35438 , \35439 );
not \U$35064 ( \35441 , \34923 );
not \U$35065 ( \35442 , \34894 );
or \U$35066 ( \35443 , \35441 , \35442 );
or \U$35067 ( \35444 , \34894 , \34923 );
nand \U$35068 ( \35445 , \35443 , \35444 );
not \U$35069 ( \35446 , \35445 );
not \U$35070 ( \35447 , \34866 );
and \U$35071 ( \35448 , \35446 , \35447 );
and \U$35072 ( \35449 , \35445 , \34866 );
nor \U$35073 ( \35450 , \35448 , \35449 );
or \U$35074 ( \35451 , \35440 , \35450 );
not \U$35075 ( \35452 , \35450 );
not \U$35076 ( \35453 , \35440 );
or \U$35077 ( \35454 , \35452 , \35453 );
xor \U$35078 ( \35455 , \35071 , \35145 );
xor \U$35079 ( \35456 , \35455 , \35162 );
nand \U$35080 ( \35457 , \35454 , \35456 );
nand \U$35081 ( \35458 , \35451 , \35457 );
and \U$35082 ( \35459 , \35434 , \35458 );
and \U$35083 ( \35460 , \35427 , \35433 );
or \U$35084 ( \35461 , \35459 , \35460 );
not \U$35085 ( \35462 , \35461 );
xor \U$35086 ( \35463 , \35190 , \35191 );
xor \U$35087 ( \35464 , \35463 , \35198 );
not \U$35088 ( \35465 , \35464 );
or \U$35089 ( \35466 , \35462 , \35465 );
or \U$35090 ( \35467 , \35464 , \35461 );
xor \U$35091 ( \35468 , \35427 , \35433 );
xor \U$35092 ( \35469 , \35468 , \35458 );
xor \U$35093 ( \35470 , \35165 , \35184 );
xor \U$35094 ( \35471 , \35470 , \35187 );
and \U$35095 ( \35472 , \35469 , \35471 );
not \U$35096 ( \35473 , \35469 );
not \U$35097 ( \35474 , \35471 );
and \U$35098 ( \35475 , \35473 , \35474 );
xnor \U$35099 ( \35476 , \35404 , \35425 );
not \U$35100 ( \35477 , \35476 );
not \U$35101 ( \35478 , \35246 );
and \U$35102 ( \35479 , \35477 , \35478 );
and \U$35103 ( \35480 , \35476 , \35246 );
nor \U$35104 ( \35481 , \35479 , \35480 );
xor \U$35105 ( \35482 , \35079 , \3218 );
xor \U$35106 ( \35483 , \35482 , \35087 );
xor \U$35107 ( \35484 , \35353 , \35374 );
xor \U$35108 ( \35485 , \35484 , \35385 );
xor \U$35109 ( \35486 , \35483 , \35485 );
xor \U$35110 ( \35487 , \35123 , \35131 );
xor \U$35111 ( \35488 , \35487 , \35139 );
xor \U$35112 ( \35489 , \35391 , \35396 );
xor \U$35113 ( \35490 , \35488 , \35489 );
and \U$35114 ( \35491 , \35486 , \35490 );
and \U$35115 ( \35492 , \35483 , \35485 );
nor \U$35116 ( \35493 , \35491 , \35492 );
xor \U$35117 ( \35494 , \35090 , \35115 );
xor \U$35118 ( \35495 , \35494 , \35142 );
not \U$35119 ( \35496 , \35495 );
and \U$35120 ( \35497 , \35493 , \35496 );
not \U$35121 ( \35498 , \35493 );
not \U$35122 ( \35499 , \35496 );
and \U$35123 ( \35500 , \35498 , \35499 );
and \U$35124 ( \35501 , \2607 , RIae76820_50);
and \U$35125 ( \35502 , RIae76910_52, \2605 );
nor \U$35126 ( \35503 , \35501 , \35502 );
and \U$35127 ( \35504 , \35503 , \2397 );
not \U$35128 ( \35505 , \35503 );
and \U$35129 ( \35506 , \35505 , \2611 );
nor \U$35130 ( \35507 , \35504 , \35506 );
and \U$35131 ( \35508 , \1939 , RIae76370_40);
and \U$35132 ( \35509 , RIae76280_38, \1937 );
nor \U$35133 ( \35510 , \35508 , \35509 );
and \U$35134 ( \35511 , \35510 , \1734 );
not \U$35135 ( \35512 , \35510 );
and \U$35136 ( \35513 , \35512 , \1735 );
nor \U$35137 ( \35514 , \35511 , \35513 );
xor \U$35138 ( \35515 , \35507 , \35514 );
and \U$35139 ( \35516 , \2224 , RIae76af0_56);
and \U$35140 ( \35517 , RIae76a00_54, \2222 );
nor \U$35141 ( \35518 , \35516 , \35517 );
and \U$35142 ( \35519 , \35518 , \2060 );
not \U$35143 ( \35520 , \35518 );
and \U$35144 ( \35521 , \35520 , \2061 );
nor \U$35145 ( \35522 , \35519 , \35521 );
and \U$35146 ( \35523 , \35515 , \35522 );
and \U$35147 ( \35524 , \35507 , \35514 );
or \U$35148 ( \35525 , \35523 , \35524 );
and \U$35149 ( \35526 , \2783 , RIae76be0_58);
and \U$35150 ( \35527 , RIae78ad0_124, \2781 );
nor \U$35151 ( \35528 , \35526 , \35527 );
not \U$35152 ( \35529 , \35528 );
not \U$35153 ( \35530 , \3089 );
and \U$35154 ( \35531 , \35529 , \35530 );
and \U$35155 ( \35532 , \35528 , \2789 );
nor \U$35156 ( \35533 , \35531 , \35532 );
xor \U$35157 ( \35534 , \35533 , \3422 );
and \U$35158 ( \35535 , \3214 , RIae78d28_129);
and \U$35159 ( \35536 , RIae78e18_131, \3212 );
nor \U$35160 ( \35537 , \35535 , \35536 );
not \U$35161 ( \35538 , \35537 );
not \U$35162 ( \35539 , \3218 );
and \U$35163 ( \35540 , \35538 , \35539 );
and \U$35164 ( \35541 , \35537 , \3218 );
nor \U$35165 ( \35542 , \35540 , \35541 );
and \U$35166 ( \35543 , \35534 , \35542 );
and \U$35167 ( \35544 , \35533 , \3422 );
or \U$35168 ( \35545 , \35543 , \35544 );
xor \U$35169 ( \35546 , \35525 , \35545 );
and \U$35170 ( \35547 , \1593 , RIae76190_36);
and \U$35171 ( \35548 , RIae760a0_34, \1591 );
nor \U$35172 ( \35549 , \35547 , \35548 );
and \U$35173 ( \35550 , \35549 , \1488 );
not \U$35174 ( \35551 , \35549 );
and \U$35175 ( \35552 , \35551 , \1498 );
nor \U$35176 ( \35553 , \35550 , \35552 );
and \U$35177 ( \35554 , \1138 , RIae76460_42);
and \U$35178 ( \35555 , RIae76550_44, \1136 );
nor \U$35179 ( \35556 , \35554 , \35555 );
and \U$35180 ( \35557 , \35556 , \1142 );
not \U$35181 ( \35558 , \35556 );
and \U$35182 ( \35559 , \35558 , \1012 );
nor \U$35183 ( \35560 , \35557 , \35559 );
xor \U$35184 ( \35561 , \35553 , \35560 );
and \U$35185 ( \35562 , \1376 , RIae76730_48);
and \U$35186 ( \35563 , RIae76640_46, \1374 );
nor \U$35187 ( \35564 , \35562 , \35563 );
and \U$35188 ( \35565 , \35564 , \1261 );
not \U$35189 ( \35566 , \35564 );
and \U$35190 ( \35567 , \35566 , \1380 );
nor \U$35191 ( \35568 , \35565 , \35567 );
and \U$35192 ( \35569 , \35561 , \35568 );
and \U$35193 ( \35570 , \35553 , \35560 );
or \U$35194 ( \35571 , \35569 , \35570 );
and \U$35195 ( \35572 , \35546 , \35571 );
and \U$35196 ( \35573 , \35525 , \35545 );
or \U$35197 ( \35574 , \35572 , \35573 );
and \U$35198 ( \35575 , \384 , RIae75fb0_32);
and \U$35199 ( \35576 , RIae75ec0_30, \382 );
nor \U$35200 ( \35577 , \35575 , \35576 );
not \U$35201 ( \35578 , \35577 );
not \U$35202 ( \35579 , \388 );
and \U$35203 ( \35580 , \35578 , \35579 );
and \U$35204 ( \35581 , \35577 , \388 );
nor \U$35205 ( \35582 , \35580 , \35581 );
and \U$35206 ( \35583 , \514 , RIae75650_12);
and \U$35207 ( \35584 , RIae75560_10, \512 );
nor \U$35208 ( \35585 , \35583 , \35584 );
not \U$35209 ( \35586 , \35585 );
not \U$35210 ( \35587 , \469 );
and \U$35211 ( \35588 , \35586 , \35587 );
and \U$35212 ( \35589 , \35585 , \471 );
nor \U$35213 ( \35590 , \35588 , \35589 );
or \U$35214 ( \35591 , \35582 , \35590 );
not \U$35215 ( \35592 , \35590 );
not \U$35216 ( \35593 , \35582 );
or \U$35217 ( \35594 , \35592 , \35593 );
not \U$35218 ( \35595 , \402 );
and \U$35219 ( \35596 , \436 , RIae75ce0_26);
and \U$35220 ( \35597 , RIae75dd0_28, \434 );
nor \U$35221 ( \35598 , \35596 , \35597 );
not \U$35222 ( \35599 , \35598 );
or \U$35223 ( \35600 , \35595 , \35599 );
or \U$35224 ( \35601 , \35598 , \402 );
nand \U$35225 ( \35602 , \35600 , \35601 );
nand \U$35226 ( \35603 , \35594 , \35602 );
nand \U$35227 ( \35604 , \35591 , \35603 );
and \U$35228 ( \35605 , \672 , RIae75290_4);
and \U$35229 ( \35606 , RIae751a0_2, \670 );
nor \U$35230 ( \35607 , \35605 , \35606 );
and \U$35231 ( \35608 , \35607 , \587 );
not \U$35232 ( \35609 , \35607 );
and \U$35233 ( \35610 , \35609 , \588 );
nor \U$35234 ( \35611 , \35608 , \35610 );
and \U$35235 ( \35612 , \883 , RIae75380_6);
and \U$35236 ( \35613 , RIae75470_8, \881 );
nor \U$35237 ( \35614 , \35612 , \35613 );
not \U$35238 ( \35615 , \35614 );
not \U$35239 ( \35616 , \787 );
and \U$35240 ( \35617 , \35615 , \35616 );
and \U$35241 ( \35618 , \35614 , \789 );
nor \U$35242 ( \35619 , \35617 , \35618 );
xor \U$35243 ( \35620 , \35611 , \35619 );
and \U$35244 ( \35621 , \558 , RIae75830_16);
and \U$35245 ( \35622 , RIae75740_14, \556 );
nor \U$35246 ( \35623 , \35621 , \35622 );
and \U$35247 ( \35624 , \35623 , \562 );
not \U$35248 ( \35625 , \35623 );
and \U$35249 ( \35626 , \35625 , \504 );
nor \U$35250 ( \35627 , \35624 , \35626 );
and \U$35251 ( \35628 , \35620 , \35627 );
and \U$35252 ( \35629 , \35611 , \35619 );
nor \U$35253 ( \35630 , \35628 , \35629 );
nor \U$35254 ( \35631 , \35604 , \35630 );
xor \U$35255 ( \35632 , \35574 , \35631 );
xor \U$35256 ( \35633 , \35334 , \35342 );
xor \U$35257 ( \35634 , \35633 , \35350 );
xor \U$35258 ( \35635 , \35361 , \35362 );
xor \U$35259 ( \35636 , \35635 , \35371 );
and \U$35260 ( \35637 , \35634 , \35636 );
xor \U$35261 ( \35638 , \35305 , \35313 );
xor \U$35262 ( \35639 , \35638 , \35321 );
xor \U$35263 ( \35640 , \35361 , \35362 );
xor \U$35264 ( \35641 , \35640 , \35371 );
and \U$35265 ( \35642 , \35639 , \35641 );
and \U$35266 ( \35643 , \35634 , \35639 );
or \U$35267 ( \35644 , \35637 , \35642 , \35643 );
and \U$35268 ( \35645 , \35632 , \35644 );
and \U$35269 ( \35646 , \35574 , \35631 );
or \U$35270 ( \35647 , \35645 , \35646 );
nor \U$35271 ( \35648 , \35500 , \35647 );
nor \U$35272 ( \35649 , \35497 , \35648 );
xor \U$35273 ( \35650 , \35481 , \35649 );
not \U$35274 ( \35651 , \35450 );
not \U$35275 ( \35652 , \35456 );
or \U$35276 ( \35653 , \35651 , \35652 );
or \U$35277 ( \35654 , \35456 , \35450 );
nand \U$35278 ( \35655 , \35653 , \35654 );
not \U$35279 ( \35656 , \35655 );
not \U$35280 ( \35657 , \35440 );
and \U$35281 ( \35658 , \35656 , \35657 );
and \U$35282 ( \35659 , \35655 , \35440 );
nor \U$35283 ( \35660 , \35658 , \35659 );
and \U$35284 ( \35661 , \35650 , \35660 );
and \U$35285 ( \35662 , \35481 , \35649 );
or \U$35286 ( \35663 , \35661 , \35662 );
nor \U$35287 ( \35664 , \35475 , \35663 );
nor \U$35288 ( \35665 , \35472 , \35664 );
not \U$35289 ( \35666 , \35665 );
nand \U$35290 ( \35667 , \35467 , \35666 );
nand \U$35291 ( \35668 , \35466 , \35667 );
xor \U$35292 ( \35669 , \34831 , \35015 );
xor \U$35293 ( \35670 , \35669 , \35201 );
and \U$35294 ( \35671 , \35668 , \35670 );
xor \U$35295 ( \35672 , \35670 , \35668 );
not \U$35296 ( \35673 , \35665 );
not \U$35297 ( \35674 , \35461 );
and \U$35298 ( \35675 , \35673 , \35674 );
and \U$35299 ( \35676 , \35665 , \35461 );
nor \U$35300 ( \35677 , \35675 , \35676 );
not \U$35301 ( \35678 , \35677 );
not \U$35302 ( \35679 , \35464 );
and \U$35303 ( \35680 , \35678 , \35679 );
and \U$35304 ( \35681 , \35677 , \35464 );
nor \U$35305 ( \35682 , \35680 , \35681 );
xor \U$35306 ( \35683 , \35481 , \35649 );
xor \U$35307 ( \35684 , \35683 , \35660 );
not \U$35308 ( \35685 , \35684 );
xor \U$35309 ( \35686 , \35327 , \35388 );
xor \U$35310 ( \35687 , \35686 , \35401 );
not \U$35311 ( \35688 , \35687 );
not \U$35312 ( \35689 , \35495 );
not \U$35313 ( \35690 , \35647 );
not \U$35314 ( \35691 , \35493 );
or \U$35315 ( \35692 , \35690 , \35691 );
or \U$35316 ( \35693 , \35493 , \35647 );
nand \U$35317 ( \35694 , \35692 , \35693 );
not \U$35318 ( \35695 , \35694 );
or \U$35319 ( \35696 , \35689 , \35695 );
or \U$35320 ( \35697 , \35694 , \35495 );
nand \U$35321 ( \35698 , \35696 , \35697 );
nand \U$35322 ( \35699 , \35688 , \35698 );
not \U$35323 ( \35700 , \35699 );
and \U$35324 ( \35701 , \35685 , \35700 );
and \U$35325 ( \35702 , \35684 , \35699 );
xor \U$35326 ( \35703 , \35272 , \35297 );
xor \U$35327 ( \35704 , \35703 , \35324 );
xor \U$35328 ( \35705 , \35574 , \35631 );
xor \U$35329 ( \35706 , \35705 , \35644 );
xor \U$35330 ( \35707 , \35704 , \35706 );
xor \U$35331 ( \35708 , \35483 , \35485 );
xor \U$35332 ( \35709 , \35708 , \35490 );
and \U$35333 ( \35710 , \35707 , \35709 );
and \U$35334 ( \35711 , \35704 , \35706 );
nor \U$35335 ( \35712 , \35710 , \35711 );
xor \U$35336 ( \35713 , \35039 , \35041 );
xor \U$35337 ( \35714 , \35713 , \35068 );
xor \U$35338 ( \35715 , \35413 , \35420 );
xor \U$35339 ( \35716 , \35714 , \35715 );
and \U$35340 ( \35717 , \35712 , \35716 );
not \U$35341 ( \35718 , \35712 );
not \U$35342 ( \35719 , \35716 );
and \U$35343 ( \35720 , \35718 , \35719 );
and \U$35344 ( \35721 , \2783 , RIae76910_52);
and \U$35345 ( \35722 , RIae76be0_58, \2781 );
nor \U$35346 ( \35723 , \35721 , \35722 );
not \U$35347 ( \35724 , \35723 );
not \U$35348 ( \35725 , \2789 );
and \U$35349 ( \35726 , \35724 , \35725 );
and \U$35350 ( \35727 , \35723 , \2789 );
nor \U$35351 ( \35728 , \35726 , \35727 );
not \U$35352 ( \35729 , \35728 );
and \U$35353 ( \35730 , \3214 , RIae78ad0_124);
and \U$35354 ( \35731 , RIae78d28_129, \3212 );
nor \U$35355 ( \35732 , \35730 , \35731 );
not \U$35356 ( \35733 , \35732 );
not \U$35357 ( \35734 , \2774 );
and \U$35358 ( \35735 , \35733 , \35734 );
and \U$35359 ( \35736 , \35732 , \3218 );
nor \U$35360 ( \35737 , \35735 , \35736 );
not \U$35361 ( \35738 , \35737 );
and \U$35362 ( \35739 , \35729 , \35738 );
and \U$35363 ( \35740 , \35737 , \35728 );
nand \U$35364 ( \35741 , RIae78e18_131, \3730 );
and \U$35365 ( \35742 , \35741 , \3422 );
not \U$35366 ( \35743 , \35741 );
and \U$35367 ( \35744 , \35743 , \3732 );
nor \U$35368 ( \35745 , \35742 , \35744 );
nor \U$35369 ( \35746 , \35740 , \35745 );
nor \U$35370 ( \35747 , \35739 , \35746 );
not \U$35371 ( \35748 , \35747 );
and \U$35372 ( \35749 , \1138 , RIae75470_8);
and \U$35373 ( \35750 , RIae76460_42, \1136 );
nor \U$35374 ( \35751 , \35749 , \35750 );
and \U$35375 ( \35752 , \35751 , \1142 );
not \U$35376 ( \35753 , \35751 );
and \U$35377 ( \35754 , \35753 , \1012 );
nor \U$35378 ( \35755 , \35752 , \35754 );
not \U$35379 ( \35756 , \35755 );
and \U$35380 ( \35757 , \1593 , RIae76640_46);
and \U$35381 ( \35758 , RIae76190_36, \1591 );
nor \U$35382 ( \35759 , \35757 , \35758 );
and \U$35383 ( \35760 , \35759 , \1488 );
not \U$35384 ( \35761 , \35759 );
and \U$35385 ( \35762 , \35761 , \1498 );
nor \U$35386 ( \35763 , \35760 , \35762 );
not \U$35387 ( \35764 , \35763 );
and \U$35388 ( \35765 , \35756 , \35764 );
and \U$35389 ( \35766 , \35763 , \35755 );
and \U$35390 ( \35767 , \1376 , RIae76550_44);
and \U$35391 ( \35768 , RIae76730_48, \1374 );
nor \U$35392 ( \35769 , \35767 , \35768 );
and \U$35393 ( \35770 , \35769 , \1261 );
not \U$35394 ( \35771 , \35769 );
and \U$35395 ( \35772 , \35771 , \1380 );
nor \U$35396 ( \35773 , \35770 , \35772 );
nor \U$35397 ( \35774 , \35766 , \35773 );
nor \U$35398 ( \35775 , \35765 , \35774 );
not \U$35399 ( \35776 , \35775 );
and \U$35400 ( \35777 , \35748 , \35776 );
and \U$35401 ( \35778 , \35747 , \35775 );
and \U$35402 ( \35779 , \1939 , RIae760a0_34);
and \U$35403 ( \35780 , RIae76370_40, \1937 );
nor \U$35404 ( \35781 , \35779 , \35780 );
and \U$35405 ( \35782 , \35781 , \1734 );
not \U$35406 ( \35783 , \35781 );
and \U$35407 ( \35784 , \35783 , \1735 );
nor \U$35408 ( \35785 , \35782 , \35784 );
not \U$35409 ( \35786 , \35785 );
and \U$35410 ( \35787 , \2224 , RIae76280_38);
and \U$35411 ( \35788 , RIae76af0_56, \2222 );
nor \U$35412 ( \35789 , \35787 , \35788 );
and \U$35413 ( \35790 , \35789 , \2060 );
not \U$35414 ( \35791 , \35789 );
and \U$35415 ( \35792 , \35791 , \2061 );
nor \U$35416 ( \35793 , \35790 , \35792 );
not \U$35417 ( \35794 , \35793 );
and \U$35418 ( \35795 , \35786 , \35794 );
and \U$35419 ( \35796 , \35793 , \35785 );
and \U$35420 ( \35797 , \2607 , RIae76a00_54);
and \U$35421 ( \35798 , RIae76820_50, \2605 );
nor \U$35422 ( \35799 , \35797 , \35798 );
and \U$35423 ( \35800 , \35799 , \2397 );
not \U$35424 ( \35801 , \35799 );
and \U$35425 ( \35802 , \35801 , \2611 );
nor \U$35426 ( \35803 , \35800 , \35802 );
nor \U$35427 ( \35804 , \35796 , \35803 );
nor \U$35428 ( \35805 , \35795 , \35804 );
nor \U$35429 ( \35806 , \35778 , \35805 );
nor \U$35430 ( \35807 , \35777 , \35806 );
not \U$35431 ( \35808 , \471 );
and \U$35432 ( \35809 , \514 , RIae75dd0_28);
and \U$35433 ( \35810 , RIae75650_12, \512 );
nor \U$35434 ( \35811 , \35809 , \35810 );
not \U$35435 ( \35812 , \35811 );
or \U$35436 ( \35813 , \35808 , \35812 );
or \U$35437 ( \35814 , \35811 , \471 );
nand \U$35438 ( \35815 , \35813 , \35814 );
not \U$35439 ( \35816 , \392 );
and \U$35440 ( \35817 , \384 , RIae75920_18);
and \U$35441 ( \35818 , RIae75fb0_32, \382 );
nor \U$35442 ( \35819 , \35817 , \35818 );
not \U$35443 ( \35820 , \35819 );
or \U$35444 ( \35821 , \35816 , \35820 );
or \U$35445 ( \35822 , \35819 , \388 );
nand \U$35446 ( \35823 , \35821 , \35822 );
xor \U$35447 ( \35824 , \35815 , \35823 );
not \U$35448 ( \35825 , \400 );
and \U$35449 ( \35826 , \436 , RIae75ec0_30);
and \U$35450 ( \35827 , RIae75ce0_26, \434 );
nor \U$35451 ( \35828 , \35826 , \35827 );
not \U$35452 ( \35829 , \35828 );
or \U$35453 ( \35830 , \35825 , \35829 );
or \U$35454 ( \35831 , \35828 , \402 );
nand \U$35455 ( \35832 , \35830 , \35831 );
and \U$35456 ( \35833 , \35824 , \35832 );
and \U$35457 ( \35834 , \35815 , \35823 );
or \U$35458 ( \35835 , \35833 , \35834 );
not \U$35459 ( \35836 , \789 );
and \U$35460 ( \35837 , \883 , RIae751a0_2);
and \U$35461 ( \35838 , RIae75380_6, \881 );
nor \U$35462 ( \35839 , \35837 , \35838 );
not \U$35463 ( \35840 , \35839 );
or \U$35464 ( \35841 , \35836 , \35840 );
or \U$35465 ( \35842 , \35839 , \787 );
nand \U$35466 ( \35843 , \35841 , \35842 );
and \U$35467 ( \35844 , \558 , RIae75560_10);
and \U$35468 ( \35845 , RIae75830_16, \556 );
nor \U$35469 ( \35846 , \35844 , \35845 );
and \U$35470 ( \35847 , \35846 , \504 );
not \U$35471 ( \35848 , \35846 );
and \U$35472 ( \35849 , \35848 , \562 );
nor \U$35473 ( \35850 , \35847 , \35849 );
xor \U$35474 ( \35851 , \35843 , \35850 );
and \U$35475 ( \35852 , \672 , RIae75740_14);
and \U$35476 ( \35853 , RIae75290_4, \670 );
nor \U$35477 ( \35854 , \35852 , \35853 );
and \U$35478 ( \35855 , \35854 , \588 );
not \U$35479 ( \35856 , \35854 );
and \U$35480 ( \35857 , \35856 , \587 );
nor \U$35481 ( \35858 , \35855 , \35857 );
and \U$35482 ( \35859 , \35851 , \35858 );
and \U$35483 ( \35860 , \35843 , \35850 );
or \U$35484 ( \35861 , \35859 , \35860 );
xor \U$35485 ( \35862 , \35835 , \35861 );
nand \U$35486 ( \35863 , RIae75a10_20, RIae78b48_125);
not \U$35487 ( \35864 , \35863 );
and \U$35488 ( \35865 , \35862 , \35864 );
and \U$35489 ( \35866 , \35835 , \35861 );
or \U$35490 ( \35867 , \35865 , \35866 );
not \U$35491 ( \35868 , \35867 );
xor \U$35492 ( \35869 , \35807 , \35868 );
not \U$35493 ( \35870 , \35590 );
not \U$35494 ( \35871 , \35602 );
or \U$35495 ( \35872 , \35870 , \35871 );
or \U$35496 ( \35873 , \35590 , \35602 );
nand \U$35497 ( \35874 , \35872 , \35873 );
not \U$35498 ( \35875 , \35874 );
not \U$35499 ( \35876 , \35582 );
and \U$35500 ( \35877 , \35875 , \35876 );
and \U$35501 ( \35878 , \35874 , \35582 );
nor \U$35502 ( \35879 , \35877 , \35878 );
nand \U$35503 ( \35880 , RIae75920_18, RIae78b48_125);
xor \U$35504 ( \35881 , \35879 , \35880 );
xor \U$35505 ( \35882 , \35611 , \35619 );
xor \U$35506 ( \35883 , \35882 , \35627 );
and \U$35507 ( \35884 , \35881 , \35883 );
and \U$35508 ( \35885 , \35879 , \35880 );
or \U$35509 ( \35886 , \35884 , \35885 );
and \U$35510 ( \35887 , \35869 , \35886 );
and \U$35511 ( \35888 , \35807 , \35868 );
or \U$35512 ( \35889 , \35887 , \35888 );
xor \U$35513 ( \35890 , \35254 , \35261 );
xor \U$35514 ( \35891 , \35890 , \35269 );
xor \U$35515 ( \35892 , \35279 , \35285 );
xor \U$35516 ( \35893 , \35892 , \35294 );
xor \U$35517 ( \35894 , \35891 , \35893 );
xor \U$35518 ( \35895 , \35553 , \35560 );
xor \U$35519 ( \35896 , \35895 , \35568 );
xor \U$35520 ( \35897 , \35533 , \3422 );
xor \U$35521 ( \35898 , \35897 , \35542 );
and \U$35522 ( \35899 , \35896 , \35898 );
xor \U$35523 ( \35900 , \35507 , \35514 );
xor \U$35524 ( \35901 , \35900 , \35522 );
xor \U$35525 ( \35902 , \35533 , \3422 );
xor \U$35526 ( \35903 , \35902 , \35542 );
and \U$35527 ( \35904 , \35901 , \35903 );
and \U$35528 ( \35905 , \35896 , \35901 );
or \U$35529 ( \35906 , \35899 , \35904 , \35905 );
and \U$35530 ( \35907 , \35894 , \35906 );
and \U$35531 ( \35908 , \35891 , \35893 );
or \U$35532 ( \35909 , \35907 , \35908 );
xor \U$35533 ( \35910 , \35889 , \35909 );
and \U$35534 ( \35911 , \35604 , \35630 );
nor \U$35535 ( \35912 , \35911 , \35631 );
xor \U$35536 ( \35913 , \35525 , \35545 );
xor \U$35537 ( \35914 , \35913 , \35571 );
and \U$35538 ( \35915 , \35912 , \35914 );
xor \U$35539 ( \35916 , \35361 , \35362 );
xor \U$35540 ( \35917 , \35916 , \35371 );
xor \U$35541 ( \35918 , \35634 , \35639 );
xor \U$35542 ( \35919 , \35917 , \35918 );
xor \U$35543 ( \35920 , \35525 , \35545 );
xor \U$35544 ( \35921 , \35920 , \35571 );
and \U$35545 ( \35922 , \35919 , \35921 );
and \U$35546 ( \35923 , \35912 , \35919 );
or \U$35547 ( \35924 , \35915 , \35922 , \35923 );
and \U$35548 ( \35925 , \35910 , \35924 );
and \U$35549 ( \35926 , \35889 , \35909 );
or \U$35550 ( \35927 , \35925 , \35926 );
nor \U$35551 ( \35928 , \35720 , \35927 );
nor \U$35552 ( \35929 , \35717 , \35928 );
nor \U$35553 ( \35930 , \35702 , \35929 );
nor \U$35554 ( \35931 , \35701 , \35930 );
not \U$35555 ( \35932 , \35931 );
not \U$35556 ( \35933 , \35471 );
not \U$35557 ( \35934 , \35663 );
not \U$35558 ( \35935 , \35469 );
and \U$35559 ( \35936 , \35934 , \35935 );
and \U$35560 ( \35937 , \35663 , \35469 );
nor \U$35561 ( \35938 , \35936 , \35937 );
not \U$35562 ( \35939 , \35938 );
or \U$35563 ( \35940 , \35933 , \35939 );
or \U$35564 ( \35941 , \35938 , \35471 );
nand \U$35565 ( \35942 , \35940 , \35941 );
nand \U$35566 ( \35943 , \35932 , \35942 );
or \U$35567 ( \35944 , \35682 , \35943 );
xnor \U$35568 ( \35945 , \35943 , \35682 );
xor \U$35569 ( \35946 , \35891 , \35893 );
xor \U$35570 ( \35947 , \35946 , \35906 );
xor \U$35571 ( \35948 , \35807 , \35868 );
xor \U$35572 ( \35949 , \35948 , \35886 );
xor \U$35573 ( \35950 , \35525 , \35545 );
xor \U$35574 ( \35951 , \35950 , \35571 );
xor \U$35575 ( \35952 , \35912 , \35919 );
xor \U$35576 ( \35953 , \35951 , \35952 );
xor \U$35577 ( \35954 , \35949 , \35953 );
xor \U$35578 ( \35955 , \35947 , \35954 );
not \U$35579 ( \35956 , \35955 );
not \U$35580 ( \35957 , \469 );
and \U$35581 ( \35958 , \514 , RIae75ce0_26);
and \U$35582 ( \35959 , RIae75dd0_28, \512 );
nor \U$35583 ( \35960 , \35958 , \35959 );
not \U$35584 ( \35961 , \35960 );
or \U$35585 ( \35962 , \35957 , \35961 );
or \U$35586 ( \35963 , \35960 , \469 );
nand \U$35587 ( \35964 , \35962 , \35963 );
not \U$35588 ( \35965 , \400 );
and \U$35589 ( \35966 , \436 , RIae75fb0_32);
and \U$35590 ( \35967 , RIae75ec0_30, \434 );
nor \U$35591 ( \35968 , \35966 , \35967 );
not \U$35592 ( \35969 , \35968 );
or \U$35593 ( \35970 , \35965 , \35969 );
or \U$35594 ( \35971 , \35968 , \402 );
nand \U$35595 ( \35972 , \35970 , \35971 );
xor \U$35596 ( \35973 , \35964 , \35972 );
and \U$35597 ( \35974 , \558 , RIae75650_12);
and \U$35598 ( \35975 , RIae75560_10, \556 );
nor \U$35599 ( \35976 , \35974 , \35975 );
and \U$35600 ( \35977 , \35976 , \504 );
not \U$35601 ( \35978 , \35976 );
and \U$35602 ( \35979 , \35978 , \562 );
nor \U$35603 ( \35980 , \35977 , \35979 );
and \U$35604 ( \35981 , \35973 , \35980 );
and \U$35605 ( \35982 , \35964 , \35972 );
or \U$35606 ( \35983 , \35981 , \35982 );
not \U$35607 ( \35984 , RIae75b00_22);
nor \U$35608 ( \35985 , \35984 , \491 );
not \U$35609 ( \35986 , \388 );
and \U$35610 ( \35987 , \384 , RIae75a10_20);
and \U$35611 ( \35988 , RIae75920_18, \382 );
nor \U$35612 ( \35989 , \35987 , \35988 );
not \U$35613 ( \35990 , \35989 );
or \U$35614 ( \35991 , \35986 , \35990 );
or \U$35615 ( \35992 , \35989 , \388 );
nand \U$35616 ( \35993 , \35991 , \35992 );
and \U$35617 ( \35994 , \35985 , \35993 );
xor \U$35618 ( \35995 , \35983 , \35994 );
and \U$35619 ( \35996 , \1138 , RIae75380_6);
and \U$35620 ( \35997 , RIae75470_8, \1136 );
nor \U$35621 ( \35998 , \35996 , \35997 );
and \U$35622 ( \35999 , \35998 , \1012 );
not \U$35623 ( \36000 , \35998 );
and \U$35624 ( \36001 , \36000 , \1142 );
nor \U$35625 ( \36002 , \35999 , \36001 );
and \U$35626 ( \36003 , \672 , RIae75830_16);
and \U$35627 ( \36004 , RIae75740_14, \670 );
nor \U$35628 ( \36005 , \36003 , \36004 );
and \U$35629 ( \36006 , \36005 , \588 );
not \U$35630 ( \36007 , \36005 );
and \U$35631 ( \36008 , \36007 , \587 );
nor \U$35632 ( \36009 , \36006 , \36008 );
xor \U$35633 ( \36010 , \36002 , \36009 );
not \U$35634 ( \36011 , \789 );
and \U$35635 ( \36012 , \883 , RIae75290_4);
and \U$35636 ( \36013 , RIae751a0_2, \881 );
nor \U$35637 ( \36014 , \36012 , \36013 );
not \U$35638 ( \36015 , \36014 );
or \U$35639 ( \36016 , \36011 , \36015 );
or \U$35640 ( \36017 , \36014 , \789 );
nand \U$35641 ( \36018 , \36016 , \36017 );
and \U$35642 ( \36019 , \36010 , \36018 );
and \U$35643 ( \36020 , \36002 , \36009 );
or \U$35644 ( \36021 , \36019 , \36020 );
and \U$35645 ( \36022 , \35995 , \36021 );
and \U$35646 ( \36023 , \35983 , \35994 );
or \U$35647 ( \36024 , \36022 , \36023 );
and \U$35648 ( \36025 , \3214 , RIae76be0_58);
and \U$35649 ( \36026 , RIae78ad0_124, \3212 );
nor \U$35650 ( \36027 , \36025 , \36026 );
not \U$35651 ( \36028 , \36027 );
not \U$35652 ( \36029 , \2774 );
and \U$35653 ( \36030 , \36028 , \36029 );
and \U$35654 ( \36031 , \36027 , \2774 );
nor \U$35655 ( \36032 , \36030 , \36031 );
not \U$35656 ( \36033 , \36032 );
not \U$35657 ( \36034 , \4251 );
and \U$35658 ( \36035 , \36033 , \36034 );
and \U$35659 ( \36036 , \36032 , \4251 );
and \U$35660 ( \36037 , \3730 , RIae78d28_129);
and \U$35661 ( \36038 , RIae78e18_131, \3728 );
nor \U$35662 ( \36039 , \36037 , \36038 );
and \U$35663 ( \36040 , \36039 , \3422 );
not \U$35664 ( \36041 , \36039 );
and \U$35665 ( \36042 , \36041 , \3732 );
nor \U$35666 ( \36043 , \36040 , \36042 );
nor \U$35667 ( \36044 , \36036 , \36043 );
nor \U$35668 ( \36045 , \36035 , \36044 );
and \U$35669 ( \36046 , \1376 , RIae76460_42);
and \U$35670 ( \36047 , RIae76550_44, \1374 );
nor \U$35671 ( \36048 , \36046 , \36047 );
and \U$35672 ( \36049 , \36048 , \1261 );
not \U$35673 ( \36050 , \36048 );
and \U$35674 ( \36051 , \36050 , \1380 );
nor \U$35675 ( \36052 , \36049 , \36051 );
not \U$35676 ( \36053 , \36052 );
and \U$35677 ( \36054 , \1593 , RIae76730_48);
and \U$35678 ( \36055 , RIae76640_46, \1591 );
nor \U$35679 ( \36056 , \36054 , \36055 );
and \U$35680 ( \36057 , \36056 , \1488 );
not \U$35681 ( \36058 , \36056 );
and \U$35682 ( \36059 , \36058 , \1498 );
nor \U$35683 ( \36060 , \36057 , \36059 );
not \U$35684 ( \36061 , \36060 );
and \U$35685 ( \36062 , \36053 , \36061 );
and \U$35686 ( \36063 , \36060 , \36052 );
and \U$35687 ( \36064 , \1939 , RIae76190_36);
and \U$35688 ( \36065 , RIae760a0_34, \1937 );
nor \U$35689 ( \36066 , \36064 , \36065 );
and \U$35690 ( \36067 , \36066 , \1734 );
not \U$35691 ( \36068 , \36066 );
and \U$35692 ( \36069 , \36068 , \1735 );
nor \U$35693 ( \36070 , \36067 , \36069 );
nor \U$35694 ( \36071 , \36063 , \36070 );
nor \U$35695 ( \36072 , \36062 , \36071 );
xor \U$35696 ( \36073 , \36045 , \36072 );
and \U$35697 ( \36074 , \2224 , RIae76370_40);
and \U$35698 ( \36075 , RIae76280_38, \2222 );
nor \U$35699 ( \36076 , \36074 , \36075 );
and \U$35700 ( \36077 , \36076 , \2060 );
not \U$35701 ( \36078 , \36076 );
and \U$35702 ( \36079 , \36078 , \2061 );
nor \U$35703 ( \36080 , \36077 , \36079 );
not \U$35704 ( \36081 , \36080 );
and \U$35705 ( \36082 , \2607 , RIae76af0_56);
and \U$35706 ( \36083 , RIae76a00_54, \2605 );
nor \U$35707 ( \36084 , \36082 , \36083 );
and \U$35708 ( \36085 , \36084 , \2397 );
not \U$35709 ( \36086 , \36084 );
and \U$35710 ( \36087 , \36086 , \2611 );
nor \U$35711 ( \36088 , \36085 , \36087 );
not \U$35712 ( \36089 , \36088 );
and \U$35713 ( \36090 , \36081 , \36089 );
and \U$35714 ( \36091 , \36088 , \36080 );
and \U$35715 ( \36092 , \2783 , RIae76820_50);
and \U$35716 ( \36093 , RIae76910_52, \2781 );
nor \U$35717 ( \36094 , \36092 , \36093 );
not \U$35718 ( \36095 , \36094 );
not \U$35719 ( \36096 , \2789 );
and \U$35720 ( \36097 , \36095 , \36096 );
and \U$35721 ( \36098 , \36094 , \3089 );
nor \U$35722 ( \36099 , \36097 , \36098 );
nor \U$35723 ( \36100 , \36091 , \36099 );
nor \U$35724 ( \36101 , \36090 , \36100 );
and \U$35725 ( \36102 , \36073 , \36101 );
and \U$35726 ( \36103 , \36045 , \36072 );
nor \U$35727 ( \36104 , \36102 , \36103 );
xor \U$35728 ( \36105 , \36024 , \36104 );
xor \U$35729 ( \36106 , \35843 , \35850 );
xor \U$35730 ( \36107 , \36106 , \35858 );
and \U$35731 ( \36108 , \35863 , \36107 );
xor \U$35732 ( \36109 , \35815 , \35823 );
xor \U$35733 ( \36110 , \36109 , \35832 );
xor \U$35734 ( \36111 , \35843 , \35850 );
xor \U$35735 ( \36112 , \36111 , \35858 );
and \U$35736 ( \36113 , \36110 , \36112 );
and \U$35737 ( \36114 , \35863 , \36110 );
or \U$35738 ( \36115 , \36108 , \36113 , \36114 );
xor \U$35739 ( \36116 , \36105 , \36115 );
not \U$35740 ( \36117 , \35775 );
xor \U$35741 ( \36118 , \35747 , \35805 );
not \U$35742 ( \36119 , \36118 );
or \U$35743 ( \36120 , \36117 , \36119 );
or \U$35744 ( \36121 , \36118 , \35775 );
nand \U$35745 ( \36122 , \36120 , \36121 );
xor \U$35746 ( \36123 , \35835 , \35861 );
not \U$35747 ( \36124 , \35863 );
xor \U$35748 ( \36125 , \36123 , \36124 );
xor \U$35749 ( \36126 , \36122 , \36125 );
and \U$35750 ( \36127 , \36116 , \36126 );
not \U$35751 ( \36128 , \36116 );
not \U$35752 ( \36129 , \36126 );
and \U$35753 ( \36130 , \36128 , \36129 );
not \U$35754 ( \36131 , \35755 );
xor \U$35755 ( \36132 , \35773 , \35763 );
not \U$35756 ( \36133 , \36132 );
or \U$35757 ( \36134 , \36131 , \36133 );
or \U$35758 ( \36135 , \36132 , \35755 );
nand \U$35759 ( \36136 , \36134 , \36135 );
not \U$35760 ( \36137 , \35728 );
xor \U$35761 ( \36138 , \35745 , \35737 );
not \U$35762 ( \36139 , \36138 );
or \U$35763 ( \36140 , \36137 , \36139 );
or \U$35764 ( \36141 , \36138 , \35728 );
nand \U$35765 ( \36142 , \36140 , \36141 );
xor \U$35766 ( \36143 , \36136 , \36142 );
not \U$35767 ( \36144 , \35785 );
xor \U$35768 ( \36145 , \35793 , \35803 );
not \U$35769 ( \36146 , \36145 );
or \U$35770 ( \36147 , \36144 , \36146 );
or \U$35771 ( \36148 , \36145 , \35785 );
nand \U$35772 ( \36149 , \36147 , \36148 );
and \U$35773 ( \36150 , \36143 , \36149 );
and \U$35774 ( \36151 , \36136 , \36142 );
or \U$35775 ( \36152 , \36150 , \36151 );
not \U$35776 ( \36153 , \36152 );
xor \U$35777 ( \36154 , \35533 , \3422 );
xor \U$35778 ( \36155 , \36154 , \35542 );
xor \U$35779 ( \36156 , \35896 , \35901 );
xor \U$35780 ( \36157 , \36155 , \36156 );
not \U$35781 ( \36158 , \36157 );
or \U$35782 ( \36159 , \36153 , \36158 );
or \U$35783 ( \36160 , \36157 , \36152 );
nand \U$35784 ( \36161 , \36159 , \36160 );
not \U$35785 ( \36162 , \36161 );
xor \U$35786 ( \36163 , \35879 , \35880 );
xor \U$35787 ( \36164 , \36163 , \35883 );
not \U$35788 ( \36165 , \36164 );
and \U$35789 ( \36166 , \36162 , \36165 );
and \U$35790 ( \36167 , \36161 , \36164 );
nor \U$35791 ( \36168 , \36166 , \36167 );
nor \U$35792 ( \36169 , \36130 , \36168 );
nor \U$35793 ( \36170 , \36127 , \36169 );
not \U$35794 ( \36171 , \36170 );
and \U$35795 ( \36172 , \35956 , \36171 );
and \U$35796 ( \36173 , \35955 , \36170 );
xor \U$35797 ( \36174 , \36136 , \36142 );
xor \U$35798 ( \36175 , \36174 , \36149 );
not \U$35799 ( \36176 , \36032 );
and \U$35800 ( \36177 , \36043 , \4251 );
not \U$35801 ( \36178 , \36043 );
and \U$35802 ( \36179 , \36178 , \3989 );
nor \U$35803 ( \36180 , \36177 , \36179 );
not \U$35804 ( \36181 , \36180 );
or \U$35805 ( \36182 , \36176 , \36181 );
or \U$35806 ( \36183 , \36180 , \36032 );
nand \U$35807 ( \36184 , \36182 , \36183 );
not \U$35808 ( \36185 , \36052 );
xor \U$35809 ( \36186 , \36060 , \36070 );
not \U$35810 ( \36187 , \36186 );
or \U$35811 ( \36188 , \36185 , \36187 );
or \U$35812 ( \36189 , \36186 , \36052 );
nand \U$35813 ( \36190 , \36188 , \36189 );
xor \U$35814 ( \36191 , \36184 , \36190 );
not \U$35815 ( \36192 , \36080 );
xor \U$35816 ( \36193 , \36088 , \36099 );
not \U$35817 ( \36194 , \36193 );
or \U$35818 ( \36195 , \36192 , \36194 );
or \U$35819 ( \36196 , \36193 , \36080 );
nand \U$35820 ( \36197 , \36195 , \36196 );
and \U$35821 ( \36198 , \36191 , \36197 );
and \U$35822 ( \36199 , \36184 , \36190 );
or \U$35823 ( \36200 , \36198 , \36199 );
xor \U$35824 ( \36201 , \36175 , \36200 );
xor \U$35825 ( \36202 , \35843 , \35850 );
xor \U$35826 ( \36203 , \36202 , \35858 );
xor \U$35827 ( \36204 , \35863 , \36110 );
xor \U$35828 ( \36205 , \36203 , \36204 );
and \U$35829 ( \36206 , \36201 , \36205 );
and \U$35830 ( \36207 , \36175 , \36200 );
nor \U$35831 ( \36208 , \36206 , \36207 );
not \U$35832 ( \36209 , \36208 );
xor \U$35833 ( \36210 , \36045 , \36072 );
xor \U$35834 ( \36211 , \36210 , \36101 );
not \U$35835 ( \36212 , \36211 );
xor \U$35836 ( \36213 , \35983 , \35994 );
xor \U$35837 ( \36214 , \36213 , \36021 );
nand \U$35838 ( \36215 , \36212 , \36214 );
not \U$35839 ( \36216 , \36215 );
and \U$35840 ( \36217 , \36209 , \36216 );
and \U$35841 ( \36218 , \36208 , \36215 );
and \U$35842 ( \36219 , \3214 , RIae76910_52);
and \U$35843 ( \36220 , RIae76be0_58, \3212 );
nor \U$35844 ( \36221 , \36219 , \36220 );
not \U$35845 ( \36222 , \36221 );
not \U$35846 ( \36223 , \2774 );
and \U$35847 ( \36224 , \36222 , \36223 );
and \U$35848 ( \36225 , \36221 , \2774 );
nor \U$35849 ( \36226 , \36224 , \36225 );
not \U$35850 ( \36227 , \36226 );
and \U$35851 ( \36228 , \3730 , RIae78ad0_124);
and \U$35852 ( \36229 , RIae78d28_129, \3728 );
nor \U$35853 ( \36230 , \36228 , \36229 );
and \U$35854 ( \36231 , \36230 , \3422 );
not \U$35855 ( \36232 , \36230 );
and \U$35856 ( \36233 , \36232 , \3732 );
nor \U$35857 ( \36234 , \36231 , \36233 );
not \U$35858 ( \36235 , \36234 );
and \U$35859 ( \36236 , \36227 , \36235 );
and \U$35860 ( \36237 , \36234 , \36226 );
nand \U$35861 ( \36238 , RIae78e18_131, \4247 );
and \U$35862 ( \36239 , \36238 , \4251 );
not \U$35863 ( \36240 , \36238 );
and \U$35864 ( \36241 , \36240 , \3989 );
nor \U$35865 ( \36242 , \36239 , \36241 );
nor \U$35866 ( \36243 , \36237 , \36242 );
nor \U$35867 ( \36244 , \36236 , \36243 );
and \U$35868 ( \36245 , \2224 , RIae760a0_34);
and \U$35869 ( \36246 , RIae76370_40, \2222 );
nor \U$35870 ( \36247 , \36245 , \36246 );
and \U$35871 ( \36248 , \36247 , \2060 );
not \U$35872 ( \36249 , \36247 );
and \U$35873 ( \36250 , \36249 , \2061 );
nor \U$35874 ( \36251 , \36248 , \36250 );
not \U$35875 ( \36252 , \36251 );
and \U$35876 ( \36253 , \2607 , RIae76280_38);
and \U$35877 ( \36254 , RIae76af0_56, \2605 );
nor \U$35878 ( \36255 , \36253 , \36254 );
and \U$35879 ( \36256 , \36255 , \2397 );
not \U$35880 ( \36257 , \36255 );
and \U$35881 ( \36258 , \36257 , \2611 );
nor \U$35882 ( \36259 , \36256 , \36258 );
not \U$35883 ( \36260 , \36259 );
and \U$35884 ( \36261 , \36252 , \36260 );
and \U$35885 ( \36262 , \36259 , \36251 );
and \U$35886 ( \36263 , \2783 , RIae76a00_54);
and \U$35887 ( \36264 , RIae76820_50, \2781 );
nor \U$35888 ( \36265 , \36263 , \36264 );
not \U$35889 ( \36266 , \36265 );
not \U$35890 ( \36267 , \3089 );
and \U$35891 ( \36268 , \36266 , \36267 );
and \U$35892 ( \36269 , \36265 , \3089 );
nor \U$35893 ( \36270 , \36268 , \36269 );
nor \U$35894 ( \36271 , \36262 , \36270 );
nor \U$35895 ( \36272 , \36261 , \36271 );
or \U$35896 ( \36273 , \36244 , \36272 );
not \U$35897 ( \36274 , \36244 );
not \U$35898 ( \36275 , \36272 );
or \U$35899 ( \36276 , \36274 , \36275 );
and \U$35900 ( \36277 , \1593 , RIae76550_44);
and \U$35901 ( \36278 , RIae76730_48, \1591 );
nor \U$35902 ( \36279 , \36277 , \36278 );
and \U$35903 ( \36280 , \36279 , \1498 );
not \U$35904 ( \36281 , \36279 );
and \U$35905 ( \36282 , \36281 , \1488 );
nor \U$35906 ( \36283 , \36280 , \36282 );
and \U$35907 ( \36284 , \1376 , RIae75470_8);
and \U$35908 ( \36285 , RIae76460_42, \1374 );
nor \U$35909 ( \36286 , \36284 , \36285 );
and \U$35910 ( \36287 , \36286 , \1380 );
not \U$35911 ( \36288 , \36286 );
and \U$35912 ( \36289 , \36288 , \1261 );
nor \U$35913 ( \36290 , \36287 , \36289 );
xor \U$35914 ( \36291 , \36283 , \36290 );
and \U$35915 ( \36292 , \1939 , RIae76640_46);
and \U$35916 ( \36293 , RIae76190_36, \1937 );
nor \U$35917 ( \36294 , \36292 , \36293 );
and \U$35918 ( \36295 , \36294 , \1735 );
not \U$35919 ( \36296 , \36294 );
and \U$35920 ( \36297 , \36296 , \1734 );
nor \U$35921 ( \36298 , \36295 , \36297 );
and \U$35922 ( \36299 , \36291 , \36298 );
and \U$35923 ( \36300 , \36283 , \36290 );
or \U$35924 ( \36301 , \36299 , \36300 );
nand \U$35925 ( \36302 , \36276 , \36301 );
nand \U$35926 ( \36303 , \36273 , \36302 );
and \U$35927 ( \36304 , \1138 , RIae751a0_2);
and \U$35928 ( \36305 , RIae75380_6, \1136 );
nor \U$35929 ( \36306 , \36304 , \36305 );
and \U$35930 ( \36307 , \36306 , \1012 );
not \U$35931 ( \36308 , \36306 );
and \U$35932 ( \36309 , \36308 , \1142 );
nor \U$35933 ( \36310 , \36307 , \36309 );
and \U$35934 ( \36311 , \672 , RIae75560_10);
and \U$35935 ( \36312 , RIae75830_16, \670 );
nor \U$35936 ( \36313 , \36311 , \36312 );
and \U$35937 ( \36314 , \36313 , \588 );
not \U$35938 ( \36315 , \36313 );
and \U$35939 ( \36316 , \36315 , \587 );
nor \U$35940 ( \36317 , \36314 , \36316 );
xor \U$35941 ( \36318 , \36310 , \36317 );
not \U$35942 ( \36319 , \789 );
and \U$35943 ( \36320 , \883 , RIae75740_14);
and \U$35944 ( \36321 , RIae75290_4, \881 );
nor \U$35945 ( \36322 , \36320 , \36321 );
not \U$35946 ( \36323 , \36322 );
or \U$35947 ( \36324 , \36319 , \36323 );
or \U$35948 ( \36325 , \36322 , \789 );
nand \U$35949 ( \36326 , \36324 , \36325 );
and \U$35950 ( \36327 , \36318 , \36326 );
and \U$35951 ( \36328 , \36310 , \36317 );
or \U$35952 ( \36329 , \36327 , \36328 );
nand \U$35953 ( \36330 , RIae75bf0_24, RIae78b48_125);
and \U$35954 ( \36331 , \384 , RIae75b00_22);
and \U$35955 ( \36332 , RIae75a10_20, \382 );
nor \U$35956 ( \36333 , \36331 , \36332 );
not \U$35957 ( \36334 , \36333 );
not \U$35958 ( \36335 , \388 );
and \U$35959 ( \36336 , \36334 , \36335 );
and \U$35960 ( \36337 , \36333 , \392 );
nor \U$35961 ( \36338 , \36336 , \36337 );
nand \U$35962 ( \36339 , \36330 , \36338 );
xor \U$35963 ( \36340 , \36329 , \36339 );
not \U$35964 ( \36341 , \400 );
and \U$35965 ( \36342 , \436 , RIae75920_18);
and \U$35966 ( \36343 , RIae75fb0_32, \434 );
nor \U$35967 ( \36344 , \36342 , \36343 );
not \U$35968 ( \36345 , \36344 );
or \U$35969 ( \36346 , \36341 , \36345 );
or \U$35970 ( \36347 , \36344 , \400 );
nand \U$35971 ( \36348 , \36346 , \36347 );
not \U$35972 ( \36349 , \471 );
and \U$35973 ( \36350 , \514 , RIae75ec0_30);
and \U$35974 ( \36351 , RIae75ce0_26, \512 );
nor \U$35975 ( \36352 , \36350 , \36351 );
not \U$35976 ( \36353 , \36352 );
or \U$35977 ( \36354 , \36349 , \36353 );
or \U$35978 ( \36355 , \36352 , \471 );
nand \U$35979 ( \36356 , \36354 , \36355 );
xor \U$35980 ( \36357 , \36348 , \36356 );
and \U$35981 ( \36358 , \558 , RIae75dd0_28);
and \U$35982 ( \36359 , RIae75650_12, \556 );
nor \U$35983 ( \36360 , \36358 , \36359 );
and \U$35984 ( \36361 , \36360 , \504 );
not \U$35985 ( \36362 , \36360 );
and \U$35986 ( \36363 , \36362 , \562 );
nor \U$35987 ( \36364 , \36361 , \36363 );
and \U$35988 ( \36365 , \36357 , \36364 );
and \U$35989 ( \36366 , \36348 , \36356 );
or \U$35990 ( \36367 , \36365 , \36366 );
and \U$35991 ( \36368 , \36340 , \36367 );
and \U$35992 ( \36369 , \36329 , \36339 );
or \U$35993 ( \36370 , \36368 , \36369 );
xor \U$35994 ( \36371 , \36303 , \36370 );
xor \U$35995 ( \36372 , \35964 , \35972 );
xor \U$35996 ( \36373 , \36372 , \35980 );
xor \U$35997 ( \36374 , \35985 , \35993 );
xor \U$35998 ( \36375 , \36373 , \36374 );
xor \U$35999 ( \36376 , \36002 , \36009 );
xor \U$36000 ( \36377 , \36376 , \36018 );
and \U$36001 ( \36378 , \36375 , \36377 );
and \U$36002 ( \36379 , \36373 , \36374 );
or \U$36003 ( \36380 , \36378 , \36379 );
and \U$36004 ( \36381 , \36371 , \36380 );
and \U$36005 ( \36382 , \36303 , \36370 );
nor \U$36006 ( \36383 , \36381 , \36382 );
nor \U$36007 ( \36384 , \36218 , \36383 );
nor \U$36008 ( \36385 , \36217 , \36384 );
nor \U$36009 ( \36386 , \36173 , \36385 );
nor \U$36010 ( \36387 , \36172 , \36386 );
xor \U$36011 ( \36388 , \35889 , \35909 );
xor \U$36012 ( \36389 , \36388 , \35924 );
xor \U$36013 ( \36390 , \36387 , \36389 );
xor \U$36014 ( \36391 , \36024 , \36104 );
and \U$36015 ( \36392 , \36391 , \36115 );
and \U$36016 ( \36393 , \36024 , \36104 );
or \U$36017 ( \36394 , \36392 , \36393 );
and \U$36018 ( \36395 , \36122 , \36125 );
xor \U$36019 ( \36396 , \36394 , \36395 );
or \U$36020 ( \36397 , \36164 , \36157 );
not \U$36021 ( \36398 , \36164 );
not \U$36022 ( \36399 , \36157 );
or \U$36023 ( \36400 , \36398 , \36399 );
nand \U$36024 ( \36401 , \36400 , \36152 );
nand \U$36025 ( \36402 , \36397 , \36401 );
and \U$36026 ( \36403 , \36396 , \36402 );
and \U$36027 ( \36404 , \36394 , \36395 );
or \U$36028 ( \36405 , \36403 , \36404 );
not \U$36029 ( \36406 , \36405 );
xor \U$36030 ( \36407 , \35891 , \35893 );
xor \U$36031 ( \36408 , \36407 , \35906 );
and \U$36032 ( \36409 , \35949 , \36408 );
xor \U$36033 ( \36410 , \35891 , \35893 );
xor \U$36034 ( \36411 , \36410 , \35906 );
and \U$36035 ( \36412 , \35953 , \36411 );
and \U$36036 ( \36413 , \35949 , \35953 );
or \U$36037 ( \36414 , \36409 , \36412 , \36413 );
not \U$36038 ( \36415 , \36414 );
or \U$36039 ( \36416 , \36406 , \36415 );
or \U$36040 ( \36417 , \36414 , \36405 );
nand \U$36041 ( \36418 , \36416 , \36417 );
not \U$36042 ( \36419 , \36418 );
xor \U$36043 ( \36420 , \35704 , \35706 );
xor \U$36044 ( \36421 , \36420 , \35709 );
not \U$36045 ( \36422 , \36421 );
and \U$36046 ( \36423 , \36419 , \36422 );
and \U$36047 ( \36424 , \36418 , \36421 );
nor \U$36048 ( \36425 , \36423 , \36424 );
xor \U$36049 ( \36426 , \36390 , \36425 );
not \U$36050 ( \36427 , \36426 );
xor \U$36051 ( \36428 , \36303 , \36370 );
xor \U$36052 ( \36429 , \36428 , \36380 );
not \U$36053 ( \36430 , \36214 );
not \U$36054 ( \36431 , \36211 );
or \U$36055 ( \36432 , \36430 , \36431 );
or \U$36056 ( \36433 , \36214 , \36211 );
nand \U$36057 ( \36434 , \36432 , \36433 );
xor \U$36058 ( \36435 , \36429 , \36434 );
xor \U$36059 ( \36436 , \36175 , \36200 );
xor \U$36060 ( \36437 , \36436 , \36205 );
and \U$36061 ( \36438 , \36435 , \36437 );
and \U$36062 ( \36439 , \36429 , \36434 );
or \U$36063 ( \36440 , \36438 , \36439 );
and \U$36064 ( \36441 , \1593 , RIae76460_42);
and \U$36065 ( \36442 , RIae76550_44, \1591 );
nor \U$36066 ( \36443 , \36441 , \36442 );
and \U$36067 ( \36444 , \36443 , \1498 );
not \U$36068 ( \36445 , \36443 );
and \U$36069 ( \36446 , \36445 , \1488 );
nor \U$36070 ( \36447 , \36444 , \36446 );
and \U$36071 ( \36448 , \1939 , RIae76730_48);
and \U$36072 ( \36449 , RIae76640_46, \1937 );
nor \U$36073 ( \36450 , \36448 , \36449 );
and \U$36074 ( \36451 , \36450 , \1735 );
not \U$36075 ( \36452 , \36450 );
and \U$36076 ( \36453 , \36452 , \1734 );
nor \U$36077 ( \36454 , \36451 , \36453 );
xor \U$36078 ( \36455 , \36447 , \36454 );
and \U$36079 ( \36456 , \2224 , RIae76190_36);
and \U$36080 ( \36457 , RIae760a0_34, \2222 );
nor \U$36081 ( \36458 , \36456 , \36457 );
and \U$36082 ( \36459 , \36458 , \2061 );
not \U$36083 ( \36460 , \36458 );
and \U$36084 ( \36461 , \36460 , \2060 );
nor \U$36085 ( \36462 , \36459 , \36461 );
and \U$36086 ( \36463 , \36455 , \36462 );
and \U$36087 ( \36464 , \36447 , \36454 );
or \U$36088 ( \36465 , \36463 , \36464 );
and \U$36089 ( \36466 , \4247 , RIae78d28_129);
and \U$36090 ( \36467 , RIae78e18_131, \4245 );
nor \U$36091 ( \36468 , \36466 , \36467 );
and \U$36092 ( \36469 , \36468 , \3989 );
not \U$36093 ( \36470 , \36468 );
and \U$36094 ( \36471 , \36470 , \4251 );
nor \U$36095 ( \36472 , \36469 , \36471 );
xor \U$36096 ( \36473 , \36472 , \4481 );
and \U$36097 ( \36474 , \3730 , RIae76be0_58);
and \U$36098 ( \36475 , RIae78ad0_124, \3728 );
nor \U$36099 ( \36476 , \36474 , \36475 );
and \U$36100 ( \36477 , \36476 , \3732 );
not \U$36101 ( \36478 , \36476 );
and \U$36102 ( \36479 , \36478 , \3422 );
nor \U$36103 ( \36480 , \36477 , \36479 );
and \U$36104 ( \36481 , \36473 , \36480 );
and \U$36105 ( \36482 , \36472 , \4481 );
or \U$36106 ( \36483 , \36481 , \36482 );
xor \U$36107 ( \36484 , \36465 , \36483 );
not \U$36108 ( \36485 , \2774 );
and \U$36109 ( \36486 , \3214 , RIae76820_50);
and \U$36110 ( \36487 , RIae76910_52, \3212 );
nor \U$36111 ( \36488 , \36486 , \36487 );
not \U$36112 ( \36489 , \36488 );
or \U$36113 ( \36490 , \36485 , \36489 );
or \U$36114 ( \36491 , \36488 , \2774 );
nand \U$36115 ( \36492 , \36490 , \36491 );
and \U$36116 ( \36493 , \2607 , RIae76370_40);
and \U$36117 ( \36494 , RIae76280_38, \2605 );
nor \U$36118 ( \36495 , \36493 , \36494 );
and \U$36119 ( \36496 , \36495 , \2611 );
not \U$36120 ( \36497 , \36495 );
and \U$36121 ( \36498 , \36497 , \2397 );
nor \U$36122 ( \36499 , \36496 , \36498 );
xor \U$36123 ( \36500 , \36492 , \36499 );
not \U$36124 ( \36501 , \2789 );
and \U$36125 ( \36502 , \2783 , RIae76af0_56);
and \U$36126 ( \36503 , RIae76a00_54, \2781 );
nor \U$36127 ( \36504 , \36502 , \36503 );
not \U$36128 ( \36505 , \36504 );
or \U$36129 ( \36506 , \36501 , \36505 );
or \U$36130 ( \36507 , \36504 , \3089 );
nand \U$36131 ( \36508 , \36506 , \36507 );
and \U$36132 ( \36509 , \36500 , \36508 );
and \U$36133 ( \36510 , \36492 , \36499 );
or \U$36134 ( \36511 , \36509 , \36510 );
and \U$36135 ( \36512 , \36484 , \36511 );
and \U$36136 ( \36513 , \36465 , \36483 );
or \U$36137 ( \36514 , \36512 , \36513 );
and \U$36138 ( \36515 , \672 , RIae75650_12);
and \U$36139 ( \36516 , RIae75560_10, \670 );
nor \U$36140 ( \36517 , \36515 , \36516 );
and \U$36141 ( \36518 , \36517 , \588 );
not \U$36142 ( \36519 , \36517 );
and \U$36143 ( \36520 , \36519 , \587 );
nor \U$36144 ( \36521 , \36518 , \36520 );
not \U$36145 ( \36522 , \469 );
and \U$36146 ( \36523 , \514 , RIae75fb0_32);
and \U$36147 ( \36524 , RIae75ec0_30, \512 );
nor \U$36148 ( \36525 , \36523 , \36524 );
not \U$36149 ( \36526 , \36525 );
or \U$36150 ( \36527 , \36522 , \36526 );
or \U$36151 ( \36528 , \36525 , \471 );
nand \U$36152 ( \36529 , \36527 , \36528 );
xor \U$36153 ( \36530 , \36521 , \36529 );
and \U$36154 ( \36531 , \558 , RIae75ce0_26);
and \U$36155 ( \36532 , RIae75dd0_28, \556 );
nor \U$36156 ( \36533 , \36531 , \36532 );
and \U$36157 ( \36534 , \36533 , \504 );
not \U$36158 ( \36535 , \36533 );
and \U$36159 ( \36536 , \36535 , \562 );
nor \U$36160 ( \36537 , \36534 , \36536 );
and \U$36161 ( \36538 , \36530 , \36537 );
and \U$36162 ( \36539 , \36521 , \36529 );
or \U$36163 ( \36540 , \36538 , \36539 );
not \U$36164 ( \36541 , \402 );
and \U$36165 ( \36542 , \436 , RIae75a10_20);
and \U$36166 ( \36543 , RIae75920_18, \434 );
nor \U$36167 ( \36544 , \36542 , \36543 );
not \U$36168 ( \36545 , \36544 );
or \U$36169 ( \36546 , \36541 , \36545 );
or \U$36170 ( \36547 , \36544 , \400 );
nand \U$36171 ( \36548 , \36546 , \36547 );
not \U$36172 ( \36549 , RIae78710_116);
nor \U$36173 ( \36550 , \36549 , \491 );
xor \U$36174 ( \36551 , \36548 , \36550 );
not \U$36175 ( \36552 , \392 );
and \U$36176 ( \36553 , \384 , RIae75bf0_24);
and \U$36177 ( \36554 , RIae75b00_22, \382 );
nor \U$36178 ( \36555 , \36553 , \36554 );
not \U$36179 ( \36556 , \36555 );
or \U$36180 ( \36557 , \36552 , \36556 );
or \U$36181 ( \36558 , \36555 , \388 );
nand \U$36182 ( \36559 , \36557 , \36558 );
and \U$36183 ( \36560 , \36551 , \36559 );
and \U$36184 ( \36561 , \36548 , \36550 );
or \U$36185 ( \36562 , \36560 , \36561 );
xor \U$36186 ( \36563 , \36540 , \36562 );
and \U$36187 ( \36564 , \1376 , RIae75380_6);
and \U$36188 ( \36565 , RIae75470_8, \1374 );
nor \U$36189 ( \36566 , \36564 , \36565 );
and \U$36190 ( \36567 , \36566 , \1380 );
not \U$36191 ( \36568 , \36566 );
and \U$36192 ( \36569 , \36568 , \1261 );
nor \U$36193 ( \36570 , \36567 , \36569 );
not \U$36194 ( \36571 , \789 );
and \U$36195 ( \36572 , \883 , RIae75830_16);
and \U$36196 ( \36573 , RIae75740_14, \881 );
nor \U$36197 ( \36574 , \36572 , \36573 );
not \U$36198 ( \36575 , \36574 );
or \U$36199 ( \36576 , \36571 , \36575 );
or \U$36200 ( \36577 , \36574 , \787 );
nand \U$36201 ( \36578 , \36576 , \36577 );
xor \U$36202 ( \36579 , \36570 , \36578 );
and \U$36203 ( \36580 , \1138 , RIae75290_4);
and \U$36204 ( \36581 , RIae751a0_2, \1136 );
nor \U$36205 ( \36582 , \36580 , \36581 );
and \U$36206 ( \36583 , \36582 , \1012 );
not \U$36207 ( \36584 , \36582 );
and \U$36208 ( \36585 , \36584 , \1142 );
nor \U$36209 ( \36586 , \36583 , \36585 );
and \U$36210 ( \36587 , \36579 , \36586 );
and \U$36211 ( \36588 , \36570 , \36578 );
or \U$36212 ( \36589 , \36587 , \36588 );
and \U$36213 ( \36590 , \36563 , \36589 );
and \U$36214 ( \36591 , \36540 , \36562 );
or \U$36215 ( \36592 , \36590 , \36591 );
xor \U$36216 ( \36593 , \36514 , \36592 );
xor \U$36217 ( \36594 , \36348 , \36356 );
xor \U$36218 ( \36595 , \36594 , \36364 );
or \U$36219 ( \36596 , \36338 , \36330 );
nand \U$36220 ( \36597 , \36596 , \36339 );
xor \U$36221 ( \36598 , \36595 , \36597 );
xor \U$36222 ( \36599 , \36310 , \36317 );
xor \U$36223 ( \36600 , \36599 , \36326 );
and \U$36224 ( \36601 , \36598 , \36600 );
and \U$36225 ( \36602 , \36595 , \36597 );
or \U$36226 ( \36603 , \36601 , \36602 );
and \U$36227 ( \36604 , \36593 , \36603 );
and \U$36228 ( \36605 , \36514 , \36592 );
nor \U$36229 ( \36606 , \36604 , \36605 );
not \U$36230 ( \36607 , \36301 );
not \U$36231 ( \36608 , \36244 );
or \U$36232 ( \36609 , \36607 , \36608 );
or \U$36233 ( \36610 , \36244 , \36301 );
nand \U$36234 ( \36611 , \36609 , \36610 );
not \U$36235 ( \36612 , \36611 );
not \U$36236 ( \36613 , \36272 );
and \U$36237 ( \36614 , \36612 , \36613 );
and \U$36238 ( \36615 , \36611 , \36272 );
nor \U$36239 ( \36616 , \36614 , \36615 );
not \U$36240 ( \36617 , \36616 );
xor \U$36241 ( \36618 , \36329 , \36339 );
xor \U$36242 ( \36619 , \36618 , \36367 );
nand \U$36243 ( \36620 , \36617 , \36619 );
or \U$36244 ( \36621 , \36606 , \36620 );
not \U$36245 ( \36622 , \36620 );
not \U$36246 ( \36623 , \36606 );
or \U$36247 ( \36624 , \36622 , \36623 );
not \U$36248 ( \36625 , \36226 );
xor \U$36249 ( \36626 , \36242 , \36234 );
not \U$36250 ( \36627 , \36626 );
or \U$36251 ( \36628 , \36625 , \36627 );
or \U$36252 ( \36629 , \36626 , \36226 );
nand \U$36253 ( \36630 , \36628 , \36629 );
xor \U$36254 ( \36631 , \36283 , \36290 );
xor \U$36255 ( \36632 , \36631 , \36298 );
xor \U$36256 ( \36633 , \36630 , \36632 );
not \U$36257 ( \36634 , \36251 );
xor \U$36258 ( \36635 , \36259 , \36270 );
not \U$36259 ( \36636 , \36635 );
or \U$36260 ( \36637 , \36634 , \36636 );
or \U$36261 ( \36638 , \36635 , \36251 );
nand \U$36262 ( \36639 , \36637 , \36638 );
and \U$36263 ( \36640 , \36633 , \36639 );
and \U$36264 ( \36641 , \36630 , \36632 );
or \U$36265 ( \36642 , \36640 , \36641 );
xor \U$36266 ( \36643 , \36373 , \36374 );
xor \U$36267 ( \36644 , \36643 , \36377 );
and \U$36268 ( \36645 , \36642 , \36644 );
xor \U$36269 ( \36646 , \36184 , \36190 );
xor \U$36270 ( \36647 , \36646 , \36197 );
xor \U$36271 ( \36648 , \36373 , \36374 );
xor \U$36272 ( \36649 , \36648 , \36377 );
and \U$36273 ( \36650 , \36647 , \36649 );
and \U$36274 ( \36651 , \36642 , \36647 );
or \U$36275 ( \36652 , \36645 , \36650 , \36651 );
nand \U$36276 ( \36653 , \36624 , \36652 );
nand \U$36277 ( \36654 , \36621 , \36653 );
xor \U$36278 ( \36655 , \36440 , \36654 );
not \U$36279 ( \36656 , \36126 );
not \U$36280 ( \36657 , \36168 );
not \U$36281 ( \36658 , \36116 );
and \U$36282 ( \36659 , \36657 , \36658 );
and \U$36283 ( \36660 , \36168 , \36116 );
nor \U$36284 ( \36661 , \36659 , \36660 );
not \U$36285 ( \36662 , \36661 );
or \U$36286 ( \36663 , \36656 , \36662 );
or \U$36287 ( \36664 , \36661 , \36126 );
nand \U$36288 ( \36665 , \36663 , \36664 );
and \U$36289 ( \36666 , \36655 , \36665 );
and \U$36290 ( \36667 , \36440 , \36654 );
or \U$36291 ( \36668 , \36666 , \36667 );
xor \U$36292 ( \36669 , \36394 , \36395 );
xor \U$36293 ( \36670 , \36669 , \36402 );
xor \U$36294 ( \36671 , \36668 , \36670 );
not \U$36295 ( \36672 , \35955 );
xor \U$36296 ( \36673 , \36385 , \36170 );
not \U$36297 ( \36674 , \36673 );
or \U$36298 ( \36675 , \36672 , \36674 );
or \U$36299 ( \36676 , \36673 , \35955 );
nand \U$36300 ( \36677 , \36675 , \36676 );
and \U$36301 ( \36678 , \36671 , \36677 );
and \U$36302 ( \36679 , \36668 , \36670 );
or \U$36303 ( \36680 , \36678 , \36679 );
not \U$36304 ( \36681 , \36680 );
and \U$36305 ( \36682 , \36427 , \36681 );
and \U$36306 ( \36683 , \36426 , \36680 );
nor \U$36307 ( \36684 , \36682 , \36683 );
not \U$36308 ( \36685 , \36215 );
xor \U$36309 ( \36686 , \36383 , \36208 );
not \U$36310 ( \36687 , \36686 );
or \U$36311 ( \36688 , \36685 , \36687 );
or \U$36312 ( \36689 , \36686 , \36215 );
nand \U$36313 ( \36690 , \36688 , \36689 );
xor \U$36314 ( \36691 , \36440 , \36654 );
xor \U$36315 ( \36692 , \36691 , \36665 );
and \U$36316 ( \36693 , \36690 , \36692 );
xor \U$36317 ( \36694 , \36514 , \36592 );
xor \U$36318 ( \36695 , \36694 , \36603 );
not \U$36319 ( \36696 , \36616 );
not \U$36320 ( \36697 , \36619 );
or \U$36321 ( \36698 , \36696 , \36697 );
or \U$36322 ( \36699 , \36619 , \36616 );
nand \U$36323 ( \36700 , \36698 , \36699 );
xor \U$36324 ( \36701 , \36695 , \36700 );
xor \U$36325 ( \36702 , \36373 , \36374 );
xor \U$36326 ( \36703 , \36702 , \36377 );
xor \U$36327 ( \36704 , \36642 , \36647 );
xor \U$36328 ( \36705 , \36703 , \36704 );
and \U$36329 ( \36706 , \36701 , \36705 );
and \U$36330 ( \36707 , \36695 , \36700 );
or \U$36331 ( \36708 , \36706 , \36707 );
not \U$36332 ( \36709 , \36708 );
xor \U$36333 ( \36710 , \36429 , \36434 );
xor \U$36334 ( \36711 , \36710 , \36437 );
not \U$36335 ( \36712 , \36711 );
or \U$36336 ( \36713 , \36709 , \36712 );
or \U$36337 ( \36714 , \36711 , \36708 );
xor \U$36338 ( \36715 , \36465 , \36483 );
xor \U$36339 ( \36716 , \36715 , \36511 );
xor \U$36340 ( \36717 , \36540 , \36562 );
xor \U$36341 ( \36718 , \36717 , \36589 );
and \U$36342 ( \36719 , \36716 , \36718 );
not \U$36343 ( \36720 , \36719 );
and \U$36344 ( \36721 , \1593 , RIae75470_8);
and \U$36345 ( \36722 , RIae76460_42, \1591 );
nor \U$36346 ( \36723 , \36721 , \36722 );
and \U$36347 ( \36724 , \36723 , \1498 );
not \U$36348 ( \36725 , \36723 );
and \U$36349 ( \36726 , \36725 , \1488 );
nor \U$36350 ( \36727 , \36724 , \36726 );
and \U$36351 ( \36728 , \1939 , RIae76550_44);
and \U$36352 ( \36729 , RIae76730_48, \1937 );
nor \U$36353 ( \36730 , \36728 , \36729 );
and \U$36354 ( \36731 , \36730 , \1735 );
not \U$36355 ( \36732 , \36730 );
and \U$36356 ( \36733 , \36732 , \1734 );
nor \U$36357 ( \36734 , \36731 , \36733 );
xor \U$36358 ( \36735 , \36727 , \36734 );
and \U$36359 ( \36736 , \2224 , RIae76640_46);
and \U$36360 ( \36737 , RIae76190_36, \2222 );
nor \U$36361 ( \36738 , \36736 , \36737 );
and \U$36362 ( \36739 , \36738 , \2061 );
not \U$36363 ( \36740 , \36738 );
and \U$36364 ( \36741 , \36740 , \2060 );
nor \U$36365 ( \36742 , \36739 , \36741 );
and \U$36366 ( \36743 , \36735 , \36742 );
and \U$36367 ( \36744 , \36727 , \36734 );
or \U$36368 ( \36745 , \36743 , \36744 );
and \U$36369 ( \36746 , \3730 , RIae76910_52);
and \U$36370 ( \36747 , RIae76be0_58, \3728 );
nor \U$36371 ( \36748 , \36746 , \36747 );
and \U$36372 ( \36749 , \36748 , \3732 );
not \U$36373 ( \36750 , \36748 );
and \U$36374 ( \36751 , \36750 , \3422 );
nor \U$36375 ( \36752 , \36749 , \36751 );
nand \U$36376 ( \36753 , RIae78e18_131, \4688 );
and \U$36377 ( \36754 , \36753 , \4481 );
not \U$36378 ( \36755 , \36753 );
and \U$36379 ( \36756 , \36755 , \4482 );
nor \U$36380 ( \36757 , \36754 , \36756 );
xor \U$36381 ( \36758 , \36752 , \36757 );
and \U$36382 ( \36759 , \4247 , RIae78ad0_124);
and \U$36383 ( \36760 , RIae78d28_129, \4245 );
nor \U$36384 ( \36761 , \36759 , \36760 );
and \U$36385 ( \36762 , \36761 , \3989 );
not \U$36386 ( \36763 , \36761 );
and \U$36387 ( \36764 , \36763 , \4251 );
nor \U$36388 ( \36765 , \36762 , \36764 );
and \U$36389 ( \36766 , \36758 , \36765 );
and \U$36390 ( \36767 , \36752 , \36757 );
or \U$36391 ( \36768 , \36766 , \36767 );
xor \U$36392 ( \36769 , \36745 , \36768 );
and \U$36393 ( \36770 , \2607 , RIae760a0_34);
and \U$36394 ( \36771 , RIae76370_40, \2605 );
nor \U$36395 ( \36772 , \36770 , \36771 );
and \U$36396 ( \36773 , \36772 , \2611 );
not \U$36397 ( \36774 , \36772 );
and \U$36398 ( \36775 , \36774 , \2397 );
nor \U$36399 ( \36776 , \36773 , \36775 );
not \U$36400 ( \36777 , \3089 );
and \U$36401 ( \36778 , \2783 , RIae76280_38);
and \U$36402 ( \36779 , RIae76af0_56, \2781 );
nor \U$36403 ( \36780 , \36778 , \36779 );
not \U$36404 ( \36781 , \36780 );
or \U$36405 ( \36782 , \36777 , \36781 );
or \U$36406 ( \36783 , \36780 , \2789 );
nand \U$36407 ( \36784 , \36782 , \36783 );
xor \U$36408 ( \36785 , \36776 , \36784 );
not \U$36409 ( \36786 , \3218 );
and \U$36410 ( \36787 , \3214 , RIae76a00_54);
and \U$36411 ( \36788 , RIae76820_50, \3212 );
nor \U$36412 ( \36789 , \36787 , \36788 );
not \U$36413 ( \36790 , \36789 );
or \U$36414 ( \36791 , \36786 , \36790 );
or \U$36415 ( \36792 , \36789 , \3218 );
nand \U$36416 ( \36793 , \36791 , \36792 );
and \U$36417 ( \36794 , \36785 , \36793 );
and \U$36418 ( \36795 , \36776 , \36784 );
or \U$36419 ( \36796 , \36794 , \36795 );
and \U$36420 ( \36797 , \36769 , \36796 );
and \U$36421 ( \36798 , \36745 , \36768 );
or \U$36422 ( \36799 , \36797 , \36798 );
and \U$36423 ( \36800 , \514 , RIae75920_18);
and \U$36424 ( \36801 , RIae75fb0_32, \512 );
nor \U$36425 ( \36802 , \36800 , \36801 );
not \U$36426 ( \36803 , \36802 );
not \U$36427 ( \36804 , \471 );
and \U$36428 ( \36805 , \36803 , \36804 );
and \U$36429 ( \36806 , \36802 , \471 );
nor \U$36430 ( \36807 , \36805 , \36806 );
and \U$36431 ( \36808 , \672 , RIae75dd0_28);
and \U$36432 ( \36809 , RIae75650_12, \670 );
nor \U$36433 ( \36810 , \36808 , \36809 );
and \U$36434 ( \36811 , \36810 , \587 );
not \U$36435 ( \36812 , \36810 );
and \U$36436 ( \36813 , \36812 , \588 );
nor \U$36437 ( \36814 , \36811 , \36813 );
or \U$36438 ( \36815 , \36807 , \36814 );
not \U$36439 ( \36816 , \36814 );
not \U$36440 ( \36817 , \36807 );
or \U$36441 ( \36818 , \36816 , \36817 );
and \U$36442 ( \36819 , \558 , RIae75ec0_30);
and \U$36443 ( \36820 , RIae75ce0_26, \556 );
nor \U$36444 ( \36821 , \36819 , \36820 );
and \U$36445 ( \36822 , \36821 , \504 );
not \U$36446 ( \36823 , \36821 );
and \U$36447 ( \36824 , \36823 , \562 );
nor \U$36448 ( \36825 , \36822 , \36824 );
nand \U$36449 ( \36826 , \36818 , \36825 );
nand \U$36450 ( \36827 , \36815 , \36826 );
and \U$36451 ( \36828 , \384 , RIae78710_116);
and \U$36452 ( \36829 , RIae75bf0_24, \382 );
nor \U$36453 ( \36830 , \36828 , \36829 );
not \U$36454 ( \36831 , \36830 );
not \U$36455 ( \36832 , \392 );
and \U$36456 ( \36833 , \36831 , \36832 );
and \U$36457 ( \36834 , \36830 , \392 );
nor \U$36458 ( \36835 , \36833 , \36834 );
nand \U$36459 ( \36836 , RIae78800_118, RIae78b48_125);
or \U$36460 ( \36837 , \36835 , \36836 );
not \U$36461 ( \36838 , \36836 );
not \U$36462 ( \36839 , \36835 );
or \U$36463 ( \36840 , \36838 , \36839 );
not \U$36464 ( \36841 , \400 );
and \U$36465 ( \36842 , \436 , RIae75b00_22);
and \U$36466 ( \36843 , RIae75a10_20, \434 );
nor \U$36467 ( \36844 , \36842 , \36843 );
not \U$36468 ( \36845 , \36844 );
or \U$36469 ( \36846 , \36841 , \36845 );
or \U$36470 ( \36847 , \36844 , \400 );
nand \U$36471 ( \36848 , \36846 , \36847 );
nand \U$36472 ( \36849 , \36840 , \36848 );
nand \U$36473 ( \36850 , \36837 , \36849 );
xor \U$36474 ( \36851 , \36827 , \36850 );
and \U$36475 ( \36852 , \1376 , RIae751a0_2);
and \U$36476 ( \36853 , RIae75380_6, \1374 );
nor \U$36477 ( \36854 , \36852 , \36853 );
and \U$36478 ( \36855 , \36854 , \1380 );
not \U$36479 ( \36856 , \36854 );
and \U$36480 ( \36857 , \36856 , \1261 );
nor \U$36481 ( \36858 , \36855 , \36857 );
not \U$36482 ( \36859 , \789 );
and \U$36483 ( \36860 , \883 , RIae75560_10);
and \U$36484 ( \36861 , RIae75830_16, \881 );
nor \U$36485 ( \36862 , \36860 , \36861 );
not \U$36486 ( \36863 , \36862 );
or \U$36487 ( \36864 , \36859 , \36863 );
or \U$36488 ( \36865 , \36862 , \789 );
nand \U$36489 ( \36866 , \36864 , \36865 );
xor \U$36490 ( \36867 , \36858 , \36866 );
and \U$36491 ( \36868 , \1138 , RIae75740_14);
and \U$36492 ( \36869 , RIae75290_4, \1136 );
nor \U$36493 ( \36870 , \36868 , \36869 );
and \U$36494 ( \36871 , \36870 , \1012 );
not \U$36495 ( \36872 , \36870 );
and \U$36496 ( \36873 , \36872 , \1142 );
nor \U$36497 ( \36874 , \36871 , \36873 );
and \U$36498 ( \36875 , \36867 , \36874 );
and \U$36499 ( \36876 , \36858 , \36866 );
or \U$36500 ( \36877 , \36875 , \36876 );
and \U$36501 ( \36878 , \36851 , \36877 );
and \U$36502 ( \36879 , \36827 , \36850 );
or \U$36503 ( \36880 , \36878 , \36879 );
xor \U$36504 ( \36881 , \36799 , \36880 );
xor \U$36505 ( \36882 , \36548 , \36550 );
xor \U$36506 ( \36883 , \36882 , \36559 );
xor \U$36507 ( \36884 , \36521 , \36529 );
xor \U$36508 ( \36885 , \36884 , \36537 );
xor \U$36509 ( \36886 , \36883 , \36885 );
xor \U$36510 ( \36887 , \36570 , \36578 );
xor \U$36511 ( \36888 , \36887 , \36586 );
and \U$36512 ( \36889 , \36886 , \36888 );
and \U$36513 ( \36890 , \36883 , \36885 );
or \U$36514 ( \36891 , \36889 , \36890 );
and \U$36515 ( \36892 , \36881 , \36891 );
and \U$36516 ( \36893 , \36799 , \36880 );
or \U$36517 ( \36894 , \36892 , \36893 );
not \U$36518 ( \36895 , \36894 );
or \U$36519 ( \36896 , \36720 , \36895 );
or \U$36520 ( \36897 , \36894 , \36719 );
xor \U$36521 ( \36898 , \36472 , \4481 );
xor \U$36522 ( \36899 , \36898 , \36480 );
xor \U$36523 ( \36900 , \36447 , \36454 );
xor \U$36524 ( \36901 , \36900 , \36462 );
and \U$36525 ( \36902 , \36899 , \36901 );
xor \U$36526 ( \36903 , \36492 , \36499 );
xor \U$36527 ( \36904 , \36903 , \36508 );
xor \U$36528 ( \36905 , \36447 , \36454 );
xor \U$36529 ( \36906 , \36905 , \36462 );
and \U$36530 ( \36907 , \36904 , \36906 );
and \U$36531 ( \36908 , \36899 , \36904 );
or \U$36532 ( \36909 , \36902 , \36907 , \36908 );
xor \U$36533 ( \36910 , \36595 , \36597 );
xor \U$36534 ( \36911 , \36910 , \36600 );
and \U$36535 ( \36912 , \36909 , \36911 );
xor \U$36536 ( \36913 , \36630 , \36632 );
xor \U$36537 ( \36914 , \36913 , \36639 );
xor \U$36538 ( \36915 , \36595 , \36597 );
xor \U$36539 ( \36916 , \36915 , \36600 );
and \U$36540 ( \36917 , \36914 , \36916 );
and \U$36541 ( \36918 , \36909 , \36914 );
or \U$36542 ( \36919 , \36912 , \36917 , \36918 );
nand \U$36543 ( \36920 , \36897 , \36919 );
nand \U$36544 ( \36921 , \36896 , \36920 );
nand \U$36545 ( \36922 , \36714 , \36921 );
nand \U$36546 ( \36923 , \36713 , \36922 );
xor \U$36547 ( \36924 , \36440 , \36654 );
xor \U$36548 ( \36925 , \36924 , \36665 );
and \U$36549 ( \36926 , \36923 , \36925 );
and \U$36550 ( \36927 , \36690 , \36923 );
or \U$36551 ( \36928 , \36693 , \36926 , \36927 );
xor \U$36552 ( \36929 , \36668 , \36670 );
xor \U$36553 ( \36930 , \36929 , \36677 );
nand \U$36554 ( \36931 , \36928 , \36930 );
or \U$36555 ( \36932 , \36684 , \36931 );
xnor \U$36556 ( \36933 , \36931 , \36684 );
xor \U$36557 ( \36934 , \36928 , \36930 );
xor \U$36558 ( \36935 , \36440 , \36654 );
xor \U$36559 ( \36936 , \36935 , \36665 );
xor \U$36560 ( \36937 , \36690 , \36923 );
xor \U$36561 ( \36938 , \36936 , \36937 );
not \U$36562 ( \36939 , \36938 );
xnor \U$36563 ( \36940 , \36921 , \36708 );
not \U$36564 ( \36941 , \36940 );
not \U$36565 ( \36942 , \36711 );
and \U$36566 ( \36943 , \36941 , \36942 );
and \U$36567 ( \36944 , \36940 , \36711 );
nor \U$36568 ( \36945 , \36943 , \36944 );
not \U$36569 ( \36946 , \36606 );
not \U$36570 ( \36947 , \36652 );
or \U$36571 ( \36948 , \36946 , \36947 );
or \U$36572 ( \36949 , \36652 , \36606 );
nand \U$36573 ( \36950 , \36948 , \36949 );
not \U$36574 ( \36951 , \36950 );
not \U$36575 ( \36952 , \36620 );
and \U$36576 ( \36953 , \36951 , \36952 );
and \U$36577 ( \36954 , \36950 , \36620 );
nor \U$36578 ( \36955 , \36953 , \36954 );
xor \U$36579 ( \36956 , \36945 , \36955 );
xor \U$36580 ( \36957 , \36695 , \36700 );
xor \U$36581 ( \36958 , \36957 , \36705 );
xor \U$36582 ( \36959 , \36716 , \36718 );
xor \U$36583 ( \36960 , \36799 , \36880 );
xor \U$36584 ( \36961 , \36960 , \36891 );
and \U$36585 ( \36962 , \36959 , \36961 );
xor \U$36586 ( \36963 , \36595 , \36597 );
xor \U$36587 ( \36964 , \36963 , \36600 );
xor \U$36588 ( \36965 , \36909 , \36914 );
xor \U$36589 ( \36966 , \36964 , \36965 );
xor \U$36590 ( \36967 , \36799 , \36880 );
xor \U$36591 ( \36968 , \36967 , \36891 );
and \U$36592 ( \36969 , \36966 , \36968 );
and \U$36593 ( \36970 , \36959 , \36966 );
or \U$36594 ( \36971 , \36962 , \36969 , \36970 );
xor \U$36595 ( \36972 , \36958 , \36971 );
and \U$36596 ( \36973 , \2607 , RIae76190_36);
and \U$36597 ( \36974 , RIae760a0_34, \2605 );
nor \U$36598 ( \36975 , \36973 , \36974 );
and \U$36599 ( \36976 , \36975 , \2611 );
not \U$36600 ( \36977 , \36975 );
and \U$36601 ( \36978 , \36977 , \2397 );
nor \U$36602 ( \36979 , \36976 , \36978 );
and \U$36603 ( \36980 , \1939 , RIae76460_42);
and \U$36604 ( \36981 , RIae76550_44, \1937 );
nor \U$36605 ( \36982 , \36980 , \36981 );
and \U$36606 ( \36983 , \36982 , \1735 );
not \U$36607 ( \36984 , \36982 );
and \U$36608 ( \36985 , \36984 , \1734 );
nor \U$36609 ( \36986 , \36983 , \36985 );
xor \U$36610 ( \36987 , \36979 , \36986 );
and \U$36611 ( \36988 , \2224 , RIae76730_48);
and \U$36612 ( \36989 , RIae76640_46, \2222 );
nor \U$36613 ( \36990 , \36988 , \36989 );
and \U$36614 ( \36991 , \36990 , \2061 );
not \U$36615 ( \36992 , \36990 );
and \U$36616 ( \36993 , \36992 , \2060 );
nor \U$36617 ( \36994 , \36991 , \36993 );
and \U$36618 ( \36995 , \36987 , \36994 );
and \U$36619 ( \36996 , \36979 , \36986 );
or \U$36620 ( \36997 , \36995 , \36996 );
and \U$36621 ( \36998 , \4688 , RIae78d28_129);
and \U$36622 ( \36999 , RIae78e18_131, \4686 );
nor \U$36623 ( \37000 , \36998 , \36999 );
and \U$36624 ( \37001 , \37000 , \4481 );
not \U$36625 ( \37002 , \37000 );
and \U$36626 ( \37003 , \37002 , \4482 );
nor \U$36627 ( \37004 , \37001 , \37003 );
xor \U$36628 ( \37005 , \37004 , \5016 );
and \U$36629 ( \37006 , \4247 , RIae76be0_58);
and \U$36630 ( \37007 , RIae78ad0_124, \4245 );
nor \U$36631 ( \37008 , \37006 , \37007 );
and \U$36632 ( \37009 , \37008 , \3989 );
not \U$36633 ( \37010 , \37008 );
and \U$36634 ( \37011 , \37010 , \4251 );
nor \U$36635 ( \37012 , \37009 , \37011 );
and \U$36636 ( \37013 , \37005 , \37012 );
and \U$36637 ( \37014 , \37004 , \5016 );
or \U$36638 ( \37015 , \37013 , \37014 );
xor \U$36639 ( \37016 , \36997 , \37015 );
and \U$36640 ( \37017 , \3730 , RIae76820_50);
and \U$36641 ( \37018 , RIae76910_52, \3728 );
nor \U$36642 ( \37019 , \37017 , \37018 );
and \U$36643 ( \37020 , \37019 , \3732 );
not \U$36644 ( \37021 , \37019 );
and \U$36645 ( \37022 , \37021 , \3422 );
nor \U$36646 ( \37023 , \37020 , \37022 );
not \U$36647 ( \37024 , \2789 );
and \U$36648 ( \37025 , \2783 , RIae76370_40);
and \U$36649 ( \37026 , RIae76280_38, \2781 );
nor \U$36650 ( \37027 , \37025 , \37026 );
not \U$36651 ( \37028 , \37027 );
or \U$36652 ( \37029 , \37024 , \37028 );
or \U$36653 ( \37030 , \37027 , \2789 );
nand \U$36654 ( \37031 , \37029 , \37030 );
xor \U$36655 ( \37032 , \37023 , \37031 );
not \U$36656 ( \37033 , \2774 );
and \U$36657 ( \37034 , \3214 , RIae76af0_56);
and \U$36658 ( \37035 , RIae76a00_54, \3212 );
nor \U$36659 ( \37036 , \37034 , \37035 );
not \U$36660 ( \37037 , \37036 );
or \U$36661 ( \37038 , \37033 , \37037 );
or \U$36662 ( \37039 , \37036 , \2774 );
nand \U$36663 ( \37040 , \37038 , \37039 );
and \U$36664 ( \37041 , \37032 , \37040 );
and \U$36665 ( \37042 , \37023 , \37031 );
or \U$36666 ( \37043 , \37041 , \37042 );
and \U$36667 ( \37044 , \37016 , \37043 );
and \U$36668 ( \37045 , \36997 , \37015 );
or \U$36669 ( \37046 , \37044 , \37045 );
not \U$36670 ( \37047 , \36835 );
not \U$36671 ( \37048 , \36848 );
or \U$36672 ( \37049 , \37047 , \37048 );
or \U$36673 ( \37050 , \36835 , \36848 );
nand \U$36674 ( \37051 , \37049 , \37050 );
not \U$36675 ( \37052 , \37051 );
not \U$36676 ( \37053 , \36836 );
and \U$36677 ( \37054 , \37052 , \37053 );
and \U$36678 ( \37055 , \37051 , \36836 );
nor \U$36679 ( \37056 , \37054 , \37055 );
not \U$36680 ( \37057 , \36814 );
not \U$36681 ( \37058 , \36825 );
or \U$36682 ( \37059 , \37057 , \37058 );
or \U$36683 ( \37060 , \36814 , \36825 );
nand \U$36684 ( \37061 , \37059 , \37060 );
not \U$36685 ( \37062 , \37061 );
not \U$36686 ( \37063 , \36807 );
and \U$36687 ( \37064 , \37062 , \37063 );
and \U$36688 ( \37065 , \37061 , \36807 );
nor \U$36689 ( \37066 , \37064 , \37065 );
nand \U$36690 ( \37067 , \37056 , \37066 );
xor \U$36691 ( \37068 , \37046 , \37067 );
and \U$36692 ( \37069 , \1138 , RIae75830_16);
and \U$36693 ( \37070 , RIae75740_14, \1136 );
nor \U$36694 ( \37071 , \37069 , \37070 );
and \U$36695 ( \37072 , \37071 , \1012 );
not \U$36696 ( \37073 , \37071 );
and \U$36697 ( \37074 , \37073 , \1142 );
nor \U$36698 ( \37075 , \37072 , \37074 );
and \U$36699 ( \37076 , \1376 , RIae75290_4);
and \U$36700 ( \37077 , RIae751a0_2, \1374 );
nor \U$36701 ( \37078 , \37076 , \37077 );
and \U$36702 ( \37079 , \37078 , \1380 );
not \U$36703 ( \37080 , \37078 );
and \U$36704 ( \37081 , \37080 , \1261 );
nor \U$36705 ( \37082 , \37079 , \37081 );
xor \U$36706 ( \37083 , \37075 , \37082 );
and \U$36707 ( \37084 , \1593 , RIae75380_6);
and \U$36708 ( \37085 , RIae75470_8, \1591 );
nor \U$36709 ( \37086 , \37084 , \37085 );
and \U$36710 ( \37087 , \37086 , \1498 );
not \U$36711 ( \37088 , \37086 );
and \U$36712 ( \37089 , \37088 , \1488 );
nor \U$36713 ( \37090 , \37087 , \37089 );
and \U$36714 ( \37091 , \37083 , \37090 );
and \U$36715 ( \37092 , \37075 , \37082 );
or \U$36716 ( \37093 , \37091 , \37092 );
and \U$36717 ( \37094 , \558 , RIae75fb0_32);
and \U$36718 ( \37095 , RIae75ec0_30, \556 );
nor \U$36719 ( \37096 , \37094 , \37095 );
and \U$36720 ( \37097 , \37096 , \504 );
not \U$36721 ( \37098 , \37096 );
and \U$36722 ( \37099 , \37098 , \562 );
nor \U$36723 ( \37100 , \37097 , \37099 );
and \U$36724 ( \37101 , \672 , RIae75ce0_26);
and \U$36725 ( \37102 , RIae75dd0_28, \670 );
nor \U$36726 ( \37103 , \37101 , \37102 );
and \U$36727 ( \37104 , \37103 , \588 );
not \U$36728 ( \37105 , \37103 );
and \U$36729 ( \37106 , \37105 , \587 );
nor \U$36730 ( \37107 , \37104 , \37106 );
xor \U$36731 ( \37108 , \37100 , \37107 );
not \U$36732 ( \37109 , \789 );
and \U$36733 ( \37110 , \883 , RIae75650_12);
and \U$36734 ( \37111 , RIae75560_10, \881 );
nor \U$36735 ( \37112 , \37110 , \37111 );
not \U$36736 ( \37113 , \37112 );
or \U$36737 ( \37114 , \37109 , \37113 );
or \U$36738 ( \37115 , \37112 , \787 );
nand \U$36739 ( \37116 , \37114 , \37115 );
and \U$36740 ( \37117 , \37108 , \37116 );
and \U$36741 ( \37118 , \37100 , \37107 );
or \U$36742 ( \37119 , \37117 , \37118 );
xor \U$36743 ( \37120 , \37093 , \37119 );
not \U$36744 ( \37121 , \392 );
and \U$36745 ( \37122 , \384 , RIae78800_118);
and \U$36746 ( \37123 , RIae78710_116, \382 );
nor \U$36747 ( \37124 , \37122 , \37123 );
not \U$36748 ( \37125 , \37124 );
or \U$36749 ( \37126 , \37121 , \37125 );
or \U$36750 ( \37127 , \37124 , \392 );
nand \U$36751 ( \37128 , \37126 , \37127 );
not \U$36752 ( \37129 , \402 );
and \U$36753 ( \37130 , \436 , RIae75bf0_24);
and \U$36754 ( \37131 , RIae75b00_22, \434 );
nor \U$36755 ( \37132 , \37130 , \37131 );
not \U$36756 ( \37133 , \37132 );
or \U$36757 ( \37134 , \37129 , \37133 );
or \U$36758 ( \37135 , \37132 , \400 );
nand \U$36759 ( \37136 , \37134 , \37135 );
xor \U$36760 ( \37137 , \37128 , \37136 );
not \U$36761 ( \37138 , \471 );
and \U$36762 ( \37139 , \514 , RIae75a10_20);
and \U$36763 ( \37140 , RIae75920_18, \512 );
nor \U$36764 ( \37141 , \37139 , \37140 );
not \U$36765 ( \37142 , \37141 );
or \U$36766 ( \37143 , \37138 , \37142 );
or \U$36767 ( \37144 , \37141 , \471 );
nand \U$36768 ( \37145 , \37143 , \37144 );
and \U$36769 ( \37146 , \37137 , \37145 );
and \U$36770 ( \37147 , \37128 , \37136 );
or \U$36771 ( \37148 , \37146 , \37147 );
and \U$36772 ( \37149 , \37120 , \37148 );
and \U$36773 ( \37150 , \37093 , \37119 );
or \U$36774 ( \37151 , \37149 , \37150 );
and \U$36775 ( \37152 , \37068 , \37151 );
and \U$36776 ( \37153 , \37046 , \37067 );
or \U$36777 ( \37154 , \37152 , \37153 );
xor \U$36778 ( \37155 , \36745 , \36768 );
xor \U$36779 ( \37156 , \37155 , \36796 );
xor \U$36780 ( \37157 , \36827 , \36850 );
xor \U$36781 ( \37158 , \37157 , \36877 );
and \U$36782 ( \37159 , \37156 , \37158 );
xor \U$36783 ( \37160 , \37154 , \37159 );
xor \U$36784 ( \37161 , \36858 , \36866 );
xor \U$36785 ( \37162 , \37161 , \36874 );
xor \U$36786 ( \37163 , \36776 , \36784 );
xor \U$36787 ( \37164 , \37163 , \36793 );
and \U$36788 ( \37165 , \37162 , \37164 );
xor \U$36789 ( \37166 , \36727 , \36734 );
xor \U$36790 ( \37167 , \37166 , \36742 );
xor \U$36791 ( \37168 , \36776 , \36784 );
xor \U$36792 ( \37169 , \37168 , \36793 );
and \U$36793 ( \37170 , \37167 , \37169 );
and \U$36794 ( \37171 , \37162 , \37167 );
or \U$36795 ( \37172 , \37165 , \37170 , \37171 );
xor \U$36796 ( \37173 , \36883 , \36885 );
xor \U$36797 ( \37174 , \37173 , \36888 );
and \U$36798 ( \37175 , \37172 , \37174 );
xor \U$36799 ( \37176 , \36447 , \36454 );
xor \U$36800 ( \37177 , \37176 , \36462 );
xor \U$36801 ( \37178 , \36899 , \36904 );
xor \U$36802 ( \37179 , \37177 , \37178 );
xor \U$36803 ( \37180 , \36883 , \36885 );
xor \U$36804 ( \37181 , \37180 , \36888 );
and \U$36805 ( \37182 , \37179 , \37181 );
and \U$36806 ( \37183 , \37172 , \37179 );
or \U$36807 ( \37184 , \37175 , \37182 , \37183 );
and \U$36808 ( \37185 , \37160 , \37184 );
and \U$36809 ( \37186 , \37154 , \37159 );
or \U$36810 ( \37187 , \37185 , \37186 );
and \U$36811 ( \37188 , \36972 , \37187 );
and \U$36812 ( \37189 , \36958 , \36971 );
nor \U$36813 ( \37190 , \37188 , \37189 );
and \U$36814 ( \37191 , \36956 , \37190 );
and \U$36815 ( \37192 , \36945 , \36955 );
or \U$36816 ( \37193 , \37191 , \37192 );
nor \U$36817 ( \37194 , \36939 , \37193 );
and \U$36818 ( \37195 , \36934 , \37194 );
xor \U$36819 ( \37196 , \37194 , \36934 );
and \U$36820 ( \37197 , \384 , RIae77bd0_92);
and \U$36821 ( \37198 , RIae77db0_96, \382 );
nor \U$36822 ( \37199 , \37197 , \37198 );
not \U$36823 ( \37200 , \37199 );
not \U$36824 ( \37201 , \388 );
and \U$36825 ( \37202 , \37200 , \37201 );
and \U$36826 ( \37203 , \37199 , \392 );
nor \U$36827 ( \37204 , \37202 , \37203 );
not \U$36828 ( \37205 , \37204 );
not \U$36829 ( \37206 , \402 );
and \U$36830 ( \37207 , \436 , RIae77ea0_98);
and \U$36831 ( \37208 , RIae789e0_122, \434 );
nor \U$36832 ( \37209 , \37207 , \37208 );
not \U$36833 ( \37210 , \37209 );
or \U$36834 ( \37211 , \37206 , \37210 );
or \U$36835 ( \37212 , \37209 , \402 );
nand \U$36836 ( \37213 , \37211 , \37212 );
not \U$36837 ( \37214 , \37213 );
or \U$36838 ( \37215 , \37205 , \37214 );
or \U$36839 ( \37216 , \37204 , \37213 );
nand \U$36840 ( \37217 , \37215 , \37216 );
not \U$36841 ( \37218 , \37217 );
nand \U$36842 ( \37219 , RIae77cc0_94, RIae78b48_125);
not \U$36843 ( \37220 , \37219 );
and \U$36844 ( \37221 , \37218 , \37220 );
and \U$36845 ( \37222 , \37217 , \37219 );
nor \U$36846 ( \37223 , \37221 , \37222 );
not \U$36847 ( \37224 , \402 );
and \U$36848 ( \37225 , \436 , RIae77db0_96);
and \U$36849 ( \37226 , RIae77ea0_98, \434 );
nor \U$36850 ( \37227 , \37225 , \37226 );
not \U$36851 ( \37228 , \37227 );
or \U$36852 ( \37229 , \37224 , \37228 );
or \U$36853 ( \37230 , \37227 , \400 );
nand \U$36854 ( \37231 , \37229 , \37230 );
not \U$36855 ( \37232 , \471 );
and \U$36856 ( \37233 , \514 , RIae789e0_122);
and \U$36857 ( \37234 , RIae788f0_120, \512 );
nor \U$36858 ( \37235 , \37233 , \37234 );
not \U$36859 ( \37236 , \37235 );
or \U$36860 ( \37237 , \37232 , \37236 );
or \U$36861 ( \37238 , \37235 , \471 );
nand \U$36862 ( \37239 , \37237 , \37238 );
xor \U$36863 ( \37240 , \37231 , \37239 );
not \U$36864 ( \37241 , \392 );
and \U$36865 ( \37242 , \384 , RIae77cc0_94);
and \U$36866 ( \37243 , RIae77bd0_92, \382 );
nor \U$36867 ( \37244 , \37242 , \37243 );
not \U$36868 ( \37245 , \37244 );
or \U$36869 ( \37246 , \37241 , \37245 );
or \U$36870 ( \37247 , \37244 , \388 );
nand \U$36871 ( \37248 , \37246 , \37247 );
and \U$36872 ( \37249 , \37240 , \37248 );
and \U$36873 ( \37250 , \37231 , \37239 );
nor \U$36874 ( \37251 , \37249 , \37250 );
or \U$36875 ( \37252 , \37223 , \37251 );
nand \U$36876 ( \37253 , \37251 , \37223 );
nand \U$36877 ( \37254 , \37252 , \37253 );
and \U$36878 ( \37255 , \2607 , RIae75380_6);
and \U$36879 ( \37256 , RIae75470_8, \2605 );
nor \U$36880 ( \37257 , \37255 , \37256 );
and \U$36881 ( \37258 , \37257 , \2611 );
not \U$36882 ( \37259 , \37257 );
and \U$36883 ( \37260 , \37259 , \2397 );
nor \U$36884 ( \37261 , \37258 , \37260 );
and \U$36885 ( \37262 , \1939 , RIae75830_16);
and \U$36886 ( \37263 , RIae75740_14, \1937 );
nor \U$36887 ( \37264 , \37262 , \37263 );
and \U$36888 ( \37265 , \37264 , \1735 );
not \U$36889 ( \37266 , \37264 );
and \U$36890 ( \37267 , \37266 , \1734 );
nor \U$36891 ( \37268 , \37265 , \37267 );
xor \U$36892 ( \37269 , \37261 , \37268 );
and \U$36893 ( \37270 , \2224 , RIae75290_4);
and \U$36894 ( \37271 , RIae751a0_2, \2222 );
nor \U$36895 ( \37272 , \37270 , \37271 );
and \U$36896 ( \37273 , \37272 , \2061 );
not \U$36897 ( \37274 , \37272 );
and \U$36898 ( \37275 , \37274 , \2060 );
nor \U$36899 ( \37276 , \37273 , \37275 );
and \U$36900 ( \37277 , \37269 , \37276 );
and \U$36901 ( \37278 , \37261 , \37268 );
or \U$36902 ( \37279 , \37277 , \37278 );
and \U$36903 ( \37280 , \672 , RIae75bf0_24);
and \U$36904 ( \37281 , RIae75b00_22, \670 );
nor \U$36905 ( \37282 , \37280 , \37281 );
and \U$36906 ( \37283 , \37282 , \588 );
not \U$36907 ( \37284 , \37282 );
and \U$36908 ( \37285 , \37284 , \587 );
nor \U$36909 ( \37286 , \37283 , \37285 );
and \U$36910 ( \37287 , \558 , RIae78800_118);
and \U$36911 ( \37288 , RIae78710_116, \556 );
nor \U$36912 ( \37289 , \37287 , \37288 );
and \U$36913 ( \37290 , \37289 , \504 );
not \U$36914 ( \37291 , \37289 );
and \U$36915 ( \37292 , \37291 , \562 );
nor \U$36916 ( \37293 , \37290 , \37292 );
xor \U$36917 ( \37294 , \37286 , \37293 );
not \U$36918 ( \37295 , \787 );
and \U$36919 ( \37296 , \883 , RIae75a10_20);
and \U$36920 ( \37297 , RIae75920_18, \881 );
nor \U$36921 ( \37298 , \37296 , \37297 );
not \U$36922 ( \37299 , \37298 );
or \U$36923 ( \37300 , \37295 , \37299 );
or \U$36924 ( \37301 , \37298 , \787 );
nand \U$36925 ( \37302 , \37300 , \37301 );
and \U$36926 ( \37303 , \37294 , \37302 );
and \U$36927 ( \37304 , \37286 , \37293 );
or \U$36928 ( \37305 , \37303 , \37304 );
xor \U$36929 ( \37306 , \37279 , \37305 );
and \U$36930 ( \37307 , \1593 , RIae75650_12);
and \U$36931 ( \37308 , RIae75560_10, \1591 );
nor \U$36932 ( \37309 , \37307 , \37308 );
and \U$36933 ( \37310 , \37309 , \1498 );
not \U$36934 ( \37311 , \37309 );
and \U$36935 ( \37312 , \37311 , \1488 );
nor \U$36936 ( \37313 , \37310 , \37312 );
and \U$36937 ( \37314 , \1138 , RIae75fb0_32);
and \U$36938 ( \37315 , RIae75ec0_30, \1136 );
nor \U$36939 ( \37316 , \37314 , \37315 );
and \U$36940 ( \37317 , \37316 , \1012 );
not \U$36941 ( \37318 , \37316 );
and \U$36942 ( \37319 , \37318 , \1142 );
nor \U$36943 ( \37320 , \37317 , \37319 );
xor \U$36944 ( \37321 , \37313 , \37320 );
and \U$36945 ( \37322 , \1376 , RIae75ce0_26);
and \U$36946 ( \37323 , RIae75dd0_28, \1374 );
nor \U$36947 ( \37324 , \37322 , \37323 );
and \U$36948 ( \37325 , \37324 , \1380 );
not \U$36949 ( \37326 , \37324 );
and \U$36950 ( \37327 , \37326 , \1261 );
nor \U$36951 ( \37328 , \37325 , \37327 );
and \U$36952 ( \37329 , \37321 , \37328 );
and \U$36953 ( \37330 , \37313 , \37320 );
or \U$36954 ( \37331 , \37329 , \37330 );
xor \U$36955 ( \37332 , \37306 , \37331 );
and \U$36956 ( \37333 , \37254 , \37332 );
and \U$36957 ( \37334 , \1593 , RIae75560_10);
and \U$36958 ( \37335 , RIae75830_16, \1591 );
nor \U$36959 ( \37336 , \37334 , \37335 );
and \U$36960 ( \37337 , \37336 , \1498 );
not \U$36961 ( \37338 , \37336 );
and \U$36962 ( \37339 , \37338 , \1488 );
nor \U$36963 ( \37340 , \37337 , \37339 );
and \U$36964 ( \37341 , \1939 , RIae75740_14);
and \U$36965 ( \37342 , RIae75290_4, \1937 );
nor \U$36966 ( \37343 , \37341 , \37342 );
and \U$36967 ( \37344 , \37343 , \1735 );
not \U$36968 ( \37345 , \37343 );
and \U$36969 ( \37346 , \37345 , \1734 );
nor \U$36970 ( \37347 , \37344 , \37346 );
xor \U$36971 ( \37348 , \37340 , \37347 );
and \U$36972 ( \37349 , \2224 , RIae751a0_2);
and \U$36973 ( \37350 , RIae75380_6, \2222 );
nor \U$36974 ( \37351 , \37349 , \37350 );
and \U$36975 ( \37352 , \37351 , \2061 );
not \U$36976 ( \37353 , \37351 );
and \U$36977 ( \37354 , \37353 , \2060 );
nor \U$36978 ( \37355 , \37352 , \37354 );
xor \U$36979 ( \37356 , \37348 , \37355 );
not \U$36980 ( \37357 , \469 );
and \U$36981 ( \37358 , \514 , RIae788f0_120);
and \U$36982 ( \37359 , RIae78800_118, \512 );
nor \U$36983 ( \37360 , \37358 , \37359 );
not \U$36984 ( \37361 , \37360 );
or \U$36985 ( \37362 , \37357 , \37361 );
or \U$36986 ( \37363 , \37360 , \471 );
nand \U$36987 ( \37364 , \37362 , \37363 );
and \U$36988 ( \37365 , \558 , RIae78710_116);
and \U$36989 ( \37366 , RIae75bf0_24, \556 );
nor \U$36990 ( \37367 , \37365 , \37366 );
and \U$36991 ( \37368 , \37367 , \504 );
not \U$36992 ( \37369 , \37367 );
and \U$36993 ( \37370 , \37369 , \562 );
nor \U$36994 ( \37371 , \37368 , \37370 );
xor \U$36995 ( \37372 , \37364 , \37371 );
and \U$36996 ( \37373 , \672 , RIae75b00_22);
and \U$36997 ( \37374 , RIae75a10_20, \670 );
nor \U$36998 ( \37375 , \37373 , \37374 );
and \U$36999 ( \37376 , \37375 , \588 );
not \U$37000 ( \37377 , \37375 );
and \U$37001 ( \37378 , \37377 , \587 );
nor \U$37002 ( \37379 , \37376 , \37378 );
xor \U$37003 ( \37380 , \37372 , \37379 );
and \U$37004 ( \37381 , \1376 , RIae75dd0_28);
and \U$37005 ( \37382 , RIae75650_12, \1374 );
nor \U$37006 ( \37383 , \37381 , \37382 );
and \U$37007 ( \37384 , \37383 , \1380 );
not \U$37008 ( \37385 , \37383 );
and \U$37009 ( \37386 , \37385 , \1261 );
nor \U$37010 ( \37387 , \37384 , \37386 );
not \U$37011 ( \37388 , \789 );
and \U$37012 ( \37389 , \883 , RIae75920_18);
and \U$37013 ( \37390 , RIae75fb0_32, \881 );
nor \U$37014 ( \37391 , \37389 , \37390 );
not \U$37015 ( \37392 , \37391 );
or \U$37016 ( \37393 , \37388 , \37392 );
or \U$37017 ( \37394 , \37391 , \789 );
nand \U$37018 ( \37395 , \37393 , \37394 );
xor \U$37019 ( \37396 , \37387 , \37395 );
and \U$37020 ( \37397 , \1138 , RIae75ec0_30);
and \U$37021 ( \37398 , RIae75ce0_26, \1136 );
nor \U$37022 ( \37399 , \37397 , \37398 );
and \U$37023 ( \37400 , \37399 , \1012 );
not \U$37024 ( \37401 , \37399 );
and \U$37025 ( \37402 , \37401 , \1142 );
nor \U$37026 ( \37403 , \37400 , \37402 );
xor \U$37027 ( \37404 , \37396 , \37403 );
xor \U$37028 ( \37405 , \37380 , \37404 );
xor \U$37029 ( \37406 , \37356 , \37405 );
xor \U$37030 ( \37407 , \37279 , \37305 );
xor \U$37031 ( \37408 , \37407 , \37331 );
and \U$37032 ( \37409 , \37406 , \37408 );
and \U$37033 ( \37410 , \37254 , \37406 );
or \U$37034 ( \37411 , \37333 , \37409 , \37410 );
and \U$37035 ( \37412 , \4688 , RIae76280_38);
and \U$37036 ( \37413 , RIae76af0_56, \4686 );
nor \U$37037 ( \37414 , \37412 , \37413 );
and \U$37038 ( \37415 , \37414 , \4481 );
not \U$37039 ( \37416 , \37414 );
and \U$37040 ( \37417 , \37416 , \4482 );
nor \U$37041 ( \37418 , \37415 , \37417 );
and \U$37042 ( \37419 , \4247 , RIae760a0_34);
and \U$37043 ( \37420 , RIae76370_40, \4245 );
nor \U$37044 ( \37421 , \37419 , \37420 );
and \U$37045 ( \37422 , \37421 , \3989 );
not \U$37046 ( \37423 , \37421 );
and \U$37047 ( \37424 , \37423 , \4251 );
nor \U$37048 ( \37425 , \37422 , \37424 );
xor \U$37049 ( \37426 , \37418 , \37425 );
and \U$37050 ( \37427 , \5399 , RIae76a00_54);
and \U$37051 ( \37428 , RIae76820_50, \5397 );
nor \U$37052 ( \37429 , \37427 , \37428 );
and \U$37053 ( \37430 , \37429 , \5016 );
not \U$37054 ( \37431 , \37429 );
and \U$37055 ( \37432 , \37431 , \5403 );
nor \U$37056 ( \37433 , \37430 , \37432 );
and \U$37057 ( \37434 , \37426 , \37433 );
and \U$37058 ( \37435 , \37418 , \37425 );
or \U$37059 ( \37436 , \37434 , \37435 );
and \U$37060 ( \37437 , \5896 , RIae76910_52);
and \U$37061 ( \37438 , RIae76be0_58, \5894 );
nor \U$37062 ( \37439 , \37437 , \37438 );
and \U$37063 ( \37440 , \37439 , \5590 );
not \U$37064 ( \37441 , \37439 );
and \U$37065 ( \37442 , \37441 , \5589 );
nor \U$37066 ( \37443 , \37440 , \37442 );
nand \U$37067 ( \37444 , RIae78e18_131, \6941 );
and \U$37068 ( \37445 , \37444 , \6314 );
not \U$37069 ( \37446 , \37444 );
and \U$37070 ( \37447 , \37446 , \6945 );
nor \U$37071 ( \37448 , \37445 , \37447 );
xor \U$37072 ( \37449 , \37443 , \37448 );
and \U$37073 ( \37450 , \6172 , RIae78ad0_124);
and \U$37074 ( \37451 , RIae78d28_129, \6170 );
nor \U$37075 ( \37452 , \37450 , \37451 );
and \U$37076 ( \37453 , \37452 , \6176 );
not \U$37077 ( \37454 , \37452 );
and \U$37078 ( \37455 , \37454 , \6175 );
nor \U$37079 ( \37456 , \37453 , \37455 );
and \U$37080 ( \37457 , \37449 , \37456 );
and \U$37081 ( \37458 , \37443 , \37448 );
or \U$37082 ( \37459 , \37457 , \37458 );
xor \U$37083 ( \37460 , \37436 , \37459 );
and \U$37084 ( \37461 , \3730 , RIae76640_46);
and \U$37085 ( \37462 , RIae76190_36, \3728 );
nor \U$37086 ( \37463 , \37461 , \37462 );
and \U$37087 ( \37464 , \37463 , \3732 );
not \U$37088 ( \37465 , \37463 );
and \U$37089 ( \37466 , \37465 , \3422 );
nor \U$37090 ( \37467 , \37464 , \37466 );
not \U$37091 ( \37468 , \3089 );
and \U$37092 ( \37469 , \2783 , RIae75470_8);
and \U$37093 ( \37470 , RIae76460_42, \2781 );
nor \U$37094 ( \37471 , \37469 , \37470 );
not \U$37095 ( \37472 , \37471 );
or \U$37096 ( \37473 , \37468 , \37472 );
or \U$37097 ( \37474 , \37471 , \2789 );
nand \U$37098 ( \37475 , \37473 , \37474 );
xor \U$37099 ( \37476 , \37467 , \37475 );
not \U$37100 ( \37477 , \3218 );
and \U$37101 ( \37478 , \3214 , RIae76550_44);
and \U$37102 ( \37479 , RIae76730_48, \3212 );
nor \U$37103 ( \37480 , \37478 , \37479 );
not \U$37104 ( \37481 , \37480 );
or \U$37105 ( \37482 , \37477 , \37481 );
or \U$37106 ( \37483 , \37480 , \3218 );
nand \U$37107 ( \37484 , \37482 , \37483 );
and \U$37108 ( \37485 , \37476 , \37484 );
and \U$37109 ( \37486 , \37467 , \37475 );
or \U$37110 ( \37487 , \37485 , \37486 );
and \U$37111 ( \37488 , \37460 , \37487 );
and \U$37112 ( \37489 , \37436 , \37459 );
or \U$37113 ( \37490 , \37488 , \37489 );
nand \U$37114 ( \37491 , RIae78440_110, RIae78b48_125);
not \U$37115 ( \37492 , \37491 );
not \U$37116 ( \37493 , RIae784b8_111);
nor \U$37117 ( \37494 , \37493 , \491 );
xor \U$37118 ( \37495 , \37492 , \37494 );
not \U$37119 ( \37496 , \388 );
and \U$37120 ( \37497 , \384 , RIae784b8_111);
and \U$37121 ( \37498 , RIae77cc0_94, \382 );
nor \U$37122 ( \37499 , \37497 , \37498 );
not \U$37123 ( \37500 , \37499 );
or \U$37124 ( \37501 , \37496 , \37500 );
or \U$37125 ( \37502 , \37499 , \388 );
nand \U$37126 ( \37503 , \37501 , \37502 );
not \U$37127 ( \37504 , \402 );
and \U$37128 ( \37505 , \436 , RIae77bd0_92);
and \U$37129 ( \37506 , RIae77db0_96, \434 );
nor \U$37130 ( \37507 , \37505 , \37506 );
not \U$37131 ( \37508 , \37507 );
or \U$37132 ( \37509 , \37504 , \37508 );
or \U$37133 ( \37510 , \37507 , \402 );
nand \U$37134 ( \37511 , \37509 , \37510 );
xor \U$37135 ( \37512 , \37503 , \37511 );
not \U$37136 ( \37513 , \469 );
and \U$37137 ( \37514 , \514 , RIae77ea0_98);
and \U$37138 ( \37515 , RIae789e0_122, \512 );
nor \U$37139 ( \37516 , \37514 , \37515 );
not \U$37140 ( \37517 , \37516 );
or \U$37141 ( \37518 , \37513 , \37517 );
or \U$37142 ( \37519 , \37516 , \469 );
nand \U$37143 ( \37520 , \37518 , \37519 );
and \U$37144 ( \37521 , \37512 , \37520 );
and \U$37145 ( \37522 , \37503 , \37511 );
or \U$37146 ( \37523 , \37521 , \37522 );
and \U$37147 ( \37524 , \37495 , \37523 );
and \U$37148 ( \37525 , \37492 , \37494 );
or \U$37149 ( \37526 , \37524 , \37525 );
xor \U$37150 ( \37527 , \37490 , \37526 );
and \U$37151 ( \37528 , \2607 , RIae751a0_2);
and \U$37152 ( \37529 , RIae75380_6, \2605 );
nor \U$37153 ( \37530 , \37528 , \37529 );
and \U$37154 ( \37531 , \37530 , \2611 );
not \U$37155 ( \37532 , \37530 );
and \U$37156 ( \37533 , \37532 , \2397 );
nor \U$37157 ( \37534 , \37531 , \37533 );
and \U$37158 ( \37535 , \1939 , RIae75560_10);
and \U$37159 ( \37536 , RIae75830_16, \1937 );
nor \U$37160 ( \37537 , \37535 , \37536 );
and \U$37161 ( \37538 , \37537 , \1735 );
not \U$37162 ( \37539 , \37537 );
and \U$37163 ( \37540 , \37539 , \1734 );
nor \U$37164 ( \37541 , \37538 , \37540 );
xor \U$37165 ( \37542 , \37534 , \37541 );
and \U$37166 ( \37543 , \2224 , RIae75740_14);
and \U$37167 ( \37544 , RIae75290_4, \2222 );
nor \U$37168 ( \37545 , \37543 , \37544 );
and \U$37169 ( \37546 , \37545 , \2061 );
not \U$37170 ( \37547 , \37545 );
and \U$37171 ( \37548 , \37547 , \2060 );
nor \U$37172 ( \37549 , \37546 , \37548 );
and \U$37173 ( \37550 , \37542 , \37549 );
and \U$37174 ( \37551 , \37534 , \37541 );
or \U$37175 ( \37552 , \37550 , \37551 );
and \U$37176 ( \37553 , \1376 , RIae75ec0_30);
and \U$37177 ( \37554 , RIae75ce0_26, \1374 );
nor \U$37178 ( \37555 , \37553 , \37554 );
and \U$37179 ( \37556 , \37555 , \1380 );
not \U$37180 ( \37557 , \37555 );
and \U$37181 ( \37558 , \37557 , \1261 );
nor \U$37182 ( \37559 , \37556 , \37558 );
and \U$37183 ( \37560 , \1138 , RIae75920_18);
and \U$37184 ( \37561 , RIae75fb0_32, \1136 );
nor \U$37185 ( \37562 , \37560 , \37561 );
and \U$37186 ( \37563 , \37562 , \1012 );
not \U$37187 ( \37564 , \37562 );
and \U$37188 ( \37565 , \37564 , \1142 );
nor \U$37189 ( \37566 , \37563 , \37565 );
xor \U$37190 ( \37567 , \37559 , \37566 );
and \U$37191 ( \37568 , \1593 , RIae75dd0_28);
and \U$37192 ( \37569 , RIae75650_12, \1591 );
nor \U$37193 ( \37570 , \37568 , \37569 );
and \U$37194 ( \37571 , \37570 , \1498 );
not \U$37195 ( \37572 , \37570 );
and \U$37196 ( \37573 , \37572 , \1488 );
nor \U$37197 ( \37574 , \37571 , \37573 );
and \U$37198 ( \37575 , \37567 , \37574 );
and \U$37199 ( \37576 , \37559 , \37566 );
or \U$37200 ( \37577 , \37575 , \37576 );
xor \U$37201 ( \37578 , \37552 , \37577 );
not \U$37202 ( \37579 , \787 );
and \U$37203 ( \37580 , \883 , RIae75b00_22);
and \U$37204 ( \37581 , RIae75a10_20, \881 );
nor \U$37205 ( \37582 , \37580 , \37581 );
not \U$37206 ( \37583 , \37582 );
or \U$37207 ( \37584 , \37579 , \37583 );
or \U$37208 ( \37585 , \37582 , \789 );
nand \U$37209 ( \37586 , \37584 , \37585 );
and \U$37210 ( \37587 , \558 , RIae788f0_120);
and \U$37211 ( \37588 , RIae78800_118, \556 );
nor \U$37212 ( \37589 , \37587 , \37588 );
and \U$37213 ( \37590 , \37589 , \504 );
not \U$37214 ( \37591 , \37589 );
and \U$37215 ( \37592 , \37591 , \562 );
nor \U$37216 ( \37593 , \37590 , \37592 );
xor \U$37217 ( \37594 , \37586 , \37593 );
and \U$37218 ( \37595 , \672 , RIae78710_116);
and \U$37219 ( \37596 , RIae75bf0_24, \670 );
nor \U$37220 ( \37597 , \37595 , \37596 );
and \U$37221 ( \37598 , \37597 , \588 );
not \U$37222 ( \37599 , \37597 );
and \U$37223 ( \37600 , \37599 , \587 );
nor \U$37224 ( \37601 , \37598 , \37600 );
and \U$37225 ( \37602 , \37594 , \37601 );
and \U$37226 ( \37603 , \37586 , \37593 );
or \U$37227 ( \37604 , \37602 , \37603 );
and \U$37228 ( \37605 , \37578 , \37604 );
and \U$37229 ( \37606 , \37552 , \37577 );
or \U$37230 ( \37607 , \37605 , \37606 );
and \U$37231 ( \37608 , \37527 , \37607 );
and \U$37232 ( \37609 , \37490 , \37526 );
or \U$37233 ( \37610 , \37608 , \37609 );
xor \U$37234 ( \37611 , \37411 , \37610 );
xor \U$37235 ( \37612 , \37231 , \37239 );
xor \U$37236 ( \37613 , \37612 , \37248 );
xor \U$37237 ( \37614 , \37286 , \37293 );
xor \U$37238 ( \37615 , \37614 , \37302 );
and \U$37239 ( \37616 , \37613 , \37615 );
xor \U$37240 ( \37617 , \37313 , \37320 );
xor \U$37241 ( \37618 , \37617 , \37328 );
xor \U$37242 ( \37619 , \37286 , \37293 );
xor \U$37243 ( \37620 , \37619 , \37302 );
and \U$37244 ( \37621 , \37618 , \37620 );
and \U$37245 ( \37622 , \37613 , \37618 );
or \U$37246 ( \37623 , \37616 , \37621 , \37622 );
and \U$37247 ( \37624 , \4688 , RIae76af0_56);
and \U$37248 ( \37625 , RIae76a00_54, \4686 );
nor \U$37249 ( \37626 , \37624 , \37625 );
and \U$37250 ( \37627 , \37626 , \4481 );
not \U$37251 ( \37628 , \37626 );
and \U$37252 ( \37629 , \37628 , \4482 );
nor \U$37253 ( \37630 , \37627 , \37629 );
and \U$37254 ( \37631 , \4247 , RIae76370_40);
and \U$37255 ( \37632 , RIae76280_38, \4245 );
nor \U$37256 ( \37633 , \37631 , \37632 );
and \U$37257 ( \37634 , \37633 , \3989 );
not \U$37258 ( \37635 , \37633 );
and \U$37259 ( \37636 , \37635 , \4251 );
nor \U$37260 ( \37637 , \37634 , \37636 );
xor \U$37261 ( \37638 , \37630 , \37637 );
and \U$37262 ( \37639 , \5399 , RIae76820_50);
and \U$37263 ( \37640 , RIae76910_52, \5397 );
nor \U$37264 ( \37641 , \37639 , \37640 );
and \U$37265 ( \37642 , \37641 , \5016 );
not \U$37266 ( \37643 , \37641 );
and \U$37267 ( \37644 , \37643 , \5403 );
nor \U$37268 ( \37645 , \37642 , \37644 );
xor \U$37269 ( \37646 , \37638 , \37645 );
xor \U$37270 ( \37647 , \37261 , \37268 );
xor \U$37271 ( \37648 , \37647 , \37276 );
xor \U$37272 ( \37649 , \37646 , \37648 );
and \U$37273 ( \37650 , \3730 , RIae76190_36);
and \U$37274 ( \37651 , RIae760a0_34, \3728 );
nor \U$37275 ( \37652 , \37650 , \37651 );
and \U$37276 ( \37653 , \37652 , \3732 );
not \U$37277 ( \37654 , \37652 );
and \U$37278 ( \37655 , \37654 , \3422 );
nor \U$37279 ( \37656 , \37653 , \37655 );
not \U$37280 ( \37657 , \3089 );
and \U$37281 ( \37658 , \2783 , RIae76460_42);
and \U$37282 ( \37659 , RIae76550_44, \2781 );
nor \U$37283 ( \37660 , \37658 , \37659 );
not \U$37284 ( \37661 , \37660 );
or \U$37285 ( \37662 , \37657 , \37661 );
or \U$37286 ( \37663 , \37660 , \2789 );
nand \U$37287 ( \37664 , \37662 , \37663 );
xor \U$37288 ( \37665 , \37656 , \37664 );
not \U$37289 ( \37666 , \3218 );
and \U$37290 ( \37667 , \3214 , RIae76730_48);
and \U$37291 ( \37668 , RIae76640_46, \3212 );
nor \U$37292 ( \37669 , \37667 , \37668 );
not \U$37293 ( \37670 , \37669 );
or \U$37294 ( \37671 , \37666 , \37670 );
or \U$37295 ( \37672 , \37669 , \2774 );
nand \U$37296 ( \37673 , \37671 , \37672 );
xor \U$37297 ( \37674 , \37665 , \37673 );
and \U$37298 ( \37675 , \37649 , \37674 );
and \U$37299 ( \37676 , \37646 , \37648 );
or \U$37300 ( \37677 , \37675 , \37676 );
xor \U$37301 ( \37678 , \37623 , \37677 );
and \U$37302 ( \37679 , \4688 , RIae76a00_54);
and \U$37303 ( \37680 , RIae76820_50, \4686 );
nor \U$37304 ( \37681 , \37679 , \37680 );
and \U$37305 ( \37682 , \37681 , \4481 );
not \U$37306 ( \37683 , \37681 );
and \U$37307 ( \37684 , \37683 , \4482 );
nor \U$37308 ( \37685 , \37682 , \37684 );
and \U$37309 ( \37686 , \3730 , RIae760a0_34);
and \U$37310 ( \37687 , RIae76370_40, \3728 );
nor \U$37311 ( \37688 , \37686 , \37687 );
and \U$37312 ( \37689 , \37688 , \3732 );
not \U$37313 ( \37690 , \37688 );
and \U$37314 ( \37691 , \37690 , \3422 );
nor \U$37315 ( \37692 , \37689 , \37691 );
xor \U$37316 ( \37693 , \37685 , \37692 );
and \U$37317 ( \37694 , \4247 , RIae76280_38);
and \U$37318 ( \37695 , RIae76af0_56, \4245 );
nor \U$37319 ( \37696 , \37694 , \37695 );
and \U$37320 ( \37697 , \37696 , \3989 );
not \U$37321 ( \37698 , \37696 );
and \U$37322 ( \37699 , \37698 , \4251 );
nor \U$37323 ( \37700 , \37697 , \37699 );
xor \U$37324 ( \37701 , \37693 , \37700 );
and \U$37325 ( \37702 , \5399 , RIae76910_52);
and \U$37326 ( \37703 , RIae76be0_58, \5397 );
nor \U$37327 ( \37704 , \37702 , \37703 );
and \U$37328 ( \37705 , \37704 , \5016 );
not \U$37329 ( \37706 , \37704 );
and \U$37330 ( \37707 , \37706 , \5403 );
nor \U$37331 ( \37708 , \37705 , \37707 );
nand \U$37332 ( \37709 , RIae78e18_131, \6172 );
and \U$37333 ( \37710 , \37709 , \6176 );
not \U$37334 ( \37711 , \37709 );
and \U$37335 ( \37712 , \37711 , \6175 );
nor \U$37336 ( \37713 , \37710 , \37712 );
xor \U$37337 ( \37714 , \37708 , \37713 );
and \U$37338 ( \37715 , \5896 , RIae78ad0_124);
and \U$37339 ( \37716 , RIae78d28_129, \5894 );
nor \U$37340 ( \37717 , \37715 , \37716 );
and \U$37341 ( \37718 , \37717 , \5590 );
not \U$37342 ( \37719 , \37717 );
and \U$37343 ( \37720 , \37719 , \5589 );
nor \U$37344 ( \37721 , \37718 , \37720 );
xor \U$37345 ( \37722 , \37714 , \37721 );
not \U$37346 ( \37723 , \2774 );
and \U$37347 ( \37724 , \3214 , RIae76640_46);
and \U$37348 ( \37725 , RIae76190_36, \3212 );
nor \U$37349 ( \37726 , \37724 , \37725 );
not \U$37350 ( \37727 , \37726 );
or \U$37351 ( \37728 , \37723 , \37727 );
or \U$37352 ( \37729 , \37726 , \2774 );
nand \U$37353 ( \37730 , \37728 , \37729 );
and \U$37354 ( \37731 , \2607 , RIae75470_8);
and \U$37355 ( \37732 , RIae76460_42, \2605 );
nor \U$37356 ( \37733 , \37731 , \37732 );
and \U$37357 ( \37734 , \37733 , \2611 );
not \U$37358 ( \37735 , \37733 );
and \U$37359 ( \37736 , \37735 , \2397 );
nor \U$37360 ( \37737 , \37734 , \37736 );
xor \U$37361 ( \37738 , \37730 , \37737 );
not \U$37362 ( \37739 , \3089 );
and \U$37363 ( \37740 , \2783 , RIae76550_44);
and \U$37364 ( \37741 , RIae76730_48, \2781 );
nor \U$37365 ( \37742 , \37740 , \37741 );
not \U$37366 ( \37743 , \37742 );
or \U$37367 ( \37744 , \37739 , \37743 );
or \U$37368 ( \37745 , \37742 , \3089 );
nand \U$37369 ( \37746 , \37744 , \37745 );
xor \U$37370 ( \37747 , \37738 , \37746 );
xor \U$37371 ( \37748 , \37722 , \37747 );
xor \U$37372 ( \37749 , \37701 , \37748 );
and \U$37373 ( \37750 , \37678 , \37749 );
and \U$37374 ( \37751 , \37623 , \37677 );
or \U$37375 ( \37752 , \37750 , \37751 );
and \U$37376 ( \37753 , \37611 , \37752 );
and \U$37377 ( \37754 , \37411 , \37610 );
or \U$37378 ( \37755 , \37753 , \37754 );
xor \U$37379 ( \37756 , \37340 , \37347 );
and \U$37380 ( \37757 , \37756 , \37355 );
and \U$37381 ( \37758 , \37340 , \37347 );
or \U$37382 ( \37759 , \37757 , \37758 );
xor \U$37383 ( \37760 , \37364 , \37371 );
and \U$37384 ( \37761 , \37760 , \37379 );
and \U$37385 ( \37762 , \37364 , \37371 );
or \U$37386 ( \37763 , \37761 , \37762 );
xor \U$37387 ( \37764 , \37759 , \37763 );
xor \U$37388 ( \37765 , \37387 , \37395 );
and \U$37389 ( \37766 , \37765 , \37403 );
and \U$37390 ( \37767 , \37387 , \37395 );
or \U$37391 ( \37768 , \37766 , \37767 );
xor \U$37392 ( \37769 , \37764 , \37768 );
xor \U$37393 ( \37770 , \37685 , \37692 );
and \U$37394 ( \37771 , \37770 , \37700 );
and \U$37395 ( \37772 , \37685 , \37692 );
or \U$37396 ( \37773 , \37771 , \37772 );
xor \U$37397 ( \37774 , \37708 , \37713 );
and \U$37398 ( \37775 , \37774 , \37721 );
and \U$37399 ( \37776 , \37708 , \37713 );
or \U$37400 ( \37777 , \37775 , \37776 );
xor \U$37401 ( \37778 , \37773 , \37777 );
xor \U$37402 ( \37779 , \37730 , \37737 );
and \U$37403 ( \37780 , \37779 , \37746 );
and \U$37404 ( \37781 , \37730 , \37737 );
or \U$37405 ( \37782 , \37780 , \37781 );
xor \U$37406 ( \37783 , \37778 , \37782 );
xor \U$37407 ( \37784 , \37769 , \37783 );
and \U$37408 ( \37785 , \558 , RIae75bf0_24);
and \U$37409 ( \37786 , RIae75b00_22, \556 );
nor \U$37410 ( \37787 , \37785 , \37786 );
and \U$37411 ( \37788 , \37787 , \504 );
not \U$37412 ( \37789 , \37787 );
and \U$37413 ( \37790 , \37789 , \562 );
nor \U$37414 ( \37791 , \37788 , \37790 );
not \U$37415 ( \37792 , \471 );
and \U$37416 ( \37793 , \514 , RIae78800_118);
and \U$37417 ( \37794 , RIae78710_116, \512 );
nor \U$37418 ( \37795 , \37793 , \37794 );
not \U$37419 ( \37796 , \37795 );
or \U$37420 ( \37797 , \37792 , \37796 );
or \U$37421 ( \37798 , \37795 , \471 );
nand \U$37422 ( \37799 , \37797 , \37798 );
xor \U$37423 ( \37800 , \37791 , \37799 );
and \U$37424 ( \37801 , \672 , RIae75a10_20);
and \U$37425 ( \37802 , RIae75920_18, \670 );
nor \U$37426 ( \37803 , \37801 , \37802 );
and \U$37427 ( \37804 , \37803 , \588 );
not \U$37428 ( \37805 , \37803 );
and \U$37429 ( \37806 , \37805 , \587 );
nor \U$37430 ( \37807 , \37804 , \37806 );
xor \U$37431 ( \37808 , \37800 , \37807 );
or \U$37432 ( \37809 , \37204 , \37219 );
not \U$37433 ( \37810 , \37219 );
not \U$37434 ( \37811 , \37204 );
or \U$37435 ( \37812 , \37810 , \37811 );
nand \U$37436 ( \37813 , \37812 , \37213 );
nand \U$37437 ( \37814 , \37809 , \37813 );
xor \U$37438 ( \37815 , \37808 , \37814 );
not \U$37439 ( \37816 , \392 );
and \U$37440 ( \37817 , \384 , RIae77db0_96);
and \U$37441 ( \37818 , RIae77ea0_98, \382 );
nor \U$37442 ( \37819 , \37817 , \37818 );
not \U$37443 ( \37820 , \37819 );
or \U$37444 ( \37821 , \37816 , \37820 );
or \U$37445 ( \37822 , \37819 , \388 );
nand \U$37446 ( \37823 , \37821 , \37822 );
not \U$37447 ( \37824 , RIae77bd0_92);
nor \U$37448 ( \37825 , \37824 , \491 );
xor \U$37449 ( \37826 , \37823 , \37825 );
not \U$37450 ( \37827 , \400 );
and \U$37451 ( \37828 , \436 , RIae789e0_122);
and \U$37452 ( \37829 , RIae788f0_120, \434 );
nor \U$37453 ( \37830 , \37828 , \37829 );
not \U$37454 ( \37831 , \37830 );
or \U$37455 ( \37832 , \37827 , \37831 );
or \U$37456 ( \37833 , \37830 , \402 );
nand \U$37457 ( \37834 , \37832 , \37833 );
xor \U$37458 ( \37835 , \37826 , \37834 );
xor \U$37459 ( \37836 , \37815 , \37835 );
and \U$37460 ( \37837 , \5399 , RIae76be0_58);
and \U$37461 ( \37838 , RIae78ad0_124, \5397 );
nor \U$37462 ( \37839 , \37837 , \37838 );
and \U$37463 ( \37840 , \37839 , \5016 );
not \U$37464 ( \37841 , \37839 );
and \U$37465 ( \37842 , \37841 , \5403 );
nor \U$37466 ( \37843 , \37840 , \37842 );
xor \U$37467 ( \37844 , \37843 , \6176 );
and \U$37468 ( \37845 , \5896 , RIae78d28_129);
and \U$37469 ( \37846 , RIae78e18_131, \5894 );
nor \U$37470 ( \37847 , \37845 , \37846 );
and \U$37471 ( \37848 , \37847 , \5590 );
not \U$37472 ( \37849 , \37847 );
and \U$37473 ( \37850 , \37849 , \5589 );
nor \U$37474 ( \37851 , \37848 , \37850 );
xor \U$37475 ( \37852 , \37844 , \37851 );
and \U$37476 ( \37853 , \1138 , RIae75ce0_26);
and \U$37477 ( \37854 , RIae75dd0_28, \1136 );
nor \U$37478 ( \37855 , \37853 , \37854 );
and \U$37479 ( \37856 , \37855 , \1012 );
not \U$37480 ( \37857 , \37855 );
and \U$37481 ( \37858 , \37857 , \1142 );
nor \U$37482 ( \37859 , \37856 , \37858 );
not \U$37483 ( \37860 , \787 );
and \U$37484 ( \37861 , \883 , RIae75fb0_32);
and \U$37485 ( \37862 , RIae75ec0_30, \881 );
nor \U$37486 ( \37863 , \37861 , \37862 );
not \U$37487 ( \37864 , \37863 );
or \U$37488 ( \37865 , \37860 , \37864 );
or \U$37489 ( \37866 , \37863 , \789 );
nand \U$37490 ( \37867 , \37865 , \37866 );
xor \U$37491 ( \37868 , \37859 , \37867 );
and \U$37492 ( \37869 , \1376 , RIae75650_12);
and \U$37493 ( \37870 , RIae75560_10, \1374 );
nor \U$37494 ( \37871 , \37869 , \37870 );
and \U$37495 ( \37872 , \37871 , \1380 );
not \U$37496 ( \37873 , \37871 );
and \U$37497 ( \37874 , \37873 , \1261 );
nor \U$37498 ( \37875 , \37872 , \37874 );
xor \U$37499 ( \37876 , \37868 , \37875 );
and \U$37500 ( \37877 , \1593 , RIae75830_16);
and \U$37501 ( \37878 , RIae75740_14, \1591 );
nor \U$37502 ( \37879 , \37877 , \37878 );
and \U$37503 ( \37880 , \37879 , \1498 );
not \U$37504 ( \37881 , \37879 );
and \U$37505 ( \37882 , \37881 , \1488 );
nor \U$37506 ( \37883 , \37880 , \37882 );
and \U$37507 ( \37884 , \1939 , RIae75290_4);
and \U$37508 ( \37885 , RIae751a0_2, \1937 );
nor \U$37509 ( \37886 , \37884 , \37885 );
and \U$37510 ( \37887 , \37886 , \1735 );
not \U$37511 ( \37888 , \37886 );
and \U$37512 ( \37889 , \37888 , \1734 );
nor \U$37513 ( \37890 , \37887 , \37889 );
xor \U$37514 ( \37891 , \37883 , \37890 );
and \U$37515 ( \37892 , \2224 , RIae75380_6);
and \U$37516 ( \37893 , RIae75470_8, \2222 );
nor \U$37517 ( \37894 , \37892 , \37893 );
and \U$37518 ( \37895 , \37894 , \2061 );
not \U$37519 ( \37896 , \37894 );
and \U$37520 ( \37897 , \37896 , \2060 );
nor \U$37521 ( \37898 , \37895 , \37897 );
xor \U$37522 ( \37899 , \37891 , \37898 );
and \U$37523 ( \37900 , \2607 , RIae76460_42);
and \U$37524 ( \37901 , RIae76550_44, \2605 );
nor \U$37525 ( \37902 , \37900 , \37901 );
and \U$37526 ( \37903 , \37902 , \2611 );
not \U$37527 ( \37904 , \37902 );
and \U$37528 ( \37905 , \37904 , \2397 );
nor \U$37529 ( \37906 , \37903 , \37905 );
not \U$37530 ( \37907 , \3089 );
and \U$37531 ( \37908 , \2783 , RIae76730_48);
and \U$37532 ( \37909 , RIae76640_46, \2781 );
nor \U$37533 ( \37910 , \37908 , \37909 );
not \U$37534 ( \37911 , \37910 );
or \U$37535 ( \37912 , \37907 , \37911 );
or \U$37536 ( \37913 , \37910 , \3089 );
nand \U$37537 ( \37914 , \37912 , \37913 );
xor \U$37538 ( \37915 , \37906 , \37914 );
not \U$37539 ( \37916 , \3218 );
and \U$37540 ( \37917 , \3214 , RIae76190_36);
and \U$37541 ( \37918 , RIae760a0_34, \3212 );
nor \U$37542 ( \37919 , \37917 , \37918 );
not \U$37543 ( \37920 , \37919 );
or \U$37544 ( \37921 , \37916 , \37920 );
or \U$37545 ( \37922 , \37919 , \2774 );
nand \U$37546 ( \37923 , \37921 , \37922 );
xor \U$37547 ( \37924 , \37915 , \37923 );
xor \U$37548 ( \37925 , \37899 , \37924 );
xor \U$37549 ( \37926 , \37876 , \37925 );
xor \U$37550 ( \37927 , \37852 , \37926 );
xor \U$37551 ( \37928 , \37836 , \37927 );
and \U$37552 ( \37929 , \37784 , \37928 );
and \U$37553 ( \37930 , \37769 , \37783 );
or \U$37554 ( \37931 , \37929 , \37930 );
xor \U$37555 ( \37932 , \37755 , \37931 );
and \U$37556 ( \37933 , \4247 , RIae76af0_56);
and \U$37557 ( \37934 , RIae76a00_54, \4245 );
nor \U$37558 ( \37935 , \37933 , \37934 );
and \U$37559 ( \37936 , \37935 , \3989 );
not \U$37560 ( \37937 , \37935 );
and \U$37561 ( \37938 , \37937 , \4251 );
nor \U$37562 ( \37939 , \37936 , \37938 );
and \U$37563 ( \37940 , \3730 , RIae76370_40);
and \U$37564 ( \37941 , RIae76280_38, \3728 );
nor \U$37565 ( \37942 , \37940 , \37941 );
and \U$37566 ( \37943 , \37942 , \3732 );
not \U$37567 ( \37944 , \37942 );
and \U$37568 ( \37945 , \37944 , \3422 );
nor \U$37569 ( \37946 , \37943 , \37945 );
xor \U$37570 ( \37947 , \37939 , \37946 );
and \U$37571 ( \37948 , \4688 , RIae76820_50);
and \U$37572 ( \37949 , RIae76910_52, \4686 );
nor \U$37573 ( \37950 , \37948 , \37949 );
and \U$37574 ( \37951 , \37950 , \4481 );
not \U$37575 ( \37952 , \37950 );
and \U$37576 ( \37953 , \37952 , \4482 );
nor \U$37577 ( \37954 , \37951 , \37953 );
and \U$37578 ( \37955 , \37947 , \37954 );
and \U$37579 ( \37956 , \37939 , \37946 );
or \U$37580 ( \37957 , \37955 , \37956 );
xor \U$37581 ( \37958 , \37843 , \6176 );
and \U$37582 ( \37959 , \37958 , \37851 );
and \U$37583 ( \37960 , \37843 , \6176 );
or \U$37584 ( \37961 , \37959 , \37960 );
xor \U$37585 ( \37962 , \37957 , \37961 );
xor \U$37586 ( \37963 , \37906 , \37914 );
and \U$37587 ( \37964 , \37963 , \37923 );
and \U$37588 ( \37965 , \37906 , \37914 );
or \U$37589 ( \37966 , \37964 , \37965 );
xor \U$37590 ( \37967 , \37962 , \37966 );
xor \U$37591 ( \37968 , \37883 , \37890 );
and \U$37592 ( \37969 , \37968 , \37898 );
and \U$37593 ( \37970 , \37883 , \37890 );
or \U$37594 ( \37971 , \37969 , \37970 );
xor \U$37595 ( \37972 , \37859 , \37867 );
and \U$37596 ( \37973 , \37972 , \37875 );
and \U$37597 ( \37974 , \37859 , \37867 );
or \U$37598 ( \37975 , \37973 , \37974 );
xor \U$37599 ( \37976 , \37971 , \37975 );
xor \U$37600 ( \37977 , \37791 , \37799 );
and \U$37601 ( \37978 , \37977 , \37807 );
and \U$37602 ( \37979 , \37791 , \37799 );
or \U$37603 ( \37980 , \37978 , \37979 );
xor \U$37604 ( \37981 , \37976 , \37980 );
xor \U$37605 ( \37982 , \37967 , \37981 );
xor \U$37606 ( \37983 , \37823 , \37825 );
and \U$37607 ( \37984 , \37983 , \37834 );
and \U$37608 ( \37985 , \37823 , \37825 );
or \U$37609 ( \37986 , \37984 , \37985 );
and \U$37610 ( \37987 , \384 , RIae77ea0_98);
and \U$37611 ( \37988 , RIae789e0_122, \382 );
nor \U$37612 ( \37989 , \37987 , \37988 );
not \U$37613 ( \37990 , \37989 );
not \U$37614 ( \37991 , \392 );
and \U$37615 ( \37992 , \37990 , \37991 );
and \U$37616 ( \37993 , \37989 , \388 );
nor \U$37617 ( \37994 , \37992 , \37993 );
nand \U$37618 ( \37995 , RIae77db0_96, RIae78b48_125);
or \U$37619 ( \37996 , \37994 , \37995 );
nand \U$37620 ( \37997 , \37995 , \37994 );
nand \U$37621 ( \37998 , \37996 , \37997 );
xor \U$37622 ( \37999 , \37986 , \37998 );
not \U$37623 ( \38000 , \402 );
and \U$37624 ( \38001 , \436 , RIae788f0_120);
and \U$37625 ( \38002 , RIae78800_118, \434 );
nor \U$37626 ( \38003 , \38001 , \38002 );
not \U$37627 ( \38004 , \38003 );
or \U$37628 ( \38005 , \38000 , \38004 );
or \U$37629 ( \38006 , \38003 , \402 );
nand \U$37630 ( \38007 , \38005 , \38006 );
not \U$37631 ( \38008 , \469 );
and \U$37632 ( \38009 , \514 , RIae78710_116);
and \U$37633 ( \38010 , RIae75bf0_24, \512 );
nor \U$37634 ( \38011 , \38009 , \38010 );
not \U$37635 ( \38012 , \38011 );
or \U$37636 ( \38013 , \38008 , \38012 );
or \U$37637 ( \38014 , \38011 , \469 );
nand \U$37638 ( \38015 , \38013 , \38014 );
xor \U$37639 ( \38016 , \38007 , \38015 );
and \U$37640 ( \38017 , \558 , RIae75b00_22);
and \U$37641 ( \38018 , RIae75a10_20, \556 );
nor \U$37642 ( \38019 , \38017 , \38018 );
and \U$37643 ( \38020 , \38019 , \504 );
not \U$37644 ( \38021 , \38019 );
and \U$37645 ( \38022 , \38021 , \562 );
nor \U$37646 ( \38023 , \38020 , \38022 );
xor \U$37647 ( \38024 , \38016 , \38023 );
xor \U$37648 ( \38025 , \37999 , \38024 );
xor \U$37649 ( \38026 , \37982 , \38025 );
xor \U$37650 ( \38027 , \37759 , \37763 );
and \U$37651 ( \38028 , \38027 , \37768 );
and \U$37652 ( \38029 , \37759 , \37763 );
or \U$37653 ( \38030 , \38028 , \38029 );
xor \U$37654 ( \38031 , \37773 , \37777 );
and \U$37655 ( \38032 , \38031 , \37782 );
and \U$37656 ( \38033 , \37773 , \37777 );
or \U$37657 ( \38034 , \38032 , \38033 );
xor \U$37658 ( \38035 , \38030 , \38034 );
xor \U$37659 ( \38036 , \37808 , \37814 );
and \U$37660 ( \38037 , \38036 , \37835 );
and \U$37661 ( \38038 , \37808 , \37814 );
or \U$37662 ( \38039 , \38037 , \38038 );
xor \U$37663 ( \38040 , \38035 , \38039 );
xor \U$37664 ( \38041 , \37859 , \37867 );
xor \U$37665 ( \38042 , \38041 , \37875 );
and \U$37666 ( \38043 , \37899 , \38042 );
xor \U$37667 ( \38044 , \37859 , \37867 );
xor \U$37668 ( \38045 , \38044 , \37875 );
and \U$37669 ( \38046 , \37924 , \38045 );
and \U$37670 ( \38047 , \37899 , \37924 );
or \U$37671 ( \38048 , \38043 , \38046 , \38047 );
not \U$37672 ( \38049 , \3218 );
and \U$37673 ( \38050 , \3214 , RIae760a0_34);
and \U$37674 ( \38051 , RIae76370_40, \3212 );
nor \U$37675 ( \38052 , \38050 , \38051 );
not \U$37676 ( \38053 , \38052 );
or \U$37677 ( \38054 , \38049 , \38053 );
or \U$37678 ( \38055 , \38052 , \2774 );
nand \U$37679 ( \38056 , \38054 , \38055 );
and \U$37680 ( \38057 , \3730 , RIae76280_38);
and \U$37681 ( \38058 , RIae76af0_56, \3728 );
nor \U$37682 ( \38059 , \38057 , \38058 );
and \U$37683 ( \38060 , \38059 , \3732 );
not \U$37684 ( \38061 , \38059 );
and \U$37685 ( \38062 , \38061 , \3422 );
nor \U$37686 ( \38063 , \38060 , \38062 );
xor \U$37687 ( \38064 , \38056 , \38063 );
and \U$37688 ( \38065 , \4247 , RIae76a00_54);
and \U$37689 ( \38066 , RIae76820_50, \4245 );
nor \U$37690 ( \38067 , \38065 , \38066 );
and \U$37691 ( \38068 , \38067 , \3989 );
not \U$37692 ( \38069 , \38067 );
and \U$37693 ( \38070 , \38069 , \4251 );
nor \U$37694 ( \38071 , \38068 , \38070 );
xor \U$37695 ( \38072 , \38064 , \38071 );
and \U$37696 ( \38073 , \4688 , RIae76910_52);
and \U$37697 ( \38074 , RIae76be0_58, \4686 );
nor \U$37698 ( \38075 , \38073 , \38074 );
and \U$37699 ( \38076 , \38075 , \4481 );
not \U$37700 ( \38077 , \38075 );
and \U$37701 ( \38078 , \38077 , \4482 );
nor \U$37702 ( \38079 , \38076 , \38078 );
nand \U$37703 ( \38080 , RIae78e18_131, \5896 );
and \U$37704 ( \38081 , \38080 , \5590 );
not \U$37705 ( \38082 , \38080 );
and \U$37706 ( \38083 , \38082 , \5589 );
nor \U$37707 ( \38084 , \38081 , \38083 );
xor \U$37708 ( \38085 , \38079 , \38084 );
and \U$37709 ( \38086 , \5399 , RIae78ad0_124);
and \U$37710 ( \38087 , RIae78d28_129, \5397 );
nor \U$37711 ( \38088 , \38086 , \38087 );
and \U$37712 ( \38089 , \38088 , \5016 );
not \U$37713 ( \38090 , \38088 );
and \U$37714 ( \38091 , \38090 , \5403 );
nor \U$37715 ( \38092 , \38089 , \38091 );
xor \U$37716 ( \38093 , \38085 , \38092 );
xor \U$37717 ( \38094 , \38072 , \38093 );
xor \U$37718 ( \38095 , \38048 , \38094 );
not \U$37719 ( \38096 , \3089 );
and \U$37720 ( \38097 , \2783 , RIae76640_46);
and \U$37721 ( \38098 , RIae76190_36, \2781 );
nor \U$37722 ( \38099 , \38097 , \38098 );
not \U$37723 ( \38100 , \38099 );
or \U$37724 ( \38101 , \38096 , \38100 );
or \U$37725 ( \38102 , \38099 , \3089 );
nand \U$37726 ( \38103 , \38101 , \38102 );
and \U$37727 ( \38104 , \2224 , RIae75470_8);
and \U$37728 ( \38105 , RIae76460_42, \2222 );
nor \U$37729 ( \38106 , \38104 , \38105 );
and \U$37730 ( \38107 , \38106 , \2061 );
not \U$37731 ( \38108 , \38106 );
and \U$37732 ( \38109 , \38108 , \2060 );
nor \U$37733 ( \38110 , \38107 , \38109 );
xor \U$37734 ( \38111 , \38103 , \38110 );
and \U$37735 ( \38112 , \2607 , RIae76550_44);
and \U$37736 ( \38113 , RIae76730_48, \2605 );
nor \U$37737 ( \38114 , \38112 , \38113 );
and \U$37738 ( \38115 , \38114 , \2611 );
not \U$37739 ( \38116 , \38114 );
and \U$37740 ( \38117 , \38116 , \2397 );
nor \U$37741 ( \38118 , \38115 , \38117 );
xor \U$37742 ( \38119 , \38111 , \38118 );
and \U$37743 ( \38120 , \1138 , RIae75dd0_28);
and \U$37744 ( \38121 , RIae75650_12, \1136 );
nor \U$37745 ( \38122 , \38120 , \38121 );
and \U$37746 ( \38123 , \38122 , \1012 );
not \U$37747 ( \38124 , \38122 );
and \U$37748 ( \38125 , \38124 , \1142 );
nor \U$37749 ( \38126 , \38123 , \38125 );
and \U$37750 ( \38127 , \672 , RIae75920_18);
and \U$37751 ( \38128 , RIae75fb0_32, \670 );
nor \U$37752 ( \38129 , \38127 , \38128 );
and \U$37753 ( \38130 , \38129 , \588 );
not \U$37754 ( \38131 , \38129 );
and \U$37755 ( \38132 , \38131 , \587 );
nor \U$37756 ( \38133 , \38130 , \38132 );
xor \U$37757 ( \38134 , \38126 , \38133 );
not \U$37758 ( \38135 , \787 );
and \U$37759 ( \38136 , \883 , RIae75ec0_30);
and \U$37760 ( \38137 , RIae75ce0_26, \881 );
nor \U$37761 ( \38138 , \38136 , \38137 );
not \U$37762 ( \38139 , \38138 );
or \U$37763 ( \38140 , \38135 , \38139 );
or \U$37764 ( \38141 , \38138 , \787 );
nand \U$37765 ( \38142 , \38140 , \38141 );
xor \U$37766 ( \38143 , \38134 , \38142 );
and \U$37767 ( \38144 , \1376 , RIae75560_10);
and \U$37768 ( \38145 , RIae75830_16, \1374 );
nor \U$37769 ( \38146 , \38144 , \38145 );
and \U$37770 ( \38147 , \38146 , \1380 );
not \U$37771 ( \38148 , \38146 );
and \U$37772 ( \38149 , \38148 , \1261 );
nor \U$37773 ( \38150 , \38147 , \38149 );
and \U$37774 ( \38151 , \1593 , RIae75740_14);
and \U$37775 ( \38152 , RIae75290_4, \1591 );
nor \U$37776 ( \38153 , \38151 , \38152 );
and \U$37777 ( \38154 , \38153 , \1498 );
not \U$37778 ( \38155 , \38153 );
and \U$37779 ( \38156 , \38155 , \1488 );
nor \U$37780 ( \38157 , \38154 , \38156 );
xor \U$37781 ( \38158 , \38150 , \38157 );
and \U$37782 ( \38159 , \1939 , RIae751a0_2);
and \U$37783 ( \38160 , RIae75380_6, \1937 );
nor \U$37784 ( \38161 , \38159 , \38160 );
and \U$37785 ( \38162 , \38161 , \1735 );
not \U$37786 ( \38163 , \38161 );
and \U$37787 ( \38164 , \38163 , \1734 );
nor \U$37788 ( \38165 , \38162 , \38164 );
xor \U$37789 ( \38166 , \38158 , \38165 );
xor \U$37790 ( \38167 , \38143 , \38166 );
xor \U$37791 ( \38168 , \38119 , \38167 );
xor \U$37792 ( \38169 , \38095 , \38168 );
xor \U$37793 ( \38170 , \38040 , \38169 );
xor \U$37794 ( \38171 , \38026 , \38170 );
and \U$37795 ( \38172 , \37932 , \38171 );
and \U$37796 ( \38173 , \37755 , \37931 );
or \U$37797 ( \38174 , \38172 , \38173 );
xor \U$37798 ( \38175 , \37967 , \37981 );
and \U$37799 ( \38176 , \38175 , \38025 );
and \U$37800 ( \38177 , \37967 , \37981 );
or \U$37801 ( \38178 , \38176 , \38177 );
xor \U$37802 ( \38179 , \38030 , \38034 );
and \U$37803 ( \38180 , \38179 , \38039 );
and \U$37804 ( \38181 , \38030 , \38034 );
or \U$37805 ( \38182 , \38180 , \38181 );
xor \U$37806 ( \38183 , \38178 , \38182 );
xor \U$37807 ( \38184 , \38048 , \38094 );
and \U$37808 ( \38185 , \38184 , \38168 );
and \U$37809 ( \38186 , \38048 , \38094 );
or \U$37810 ( \38187 , \38185 , \38186 );
xor \U$37811 ( \38188 , \38183 , \38187 );
xor \U$37812 ( \38189 , \38103 , \38110 );
xor \U$37813 ( \38190 , \38189 , \38118 );
and \U$37814 ( \38191 , \38143 , \38190 );
xor \U$37815 ( \38192 , \38103 , \38110 );
xor \U$37816 ( \38193 , \38192 , \38118 );
and \U$37817 ( \38194 , \38166 , \38193 );
and \U$37818 ( \38195 , \38143 , \38166 );
or \U$37819 ( \38196 , \38191 , \38194 , \38195 );
and \U$37820 ( \38197 , \38072 , \38093 );
xor \U$37821 ( \38198 , \38196 , \38197 );
and \U$37822 ( \38199 , \4247 , RIae76820_50);
and \U$37823 ( \38200 , RIae76910_52, \4245 );
nor \U$37824 ( \38201 , \38199 , \38200 );
and \U$37825 ( \38202 , \38201 , \3989 );
not \U$37826 ( \38203 , \38201 );
and \U$37827 ( \38204 , \38203 , \4251 );
nor \U$37828 ( \38205 , \38202 , \38204 );
not \U$37829 ( \38206 , \2774 );
and \U$37830 ( \38207 , \3214 , RIae76370_40);
and \U$37831 ( \38208 , RIae76280_38, \3212 );
nor \U$37832 ( \38209 , \38207 , \38208 );
not \U$37833 ( \38210 , \38209 );
or \U$37834 ( \38211 , \38206 , \38210 );
or \U$37835 ( \38212 , \38209 , \3218 );
nand \U$37836 ( \38213 , \38211 , \38212 );
xor \U$37837 ( \38214 , \38205 , \38213 );
and \U$37838 ( \38215 , \3730 , RIae76af0_56);
and \U$37839 ( \38216 , RIae76a00_54, \3728 );
nor \U$37840 ( \38217 , \38215 , \38216 );
and \U$37841 ( \38218 , \38217 , \3732 );
not \U$37842 ( \38219 , \38217 );
and \U$37843 ( \38220 , \38219 , \3422 );
nor \U$37844 ( \38221 , \38218 , \38220 );
xor \U$37845 ( \38222 , \38214 , \38221 );
and \U$37846 ( \38223 , \5399 , RIae78d28_129);
and \U$37847 ( \38224 , RIae78e18_131, \5397 );
nor \U$37848 ( \38225 , \38223 , \38224 );
and \U$37849 ( \38226 , \38225 , \5016 );
not \U$37850 ( \38227 , \38225 );
and \U$37851 ( \38228 , \38227 , \5403 );
nor \U$37852 ( \38229 , \38226 , \38228 );
xor \U$37853 ( \38230 , \38229 , \5590 );
and \U$37854 ( \38231 , \4688 , RIae76be0_58);
and \U$37855 ( \38232 , RIae78ad0_124, \4686 );
nor \U$37856 ( \38233 , \38231 , \38232 );
and \U$37857 ( \38234 , \38233 , \4481 );
not \U$37858 ( \38235 , \38233 );
and \U$37859 ( \38236 , \38235 , \4482 );
nor \U$37860 ( \38237 , \38234 , \38236 );
xor \U$37861 ( \38238 , \38230 , \38237 );
not \U$37862 ( \38239 , \3089 );
and \U$37863 ( \38240 , \2783 , RIae76190_36);
and \U$37864 ( \38241 , RIae760a0_34, \2781 );
nor \U$37865 ( \38242 , \38240 , \38241 );
not \U$37866 ( \38243 , \38242 );
or \U$37867 ( \38244 , \38239 , \38243 );
or \U$37868 ( \38245 , \38242 , \2789 );
nand \U$37869 ( \38246 , \38244 , \38245 );
and \U$37870 ( \38247 , \2224 , RIae76460_42);
and \U$37871 ( \38248 , RIae76550_44, \2222 );
nor \U$37872 ( \38249 , \38247 , \38248 );
and \U$37873 ( \38250 , \38249 , \2061 );
not \U$37874 ( \38251 , \38249 );
and \U$37875 ( \38252 , \38251 , \2060 );
nor \U$37876 ( \38253 , \38250 , \38252 );
xor \U$37877 ( \38254 , \38246 , \38253 );
and \U$37878 ( \38255 , \2607 , RIae76730_48);
and \U$37879 ( \38256 , RIae76640_46, \2605 );
nor \U$37880 ( \38257 , \38255 , \38256 );
and \U$37881 ( \38258 , \38257 , \2611 );
not \U$37882 ( \38259 , \38257 );
and \U$37883 ( \38260 , \38259 , \2396 );
nor \U$37884 ( \38261 , \38258 , \38260 );
xor \U$37885 ( \38262 , \38254 , \38261 );
xor \U$37886 ( \38263 , \38238 , \38262 );
xor \U$37887 ( \38264 , \38222 , \38263 );
xor \U$37888 ( \38265 , \38198 , \38264 );
xor \U$37889 ( \38266 , \38103 , \38110 );
and \U$37890 ( \38267 , \38266 , \38118 );
and \U$37891 ( \38268 , \38103 , \38110 );
or \U$37892 ( \38269 , \38267 , \38268 );
xor \U$37893 ( \38270 , \38079 , \38084 );
and \U$37894 ( \38271 , \38270 , \38092 );
and \U$37895 ( \38272 , \38079 , \38084 );
or \U$37896 ( \38273 , \38271 , \38272 );
xor \U$37897 ( \38274 , \38269 , \38273 );
xor \U$37898 ( \38275 , \38056 , \38063 );
and \U$37899 ( \38276 , \38275 , \38071 );
and \U$37900 ( \38277 , \38056 , \38063 );
or \U$37901 ( \38278 , \38276 , \38277 );
xor \U$37902 ( \38279 , \38274 , \38278 );
xor \U$37903 ( \38280 , \38126 , \38133 );
and \U$37904 ( \38281 , \38280 , \38142 );
and \U$37905 ( \38282 , \38126 , \38133 );
or \U$37906 ( \38283 , \38281 , \38282 );
xor \U$37907 ( \38284 , \38007 , \38015 );
and \U$37908 ( \38285 , \38284 , \38023 );
and \U$37909 ( \38286 , \38007 , \38015 );
or \U$37910 ( \38287 , \38285 , \38286 );
xor \U$37911 ( \38288 , \38283 , \38287 );
xor \U$37912 ( \38289 , \38150 , \38157 );
and \U$37913 ( \38290 , \38289 , \38165 );
and \U$37914 ( \38291 , \38150 , \38157 );
or \U$37915 ( \38292 , \38290 , \38291 );
xor \U$37916 ( \38293 , \38288 , \38292 );
not \U$37917 ( \38294 , \388 );
and \U$37918 ( \38295 , \384 , RIae789e0_122);
and \U$37919 ( \38296 , RIae788f0_120, \382 );
nor \U$37920 ( \38297 , \38295 , \38296 );
not \U$37921 ( \38298 , \38297 );
or \U$37922 ( \38299 , \38294 , \38298 );
or \U$37923 ( \38300 , \38297 , \388 );
nand \U$37924 ( \38301 , \38299 , \38300 );
not \U$37925 ( \38302 , RIae77ea0_98);
nor \U$37926 ( \38303 , \38302 , \491 );
xor \U$37927 ( \38304 , \38301 , \38303 );
xor \U$37928 ( \38305 , \38304 , \37997 );
and \U$37929 ( \38306 , \1376 , RIae75830_16);
and \U$37930 ( \38307 , RIae75740_14, \1374 );
nor \U$37931 ( \38308 , \38306 , \38307 );
and \U$37932 ( \38309 , \38308 , \1380 );
not \U$37933 ( \38310 , \38308 );
and \U$37934 ( \38311 , \38310 , \1261 );
nor \U$37935 ( \38312 , \38309 , \38311 );
and \U$37936 ( \38313 , \1593 , RIae75290_4);
and \U$37937 ( \38314 , RIae751a0_2, \1591 );
nor \U$37938 ( \38315 , \38313 , \38314 );
and \U$37939 ( \38316 , \38315 , \1498 );
not \U$37940 ( \38317 , \38315 );
and \U$37941 ( \38318 , \38317 , \1488 );
nor \U$37942 ( \38319 , \38316 , \38318 );
xor \U$37943 ( \38320 , \38312 , \38319 );
and \U$37944 ( \38321 , \1939 , RIae75380_6);
and \U$37945 ( \38322 , RIae75470_8, \1937 );
nor \U$37946 ( \38323 , \38321 , \38322 );
and \U$37947 ( \38324 , \38323 , \1735 );
not \U$37948 ( \38325 , \38323 );
and \U$37949 ( \38326 , \38325 , \1734 );
nor \U$37950 ( \38327 , \38324 , \38326 );
xor \U$37951 ( \38328 , \38320 , \38327 );
and \U$37952 ( \38329 , \558 , RIae75a10_20);
and \U$37953 ( \38330 , RIae75920_18, \556 );
nor \U$37954 ( \38331 , \38329 , \38330 );
and \U$37955 ( \38332 , \38331 , \504 );
not \U$37956 ( \38333 , \38331 );
and \U$37957 ( \38334 , \38333 , \562 );
nor \U$37958 ( \38335 , \38332 , \38334 );
not \U$37959 ( \38336 , \400 );
and \U$37960 ( \38337 , \436 , RIae78800_118);
and \U$37961 ( \38338 , RIae78710_116, \434 );
nor \U$37962 ( \38339 , \38337 , \38338 );
not \U$37963 ( \38340 , \38339 );
or \U$37964 ( \38341 , \38336 , \38340 );
or \U$37965 ( \38342 , \38339 , \400 );
nand \U$37966 ( \38343 , \38341 , \38342 );
xor \U$37967 ( \38344 , \38335 , \38343 );
not \U$37968 ( \38345 , \471 );
and \U$37969 ( \38346 , \514 , RIae75bf0_24);
and \U$37970 ( \38347 , RIae75b00_22, \512 );
nor \U$37971 ( \38348 , \38346 , \38347 );
not \U$37972 ( \38349 , \38348 );
or \U$37973 ( \38350 , \38345 , \38349 );
or \U$37974 ( \38351 , \38348 , \469 );
nand \U$37975 ( \38352 , \38350 , \38351 );
xor \U$37976 ( \38353 , \38344 , \38352 );
not \U$37977 ( \38354 , \787 );
and \U$37978 ( \38355 , \883 , RIae75ce0_26);
and \U$37979 ( \38356 , RIae75dd0_28, \881 );
nor \U$37980 ( \38357 , \38355 , \38356 );
not \U$37981 ( \38358 , \38357 );
or \U$37982 ( \38359 , \38354 , \38358 );
or \U$37983 ( \38360 , \38357 , \789 );
nand \U$37984 ( \38361 , \38359 , \38360 );
and \U$37985 ( \38362 , \672 , RIae75fb0_32);
and \U$37986 ( \38363 , RIae75ec0_30, \670 );
nor \U$37987 ( \38364 , \38362 , \38363 );
and \U$37988 ( \38365 , \38364 , \588 );
not \U$37989 ( \38366 , \38364 );
and \U$37990 ( \38367 , \38366 , \587 );
nor \U$37991 ( \38368 , \38365 , \38367 );
xor \U$37992 ( \38369 , \38361 , \38368 );
and \U$37993 ( \38370 , \1138 , RIae75650_12);
and \U$37994 ( \38371 , RIae75560_10, \1136 );
nor \U$37995 ( \38372 , \38370 , \38371 );
and \U$37996 ( \38373 , \38372 , \1012 );
not \U$37997 ( \38374 , \38372 );
and \U$37998 ( \38375 , \38374 , \1142 );
nor \U$37999 ( \38376 , \38373 , \38375 );
xor \U$38000 ( \38377 , \38369 , \38376 );
xor \U$38001 ( \38378 , \38353 , \38377 );
xor \U$38002 ( \38379 , \38328 , \38378 );
xor \U$38003 ( \38380 , \38305 , \38379 );
xor \U$38004 ( \38381 , \38293 , \38380 );
xor \U$38005 ( \38382 , \38279 , \38381 );
xor \U$38006 ( \38383 , \38265 , \38382 );
xor \U$38007 ( \38384 , \38188 , \38383 );
xor \U$38008 ( \38385 , \38174 , \38384 );
xor \U$38009 ( \38386 , \37685 , \37692 );
xor \U$38010 ( \38387 , \38386 , \37700 );
and \U$38011 ( \38388 , \37722 , \38387 );
xor \U$38012 ( \38389 , \37685 , \37692 );
xor \U$38013 ( \38390 , \38389 , \37700 );
and \U$38014 ( \38391 , \37747 , \38390 );
and \U$38015 ( \38392 , \37722 , \37747 );
or \U$38016 ( \38393 , \38388 , \38391 , \38392 );
xor \U$38017 ( \38394 , \37939 , \37946 );
xor \U$38018 ( \38395 , \38394 , \37954 );
xor \U$38019 ( \38396 , \38393 , \38395 );
xor \U$38020 ( \38397 , \37340 , \37347 );
xor \U$38021 ( \38398 , \38397 , \37355 );
and \U$38022 ( \38399 , \37380 , \38398 );
xor \U$38023 ( \38400 , \37340 , \37347 );
xor \U$38024 ( \38401 , \38400 , \37355 );
and \U$38025 ( \38402 , \37404 , \38401 );
and \U$38026 ( \38403 , \37380 , \37404 );
or \U$38027 ( \38404 , \38399 , \38402 , \38403 );
and \U$38028 ( \38405 , \38396 , \38404 );
and \U$38029 ( \38406 , \38393 , \38395 );
or \U$38030 ( \38407 , \38405 , \38406 );
xor \U$38031 ( \38408 , \37656 , \37664 );
and \U$38032 ( \38409 , \38408 , \37673 );
and \U$38033 ( \38410 , \37656 , \37664 );
or \U$38034 ( \38411 , \38409 , \38410 );
and \U$38035 ( \38412 , \5896 , RIae76be0_58);
and \U$38036 ( \38413 , RIae78ad0_124, \5894 );
nor \U$38037 ( \38414 , \38412 , \38413 );
and \U$38038 ( \38415 , \38414 , \5590 );
not \U$38039 ( \38416 , \38414 );
and \U$38040 ( \38417 , \38416 , \5589 );
nor \U$38041 ( \38418 , \38415 , \38417 );
xor \U$38042 ( \38419 , \38418 , \6314 );
and \U$38043 ( \38420 , \6172 , RIae78d28_129);
and \U$38044 ( \38421 , RIae78e18_131, \6170 );
nor \U$38045 ( \38422 , \38420 , \38421 );
and \U$38046 ( \38423 , \38422 , \6176 );
not \U$38047 ( \38424 , \38422 );
and \U$38048 ( \38425 , \38424 , \6175 );
nor \U$38049 ( \38426 , \38423 , \38425 );
and \U$38050 ( \38427 , \38419 , \38426 );
and \U$38051 ( \38428 , \38418 , \6314 );
or \U$38052 ( \38429 , \38427 , \38428 );
xor \U$38053 ( \38430 , \38411 , \38429 );
xor \U$38054 ( \38431 , \37630 , \37637 );
and \U$38055 ( \38432 , \38431 , \37645 );
and \U$38056 ( \38433 , \37630 , \37637 );
or \U$38057 ( \38434 , \38432 , \38433 );
and \U$38058 ( \38435 , \38430 , \38434 );
and \U$38059 ( \38436 , \38411 , \38429 );
or \U$38060 ( \38437 , \38435 , \38436 );
xor \U$38061 ( \38438 , \38437 , \37253 );
xor \U$38062 ( \38439 , \37279 , \37305 );
and \U$38063 ( \38440 , \38439 , \37331 );
and \U$38064 ( \38441 , \37279 , \37305 );
or \U$38065 ( \38442 , \38440 , \38441 );
and \U$38066 ( \38443 , \38438 , \38442 );
and \U$38067 ( \38444 , \38437 , \37253 );
or \U$38068 ( \38445 , \38443 , \38444 );
xor \U$38069 ( \38446 , \38407 , \38445 );
xor \U$38070 ( \38447 , \37808 , \37814 );
xor \U$38071 ( \38448 , \38447 , \37835 );
and \U$38072 ( \38449 , \37852 , \38448 );
xor \U$38073 ( \38450 , \37808 , \37814 );
xor \U$38074 ( \38451 , \38450 , \37835 );
and \U$38075 ( \38452 , \37926 , \38451 );
and \U$38076 ( \38453 , \37852 , \37926 );
or \U$38077 ( \38454 , \38449 , \38452 , \38453 );
and \U$38078 ( \38455 , \38446 , \38454 );
and \U$38079 ( \38456 , \38407 , \38445 );
or \U$38080 ( \38457 , \38455 , \38456 );
xor \U$38081 ( \38458 , \37971 , \37975 );
and \U$38082 ( \38459 , \38458 , \37980 );
and \U$38083 ( \38460 , \37971 , \37975 );
or \U$38084 ( \38461 , \38459 , \38460 );
xor \U$38085 ( \38462 , \37957 , \37961 );
and \U$38086 ( \38463 , \38462 , \37966 );
and \U$38087 ( \38464 , \37957 , \37961 );
or \U$38088 ( \38465 , \38463 , \38464 );
xor \U$38089 ( \38466 , \38461 , \38465 );
xor \U$38090 ( \38467 , \37986 , \37998 );
and \U$38091 ( \38468 , \38467 , \38024 );
and \U$38092 ( \38469 , \37986 , \37998 );
or \U$38093 ( \38470 , \38468 , \38469 );
xor \U$38094 ( \38471 , \38466 , \38470 );
xor \U$38095 ( \38472 , \38457 , \38471 );
xor \U$38096 ( \38473 , \37967 , \37981 );
xor \U$38097 ( \38474 , \38473 , \38025 );
and \U$38098 ( \38475 , \38040 , \38474 );
xor \U$38099 ( \38476 , \37967 , \37981 );
xor \U$38100 ( \38477 , \38476 , \38025 );
and \U$38101 ( \38478 , \38169 , \38477 );
and \U$38102 ( \38479 , \38040 , \38169 );
or \U$38103 ( \38480 , \38475 , \38478 , \38479 );
xor \U$38104 ( \38481 , \38472 , \38480 );
xor \U$38105 ( \38482 , \38385 , \38481 );
xor \U$38106 ( \38483 , \38437 , \37253 );
xor \U$38107 ( \38484 , \38483 , \38442 );
xor \U$38108 ( \38485 , \37769 , \37783 );
xor \U$38109 ( \38486 , \38485 , \37928 );
and \U$38110 ( \38487 , \38484 , \38486 );
xor \U$38111 ( \38488 , \37411 , \37610 );
xor \U$38112 ( \38489 , \38488 , \37752 );
xor \U$38113 ( \38490 , \37769 , \37783 );
xor \U$38114 ( \38491 , \38490 , \37928 );
and \U$38115 ( \38492 , \38489 , \38491 );
and \U$38116 ( \38493 , \38484 , \38489 );
or \U$38117 ( \38494 , \38487 , \38492 , \38493 );
xor \U$38118 ( \38495 , \38407 , \38445 );
xor \U$38119 ( \38496 , \38495 , \38454 );
xor \U$38120 ( \38497 , \38494 , \38496 );
xor \U$38121 ( \38498 , \37586 , \37593 );
xor \U$38122 ( \38499 , \38498 , \37601 );
xor \U$38123 ( \38500 , \37534 , \37541 );
xor \U$38124 ( \38501 , \38500 , \37549 );
and \U$38125 ( \38502 , \38499 , \38501 );
xor \U$38126 ( \38503 , \37559 , \37566 );
xor \U$38127 ( \38504 , \38503 , \37574 );
xor \U$38128 ( \38505 , \37534 , \37541 );
xor \U$38129 ( \38506 , \38505 , \37549 );
and \U$38130 ( \38507 , \38504 , \38506 );
and \U$38131 ( \38508 , \38499 , \38504 );
or \U$38132 ( \38509 , \38502 , \38507 , \38508 );
xor \U$38133 ( \38510 , \38418 , \6314 );
xor \U$38134 ( \38511 , \38510 , \38426 );
xor \U$38135 ( \38512 , \38509 , \38511 );
xor \U$38136 ( \38513 , \37467 , \37475 );
xor \U$38137 ( \38514 , \38513 , \37484 );
xor \U$38138 ( \38515 , \37443 , \37448 );
xor \U$38139 ( \38516 , \38515 , \37456 );
and \U$38140 ( \38517 , \38514 , \38516 );
xor \U$38141 ( \38518 , \37418 , \37425 );
xor \U$38142 ( \38519 , \38518 , \37433 );
xor \U$38143 ( \38520 , \37443 , \37448 );
xor \U$38144 ( \38521 , \38520 , \37456 );
and \U$38145 ( \38522 , \38519 , \38521 );
and \U$38146 ( \38523 , \38514 , \38519 );
or \U$38147 ( \38524 , \38517 , \38522 , \38523 );
and \U$38148 ( \38525 , \38512 , \38524 );
and \U$38149 ( \38526 , \38509 , \38511 );
or \U$38150 ( \38527 , \38525 , \38526 );
and \U$38151 ( \38528 , \5399 , RIae76af0_56);
and \U$38152 ( \38529 , RIae76a00_54, \5397 );
nor \U$38153 ( \38530 , \38528 , \38529 );
and \U$38154 ( \38531 , \38530 , \5016 );
not \U$38155 ( \38532 , \38530 );
and \U$38156 ( \38533 , \38532 , \5403 );
nor \U$38157 ( \38534 , \38531 , \38533 );
and \U$38158 ( \38535 , \4688 , RIae76370_40);
and \U$38159 ( \38536 , RIae76280_38, \4686 );
nor \U$38160 ( \38537 , \38535 , \38536 );
and \U$38161 ( \38538 , \38537 , \4481 );
not \U$38162 ( \38539 , \38537 );
and \U$38163 ( \38540 , \38539 , \4482 );
nor \U$38164 ( \38541 , \38538 , \38540 );
xor \U$38165 ( \38542 , \38534 , \38541 );
and \U$38166 ( \38543 , \5896 , RIae76820_50);
and \U$38167 ( \38544 , RIae76910_52, \5894 );
nor \U$38168 ( \38545 , \38543 , \38544 );
and \U$38169 ( \38546 , \38545 , \5590 );
not \U$38170 ( \38547 , \38545 );
and \U$38171 ( \38548 , \38547 , \5589 );
nor \U$38172 ( \38549 , \38546 , \38548 );
and \U$38173 ( \38550 , \38542 , \38549 );
and \U$38174 ( \38551 , \38534 , \38541 );
or \U$38175 ( \38552 , \38550 , \38551 );
and \U$38176 ( \38553 , \6941 , RIae78d28_129);
and \U$38177 ( \38554 , RIae78e18_131, \6939 );
nor \U$38178 ( \38555 , \38553 , \38554 );
and \U$38179 ( \38556 , \38555 , \6314 );
not \U$38180 ( \38557 , \38555 );
and \U$38181 ( \38558 , \38557 , \6945 );
nor \U$38182 ( \38559 , \38556 , \38558 );
xor \U$38183 ( \38560 , \38559 , \7206 );
and \U$38184 ( \38561 , \6172 , RIae76be0_58);
and \U$38185 ( \38562 , RIae78ad0_124, \6170 );
nor \U$38186 ( \38563 , \38561 , \38562 );
and \U$38187 ( \38564 , \38563 , \6176 );
not \U$38188 ( \38565 , \38563 );
and \U$38189 ( \38566 , \38565 , \6175 );
nor \U$38190 ( \38567 , \38564 , \38566 );
and \U$38191 ( \38568 , \38560 , \38567 );
and \U$38192 ( \38569 , \38559 , \7206 );
or \U$38193 ( \38570 , \38568 , \38569 );
xor \U$38194 ( \38571 , \38552 , \38570 );
and \U$38195 ( \38572 , \4247 , RIae76190_36);
and \U$38196 ( \38573 , RIae760a0_34, \4245 );
nor \U$38197 ( \38574 , \38572 , \38573 );
and \U$38198 ( \38575 , \38574 , \3989 );
not \U$38199 ( \38576 , \38574 );
and \U$38200 ( \38577 , \38576 , \4251 );
nor \U$38201 ( \38578 , \38575 , \38577 );
not \U$38202 ( \38579 , \2774 );
and \U$38203 ( \38580 , \3214 , RIae76460_42);
and \U$38204 ( \38581 , RIae76550_44, \3212 );
nor \U$38205 ( \38582 , \38580 , \38581 );
not \U$38206 ( \38583 , \38582 );
or \U$38207 ( \38584 , \38579 , \38583 );
or \U$38208 ( \38585 , \38582 , \3218 );
nand \U$38209 ( \38586 , \38584 , \38585 );
xor \U$38210 ( \38587 , \38578 , \38586 );
and \U$38211 ( \38588 , \3730 , RIae76730_48);
and \U$38212 ( \38589 , RIae76640_46, \3728 );
nor \U$38213 ( \38590 , \38588 , \38589 );
and \U$38214 ( \38591 , \38590 , \3732 );
not \U$38215 ( \38592 , \38590 );
and \U$38216 ( \38593 , \38592 , \3422 );
nor \U$38217 ( \38594 , \38591 , \38593 );
and \U$38218 ( \38595 , \38587 , \38594 );
and \U$38219 ( \38596 , \38578 , \38586 );
or \U$38220 ( \38597 , \38595 , \38596 );
and \U$38221 ( \38598 , \38571 , \38597 );
and \U$38222 ( \38599 , \38552 , \38570 );
or \U$38223 ( \38600 , \38598 , \38599 );
not \U$38224 ( \38601 , \400 );
and \U$38225 ( \38602 , \436 , RIae77cc0_94);
and \U$38226 ( \38603 , RIae77bd0_92, \434 );
nor \U$38227 ( \38604 , \38602 , \38603 );
not \U$38228 ( \38605 , \38604 );
or \U$38229 ( \38606 , \38601 , \38605 );
or \U$38230 ( \38607 , \38604 , \402 );
nand \U$38231 ( \38608 , \38606 , \38607 );
not \U$38232 ( \38609 , \469 );
and \U$38233 ( \38610 , \514 , RIae77db0_96);
and \U$38234 ( \38611 , RIae77ea0_98, \512 );
nor \U$38235 ( \38612 , \38610 , \38611 );
not \U$38236 ( \38613 , \38612 );
or \U$38237 ( \38614 , \38609 , \38613 );
or \U$38238 ( \38615 , \38612 , \471 );
nand \U$38239 ( \38616 , \38614 , \38615 );
xor \U$38240 ( \38617 , \38608 , \38616 );
and \U$38241 ( \38618 , \558 , RIae789e0_122);
and \U$38242 ( \38619 , RIae788f0_120, \556 );
nor \U$38243 ( \38620 , \38618 , \38619 );
and \U$38244 ( \38621 , \38620 , \504 );
not \U$38245 ( \38622 , \38620 );
and \U$38246 ( \38623 , \38622 , \562 );
nor \U$38247 ( \38624 , \38621 , \38623 );
and \U$38248 ( \38625 , \38617 , \38624 );
and \U$38249 ( \38626 , \38608 , \38616 );
or \U$38250 ( \38627 , \38625 , \38626 );
xor \U$38251 ( \38628 , \38627 , \37491 );
xor \U$38252 ( \38629 , \37503 , \37511 );
xor \U$38253 ( \38630 , \38629 , \37520 );
and \U$38254 ( \38631 , \38628 , \38630 );
and \U$38255 ( \38632 , \38627 , \37491 );
or \U$38256 ( \38633 , \38631 , \38632 );
xor \U$38257 ( \38634 , \38600 , \38633 );
and \U$38258 ( \38635 , \1939 , RIae75650_12);
and \U$38259 ( \38636 , RIae75560_10, \1937 );
nor \U$38260 ( \38637 , \38635 , \38636 );
and \U$38261 ( \38638 , \38637 , \1735 );
not \U$38262 ( \38639 , \38637 );
and \U$38263 ( \38640 , \38639 , \1734 );
nor \U$38264 ( \38641 , \38638 , \38640 );
and \U$38265 ( \38642 , \1376 , RIae75fb0_32);
and \U$38266 ( \38643 , RIae75ec0_30, \1374 );
nor \U$38267 ( \38644 , \38642 , \38643 );
and \U$38268 ( \38645 , \38644 , \1380 );
not \U$38269 ( \38646 , \38644 );
and \U$38270 ( \38647 , \38646 , \1261 );
nor \U$38271 ( \38648 , \38645 , \38647 );
xor \U$38272 ( \38649 , \38641 , \38648 );
and \U$38273 ( \38650 , \1593 , RIae75ce0_26);
and \U$38274 ( \38651 , RIae75dd0_28, \1591 );
nor \U$38275 ( \38652 , \38650 , \38651 );
and \U$38276 ( \38653 , \38652 , \1498 );
not \U$38277 ( \38654 , \38652 );
and \U$38278 ( \38655 , \38654 , \1488 );
nor \U$38279 ( \38656 , \38653 , \38655 );
and \U$38280 ( \38657 , \38649 , \38656 );
and \U$38281 ( \38658 , \38641 , \38648 );
or \U$38282 ( \38659 , \38657 , \38658 );
and \U$38283 ( \38660 , \1138 , RIae75a10_20);
and \U$38284 ( \38661 , RIae75920_18, \1136 );
nor \U$38285 ( \38662 , \38660 , \38661 );
and \U$38286 ( \38663 , \38662 , \1012 );
not \U$38287 ( \38664 , \38662 );
and \U$38288 ( \38665 , \38664 , \1142 );
nor \U$38289 ( \38666 , \38663 , \38665 );
and \U$38290 ( \38667 , \672 , RIae78800_118);
and \U$38291 ( \38668 , RIae78710_116, \670 );
nor \U$38292 ( \38669 , \38667 , \38668 );
and \U$38293 ( \38670 , \38669 , \588 );
not \U$38294 ( \38671 , \38669 );
and \U$38295 ( \38672 , \38671 , \587 );
nor \U$38296 ( \38673 , \38670 , \38672 );
xor \U$38297 ( \38674 , \38666 , \38673 );
not \U$38298 ( \38675 , \787 );
and \U$38299 ( \38676 , \883 , RIae75bf0_24);
and \U$38300 ( \38677 , RIae75b00_22, \881 );
nor \U$38301 ( \38678 , \38676 , \38677 );
not \U$38302 ( \38679 , \38678 );
or \U$38303 ( \38680 , \38675 , \38679 );
or \U$38304 ( \38681 , \38678 , \789 );
nand \U$38305 ( \38682 , \38680 , \38681 );
and \U$38306 ( \38683 , \38674 , \38682 );
and \U$38307 ( \38684 , \38666 , \38673 );
or \U$38308 ( \38685 , \38683 , \38684 );
xor \U$38309 ( \38686 , \38659 , \38685 );
and \U$38310 ( \38687 , \2224 , RIae75830_16);
and \U$38311 ( \38688 , RIae75740_14, \2222 );
nor \U$38312 ( \38689 , \38687 , \38688 );
and \U$38313 ( \38690 , \38689 , \2061 );
not \U$38314 ( \38691 , \38689 );
and \U$38315 ( \38692 , \38691 , \2060 );
nor \U$38316 ( \38693 , \38690 , \38692 );
and \U$38317 ( \38694 , \2607 , RIae75290_4);
and \U$38318 ( \38695 , RIae751a0_2, \2605 );
nor \U$38319 ( \38696 , \38694 , \38695 );
and \U$38320 ( \38697 , \38696 , \2611 );
not \U$38321 ( \38698 , \38696 );
and \U$38322 ( \38699 , \38698 , \2397 );
nor \U$38323 ( \38700 , \38697 , \38699 );
xor \U$38324 ( \38701 , \38693 , \38700 );
not \U$38325 ( \38702 , \2789 );
and \U$38326 ( \38703 , \2783 , RIae75380_6);
and \U$38327 ( \38704 , RIae75470_8, \2781 );
nor \U$38328 ( \38705 , \38703 , \38704 );
not \U$38329 ( \38706 , \38705 );
or \U$38330 ( \38707 , \38702 , \38706 );
or \U$38331 ( \38708 , \38705 , \3089 );
nand \U$38332 ( \38709 , \38707 , \38708 );
and \U$38333 ( \38710 , \38701 , \38709 );
and \U$38334 ( \38711 , \38693 , \38700 );
or \U$38335 ( \38712 , \38710 , \38711 );
and \U$38336 ( \38713 , \38686 , \38712 );
and \U$38337 ( \38714 , \38659 , \38685 );
or \U$38338 ( \38715 , \38713 , \38714 );
and \U$38339 ( \38716 , \38634 , \38715 );
and \U$38340 ( \38717 , \38600 , \38633 );
or \U$38341 ( \38718 , \38716 , \38717 );
xor \U$38342 ( \38719 , \38527 , \38718 );
xor \U$38343 ( \38720 , \37492 , \37494 );
xor \U$38344 ( \38721 , \38720 , \37523 );
xor \U$38345 ( \38722 , \37646 , \37648 );
xor \U$38346 ( \38723 , \38722 , \37674 );
and \U$38347 ( \38724 , \38721 , \38723 );
xor \U$38348 ( \38725 , \37286 , \37293 );
xor \U$38349 ( \38726 , \38725 , \37302 );
xor \U$38350 ( \38727 , \37613 , \37618 );
xor \U$38351 ( \38728 , \38726 , \38727 );
xor \U$38352 ( \38729 , \37646 , \37648 );
xor \U$38353 ( \38730 , \38729 , \37674 );
and \U$38354 ( \38731 , \38728 , \38730 );
and \U$38355 ( \38732 , \38721 , \38728 );
or \U$38356 ( \38733 , \38724 , \38731 , \38732 );
and \U$38357 ( \38734 , \38719 , \38733 );
and \U$38358 ( \38735 , \38527 , \38718 );
or \U$38359 ( \38736 , \38734 , \38735 );
xor \U$38360 ( \38737 , \38393 , \38395 );
xor \U$38361 ( \38738 , \38737 , \38404 );
xor \U$38362 ( \38739 , \38736 , \38738 );
xor \U$38363 ( \38740 , \38411 , \38429 );
xor \U$38364 ( \38741 , \38740 , \38434 );
xor \U$38365 ( \38742 , \37623 , \37677 );
xor \U$38366 ( \38743 , \38742 , \37749 );
and \U$38367 ( \38744 , \38741 , \38743 );
xor \U$38368 ( \38745 , \37279 , \37305 );
xor \U$38369 ( \38746 , \38745 , \37331 );
xor \U$38370 ( \38747 , \37254 , \37406 );
xor \U$38371 ( \38748 , \38746 , \38747 );
xor \U$38372 ( \38749 , \37623 , \37677 );
xor \U$38373 ( \38750 , \38749 , \37749 );
and \U$38374 ( \38751 , \38748 , \38750 );
and \U$38375 ( \38752 , \38741 , \38748 );
or \U$38376 ( \38753 , \38744 , \38751 , \38752 );
and \U$38377 ( \38754 , \38739 , \38753 );
and \U$38378 ( \38755 , \38736 , \38738 );
or \U$38379 ( \38756 , \38754 , \38755 );
and \U$38380 ( \38757 , \38497 , \38756 );
and \U$38381 ( \38758 , \38494 , \38496 );
or \U$38382 ( \38759 , \38757 , \38758 );
xor \U$38383 ( \38760 , \37755 , \37931 );
xor \U$38384 ( \38761 , \38760 , \38171 );
not \U$38385 ( \38762 , \38761 );
xor \U$38386 ( \38763 , \38494 , \38496 );
xor \U$38387 ( \38764 , \38763 , \38756 );
not \U$38388 ( \38765 , \38764 );
or \U$38389 ( \38766 , \38762 , \38765 );
or \U$38390 ( \38767 , \38764 , \38761 );
xor \U$38391 ( \38768 , \38641 , \38648 );
xor \U$38392 ( \38769 , \38768 , \38656 );
xor \U$38393 ( \38770 , \38578 , \38586 );
xor \U$38394 ( \38771 , \38770 , \38594 );
and \U$38395 ( \38772 , \38769 , \38771 );
xor \U$38396 ( \38773 , \38693 , \38700 );
xor \U$38397 ( \38774 , \38773 , \38709 );
xor \U$38398 ( \38775 , \38578 , \38586 );
xor \U$38399 ( \38776 , \38775 , \38594 );
and \U$38400 ( \38777 , \38774 , \38776 );
and \U$38401 ( \38778 , \38769 , \38774 );
or \U$38402 ( \38779 , \38772 , \38777 , \38778 );
xor \U$38403 ( \38780 , \38608 , \38616 );
xor \U$38404 ( \38781 , \38780 , \38624 );
not \U$38405 ( \38782 , RIae78620_114);
nor \U$38406 ( \38783 , \38782 , \491 );
xor \U$38407 ( \38784 , \38781 , \38783 );
xor \U$38408 ( \38785 , \38666 , \38673 );
xor \U$38409 ( \38786 , \38785 , \38682 );
and \U$38410 ( \38787 , \38784 , \38786 );
and \U$38411 ( \38788 , \38781 , \38783 );
or \U$38412 ( \38789 , \38787 , \38788 );
xor \U$38413 ( \38790 , \38779 , \38789 );
xor \U$38414 ( \38791 , \37443 , \37448 );
xor \U$38415 ( \38792 , \38791 , \37456 );
xor \U$38416 ( \38793 , \38514 , \38519 );
xor \U$38417 ( \38794 , \38792 , \38793 );
and \U$38418 ( \38795 , \38790 , \38794 );
and \U$38419 ( \38796 , \38779 , \38789 );
or \U$38420 ( \38797 , \38795 , \38796 );
and \U$38421 ( \38798 , \2607 , RIae75740_14);
and \U$38422 ( \38799 , RIae75290_4, \2605 );
nor \U$38423 ( \38800 , \38798 , \38799 );
and \U$38424 ( \38801 , \38800 , \2611 );
not \U$38425 ( \38802 , \38800 );
and \U$38426 ( \38803 , \38802 , \2397 );
nor \U$38427 ( \38804 , \38801 , \38803 );
and \U$38428 ( \38805 , \2224 , RIae75560_10);
and \U$38429 ( \38806 , RIae75830_16, \2222 );
nor \U$38430 ( \38807 , \38805 , \38806 );
and \U$38431 ( \38808 , \38807 , \2061 );
not \U$38432 ( \38809 , \38807 );
and \U$38433 ( \38810 , \38809 , \2060 );
nor \U$38434 ( \38811 , \38808 , \38810 );
xor \U$38435 ( \38812 , \38804 , \38811 );
not \U$38436 ( \38813 , \2789 );
and \U$38437 ( \38814 , \2783 , RIae751a0_2);
and \U$38438 ( \38815 , RIae75380_6, \2781 );
nor \U$38439 ( \38816 , \38814 , \38815 );
not \U$38440 ( \38817 , \38816 );
or \U$38441 ( \38818 , \38813 , \38817 );
or \U$38442 ( \38819 , \38816 , \3089 );
nand \U$38443 ( \38820 , \38818 , \38819 );
and \U$38444 ( \38821 , \38812 , \38820 );
and \U$38445 ( \38822 , \38804 , \38811 );
or \U$38446 ( \38823 , \38821 , \38822 );
and \U$38447 ( \38824 , \1593 , RIae75ec0_30);
and \U$38448 ( \38825 , RIae75ce0_26, \1591 );
nor \U$38449 ( \38826 , \38824 , \38825 );
and \U$38450 ( \38827 , \38826 , \1498 );
not \U$38451 ( \38828 , \38826 );
and \U$38452 ( \38829 , \38828 , \1488 );
nor \U$38453 ( \38830 , \38827 , \38829 );
and \U$38454 ( \38831 , \1376 , RIae75920_18);
and \U$38455 ( \38832 , RIae75fb0_32, \1374 );
nor \U$38456 ( \38833 , \38831 , \38832 );
and \U$38457 ( \38834 , \38833 , \1380 );
not \U$38458 ( \38835 , \38833 );
and \U$38459 ( \38836 , \38835 , \1261 );
nor \U$38460 ( \38837 , \38834 , \38836 );
xor \U$38461 ( \38838 , \38830 , \38837 );
and \U$38462 ( \38839 , \1939 , RIae75dd0_28);
and \U$38463 ( \38840 , RIae75650_12, \1937 );
nor \U$38464 ( \38841 , \38839 , \38840 );
and \U$38465 ( \38842 , \38841 , \1735 );
not \U$38466 ( \38843 , \38841 );
and \U$38467 ( \38844 , \38843 , \1734 );
nor \U$38468 ( \38845 , \38842 , \38844 );
and \U$38469 ( \38846 , \38838 , \38845 );
and \U$38470 ( \38847 , \38830 , \38837 );
or \U$38471 ( \38848 , \38846 , \38847 );
xor \U$38472 ( \38849 , \38823 , \38848 );
and \U$38473 ( \38850 , \1138 , RIae75b00_22);
and \U$38474 ( \38851 , RIae75a10_20, \1136 );
nor \U$38475 ( \38852 , \38850 , \38851 );
and \U$38476 ( \38853 , \38852 , \1012 );
not \U$38477 ( \38854 , \38852 );
and \U$38478 ( \38855 , \38854 , \1142 );
nor \U$38479 ( \38856 , \38853 , \38855 );
and \U$38480 ( \38857 , \672 , RIae788f0_120);
and \U$38481 ( \38858 , RIae78800_118, \670 );
nor \U$38482 ( \38859 , \38857 , \38858 );
and \U$38483 ( \38860 , \38859 , \588 );
not \U$38484 ( \38861 , \38859 );
and \U$38485 ( \38862 , \38861 , \587 );
nor \U$38486 ( \38863 , \38860 , \38862 );
xor \U$38487 ( \38864 , \38856 , \38863 );
not \U$38488 ( \38865 , \789 );
and \U$38489 ( \38866 , \883 , RIae78710_116);
and \U$38490 ( \38867 , RIae75bf0_24, \881 );
nor \U$38491 ( \38868 , \38866 , \38867 );
not \U$38492 ( \38869 , \38868 );
or \U$38493 ( \38870 , \38865 , \38869 );
or \U$38494 ( \38871 , \38868 , \789 );
nand \U$38495 ( \38872 , \38870 , \38871 );
and \U$38496 ( \38873 , \38864 , \38872 );
and \U$38497 ( \38874 , \38856 , \38863 );
or \U$38498 ( \38875 , \38873 , \38874 );
and \U$38499 ( \38876 , \38849 , \38875 );
and \U$38500 ( \38877 , \38823 , \38848 );
or \U$38501 ( \38878 , \38876 , \38877 );
nand \U$38502 ( \38879 , RIae78260_106, RIae78b48_125);
and \U$38503 ( \38880 , \384 , RIae78620_114);
and \U$38504 ( \38881 , RIae78440_110, \382 );
nor \U$38505 ( \38882 , \38880 , \38881 );
not \U$38506 ( \38883 , \38882 );
not \U$38507 ( \38884 , \392 );
and \U$38508 ( \38885 , \38883 , \38884 );
and \U$38509 ( \38886 , \38882 , \392 );
nor \U$38510 ( \38887 , \38885 , \38886 );
nand \U$38511 ( \38888 , \38879 , \38887 );
not \U$38512 ( \38889 , \392 );
and \U$38513 ( \38890 , \384 , RIae78440_110);
and \U$38514 ( \38891 , RIae784b8_111, \382 );
nor \U$38515 ( \38892 , \38890 , \38891 );
not \U$38516 ( \38893 , \38892 );
or \U$38517 ( \38894 , \38889 , \38893 );
or \U$38518 ( \38895 , \38892 , \388 );
nand \U$38519 ( \38896 , \38894 , \38895 );
xor \U$38520 ( \38897 , \38888 , \38896 );
not \U$38521 ( \38898 , \402 );
and \U$38522 ( \38899 , \436 , RIae784b8_111);
and \U$38523 ( \38900 , RIae77cc0_94, \434 );
nor \U$38524 ( \38901 , \38899 , \38900 );
not \U$38525 ( \38902 , \38901 );
or \U$38526 ( \38903 , \38898 , \38902 );
or \U$38527 ( \38904 , \38901 , \402 );
nand \U$38528 ( \38905 , \38903 , \38904 );
not \U$38529 ( \38906 , \471 );
and \U$38530 ( \38907 , \514 , RIae77bd0_92);
and \U$38531 ( \38908 , RIae77db0_96, \512 );
nor \U$38532 ( \38909 , \38907 , \38908 );
not \U$38533 ( \38910 , \38909 );
or \U$38534 ( \38911 , \38906 , \38910 );
or \U$38535 ( \38912 , \38909 , \471 );
nand \U$38536 ( \38913 , \38911 , \38912 );
xor \U$38537 ( \38914 , \38905 , \38913 );
and \U$38538 ( \38915 , \558 , RIae77ea0_98);
and \U$38539 ( \38916 , RIae789e0_122, \556 );
nor \U$38540 ( \38917 , \38915 , \38916 );
and \U$38541 ( \38918 , \38917 , \504 );
not \U$38542 ( \38919 , \38917 );
and \U$38543 ( \38920 , \38919 , \562 );
nor \U$38544 ( \38921 , \38918 , \38920 );
and \U$38545 ( \38922 , \38914 , \38921 );
and \U$38546 ( \38923 , \38905 , \38913 );
or \U$38547 ( \38924 , \38922 , \38923 );
and \U$38548 ( \38925 , \38897 , \38924 );
and \U$38549 ( \38926 , \38888 , \38896 );
or \U$38550 ( \38927 , \38925 , \38926 );
xor \U$38551 ( \38928 , \38878 , \38927 );
not \U$38552 ( \38929 , \2774 );
and \U$38553 ( \38930 , \3214 , RIae75470_8);
and \U$38554 ( \38931 , RIae76460_42, \3212 );
nor \U$38555 ( \38932 , \38930 , \38931 );
not \U$38556 ( \38933 , \38932 );
or \U$38557 ( \38934 , \38929 , \38933 );
or \U$38558 ( \38935 , \38932 , \2774 );
nand \U$38559 ( \38936 , \38934 , \38935 );
and \U$38560 ( \38937 , \3730 , RIae76550_44);
and \U$38561 ( \38938 , RIae76730_48, \3728 );
nor \U$38562 ( \38939 , \38937 , \38938 );
and \U$38563 ( \38940 , \38939 , \3732 );
not \U$38564 ( \38941 , \38939 );
and \U$38565 ( \38942 , \38941 , \3422 );
nor \U$38566 ( \38943 , \38940 , \38942 );
xor \U$38567 ( \38944 , \38936 , \38943 );
and \U$38568 ( \38945 , \4247 , RIae76640_46);
and \U$38569 ( \38946 , RIae76190_36, \4245 );
nor \U$38570 ( \38947 , \38945 , \38946 );
and \U$38571 ( \38948 , \38947 , \3989 );
not \U$38572 ( \38949 , \38947 );
and \U$38573 ( \38950 , \38949 , \4251 );
nor \U$38574 ( \38951 , \38948 , \38950 );
and \U$38575 ( \38952 , \38944 , \38951 );
and \U$38576 ( \38953 , \38936 , \38943 );
or \U$38577 ( \38954 , \38952 , \38953 );
and \U$38578 ( \38955 , \6172 , RIae76910_52);
and \U$38579 ( \38956 , RIae76be0_58, \6170 );
nor \U$38580 ( \38957 , \38955 , \38956 );
and \U$38581 ( \38958 , \38957 , \6175 );
not \U$38582 ( \38959 , \38957 );
and \U$38583 ( \38960 , \38959 , \6176 );
nor \U$38584 ( \38961 , \38958 , \38960 );
and \U$38585 ( \38962 , \6941 , RIae78ad0_124);
and \U$38586 ( \38963 , RIae78d28_129, \6939 );
nor \U$38587 ( \38964 , \38962 , \38963 );
and \U$38588 ( \38965 , \38964 , \6945 );
not \U$38589 ( \38966 , \38964 );
and \U$38590 ( \38967 , \38966 , \6314 );
nor \U$38591 ( \38968 , \38965 , \38967 );
or \U$38592 ( \38969 , \38961 , \38968 );
not \U$38593 ( \38970 , \38968 );
not \U$38594 ( \38971 , \38961 );
or \U$38595 ( \38972 , \38970 , \38971 );
nand \U$38596 ( \38973 , RIae78e18_131, \7633 );
and \U$38597 ( \38974 , \38973 , \7206 );
not \U$38598 ( \38975 , \38973 );
and \U$38599 ( \38976 , \38975 , \7205 );
nor \U$38600 ( \38977 , \38974 , \38976 );
nand \U$38601 ( \38978 , \38972 , \38977 );
nand \U$38602 ( \38979 , \38969 , \38978 );
xor \U$38603 ( \38980 , \38954 , \38979 );
and \U$38604 ( \38981 , \5896 , RIae76a00_54);
and \U$38605 ( \38982 , RIae76820_50, \5894 );
nor \U$38606 ( \38983 , \38981 , \38982 );
and \U$38607 ( \38984 , \38983 , \5590 );
not \U$38608 ( \38985 , \38983 );
and \U$38609 ( \38986 , \38985 , \5589 );
nor \U$38610 ( \38987 , \38984 , \38986 );
and \U$38611 ( \38988 , \4688 , RIae760a0_34);
and \U$38612 ( \38989 , RIae76370_40, \4686 );
nor \U$38613 ( \38990 , \38988 , \38989 );
and \U$38614 ( \38991 , \38990 , \4481 );
not \U$38615 ( \38992 , \38990 );
and \U$38616 ( \38993 , \38992 , \4482 );
nor \U$38617 ( \38994 , \38991 , \38993 );
xor \U$38618 ( \38995 , \38987 , \38994 );
and \U$38619 ( \38996 , \5399 , RIae76280_38);
and \U$38620 ( \38997 , RIae76af0_56, \5397 );
nor \U$38621 ( \38998 , \38996 , \38997 );
and \U$38622 ( \38999 , \38998 , \5016 );
not \U$38623 ( \39000 , \38998 );
and \U$38624 ( \39001 , \39000 , \5403 );
nor \U$38625 ( \39002 , \38999 , \39001 );
and \U$38626 ( \39003 , \38995 , \39002 );
and \U$38627 ( \39004 , \38987 , \38994 );
or \U$38628 ( \39005 , \39003 , \39004 );
and \U$38629 ( \39006 , \38980 , \39005 );
and \U$38630 ( \39007 , \38954 , \38979 );
or \U$38631 ( \39008 , \39006 , \39007 );
and \U$38632 ( \39009 , \38928 , \39008 );
and \U$38633 ( \39010 , \38878 , \38927 );
or \U$38634 ( \39011 , \39009 , \39010 );
xor \U$38635 ( \39012 , \38797 , \39011 );
xor \U$38636 ( \39013 , \38659 , \38685 );
xor \U$38637 ( \39014 , \39013 , \38712 );
xor \U$38638 ( \39015 , \38627 , \37491 );
xor \U$38639 ( \39016 , \39015 , \38630 );
and \U$38640 ( \39017 , \39014 , \39016 );
xor \U$38641 ( \39018 , \37534 , \37541 );
xor \U$38642 ( \39019 , \39018 , \37549 );
xor \U$38643 ( \39020 , \38499 , \38504 );
xor \U$38644 ( \39021 , \39019 , \39020 );
xor \U$38645 ( \39022 , \38627 , \37491 );
xor \U$38646 ( \39023 , \39022 , \38630 );
and \U$38647 ( \39024 , \39021 , \39023 );
and \U$38648 ( \39025 , \39014 , \39021 );
or \U$38649 ( \39026 , \39017 , \39024 , \39025 );
and \U$38650 ( \39027 , \39012 , \39026 );
and \U$38651 ( \39028 , \38797 , \39011 );
or \U$38652 ( \39029 , \39027 , \39028 );
xor \U$38653 ( \39030 , \37490 , \37526 );
xor \U$38654 ( \39031 , \39030 , \37607 );
xor \U$38655 ( \39032 , \39029 , \39031 );
xor \U$38656 ( \39033 , \37552 , \37577 );
xor \U$38657 ( \39034 , \39033 , \37604 );
xor \U$38658 ( \39035 , \37436 , \37459 );
xor \U$38659 ( \39036 , \39035 , \37487 );
xor \U$38660 ( \39037 , \39034 , \39036 );
xor \U$38661 ( \39038 , \37646 , \37648 );
xor \U$38662 ( \39039 , \39038 , \37674 );
xor \U$38663 ( \39040 , \38721 , \38728 );
xor \U$38664 ( \39041 , \39039 , \39040 );
and \U$38665 ( \39042 , \39037 , \39041 );
and \U$38666 ( \39043 , \39034 , \39036 );
or \U$38667 ( \39044 , \39042 , \39043 );
and \U$38668 ( \39045 , \39032 , \39044 );
and \U$38669 ( \39046 , \39029 , \39031 );
or \U$38670 ( \39047 , \39045 , \39046 );
xor \U$38671 ( \39048 , \38736 , \38738 );
xor \U$38672 ( \39049 , \39048 , \38753 );
and \U$38673 ( \39050 , \39047 , \39049 );
xor \U$38674 ( \39051 , \37769 , \37783 );
xor \U$38675 ( \39052 , \39051 , \37928 );
xor \U$38676 ( \39053 , \38484 , \38489 );
xor \U$38677 ( \39054 , \39052 , \39053 );
xor \U$38678 ( \39055 , \38736 , \38738 );
xor \U$38679 ( \39056 , \39055 , \38753 );
and \U$38680 ( \39057 , \39054 , \39056 );
and \U$38681 ( \39058 , \39047 , \39054 );
or \U$38682 ( \39059 , \39050 , \39057 , \39058 );
nand \U$38683 ( \39060 , \38767 , \39059 );
nand \U$38684 ( \39061 , \38766 , \39060 );
xor \U$38685 ( \39062 , \38759 , \39061 );
xor \U$38686 ( \39063 , \38482 , \39062 );
not \U$38687 ( \39064 , \39063 );
xnor \U$38688 ( \39065 , \38764 , \39059 );
not \U$38689 ( \39066 , \39065 );
not \U$38690 ( \39067 , \38761 );
and \U$38691 ( \39068 , \39066 , \39067 );
and \U$38692 ( \39069 , \39065 , \38761 );
nor \U$38693 ( \39070 , \39068 , \39069 );
not \U$38694 ( \39071 , \39070 );
xor \U$38695 ( \39072 , \38905 , \38913 );
xor \U$38696 ( \39073 , \39072 , \38921 );
xor \U$38697 ( \39074 , \38856 , \38863 );
xor \U$38698 ( \39075 , \39074 , \38872 );
and \U$38699 ( \39076 , \39073 , \39075 );
xor \U$38700 ( \39077 , \38830 , \38837 );
xor \U$38701 ( \39078 , \39077 , \38845 );
xor \U$38702 ( \39079 , \38856 , \38863 );
xor \U$38703 ( \39080 , \39079 , \38872 );
and \U$38704 ( \39081 , \39078 , \39080 );
and \U$38705 ( \39082 , \39073 , \39078 );
or \U$38706 ( \39083 , \39076 , \39081 , \39082 );
xor \U$38707 ( \39084 , \38534 , \38541 );
xor \U$38708 ( \39085 , \39084 , \38549 );
xor \U$38709 ( \39086 , \39083 , \39085 );
xor \U$38710 ( \39087 , \38804 , \38811 );
xor \U$38711 ( \39088 , \39087 , \38820 );
xor \U$38712 ( \39089 , \38936 , \38943 );
xor \U$38713 ( \39090 , \39089 , \38951 );
xor \U$38714 ( \39091 , \39088 , \39090 );
xor \U$38715 ( \39092 , \38987 , \38994 );
xor \U$38716 ( \39093 , \39092 , \39002 );
and \U$38717 ( \39094 , \39091 , \39093 );
and \U$38718 ( \39095 , \39088 , \39090 );
or \U$38719 ( \39096 , \39094 , \39095 );
and \U$38720 ( \39097 , \39086 , \39096 );
and \U$38721 ( \39098 , \39083 , \39085 );
or \U$38722 ( \39099 , \39097 , \39098 );
and \U$38723 ( \39100 , \5896 , RIae76af0_56);
and \U$38724 ( \39101 , RIae76a00_54, \5894 );
nor \U$38725 ( \39102 , \39100 , \39101 );
and \U$38726 ( \39103 , \39102 , \5589 );
not \U$38727 ( \39104 , \39102 );
and \U$38728 ( \39105 , \39104 , \5590 );
nor \U$38729 ( \39106 , \39103 , \39105 );
and \U$38730 ( \39107 , \6172 , RIae76820_50);
and \U$38731 ( \39108 , RIae76910_52, \6170 );
nor \U$38732 ( \39109 , \39107 , \39108 );
and \U$38733 ( \39110 , \39109 , \6175 );
not \U$38734 ( \39111 , \39109 );
and \U$38735 ( \39112 , \39111 , \6176 );
nor \U$38736 ( \39113 , \39110 , \39112 );
xor \U$38737 ( \39114 , \39106 , \39113 );
and \U$38738 ( \39115 , \5399 , RIae76370_40);
and \U$38739 ( \39116 , RIae76280_38, \5397 );
nor \U$38740 ( \39117 , \39115 , \39116 );
and \U$38741 ( \39118 , \39117 , \5403 );
not \U$38742 ( \39119 , \39117 );
and \U$38743 ( \39120 , \39119 , \5016 );
nor \U$38744 ( \39121 , \39118 , \39120 );
and \U$38745 ( \39122 , \39114 , \39121 );
and \U$38746 ( \39123 , \39106 , \39113 );
nor \U$38747 ( \39124 , \39122 , \39123 );
and \U$38748 ( \39125 , \6941 , RIae76be0_58);
and \U$38749 ( \39126 , RIae78ad0_124, \6939 );
nor \U$38750 ( \39127 , \39125 , \39126 );
and \U$38751 ( \39128 , \39127 , \6945 );
not \U$38752 ( \39129 , \39127 );
and \U$38753 ( \39130 , \39129 , \6314 );
nor \U$38754 ( \39131 , \39128 , \39130 );
or \U$38755 ( \39132 , \39131 , \8019 );
not \U$38756 ( \39133 , \8019 );
not \U$38757 ( \39134 , \39131 );
or \U$38758 ( \39135 , \39133 , \39134 );
and \U$38759 ( \39136 , \7633 , RIae78d28_129);
and \U$38760 ( \39137 , RIae78e18_131, \7631 );
nor \U$38761 ( \39138 , \39136 , \39137 );
and \U$38762 ( \39139 , \39138 , \7206 );
not \U$38763 ( \39140 , \39138 );
and \U$38764 ( \39141 , \39140 , \7205 );
nor \U$38765 ( \39142 , \39139 , \39141 );
nand \U$38766 ( \39143 , \39135 , \39142 );
nand \U$38767 ( \39144 , \39132 , \39143 );
xor \U$38768 ( \39145 , \39124 , \39144 );
and \U$38769 ( \39146 , \3730 , RIae76460_42);
and \U$38770 ( \39147 , RIae76550_44, \3728 );
nor \U$38771 ( \39148 , \39146 , \39147 );
and \U$38772 ( \39149 , \39148 , \3422 );
not \U$38773 ( \39150 , \39148 );
and \U$38774 ( \39151 , \39150 , \3732 );
nor \U$38775 ( \39152 , \39149 , \39151 );
and \U$38776 ( \39153 , \4247 , RIae76730_48);
and \U$38777 ( \39154 , RIae76640_46, \4245 );
nor \U$38778 ( \39155 , \39153 , \39154 );
and \U$38779 ( \39156 , \39155 , \4251 );
not \U$38780 ( \39157 , \39155 );
and \U$38781 ( \39158 , \39157 , \3989 );
nor \U$38782 ( \39159 , \39156 , \39158 );
or \U$38783 ( \39160 , \39152 , \39159 );
not \U$38784 ( \39161 , \39159 );
not \U$38785 ( \39162 , \39152 );
or \U$38786 ( \39163 , \39161 , \39162 );
and \U$38787 ( \39164 , \4688 , RIae76190_36);
and \U$38788 ( \39165 , RIae760a0_34, \4686 );
nor \U$38789 ( \39166 , \39164 , \39165 );
and \U$38790 ( \39167 , \39166 , \4481 );
not \U$38791 ( \39168 , \39166 );
and \U$38792 ( \39169 , \39168 , \4482 );
nor \U$38793 ( \39170 , \39167 , \39169 );
nand \U$38794 ( \39171 , \39163 , \39170 );
nand \U$38795 ( \39172 , \39160 , \39171 );
and \U$38796 ( \39173 , \39145 , \39172 );
and \U$38797 ( \39174 , \39124 , \39144 );
nor \U$38798 ( \39175 , \39173 , \39174 );
and \U$38799 ( \39176 , \2783 , RIae75290_4);
and \U$38800 ( \39177 , RIae751a0_2, \2781 );
nor \U$38801 ( \39178 , \39176 , \39177 );
not \U$38802 ( \39179 , \39178 );
not \U$38803 ( \39180 , \2789 );
and \U$38804 ( \39181 , \39179 , \39180 );
and \U$38805 ( \39182 , \39178 , \2789 );
nor \U$38806 ( \39183 , \39181 , \39182 );
and \U$38807 ( \39184 , \2607 , RIae75830_16);
and \U$38808 ( \39185 , RIae75740_14, \2605 );
nor \U$38809 ( \39186 , \39184 , \39185 );
and \U$38810 ( \39187 , \39186 , \2397 );
not \U$38811 ( \39188 , \39186 );
and \U$38812 ( \39189 , \39188 , \2611 );
nor \U$38813 ( \39190 , \39187 , \39189 );
xor \U$38814 ( \39191 , \39183 , \39190 );
and \U$38815 ( \39192 , \3214 , RIae75380_6);
and \U$38816 ( \39193 , RIae75470_8, \3212 );
nor \U$38817 ( \39194 , \39192 , \39193 );
not \U$38818 ( \39195 , \39194 );
not \U$38819 ( \39196 , \2774 );
and \U$38820 ( \39197 , \39195 , \39196 );
and \U$38821 ( \39198 , \39194 , \2774 );
nor \U$38822 ( \39199 , \39197 , \39198 );
and \U$38823 ( \39200 , \39191 , \39199 );
and \U$38824 ( \39201 , \39183 , \39190 );
or \U$38825 ( \39202 , \39200 , \39201 );
and \U$38826 ( \39203 , \1138 , RIae75bf0_24);
and \U$38827 ( \39204 , RIae75b00_22, \1136 );
nor \U$38828 ( \39205 , \39203 , \39204 );
and \U$38829 ( \39206 , \39205 , \1142 );
not \U$38830 ( \39207 , \39205 );
and \U$38831 ( \39208 , \39207 , \1012 );
nor \U$38832 ( \39209 , \39206 , \39208 );
and \U$38833 ( \39210 , \883 , RIae78800_118);
and \U$38834 ( \39211 , RIae78710_116, \881 );
nor \U$38835 ( \39212 , \39210 , \39211 );
not \U$38836 ( \39213 , \39212 );
not \U$38837 ( \39214 , \789 );
and \U$38838 ( \39215 , \39213 , \39214 );
and \U$38839 ( \39216 , \39212 , \787 );
nor \U$38840 ( \39217 , \39215 , \39216 );
xor \U$38841 ( \39218 , \39209 , \39217 );
and \U$38842 ( \39219 , \1376 , RIae75a10_20);
and \U$38843 ( \39220 , RIae75920_18, \1374 );
nor \U$38844 ( \39221 , \39219 , \39220 );
and \U$38845 ( \39222 , \39221 , \1261 );
not \U$38846 ( \39223 , \39221 );
and \U$38847 ( \39224 , \39223 , \1380 );
nor \U$38848 ( \39225 , \39222 , \39224 );
and \U$38849 ( \39226 , \39218 , \39225 );
and \U$38850 ( \39227 , \39209 , \39217 );
or \U$38851 ( \39228 , \39226 , \39227 );
xor \U$38852 ( \39229 , \39202 , \39228 );
and \U$38853 ( \39230 , \1939 , RIae75ce0_26);
and \U$38854 ( \39231 , RIae75dd0_28, \1937 );
nor \U$38855 ( \39232 , \39230 , \39231 );
and \U$38856 ( \39233 , \39232 , \1734 );
not \U$38857 ( \39234 , \39232 );
and \U$38858 ( \39235 , \39234 , \1735 );
nor \U$38859 ( \39236 , \39233 , \39235 );
and \U$38860 ( \39237 , \1593 , RIae75fb0_32);
and \U$38861 ( \39238 , RIae75ec0_30, \1591 );
nor \U$38862 ( \39239 , \39237 , \39238 );
and \U$38863 ( \39240 , \39239 , \1488 );
not \U$38864 ( \39241 , \39239 );
and \U$38865 ( \39242 , \39241 , \1498 );
nor \U$38866 ( \39243 , \39240 , \39242 );
xor \U$38867 ( \39244 , \39236 , \39243 );
and \U$38868 ( \39245 , \2224 , RIae75650_12);
and \U$38869 ( \39246 , RIae75560_10, \2222 );
nor \U$38870 ( \39247 , \39245 , \39246 );
and \U$38871 ( \39248 , \39247 , \2060 );
not \U$38872 ( \39249 , \39247 );
and \U$38873 ( \39250 , \39249 , \2061 );
nor \U$38874 ( \39251 , \39248 , \39250 );
and \U$38875 ( \39252 , \39244 , \39251 );
and \U$38876 ( \39253 , \39236 , \39243 );
or \U$38877 ( \39254 , \39252 , \39253 );
and \U$38878 ( \39255 , \39229 , \39254 );
and \U$38879 ( \39256 , \39202 , \39228 );
or \U$38880 ( \39257 , \39255 , \39256 );
or \U$38881 ( \39258 , \39175 , \39257 );
not \U$38882 ( \39259 , \39175 );
not \U$38883 ( \39260 , \39257 );
or \U$38884 ( \39261 , \39259 , \39260 );
and \U$38885 ( \39262 , \436 , RIae78440_110);
and \U$38886 ( \39263 , RIae784b8_111, \434 );
nor \U$38887 ( \39264 , \39262 , \39263 );
not \U$38888 ( \39265 , \39264 );
not \U$38889 ( \39266 , \402 );
and \U$38890 ( \39267 , \39265 , \39266 );
and \U$38891 ( \39268 , \39264 , \402 );
nor \U$38892 ( \39269 , \39267 , \39268 );
nand \U$38893 ( \39270 , RIae78080_102, RIae78b48_125);
or \U$38894 ( \39271 , \39269 , \39270 );
not \U$38895 ( \39272 , \39270 );
not \U$38896 ( \39273 , \39269 );
or \U$38897 ( \39274 , \39272 , \39273 );
not \U$38898 ( \39275 , \392 );
and \U$38899 ( \39276 , \384 , RIae78260_106);
and \U$38900 ( \39277 , RIae78620_114, \382 );
nor \U$38901 ( \39278 , \39276 , \39277 );
not \U$38902 ( \39279 , \39278 );
or \U$38903 ( \39280 , \39275 , \39279 );
or \U$38904 ( \39281 , \39278 , \388 );
nand \U$38905 ( \39282 , \39280 , \39281 );
nand \U$38906 ( \39283 , \39274 , \39282 );
nand \U$38907 ( \39284 , \39271 , \39283 );
or \U$38908 ( \39285 , \38887 , \38879 );
nand \U$38909 ( \39286 , \39285 , \38888 );
xor \U$38910 ( \39287 , \39284 , \39286 );
and \U$38911 ( \39288 , \514 , RIae77cc0_94);
and \U$38912 ( \39289 , RIae77bd0_92, \512 );
nor \U$38913 ( \39290 , \39288 , \39289 );
not \U$38914 ( \39291 , \39290 );
not \U$38915 ( \39292 , \471 );
and \U$38916 ( \39293 , \39291 , \39292 );
and \U$38917 ( \39294 , \39290 , \471 );
nor \U$38918 ( \39295 , \39293 , \39294 );
and \U$38919 ( \39296 , \558 , RIae77db0_96);
and \U$38920 ( \39297 , RIae77ea0_98, \556 );
nor \U$38921 ( \39298 , \39296 , \39297 );
and \U$38922 ( \39299 , \39298 , \562 );
not \U$38923 ( \39300 , \39298 );
and \U$38924 ( \39301 , \39300 , \504 );
nor \U$38925 ( \39302 , \39299 , \39301 );
or \U$38926 ( \39303 , \39295 , \39302 );
not \U$38927 ( \39304 , \39302 );
not \U$38928 ( \39305 , \39295 );
or \U$38929 ( \39306 , \39304 , \39305 );
and \U$38930 ( \39307 , \672 , RIae789e0_122);
and \U$38931 ( \39308 , RIae788f0_120, \670 );
nor \U$38932 ( \39309 , \39307 , \39308 );
and \U$38933 ( \39310 , \39309 , \588 );
not \U$38934 ( \39311 , \39309 );
and \U$38935 ( \39312 , \39311 , \587 );
nor \U$38936 ( \39313 , \39310 , \39312 );
nand \U$38937 ( \39314 , \39306 , \39313 );
nand \U$38938 ( \39315 , \39303 , \39314 );
and \U$38939 ( \39316 , \39287 , \39315 );
and \U$38940 ( \39317 , \39284 , \39286 );
or \U$38941 ( \39318 , \39316 , \39317 );
nand \U$38942 ( \39319 , \39261 , \39318 );
nand \U$38943 ( \39320 , \39258 , \39319 );
xor \U$38944 ( \39321 , \39099 , \39320 );
xor \U$38945 ( \39322 , \38559 , \7206 );
xor \U$38946 ( \39323 , \39322 , \38567 );
xor \U$38947 ( \39324 , \38781 , \38783 );
xor \U$38948 ( \39325 , \39324 , \38786 );
and \U$38949 ( \39326 , \39323 , \39325 );
xor \U$38950 ( \39327 , \38578 , \38586 );
xor \U$38951 ( \39328 , \39327 , \38594 );
xor \U$38952 ( \39329 , \38769 , \38774 );
xor \U$38953 ( \39330 , \39328 , \39329 );
xor \U$38954 ( \39331 , \38781 , \38783 );
xor \U$38955 ( \39332 , \39331 , \38786 );
and \U$38956 ( \39333 , \39330 , \39332 );
and \U$38957 ( \39334 , \39323 , \39330 );
or \U$38958 ( \39335 , \39326 , \39333 , \39334 );
and \U$38959 ( \39336 , \39321 , \39335 );
and \U$38960 ( \39337 , \39099 , \39320 );
or \U$38961 ( \39338 , \39336 , \39337 );
xor \U$38962 ( \39339 , \38509 , \38511 );
xor \U$38963 ( \39340 , \39339 , \38524 );
xor \U$38964 ( \39341 , \39338 , \39340 );
xor \U$38965 ( \39342 , \38888 , \38896 );
xor \U$38966 ( \39343 , \39342 , \38924 );
xor \U$38967 ( \39344 , \38954 , \38979 );
xor \U$38968 ( \39345 , \39344 , \39005 );
and \U$38969 ( \39346 , \39343 , \39345 );
xor \U$38970 ( \39347 , \38823 , \38848 );
xor \U$38971 ( \39348 , \39347 , \38875 );
xor \U$38972 ( \39349 , \38954 , \38979 );
xor \U$38973 ( \39350 , \39349 , \39005 );
and \U$38974 ( \39351 , \39348 , \39350 );
and \U$38975 ( \39352 , \39343 , \39348 );
or \U$38976 ( \39353 , \39346 , \39351 , \39352 );
xor \U$38977 ( \39354 , \38552 , \38570 );
xor \U$38978 ( \39355 , \39354 , \38597 );
xor \U$38979 ( \39356 , \39353 , \39355 );
xor \U$38980 ( \39357 , \38627 , \37491 );
xor \U$38981 ( \39358 , \39357 , \38630 );
xor \U$38982 ( \39359 , \39014 , \39021 );
xor \U$38983 ( \39360 , \39358 , \39359 );
and \U$38984 ( \39361 , \39356 , \39360 );
and \U$38985 ( \39362 , \39353 , \39355 );
or \U$38986 ( \39363 , \39361 , \39362 );
and \U$38987 ( \39364 , \39341 , \39363 );
and \U$38988 ( \39365 , \39338 , \39340 );
or \U$38989 ( \39366 , \39364 , \39365 );
xor \U$38990 ( \39367 , \37623 , \37677 );
xor \U$38991 ( \39368 , \39367 , \37749 );
xor \U$38992 ( \39369 , \38741 , \38748 );
xor \U$38993 ( \39370 , \39368 , \39369 );
xor \U$38994 ( \39371 , \39366 , \39370 );
xor \U$38995 ( \39372 , \38600 , \38633 );
xor \U$38996 ( \39373 , \39372 , \38715 );
xor \U$38997 ( \39374 , \39034 , \39036 );
xor \U$38998 ( \39375 , \39374 , \39041 );
and \U$38999 ( \39376 , \39373 , \39375 );
xor \U$39000 ( \39377 , \38797 , \39011 );
xor \U$39001 ( \39378 , \39377 , \39026 );
xor \U$39002 ( \39379 , \39034 , \39036 );
xor \U$39003 ( \39380 , \39379 , \39041 );
and \U$39004 ( \39381 , \39378 , \39380 );
and \U$39005 ( \39382 , \39373 , \39378 );
or \U$39006 ( \39383 , \39376 , \39381 , \39382 );
and \U$39007 ( \39384 , \39371 , \39383 );
and \U$39008 ( \39385 , \39366 , \39370 );
or \U$39009 ( \39386 , \39384 , \39385 );
xor \U$39010 ( \39387 , \38527 , \38718 );
xor \U$39011 ( \39388 , \39387 , \38733 );
xor \U$39012 ( \39389 , \39029 , \39031 );
xor \U$39013 ( \39390 , \39389 , \39044 );
and \U$39014 ( \39391 , \39388 , \39390 );
xor \U$39015 ( \39392 , \39386 , \39391 );
xor \U$39016 ( \39393 , \38736 , \38738 );
xor \U$39017 ( \39394 , \39393 , \38753 );
xor \U$39018 ( \39395 , \39047 , \39054 );
xor \U$39019 ( \39396 , \39394 , \39395 );
and \U$39020 ( \39397 , \39392 , \39396 );
and \U$39021 ( \39398 , \39386 , \39391 );
or \U$39022 ( \39399 , \39397 , \39398 );
nand \U$39023 ( \39400 , \39071 , \39399 );
or \U$39024 ( \39401 , \39064 , \39400 );
not \U$39025 ( \39402 , \39063 );
not \U$39026 ( \39403 , \39400 );
and \U$39027 ( \39404 , \39402 , \39403 );
and \U$39028 ( \39405 , \39063 , \39400 );
nor \U$39029 ( \39406 , \39404 , \39405 );
not \U$39030 ( \39407 , \39399 );
not \U$39031 ( \39408 , \39070 );
or \U$39032 ( \39409 , \39407 , \39408 );
or \U$39033 ( \39410 , \39070 , \39399 );
nand \U$39034 ( \39411 , \39409 , \39410 );
xor \U$39035 ( \39412 , \38878 , \38927 );
xor \U$39036 ( \39413 , \39412 , \39008 );
xor \U$39037 ( \39414 , \39099 , \39320 );
xor \U$39038 ( \39415 , \39414 , \39335 );
and \U$39039 ( \39416 , \39413 , \39415 );
xor \U$39040 ( \39417 , \39353 , \39355 );
xor \U$39041 ( \39418 , \39417 , \39360 );
xor \U$39042 ( \39419 , \39099 , \39320 );
xor \U$39043 ( \39420 , \39419 , \39335 );
and \U$39044 ( \39421 , \39418 , \39420 );
and \U$39045 ( \39422 , \39413 , \39418 );
or \U$39046 ( \39423 , \39416 , \39421 , \39422 );
and \U$39047 ( \39424 , \6941 , RIae76910_52);
and \U$39048 ( \39425 , RIae76be0_58, \6939 );
nor \U$39049 ( \39426 , \39424 , \39425 );
and \U$39050 ( \39427 , \39426 , \6945 );
not \U$39051 ( \39428 , \39426 );
and \U$39052 ( \39429 , \39428 , \6314 );
nor \U$39053 ( \39430 , \39427 , \39429 );
nand \U$39054 ( \39431 , RIae78e18_131, \8371 );
and \U$39055 ( \39432 , \39431 , \8019 );
not \U$39056 ( \39433 , \39431 );
and \U$39057 ( \39434 , \39433 , \8020 );
nor \U$39058 ( \39435 , \39432 , \39434 );
xor \U$39059 ( \39436 , \39430 , \39435 );
and \U$39060 ( \39437 , \7633 , RIae78ad0_124);
and \U$39061 ( \39438 , RIae78d28_129, \7631 );
nor \U$39062 ( \39439 , \39437 , \39438 );
and \U$39063 ( \39440 , \39439 , \7205 );
not \U$39064 ( \39441 , \39439 );
and \U$39065 ( \39442 , \39441 , \7206 );
nor \U$39066 ( \39443 , \39440 , \39442 );
and \U$39067 ( \39444 , \39436 , \39443 );
and \U$39068 ( \39445 , \39430 , \39435 );
or \U$39069 ( \39446 , \39444 , \39445 );
and \U$39070 ( \39447 , \5896 , RIae76280_38);
and \U$39071 ( \39448 , RIae76af0_56, \5894 );
nor \U$39072 ( \39449 , \39447 , \39448 );
and \U$39073 ( \39450 , \39449 , \5590 );
not \U$39074 ( \39451 , \39449 );
and \U$39075 ( \39452 , \39451 , \5589 );
nor \U$39076 ( \39453 , \39450 , \39452 );
and \U$39077 ( \39454 , \6172 , RIae76a00_54);
and \U$39078 ( \39455 , RIae76820_50, \6170 );
nor \U$39079 ( \39456 , \39454 , \39455 );
and \U$39080 ( \39457 , \39456 , \6176 );
not \U$39081 ( \39458 , \39456 );
and \U$39082 ( \39459 , \39458 , \6175 );
nor \U$39083 ( \39460 , \39457 , \39459 );
xor \U$39084 ( \39461 , \39453 , \39460 );
and \U$39085 ( \39462 , \5399 , RIae760a0_34);
and \U$39086 ( \39463 , RIae76370_40, \5397 );
nor \U$39087 ( \39464 , \39462 , \39463 );
and \U$39088 ( \39465 , \39464 , \5016 );
not \U$39089 ( \39466 , \39464 );
and \U$39090 ( \39467 , \39466 , \5403 );
nor \U$39091 ( \39468 , \39465 , \39467 );
and \U$39092 ( \39469 , \39461 , \39468 );
and \U$39093 ( \39470 , \39453 , \39460 );
nor \U$39094 ( \39471 , \39469 , \39470 );
xor \U$39095 ( \39472 , \39446 , \39471 );
and \U$39096 ( \39473 , \4688 , RIae76640_46);
and \U$39097 ( \39474 , RIae76190_36, \4686 );
nor \U$39098 ( \39475 , \39473 , \39474 );
and \U$39099 ( \39476 , \39475 , \4482 );
not \U$39100 ( \39477 , \39475 );
and \U$39101 ( \39478 , \39477 , \4481 );
nor \U$39102 ( \39479 , \39476 , \39478 );
and \U$39103 ( \39480 , \3730 , RIae75470_8);
and \U$39104 ( \39481 , RIae76460_42, \3728 );
nor \U$39105 ( \39482 , \39480 , \39481 );
and \U$39106 ( \39483 , \39482 , \3422 );
not \U$39107 ( \39484 , \39482 );
and \U$39108 ( \39485 , \39484 , \3732 );
nor \U$39109 ( \39486 , \39483 , \39485 );
xor \U$39110 ( \39487 , \39479 , \39486 );
and \U$39111 ( \39488 , \4247 , RIae76550_44);
and \U$39112 ( \39489 , RIae76730_48, \4245 );
nor \U$39113 ( \39490 , \39488 , \39489 );
and \U$39114 ( \39491 , \39490 , \4251 );
not \U$39115 ( \39492 , \39490 );
and \U$39116 ( \39493 , \39492 , \3989 );
nor \U$39117 ( \39494 , \39491 , \39493 );
and \U$39118 ( \39495 , \39487 , \39494 );
and \U$39119 ( \39496 , \39479 , \39486 );
or \U$39120 ( \39497 , \39495 , \39496 );
and \U$39121 ( \39498 , \39472 , \39497 );
and \U$39122 ( \39499 , \39446 , \39471 );
nor \U$39123 ( \39500 , \39498 , \39499 );
and \U$39124 ( \39501 , \1593 , RIae75920_18);
and \U$39125 ( \39502 , RIae75fb0_32, \1591 );
nor \U$39126 ( \39503 , \39501 , \39502 );
and \U$39127 ( \39504 , \39503 , \1488 );
not \U$39128 ( \39505 , \39503 );
and \U$39129 ( \39506 , \39505 , \1498 );
nor \U$39130 ( \39507 , \39504 , \39506 );
and \U$39131 ( \39508 , \1939 , RIae75ec0_30);
and \U$39132 ( \39509 , RIae75ce0_26, \1937 );
nor \U$39133 ( \39510 , \39508 , \39509 );
and \U$39134 ( \39511 , \39510 , \1734 );
not \U$39135 ( \39512 , \39510 );
and \U$39136 ( \39513 , \39512 , \1735 );
nor \U$39137 ( \39514 , \39511 , \39513 );
xor \U$39138 ( \39515 , \39507 , \39514 );
and \U$39139 ( \39516 , \2224 , RIae75dd0_28);
and \U$39140 ( \39517 , RIae75650_12, \2222 );
nor \U$39141 ( \39518 , \39516 , \39517 );
and \U$39142 ( \39519 , \39518 , \2060 );
not \U$39143 ( \39520 , \39518 );
and \U$39144 ( \39521 , \39520 , \2061 );
nor \U$39145 ( \39522 , \39519 , \39521 );
and \U$39146 ( \39523 , \39515 , \39522 );
and \U$39147 ( \39524 , \39507 , \39514 );
or \U$39148 ( \39525 , \39523 , \39524 );
and \U$39149 ( \39526 , \3214 , RIae751a0_2);
and \U$39150 ( \39527 , RIae75380_6, \3212 );
nor \U$39151 ( \39528 , \39526 , \39527 );
not \U$39152 ( \39529 , \39528 );
not \U$39153 ( \39530 , \2774 );
and \U$39154 ( \39531 , \39529 , \39530 );
and \U$39155 ( \39532 , \39528 , \2774 );
nor \U$39156 ( \39533 , \39531 , \39532 );
and \U$39157 ( \39534 , \2607 , RIae75560_10);
and \U$39158 ( \39535 , RIae75830_16, \2605 );
nor \U$39159 ( \39536 , \39534 , \39535 );
and \U$39160 ( \39537 , \39536 , \2397 );
not \U$39161 ( \39538 , \39536 );
and \U$39162 ( \39539 , \39538 , \2611 );
nor \U$39163 ( \39540 , \39537 , \39539 );
xor \U$39164 ( \39541 , \39533 , \39540 );
and \U$39165 ( \39542 , \2783 , RIae75740_14);
and \U$39166 ( \39543 , RIae75290_4, \2781 );
nor \U$39167 ( \39544 , \39542 , \39543 );
not \U$39168 ( \39545 , \39544 );
not \U$39169 ( \39546 , \2789 );
and \U$39170 ( \39547 , \39545 , \39546 );
and \U$39171 ( \39548 , \39544 , \2789 );
nor \U$39172 ( \39549 , \39547 , \39548 );
and \U$39173 ( \39550 , \39541 , \39549 );
and \U$39174 ( \39551 , \39533 , \39540 );
or \U$39175 ( \39552 , \39550 , \39551 );
xor \U$39176 ( \39553 , \39525 , \39552 );
and \U$39177 ( \39554 , \883 , RIae788f0_120);
and \U$39178 ( \39555 , RIae78800_118, \881 );
nor \U$39179 ( \39556 , \39554 , \39555 );
not \U$39180 ( \39557 , \39556 );
not \U$39181 ( \39558 , \787 );
and \U$39182 ( \39559 , \39557 , \39558 );
and \U$39183 ( \39560 , \39556 , \787 );
nor \U$39184 ( \39561 , \39559 , \39560 );
and \U$39185 ( \39562 , \1138 , RIae78710_116);
and \U$39186 ( \39563 , RIae75bf0_24, \1136 );
nor \U$39187 ( \39564 , \39562 , \39563 );
and \U$39188 ( \39565 , \39564 , \1142 );
not \U$39189 ( \39566 , \39564 );
and \U$39190 ( \39567 , \39566 , \1012 );
nor \U$39191 ( \39568 , \39565 , \39567 );
xor \U$39192 ( \39569 , \39561 , \39568 );
and \U$39193 ( \39570 , \1376 , RIae75b00_22);
and \U$39194 ( \39571 , RIae75a10_20, \1374 );
nor \U$39195 ( \39572 , \39570 , \39571 );
and \U$39196 ( \39573 , \39572 , \1261 );
not \U$39197 ( \39574 , \39572 );
and \U$39198 ( \39575 , \39574 , \1380 );
nor \U$39199 ( \39576 , \39573 , \39575 );
and \U$39200 ( \39577 , \39569 , \39576 );
and \U$39201 ( \39578 , \39561 , \39568 );
or \U$39202 ( \39579 , \39577 , \39578 );
and \U$39203 ( \39580 , \39553 , \39579 );
and \U$39204 ( \39581 , \39525 , \39552 );
nor \U$39205 ( \39582 , \39580 , \39581 );
and \U$39206 ( \39583 , \39500 , \39582 );
not \U$39207 ( \39584 , \39582 );
not \U$39208 ( \39585 , \39500 );
and \U$39209 ( \39586 , \39584 , \39585 );
and \U$39210 ( \39587 , \514 , RIae784b8_111);
and \U$39211 ( \39588 , RIae77cc0_94, \512 );
nor \U$39212 ( \39589 , \39587 , \39588 );
not \U$39213 ( \39590 , \39589 );
not \U$39214 ( \39591 , \471 );
and \U$39215 ( \39592 , \39590 , \39591 );
and \U$39216 ( \39593 , \39589 , \469 );
nor \U$39217 ( \39594 , \39592 , \39593 );
and \U$39218 ( \39595 , \558 , RIae77bd0_92);
and \U$39219 ( \39596 , RIae77db0_96, \556 );
nor \U$39220 ( \39597 , \39595 , \39596 );
and \U$39221 ( \39598 , \39597 , \562 );
not \U$39222 ( \39599 , \39597 );
and \U$39223 ( \39600 , \39599 , \504 );
nor \U$39224 ( \39601 , \39598 , \39600 );
xor \U$39225 ( \39602 , \39594 , \39601 );
and \U$39226 ( \39603 , \672 , RIae77ea0_98);
and \U$39227 ( \39604 , RIae789e0_122, \670 );
nor \U$39228 ( \39605 , \39603 , \39604 );
and \U$39229 ( \39606 , \39605 , \587 );
not \U$39230 ( \39607 , \39605 );
and \U$39231 ( \39608 , \39607 , \588 );
nor \U$39232 ( \39609 , \39606 , \39608 );
and \U$39233 ( \39610 , \39602 , \39609 );
and \U$39234 ( \39611 , \39594 , \39601 );
or \U$39235 ( \39612 , \39610 , \39611 );
and \U$39236 ( \39613 , \436 , RIae78620_114);
and \U$39237 ( \39614 , RIae78440_110, \434 );
nor \U$39238 ( \39615 , \39613 , \39614 );
not \U$39239 ( \39616 , \39615 );
not \U$39240 ( \39617 , \402 );
and \U$39241 ( \39618 , \39616 , \39617 );
and \U$39242 ( \39619 , \39615 , \400 );
nor \U$39243 ( \39620 , \39618 , \39619 );
nand \U$39244 ( \39621 , RIae77f90_100, RIae78b48_125);
xor \U$39245 ( \39622 , \39620 , \39621 );
and \U$39246 ( \39623 , \384 , RIae78080_102);
and \U$39247 ( \39624 , RIae78260_106, \382 );
nor \U$39248 ( \39625 , \39623 , \39624 );
not \U$39249 ( \39626 , \39625 );
not \U$39250 ( \39627 , \392 );
and \U$39251 ( \39628 , \39626 , \39627 );
and \U$39252 ( \39629 , \39625 , \388 );
nor \U$39253 ( \39630 , \39628 , \39629 );
and \U$39254 ( \39631 , \39622 , \39630 );
and \U$39255 ( \39632 , \39620 , \39621 );
or \U$39256 ( \39633 , \39631 , \39632 );
xor \U$39257 ( \39634 , \39612 , \39633 );
not \U$39258 ( \39635 , \39269 );
not \U$39259 ( \39636 , \39282 );
or \U$39260 ( \39637 , \39635 , \39636 );
or \U$39261 ( \39638 , \39269 , \39282 );
nand \U$39262 ( \39639 , \39637 , \39638 );
not \U$39263 ( \39640 , \39639 );
not \U$39264 ( \39641 , \39270 );
and \U$39265 ( \39642 , \39640 , \39641 );
and \U$39266 ( \39643 , \39639 , \39270 );
nor \U$39267 ( \39644 , \39642 , \39643 );
and \U$39268 ( \39645 , \39634 , \39644 );
and \U$39269 ( \39646 , \39612 , \39633 );
or \U$39270 ( \39647 , \39645 , \39646 );
nor \U$39271 ( \39648 , \39586 , \39647 );
nor \U$39272 ( \39649 , \39583 , \39648 );
not \U$39273 ( \39650 , \39159 );
not \U$39274 ( \39651 , \39170 );
or \U$39275 ( \39652 , \39650 , \39651 );
or \U$39276 ( \39653 , \39159 , \39170 );
nand \U$39277 ( \39654 , \39652 , \39653 );
not \U$39278 ( \39655 , \39654 );
not \U$39279 ( \39656 , \39152 );
and \U$39280 ( \39657 , \39655 , \39656 );
and \U$39281 ( \39658 , \39654 , \39152 );
nor \U$39282 ( \39659 , \39657 , \39658 );
xor \U$39283 ( \39660 , \39183 , \39190 );
xor \U$39284 ( \39661 , \39660 , \39199 );
xor \U$39285 ( \39662 , \39659 , \39661 );
xor \U$39286 ( \39663 , \39106 , \39113 );
xor \U$39287 ( \39664 , \39663 , \39121 );
and \U$39288 ( \39665 , \39662 , \39664 );
and \U$39289 ( \39666 , \39659 , \39661 );
or \U$39290 ( \39667 , \39665 , \39666 );
not \U$39291 ( \39668 , \39667 );
not \U$39292 ( \39669 , \38977 );
not \U$39293 ( \39670 , \38968 );
or \U$39294 ( \39671 , \39669 , \39670 );
or \U$39295 ( \39672 , \38968 , \38977 );
nand \U$39296 ( \39673 , \39671 , \39672 );
not \U$39297 ( \39674 , \39673 );
not \U$39298 ( \39675 , \38961 );
and \U$39299 ( \39676 , \39674 , \39675 );
and \U$39300 ( \39677 , \39673 , \38961 );
nor \U$39301 ( \39678 , \39676 , \39677 );
not \U$39302 ( \39679 , \39678 );
and \U$39303 ( \39680 , \39668 , \39679 );
and \U$39304 ( \39681 , \39667 , \39678 );
not \U$39305 ( \39682 , \39302 );
not \U$39306 ( \39683 , \39313 );
or \U$39307 ( \39684 , \39682 , \39683 );
or \U$39308 ( \39685 , \39302 , \39313 );
nand \U$39309 ( \39686 , \39684 , \39685 );
not \U$39310 ( \39687 , \39686 );
not \U$39311 ( \39688 , \39295 );
and \U$39312 ( \39689 , \39687 , \39688 );
and \U$39313 ( \39690 , \39686 , \39295 );
nor \U$39314 ( \39691 , \39689 , \39690 );
xor \U$39315 ( \39692 , \39209 , \39217 );
xor \U$39316 ( \39693 , \39692 , \39225 );
xor \U$39317 ( \39694 , \39691 , \39693 );
xor \U$39318 ( \39695 , \39236 , \39243 );
xor \U$39319 ( \39696 , \39695 , \39251 );
and \U$39320 ( \39697 , \39694 , \39696 );
and \U$39321 ( \39698 , \39691 , \39693 );
or \U$39322 ( \39699 , \39697 , \39698 );
nor \U$39323 ( \39700 , \39681 , \39699 );
nor \U$39324 ( \39701 , \39680 , \39700 );
or \U$39325 ( \39702 , \39649 , \39701 );
not \U$39326 ( \39703 , \39701 );
not \U$39327 ( \39704 , \39649 );
or \U$39328 ( \39705 , \39703 , \39704 );
xor \U$39329 ( \39706 , \39284 , \39286 );
xor \U$39330 ( \39707 , \39706 , \39315 );
xor \U$39331 ( \39708 , \39088 , \39090 );
xor \U$39332 ( \39709 , \39708 , \39093 );
and \U$39333 ( \39710 , \39707 , \39709 );
xor \U$39334 ( \39711 , \38856 , \38863 );
xor \U$39335 ( \39712 , \39711 , \38872 );
xor \U$39336 ( \39713 , \39073 , \39078 );
xor \U$39337 ( \39714 , \39712 , \39713 );
xor \U$39338 ( \39715 , \39088 , \39090 );
xor \U$39339 ( \39716 , \39715 , \39093 );
and \U$39340 ( \39717 , \39714 , \39716 );
and \U$39341 ( \39718 , \39707 , \39714 );
or \U$39342 ( \39719 , \39710 , \39717 , \39718 );
nand \U$39343 ( \39720 , \39705 , \39719 );
nand \U$39344 ( \39721 , \39702 , \39720 );
xor \U$39345 ( \39722 , \38779 , \38789 );
xor \U$39346 ( \39723 , \39722 , \38794 );
xor \U$39347 ( \39724 , \39721 , \39723 );
xor \U$39348 ( \39725 , \38954 , \38979 );
xor \U$39349 ( \39726 , \39725 , \39005 );
xor \U$39350 ( \39727 , \39343 , \39348 );
xor \U$39351 ( \39728 , \39726 , \39727 );
xor \U$39352 ( \39729 , \39083 , \39085 );
xor \U$39353 ( \39730 , \39729 , \39096 );
and \U$39354 ( \39731 , \39728 , \39730 );
xor \U$39355 ( \39732 , \38781 , \38783 );
xor \U$39356 ( \39733 , \39732 , \38786 );
xor \U$39357 ( \39734 , \39323 , \39330 );
xor \U$39358 ( \39735 , \39733 , \39734 );
xor \U$39359 ( \39736 , \39083 , \39085 );
xor \U$39360 ( \39737 , \39736 , \39096 );
and \U$39361 ( \39738 , \39735 , \39737 );
and \U$39362 ( \39739 , \39728 , \39735 );
or \U$39363 ( \39740 , \39731 , \39738 , \39739 );
and \U$39364 ( \39741 , \39724 , \39740 );
and \U$39365 ( \39742 , \39721 , \39723 );
or \U$39366 ( \39743 , \39741 , \39742 );
xor \U$39367 ( \39744 , \39423 , \39743 );
xor \U$39368 ( \39745 , \39034 , \39036 );
xor \U$39369 ( \39746 , \39745 , \39041 );
xor \U$39370 ( \39747 , \39373 , \39378 );
xor \U$39371 ( \39748 , \39746 , \39747 );
and \U$39372 ( \39749 , \39744 , \39748 );
and \U$39373 ( \39750 , \39423 , \39743 );
or \U$39374 ( \39751 , \39749 , \39750 );
xor \U$39375 ( \39752 , \39388 , \39390 );
xor \U$39376 ( \39753 , \39751 , \39752 );
xor \U$39377 ( \39754 , \39366 , \39370 );
xor \U$39378 ( \39755 , \39754 , \39383 );
and \U$39379 ( \39756 , \39753 , \39755 );
and \U$39380 ( \39757 , \39751 , \39752 );
or \U$39381 ( \39758 , \39756 , \39757 );
xor \U$39382 ( \39759 , \39386 , \39391 );
xor \U$39383 ( \39760 , \39759 , \39396 );
and \U$39384 ( \39761 , \39758 , \39760 );
and \U$39385 ( \39762 , \39411 , \39761 );
xor \U$39386 ( \39763 , \39761 , \39411 );
xor \U$39387 ( \39764 , \39758 , \39760 );
not \U$39388 ( \39765 , \39764 );
xor \U$39389 ( \39766 , \39423 , \39743 );
xor \U$39390 ( \39767 , \39766 , \39748 );
xor \U$39391 ( \39768 , \39338 , \39340 );
xor \U$39392 ( \39769 , \39768 , \39363 );
xor \U$39393 ( \39770 , \39767 , \39769 );
not \U$39394 ( \39771 , \39678 );
xor \U$39395 ( \39772 , \39699 , \39667 );
not \U$39396 ( \39773 , \39772 );
or \U$39397 ( \39774 , \39771 , \39773 );
or \U$39398 ( \39775 , \39772 , \39678 );
nand \U$39399 ( \39776 , \39774 , \39775 );
not \U$39400 ( \39777 , \39647 );
xor \U$39401 ( \39778 , \39582 , \39500 );
not \U$39402 ( \39779 , \39778 );
or \U$39403 ( \39780 , \39777 , \39779 );
or \U$39404 ( \39781 , \39778 , \39647 );
nand \U$39405 ( \39782 , \39780 , \39781 );
xor \U$39406 ( \39783 , \39776 , \39782 );
xor \U$39407 ( \39784 , \39088 , \39090 );
xor \U$39408 ( \39785 , \39784 , \39093 );
xor \U$39409 ( \39786 , \39707 , \39714 );
xor \U$39410 ( \39787 , \39785 , \39786 );
and \U$39411 ( \39788 , \39783 , \39787 );
and \U$39412 ( \39789 , \39776 , \39782 );
nor \U$39413 ( \39790 , \39788 , \39789 );
xor \U$39414 ( \39791 , \39124 , \39144 );
xor \U$39415 ( \39792 , \39791 , \39172 );
xor \U$39416 ( \39793 , \39202 , \39228 );
xor \U$39417 ( \39794 , \39793 , \39254 );
not \U$39418 ( \39795 , \39794 );
and \U$39419 ( \39796 , \39792 , \39795 );
not \U$39420 ( \39797 , \39792 );
not \U$39421 ( \39798 , \39795 );
and \U$39422 ( \39799 , \39797 , \39798 );
xor \U$39423 ( \39800 , \39612 , \39633 );
xor \U$39424 ( \39801 , \39800 , \39644 );
xor \U$39425 ( \39802 , \39446 , \39471 );
xor \U$39426 ( \39803 , \39802 , \39497 );
xor \U$39427 ( \39804 , \39801 , \39803 );
xor \U$39428 ( \39805 , \39525 , \39552 );
xor \U$39429 ( \39806 , \39805 , \39579 );
and \U$39430 ( \39807 , \39804 , \39806 );
and \U$39431 ( \39808 , \39801 , \39803 );
or \U$39432 ( \39809 , \39807 , \39808 );
nor \U$39433 ( \39810 , \39799 , \39809 );
nor \U$39434 ( \39811 , \39796 , \39810 );
or \U$39435 ( \39812 , \39790 , \39811 );
not \U$39436 ( \39813 , \39811 );
not \U$39437 ( \39814 , \39790 );
or \U$39438 ( \39815 , \39813 , \39814 );
xor \U$39439 ( \39816 , \39594 , \39601 );
xor \U$39440 ( \39817 , \39816 , \39609 );
xor \U$39441 ( \39818 , \39561 , \39568 );
xor \U$39442 ( \39819 , \39818 , \39576 );
xor \U$39443 ( \39820 , \39817 , \39819 );
xor \U$39444 ( \39821 , \39620 , \39621 );
xor \U$39445 ( \39822 , \39821 , \39630 );
and \U$39446 ( \39823 , \39820 , \39822 );
and \U$39447 ( \39824 , \39817 , \39819 );
nor \U$39448 ( \39825 , \39823 , \39824 );
xor \U$39449 ( \39826 , \39453 , \39460 );
xor \U$39450 ( \39827 , \39826 , \39468 );
not \U$39451 ( \39828 , \39827 );
xor \U$39452 ( \39829 , \39430 , \39435 );
xor \U$39453 ( \39830 , \39829 , \39443 );
nor \U$39454 ( \39831 , \39828 , \39830 );
xor \U$39455 ( \39832 , \39825 , \39831 );
xor \U$39456 ( \39833 , \39507 , \39514 );
xor \U$39457 ( \39834 , \39833 , \39522 );
xor \U$39458 ( \39835 , \39533 , \39540 );
xor \U$39459 ( \39836 , \39835 , \39549 );
xor \U$39460 ( \39837 , \39834 , \39836 );
xor \U$39461 ( \39838 , \39479 , \39486 );
xor \U$39462 ( \39839 , \39838 , \39494 );
and \U$39463 ( \39840 , \39837 , \39839 );
and \U$39464 ( \39841 , \39834 , \39836 );
nor \U$39465 ( \39842 , \39840 , \39841 );
and \U$39466 ( \39843 , \39832 , \39842 );
and \U$39467 ( \39844 , \39825 , \39831 );
or \U$39468 ( \39845 , \39843 , \39844 );
not \U$39469 ( \39846 , \402 );
and \U$39470 ( \39847 , \436 , RIae78260_106);
and \U$39471 ( \39848 , RIae78620_114, \434 );
nor \U$39472 ( \39849 , \39847 , \39848 );
not \U$39473 ( \39850 , \39849 );
or \U$39474 ( \39851 , \39846 , \39850 );
or \U$39475 ( \39852 , \39849 , \400 );
nand \U$39476 ( \39853 , \39851 , \39852 );
not \U$39477 ( \39854 , \392 );
and \U$39478 ( \39855 , \384 , RIae77f90_100);
and \U$39479 ( \39856 , RIae78080_102, \382 );
nor \U$39480 ( \39857 , \39855 , \39856 );
not \U$39481 ( \39858 , \39857 );
or \U$39482 ( \39859 , \39854 , \39858 );
or \U$39483 ( \39860 , \39857 , \392 );
nand \U$39484 ( \39861 , \39859 , \39860 );
xor \U$39485 ( \39862 , \39853 , \39861 );
not \U$39486 ( \39863 , \471 );
and \U$39487 ( \39864 , \514 , RIae78440_110);
and \U$39488 ( \39865 , RIae784b8_111, \512 );
nor \U$39489 ( \39866 , \39864 , \39865 );
not \U$39490 ( \39867 , \39866 );
or \U$39491 ( \39868 , \39863 , \39867 );
or \U$39492 ( \39869 , \39866 , \469 );
nand \U$39493 ( \39870 , \39868 , \39869 );
and \U$39494 ( \39871 , \39862 , \39870 );
and \U$39495 ( \39872 , \39853 , \39861 );
or \U$39496 ( \39873 , \39871 , \39872 );
not \U$39497 ( \39874 , \787 );
and \U$39498 ( \39875 , \883 , RIae789e0_122);
and \U$39499 ( \39876 , RIae788f0_120, \881 );
nor \U$39500 ( \39877 , \39875 , \39876 );
not \U$39501 ( \39878 , \39877 );
or \U$39502 ( \39879 , \39874 , \39878 );
or \U$39503 ( \39880 , \39877 , \789 );
nand \U$39504 ( \39881 , \39879 , \39880 );
and \U$39505 ( \39882 , \558 , RIae77cc0_94);
and \U$39506 ( \39883 , RIae77bd0_92, \556 );
nor \U$39507 ( \39884 , \39882 , \39883 );
and \U$39508 ( \39885 , \39884 , \504 );
not \U$39509 ( \39886 , \39884 );
and \U$39510 ( \39887 , \39886 , \562 );
nor \U$39511 ( \39888 , \39885 , \39887 );
xor \U$39512 ( \39889 , \39881 , \39888 );
and \U$39513 ( \39890 , \672 , RIae77db0_96);
and \U$39514 ( \39891 , RIae77ea0_98, \670 );
nor \U$39515 ( \39892 , \39890 , \39891 );
and \U$39516 ( \39893 , \39892 , \588 );
not \U$39517 ( \39894 , \39892 );
and \U$39518 ( \39895 , \39894 , \587 );
nor \U$39519 ( \39896 , \39893 , \39895 );
and \U$39520 ( \39897 , \39889 , \39896 );
and \U$39521 ( \39898 , \39881 , \39888 );
or \U$39522 ( \39899 , \39897 , \39898 );
nor \U$39523 ( \39900 , \39873 , \39899 );
not \U$39524 ( \39901 , \39900 );
not \U$39525 ( \39902 , \39901 );
and \U$39526 ( \39903 , \1138 , RIae78800_118);
and \U$39527 ( \39904 , RIae78710_116, \1136 );
nor \U$39528 ( \39905 , \39903 , \39904 );
and \U$39529 ( \39906 , \39905 , \1142 );
not \U$39530 ( \39907 , \39905 );
and \U$39531 ( \39908 , \39907 , \1012 );
nor \U$39532 ( \39909 , \39906 , \39908 );
and \U$39533 ( \39910 , \1376 , RIae75bf0_24);
and \U$39534 ( \39911 , RIae75b00_22, \1374 );
nor \U$39535 ( \39912 , \39910 , \39911 );
and \U$39536 ( \39913 , \39912 , \1261 );
not \U$39537 ( \39914 , \39912 );
and \U$39538 ( \39915 , \39914 , \1380 );
nor \U$39539 ( \39916 , \39913 , \39915 );
xor \U$39540 ( \39917 , \39909 , \39916 );
and \U$39541 ( \39918 , \1593 , RIae75a10_20);
and \U$39542 ( \39919 , RIae75920_18, \1591 );
nor \U$39543 ( \39920 , \39918 , \39919 );
and \U$39544 ( \39921 , \39920 , \1488 );
not \U$39545 ( \39922 , \39920 );
and \U$39546 ( \39923 , \39922 , \1498 );
nor \U$39547 ( \39924 , \39921 , \39923 );
and \U$39548 ( \39925 , \39917 , \39924 );
and \U$39549 ( \39926 , \39909 , \39916 );
or \U$39550 ( \39927 , \39925 , \39926 );
and \U$39551 ( \39928 , \2224 , RIae75ce0_26);
and \U$39552 ( \39929 , RIae75dd0_28, \2222 );
nor \U$39553 ( \39930 , \39928 , \39929 );
and \U$39554 ( \39931 , \39930 , \2060 );
not \U$39555 ( \39932 , \39930 );
and \U$39556 ( \39933 , \39932 , \2061 );
nor \U$39557 ( \39934 , \39931 , \39933 );
and \U$39558 ( \39935 , \1939 , RIae75fb0_32);
and \U$39559 ( \39936 , RIae75ec0_30, \1937 );
nor \U$39560 ( \39937 , \39935 , \39936 );
and \U$39561 ( \39938 , \39937 , \1734 );
not \U$39562 ( \39939 , \39937 );
and \U$39563 ( \39940 , \39939 , \1735 );
nor \U$39564 ( \39941 , \39938 , \39940 );
xor \U$39565 ( \39942 , \39934 , \39941 );
and \U$39566 ( \39943 , \2607 , RIae75650_12);
and \U$39567 ( \39944 , RIae75560_10, \2605 );
nor \U$39568 ( \39945 , \39943 , \39944 );
and \U$39569 ( \39946 , \39945 , \2397 );
not \U$39570 ( \39947 , \39945 );
and \U$39571 ( \39948 , \39947 , \2611 );
nor \U$39572 ( \39949 , \39946 , \39948 );
and \U$39573 ( \39950 , \39942 , \39949 );
and \U$39574 ( \39951 , \39934 , \39941 );
or \U$39575 ( \39952 , \39950 , \39951 );
xor \U$39576 ( \39953 , \39927 , \39952 );
and \U$39577 ( \39954 , \2783 , RIae75830_16);
and \U$39578 ( \39955 , RIae75740_14, \2781 );
nor \U$39579 ( \39956 , \39954 , \39955 );
not \U$39580 ( \39957 , \39956 );
not \U$39581 ( \39958 , \3089 );
and \U$39582 ( \39959 , \39957 , \39958 );
and \U$39583 ( \39960 , \39956 , \3089 );
nor \U$39584 ( \39961 , \39959 , \39960 );
and \U$39585 ( \39962 , \3214 , RIae75290_4);
and \U$39586 ( \39963 , RIae751a0_2, \3212 );
nor \U$39587 ( \39964 , \39962 , \39963 );
not \U$39588 ( \39965 , \39964 );
not \U$39589 ( \39966 , \3218 );
and \U$39590 ( \39967 , \39965 , \39966 );
and \U$39591 ( \39968 , \39964 , \2774 );
nor \U$39592 ( \39969 , \39967 , \39968 );
xor \U$39593 ( \39970 , \39961 , \39969 );
and \U$39594 ( \39971 , \3730 , RIae75380_6);
and \U$39595 ( \39972 , RIae75470_8, \3728 );
nor \U$39596 ( \39973 , \39971 , \39972 );
and \U$39597 ( \39974 , \39973 , \3422 );
not \U$39598 ( \39975 , \39973 );
and \U$39599 ( \39976 , \39975 , \3732 );
nor \U$39600 ( \39977 , \39974 , \39976 );
and \U$39601 ( \39978 , \39970 , \39977 );
and \U$39602 ( \39979 , \39961 , \39969 );
or \U$39603 ( \39980 , \39978 , \39979 );
and \U$39604 ( \39981 , \39953 , \39980 );
and \U$39605 ( \39982 , \39927 , \39952 );
nor \U$39606 ( \39983 , \39981 , \39982 );
not \U$39607 ( \39984 , \39983 );
or \U$39608 ( \39985 , \39902 , \39984 );
or \U$39609 ( \39986 , \39983 , \39901 );
and \U$39610 ( \39987 , \7633 , RIae76be0_58);
and \U$39611 ( \39988 , RIae78ad0_124, \7631 );
nor \U$39612 ( \39989 , \39987 , \39988 );
and \U$39613 ( \39990 , \39989 , \7205 );
not \U$39614 ( \39991 , \39989 );
and \U$39615 ( \39992 , \39991 , \7206 );
nor \U$39616 ( \39993 , \39990 , \39992 );
not \U$39617 ( \39994 , \39993 );
not \U$39618 ( \39995 , \8789 );
and \U$39619 ( \39996 , \39994 , \39995 );
and \U$39620 ( \39997 , \39993 , \8789 );
and \U$39621 ( \39998 , \8371 , RIae78d28_129);
and \U$39622 ( \39999 , RIae78e18_131, \8369 );
nor \U$39623 ( \40000 , \39998 , \39999 );
and \U$39624 ( \40001 , \40000 , \8019 );
not \U$39625 ( \40002 , \40000 );
and \U$39626 ( \40003 , \40002 , \8020 );
nor \U$39627 ( \40004 , \40001 , \40003 );
nor \U$39628 ( \40005 , \39997 , \40004 );
nor \U$39629 ( \40006 , \39996 , \40005 );
and \U$39630 ( \40007 , \5896 , RIae76370_40);
and \U$39631 ( \40008 , RIae76280_38, \5894 );
nor \U$39632 ( \40009 , \40007 , \40008 );
and \U$39633 ( \40010 , \40009 , \5589 );
not \U$39634 ( \40011 , \40009 );
and \U$39635 ( \40012 , \40011 , \5590 );
nor \U$39636 ( \40013 , \40010 , \40012 );
not \U$39637 ( \40014 , \40013 );
and \U$39638 ( \40015 , \6941 , RIae76820_50);
and \U$39639 ( \40016 , RIae76910_52, \6939 );
nor \U$39640 ( \40017 , \40015 , \40016 );
and \U$39641 ( \40018 , \40017 , \6945 );
not \U$39642 ( \40019 , \40017 );
and \U$39643 ( \40020 , \40019 , \6314 );
nor \U$39644 ( \40021 , \40018 , \40020 );
not \U$39645 ( \40022 , \40021 );
and \U$39646 ( \40023 , \40014 , \40022 );
and \U$39647 ( \40024 , \40021 , \40013 );
and \U$39648 ( \40025 , \6172 , RIae76af0_56);
and \U$39649 ( \40026 , RIae76a00_54, \6170 );
nor \U$39650 ( \40027 , \40025 , \40026 );
and \U$39651 ( \40028 , \40027 , \6175 );
not \U$39652 ( \40029 , \40027 );
and \U$39653 ( \40030 , \40029 , \6176 );
nor \U$39654 ( \40031 , \40028 , \40030 );
nor \U$39655 ( \40032 , \40024 , \40031 );
nor \U$39656 ( \40033 , \40023 , \40032 );
xor \U$39657 ( \40034 , \40006 , \40033 );
and \U$39658 ( \40035 , \4688 , RIae76730_48);
and \U$39659 ( \40036 , RIae76640_46, \4686 );
nor \U$39660 ( \40037 , \40035 , \40036 );
and \U$39661 ( \40038 , \40037 , \4481 );
not \U$39662 ( \40039 , \40037 );
and \U$39663 ( \40040 , \40039 , \4482 );
nor \U$39664 ( \40041 , \40038 , \40040 );
and \U$39665 ( \40042 , \5399 , RIae76190_36);
and \U$39666 ( \40043 , RIae760a0_34, \5397 );
nor \U$39667 ( \40044 , \40042 , \40043 );
and \U$39668 ( \40045 , \40044 , \5016 );
not \U$39669 ( \40046 , \40044 );
and \U$39670 ( \40047 , \40046 , \5403 );
nor \U$39671 ( \40048 , \40045 , \40047 );
xor \U$39672 ( \40049 , \40041 , \40048 );
and \U$39673 ( \40050 , \4247 , RIae76460_42);
and \U$39674 ( \40051 , RIae76550_44, \4245 );
nor \U$39675 ( \40052 , \40050 , \40051 );
and \U$39676 ( \40053 , \40052 , \3989 );
not \U$39677 ( \40054 , \40052 );
and \U$39678 ( \40055 , \40054 , \4251 );
nor \U$39679 ( \40056 , \40053 , \40055 );
and \U$39680 ( \40057 , \40049 , \40056 );
and \U$39681 ( \40058 , \40041 , \40048 );
nor \U$39682 ( \40059 , \40057 , \40058 );
and \U$39683 ( \40060 , \40034 , \40059 );
and \U$39684 ( \40061 , \40006 , \40033 );
nor \U$39685 ( \40062 , \40060 , \40061 );
nand \U$39686 ( \40063 , \39986 , \40062 );
nand \U$39687 ( \40064 , \39985 , \40063 );
xor \U$39688 ( \40065 , \39845 , \40064 );
and \U$39689 ( \40066 , \39142 , \8020 );
not \U$39690 ( \40067 , \39142 );
and \U$39691 ( \40068 , \40067 , \8019 );
nor \U$39692 ( \40069 , \40066 , \40068 );
not \U$39693 ( \40070 , \40069 );
not \U$39694 ( \40071 , \39131 );
and \U$39695 ( \40072 , \40070 , \40071 );
and \U$39696 ( \40073 , \40069 , \39131 );
nor \U$39697 ( \40074 , \40072 , \40073 );
xor \U$39698 ( \40075 , \39659 , \39661 );
xor \U$39699 ( \40076 , \40075 , \39664 );
xor \U$39700 ( \40077 , \40074 , \40076 );
xor \U$39701 ( \40078 , \39691 , \39693 );
xor \U$39702 ( \40079 , \40078 , \39696 );
and \U$39703 ( \40080 , \40077 , \40079 );
and \U$39704 ( \40081 , \40074 , \40076 );
nor \U$39705 ( \40082 , \40080 , \40081 );
and \U$39706 ( \40083 , \40065 , \40082 );
and \U$39707 ( \40084 , \39845 , \40064 );
or \U$39708 ( \40085 , \40083 , \40084 );
nand \U$39709 ( \40086 , \39815 , \40085 );
nand \U$39710 ( \40087 , \39812 , \40086 );
xnor \U$39711 ( \40088 , \39701 , \39649 );
not \U$39712 ( \40089 , \40088 );
not \U$39713 ( \40090 , \39719 );
and \U$39714 ( \40091 , \40089 , \40090 );
and \U$39715 ( \40092 , \40088 , \39719 );
nor \U$39716 ( \40093 , \40091 , \40092 );
xnor \U$39717 ( \40094 , \39175 , \39257 );
not \U$39718 ( \40095 , \40094 );
not \U$39719 ( \40096 , \39318 );
and \U$39720 ( \40097 , \40095 , \40096 );
and \U$39721 ( \40098 , \40094 , \39318 );
nor \U$39722 ( \40099 , \40097 , \40098 );
or \U$39723 ( \40100 , \40093 , \40099 );
not \U$39724 ( \40101 , \40099 );
not \U$39725 ( \40102 , \40093 );
or \U$39726 ( \40103 , \40101 , \40102 );
xor \U$39727 ( \40104 , \39083 , \39085 );
xor \U$39728 ( \40105 , \40104 , \39096 );
xor \U$39729 ( \40106 , \39728 , \39735 );
xor \U$39730 ( \40107 , \40105 , \40106 );
nand \U$39731 ( \40108 , \40103 , \40107 );
nand \U$39732 ( \40109 , \40100 , \40108 );
xor \U$39733 ( \40110 , \40087 , \40109 );
xor \U$39734 ( \40111 , \39099 , \39320 );
xor \U$39735 ( \40112 , \40111 , \39335 );
xor \U$39736 ( \40113 , \39413 , \39418 );
xor \U$39737 ( \40114 , \40112 , \40113 );
and \U$39738 ( \40115 , \40110 , \40114 );
and \U$39739 ( \40116 , \40087 , \40109 );
or \U$39740 ( \40117 , \40115 , \40116 );
and \U$39741 ( \40118 , \39770 , \40117 );
and \U$39742 ( \40119 , \39767 , \39769 );
nor \U$39743 ( \40120 , \40118 , \40119 );
not \U$39744 ( \40121 , \40120 );
xor \U$39745 ( \40122 , \39751 , \39752 );
xor \U$39746 ( \40123 , \40122 , \39755 );
nand \U$39747 ( \40124 , \40121 , \40123 );
or \U$39748 ( \40125 , \39765 , \40124 );
not \U$39749 ( \40126 , \39764 );
not \U$39750 ( \40127 , \40124 );
and \U$39751 ( \40128 , \40126 , \40127 );
and \U$39752 ( \40129 , \39764 , \40124 );
nor \U$39753 ( \40130 , \40128 , \40129 );
not \U$39754 ( \40131 , \40120 );
not \U$39755 ( \40132 , \40123 );
or \U$39756 ( \40133 , \40131 , \40132 );
or \U$39757 ( \40134 , \40123 , \40120 );
nand \U$39758 ( \40135 , \40133 , \40134 );
xor \U$39759 ( \40136 , \39767 , \39769 );
xor \U$39760 ( \40137 , \40136 , \40117 );
not \U$39761 ( \40138 , \40137 );
xor \U$39762 ( \40139 , \40087 , \40109 );
xor \U$39763 ( \40140 , \40139 , \40114 );
xor \U$39764 ( \40141 , \39721 , \39723 );
xor \U$39765 ( \40142 , \40141 , \39740 );
and \U$39766 ( \40143 , \40140 , \40142 );
not \U$39767 ( \40144 , \40140 );
not \U$39768 ( \40145 , \40142 );
and \U$39769 ( \40146 , \40144 , \40145 );
not \U$39770 ( \40147 , \39794 );
not \U$39771 ( \40148 , \39792 );
not \U$39772 ( \40149 , \39809 );
or \U$39773 ( \40150 , \40148 , \40149 );
or \U$39774 ( \40151 , \39809 , \39792 );
nand \U$39775 ( \40152 , \40150 , \40151 );
not \U$39776 ( \40153 , \40152 );
or \U$39777 ( \40154 , \40147 , \40153 );
or \U$39778 ( \40155 , \40152 , \39794 );
nand \U$39779 ( \40156 , \40154 , \40155 );
xor \U$39780 ( \40157 , \39845 , \40064 );
xor \U$39781 ( \40158 , \40157 , \40082 );
xor \U$39782 ( \40159 , \40156 , \40158 );
xor \U$39783 ( \40160 , \39776 , \39782 );
xor \U$39784 ( \40161 , \40160 , \39787 );
and \U$39785 ( \40162 , \40159 , \40161 );
and \U$39786 ( \40163 , \40156 , \40158 );
nor \U$39787 ( \40164 , \40162 , \40163 );
xor \U$39788 ( \40165 , \39927 , \39952 );
xor \U$39789 ( \40166 , \40165 , \39980 );
not \U$39790 ( \40167 , \40166 );
and \U$39791 ( \40168 , \39873 , \39899 );
nor \U$39792 ( \40169 , \40168 , \39900 );
not \U$39793 ( \40170 , \40169 );
and \U$39794 ( \40171 , \40167 , \40170 );
and \U$39795 ( \40172 , \40166 , \40169 );
xor \U$39796 ( \40173 , \40006 , \40033 );
xor \U$39797 ( \40174 , \40173 , \40059 );
nor \U$39798 ( \40175 , \40172 , \40174 );
nor \U$39799 ( \40176 , \40171 , \40175 );
xor \U$39800 ( \40177 , \39801 , \39803 );
xor \U$39801 ( \40178 , \40177 , \39806 );
and \U$39802 ( \40179 , \40176 , \40178 );
xor \U$39803 ( \40180 , \40074 , \40076 );
xor \U$39804 ( \40181 , \40180 , \40079 );
xor \U$39805 ( \40182 , \39801 , \39803 );
xor \U$39806 ( \40183 , \40182 , \39806 );
and \U$39807 ( \40184 , \40181 , \40183 );
and \U$39808 ( \40185 , \40176 , \40181 );
or \U$39809 ( \40186 , \40179 , \40184 , \40185 );
not \U$39810 ( \40187 , \40186 );
xnor \U$39811 ( \40188 , \39983 , \40062 );
not \U$39812 ( \40189 , \40188 );
not \U$39813 ( \40190 , \39901 );
and \U$39814 ( \40191 , \40189 , \40190 );
and \U$39815 ( \40192 , \40188 , \39901 );
nor \U$39816 ( \40193 , \40191 , \40192 );
not \U$39817 ( \40194 , \40193 );
xor \U$39818 ( \40195 , \39825 , \39831 );
xor \U$39819 ( \40196 , \40195 , \39842 );
nand \U$39820 ( \40197 , \40194 , \40196 );
not \U$39821 ( \40198 , \40197 );
and \U$39822 ( \40199 , \40187 , \40198 );
and \U$39823 ( \40200 , \40186 , \40197 );
not \U$39824 ( \40201 , RIae78170_104);
nor \U$39825 ( \40202 , \40201 , \491 );
xor \U$39826 ( \40203 , \39881 , \39888 );
xor \U$39827 ( \40204 , \40203 , \39896 );
and \U$39828 ( \40205 , \40202 , \40204 );
xor \U$39829 ( \40206 , \39853 , \39861 );
xor \U$39830 ( \40207 , \40206 , \39870 );
xor \U$39831 ( \40208 , \39881 , \39888 );
xor \U$39832 ( \40209 , \40208 , \39896 );
and \U$39833 ( \40210 , \40207 , \40209 );
and \U$39834 ( \40211 , \40202 , \40207 );
or \U$39835 ( \40212 , \40205 , \40210 , \40211 );
not \U$39836 ( \40213 , \40212 );
not \U$39837 ( \40214 , \40213 );
xor \U$39838 ( \40215 , \39934 , \39941 );
xor \U$39839 ( \40216 , \40215 , \39949 );
not \U$39840 ( \40217 , \40216 );
xor \U$39841 ( \40218 , \39961 , \39969 );
xor \U$39842 ( \40219 , \40218 , \39977 );
not \U$39843 ( \40220 , \40219 );
and \U$39844 ( \40221 , \40217 , \40220 );
and \U$39845 ( \40222 , \40219 , \40216 );
xor \U$39846 ( \40223 , \39909 , \39916 );
xor \U$39847 ( \40224 , \40223 , \39924 );
nor \U$39848 ( \40225 , \40222 , \40224 );
nor \U$39849 ( \40226 , \40221 , \40225 );
not \U$39850 ( \40227 , \40226 );
and \U$39851 ( \40228 , \40214 , \40227 );
and \U$39852 ( \40229 , \40226 , \40213 );
not \U$39853 ( \40230 , \39993 );
and \U$39854 ( \40231 , \40004 , \8789 );
not \U$39855 ( \40232 , \40004 );
and \U$39856 ( \40233 , \40232 , \8799 );
nor \U$39857 ( \40234 , \40231 , \40233 );
not \U$39858 ( \40235 , \40234 );
or \U$39859 ( \40236 , \40230 , \40235 );
or \U$39860 ( \40237 , \40234 , \39993 );
nand \U$39861 ( \40238 , \40236 , \40237 );
xor \U$39862 ( \40239 , \40041 , \40048 );
xor \U$39863 ( \40240 , \40239 , \40056 );
xor \U$39864 ( \40241 , \40238 , \40240 );
not \U$39865 ( \40242 , \40013 );
xor \U$39866 ( \40243 , \40031 , \40021 );
not \U$39867 ( \40244 , \40243 );
or \U$39868 ( \40245 , \40242 , \40244 );
or \U$39869 ( \40246 , \40243 , \40013 );
nand \U$39870 ( \40247 , \40245 , \40246 );
and \U$39871 ( \40248 , \40241 , \40247 );
and \U$39872 ( \40249 , \40238 , \40240 );
nor \U$39873 ( \40250 , \40248 , \40249 );
nor \U$39874 ( \40251 , \40229 , \40250 );
nor \U$39875 ( \40252 , \40228 , \40251 );
and \U$39876 ( \40253 , \6941 , RIae76a00_54);
and \U$39877 ( \40254 , RIae76820_50, \6939 );
nor \U$39878 ( \40255 , \40253 , \40254 );
and \U$39879 ( \40256 , \40255 , \6314 );
not \U$39880 ( \40257 , \40255 );
and \U$39881 ( \40258 , \40257 , \6945 );
nor \U$39882 ( \40259 , \40256 , \40258 );
and \U$39883 ( \40260 , \5896 , RIae760a0_34);
and \U$39884 ( \40261 , RIae76370_40, \5894 );
nor \U$39885 ( \40262 , \40260 , \40261 );
and \U$39886 ( \40263 , \40262 , \5590 );
not \U$39887 ( \40264 , \40262 );
and \U$39888 ( \40265 , \40264 , \5589 );
nor \U$39889 ( \40266 , \40263 , \40265 );
xor \U$39890 ( \40267 , \40259 , \40266 );
and \U$39891 ( \40268 , \6172 , RIae76280_38);
and \U$39892 ( \40269 , RIae76af0_56, \6170 );
nor \U$39893 ( \40270 , \40268 , \40269 );
and \U$39894 ( \40271 , \40270 , \6176 );
not \U$39895 ( \40272 , \40270 );
and \U$39896 ( \40273 , \40272 , \6175 );
nor \U$39897 ( \40274 , \40271 , \40273 );
and \U$39898 ( \40275 , \40267 , \40274 );
and \U$39899 ( \40276 , \40259 , \40266 );
or \U$39900 ( \40277 , \40275 , \40276 );
and \U$39901 ( \40278 , \4247 , RIae75470_8);
and \U$39902 ( \40279 , RIae76460_42, \4245 );
nor \U$39903 ( \40280 , \40278 , \40279 );
and \U$39904 ( \40281 , \40280 , \3989 );
not \U$39905 ( \40282 , \40280 );
and \U$39906 ( \40283 , \40282 , \4251 );
nor \U$39907 ( \40284 , \40281 , \40283 );
and \U$39908 ( \40285 , \4688 , RIae76550_44);
and \U$39909 ( \40286 , RIae76730_48, \4686 );
nor \U$39910 ( \40287 , \40285 , \40286 );
and \U$39911 ( \40288 , \40287 , \4481 );
not \U$39912 ( \40289 , \40287 );
and \U$39913 ( \40290 , \40289 , \4482 );
nor \U$39914 ( \40291 , \40288 , \40290 );
xor \U$39915 ( \40292 , \40284 , \40291 );
and \U$39916 ( \40293 , \5399 , RIae76640_46);
and \U$39917 ( \40294 , RIae76190_36, \5397 );
nor \U$39918 ( \40295 , \40293 , \40294 );
and \U$39919 ( \40296 , \40295 , \5016 );
not \U$39920 ( \40297 , \40295 );
and \U$39921 ( \40298 , \40297 , \5403 );
nor \U$39922 ( \40299 , \40296 , \40298 );
and \U$39923 ( \40300 , \40292 , \40299 );
and \U$39924 ( \40301 , \40284 , \40291 );
or \U$39925 ( \40302 , \40300 , \40301 );
xor \U$39926 ( \40303 , \40277 , \40302 );
and \U$39927 ( \40304 , \7633 , RIae76910_52);
and \U$39928 ( \40305 , RIae76be0_58, \7631 );
nor \U$39929 ( \40306 , \40304 , \40305 );
and \U$39930 ( \40307 , \40306 , \7206 );
not \U$39931 ( \40308 , \40306 );
and \U$39932 ( \40309 , \40308 , \7205 );
nor \U$39933 ( \40310 , \40307 , \40309 );
nand \U$39934 ( \40311 , RIae78e18_131, \8966 );
and \U$39935 ( \40312 , \40311 , \8799 );
not \U$39936 ( \40313 , \40311 );
and \U$39937 ( \40314 , \40313 , \8789 );
nor \U$39938 ( \40315 , \40312 , \40314 );
xor \U$39939 ( \40316 , \40310 , \40315 );
and \U$39940 ( \40317 , \8371 , RIae78ad0_124);
and \U$39941 ( \40318 , RIae78d28_129, \8369 );
nor \U$39942 ( \40319 , \40317 , \40318 );
and \U$39943 ( \40320 , \40319 , \8020 );
not \U$39944 ( \40321 , \40319 );
and \U$39945 ( \40322 , \40321 , \8019 );
nor \U$39946 ( \40323 , \40320 , \40322 );
and \U$39947 ( \40324 , \40316 , \40323 );
and \U$39948 ( \40325 , \40310 , \40315 );
or \U$39949 ( \40326 , \40324 , \40325 );
and \U$39950 ( \40327 , \40303 , \40326 );
and \U$39951 ( \40328 , \40277 , \40302 );
nor \U$39952 ( \40329 , \40327 , \40328 );
not \U$39953 ( \40330 , \40329 );
not \U$39954 ( \40331 , \3089 );
and \U$39955 ( \40332 , \2783 , RIae75560_10);
and \U$39956 ( \40333 , RIae75830_16, \2781 );
nor \U$39957 ( \40334 , \40332 , \40333 );
not \U$39958 ( \40335 , \40334 );
or \U$39959 ( \40336 , \40331 , \40335 );
or \U$39960 ( \40337 , \40334 , \3089 );
nand \U$39961 ( \40338 , \40336 , \40337 );
not \U$39962 ( \40339 , \2774 );
and \U$39963 ( \40340 , \3214 , RIae75740_14);
and \U$39964 ( \40341 , RIae75290_4, \3212 );
nor \U$39965 ( \40342 , \40340 , \40341 );
not \U$39966 ( \40343 , \40342 );
or \U$39967 ( \40344 , \40339 , \40343 );
or \U$39968 ( \40345 , \40342 , \3218 );
nand \U$39969 ( \40346 , \40344 , \40345 );
xor \U$39970 ( \40347 , \40338 , \40346 );
and \U$39971 ( \40348 , \3730 , RIae751a0_2);
and \U$39972 ( \40349 , RIae75380_6, \3728 );
nor \U$39973 ( \40350 , \40348 , \40349 );
and \U$39974 ( \40351 , \40350 , \3732 );
not \U$39975 ( \40352 , \40350 );
and \U$39976 ( \40353 , \40352 , \3422 );
nor \U$39977 ( \40354 , \40351 , \40353 );
and \U$39978 ( \40355 , \40347 , \40354 );
and \U$39979 ( \40356 , \40338 , \40346 );
or \U$39980 ( \40357 , \40355 , \40356 );
and \U$39981 ( \40358 , \1939 , RIae75920_18);
and \U$39982 ( \40359 , RIae75fb0_32, \1937 );
nor \U$39983 ( \40360 , \40358 , \40359 );
and \U$39984 ( \40361 , \40360 , \1735 );
not \U$39985 ( \40362 , \40360 );
and \U$39986 ( \40363 , \40362 , \1734 );
nor \U$39987 ( \40364 , \40361 , \40363 );
and \U$39988 ( \40365 , \2224 , RIae75ec0_30);
and \U$39989 ( \40366 , RIae75ce0_26, \2222 );
nor \U$39990 ( \40367 , \40365 , \40366 );
and \U$39991 ( \40368 , \40367 , \2061 );
not \U$39992 ( \40369 , \40367 );
and \U$39993 ( \40370 , \40369 , \2060 );
nor \U$39994 ( \40371 , \40368 , \40370 );
xor \U$39995 ( \40372 , \40364 , \40371 );
and \U$39996 ( \40373 , \2607 , RIae75dd0_28);
and \U$39997 ( \40374 , RIae75650_12, \2605 );
nor \U$39998 ( \40375 , \40373 , \40374 );
and \U$39999 ( \40376 , \40375 , \2611 );
not \U$40000 ( \40377 , \40375 );
and \U$40001 ( \40378 , \40377 , \2397 );
nor \U$40002 ( \40379 , \40376 , \40378 );
and \U$40003 ( \40380 , \40372 , \40379 );
and \U$40004 ( \40381 , \40364 , \40371 );
or \U$40005 ( \40382 , \40380 , \40381 );
xor \U$40006 ( \40383 , \40357 , \40382 );
and \U$40007 ( \40384 , \1593 , RIae75b00_22);
and \U$40008 ( \40385 , RIae75a10_20, \1591 );
nor \U$40009 ( \40386 , \40384 , \40385 );
and \U$40010 ( \40387 , \40386 , \1498 );
not \U$40011 ( \40388 , \40386 );
and \U$40012 ( \40389 , \40388 , \1488 );
nor \U$40013 ( \40390 , \40387 , \40389 );
and \U$40014 ( \40391 , \1138 , RIae788f0_120);
and \U$40015 ( \40392 , RIae78800_118, \1136 );
nor \U$40016 ( \40393 , \40391 , \40392 );
and \U$40017 ( \40394 , \40393 , \1012 );
not \U$40018 ( \40395 , \40393 );
and \U$40019 ( \40396 , \40395 , \1142 );
nor \U$40020 ( \40397 , \40394 , \40396 );
xor \U$40021 ( \40398 , \40390 , \40397 );
and \U$40022 ( \40399 , \1376 , RIae78710_116);
and \U$40023 ( \40400 , RIae75bf0_24, \1374 );
nor \U$40024 ( \40401 , \40399 , \40400 );
and \U$40025 ( \40402 , \40401 , \1380 );
not \U$40026 ( \40403 , \40401 );
and \U$40027 ( \40404 , \40403 , \1261 );
nor \U$40028 ( \40405 , \40402 , \40404 );
and \U$40029 ( \40406 , \40398 , \40405 );
and \U$40030 ( \40407 , \40390 , \40397 );
or \U$40031 ( \40408 , \40406 , \40407 );
and \U$40032 ( \40409 , \40383 , \40408 );
and \U$40033 ( \40410 , \40357 , \40382 );
nor \U$40034 ( \40411 , \40409 , \40410 );
not \U$40035 ( \40412 , \40411 );
and \U$40036 ( \40413 , \40330 , \40412 );
and \U$40037 ( \40414 , \40329 , \40411 );
and \U$40038 ( \40415 , \384 , RIae78170_104);
and \U$40039 ( \40416 , RIae77f90_100, \382 );
nor \U$40040 ( \40417 , \40415 , \40416 );
not \U$40041 ( \40418 , \40417 );
not \U$40042 ( \40419 , \388 );
and \U$40043 ( \40420 , \40418 , \40419 );
and \U$40044 ( \40421 , \40417 , \392 );
nor \U$40045 ( \40422 , \40420 , \40421 );
not \U$40046 ( \40423 , \40422 );
and \U$40047 ( \40424 , \514 , RIae78620_114);
and \U$40048 ( \40425 , RIae78440_110, \512 );
nor \U$40049 ( \40426 , \40424 , \40425 );
not \U$40050 ( \40427 , \40426 );
not \U$40051 ( \40428 , \471 );
and \U$40052 ( \40429 , \40427 , \40428 );
and \U$40053 ( \40430 , \40426 , \469 );
nor \U$40054 ( \40431 , \40429 , \40430 );
not \U$40055 ( \40432 , \40431 );
and \U$40056 ( \40433 , \40423 , \40432 );
and \U$40057 ( \40434 , \40431 , \40422 );
and \U$40058 ( \40435 , \436 , RIae78080_102);
and \U$40059 ( \40436 , RIae78260_106, \434 );
nor \U$40060 ( \40437 , \40435 , \40436 );
not \U$40061 ( \40438 , \40437 );
not \U$40062 ( \40439 , \400 );
and \U$40063 ( \40440 , \40438 , \40439 );
and \U$40064 ( \40441 , \40437 , \402 );
nor \U$40065 ( \40442 , \40440 , \40441 );
nor \U$40066 ( \40443 , \40434 , \40442 );
nor \U$40067 ( \40444 , \40433 , \40443 );
not \U$40068 ( \40445 , \40444 );
nand \U$40069 ( \40446 , RIae78350_108, RIae78b48_125);
not \U$40070 ( \40447 , \40446 );
and \U$40071 ( \40448 , \40445 , \40447 );
and \U$40072 ( \40449 , \40444 , \40446 );
and \U$40073 ( \40450 , \558 , RIae784b8_111);
and \U$40074 ( \40451 , RIae77cc0_94, \556 );
nor \U$40075 ( \40452 , \40450 , \40451 );
and \U$40076 ( \40453 , \40452 , \504 );
not \U$40077 ( \40454 , \40452 );
and \U$40078 ( \40455 , \40454 , \562 );
nor \U$40079 ( \40456 , \40453 , \40455 );
and \U$40080 ( \40457 , \672 , RIae77bd0_92);
and \U$40081 ( \40458 , RIae77db0_96, \670 );
nor \U$40082 ( \40459 , \40457 , \40458 );
and \U$40083 ( \40460 , \40459 , \588 );
not \U$40084 ( \40461 , \40459 );
and \U$40085 ( \40462 , \40461 , \587 );
nor \U$40086 ( \40463 , \40460 , \40462 );
xor \U$40087 ( \40464 , \40456 , \40463 );
not \U$40088 ( \40465 , \789 );
and \U$40089 ( \40466 , \883 , RIae77ea0_98);
and \U$40090 ( \40467 , RIae789e0_122, \881 );
nor \U$40091 ( \40468 , \40466 , \40467 );
not \U$40092 ( \40469 , \40468 );
or \U$40093 ( \40470 , \40465 , \40469 );
or \U$40094 ( \40471 , \40468 , \787 );
nand \U$40095 ( \40472 , \40470 , \40471 );
and \U$40096 ( \40473 , \40464 , \40472 );
and \U$40097 ( \40474 , \40456 , \40463 );
or \U$40098 ( \40475 , \40473 , \40474 );
not \U$40099 ( \40476 , \40475 );
nor \U$40100 ( \40477 , \40449 , \40476 );
nor \U$40101 ( \40478 , \40448 , \40477 );
nor \U$40102 ( \40479 , \40414 , \40478 );
nor \U$40103 ( \40480 , \40413 , \40479 );
xor \U$40104 ( \40481 , \40252 , \40480 );
xor \U$40105 ( \40482 , \39834 , \39836 );
xor \U$40106 ( \40483 , \40482 , \39839 );
not \U$40107 ( \40484 , \40483 );
not \U$40108 ( \40485 , \39830 );
not \U$40109 ( \40486 , \39827 );
and \U$40110 ( \40487 , \40485 , \40486 );
and \U$40111 ( \40488 , \39830 , \39827 );
nor \U$40112 ( \40489 , \40487 , \40488 );
not \U$40113 ( \40490 , \40489 );
and \U$40114 ( \40491 , \40484 , \40490 );
and \U$40115 ( \40492 , \40483 , \40489 );
xor \U$40116 ( \40493 , \39817 , \39819 );
xor \U$40117 ( \40494 , \40493 , \39822 );
nor \U$40118 ( \40495 , \40492 , \40494 );
nor \U$40119 ( \40496 , \40491 , \40495 );
and \U$40120 ( \40497 , \40481 , \40496 );
and \U$40121 ( \40498 , \40252 , \40480 );
or \U$40122 ( \40499 , \40497 , \40498 );
nor \U$40123 ( \40500 , \40200 , \40499 );
nor \U$40124 ( \40501 , \40199 , \40500 );
xor \U$40125 ( \40502 , \40164 , \40501 );
xnor \U$40126 ( \40503 , \40099 , \40093 );
not \U$40127 ( \40504 , \40503 );
not \U$40128 ( \40505 , \40107 );
and \U$40129 ( \40506 , \40504 , \40505 );
and \U$40130 ( \40507 , \40503 , \40107 );
nor \U$40131 ( \40508 , \40506 , \40507 );
and \U$40132 ( \40509 , \40502 , \40508 );
and \U$40133 ( \40510 , \40164 , \40501 );
or \U$40134 ( \40511 , \40509 , \40510 );
nor \U$40135 ( \40512 , \40146 , \40511 );
nor \U$40136 ( \40513 , \40143 , \40512 );
nor \U$40137 ( \40514 , \40138 , \40513 );
and \U$40138 ( \40515 , \40135 , \40514 );
xor \U$40139 ( \40516 , \40514 , \40135 );
not \U$40140 ( \40517 , \40137 );
not \U$40141 ( \40518 , \40513 );
and \U$40142 ( \40519 , \40517 , \40518 );
and \U$40143 ( \40520 , \40137 , \40513 );
nor \U$40144 ( \40521 , \40519 , \40520 );
xor \U$40145 ( \40522 , \40156 , \40158 );
xor \U$40146 ( \40523 , \40522 , \40161 );
xor \U$40147 ( \40524 , \40310 , \40315 );
xor \U$40148 ( \40525 , \40524 , \40323 );
xor \U$40149 ( \40526 , \40259 , \40266 );
xor \U$40150 ( \40527 , \40526 , \40274 );
and \U$40151 ( \40528 , \40525 , \40527 );
xor \U$40152 ( \40529 , \40284 , \40291 );
xor \U$40153 ( \40530 , \40529 , \40299 );
xor \U$40154 ( \40531 , \40259 , \40266 );
xor \U$40155 ( \40532 , \40531 , \40274 );
and \U$40156 ( \40533 , \40530 , \40532 );
and \U$40157 ( \40534 , \40525 , \40530 );
or \U$40158 ( \40535 , \40528 , \40533 , \40534 );
xor \U$40159 ( \40536 , \40456 , \40463 );
xor \U$40160 ( \40537 , \40536 , \40472 );
xor \U$40161 ( \40538 , \40537 , \40446 );
not \U$40162 ( \40539 , \40422 );
xor \U$40163 ( \40540 , \40442 , \40431 );
not \U$40164 ( \40541 , \40540 );
or \U$40165 ( \40542 , \40539 , \40541 );
or \U$40166 ( \40543 , \40540 , \40422 );
nand \U$40167 ( \40544 , \40542 , \40543 );
and \U$40168 ( \40545 , \40538 , \40544 );
and \U$40169 ( \40546 , \40537 , \40446 );
or \U$40170 ( \40547 , \40545 , \40546 );
xor \U$40171 ( \40548 , \40535 , \40547 );
xor \U$40172 ( \40549 , \40390 , \40397 );
xor \U$40173 ( \40550 , \40549 , \40405 );
xor \U$40174 ( \40551 , \40364 , \40371 );
xor \U$40175 ( \40552 , \40551 , \40379 );
and \U$40176 ( \40553 , \40550 , \40552 );
xor \U$40177 ( \40554 , \40338 , \40346 );
xor \U$40178 ( \40555 , \40554 , \40354 );
xor \U$40179 ( \40556 , \40364 , \40371 );
xor \U$40180 ( \40557 , \40556 , \40379 );
and \U$40181 ( \40558 , \40555 , \40557 );
and \U$40182 ( \40559 , \40550 , \40555 );
or \U$40183 ( \40560 , \40553 , \40558 , \40559 );
and \U$40184 ( \40561 , \40548 , \40560 );
and \U$40185 ( \40562 , \40535 , \40547 );
or \U$40186 ( \40563 , \40561 , \40562 );
and \U$40187 ( \40564 , \5896 , RIae76190_36);
and \U$40188 ( \40565 , RIae760a0_34, \5894 );
nor \U$40189 ( \40566 , \40564 , \40565 );
and \U$40190 ( \40567 , \40566 , \5590 );
not \U$40191 ( \40568 , \40566 );
and \U$40192 ( \40569 , \40568 , \5589 );
nor \U$40193 ( \40570 , \40567 , \40569 );
and \U$40194 ( \40571 , \4688 , RIae76460_42);
and \U$40195 ( \40572 , RIae76550_44, \4686 );
nor \U$40196 ( \40573 , \40571 , \40572 );
and \U$40197 ( \40574 , \40573 , \4481 );
not \U$40198 ( \40575 , \40573 );
and \U$40199 ( \40576 , \40575 , \4482 );
nor \U$40200 ( \40577 , \40574 , \40576 );
xor \U$40201 ( \40578 , \40570 , \40577 );
and \U$40202 ( \40579 , \5399 , RIae76730_48);
and \U$40203 ( \40580 , RIae76640_46, \5397 );
nor \U$40204 ( \40581 , \40579 , \40580 );
and \U$40205 ( \40582 , \40581 , \5016 );
not \U$40206 ( \40583 , \40581 );
and \U$40207 ( \40584 , \40583 , \5403 );
nor \U$40208 ( \40585 , \40582 , \40584 );
and \U$40209 ( \40586 , \40578 , \40585 );
and \U$40210 ( \40587 , \40570 , \40577 );
or \U$40211 ( \40588 , \40586 , \40587 );
and \U$40212 ( \40589 , \8966 , RIae78d28_129);
and \U$40213 ( \40590 , RIae78e18_131, \8964 );
nor \U$40214 ( \40591 , \40589 , \40590 );
and \U$40215 ( \40592 , \40591 , \8799 );
not \U$40216 ( \40593 , \40591 );
and \U$40217 ( \40594 , \40593 , \8789 );
nor \U$40218 ( \40595 , \40592 , \40594 );
xor \U$40219 ( \40596 , \40595 , \9273 );
and \U$40220 ( \40597 , \8371 , RIae76be0_58);
and \U$40221 ( \40598 , RIae78ad0_124, \8369 );
nor \U$40222 ( \40599 , \40597 , \40598 );
and \U$40223 ( \40600 , \40599 , \8020 );
not \U$40224 ( \40601 , \40599 );
and \U$40225 ( \40602 , \40601 , \8019 );
nor \U$40226 ( \40603 , \40600 , \40602 );
and \U$40227 ( \40604 , \40596 , \40603 );
and \U$40228 ( \40605 , \40595 , \9273 );
or \U$40229 ( \40606 , \40604 , \40605 );
xor \U$40230 ( \40607 , \40588 , \40606 );
and \U$40231 ( \40608 , \7633 , RIae76820_50);
and \U$40232 ( \40609 , RIae76910_52, \7631 );
nor \U$40233 ( \40610 , \40608 , \40609 );
and \U$40234 ( \40611 , \40610 , \7206 );
not \U$40235 ( \40612 , \40610 );
and \U$40236 ( \40613 , \40612 , \7205 );
nor \U$40237 ( \40614 , \40611 , \40613 );
and \U$40238 ( \40615 , \6172 , RIae76370_40);
and \U$40239 ( \40616 , RIae76280_38, \6170 );
nor \U$40240 ( \40617 , \40615 , \40616 );
and \U$40241 ( \40618 , \40617 , \6176 );
not \U$40242 ( \40619 , \40617 );
and \U$40243 ( \40620 , \40619 , \6175 );
nor \U$40244 ( \40621 , \40618 , \40620 );
xor \U$40245 ( \40622 , \40614 , \40621 );
and \U$40246 ( \40623 , \6941 , RIae76af0_56);
and \U$40247 ( \40624 , RIae76a00_54, \6939 );
nor \U$40248 ( \40625 , \40623 , \40624 );
and \U$40249 ( \40626 , \40625 , \6314 );
not \U$40250 ( \40627 , \40625 );
and \U$40251 ( \40628 , \40627 , \6945 );
nor \U$40252 ( \40629 , \40626 , \40628 );
and \U$40253 ( \40630 , \40622 , \40629 );
and \U$40254 ( \40631 , \40614 , \40621 );
or \U$40255 ( \40632 , \40630 , \40631 );
and \U$40256 ( \40633 , \40607 , \40632 );
and \U$40257 ( \40634 , \40588 , \40606 );
or \U$40258 ( \40635 , \40633 , \40634 );
and \U$40259 ( \40636 , \1138 , RIae789e0_122);
and \U$40260 ( \40637 , RIae788f0_120, \1136 );
nor \U$40261 ( \40638 , \40636 , \40637 );
and \U$40262 ( \40639 , \40638 , \1012 );
not \U$40263 ( \40640 , \40638 );
and \U$40264 ( \40641 , \40640 , \1142 );
nor \U$40265 ( \40642 , \40639 , \40641 );
and \U$40266 ( \40643 , \672 , RIae77cc0_94);
and \U$40267 ( \40644 , RIae77bd0_92, \670 );
nor \U$40268 ( \40645 , \40643 , \40644 );
and \U$40269 ( \40646 , \40645 , \588 );
not \U$40270 ( \40647 , \40645 );
and \U$40271 ( \40648 , \40647 , \587 );
nor \U$40272 ( \40649 , \40646 , \40648 );
xor \U$40273 ( \40650 , \40642 , \40649 );
not \U$40274 ( \40651 , \789 );
and \U$40275 ( \40652 , \883 , RIae77db0_96);
and \U$40276 ( \40653 , RIae77ea0_98, \881 );
nor \U$40277 ( \40654 , \40652 , \40653 );
not \U$40278 ( \40655 , \40654 );
or \U$40279 ( \40656 , \40651 , \40655 );
or \U$40280 ( \40657 , \40654 , \787 );
nand \U$40281 ( \40658 , \40656 , \40657 );
and \U$40282 ( \40659 , \40650 , \40658 );
and \U$40283 ( \40660 , \40642 , \40649 );
or \U$40284 ( \40661 , \40659 , \40660 );
not \U$40285 ( \40662 , RIae77360_74);
nor \U$40286 ( \40663 , \40662 , \491 );
not \U$40287 ( \40664 , \388 );
and \U$40288 ( \40665 , \384 , RIae78350_108);
and \U$40289 ( \40666 , RIae78170_104, \382 );
nor \U$40290 ( \40667 , \40665 , \40666 );
not \U$40291 ( \40668 , \40667 );
or \U$40292 ( \40669 , \40664 , \40668 );
or \U$40293 ( \40670 , \40667 , \392 );
nand \U$40294 ( \40671 , \40669 , \40670 );
and \U$40295 ( \40672 , \40663 , \40671 );
xor \U$40296 ( \40673 , \40661 , \40672 );
not \U$40297 ( \40674 , \402 );
and \U$40298 ( \40675 , \436 , RIae77f90_100);
and \U$40299 ( \40676 , RIae78080_102, \434 );
nor \U$40300 ( \40677 , \40675 , \40676 );
not \U$40301 ( \40678 , \40677 );
or \U$40302 ( \40679 , \40674 , \40678 );
or \U$40303 ( \40680 , \40677 , \402 );
nand \U$40304 ( \40681 , \40679 , \40680 );
not \U$40305 ( \40682 , \471 );
and \U$40306 ( \40683 , \514 , RIae78260_106);
and \U$40307 ( \40684 , RIae78620_114, \512 );
nor \U$40308 ( \40685 , \40683 , \40684 );
not \U$40309 ( \40686 , \40685 );
or \U$40310 ( \40687 , \40682 , \40686 );
or \U$40311 ( \40688 , \40685 , \469 );
nand \U$40312 ( \40689 , \40687 , \40688 );
xor \U$40313 ( \40690 , \40681 , \40689 );
and \U$40314 ( \40691 , \558 , RIae78440_110);
and \U$40315 ( \40692 , RIae784b8_111, \556 );
nor \U$40316 ( \40693 , \40691 , \40692 );
and \U$40317 ( \40694 , \40693 , \504 );
not \U$40318 ( \40695 , \40693 );
and \U$40319 ( \40696 , \40695 , \562 );
nor \U$40320 ( \40697 , \40694 , \40696 );
and \U$40321 ( \40698 , \40690 , \40697 );
and \U$40322 ( \40699 , \40681 , \40689 );
or \U$40323 ( \40700 , \40698 , \40699 );
and \U$40324 ( \40701 , \40673 , \40700 );
and \U$40325 ( \40702 , \40661 , \40672 );
or \U$40326 ( \40703 , \40701 , \40702 );
xor \U$40327 ( \40704 , \40635 , \40703 );
not \U$40328 ( \40705 , \2789 );
and \U$40329 ( \40706 , \2783 , RIae75650_12);
and \U$40330 ( \40707 , RIae75560_10, \2781 );
nor \U$40331 ( \40708 , \40706 , \40707 );
not \U$40332 ( \40709 , \40708 );
or \U$40333 ( \40710 , \40705 , \40709 );
or \U$40334 ( \40711 , \40708 , \3089 );
nand \U$40335 ( \40712 , \40710 , \40711 );
and \U$40336 ( \40713 , \2224 , RIae75fb0_32);
and \U$40337 ( \40714 , RIae75ec0_30, \2222 );
nor \U$40338 ( \40715 , \40713 , \40714 );
and \U$40339 ( \40716 , \40715 , \2061 );
not \U$40340 ( \40717 , \40715 );
and \U$40341 ( \40718 , \40717 , \2060 );
nor \U$40342 ( \40719 , \40716 , \40718 );
xor \U$40343 ( \40720 , \40712 , \40719 );
and \U$40344 ( \40721 , \2607 , RIae75ce0_26);
and \U$40345 ( \40722 , RIae75dd0_28, \2605 );
nor \U$40346 ( \40723 , \40721 , \40722 );
and \U$40347 ( \40724 , \40723 , \2611 );
not \U$40348 ( \40725 , \40723 );
and \U$40349 ( \40726 , \40725 , \2397 );
nor \U$40350 ( \40727 , \40724 , \40726 );
and \U$40351 ( \40728 , \40720 , \40727 );
and \U$40352 ( \40729 , \40712 , \40719 );
or \U$40353 ( \40730 , \40728 , \40729 );
and \U$40354 ( \40731 , \1376 , RIae78800_118);
and \U$40355 ( \40732 , RIae78710_116, \1374 );
nor \U$40356 ( \40733 , \40731 , \40732 );
and \U$40357 ( \40734 , \40733 , \1380 );
not \U$40358 ( \40735 , \40733 );
and \U$40359 ( \40736 , \40735 , \1261 );
nor \U$40360 ( \40737 , \40734 , \40736 );
and \U$40361 ( \40738 , \1593 , RIae75bf0_24);
and \U$40362 ( \40739 , RIae75b00_22, \1591 );
nor \U$40363 ( \40740 , \40738 , \40739 );
and \U$40364 ( \40741 , \40740 , \1498 );
not \U$40365 ( \40742 , \40740 );
and \U$40366 ( \40743 , \40742 , \1488 );
nor \U$40367 ( \40744 , \40741 , \40743 );
xor \U$40368 ( \40745 , \40737 , \40744 );
and \U$40369 ( \40746 , \1939 , RIae75a10_20);
and \U$40370 ( \40747 , RIae75920_18, \1937 );
nor \U$40371 ( \40748 , \40746 , \40747 );
and \U$40372 ( \40749 , \40748 , \1735 );
not \U$40373 ( \40750 , \40748 );
and \U$40374 ( \40751 , \40750 , \1734 );
nor \U$40375 ( \40752 , \40749 , \40751 );
and \U$40376 ( \40753 , \40745 , \40752 );
and \U$40377 ( \40754 , \40737 , \40744 );
or \U$40378 ( \40755 , \40753 , \40754 );
xor \U$40379 ( \40756 , \40730 , \40755 );
not \U$40380 ( \40757 , \2774 );
and \U$40381 ( \40758 , \3214 , RIae75830_16);
and \U$40382 ( \40759 , RIae75740_14, \3212 );
nor \U$40383 ( \40760 , \40758 , \40759 );
not \U$40384 ( \40761 , \40760 );
or \U$40385 ( \40762 , \40757 , \40761 );
or \U$40386 ( \40763 , \40760 , \3218 );
nand \U$40387 ( \40764 , \40762 , \40763 );
and \U$40388 ( \40765 , \3730 , RIae75290_4);
and \U$40389 ( \40766 , RIae751a0_2, \3728 );
nor \U$40390 ( \40767 , \40765 , \40766 );
and \U$40391 ( \40768 , \40767 , \3732 );
not \U$40392 ( \40769 , \40767 );
and \U$40393 ( \40770 , \40769 , \3422 );
nor \U$40394 ( \40771 , \40768 , \40770 );
xor \U$40395 ( \40772 , \40764 , \40771 );
and \U$40396 ( \40773 , \4247 , RIae75380_6);
and \U$40397 ( \40774 , RIae75470_8, \4245 );
nor \U$40398 ( \40775 , \40773 , \40774 );
and \U$40399 ( \40776 , \40775 , \3989 );
not \U$40400 ( \40777 , \40775 );
and \U$40401 ( \40778 , \40777 , \4251 );
nor \U$40402 ( \40779 , \40776 , \40778 );
and \U$40403 ( \40780 , \40772 , \40779 );
and \U$40404 ( \40781 , \40764 , \40771 );
or \U$40405 ( \40782 , \40780 , \40781 );
and \U$40406 ( \40783 , \40756 , \40782 );
and \U$40407 ( \40784 , \40730 , \40755 );
or \U$40408 ( \40785 , \40783 , \40784 );
and \U$40409 ( \40786 , \40704 , \40785 );
and \U$40410 ( \40787 , \40635 , \40703 );
or \U$40411 ( \40788 , \40786 , \40787 );
xor \U$40412 ( \40789 , \40563 , \40788 );
xor \U$40413 ( \40790 , \40238 , \40240 );
xor \U$40414 ( \40791 , \40790 , \40247 );
xor \U$40415 ( \40792 , \39881 , \39888 );
xor \U$40416 ( \40793 , \40792 , \39896 );
xor \U$40417 ( \40794 , \40202 , \40207 );
xor \U$40418 ( \40795 , \40793 , \40794 );
xor \U$40419 ( \40796 , \40791 , \40795 );
not \U$40420 ( \40797 , \40219 );
xor \U$40421 ( \40798 , \40224 , \40216 );
not \U$40422 ( \40799 , \40798 );
or \U$40423 ( \40800 , \40797 , \40799 );
or \U$40424 ( \40801 , \40798 , \40219 );
nand \U$40425 ( \40802 , \40800 , \40801 );
and \U$40426 ( \40803 , \40796 , \40802 );
and \U$40427 ( \40804 , \40791 , \40795 );
or \U$40428 ( \40805 , \40803 , \40804 );
and \U$40429 ( \40806 , \40789 , \40805 );
and \U$40430 ( \40807 , \40563 , \40788 );
or \U$40431 ( \40808 , \40806 , \40807 );
not \U$40432 ( \40809 , \40329 );
xor \U$40433 ( \40810 , \40478 , \40411 );
not \U$40434 ( \40811 , \40810 );
or \U$40435 ( \40812 , \40809 , \40811 );
or \U$40436 ( \40813 , \40810 , \40329 );
nand \U$40437 ( \40814 , \40812 , \40813 );
not \U$40438 ( \40815 , \40213 );
xor \U$40439 ( \40816 , \40226 , \40250 );
not \U$40440 ( \40817 , \40816 );
or \U$40441 ( \40818 , \40815 , \40817 );
or \U$40442 ( \40819 , \40816 , \40213 );
nand \U$40443 ( \40820 , \40818 , \40819 );
and \U$40444 ( \40821 , \40814 , \40820 );
xor \U$40445 ( \40822 , \40808 , \40821 );
not \U$40446 ( \40823 , \40169 );
xor \U$40447 ( \40824 , \40174 , \40166 );
not \U$40448 ( \40825 , \40824 );
or \U$40449 ( \40826 , \40823 , \40825 );
or \U$40450 ( \40827 , \40824 , \40169 );
nand \U$40451 ( \40828 , \40826 , \40827 );
xor \U$40452 ( \40829 , \40357 , \40382 );
xor \U$40453 ( \40830 , \40829 , \40408 );
xor \U$40454 ( \40831 , \40277 , \40302 );
xor \U$40455 ( \40832 , \40831 , \40326 );
xor \U$40456 ( \40833 , \40830 , \40832 );
not \U$40457 ( \40834 , \40446 );
not \U$40458 ( \40835 , \40475 );
not \U$40459 ( \40836 , \40444 );
or \U$40460 ( \40837 , \40835 , \40836 );
or \U$40461 ( \40838 , \40444 , \40475 );
nand \U$40462 ( \40839 , \40837 , \40838 );
not \U$40463 ( \40840 , \40839 );
or \U$40464 ( \40841 , \40834 , \40840 );
or \U$40465 ( \40842 , \40839 , \40446 );
nand \U$40466 ( \40843 , \40841 , \40842 );
and \U$40467 ( \40844 , \40833 , \40843 );
and \U$40468 ( \40845 , \40830 , \40832 );
or \U$40469 ( \40846 , \40844 , \40845 );
xor \U$40470 ( \40847 , \40828 , \40846 );
not \U$40471 ( \40848 , \40489 );
xor \U$40472 ( \40849 , \40483 , \40494 );
not \U$40473 ( \40850 , \40849 );
or \U$40474 ( \40851 , \40848 , \40850 );
or \U$40475 ( \40852 , \40849 , \40489 );
nand \U$40476 ( \40853 , \40851 , \40852 );
and \U$40477 ( \40854 , \40847 , \40853 );
and \U$40478 ( \40855 , \40828 , \40846 );
or \U$40479 ( \40856 , \40854 , \40855 );
and \U$40480 ( \40857 , \40822 , \40856 );
and \U$40481 ( \40858 , \40808 , \40821 );
or \U$40482 ( \40859 , \40857 , \40858 );
and \U$40483 ( \40860 , \40523 , \40859 );
not \U$40484 ( \40861 , \40523 );
not \U$40485 ( \40862 , \40859 );
and \U$40486 ( \40863 , \40861 , \40862 );
not \U$40487 ( \40864 , \40196 );
not \U$40488 ( \40865 , \40193 );
and \U$40489 ( \40866 , \40864 , \40865 );
and \U$40490 ( \40867 , \40196 , \40193 );
nor \U$40491 ( \40868 , \40866 , \40867 );
xor \U$40492 ( \40869 , \40252 , \40480 );
xor \U$40493 ( \40870 , \40869 , \40496 );
and \U$40494 ( \40871 , \40868 , \40870 );
xor \U$40495 ( \40872 , \39801 , \39803 );
xor \U$40496 ( \40873 , \40872 , \39806 );
xor \U$40497 ( \40874 , \40176 , \40181 );
xor \U$40498 ( \40875 , \40873 , \40874 );
xor \U$40499 ( \40876 , \40252 , \40480 );
xor \U$40500 ( \40877 , \40876 , \40496 );
and \U$40501 ( \40878 , \40875 , \40877 );
and \U$40502 ( \40879 , \40868 , \40875 );
or \U$40503 ( \40880 , \40871 , \40878 , \40879 );
nor \U$40504 ( \40881 , \40863 , \40880 );
nor \U$40505 ( \40882 , \40860 , \40881 );
not \U$40506 ( \40883 , \39811 );
not \U$40507 ( \40884 , \40085 );
or \U$40508 ( \40885 , \40883 , \40884 );
or \U$40509 ( \40886 , \39811 , \40085 );
nand \U$40510 ( \40887 , \40885 , \40886 );
not \U$40511 ( \40888 , \40887 );
not \U$40512 ( \40889 , \39790 );
and \U$40513 ( \40890 , \40888 , \40889 );
and \U$40514 ( \40891 , \40887 , \39790 );
nor \U$40515 ( \40892 , \40890 , \40891 );
xor \U$40516 ( \40893 , \40882 , \40892 );
xor \U$40517 ( \40894 , \40164 , \40501 );
xor \U$40518 ( \40895 , \40894 , \40508 );
and \U$40519 ( \40896 , \40893 , \40895 );
and \U$40520 ( \40897 , \40882 , \40892 );
or \U$40521 ( \40898 , \40896 , \40897 );
not \U$40522 ( \40899 , \40898 );
not \U$40523 ( \40900 , \40140 );
not \U$40524 ( \40901 , \40511 );
not \U$40525 ( \40902 , \40142 );
and \U$40526 ( \40903 , \40901 , \40902 );
and \U$40527 ( \40904 , \40511 , \40142 );
nor \U$40528 ( \40905 , \40903 , \40904 );
not \U$40529 ( \40906 , \40905 );
or \U$40530 ( \40907 , \40900 , \40906 );
or \U$40531 ( \40908 , \40905 , \40140 );
nand \U$40532 ( \40909 , \40907 , \40908 );
nand \U$40533 ( \40910 , \40899 , \40909 );
or \U$40534 ( \40911 , \40521 , \40910 );
xnor \U$40535 ( \40912 , \40910 , \40521 );
xor \U$40536 ( \40913 , \40882 , \40892 );
xor \U$40537 ( \40914 , \40913 , \40895 );
not \U$40538 ( \40915 , \40914 );
not \U$40539 ( \40916 , \40197 );
xor \U$40540 ( \40917 , \40499 , \40186 );
not \U$40541 ( \40918 , \40917 );
or \U$40542 ( \40919 , \40916 , \40918 );
or \U$40543 ( \40920 , \40917 , \40197 );
nand \U$40544 ( \40921 , \40919 , \40920 );
not \U$40545 ( \40922 , \40921 );
not \U$40546 ( \40923 , \40523 );
not \U$40547 ( \40924 , \40880 );
not \U$40548 ( \40925 , \40859 );
and \U$40549 ( \40926 , \40924 , \40925 );
and \U$40550 ( \40927 , \40880 , \40859 );
nor \U$40551 ( \40928 , \40926 , \40927 );
not \U$40552 ( \40929 , \40928 );
or \U$40553 ( \40930 , \40923 , \40929 );
or \U$40554 ( \40931 , \40928 , \40523 );
nand \U$40555 ( \40932 , \40930 , \40931 );
not \U$40556 ( \40933 , \40932 );
or \U$40557 ( \40934 , \40922 , \40933 );
or \U$40558 ( \40935 , \40932 , \40921 );
xor \U$40559 ( \40936 , \40595 , \9273 );
xor \U$40560 ( \40937 , \40936 , \40603 );
xor \U$40561 ( \40938 , \40570 , \40577 );
xor \U$40562 ( \40939 , \40938 , \40585 );
and \U$40563 ( \40940 , \40937 , \40939 );
xor \U$40564 ( \40941 , \40614 , \40621 );
xor \U$40565 ( \40942 , \40941 , \40629 );
xor \U$40566 ( \40943 , \40570 , \40577 );
xor \U$40567 ( \40944 , \40943 , \40585 );
and \U$40568 ( \40945 , \40942 , \40944 );
and \U$40569 ( \40946 , \40937 , \40942 );
or \U$40570 ( \40947 , \40940 , \40945 , \40946 );
xor \U$40571 ( \40948 , \40663 , \40671 );
xor \U$40572 ( \40949 , \40681 , \40689 );
xor \U$40573 ( \40950 , \40949 , \40697 );
and \U$40574 ( \40951 , \40948 , \40950 );
xor \U$40575 ( \40952 , \40642 , \40649 );
xor \U$40576 ( \40953 , \40952 , \40658 );
xor \U$40577 ( \40954 , \40681 , \40689 );
xor \U$40578 ( \40955 , \40954 , \40697 );
and \U$40579 ( \40956 , \40953 , \40955 );
and \U$40580 ( \40957 , \40948 , \40953 );
or \U$40581 ( \40958 , \40951 , \40956 , \40957 );
xor \U$40582 ( \40959 , \40947 , \40958 );
xor \U$40583 ( \40960 , \40712 , \40719 );
xor \U$40584 ( \40961 , \40960 , \40727 );
xor \U$40585 ( \40962 , \40737 , \40744 );
xor \U$40586 ( \40963 , \40962 , \40752 );
xor \U$40587 ( \40964 , \40961 , \40963 );
xor \U$40588 ( \40965 , \40764 , \40771 );
xor \U$40589 ( \40966 , \40965 , \40779 );
and \U$40590 ( \40967 , \40964 , \40966 );
and \U$40591 ( \40968 , \40961 , \40963 );
or \U$40592 ( \40969 , \40967 , \40968 );
and \U$40593 ( \40970 , \40959 , \40969 );
and \U$40594 ( \40971 , \40947 , \40958 );
or \U$40595 ( \40972 , \40970 , \40971 );
and \U$40596 ( \40973 , \7633 , RIae76a00_54);
and \U$40597 ( \40974 , RIae76820_50, \7631 );
nor \U$40598 ( \40975 , \40973 , \40974 );
and \U$40599 ( \40976 , \40975 , \7206 );
not \U$40600 ( \40977 , \40975 );
and \U$40601 ( \40978 , \40977 , \7205 );
nor \U$40602 ( \40979 , \40976 , \40978 );
and \U$40603 ( \40980 , \6172 , RIae760a0_34);
and \U$40604 ( \40981 , RIae76370_40, \6170 );
nor \U$40605 ( \40982 , \40980 , \40981 );
and \U$40606 ( \40983 , \40982 , \6176 );
not \U$40607 ( \40984 , \40982 );
and \U$40608 ( \40985 , \40984 , \6175 );
nor \U$40609 ( \40986 , \40983 , \40985 );
xor \U$40610 ( \40987 , \40979 , \40986 );
and \U$40611 ( \40988 , \6941 , RIae76280_38);
and \U$40612 ( \40989 , RIae76af0_56, \6939 );
nor \U$40613 ( \40990 , \40988 , \40989 );
and \U$40614 ( \40991 , \40990 , \6314 );
not \U$40615 ( \40992 , \40990 );
and \U$40616 ( \40993 , \40992 , \6945 );
nor \U$40617 ( \40994 , \40991 , \40993 );
and \U$40618 ( \40995 , \40987 , \40994 );
and \U$40619 ( \40996 , \40979 , \40986 );
or \U$40620 ( \40997 , \40995 , \40996 );
and \U$40621 ( \40998 , \8371 , RIae76910_52);
and \U$40622 ( \40999 , RIae76be0_58, \8369 );
nor \U$40623 ( \41000 , \40998 , \40999 );
and \U$40624 ( \41001 , \41000 , \8020 );
not \U$40625 ( \41002 , \41000 );
and \U$40626 ( \41003 , \41002 , \8019 );
nor \U$40627 ( \41004 , \41001 , \41003 );
nand \U$40628 ( \41005 , RIae78e18_131, \9760 );
and \U$40629 ( \41006 , \41005 , \9273 );
not \U$40630 ( \41007 , \41005 );
and \U$40631 ( \41008 , \41007 , \9764 );
nor \U$40632 ( \41009 , \41006 , \41008 );
xor \U$40633 ( \41010 , \41004 , \41009 );
and \U$40634 ( \41011 , \8966 , RIae78ad0_124);
and \U$40635 ( \41012 , RIae78d28_129, \8964 );
nor \U$40636 ( \41013 , \41011 , \41012 );
and \U$40637 ( \41014 , \41013 , \8799 );
not \U$40638 ( \41015 , \41013 );
and \U$40639 ( \41016 , \41015 , \8789 );
nor \U$40640 ( \41017 , \41014 , \41016 );
and \U$40641 ( \41018 , \41010 , \41017 );
and \U$40642 ( \41019 , \41004 , \41009 );
or \U$40643 ( \41020 , \41018 , \41019 );
xor \U$40644 ( \41021 , \40997 , \41020 );
and \U$40645 ( \41022 , \5896 , RIae76640_46);
and \U$40646 ( \41023 , RIae76190_36, \5894 );
nor \U$40647 ( \41024 , \41022 , \41023 );
and \U$40648 ( \41025 , \41024 , \5590 );
not \U$40649 ( \41026 , \41024 );
and \U$40650 ( \41027 , \41026 , \5589 );
nor \U$40651 ( \41028 , \41025 , \41027 );
and \U$40652 ( \41029 , \4688 , RIae75470_8);
and \U$40653 ( \41030 , RIae76460_42, \4686 );
nor \U$40654 ( \41031 , \41029 , \41030 );
and \U$40655 ( \41032 , \41031 , \4481 );
not \U$40656 ( \41033 , \41031 );
and \U$40657 ( \41034 , \41033 , \4482 );
nor \U$40658 ( \41035 , \41032 , \41034 );
xor \U$40659 ( \41036 , \41028 , \41035 );
and \U$40660 ( \41037 , \5399 , RIae76550_44);
and \U$40661 ( \41038 , RIae76730_48, \5397 );
nor \U$40662 ( \41039 , \41037 , \41038 );
and \U$40663 ( \41040 , \41039 , \5016 );
not \U$40664 ( \41041 , \41039 );
and \U$40665 ( \41042 , \41041 , \5403 );
nor \U$40666 ( \41043 , \41040 , \41042 );
and \U$40667 ( \41044 , \41036 , \41043 );
and \U$40668 ( \41045 , \41028 , \41035 );
or \U$40669 ( \41046 , \41044 , \41045 );
and \U$40670 ( \41047 , \41021 , \41046 );
and \U$40671 ( \41048 , \40997 , \41020 );
or \U$40672 ( \41049 , \41047 , \41048 );
not \U$40673 ( \41050 , \469 );
and \U$40674 ( \41051 , \514 , RIae78080_102);
and \U$40675 ( \41052 , RIae78260_106, \512 );
nor \U$40676 ( \41053 , \41051 , \41052 );
not \U$40677 ( \41054 , \41053 );
or \U$40678 ( \41055 , \41050 , \41054 );
or \U$40679 ( \41056 , \41053 , \471 );
nand \U$40680 ( \41057 , \41055 , \41056 );
not \U$40681 ( \41058 , \400 );
and \U$40682 ( \41059 , \436 , RIae78170_104);
and \U$40683 ( \41060 , RIae77f90_100, \434 );
nor \U$40684 ( \41061 , \41059 , \41060 );
not \U$40685 ( \41062 , \41061 );
or \U$40686 ( \41063 , \41058 , \41062 );
or \U$40687 ( \41064 , \41061 , \402 );
nand \U$40688 ( \41065 , \41063 , \41064 );
xor \U$40689 ( \41066 , \41057 , \41065 );
and \U$40690 ( \41067 , \558 , RIae78620_114);
and \U$40691 ( \41068 , RIae78440_110, \556 );
nor \U$40692 ( \41069 , \41067 , \41068 );
and \U$40693 ( \41070 , \41069 , \504 );
not \U$40694 ( \41071 , \41069 );
and \U$40695 ( \41072 , \41071 , \562 );
nor \U$40696 ( \41073 , \41070 , \41072 );
and \U$40697 ( \41074 , \41066 , \41073 );
and \U$40698 ( \41075 , \41057 , \41065 );
or \U$40699 ( \41076 , \41074 , \41075 );
nand \U$40700 ( \41077 , RIae77270_72, RIae78b48_125);
and \U$40701 ( \41078 , \384 , RIae77360_74);
and \U$40702 ( \41079 , RIae78350_108, \382 );
nor \U$40703 ( \41080 , \41078 , \41079 );
not \U$40704 ( \41081 , \41080 );
not \U$40705 ( \41082 , \392 );
and \U$40706 ( \41083 , \41081 , \41082 );
and \U$40707 ( \41084 , \41080 , \392 );
nor \U$40708 ( \41085 , \41083 , \41084 );
nand \U$40709 ( \41086 , \41077 , \41085 );
xor \U$40710 ( \41087 , \41076 , \41086 );
and \U$40711 ( \41088 , \1138 , RIae77ea0_98);
and \U$40712 ( \41089 , RIae789e0_122, \1136 );
nor \U$40713 ( \41090 , \41088 , \41089 );
and \U$40714 ( \41091 , \41090 , \1012 );
not \U$40715 ( \41092 , \41090 );
and \U$40716 ( \41093 , \41092 , \1142 );
nor \U$40717 ( \41094 , \41091 , \41093 );
and \U$40718 ( \41095 , \672 , RIae784b8_111);
and \U$40719 ( \41096 , RIae77cc0_94, \670 );
nor \U$40720 ( \41097 , \41095 , \41096 );
and \U$40721 ( \41098 , \41097 , \588 );
not \U$40722 ( \41099 , \41097 );
and \U$40723 ( \41100 , \41099 , \587 );
nor \U$40724 ( \41101 , \41098 , \41100 );
xor \U$40725 ( \41102 , \41094 , \41101 );
not \U$40726 ( \41103 , \789 );
and \U$40727 ( \41104 , \883 , RIae77bd0_92);
and \U$40728 ( \41105 , RIae77db0_96, \881 );
nor \U$40729 ( \41106 , \41104 , \41105 );
not \U$40730 ( \41107 , \41106 );
or \U$40731 ( \41108 , \41103 , \41107 );
or \U$40732 ( \41109 , \41106 , \789 );
nand \U$40733 ( \41110 , \41108 , \41109 );
and \U$40734 ( \41111 , \41102 , \41110 );
and \U$40735 ( \41112 , \41094 , \41101 );
or \U$40736 ( \41113 , \41111 , \41112 );
and \U$40737 ( \41114 , \41087 , \41113 );
and \U$40738 ( \41115 , \41076 , \41086 );
or \U$40739 ( \41116 , \41114 , \41115 );
xor \U$40740 ( \41117 , \41049 , \41116 );
and \U$40741 ( \41118 , \4247 , RIae751a0_2);
and \U$40742 ( \41119 , RIae75380_6, \4245 );
nor \U$40743 ( \41120 , \41118 , \41119 );
and \U$40744 ( \41121 , \41120 , \3989 );
not \U$40745 ( \41122 , \41120 );
and \U$40746 ( \41123 , \41122 , \4251 );
nor \U$40747 ( \41124 , \41121 , \41123 );
not \U$40748 ( \41125 , \3218 );
and \U$40749 ( \41126 , \3214 , RIae75560_10);
and \U$40750 ( \41127 , RIae75830_16, \3212 );
nor \U$40751 ( \41128 , \41126 , \41127 );
not \U$40752 ( \41129 , \41128 );
or \U$40753 ( \41130 , \41125 , \41129 );
or \U$40754 ( \41131 , \41128 , \2774 );
nand \U$40755 ( \41132 , \41130 , \41131 );
xor \U$40756 ( \41133 , \41124 , \41132 );
and \U$40757 ( \41134 , \3730 , RIae75740_14);
and \U$40758 ( \41135 , RIae75290_4, \3728 );
nor \U$40759 ( \41136 , \41134 , \41135 );
and \U$40760 ( \41137 , \41136 , \3732 );
not \U$40761 ( \41138 , \41136 );
and \U$40762 ( \41139 , \41138 , \3421 );
nor \U$40763 ( \41140 , \41137 , \41139 );
and \U$40764 ( \41141 , \41133 , \41140 );
and \U$40765 ( \41142 , \41124 , \41132 );
or \U$40766 ( \41143 , \41141 , \41142 );
and \U$40767 ( \41144 , \2607 , RIae75ec0_30);
and \U$40768 ( \41145 , RIae75ce0_26, \2605 );
nor \U$40769 ( \41146 , \41144 , \41145 );
and \U$40770 ( \41147 , \41146 , \2611 );
not \U$40771 ( \41148 , \41146 );
and \U$40772 ( \41149 , \41148 , \2397 );
nor \U$40773 ( \41150 , \41147 , \41149 );
and \U$40774 ( \41151 , \2224 , RIae75920_18);
and \U$40775 ( \41152 , RIae75fb0_32, \2222 );
nor \U$40776 ( \41153 , \41151 , \41152 );
and \U$40777 ( \41154 , \41153 , \2061 );
not \U$40778 ( \41155 , \41153 );
and \U$40779 ( \41156 , \41155 , \2060 );
nor \U$40780 ( \41157 , \41154 , \41156 );
xor \U$40781 ( \41158 , \41150 , \41157 );
not \U$40782 ( \41159 , \3089 );
and \U$40783 ( \41160 , \2783 , RIae75dd0_28);
and \U$40784 ( \41161 , RIae75650_12, \2781 );
nor \U$40785 ( \41162 , \41160 , \41161 );
not \U$40786 ( \41163 , \41162 );
or \U$40787 ( \41164 , \41159 , \41163 );
or \U$40788 ( \41165 , \41162 , \2789 );
nand \U$40789 ( \41166 , \41164 , \41165 );
and \U$40790 ( \41167 , \41158 , \41166 );
and \U$40791 ( \41168 , \41150 , \41157 );
or \U$40792 ( \41169 , \41167 , \41168 );
xor \U$40793 ( \41170 , \41143 , \41169 );
and \U$40794 ( \41171 , \1939 , RIae75b00_22);
and \U$40795 ( \41172 , RIae75a10_20, \1937 );
nor \U$40796 ( \41173 , \41171 , \41172 );
and \U$40797 ( \41174 , \41173 , \1735 );
not \U$40798 ( \41175 , \41173 );
and \U$40799 ( \41176 , \41175 , \1734 );
nor \U$40800 ( \41177 , \41174 , \41176 );
and \U$40801 ( \41178 , \1376 , RIae788f0_120);
and \U$40802 ( \41179 , RIae78800_118, \1374 );
nor \U$40803 ( \41180 , \41178 , \41179 );
and \U$40804 ( \41181 , \41180 , \1380 );
not \U$40805 ( \41182 , \41180 );
and \U$40806 ( \41183 , \41182 , \1261 );
nor \U$40807 ( \41184 , \41181 , \41183 );
xor \U$40808 ( \41185 , \41177 , \41184 );
and \U$40809 ( \41186 , \1593 , RIae78710_116);
and \U$40810 ( \41187 , RIae75bf0_24, \1591 );
nor \U$40811 ( \41188 , \41186 , \41187 );
and \U$40812 ( \41189 , \41188 , \1498 );
not \U$40813 ( \41190 , \41188 );
and \U$40814 ( \41191 , \41190 , \1488 );
nor \U$40815 ( \41192 , \41189 , \41191 );
and \U$40816 ( \41193 , \41185 , \41192 );
and \U$40817 ( \41194 , \41177 , \41184 );
or \U$40818 ( \41195 , \41193 , \41194 );
and \U$40819 ( \41196 , \41170 , \41195 );
and \U$40820 ( \41197 , \41143 , \41169 );
or \U$40821 ( \41198 , \41196 , \41197 );
and \U$40822 ( \41199 , \41117 , \41198 );
and \U$40823 ( \41200 , \41049 , \41116 );
or \U$40824 ( \41201 , \41199 , \41200 );
xor \U$40825 ( \41202 , \40972 , \41201 );
xor \U$40826 ( \41203 , \40364 , \40371 );
xor \U$40827 ( \41204 , \41203 , \40379 );
xor \U$40828 ( \41205 , \40550 , \40555 );
xor \U$40829 ( \41206 , \41204 , \41205 );
xor \U$40830 ( \41207 , \40537 , \40446 );
xor \U$40831 ( \41208 , \41207 , \40544 );
and \U$40832 ( \41209 , \41206 , \41208 );
xor \U$40833 ( \41210 , \40259 , \40266 );
xor \U$40834 ( \41211 , \41210 , \40274 );
xor \U$40835 ( \41212 , \40525 , \40530 );
xor \U$40836 ( \41213 , \41211 , \41212 );
xor \U$40837 ( \41214 , \40537 , \40446 );
xor \U$40838 ( \41215 , \41214 , \40544 );
and \U$40839 ( \41216 , \41213 , \41215 );
and \U$40840 ( \41217 , \41206 , \41213 );
or \U$40841 ( \41218 , \41209 , \41216 , \41217 );
and \U$40842 ( \41219 , \41202 , \41218 );
and \U$40843 ( \41220 , \40972 , \41201 );
or \U$40844 ( \41221 , \41219 , \41220 );
xor \U$40845 ( \41222 , \40635 , \40703 );
xor \U$40846 ( \41223 , \41222 , \40785 );
xor \U$40847 ( \41224 , \40535 , \40547 );
xor \U$40848 ( \41225 , \41224 , \40560 );
and \U$40849 ( \41226 , \41223 , \41225 );
xor \U$40850 ( \41227 , \41221 , \41226 );
xor \U$40851 ( \41228 , \40730 , \40755 );
xor \U$40852 ( \41229 , \41228 , \40782 );
xor \U$40853 ( \41230 , \40661 , \40672 );
xor \U$40854 ( \41231 , \41230 , \40700 );
xor \U$40855 ( \41232 , \41229 , \41231 );
xor \U$40856 ( \41233 , \40588 , \40606 );
xor \U$40857 ( \41234 , \41233 , \40632 );
and \U$40858 ( \41235 , \41232 , \41234 );
and \U$40859 ( \41236 , \41229 , \41231 );
or \U$40860 ( \41237 , \41235 , \41236 );
xor \U$40861 ( \41238 , \40830 , \40832 );
xor \U$40862 ( \41239 , \41238 , \40843 );
and \U$40863 ( \41240 , \41237 , \41239 );
xor \U$40864 ( \41241 , \40791 , \40795 );
xor \U$40865 ( \41242 , \41241 , \40802 );
xor \U$40866 ( \41243 , \40830 , \40832 );
xor \U$40867 ( \41244 , \41243 , \40843 );
and \U$40868 ( \41245 , \41242 , \41244 );
and \U$40869 ( \41246 , \41237 , \41242 );
or \U$40870 ( \41247 , \41240 , \41245 , \41246 );
and \U$40871 ( \41248 , \41227 , \41247 );
and \U$40872 ( \41249 , \41221 , \41226 );
or \U$40873 ( \41250 , \41248 , \41249 );
xor \U$40874 ( \41251 , \40814 , \40820 );
xor \U$40875 ( \41252 , \40563 , \40788 );
xor \U$40876 ( \41253 , \41252 , \40805 );
and \U$40877 ( \41254 , \41251 , \41253 );
xor \U$40878 ( \41255 , \40828 , \40846 );
xor \U$40879 ( \41256 , \41255 , \40853 );
xor \U$40880 ( \41257 , \40563 , \40788 );
xor \U$40881 ( \41258 , \41257 , \40805 );
and \U$40882 ( \41259 , \41256 , \41258 );
and \U$40883 ( \41260 , \41251 , \41256 );
or \U$40884 ( \41261 , \41254 , \41259 , \41260 );
and \U$40885 ( \41262 , \41250 , \41261 );
not \U$40886 ( \41263 , \41250 );
not \U$40887 ( \41264 , \41261 );
and \U$40888 ( \41265 , \41263 , \41264 );
xor \U$40889 ( \41266 , \40252 , \40480 );
xor \U$40890 ( \41267 , \41266 , \40496 );
xor \U$40891 ( \41268 , \40868 , \40875 );
xor \U$40892 ( \41269 , \41267 , \41268 );
nor \U$40893 ( \41270 , \41265 , \41269 );
nor \U$40894 ( \41271 , \41262 , \41270 );
not \U$40895 ( \41272 , \41271 );
nand \U$40896 ( \41273 , \40935 , \41272 );
nand \U$40897 ( \41274 , \40934 , \41273 );
not \U$40898 ( \41275 , \41274 );
and \U$40899 ( \41276 , \40915 , \41275 );
and \U$40900 ( \41277 , \40914 , \41274 );
nor \U$40901 ( \41278 , \41276 , \41277 );
not \U$40902 ( \41279 , \41271 );
not \U$40903 ( \41280 , \40921 );
and \U$40904 ( \41281 , \41279 , \41280 );
and \U$40905 ( \41282 , \41271 , \40921 );
nor \U$40906 ( \41283 , \41281 , \41282 );
not \U$40907 ( \41284 , \41283 );
not \U$40908 ( \41285 , \40932 );
and \U$40909 ( \41286 , \41284 , \41285 );
and \U$40910 ( \41287 , \41283 , \40932 );
nor \U$40911 ( \41288 , \41286 , \41287 );
not \U$40912 ( \41289 , \41288 );
xor \U$40913 ( \41290 , \41028 , \41035 );
xor \U$40914 ( \41291 , \41290 , \41043 );
xor \U$40915 ( \41292 , \41004 , \41009 );
xor \U$40916 ( \41293 , \41292 , \41017 );
and \U$40917 ( \41294 , \41291 , \41293 );
xor \U$40918 ( \41295 , \40979 , \40986 );
xor \U$40919 ( \41296 , \41295 , \40994 );
xor \U$40920 ( \41297 , \41004 , \41009 );
xor \U$40921 ( \41298 , \41297 , \41017 );
and \U$40922 ( \41299 , \41296 , \41298 );
and \U$40923 ( \41300 , \41291 , \41296 );
or \U$40924 ( \41301 , \41294 , \41299 , \41300 );
or \U$40925 ( \41302 , \41085 , \41077 );
nand \U$40926 ( \41303 , \41302 , \41086 );
xor \U$40927 ( \41304 , \41057 , \41065 );
xor \U$40928 ( \41305 , \41304 , \41073 );
and \U$40929 ( \41306 , \41303 , \41305 );
xor \U$40930 ( \41307 , \41094 , \41101 );
xor \U$40931 ( \41308 , \41307 , \41110 );
xor \U$40932 ( \41309 , \41057 , \41065 );
xor \U$40933 ( \41310 , \41309 , \41073 );
and \U$40934 ( \41311 , \41308 , \41310 );
and \U$40935 ( \41312 , \41303 , \41308 );
or \U$40936 ( \41313 , \41306 , \41311 , \41312 );
xor \U$40937 ( \41314 , \41301 , \41313 );
xor \U$40938 ( \41315 , \41177 , \41184 );
xor \U$40939 ( \41316 , \41315 , \41192 );
xor \U$40940 ( \41317 , \41124 , \41132 );
xor \U$40941 ( \41318 , \41317 , \41140 );
and \U$40942 ( \41319 , \41316 , \41318 );
xor \U$40943 ( \41320 , \41150 , \41157 );
xor \U$40944 ( \41321 , \41320 , \41166 );
xor \U$40945 ( \41322 , \41124 , \41132 );
xor \U$40946 ( \41323 , \41322 , \41140 );
and \U$40947 ( \41324 , \41321 , \41323 );
and \U$40948 ( \41325 , \41316 , \41321 );
or \U$40949 ( \41326 , \41319 , \41324 , \41325 );
and \U$40950 ( \41327 , \41314 , \41326 );
and \U$40951 ( \41328 , \41301 , \41313 );
or \U$40952 ( \41329 , \41327 , \41328 );
and \U$40953 ( \41330 , \4688 , RIae75380_6);
and \U$40954 ( \41331 , RIae75470_8, \4686 );
nor \U$40955 ( \41332 , \41330 , \41331 );
and \U$40956 ( \41333 , \41332 , \4481 );
not \U$40957 ( \41334 , \41332 );
and \U$40958 ( \41335 , \41334 , \4482 );
nor \U$40959 ( \41336 , \41333 , \41335 );
and \U$40960 ( \41337 , \3730 , RIae75830_16);
and \U$40961 ( \41338 , RIae75740_14, \3728 );
nor \U$40962 ( \41339 , \41337 , \41338 );
and \U$40963 ( \41340 , \41339 , \3732 );
not \U$40964 ( \41341 , \41339 );
and \U$40965 ( \41342 , \41341 , \3422 );
nor \U$40966 ( \41343 , \41340 , \41342 );
xor \U$40967 ( \41344 , \41336 , \41343 );
and \U$40968 ( \41345 , \4247 , RIae75290_4);
and \U$40969 ( \41346 , RIae751a0_2, \4245 );
nor \U$40970 ( \41347 , \41345 , \41346 );
and \U$40971 ( \41348 , \41347 , \3989 );
not \U$40972 ( \41349 , \41347 );
and \U$40973 ( \41350 , \41349 , \4251 );
nor \U$40974 ( \41351 , \41348 , \41350 );
and \U$40975 ( \41352 , \41344 , \41351 );
and \U$40976 ( \41353 , \41336 , \41343 );
or \U$40977 ( \41354 , \41352 , \41353 );
and \U$40978 ( \41355 , \1593 , RIae78800_118);
and \U$40979 ( \41356 , RIae78710_116, \1591 );
nor \U$40980 ( \41357 , \41355 , \41356 );
and \U$40981 ( \41358 , \41357 , \1488 );
not \U$40982 ( \41359 , \41357 );
and \U$40983 ( \41360 , \41359 , \1498 );
nor \U$40984 ( \41361 , \41358 , \41360 );
and \U$40985 ( \41362 , \1939 , RIae75bf0_24);
and \U$40986 ( \41363 , RIae75b00_22, \1937 );
nor \U$40987 ( \41364 , \41362 , \41363 );
and \U$40988 ( \41365 , \41364 , \1734 );
not \U$40989 ( \41366 , \41364 );
and \U$40990 ( \41367 , \41366 , \1735 );
nor \U$40991 ( \41368 , \41365 , \41367 );
or \U$40992 ( \41369 , \41361 , \41368 );
not \U$40993 ( \41370 , \41368 );
not \U$40994 ( \41371 , \41361 );
or \U$40995 ( \41372 , \41370 , \41371 );
and \U$40996 ( \41373 , \2224 , RIae75a10_20);
and \U$40997 ( \41374 , RIae75920_18, \2222 );
nor \U$40998 ( \41375 , \41373 , \41374 );
and \U$40999 ( \41376 , \41375 , \2061 );
not \U$41000 ( \41377 , \41375 );
and \U$41001 ( \41378 , \41377 , \2060 );
nor \U$41002 ( \41379 , \41376 , \41378 );
nand \U$41003 ( \41380 , \41372 , \41379 );
nand \U$41004 ( \41381 , \41369 , \41380 );
xor \U$41005 ( \41382 , \41354 , \41381 );
and \U$41006 ( \41383 , \2783 , RIae75ce0_26);
and \U$41007 ( \41384 , RIae75dd0_28, \2781 );
nor \U$41008 ( \41385 , \41383 , \41384 );
not \U$41009 ( \41386 , \41385 );
not \U$41010 ( \41387 , \2789 );
and \U$41011 ( \41388 , \41386 , \41387 );
and \U$41012 ( \41389 , \41385 , \2789 );
nor \U$41013 ( \41390 , \41388 , \41389 );
and \U$41014 ( \41391 , \3214 , RIae75650_12);
and \U$41015 ( \41392 , RIae75560_10, \3212 );
nor \U$41016 ( \41393 , \41391 , \41392 );
not \U$41017 ( \41394 , \41393 );
not \U$41018 ( \41395 , \2774 );
and \U$41019 ( \41396 , \41394 , \41395 );
and \U$41020 ( \41397 , \41393 , \3218 );
nor \U$41021 ( \41398 , \41396 , \41397 );
xor \U$41022 ( \41399 , \41390 , \41398 );
and \U$41023 ( \41400 , \2607 , RIae75fb0_32);
and \U$41024 ( \41401 , RIae75ec0_30, \2605 );
nor \U$41025 ( \41402 , \41400 , \41401 );
and \U$41026 ( \41403 , \41402 , \2397 );
not \U$41027 ( \41404 , \41402 );
and \U$41028 ( \41405 , \41404 , \2611 );
nor \U$41029 ( \41406 , \41403 , \41405 );
and \U$41030 ( \41407 , \41399 , \41406 );
and \U$41031 ( \41408 , \41390 , \41398 );
nor \U$41032 ( \41409 , \41407 , \41408 );
and \U$41033 ( \41410 , \41382 , \41409 );
and \U$41034 ( \41411 , \41354 , \41381 );
or \U$41035 ( \41412 , \41410 , \41411 );
and \U$41036 ( \41413 , \436 , RIae78350_108);
and \U$41037 ( \41414 , RIae78170_104, \434 );
nor \U$41038 ( \41415 , \41413 , \41414 );
not \U$41039 ( \41416 , \41415 );
not \U$41040 ( \41417 , \400 );
and \U$41041 ( \41418 , \41416 , \41417 );
and \U$41042 ( \41419 , \41415 , \400 );
nor \U$41043 ( \41420 , \41418 , \41419 );
nand \U$41044 ( \41421 , RIae77090_68, RIae78b48_125);
xor \U$41045 ( \41422 , \41420 , \41421 );
and \U$41046 ( \41423 , \384 , RIae77270_72);
and \U$41047 ( \41424 , RIae77360_74, \382 );
nor \U$41048 ( \41425 , \41423 , \41424 );
not \U$41049 ( \41426 , \41425 );
not \U$41050 ( \41427 , \392 );
and \U$41051 ( \41428 , \41426 , \41427 );
and \U$41052 ( \41429 , \41425 , \392 );
nor \U$41053 ( \41430 , \41428 , \41429 );
and \U$41054 ( \41431 , \41422 , \41430 );
and \U$41055 ( \41432 , \41420 , \41421 );
or \U$41056 ( \41433 , \41431 , \41432 );
and \U$41057 ( \41434 , \883 , RIae77cc0_94);
and \U$41058 ( \41435 , RIae77bd0_92, \881 );
nor \U$41059 ( \41436 , \41434 , \41435 );
not \U$41060 ( \41437 , \41436 );
not \U$41061 ( \41438 , \787 );
and \U$41062 ( \41439 , \41437 , \41438 );
and \U$41063 ( \41440 , \41436 , \789 );
nor \U$41064 ( \41441 , \41439 , \41440 );
and \U$41065 ( \41442 , \1138 , RIae77db0_96);
and \U$41066 ( \41443 , RIae77ea0_98, \1136 );
nor \U$41067 ( \41444 , \41442 , \41443 );
and \U$41068 ( \41445 , \41444 , \1142 );
not \U$41069 ( \41446 , \41444 );
and \U$41070 ( \41447 , \41446 , \1012 );
nor \U$41071 ( \41448 , \41445 , \41447 );
xor \U$41072 ( \41449 , \41441 , \41448 );
and \U$41073 ( \41450 , \1376 , RIae789e0_122);
and \U$41074 ( \41451 , RIae788f0_120, \1374 );
nor \U$41075 ( \41452 , \41450 , \41451 );
and \U$41076 ( \41453 , \41452 , \1261 );
not \U$41077 ( \41454 , \41452 );
and \U$41078 ( \41455 , \41454 , \1380 );
nor \U$41079 ( \41456 , \41453 , \41455 );
and \U$41080 ( \41457 , \41449 , \41456 );
and \U$41081 ( \41458 , \41441 , \41448 );
or \U$41082 ( \41459 , \41457 , \41458 );
xor \U$41083 ( \41460 , \41433 , \41459 );
and \U$41084 ( \41461 , \672 , RIae78440_110);
and \U$41085 ( \41462 , RIae784b8_111, \670 );
nor \U$41086 ( \41463 , \41461 , \41462 );
and \U$41087 ( \41464 , \41463 , \587 );
not \U$41088 ( \41465 , \41463 );
and \U$41089 ( \41466 , \41465 , \588 );
nor \U$41090 ( \41467 , \41464 , \41466 );
and \U$41091 ( \41468 , \514 , RIae77f90_100);
and \U$41092 ( \41469 , RIae78080_102, \512 );
nor \U$41093 ( \41470 , \41468 , \41469 );
not \U$41094 ( \41471 , \41470 );
not \U$41095 ( \41472 , \469 );
and \U$41096 ( \41473 , \41471 , \41472 );
and \U$41097 ( \41474 , \41470 , \471 );
nor \U$41098 ( \41475 , \41473 , \41474 );
xor \U$41099 ( \41476 , \41467 , \41475 );
and \U$41100 ( \41477 , \558 , RIae78260_106);
and \U$41101 ( \41478 , RIae78620_114, \556 );
nor \U$41102 ( \41479 , \41477 , \41478 );
and \U$41103 ( \41480 , \41479 , \562 );
not \U$41104 ( \41481 , \41479 );
and \U$41105 ( \41482 , \41481 , \504 );
nor \U$41106 ( \41483 , \41480 , \41482 );
and \U$41107 ( \41484 , \41476 , \41483 );
and \U$41108 ( \41485 , \41467 , \41475 );
or \U$41109 ( \41486 , \41484 , \41485 );
and \U$41110 ( \41487 , \41460 , \41486 );
and \U$41111 ( \41488 , \41433 , \41459 );
nor \U$41112 ( \41489 , \41487 , \41488 );
xor \U$41113 ( \41490 , \41412 , \41489 );
and \U$41114 ( \41491 , \6172 , RIae76190_36);
and \U$41115 ( \41492 , RIae760a0_34, \6170 );
nor \U$41116 ( \41493 , \41491 , \41492 );
and \U$41117 ( \41494 , \41493 , \6175 );
not \U$41118 ( \41495 , \41493 );
and \U$41119 ( \41496 , \41495 , \6176 );
nor \U$41120 ( \41497 , \41494 , \41496 );
and \U$41121 ( \41498 , \5399 , RIae76460_42);
and \U$41122 ( \41499 , RIae76550_44, \5397 );
nor \U$41123 ( \41500 , \41498 , \41499 );
and \U$41124 ( \41501 , \41500 , \5403 );
not \U$41125 ( \41502 , \41500 );
and \U$41126 ( \41503 , \41502 , \5016 );
nor \U$41127 ( \41504 , \41501 , \41503 );
xor \U$41128 ( \41505 , \41497 , \41504 );
and \U$41129 ( \41506 , \5896 , RIae76730_48);
and \U$41130 ( \41507 , RIae76640_46, \5894 );
nor \U$41131 ( \41508 , \41506 , \41507 );
and \U$41132 ( \41509 , \41508 , \5589 );
not \U$41133 ( \41510 , \41508 );
and \U$41134 ( \41511 , \41510 , \5590 );
nor \U$41135 ( \41512 , \41509 , \41511 );
and \U$41136 ( \41513 , \41505 , \41512 );
and \U$41137 ( \41514 , \41497 , \41504 );
or \U$41138 ( \41515 , \41513 , \41514 );
and \U$41139 ( \41516 , \7633 , RIae76af0_56);
and \U$41140 ( \41517 , RIae76a00_54, \7631 );
nor \U$41141 ( \41518 , \41516 , \41517 );
and \U$41142 ( \41519 , \41518 , \7205 );
not \U$41143 ( \41520 , \41518 );
and \U$41144 ( \41521 , \41520 , \7206 );
nor \U$41145 ( \41522 , \41519 , \41521 );
and \U$41146 ( \41523 , \6941 , RIae76370_40);
and \U$41147 ( \41524 , RIae76280_38, \6939 );
nor \U$41148 ( \41525 , \41523 , \41524 );
and \U$41149 ( \41526 , \41525 , \6945 );
not \U$41150 ( \41527 , \41525 );
and \U$41151 ( \41528 , \41527 , \6314 );
nor \U$41152 ( \41529 , \41526 , \41528 );
xor \U$41153 ( \41530 , \41522 , \41529 );
and \U$41154 ( \41531 , \8371 , RIae76820_50);
and \U$41155 ( \41532 , RIae76910_52, \8369 );
nor \U$41156 ( \41533 , \41531 , \41532 );
and \U$41157 ( \41534 , \41533 , \8019 );
not \U$41158 ( \41535 , \41533 );
and \U$41159 ( \41536 , \41535 , \8020 );
nor \U$41160 ( \41537 , \41534 , \41536 );
and \U$41161 ( \41538 , \41530 , \41537 );
and \U$41162 ( \41539 , \41522 , \41529 );
or \U$41163 ( \41540 , \41538 , \41539 );
xor \U$41164 ( \41541 , \41515 , \41540 );
and \U$41165 ( \41542 , \9760 , RIae78d28_129);
and \U$41166 ( \41543 , RIae78e18_131, \9758 );
nor \U$41167 ( \41544 , \41542 , \41543 );
and \U$41168 ( \41545 , \41544 , \9764 );
not \U$41169 ( \41546 , \41544 );
and \U$41170 ( \41547 , \41546 , \9273 );
nor \U$41171 ( \41548 , \41545 , \41547 );
xor \U$41172 ( \41549 , \41548 , \10118 );
and \U$41173 ( \41550 , \8966 , RIae76be0_58);
and \U$41174 ( \41551 , RIae78ad0_124, \8964 );
nor \U$41175 ( \41552 , \41550 , \41551 );
and \U$41176 ( \41553 , \41552 , \8789 );
not \U$41177 ( \41554 , \41552 );
and \U$41178 ( \41555 , \41554 , \8799 );
nor \U$41179 ( \41556 , \41553 , \41555 );
and \U$41180 ( \41557 , \41549 , \41556 );
and \U$41181 ( \41558 , \41548 , \10118 );
or \U$41182 ( \41559 , \41557 , \41558 );
and \U$41183 ( \41560 , \41541 , \41559 );
and \U$41184 ( \41561 , \41515 , \41540 );
nor \U$41185 ( \41562 , \41560 , \41561 );
and \U$41186 ( \41563 , \41490 , \41562 );
and \U$41187 ( \41564 , \41412 , \41489 );
or \U$41188 ( \41565 , \41563 , \41564 );
xor \U$41189 ( \41566 , \41329 , \41565 );
xor \U$41190 ( \41567 , \40570 , \40577 );
xor \U$41191 ( \41568 , \41567 , \40585 );
xor \U$41192 ( \41569 , \40937 , \40942 );
xor \U$41193 ( \41570 , \41568 , \41569 );
xor \U$41194 ( \41571 , \40961 , \40963 );
xor \U$41195 ( \41572 , \41571 , \40966 );
and \U$41196 ( \41573 , \41570 , \41572 );
xor \U$41197 ( \41574 , \40681 , \40689 );
xor \U$41198 ( \41575 , \41574 , \40697 );
xor \U$41199 ( \41576 , \40948 , \40953 );
xor \U$41200 ( \41577 , \41575 , \41576 );
xor \U$41201 ( \41578 , \40961 , \40963 );
xor \U$41202 ( \41579 , \41578 , \40966 );
and \U$41203 ( \41580 , \41577 , \41579 );
and \U$41204 ( \41581 , \41570 , \41577 );
or \U$41205 ( \41582 , \41573 , \41580 , \41581 );
and \U$41206 ( \41583 , \41566 , \41582 );
and \U$41207 ( \41584 , \41329 , \41565 );
or \U$41208 ( \41585 , \41583 , \41584 );
xor \U$41209 ( \41586 , \41049 , \41116 );
xor \U$41210 ( \41587 , \41586 , \41198 );
xor \U$41211 ( \41588 , \40947 , \40958 );
xor \U$41212 ( \41589 , \41588 , \40969 );
and \U$41213 ( \41590 , \41587 , \41589 );
xor \U$41214 ( \41591 , \41585 , \41590 );
xor \U$41215 ( \41592 , \41143 , \41169 );
xor \U$41216 ( \41593 , \41592 , \41195 );
xor \U$41217 ( \41594 , \41076 , \41086 );
xor \U$41218 ( \41595 , \41594 , \41113 );
xor \U$41219 ( \41596 , \41593 , \41595 );
xor \U$41220 ( \41597 , \40997 , \41020 );
xor \U$41221 ( \41598 , \41597 , \41046 );
and \U$41222 ( \41599 , \41596 , \41598 );
and \U$41223 ( \41600 , \41593 , \41595 );
or \U$41224 ( \41601 , \41599 , \41600 );
xor \U$41225 ( \41602 , \41229 , \41231 );
xor \U$41226 ( \41603 , \41602 , \41234 );
and \U$41227 ( \41604 , \41601 , \41603 );
xor \U$41228 ( \41605 , \40537 , \40446 );
xor \U$41229 ( \41606 , \41605 , \40544 );
xor \U$41230 ( \41607 , \41206 , \41213 );
xor \U$41231 ( \41608 , \41606 , \41607 );
xor \U$41232 ( \41609 , \41229 , \41231 );
xor \U$41233 ( \41610 , \41609 , \41234 );
and \U$41234 ( \41611 , \41608 , \41610 );
and \U$41235 ( \41612 , \41601 , \41608 );
or \U$41236 ( \41613 , \41604 , \41611 , \41612 );
and \U$41237 ( \41614 , \41591 , \41613 );
and \U$41238 ( \41615 , \41585 , \41590 );
or \U$41239 ( \41616 , \41614 , \41615 );
xor \U$41240 ( \41617 , \41223 , \41225 );
xor \U$41241 ( \41618 , \40972 , \41201 );
xor \U$41242 ( \41619 , \41618 , \41218 );
and \U$41243 ( \41620 , \41617 , \41619 );
xor \U$41244 ( \41621 , \40830 , \40832 );
xor \U$41245 ( \41622 , \41621 , \40843 );
xor \U$41246 ( \41623 , \41237 , \41242 );
xor \U$41247 ( \41624 , \41622 , \41623 );
xor \U$41248 ( \41625 , \40972 , \41201 );
xor \U$41249 ( \41626 , \41625 , \41218 );
and \U$41250 ( \41627 , \41624 , \41626 );
and \U$41251 ( \41628 , \41617 , \41624 );
or \U$41252 ( \41629 , \41620 , \41627 , \41628 );
xor \U$41253 ( \41630 , \41616 , \41629 );
xor \U$41254 ( \41631 , \40563 , \40788 );
xor \U$41255 ( \41632 , \41631 , \40805 );
xor \U$41256 ( \41633 , \41251 , \41256 );
xor \U$41257 ( \41634 , \41632 , \41633 );
and \U$41258 ( \41635 , \41630 , \41634 );
and \U$41259 ( \41636 , \41616 , \41629 );
or \U$41260 ( \41637 , \41635 , \41636 );
xor \U$41261 ( \41638 , \40808 , \40821 );
xor \U$41262 ( \41639 , \41638 , \40856 );
xor \U$41263 ( \41640 , \41637 , \41639 );
not \U$41264 ( \41641 , \41269 );
xor \U$41265 ( \41642 , \41261 , \41250 );
not \U$41266 ( \41643 , \41642 );
or \U$41267 ( \41644 , \41641 , \41643 );
or \U$41268 ( \41645 , \41642 , \41269 );
nand \U$41269 ( \41646 , \41644 , \41645 );
and \U$41270 ( \41647 , \41640 , \41646 );
and \U$41271 ( \41648 , \41637 , \41639 );
or \U$41272 ( \41649 , \41647 , \41648 );
nand \U$41273 ( \41650 , \41289 , \41649 );
or \U$41274 ( \41651 , \41278 , \41650 );
xnor \U$41275 ( \41652 , \41650 , \41278 );
xor \U$41276 ( \41653 , \41412 , \41489 );
xor \U$41277 ( \41654 , \41653 , \41562 );
xor \U$41278 ( \41655 , \41301 , \41313 );
xor \U$41279 ( \41656 , \41655 , \41326 );
xor \U$41280 ( \41657 , \41654 , \41656 );
not \U$41281 ( \41658 , \41657 );
xor \U$41282 ( \41659 , \41548 , \10118 );
xor \U$41283 ( \41660 , \41659 , \41556 );
xor \U$41284 ( \41661 , \41497 , \41504 );
xor \U$41285 ( \41662 , \41661 , \41512 );
and \U$41286 ( \41663 , \41660 , \41662 );
xor \U$41287 ( \41664 , \41522 , \41529 );
xor \U$41288 ( \41665 , \41664 , \41537 );
xor \U$41289 ( \41666 , \41497 , \41504 );
xor \U$41290 ( \41667 , \41666 , \41512 );
and \U$41291 ( \41668 , \41665 , \41667 );
and \U$41292 ( \41669 , \41660 , \41665 );
or \U$41293 ( \41670 , \41663 , \41668 , \41669 );
xor \U$41294 ( \41671 , \41467 , \41475 );
xor \U$41295 ( \41672 , \41671 , \41483 );
xor \U$41296 ( \41673 , \41441 , \41448 );
xor \U$41297 ( \41674 , \41673 , \41456 );
and \U$41298 ( \41675 , \41672 , \41674 );
xor \U$41299 ( \41676 , \41420 , \41421 );
xor \U$41300 ( \41677 , \41676 , \41430 );
xor \U$41301 ( \41678 , \41441 , \41448 );
xor \U$41302 ( \41679 , \41678 , \41456 );
and \U$41303 ( \41680 , \41677 , \41679 );
and \U$41304 ( \41681 , \41672 , \41677 );
or \U$41305 ( \41682 , \41675 , \41680 , \41681 );
or \U$41306 ( \41683 , \41670 , \41682 );
not \U$41307 ( \41684 , \41682 );
not \U$41308 ( \41685 , \41670 );
or \U$41309 ( \41686 , \41684 , \41685 );
not \U$41310 ( \41687 , \41368 );
not \U$41311 ( \41688 , \41379 );
or \U$41312 ( \41689 , \41687 , \41688 );
or \U$41313 ( \41690 , \41368 , \41379 );
nand \U$41314 ( \41691 , \41689 , \41690 );
not \U$41315 ( \41692 , \41691 );
not \U$41316 ( \41693 , \41361 );
and \U$41317 ( \41694 , \41692 , \41693 );
and \U$41318 ( \41695 , \41691 , \41361 );
nor \U$41319 ( \41696 , \41694 , \41695 );
xor \U$41320 ( \41697 , \41390 , \41398 );
xor \U$41321 ( \41698 , \41697 , \41406 );
or \U$41322 ( \41699 , \41696 , \41698 );
not \U$41323 ( \41700 , \41698 );
not \U$41324 ( \41701 , \41696 );
or \U$41325 ( \41702 , \41700 , \41701 );
xor \U$41326 ( \41703 , \41336 , \41343 );
xor \U$41327 ( \41704 , \41703 , \41351 );
nand \U$41328 ( \41705 , \41702 , \41704 );
nand \U$41329 ( \41706 , \41699 , \41705 );
nand \U$41330 ( \41707 , \41686 , \41706 );
nand \U$41331 ( \41708 , \41683 , \41707 );
and \U$41332 ( \41709 , \8966 , RIae76910_52);
and \U$41333 ( \41710 , RIae76be0_58, \8964 );
nor \U$41334 ( \41711 , \41709 , \41710 );
and \U$41335 ( \41712 , \41711 , \8789 );
not \U$41336 ( \41713 , \41711 );
and \U$41337 ( \41714 , \41713 , \8799 );
nor \U$41338 ( \41715 , \41712 , \41714 );
not \U$41339 ( \41716 , \41715 );
and \U$41340 ( \41717 , \9760 , RIae78ad0_124);
and \U$41341 ( \41718 , RIae78d28_129, \9758 );
nor \U$41342 ( \41719 , \41717 , \41718 );
and \U$41343 ( \41720 , \41719 , \9272 );
not \U$41344 ( \41721 , \41719 );
and \U$41345 ( \41722 , \41721 , \9273 );
nor \U$41346 ( \41723 , \41720 , \41722 );
not \U$41347 ( \41724 , \41723 );
and \U$41348 ( \41725 , \41716 , \41724 );
and \U$41349 ( \41726 , \41723 , \41715 );
nand \U$41350 ( \41727 , RIae78e18_131, \10548 );
and \U$41351 ( \41728 , \41727 , \10118 );
not \U$41352 ( \41729 , \41727 );
and \U$41353 ( \41730 , \41729 , \10421 );
nor \U$41354 ( \41731 , \41728 , \41730 );
nor \U$41355 ( \41732 , \41726 , \41731 );
nor \U$41356 ( \41733 , \41725 , \41732 );
and \U$41357 ( \41734 , \5399 , RIae75470_8);
and \U$41358 ( \41735 , RIae76460_42, \5397 );
nor \U$41359 ( \41736 , \41734 , \41735 );
and \U$41360 ( \41737 , \41736 , \5403 );
not \U$41361 ( \41738 , \41736 );
and \U$41362 ( \41739 , \41738 , \5016 );
nor \U$41363 ( \41740 , \41737 , \41739 );
not \U$41364 ( \41741 , \41740 );
and \U$41365 ( \41742 , \5896 , RIae76550_44);
and \U$41366 ( \41743 , RIae76730_48, \5894 );
nor \U$41367 ( \41744 , \41742 , \41743 );
and \U$41368 ( \41745 , \41744 , \5589 );
not \U$41369 ( \41746 , \41744 );
and \U$41370 ( \41747 , \41746 , \5590 );
nor \U$41371 ( \41748 , \41745 , \41747 );
not \U$41372 ( \41749 , \41748 );
and \U$41373 ( \41750 , \41741 , \41749 );
and \U$41374 ( \41751 , \41748 , \41740 );
and \U$41375 ( \41752 , \6172 , RIae76640_46);
and \U$41376 ( \41753 , RIae76190_36, \6170 );
nor \U$41377 ( \41754 , \41752 , \41753 );
and \U$41378 ( \41755 , \41754 , \6175 );
not \U$41379 ( \41756 , \41754 );
and \U$41380 ( \41757 , \41756 , \6176 );
nor \U$41381 ( \41758 , \41755 , \41757 );
nor \U$41382 ( \41759 , \41751 , \41758 );
nor \U$41383 ( \41760 , \41750 , \41759 );
or \U$41384 ( \41761 , \41733 , \41760 );
not \U$41385 ( \41762 , \41733 );
not \U$41386 ( \41763 , \41760 );
or \U$41387 ( \41764 , \41762 , \41763 );
and \U$41388 ( \41765 , \8371 , RIae76a00_54);
and \U$41389 ( \41766 , RIae76820_50, \8369 );
nor \U$41390 ( \41767 , \41765 , \41766 );
and \U$41391 ( \41768 , \41767 , \8020 );
not \U$41392 ( \41769 , \41767 );
and \U$41393 ( \41770 , \41769 , \8019 );
nor \U$41394 ( \41771 , \41768 , \41770 );
and \U$41395 ( \41772 , \6941 , RIae760a0_34);
and \U$41396 ( \41773 , RIae76370_40, \6939 );
nor \U$41397 ( \41774 , \41772 , \41773 );
and \U$41398 ( \41775 , \41774 , \6314 );
not \U$41399 ( \41776 , \41774 );
and \U$41400 ( \41777 , \41776 , \6945 );
nor \U$41401 ( \41778 , \41775 , \41777 );
xor \U$41402 ( \41779 , \41771 , \41778 );
and \U$41403 ( \41780 , \7633 , RIae76280_38);
and \U$41404 ( \41781 , RIae76af0_56, \7631 );
nor \U$41405 ( \41782 , \41780 , \41781 );
and \U$41406 ( \41783 , \41782 , \7206 );
not \U$41407 ( \41784 , \41782 );
and \U$41408 ( \41785 , \41784 , \7205 );
nor \U$41409 ( \41786 , \41783 , \41785 );
and \U$41410 ( \41787 , \41779 , \41786 );
and \U$41411 ( \41788 , \41771 , \41778 );
or \U$41412 ( \41789 , \41787 , \41788 );
nand \U$41413 ( \41790 , \41764 , \41789 );
nand \U$41414 ( \41791 , \41761 , \41790 );
and \U$41415 ( \41792 , \436 , RIae77360_74);
and \U$41416 ( \41793 , RIae78350_108, \434 );
nor \U$41417 ( \41794 , \41792 , \41793 );
not \U$41418 ( \41795 , \41794 );
not \U$41419 ( \41796 , \400 );
and \U$41420 ( \41797 , \41795 , \41796 );
and \U$41421 ( \41798 , \41794 , \402 );
nor \U$41422 ( \41799 , \41797 , \41798 );
nand \U$41423 ( \41800 , RIae77108_69, RIae78b48_125);
xor \U$41424 ( \41801 , \41799 , \41800 );
and \U$41425 ( \41802 , \384 , RIae77090_68);
and \U$41426 ( \41803 , RIae77270_72, \382 );
nor \U$41427 ( \41804 , \41802 , \41803 );
not \U$41428 ( \41805 , \41804 );
not \U$41429 ( \41806 , \392 );
and \U$41430 ( \41807 , \41805 , \41806 );
and \U$41431 ( \41808 , \41804 , \388 );
nor \U$41432 ( \41809 , \41807 , \41808 );
and \U$41433 ( \41810 , \41801 , \41809 );
and \U$41434 ( \41811 , \41799 , \41800 );
or \U$41435 ( \41812 , \41810 , \41811 );
and \U$41436 ( \41813 , \1138 , RIae77bd0_92);
and \U$41437 ( \41814 , RIae77db0_96, \1136 );
nor \U$41438 ( \41815 , \41813 , \41814 );
and \U$41439 ( \41816 , \41815 , \1012 );
not \U$41440 ( \41817 , \41815 );
and \U$41441 ( \41818 , \41817 , \1142 );
nor \U$41442 ( \41819 , \41816 , \41818 );
and \U$41443 ( \41820 , \1376 , RIae77ea0_98);
and \U$41444 ( \41821 , RIae789e0_122, \1374 );
nor \U$41445 ( \41822 , \41820 , \41821 );
and \U$41446 ( \41823 , \41822 , \1380 );
not \U$41447 ( \41824 , \41822 );
and \U$41448 ( \41825 , \41824 , \1261 );
nor \U$41449 ( \41826 , \41823 , \41825 );
xor \U$41450 ( \41827 , \41819 , \41826 );
not \U$41451 ( \41828 , \789 );
and \U$41452 ( \41829 , \883 , RIae784b8_111);
and \U$41453 ( \41830 , RIae77cc0_94, \881 );
nor \U$41454 ( \41831 , \41829 , \41830 );
not \U$41455 ( \41832 , \41831 );
or \U$41456 ( \41833 , \41828 , \41832 );
or \U$41457 ( \41834 , \41831 , \787 );
nand \U$41458 ( \41835 , \41833 , \41834 );
and \U$41459 ( \41836 , \41827 , \41835 );
and \U$41460 ( \41837 , \41819 , \41826 );
nor \U$41461 ( \41838 , \41836 , \41837 );
xor \U$41462 ( \41839 , \41812 , \41838 );
and \U$41463 ( \41840 , \514 , RIae78170_104);
and \U$41464 ( \41841 , RIae77f90_100, \512 );
nor \U$41465 ( \41842 , \41840 , \41841 );
not \U$41466 ( \41843 , \41842 );
not \U$41467 ( \41844 , \471 );
and \U$41468 ( \41845 , \41843 , \41844 );
and \U$41469 ( \41846 , \41842 , \471 );
nor \U$41470 ( \41847 , \41845 , \41846 );
and \U$41471 ( \41848 , \558 , RIae78080_102);
and \U$41472 ( \41849 , RIae78260_106, \556 );
nor \U$41473 ( \41850 , \41848 , \41849 );
and \U$41474 ( \41851 , \41850 , \562 );
not \U$41475 ( \41852 , \41850 );
and \U$41476 ( \41853 , \41852 , \504 );
nor \U$41477 ( \41854 , \41851 , \41853 );
xor \U$41478 ( \41855 , \41847 , \41854 );
and \U$41479 ( \41856 , \672 , RIae78620_114);
and \U$41480 ( \41857 , RIae78440_110, \670 );
nor \U$41481 ( \41858 , \41856 , \41857 );
and \U$41482 ( \41859 , \41858 , \587 );
not \U$41483 ( \41860 , \41858 );
and \U$41484 ( \41861 , \41860 , \588 );
nor \U$41485 ( \41862 , \41859 , \41861 );
and \U$41486 ( \41863 , \41855 , \41862 );
and \U$41487 ( \41864 , \41847 , \41854 );
or \U$41488 ( \41865 , \41863 , \41864 );
and \U$41489 ( \41866 , \41839 , \41865 );
and \U$41490 ( \41867 , \41812 , \41838 );
nor \U$41491 ( \41868 , \41866 , \41867 );
xor \U$41492 ( \41869 , \41791 , \41868 );
not \U$41493 ( \41870 , \2789 );
and \U$41494 ( \41871 , \2783 , RIae75ec0_30);
and \U$41495 ( \41872 , RIae75ce0_26, \2781 );
nor \U$41496 ( \41873 , \41871 , \41872 );
not \U$41497 ( \41874 , \41873 );
or \U$41498 ( \41875 , \41870 , \41874 );
or \U$41499 ( \41876 , \41873 , \2789 );
nand \U$41500 ( \41877 , \41875 , \41876 );
not \U$41501 ( \41878 , \3218 );
and \U$41502 ( \41879 , \3214 , RIae75dd0_28);
and \U$41503 ( \41880 , RIae75650_12, \3212 );
nor \U$41504 ( \41881 , \41879 , \41880 );
not \U$41505 ( \41882 , \41881 );
or \U$41506 ( \41883 , \41878 , \41882 );
or \U$41507 ( \41884 , \41881 , \3218 );
nand \U$41508 ( \41885 , \41883 , \41884 );
xor \U$41509 ( \41886 , \41877 , \41885 );
and \U$41510 ( \41887 , \2607 , RIae75920_18);
and \U$41511 ( \41888 , RIae75fb0_32, \2605 );
nor \U$41512 ( \41889 , \41887 , \41888 );
and \U$41513 ( \41890 , \41889 , \2611 );
not \U$41514 ( \41891 , \41889 );
and \U$41515 ( \41892 , \41891 , \2397 );
nor \U$41516 ( \41893 , \41890 , \41892 );
and \U$41517 ( \41894 , \41886 , \41893 );
and \U$41518 ( \41895 , \41877 , \41885 );
nor \U$41519 ( \41896 , \41894 , \41895 );
and \U$41520 ( \41897 , \4247 , RIae75740_14);
and \U$41521 ( \41898 , RIae75290_4, \4245 );
nor \U$41522 ( \41899 , \41897 , \41898 );
and \U$41523 ( \41900 , \41899 , \3989 );
not \U$41524 ( \41901 , \41899 );
and \U$41525 ( \41902 , \41901 , \4251 );
nor \U$41526 ( \41903 , \41900 , \41902 );
and \U$41527 ( \41904 , \4688 , RIae751a0_2);
and \U$41528 ( \41905 , RIae75380_6, \4686 );
nor \U$41529 ( \41906 , \41904 , \41905 );
and \U$41530 ( \41907 , \41906 , \4481 );
not \U$41531 ( \41908 , \41906 );
and \U$41532 ( \41909 , \41908 , \4482 );
nor \U$41533 ( \41910 , \41907 , \41909 );
xor \U$41534 ( \41911 , \41903 , \41910 );
and \U$41535 ( \41912 , \3730 , RIae75560_10);
and \U$41536 ( \41913 , RIae75830_16, \3728 );
nor \U$41537 ( \41914 , \41912 , \41913 );
and \U$41538 ( \41915 , \41914 , \3732 );
not \U$41539 ( \41916 , \41914 );
and \U$41540 ( \41917 , \41916 , \3422 );
nor \U$41541 ( \41918 , \41915 , \41917 );
and \U$41542 ( \41919 , \41911 , \41918 );
and \U$41543 ( \41920 , \41903 , \41910 );
nor \U$41544 ( \41921 , \41919 , \41920 );
xor \U$41545 ( \41922 , \41896 , \41921 );
and \U$41546 ( \41923 , \1939 , RIae78710_116);
and \U$41547 ( \41924 , RIae75bf0_24, \1937 );
nor \U$41548 ( \41925 , \41923 , \41924 );
and \U$41549 ( \41926 , \41925 , \1735 );
not \U$41550 ( \41927 , \41925 );
and \U$41551 ( \41928 , \41927 , \1734 );
nor \U$41552 ( \41929 , \41926 , \41928 );
and \U$41553 ( \41930 , \2224 , RIae75b00_22);
and \U$41554 ( \41931 , RIae75a10_20, \2222 );
nor \U$41555 ( \41932 , \41930 , \41931 );
and \U$41556 ( \41933 , \41932 , \2061 );
not \U$41557 ( \41934 , \41932 );
and \U$41558 ( \41935 , \41934 , \2060 );
nor \U$41559 ( \41936 , \41933 , \41935 );
xor \U$41560 ( \41937 , \41929 , \41936 );
and \U$41561 ( \41938 , \1593 , RIae788f0_120);
and \U$41562 ( \41939 , RIae78800_118, \1591 );
nor \U$41563 ( \41940 , \41938 , \41939 );
and \U$41564 ( \41941 , \41940 , \1498 );
not \U$41565 ( \41942 , \41940 );
and \U$41566 ( \41943 , \41942 , \1488 );
nor \U$41567 ( \41944 , \41941 , \41943 );
and \U$41568 ( \41945 , \41937 , \41944 );
and \U$41569 ( \41946 , \41929 , \41936 );
nor \U$41570 ( \41947 , \41945 , \41946 );
and \U$41571 ( \41948 , \41922 , \41947 );
and \U$41572 ( \41949 , \41896 , \41921 );
nor \U$41573 ( \41950 , \41948 , \41949 );
and \U$41574 ( \41951 , \41869 , \41950 );
and \U$41575 ( \41952 , \41791 , \41868 );
or \U$41576 ( \41953 , \41951 , \41952 );
xor \U$41577 ( \41954 , \41708 , \41953 );
xor \U$41578 ( \41955 , \41004 , \41009 );
xor \U$41579 ( \41956 , \41955 , \41017 );
xor \U$41580 ( \41957 , \41291 , \41296 );
xor \U$41581 ( \41958 , \41956 , \41957 );
not \U$41582 ( \41959 , \41958 );
xor \U$41583 ( \41960 , \41057 , \41065 );
xor \U$41584 ( \41961 , \41960 , \41073 );
xor \U$41585 ( \41962 , \41303 , \41308 );
xor \U$41586 ( \41963 , \41961 , \41962 );
not \U$41587 ( \41964 , \41963 );
or \U$41588 ( \41965 , \41959 , \41964 );
or \U$41589 ( \41966 , \41963 , \41958 );
xor \U$41590 ( \41967 , \41124 , \41132 );
xor \U$41591 ( \41968 , \41967 , \41140 );
xor \U$41592 ( \41969 , \41316 , \41321 );
xor \U$41593 ( \41970 , \41968 , \41969 );
nand \U$41594 ( \41971 , \41966 , \41970 );
nand \U$41595 ( \41972 , \41965 , \41971 );
xor \U$41596 ( \41973 , \41954 , \41972 );
not \U$41597 ( \41974 , \41973 );
or \U$41598 ( \41975 , \41658 , \41974 );
or \U$41599 ( \41976 , \41973 , \41657 );
xor \U$41600 ( \41977 , \41593 , \41595 );
xor \U$41601 ( \41978 , \41977 , \41598 );
xor \U$41602 ( \41979 , \41433 , \41459 );
xor \U$41603 ( \41980 , \41979 , \41486 );
xor \U$41604 ( \41981 , \41515 , \41540 );
xor \U$41605 ( \41982 , \41981 , \41559 );
or \U$41606 ( \41983 , \41980 , \41982 );
not \U$41607 ( \41984 , \41982 );
not \U$41608 ( \41985 , \41980 );
or \U$41609 ( \41986 , \41984 , \41985 );
xor \U$41610 ( \41987 , \41354 , \41381 );
xor \U$41611 ( \41988 , \41987 , \41409 );
nand \U$41612 ( \41989 , \41986 , \41988 );
nand \U$41613 ( \41990 , \41983 , \41989 );
xor \U$41614 ( \41991 , \40961 , \40963 );
xor \U$41615 ( \41992 , \41991 , \40966 );
xor \U$41616 ( \41993 , \41570 , \41577 );
xor \U$41617 ( \41994 , \41992 , \41993 );
xor \U$41618 ( \41995 , \41990 , \41994 );
xor \U$41619 ( \41996 , \41978 , \41995 );
nand \U$41620 ( \41997 , \41976 , \41996 );
nand \U$41621 ( \41998 , \41975 , \41997 );
not \U$41622 ( \41999 , \41988 );
not \U$41623 ( \42000 , \41982 );
or \U$41624 ( \42001 , \41999 , \42000 );
or \U$41625 ( \42002 , \41982 , \41988 );
nand \U$41626 ( \42003 , \42001 , \42002 );
not \U$41627 ( \42004 , \42003 );
not \U$41628 ( \42005 , \41980 );
and \U$41629 ( \42006 , \42004 , \42005 );
and \U$41630 ( \42007 , \42003 , \41980 );
nor \U$41631 ( \42008 , \42006 , \42007 );
not \U$41632 ( \42009 , \41789 );
not \U$41633 ( \42010 , \41760 );
or \U$41634 ( \42011 , \42009 , \42010 );
or \U$41635 ( \42012 , \41760 , \41789 );
nand \U$41636 ( \42013 , \42011 , \42012 );
not \U$41637 ( \42014 , \42013 );
not \U$41638 ( \42015 , \41733 );
and \U$41639 ( \42016 , \42014 , \42015 );
and \U$41640 ( \42017 , \42013 , \41733 );
nor \U$41641 ( \42018 , \42016 , \42017 );
not \U$41642 ( \42019 , \42018 );
xor \U$41643 ( \42020 , \41896 , \41921 );
xor \U$41644 ( \42021 , \42020 , \41947 );
not \U$41645 ( \42022 , \42021 );
and \U$41646 ( \42023 , \42019 , \42022 );
and \U$41647 ( \42024 , \42021 , \42018 );
xor \U$41648 ( \42025 , \41812 , \41838 );
xor \U$41649 ( \42026 , \42025 , \41865 );
nor \U$41650 ( \42027 , \42024 , \42026 );
nor \U$41651 ( \42028 , \42023 , \42027 );
xor \U$41652 ( \42029 , \42008 , \42028 );
xnor \U$41653 ( \42030 , \41970 , \41958 );
not \U$41654 ( \42031 , \42030 );
not \U$41655 ( \42032 , \41963 );
and \U$41656 ( \42033 , \42031 , \42032 );
and \U$41657 ( \42034 , \42030 , \41963 );
nor \U$41658 ( \42035 , \42033 , \42034 );
and \U$41659 ( \42036 , \42029 , \42035 );
and \U$41660 ( \42037 , \42008 , \42028 );
or \U$41661 ( \42038 , \42036 , \42037 );
xor \U$41662 ( \42039 , \41791 , \41868 );
xor \U$41663 ( \42040 , \42039 , \41950 );
not \U$41664 ( \42041 , \42040 );
not \U$41665 ( \42042 , \41706 );
not \U$41666 ( \42043 , \41682 );
or \U$41667 ( \42044 , \42042 , \42043 );
or \U$41668 ( \42045 , \41682 , \41706 );
nand \U$41669 ( \42046 , \42044 , \42045 );
not \U$41670 ( \42047 , \42046 );
not \U$41671 ( \42048 , \41670 );
and \U$41672 ( \42049 , \42047 , \42048 );
and \U$41673 ( \42050 , \42046 , \41670 );
nor \U$41674 ( \42051 , \42049 , \42050 );
nor \U$41675 ( \42052 , \42041 , \42051 );
not \U$41676 ( \42053 , \42052 );
or \U$41677 ( \42054 , \42038 , \42053 );
not \U$41678 ( \42055 , \42053 );
not \U$41679 ( \42056 , \42038 );
or \U$41680 ( \42057 , \42055 , \42056 );
and \U$41681 ( \42058 , \4247 , RIae75830_16);
and \U$41682 ( \42059 , RIae75740_14, \4245 );
nor \U$41683 ( \42060 , \42058 , \42059 );
and \U$41684 ( \42061 , \42060 , \3989 );
not \U$41685 ( \42062 , \42060 );
and \U$41686 ( \42063 , \42062 , \4251 );
nor \U$41687 ( \42064 , \42061 , \42063 );
and \U$41688 ( \42065 , \4688 , RIae75290_4);
and \U$41689 ( \42066 , RIae751a0_2, \4686 );
nor \U$41690 ( \42067 , \42065 , \42066 );
and \U$41691 ( \42068 , \42067 , \4481 );
not \U$41692 ( \42069 , \42067 );
and \U$41693 ( \42070 , \42069 , \4482 );
nor \U$41694 ( \42071 , \42068 , \42070 );
xor \U$41695 ( \42072 , \42064 , \42071 );
and \U$41696 ( \42073 , \5399 , RIae75380_6);
and \U$41697 ( \42074 , RIae75470_8, \5397 );
nor \U$41698 ( \42075 , \42073 , \42074 );
and \U$41699 ( \42076 , \42075 , \5016 );
not \U$41700 ( \42077 , \42075 );
and \U$41701 ( \42078 , \42077 , \5403 );
nor \U$41702 ( \42079 , \42076 , \42078 );
and \U$41703 ( \42080 , \42072 , \42079 );
and \U$41704 ( \42081 , \42064 , \42071 );
or \U$41705 ( \42082 , \42080 , \42081 );
and \U$41706 ( \42083 , \3730 , RIae75650_12);
and \U$41707 ( \42084 , RIae75560_10, \3728 );
nor \U$41708 ( \42085 , \42083 , \42084 );
and \U$41709 ( \42086 , \42085 , \3732 );
not \U$41710 ( \42087 , \42085 );
and \U$41711 ( \42088 , \42087 , \3422 );
nor \U$41712 ( \42089 , \42086 , \42088 );
not \U$41713 ( \42090 , \2789 );
and \U$41714 ( \42091 , \2783 , RIae75fb0_32);
and \U$41715 ( \42092 , RIae75ec0_30, \2781 );
nor \U$41716 ( \42093 , \42091 , \42092 );
not \U$41717 ( \42094 , \42093 );
or \U$41718 ( \42095 , \42090 , \42094 );
or \U$41719 ( \42096 , \42093 , \2789 );
nand \U$41720 ( \42097 , \42095 , \42096 );
xor \U$41721 ( \42098 , \42089 , \42097 );
not \U$41722 ( \42099 , \3218 );
and \U$41723 ( \42100 , \3214 , RIae75ce0_26);
and \U$41724 ( \42101 , RIae75dd0_28, \3212 );
nor \U$41725 ( \42102 , \42100 , \42101 );
not \U$41726 ( \42103 , \42102 );
or \U$41727 ( \42104 , \42099 , \42103 );
or \U$41728 ( \42105 , \42102 , \3218 );
nand \U$41729 ( \42106 , \42104 , \42105 );
and \U$41730 ( \42107 , \42098 , \42106 );
and \U$41731 ( \42108 , \42089 , \42097 );
or \U$41732 ( \42109 , \42107 , \42108 );
xor \U$41733 ( \42110 , \42082 , \42109 );
and \U$41734 ( \42111 , \2224 , RIae75bf0_24);
and \U$41735 ( \42112 , RIae75b00_22, \2222 );
nor \U$41736 ( \42113 , \42111 , \42112 );
and \U$41737 ( \42114 , \42113 , \2061 );
not \U$41738 ( \42115 , \42113 );
and \U$41739 ( \42116 , \42115 , \2060 );
nor \U$41740 ( \42117 , \42114 , \42116 );
and \U$41741 ( \42118 , \1939 , RIae78800_118);
and \U$41742 ( \42119 , RIae78710_116, \1937 );
nor \U$41743 ( \42120 , \42118 , \42119 );
and \U$41744 ( \42121 , \42120 , \1735 );
not \U$41745 ( \42122 , \42120 );
and \U$41746 ( \42123 , \42122 , \1734 );
nor \U$41747 ( \42124 , \42121 , \42123 );
xor \U$41748 ( \42125 , \42117 , \42124 );
and \U$41749 ( \42126 , \2607 , RIae75a10_20);
and \U$41750 ( \42127 , RIae75920_18, \2605 );
nor \U$41751 ( \42128 , \42126 , \42127 );
and \U$41752 ( \42129 , \42128 , \2611 );
not \U$41753 ( \42130 , \42128 );
and \U$41754 ( \42131 , \42130 , \2396 );
nor \U$41755 ( \42132 , \42129 , \42131 );
and \U$41756 ( \42133 , \42125 , \42132 );
and \U$41757 ( \42134 , \42117 , \42124 );
or \U$41758 ( \42135 , \42133 , \42134 );
and \U$41759 ( \42136 , \42110 , \42135 );
and \U$41760 ( \42137 , \42082 , \42109 );
nor \U$41761 ( \42138 , \42136 , \42137 );
and \U$41762 ( \42139 , \8966 , RIae76820_50);
and \U$41763 ( \42140 , RIae76910_52, \8964 );
nor \U$41764 ( \42141 , \42139 , \42140 );
and \U$41765 ( \42142 , \42141 , \8799 );
not \U$41766 ( \42143 , \42141 );
and \U$41767 ( \42144 , \42143 , \8789 );
nor \U$41768 ( \42145 , \42142 , \42144 );
and \U$41769 ( \42146 , \7633 , RIae76370_40);
and \U$41770 ( \42147 , RIae76280_38, \7631 );
nor \U$41771 ( \42148 , \42146 , \42147 );
and \U$41772 ( \42149 , \42148 , \7206 );
not \U$41773 ( \42150 , \42148 );
and \U$41774 ( \42151 , \42150 , \7205 );
nor \U$41775 ( \42152 , \42149 , \42151 );
xor \U$41776 ( \42153 , \42145 , \42152 );
and \U$41777 ( \42154 , \8371 , RIae76af0_56);
and \U$41778 ( \42155 , RIae76a00_54, \8369 );
nor \U$41779 ( \42156 , \42154 , \42155 );
and \U$41780 ( \42157 , \42156 , \8020 );
not \U$41781 ( \42158 , \42156 );
and \U$41782 ( \42159 , \42158 , \8019 );
nor \U$41783 ( \42160 , \42157 , \42159 );
and \U$41784 ( \42161 , \42153 , \42160 );
and \U$41785 ( \42162 , \42145 , \42152 );
or \U$41786 ( \42163 , \42161 , \42162 );
and \U$41787 ( \42164 , \9760 , RIae76be0_58);
and \U$41788 ( \42165 , RIae78ad0_124, \9758 );
nor \U$41789 ( \42166 , \42164 , \42165 );
and \U$41790 ( \42167 , \42166 , \9273 );
not \U$41791 ( \42168 , \42166 );
and \U$41792 ( \42169 , \42168 , \9764 );
nor \U$41793 ( \42170 , \42167 , \42169 );
xor \U$41794 ( \42171 , \42170 , \10936 );
and \U$41795 ( \42172 , \10548 , RIae78d28_129);
and \U$41796 ( \42173 , RIae78e18_131, \10546 );
nor \U$41797 ( \42174 , \42172 , \42173 );
and \U$41798 ( \42175 , \42174 , \10421 );
not \U$41799 ( \42176 , \42174 );
and \U$41800 ( \42177 , \42176 , \10118 );
nor \U$41801 ( \42178 , \42175 , \42177 );
and \U$41802 ( \42179 , \42171 , \42178 );
and \U$41803 ( \42180 , \42170 , \10936 );
or \U$41804 ( \42181 , \42179 , \42180 );
xor \U$41805 ( \42182 , \42163 , \42181 );
and \U$41806 ( \42183 , \6172 , RIae76730_48);
and \U$41807 ( \42184 , RIae76640_46, \6170 );
nor \U$41808 ( \42185 , \42183 , \42184 );
and \U$41809 ( \42186 , \42185 , \6176 );
not \U$41810 ( \42187 , \42185 );
and \U$41811 ( \42188 , \42187 , \6175 );
nor \U$41812 ( \42189 , \42186 , \42188 );
and \U$41813 ( \42190 , \5896 , RIae76460_42);
and \U$41814 ( \42191 , RIae76550_44, \5894 );
nor \U$41815 ( \42192 , \42190 , \42191 );
and \U$41816 ( \42193 , \42192 , \5590 );
not \U$41817 ( \42194 , \42192 );
and \U$41818 ( \42195 , \42194 , \5589 );
nor \U$41819 ( \42196 , \42193 , \42195 );
xor \U$41820 ( \42197 , \42189 , \42196 );
and \U$41821 ( \42198 , \6941 , RIae76190_36);
and \U$41822 ( \42199 , RIae760a0_34, \6939 );
nor \U$41823 ( \42200 , \42198 , \42199 );
and \U$41824 ( \42201 , \42200 , \6314 );
not \U$41825 ( \42202 , \42200 );
and \U$41826 ( \42203 , \42202 , \6945 );
nor \U$41827 ( \42204 , \42201 , \42203 );
and \U$41828 ( \42205 , \42197 , \42204 );
and \U$41829 ( \42206 , \42189 , \42196 );
or \U$41830 ( \42207 , \42205 , \42206 );
and \U$41831 ( \42208 , \42182 , \42207 );
and \U$41832 ( \42209 , \42163 , \42181 );
nor \U$41833 ( \42210 , \42208 , \42209 );
xor \U$41834 ( \42211 , \42138 , \42210 );
and \U$41835 ( \42212 , \1593 , RIae789e0_122);
and \U$41836 ( \42213 , RIae788f0_120, \1591 );
nor \U$41837 ( \42214 , \42212 , \42213 );
and \U$41838 ( \42215 , \42214 , \1498 );
not \U$41839 ( \42216 , \42214 );
and \U$41840 ( \42217 , \42216 , \1488 );
nor \U$41841 ( \42218 , \42215 , \42217 );
and \U$41842 ( \42219 , \1138 , RIae77cc0_94);
and \U$41843 ( \42220 , RIae77bd0_92, \1136 );
nor \U$41844 ( \42221 , \42219 , \42220 );
and \U$41845 ( \42222 , \42221 , \1012 );
not \U$41846 ( \42223 , \42221 );
and \U$41847 ( \42224 , \42223 , \1142 );
nor \U$41848 ( \42225 , \42222 , \42224 );
xor \U$41849 ( \42226 , \42218 , \42225 );
and \U$41850 ( \42227 , \1376 , RIae77db0_96);
and \U$41851 ( \42228 , RIae77ea0_98, \1374 );
nor \U$41852 ( \42229 , \42227 , \42228 );
and \U$41853 ( \42230 , \42229 , \1380 );
not \U$41854 ( \42231 , \42229 );
and \U$41855 ( \42232 , \42231 , \1261 );
nor \U$41856 ( \42233 , \42230 , \42232 );
and \U$41857 ( \42234 , \42226 , \42233 );
and \U$41858 ( \42235 , \42218 , \42225 );
or \U$41859 ( \42236 , \42234 , \42235 );
not \U$41860 ( \42237 , \392 );
and \U$41861 ( \42238 , \384 , RIae77108_69);
and \U$41862 ( \42239 , RIae77090_68, \382 );
nor \U$41863 ( \42240 , \42238 , \42239 );
not \U$41864 ( \42241 , \42240 );
or \U$41865 ( \42242 , \42237 , \42241 );
or \U$41866 ( \42243 , \42240 , \388 );
nand \U$41867 ( \42244 , \42242 , \42243 );
not \U$41868 ( \42245 , \400 );
and \U$41869 ( \42246 , \436 , RIae77270_72);
and \U$41870 ( \42247 , RIae77360_74, \434 );
nor \U$41871 ( \42248 , \42246 , \42247 );
not \U$41872 ( \42249 , \42248 );
or \U$41873 ( \42250 , \42245 , \42249 );
or \U$41874 ( \42251 , \42248 , \402 );
nand \U$41875 ( \42252 , \42250 , \42251 );
xor \U$41876 ( \42253 , \42244 , \42252 );
not \U$41877 ( \42254 , \469 );
and \U$41878 ( \42255 , \514 , RIae78350_108);
and \U$41879 ( \42256 , RIae78170_104, \512 );
nor \U$41880 ( \42257 , \42255 , \42256 );
not \U$41881 ( \42258 , \42257 );
or \U$41882 ( \42259 , \42254 , \42258 );
or \U$41883 ( \42260 , \42257 , \471 );
nand \U$41884 ( \42261 , \42259 , \42260 );
and \U$41885 ( \42262 , \42253 , \42261 );
and \U$41886 ( \42263 , \42244 , \42252 );
or \U$41887 ( \42264 , \42262 , \42263 );
xor \U$41888 ( \42265 , \42236 , \42264 );
and \U$41889 ( \42266 , \672 , RIae78260_106);
and \U$41890 ( \42267 , RIae78620_114, \670 );
nor \U$41891 ( \42268 , \42266 , \42267 );
and \U$41892 ( \42269 , \42268 , \588 );
not \U$41893 ( \42270 , \42268 );
and \U$41894 ( \42271 , \42270 , \587 );
nor \U$41895 ( \42272 , \42269 , \42271 );
and \U$41896 ( \42273 , \558 , RIae77f90_100);
and \U$41897 ( \42274 , RIae78080_102, \556 );
nor \U$41898 ( \42275 , \42273 , \42274 );
and \U$41899 ( \42276 , \42275 , \504 );
not \U$41900 ( \42277 , \42275 );
and \U$41901 ( \42278 , \42277 , \562 );
nor \U$41902 ( \42279 , \42276 , \42278 );
xor \U$41903 ( \42280 , \42272 , \42279 );
not \U$41904 ( \42281 , \789 );
and \U$41905 ( \42282 , \883 , RIae78440_110);
and \U$41906 ( \42283 , RIae784b8_111, \881 );
nor \U$41907 ( \42284 , \42282 , \42283 );
not \U$41908 ( \42285 , \42284 );
or \U$41909 ( \42286 , \42281 , \42285 );
or \U$41910 ( \42287 , \42284 , \789 );
nand \U$41911 ( \42288 , \42286 , \42287 );
and \U$41912 ( \42289 , \42280 , \42288 );
and \U$41913 ( \42290 , \42272 , \42279 );
or \U$41914 ( \42291 , \42289 , \42290 );
and \U$41915 ( \42292 , \42265 , \42291 );
and \U$41916 ( \42293 , \42236 , \42264 );
nor \U$41917 ( \42294 , \42292 , \42293 );
and \U$41918 ( \42295 , \42211 , \42294 );
and \U$41919 ( \42296 , \42138 , \42210 );
or \U$41920 ( \42297 , \42295 , \42296 );
xor \U$41921 ( \42298 , \41799 , \41800 );
xor \U$41922 ( \42299 , \42298 , \41809 );
xor \U$41923 ( \42300 , \41847 , \41854 );
xor \U$41924 ( \42301 , \42300 , \41862 );
nand \U$41925 ( \42302 , \42299 , \42301 );
xor \U$41926 ( \42303 , \41903 , \41910 );
xor \U$41927 ( \42304 , \42303 , \41918 );
xor \U$41928 ( \42305 , \41771 , \41778 );
xor \U$41929 ( \42306 , \42305 , \41786 );
and \U$41930 ( \42307 , \42304 , \42306 );
not \U$41931 ( \42308 , \41740 );
xor \U$41932 ( \42309 , \41748 , \41758 );
not \U$41933 ( \42310 , \42309 );
or \U$41934 ( \42311 , \42308 , \42310 );
or \U$41935 ( \42312 , \42309 , \41740 );
nand \U$41936 ( \42313 , \42311 , \42312 );
xor \U$41937 ( \42314 , \41771 , \41778 );
xor \U$41938 ( \42315 , \42314 , \41786 );
and \U$41939 ( \42316 , \42313 , \42315 );
and \U$41940 ( \42317 , \42304 , \42313 );
or \U$41941 ( \42318 , \42307 , \42316 , \42317 );
xor \U$41942 ( \42319 , \42302 , \42318 );
xor \U$41943 ( \42320 , \41819 , \41826 );
xor \U$41944 ( \42321 , \42320 , \41835 );
xor \U$41945 ( \42322 , \41929 , \41936 );
xor \U$41946 ( \42323 , \42322 , \41944 );
xor \U$41947 ( \42324 , \42321 , \42323 );
xor \U$41948 ( \42325 , \41877 , \41885 );
xor \U$41949 ( \42326 , \42325 , \41893 );
and \U$41950 ( \42327 , \42324 , \42326 );
and \U$41951 ( \42328 , \42321 , \42323 );
or \U$41952 ( \42329 , \42327 , \42328 );
and \U$41953 ( \42330 , \42319 , \42329 );
and \U$41954 ( \42331 , \42302 , \42318 );
nor \U$41955 ( \42332 , \42330 , \42331 );
xor \U$41956 ( \42333 , \42297 , \42332 );
not \U$41957 ( \42334 , \41698 );
not \U$41958 ( \42335 , \41704 );
or \U$41959 ( \42336 , \42334 , \42335 );
or \U$41960 ( \42337 , \41698 , \41704 );
nand \U$41961 ( \42338 , \42336 , \42337 );
not \U$41962 ( \42339 , \42338 );
not \U$41963 ( \42340 , \41696 );
and \U$41964 ( \42341 , \42339 , \42340 );
and \U$41965 ( \42342 , \42338 , \41696 );
nor \U$41966 ( \42343 , \42341 , \42342 );
xor \U$41967 ( \42344 , \41441 , \41448 );
xor \U$41968 ( \42345 , \42344 , \41456 );
xor \U$41969 ( \42346 , \41672 , \41677 );
xor \U$41970 ( \42347 , \42345 , \42346 );
xor \U$41971 ( \42348 , \42343 , \42347 );
xor \U$41972 ( \42349 , \41497 , \41504 );
xor \U$41973 ( \42350 , \42349 , \41512 );
xor \U$41974 ( \42351 , \41660 , \41665 );
xor \U$41975 ( \42352 , \42350 , \42351 );
and \U$41976 ( \42353 , \42348 , \42352 );
and \U$41977 ( \42354 , \42343 , \42347 );
or \U$41978 ( \42355 , \42353 , \42354 );
and \U$41979 ( \42356 , \42333 , \42355 );
and \U$41980 ( \42357 , \42297 , \42332 );
nor \U$41981 ( \42358 , \42356 , \42357 );
nand \U$41982 ( \42359 , \42057 , \42358 );
nand \U$41983 ( \42360 , \42054 , \42359 );
xor \U$41984 ( \42361 , \41998 , \42360 );
xor \U$41985 ( \42362 , \41329 , \41565 );
xor \U$41986 ( \42363 , \42362 , \41582 );
xor \U$41987 ( \42364 , \41587 , \41589 );
xor \U$41988 ( \42365 , \41229 , \41231 );
xor \U$41989 ( \42366 , \42365 , \41234 );
xor \U$41990 ( \42367 , \41601 , \41608 );
xor \U$41991 ( \42368 , \42366 , \42367 );
xor \U$41992 ( \42369 , \42364 , \42368 );
xor \U$41993 ( \42370 , \42363 , \42369 );
and \U$41994 ( \42371 , \42361 , \42370 );
and \U$41995 ( \42372 , \41998 , \42360 );
or \U$41996 ( \42373 , \42371 , \42372 );
xor \U$41997 ( \42374 , \41585 , \41590 );
xor \U$41998 ( \42375 , \42374 , \41613 );
xor \U$41999 ( \42376 , \42373 , \42375 );
xor \U$42000 ( \42377 , \41708 , \41953 );
and \U$42001 ( \42378 , \42377 , \41972 );
and \U$42002 ( \42379 , \41708 , \41953 );
or \U$42003 ( \42380 , \42378 , \42379 );
and \U$42004 ( \42381 , \41654 , \41656 );
xor \U$42005 ( \42382 , \42380 , \42381 );
xor \U$42006 ( \42383 , \41593 , \41595 );
xor \U$42007 ( \42384 , \42383 , \41598 );
and \U$42008 ( \42385 , \41990 , \42384 );
xor \U$42009 ( \42386 , \41593 , \41595 );
xor \U$42010 ( \42387 , \42386 , \41598 );
and \U$42011 ( \42388 , \41994 , \42387 );
and \U$42012 ( \42389 , \41990 , \41994 );
or \U$42013 ( \42390 , \42385 , \42388 , \42389 );
and \U$42014 ( \42391 , \42382 , \42390 );
and \U$42015 ( \42392 , \42380 , \42381 );
or \U$42016 ( \42393 , \42391 , \42392 );
xor \U$42017 ( \42394 , \41329 , \41565 );
xor \U$42018 ( \42395 , \42394 , \41582 );
and \U$42019 ( \42396 , \42364 , \42395 );
xor \U$42020 ( \42397 , \41329 , \41565 );
xor \U$42021 ( \42398 , \42397 , \41582 );
and \U$42022 ( \42399 , \42368 , \42398 );
and \U$42023 ( \42400 , \42364 , \42368 );
or \U$42024 ( \42401 , \42396 , \42399 , \42400 );
xor \U$42025 ( \42402 , \42393 , \42401 );
xor \U$42026 ( \42403 , \40972 , \41201 );
xor \U$42027 ( \42404 , \42403 , \41218 );
xor \U$42028 ( \42405 , \41617 , \41624 );
xor \U$42029 ( \42406 , \42404 , \42405 );
xor \U$42030 ( \42407 , \42402 , \42406 );
and \U$42031 ( \42408 , \42376 , \42407 );
and \U$42032 ( \42409 , \42373 , \42375 );
or \U$42033 ( \42410 , \42408 , \42409 );
xor \U$42034 ( \42411 , \42393 , \42401 );
and \U$42035 ( \42412 , \42411 , \42406 );
and \U$42036 ( \42413 , \42393 , \42401 );
or \U$42037 ( \42414 , \42412 , \42413 );
xor \U$42038 ( \42415 , \41221 , \41226 );
xor \U$42039 ( \42416 , \42415 , \41247 );
xor \U$42040 ( \42417 , \42414 , \42416 );
xor \U$42041 ( \42418 , \41616 , \41629 );
xor \U$42042 ( \42419 , \42418 , \41634 );
xor \U$42043 ( \42420 , \42417 , \42419 );
and \U$42044 ( \42421 , \42410 , \42420 );
not \U$42045 ( \42422 , \42421 );
xor \U$42046 ( \42423 , \42414 , \42416 );
and \U$42047 ( \42424 , \42423 , \42419 );
and \U$42048 ( \42425 , \42414 , \42416 );
or \U$42049 ( \42426 , \42424 , \42425 );
xor \U$42050 ( \42427 , \41637 , \41639 );
xor \U$42051 ( \42428 , \42427 , \41646 );
xor \U$42052 ( \42429 , \42426 , \42428 );
not \U$42053 ( \42430 , \42429 );
or \U$42054 ( \42431 , \42422 , \42430 );
xor \U$42055 ( \42432 , \42410 , \42420 );
xor \U$42056 ( \42433 , \42373 , \42375 );
xor \U$42057 ( \42434 , \42433 , \42407 );
not \U$42058 ( \42435 , \42434 );
xor \U$42059 ( \42436 , \41998 , \42360 );
xor \U$42060 ( \42437 , \42436 , \42370 );
xor \U$42061 ( \42438 , \42380 , \42381 );
xor \U$42062 ( \42439 , \42438 , \42390 );
and \U$42063 ( \42440 , \42437 , \42439 );
not \U$42064 ( \42441 , \42437 );
not \U$42065 ( \42442 , \42439 );
and \U$42066 ( \42443 , \42441 , \42442 );
xor \U$42067 ( \42444 , \42297 , \42332 );
xor \U$42068 ( \42445 , \42444 , \42355 );
not \U$42069 ( \42446 , \42051 );
not \U$42070 ( \42447 , \42040 );
and \U$42071 ( \42448 , \42446 , \42447 );
and \U$42072 ( \42449 , \42051 , \42040 );
nor \U$42073 ( \42450 , \42448 , \42449 );
xor \U$42074 ( \42451 , \42445 , \42450 );
xor \U$42075 ( \42452 , \42008 , \42028 );
xor \U$42076 ( \42453 , \42452 , \42035 );
and \U$42077 ( \42454 , \42451 , \42453 );
and \U$42078 ( \42455 , \42445 , \42450 );
or \U$42079 ( \42456 , \42454 , \42455 );
xor \U$42080 ( \42457 , \42064 , \42071 );
xor \U$42081 ( \42458 , \42457 , \42079 );
xor \U$42082 ( \42459 , \42189 , \42196 );
xor \U$42083 ( \42460 , \42459 , \42204 );
and \U$42084 ( \42461 , \42458 , \42460 );
xor \U$42085 ( \42462 , \42145 , \42152 );
xor \U$42086 ( \42463 , \42462 , \42160 );
xor \U$42087 ( \42464 , \42189 , \42196 );
xor \U$42088 ( \42465 , \42464 , \42204 );
and \U$42089 ( \42466 , \42463 , \42465 );
and \U$42090 ( \42467 , \42458 , \42463 );
or \U$42091 ( \42468 , \42461 , \42466 , \42467 );
not \U$42092 ( \42469 , RIae76cd0_60);
nor \U$42093 ( \42470 , \42469 , \491 );
xor \U$42094 ( \42471 , \42272 , \42279 );
xor \U$42095 ( \42472 , \42471 , \42288 );
and \U$42096 ( \42473 , \42470 , \42472 );
xor \U$42097 ( \42474 , \42244 , \42252 );
xor \U$42098 ( \42475 , \42474 , \42261 );
xor \U$42099 ( \42476 , \42272 , \42279 );
xor \U$42100 ( \42477 , \42476 , \42288 );
and \U$42101 ( \42478 , \42475 , \42477 );
and \U$42102 ( \42479 , \42470 , \42475 );
or \U$42103 ( \42480 , \42473 , \42478 , \42479 );
xor \U$42104 ( \42481 , \42468 , \42480 );
xor \U$42105 ( \42482 , \42218 , \42225 );
xor \U$42106 ( \42483 , \42482 , \42233 );
xor \U$42107 ( \42484 , \42117 , \42124 );
xor \U$42108 ( \42485 , \42484 , \42132 );
xor \U$42109 ( \42486 , \42483 , \42485 );
xor \U$42110 ( \42487 , \42089 , \42097 );
xor \U$42111 ( \42488 , \42487 , \42106 );
and \U$42112 ( \42489 , \42486 , \42488 );
and \U$42113 ( \42490 , \42483 , \42485 );
or \U$42114 ( \42491 , \42489 , \42490 );
and \U$42115 ( \42492 , \42481 , \42491 );
and \U$42116 ( \42493 , \42468 , \42480 );
or \U$42117 ( \42494 , \42492 , \42493 );
and \U$42118 ( \42495 , \672 , RIae78080_102);
and \U$42119 ( \42496 , RIae78260_106, \670 );
nor \U$42120 ( \42497 , \42495 , \42496 );
and \U$42121 ( \42498 , \42497 , \588 );
not \U$42122 ( \42499 , \42497 );
and \U$42123 ( \42500 , \42499 , \587 );
nor \U$42124 ( \42501 , \42498 , \42500 );
and \U$42125 ( \42502 , \558 , RIae78170_104);
and \U$42126 ( \42503 , RIae77f90_100, \556 );
nor \U$42127 ( \42504 , \42502 , \42503 );
and \U$42128 ( \42505 , \42504 , \504 );
not \U$42129 ( \42506 , \42504 );
and \U$42130 ( \42507 , \42506 , \562 );
nor \U$42131 ( \42508 , \42505 , \42507 );
xor \U$42132 ( \42509 , \42501 , \42508 );
not \U$42133 ( \42510 , \789 );
and \U$42134 ( \42511 , \883 , RIae78620_114);
and \U$42135 ( \42512 , RIae78440_110, \881 );
nor \U$42136 ( \42513 , \42511 , \42512 );
not \U$42137 ( \42514 , \42513 );
or \U$42138 ( \42515 , \42510 , \42514 );
or \U$42139 ( \42516 , \42513 , \789 );
nand \U$42140 ( \42517 , \42515 , \42516 );
and \U$42141 ( \42518 , \42509 , \42517 );
and \U$42142 ( \42519 , \42501 , \42508 );
or \U$42143 ( \42520 , \42518 , \42519 );
and \U$42144 ( \42521 , \384 , RIae76cd0_60);
and \U$42145 ( \42522 , RIae77108_69, \382 );
nor \U$42146 ( \42523 , \42521 , \42522 );
not \U$42147 ( \42524 , \42523 );
not \U$42148 ( \42525 , \392 );
and \U$42149 ( \42526 , \42524 , \42525 );
and \U$42150 ( \42527 , \42523 , \388 );
nor \U$42151 ( \42528 , \42526 , \42527 );
and \U$42152 ( \42529 , \436 , RIae77090_68);
and \U$42153 ( \42530 , RIae77270_72, \434 );
nor \U$42154 ( \42531 , \42529 , \42530 );
not \U$42155 ( \42532 , \42531 );
not \U$42156 ( \42533 , \402 );
and \U$42157 ( \42534 , \42532 , \42533 );
and \U$42158 ( \42535 , \42531 , \402 );
nor \U$42159 ( \42536 , \42534 , \42535 );
or \U$42160 ( \42537 , \42528 , \42536 );
not \U$42161 ( \42538 , \42536 );
not \U$42162 ( \42539 , \42528 );
or \U$42163 ( \42540 , \42538 , \42539 );
not \U$42164 ( \42541 , \471 );
and \U$42165 ( \42542 , \514 , RIae77360_74);
and \U$42166 ( \42543 , RIae78350_108, \512 );
nor \U$42167 ( \42544 , \42542 , \42543 );
not \U$42168 ( \42545 , \42544 );
or \U$42169 ( \42546 , \42541 , \42545 );
or \U$42170 ( \42547 , \42544 , \471 );
nand \U$42171 ( \42548 , \42546 , \42547 );
nand \U$42172 ( \42549 , \42540 , \42548 );
nand \U$42173 ( \42550 , \42537 , \42549 );
xor \U$42174 ( \42551 , \42520 , \42550 );
and \U$42175 ( \42552 , \1593 , RIae77ea0_98);
and \U$42176 ( \42553 , RIae789e0_122, \1591 );
nor \U$42177 ( \42554 , \42552 , \42553 );
and \U$42178 ( \42555 , \42554 , \1498 );
not \U$42179 ( \42556 , \42554 );
and \U$42180 ( \42557 , \42556 , \1488 );
nor \U$42181 ( \42558 , \42555 , \42557 );
and \U$42182 ( \42559 , \1138 , RIae784b8_111);
and \U$42183 ( \42560 , RIae77cc0_94, \1136 );
nor \U$42184 ( \42561 , \42559 , \42560 );
and \U$42185 ( \42562 , \42561 , \1012 );
not \U$42186 ( \42563 , \42561 );
and \U$42187 ( \42564 , \42563 , \1142 );
nor \U$42188 ( \42565 , \42562 , \42564 );
xor \U$42189 ( \42566 , \42558 , \42565 );
and \U$42190 ( \42567 , \1376 , RIae77bd0_92);
and \U$42191 ( \42568 , RIae77db0_96, \1374 );
nor \U$42192 ( \42569 , \42567 , \42568 );
and \U$42193 ( \42570 , \42569 , \1380 );
not \U$42194 ( \42571 , \42569 );
and \U$42195 ( \42572 , \42571 , \1261 );
nor \U$42196 ( \42573 , \42570 , \42572 );
and \U$42197 ( \42574 , \42566 , \42573 );
and \U$42198 ( \42575 , \42558 , \42565 );
or \U$42199 ( \42576 , \42574 , \42575 );
and \U$42200 ( \42577 , \42551 , \42576 );
and \U$42201 ( \42578 , \42520 , \42550 );
or \U$42202 ( \42579 , \42577 , \42578 );
and \U$42203 ( \42580 , \8966 , RIae76a00_54);
and \U$42204 ( \42581 , RIae76820_50, \8964 );
nor \U$42205 ( \42582 , \42580 , \42581 );
and \U$42206 ( \42583 , \42582 , \8799 );
not \U$42207 ( \42584 , \42582 );
and \U$42208 ( \42585 , \42584 , \8789 );
nor \U$42209 ( \42586 , \42583 , \42585 );
and \U$42210 ( \42587 , \7633 , RIae760a0_34);
and \U$42211 ( \42588 , RIae76370_40, \7631 );
nor \U$42212 ( \42589 , \42587 , \42588 );
and \U$42213 ( \42590 , \42589 , \7206 );
not \U$42214 ( \42591 , \42589 );
and \U$42215 ( \42592 , \42591 , \7205 );
nor \U$42216 ( \42593 , \42590 , \42592 );
xor \U$42217 ( \42594 , \42586 , \42593 );
and \U$42218 ( \42595 , \8371 , RIae76280_38);
and \U$42219 ( \42596 , RIae76af0_56, \8369 );
nor \U$42220 ( \42597 , \42595 , \42596 );
and \U$42221 ( \42598 , \42597 , \8020 );
not \U$42222 ( \42599 , \42597 );
and \U$42223 ( \42600 , \42599 , \8019 );
nor \U$42224 ( \42601 , \42598 , \42600 );
and \U$42225 ( \42602 , \42594 , \42601 );
and \U$42226 ( \42603 , \42586 , \42593 );
or \U$42227 ( \42604 , \42602 , \42603 );
and \U$42228 ( \42605 , \9760 , RIae76910_52);
and \U$42229 ( \42606 , RIae76be0_58, \9758 );
nor \U$42230 ( \42607 , \42605 , \42606 );
and \U$42231 ( \42608 , \42607 , \9273 );
not \U$42232 ( \42609 , \42607 );
and \U$42233 ( \42610 , \42609 , \9764 );
nor \U$42234 ( \42611 , \42608 , \42610 );
nand \U$42235 ( \42612 , RIae78e18_131, \11470 );
and \U$42236 ( \42613 , \42612 , \10936 );
not \U$42237 ( \42614 , \42612 );
and \U$42238 ( \42615 , \42614 , \11474 );
nor \U$42239 ( \42616 , \42613 , \42615 );
xor \U$42240 ( \42617 , \42611 , \42616 );
and \U$42241 ( \42618 , \10548 , RIae78ad0_124);
and \U$42242 ( \42619 , RIae78d28_129, \10546 );
nor \U$42243 ( \42620 , \42618 , \42619 );
and \U$42244 ( \42621 , \42620 , \10421 );
not \U$42245 ( \42622 , \42620 );
and \U$42246 ( \42623 , \42622 , \10118 );
nor \U$42247 ( \42624 , \42621 , \42623 );
and \U$42248 ( \42625 , \42617 , \42624 );
and \U$42249 ( \42626 , \42611 , \42616 );
or \U$42250 ( \42627 , \42625 , \42626 );
xor \U$42251 ( \42628 , \42604 , \42627 );
and \U$42252 ( \42629 , \6941 , RIae76640_46);
and \U$42253 ( \42630 , RIae76190_36, \6939 );
nor \U$42254 ( \42631 , \42629 , \42630 );
and \U$42255 ( \42632 , \42631 , \6314 );
not \U$42256 ( \42633 , \42631 );
and \U$42257 ( \42634 , \42633 , \6945 );
nor \U$42258 ( \42635 , \42632 , \42634 );
and \U$42259 ( \42636 , \5896 , RIae75470_8);
and \U$42260 ( \42637 , RIae76460_42, \5894 );
nor \U$42261 ( \42638 , \42636 , \42637 );
and \U$42262 ( \42639 , \42638 , \5590 );
not \U$42263 ( \42640 , \42638 );
and \U$42264 ( \42641 , \42640 , \5589 );
nor \U$42265 ( \42642 , \42639 , \42641 );
xor \U$42266 ( \42643 , \42635 , \42642 );
and \U$42267 ( \42644 , \6172 , RIae76550_44);
and \U$42268 ( \42645 , RIae76730_48, \6170 );
nor \U$42269 ( \42646 , \42644 , \42645 );
and \U$42270 ( \42647 , \42646 , \6176 );
not \U$42271 ( \42648 , \42646 );
and \U$42272 ( \42649 , \42648 , \6175 );
nor \U$42273 ( \42650 , \42647 , \42649 );
and \U$42274 ( \42651 , \42643 , \42650 );
and \U$42275 ( \42652 , \42635 , \42642 );
or \U$42276 ( \42653 , \42651 , \42652 );
and \U$42277 ( \42654 , \42628 , \42653 );
and \U$42278 ( \42655 , \42604 , \42627 );
or \U$42279 ( \42656 , \42654 , \42655 );
xor \U$42280 ( \42657 , \42579 , \42656 );
and \U$42281 ( \42658 , \4247 , RIae75560_10);
and \U$42282 ( \42659 , RIae75830_16, \4245 );
nor \U$42283 ( \42660 , \42658 , \42659 );
and \U$42284 ( \42661 , \42660 , \3989 );
not \U$42285 ( \42662 , \42660 );
and \U$42286 ( \42663 , \42662 , \4251 );
nor \U$42287 ( \42664 , \42661 , \42663 );
and \U$42288 ( \42665 , \4688 , RIae75740_14);
and \U$42289 ( \42666 , RIae75290_4, \4686 );
nor \U$42290 ( \42667 , \42665 , \42666 );
and \U$42291 ( \42668 , \42667 , \4481 );
not \U$42292 ( \42669 , \42667 );
and \U$42293 ( \42670 , \42669 , \4482 );
nor \U$42294 ( \42671 , \42668 , \42670 );
xor \U$42295 ( \42672 , \42664 , \42671 );
and \U$42296 ( \42673 , \5399 , RIae751a0_2);
and \U$42297 ( \42674 , RIae75380_6, \5397 );
nor \U$42298 ( \42675 , \42673 , \42674 );
and \U$42299 ( \42676 , \42675 , \5016 );
not \U$42300 ( \42677 , \42675 );
and \U$42301 ( \42678 , \42677 , \5403 );
nor \U$42302 ( \42679 , \42676 , \42678 );
and \U$42303 ( \42680 , \42672 , \42679 );
and \U$42304 ( \42681 , \42664 , \42671 );
or \U$42305 ( \42682 , \42680 , \42681 );
and \U$42306 ( \42683 , \1939 , RIae788f0_120);
and \U$42307 ( \42684 , RIae78800_118, \1937 );
nor \U$42308 ( \42685 , \42683 , \42684 );
and \U$42309 ( \42686 , \42685 , \1735 );
not \U$42310 ( \42687 , \42685 );
and \U$42311 ( \42688 , \42687 , \1734 );
nor \U$42312 ( \42689 , \42686 , \42688 );
and \U$42313 ( \42690 , \2224 , RIae78710_116);
and \U$42314 ( \42691 , RIae75bf0_24, \2222 );
nor \U$42315 ( \42692 , \42690 , \42691 );
and \U$42316 ( \42693 , \42692 , \2061 );
not \U$42317 ( \42694 , \42692 );
and \U$42318 ( \42695 , \42694 , \2060 );
nor \U$42319 ( \42696 , \42693 , \42695 );
xor \U$42320 ( \42697 , \42689 , \42696 );
and \U$42321 ( \42698 , \2607 , RIae75b00_22);
and \U$42322 ( \42699 , RIae75a10_20, \2605 );
nor \U$42323 ( \42700 , \42698 , \42699 );
and \U$42324 ( \42701 , \42700 , \2611 );
not \U$42325 ( \42702 , \42700 );
and \U$42326 ( \42703 , \42702 , \2397 );
nor \U$42327 ( \42704 , \42701 , \42703 );
and \U$42328 ( \42705 , \42697 , \42704 );
and \U$42329 ( \42706 , \42689 , \42696 );
or \U$42330 ( \42707 , \42705 , \42706 );
xor \U$42331 ( \42708 , \42682 , \42707 );
and \U$42332 ( \42709 , \3730 , RIae75dd0_28);
and \U$42333 ( \42710 , RIae75650_12, \3728 );
nor \U$42334 ( \42711 , \42709 , \42710 );
and \U$42335 ( \42712 , \42711 , \3732 );
not \U$42336 ( \42713 , \42711 );
and \U$42337 ( \42714 , \42713 , \3422 );
nor \U$42338 ( \42715 , \42712 , \42714 );
not \U$42339 ( \42716 , \2789 );
and \U$42340 ( \42717 , \2783 , RIae75920_18);
and \U$42341 ( \42718 , RIae75fb0_32, \2781 );
nor \U$42342 ( \42719 , \42717 , \42718 );
not \U$42343 ( \42720 , \42719 );
or \U$42344 ( \42721 , \42716 , \42720 );
or \U$42345 ( \42722 , \42719 , \2789 );
nand \U$42346 ( \42723 , \42721 , \42722 );
xor \U$42347 ( \42724 , \42715 , \42723 );
not \U$42348 ( \42725 , \3218 );
and \U$42349 ( \42726 , \3214 , RIae75ec0_30);
and \U$42350 ( \42727 , RIae75ce0_26, \3212 );
nor \U$42351 ( \42728 , \42726 , \42727 );
not \U$42352 ( \42729 , \42728 );
or \U$42353 ( \42730 , \42725 , \42729 );
or \U$42354 ( \42731 , \42728 , \2774 );
nand \U$42355 ( \42732 , \42730 , \42731 );
and \U$42356 ( \42733 , \42724 , \42732 );
and \U$42357 ( \42734 , \42715 , \42723 );
or \U$42358 ( \42735 , \42733 , \42734 );
and \U$42359 ( \42736 , \42708 , \42735 );
and \U$42360 ( \42737 , \42682 , \42707 );
or \U$42361 ( \42738 , \42736 , \42737 );
and \U$42362 ( \42739 , \42657 , \42738 );
and \U$42363 ( \42740 , \42579 , \42656 );
or \U$42364 ( \42741 , \42739 , \42740 );
xor \U$42365 ( \42742 , \42494 , \42741 );
not \U$42366 ( \42743 , \41715 );
xor \U$42367 ( \42744 , \41731 , \41723 );
not \U$42368 ( \42745 , \42744 );
or \U$42369 ( \42746 , \42743 , \42745 );
or \U$42370 ( \42747 , \42744 , \41715 );
nand \U$42371 ( \42748 , \42746 , \42747 );
xor \U$42372 ( \42749 , \42321 , \42323 );
xor \U$42373 ( \42750 , \42749 , \42326 );
and \U$42374 ( \42751 , \42748 , \42750 );
xor \U$42375 ( \42752 , \41771 , \41778 );
xor \U$42376 ( \42753 , \42752 , \41786 );
xor \U$42377 ( \42754 , \42304 , \42313 );
xor \U$42378 ( \42755 , \42753 , \42754 );
xor \U$42379 ( \42756 , \42321 , \42323 );
xor \U$42380 ( \42757 , \42756 , \42326 );
and \U$42381 ( \42758 , \42755 , \42757 );
and \U$42382 ( \42759 , \42748 , \42755 );
or \U$42383 ( \42760 , \42751 , \42758 , \42759 );
and \U$42384 ( \42761 , \42742 , \42760 );
and \U$42385 ( \42762 , \42494 , \42741 );
nor \U$42386 ( \42763 , \42761 , \42762 );
xor \U$42387 ( \42764 , \42138 , \42210 );
xor \U$42388 ( \42765 , \42764 , \42294 );
not \U$42389 ( \42766 , \42765 );
xor \U$42390 ( \42767 , \42302 , \42318 );
xor \U$42391 ( \42768 , \42767 , \42329 );
nand \U$42392 ( \42769 , \42766 , \42768 );
xor \U$42393 ( \42770 , \42763 , \42769 );
not \U$42394 ( \42771 , \42021 );
xor \U$42395 ( \42772 , \42026 , \42018 );
not \U$42396 ( \42773 , \42772 );
or \U$42397 ( \42774 , \42771 , \42773 );
or \U$42398 ( \42775 , \42772 , \42021 );
nand \U$42399 ( \42776 , \42774 , \42775 );
xor \U$42400 ( \42777 , \42236 , \42264 );
xor \U$42401 ( \42778 , \42777 , \42291 );
or \U$42402 ( \42779 , \42299 , \42301 );
nand \U$42403 ( \42780 , \42779 , \42302 );
xor \U$42404 ( \42781 , \42778 , \42780 );
xor \U$42405 ( \42782 , \42082 , \42109 );
xor \U$42406 ( \42783 , \42782 , \42135 );
and \U$42407 ( \42784 , \42781 , \42783 );
and \U$42408 ( \42785 , \42778 , \42780 );
or \U$42409 ( \42786 , \42784 , \42785 );
and \U$42410 ( \42787 , \42776 , \42786 );
not \U$42411 ( \42788 , \42776 );
not \U$42412 ( \42789 , \42786 );
and \U$42413 ( \42790 , \42788 , \42789 );
xor \U$42414 ( \42791 , \42343 , \42347 );
xor \U$42415 ( \42792 , \42791 , \42352 );
nor \U$42416 ( \42793 , \42790 , \42792 );
nor \U$42417 ( \42794 , \42787 , \42793 );
and \U$42418 ( \42795 , \42770 , \42794 );
and \U$42419 ( \42796 , \42763 , \42769 );
or \U$42420 ( \42797 , \42795 , \42796 );
xor \U$42421 ( \42798 , \42456 , \42797 );
xnor \U$42422 ( \42799 , \41973 , \41996 );
not \U$42423 ( \42800 , \42799 );
not \U$42424 ( \42801 , \41657 );
and \U$42425 ( \42802 , \42800 , \42801 );
and \U$42426 ( \42803 , \42799 , \41657 );
nor \U$42427 ( \42804 , \42802 , \42803 );
and \U$42428 ( \42805 , \42798 , \42804 );
and \U$42429 ( \42806 , \42456 , \42797 );
or \U$42430 ( \42807 , \42805 , \42806 );
nor \U$42431 ( \42808 , \42443 , \42807 );
nor \U$42432 ( \42809 , \42440 , \42808 );
nor \U$42433 ( \42810 , \42435 , \42809 );
and \U$42434 ( \42811 , \42432 , \42810 );
xor \U$42435 ( \42812 , \42810 , \42432 );
not \U$42436 ( \42813 , \42434 );
not \U$42437 ( \42814 , \42809 );
and \U$42438 ( \42815 , \42813 , \42814 );
and \U$42439 ( \42816 , \42434 , \42809 );
nor \U$42440 ( \42817 , \42815 , \42816 );
not \U$42441 ( \42818 , \42765 );
not \U$42442 ( \42819 , \42768 );
or \U$42443 ( \42820 , \42818 , \42819 );
or \U$42444 ( \42821 , \42768 , \42765 );
nand \U$42445 ( \42822 , \42820 , \42821 );
xor \U$42446 ( \42823 , \42494 , \42741 );
xor \U$42447 ( \42824 , \42823 , \42760 );
xor \U$42448 ( \42825 , \42822 , \42824 );
not \U$42449 ( \42826 , \42792 );
xor \U$42450 ( \42827 , \42786 , \42776 );
not \U$42451 ( \42828 , \42827 );
or \U$42452 ( \42829 , \42826 , \42828 );
or \U$42453 ( \42830 , \42827 , \42792 );
nand \U$42454 ( \42831 , \42829 , \42830 );
and \U$42455 ( \42832 , \42825 , \42831 );
and \U$42456 ( \42833 , \42822 , \42824 );
nor \U$42457 ( \42834 , \42832 , \42833 );
xor \U$42458 ( \42835 , \42520 , \42550 );
xor \U$42459 ( \42836 , \42835 , \42576 );
xor \U$42460 ( \42837 , \42682 , \42707 );
xor \U$42461 ( \42838 , \42837 , \42735 );
and \U$42462 ( \42839 , \42836 , \42838 );
xor \U$42463 ( \42840 , \42272 , \42279 );
xor \U$42464 ( \42841 , \42840 , \42288 );
xor \U$42465 ( \42842 , \42470 , \42475 );
xor \U$42466 ( \42843 , \42841 , \42842 );
xor \U$42467 ( \42844 , \42682 , \42707 );
xor \U$42468 ( \42845 , \42844 , \42735 );
and \U$42469 ( \42846 , \42843 , \42845 );
and \U$42470 ( \42847 , \42836 , \42843 );
or \U$42471 ( \42848 , \42839 , \42846 , \42847 );
xor \U$42472 ( \42849 , \42163 , \42181 );
xor \U$42473 ( \42850 , \42849 , \42207 );
xor \U$42474 ( \42851 , \42848 , \42850 );
xor \U$42475 ( \42852 , \42778 , \42780 );
xor \U$42476 ( \42853 , \42852 , \42783 );
and \U$42477 ( \42854 , \42851 , \42853 );
and \U$42478 ( \42855 , \42848 , \42850 );
or \U$42479 ( \42856 , \42854 , \42855 );
xor \U$42480 ( \42857 , \42501 , \42508 );
xor \U$42481 ( \42858 , \42857 , \42517 );
xor \U$42482 ( \42859 , \42558 , \42565 );
xor \U$42483 ( \42860 , \42859 , \42573 );
xor \U$42484 ( \42861 , \42858 , \42860 );
xor \U$42485 ( \42862 , \42689 , \42696 );
xor \U$42486 ( \42863 , \42862 , \42704 );
and \U$42487 ( \42864 , \42861 , \42863 );
and \U$42488 ( \42865 , \42858 , \42860 );
or \U$42489 ( \42866 , \42864 , \42865 );
nand \U$42490 ( \42867 , RIae76dc0_62, RIae78b48_125);
not \U$42491 ( \42868 , \42536 );
not \U$42492 ( \42869 , \42548 );
or \U$42493 ( \42870 , \42868 , \42869 );
or \U$42494 ( \42871 , \42536 , \42548 );
nand \U$42495 ( \42872 , \42870 , \42871 );
not \U$42496 ( \42873 , \42872 );
not \U$42497 ( \42874 , \42528 );
and \U$42498 ( \42875 , \42873 , \42874 );
and \U$42499 ( \42876 , \42872 , \42528 );
nor \U$42500 ( \42877 , \42875 , \42876 );
nand \U$42501 ( \42878 , \42867 , \42877 );
xor \U$42502 ( \42879 , \42866 , \42878 );
xor \U$42503 ( \42880 , \42715 , \42723 );
xor \U$42504 ( \42881 , \42880 , \42732 );
xor \U$42505 ( \42882 , \42635 , \42642 );
xor \U$42506 ( \42883 , \42882 , \42650 );
and \U$42507 ( \42884 , \42881 , \42883 );
xor \U$42508 ( \42885 , \42664 , \42671 );
xor \U$42509 ( \42886 , \42885 , \42679 );
xor \U$42510 ( \42887 , \42635 , \42642 );
xor \U$42511 ( \42888 , \42887 , \42650 );
and \U$42512 ( \42889 , \42886 , \42888 );
and \U$42513 ( \42890 , \42881 , \42886 );
or \U$42514 ( \42891 , \42884 , \42889 , \42890 );
and \U$42515 ( \42892 , \42879 , \42891 );
and \U$42516 ( \42893 , \42866 , \42878 );
or \U$42517 ( \42894 , \42892 , \42893 );
and \U$42518 ( \42895 , \5896 , RIae75380_6);
and \U$42519 ( \42896 , RIae75470_8, \5894 );
nor \U$42520 ( \42897 , \42895 , \42896 );
and \U$42521 ( \42898 , \42897 , \5590 );
not \U$42522 ( \42899 , \42897 );
and \U$42523 ( \42900 , \42899 , \5589 );
nor \U$42524 ( \42901 , \42898 , \42900 );
and \U$42525 ( \42902 , \4688 , RIae75830_16);
and \U$42526 ( \42903 , RIae75740_14, \4686 );
nor \U$42527 ( \42904 , \42902 , \42903 );
and \U$42528 ( \42905 , \42904 , \4481 );
not \U$42529 ( \42906 , \42904 );
and \U$42530 ( \42907 , \42906 , \4482 );
nor \U$42531 ( \42908 , \42905 , \42907 );
xor \U$42532 ( \42909 , \42901 , \42908 );
and \U$42533 ( \42910 , \5399 , RIae75290_4);
and \U$42534 ( \42911 , RIae751a0_2, \5397 );
nor \U$42535 ( \42912 , \42910 , \42911 );
and \U$42536 ( \42913 , \42912 , \5016 );
not \U$42537 ( \42914 , \42912 );
and \U$42538 ( \42915 , \42914 , \5403 );
nor \U$42539 ( \42916 , \42913 , \42915 );
and \U$42540 ( \42917 , \42909 , \42916 );
and \U$42541 ( \42918 , \42901 , \42908 );
or \U$42542 ( \42919 , \42917 , \42918 );
not \U$42543 ( \42920 , \3089 );
and \U$42544 ( \42921 , \2783 , RIae75a10_20);
and \U$42545 ( \42922 , RIae75920_18, \2781 );
nor \U$42546 ( \42923 , \42921 , \42922 );
not \U$42547 ( \42924 , \42923 );
or \U$42548 ( \42925 , \42920 , \42924 );
or \U$42549 ( \42926 , \42923 , \2789 );
nand \U$42550 ( \42927 , \42925 , \42926 );
and \U$42551 ( \42928 , \2224 , RIae78800_118);
and \U$42552 ( \42929 , RIae78710_116, \2222 );
nor \U$42553 ( \42930 , \42928 , \42929 );
and \U$42554 ( \42931 , \42930 , \2061 );
not \U$42555 ( \42932 , \42930 );
and \U$42556 ( \42933 , \42932 , \2060 );
nor \U$42557 ( \42934 , \42931 , \42933 );
xor \U$42558 ( \42935 , \42927 , \42934 );
and \U$42559 ( \42936 , \2607 , RIae75bf0_24);
and \U$42560 ( \42937 , RIae75b00_22, \2605 );
nor \U$42561 ( \42938 , \42936 , \42937 );
and \U$42562 ( \42939 , \42938 , \2611 );
not \U$42563 ( \42940 , \42938 );
and \U$42564 ( \42941 , \42940 , \2397 );
nor \U$42565 ( \42942 , \42939 , \42941 );
and \U$42566 ( \42943 , \42935 , \42942 );
and \U$42567 ( \42944 , \42927 , \42934 );
or \U$42568 ( \42945 , \42943 , \42944 );
xor \U$42569 ( \42946 , \42919 , \42945 );
and \U$42570 ( \42947 , \3730 , RIae75ce0_26);
and \U$42571 ( \42948 , RIae75dd0_28, \3728 );
nor \U$42572 ( \42949 , \42947 , \42948 );
and \U$42573 ( \42950 , \42949 , \3732 );
not \U$42574 ( \42951 , \42949 );
and \U$42575 ( \42952 , \42951 , \3422 );
nor \U$42576 ( \42953 , \42950 , \42952 );
not \U$42577 ( \42954 , \3218 );
and \U$42578 ( \42955 , \3214 , RIae75fb0_32);
and \U$42579 ( \42956 , RIae75ec0_30, \3212 );
nor \U$42580 ( \42957 , \42955 , \42956 );
not \U$42581 ( \42958 , \42957 );
or \U$42582 ( \42959 , \42954 , \42958 );
or \U$42583 ( \42960 , \42957 , \3218 );
nand \U$42584 ( \42961 , \42959 , \42960 );
xor \U$42585 ( \42962 , \42953 , \42961 );
and \U$42586 ( \42963 , \4247 , RIae75650_12);
and \U$42587 ( \42964 , RIae75560_10, \4245 );
nor \U$42588 ( \42965 , \42963 , \42964 );
and \U$42589 ( \42966 , \42965 , \3989 );
not \U$42590 ( \42967 , \42965 );
and \U$42591 ( \42968 , \42967 , \4251 );
nor \U$42592 ( \42969 , \42966 , \42968 );
and \U$42593 ( \42970 , \42962 , \42969 );
and \U$42594 ( \42971 , \42953 , \42961 );
or \U$42595 ( \42972 , \42970 , \42971 );
and \U$42596 ( \42973 , \42946 , \42972 );
and \U$42597 ( \42974 , \42919 , \42945 );
or \U$42598 ( \42975 , \42973 , \42974 );
and \U$42599 ( \42976 , \1138 , RIae78440_110);
and \U$42600 ( \42977 , RIae784b8_111, \1136 );
nor \U$42601 ( \42978 , \42976 , \42977 );
and \U$42602 ( \42979 , \42978 , \1012 );
not \U$42603 ( \42980 , \42978 );
and \U$42604 ( \42981 , \42980 , \1142 );
nor \U$42605 ( \42982 , \42979 , \42981 );
and \U$42606 ( \42983 , \672 , RIae77f90_100);
and \U$42607 ( \42984 , RIae78080_102, \670 );
nor \U$42608 ( \42985 , \42983 , \42984 );
and \U$42609 ( \42986 , \42985 , \588 );
not \U$42610 ( \42987 , \42985 );
and \U$42611 ( \42988 , \42987 , \587 );
nor \U$42612 ( \42989 , \42986 , \42988 );
xor \U$42613 ( \42990 , \42982 , \42989 );
not \U$42614 ( \42991 , \787 );
and \U$42615 ( \42992 , \883 , RIae78260_106);
and \U$42616 ( \42993 , RIae78620_114, \881 );
nor \U$42617 ( \42994 , \42992 , \42993 );
not \U$42618 ( \42995 , \42994 );
or \U$42619 ( \42996 , \42991 , \42995 );
or \U$42620 ( \42997 , \42994 , \787 );
nand \U$42621 ( \42998 , \42996 , \42997 );
and \U$42622 ( \42999 , \42990 , \42998 );
and \U$42623 ( \43000 , \42982 , \42989 );
or \U$42624 ( \43001 , \42999 , \43000 );
and \U$42625 ( \43002 , \558 , RIae78350_108);
and \U$42626 ( \43003 , RIae78170_104, \556 );
nor \U$42627 ( \43004 , \43002 , \43003 );
and \U$42628 ( \43005 , \43004 , \504 );
not \U$42629 ( \43006 , \43004 );
and \U$42630 ( \43007 , \43006 , \562 );
nor \U$42631 ( \43008 , \43005 , \43007 );
not \U$42632 ( \43009 , \400 );
and \U$42633 ( \43010 , \436 , RIae77108_69);
and \U$42634 ( \43011 , RIae77090_68, \434 );
nor \U$42635 ( \43012 , \43010 , \43011 );
not \U$42636 ( \43013 , \43012 );
or \U$42637 ( \43014 , \43009 , \43013 );
or \U$42638 ( \43015 , \43012 , \400 );
nand \U$42639 ( \43016 , \43014 , \43015 );
xor \U$42640 ( \43017 , \43008 , \43016 );
not \U$42641 ( \43018 , \469 );
and \U$42642 ( \43019 , \514 , RIae77270_72);
and \U$42643 ( \43020 , RIae77360_74, \512 );
nor \U$42644 ( \43021 , \43019 , \43020 );
not \U$42645 ( \43022 , \43021 );
or \U$42646 ( \43023 , \43018 , \43022 );
or \U$42647 ( \43024 , \43021 , \471 );
nand \U$42648 ( \43025 , \43023 , \43024 );
and \U$42649 ( \43026 , \43017 , \43025 );
and \U$42650 ( \43027 , \43008 , \43016 );
or \U$42651 ( \43028 , \43026 , \43027 );
xor \U$42652 ( \43029 , \43001 , \43028 );
and \U$42653 ( \43030 , \1939 , RIae789e0_122);
and \U$42654 ( \43031 , RIae788f0_120, \1937 );
nor \U$42655 ( \43032 , \43030 , \43031 );
and \U$42656 ( \43033 , \43032 , \1735 );
not \U$42657 ( \43034 , \43032 );
and \U$42658 ( \43035 , \43034 , \1734 );
nor \U$42659 ( \43036 , \43033 , \43035 );
and \U$42660 ( \43037 , \1376 , RIae77cc0_94);
and \U$42661 ( \43038 , RIae77bd0_92, \1374 );
nor \U$42662 ( \43039 , \43037 , \43038 );
and \U$42663 ( \43040 , \43039 , \1380 );
not \U$42664 ( \43041 , \43039 );
and \U$42665 ( \43042 , \43041 , \1261 );
nor \U$42666 ( \43043 , \43040 , \43042 );
xor \U$42667 ( \43044 , \43036 , \43043 );
and \U$42668 ( \43045 , \1593 , RIae77db0_96);
and \U$42669 ( \43046 , RIae77ea0_98, \1591 );
nor \U$42670 ( \43047 , \43045 , \43046 );
and \U$42671 ( \43048 , \43047 , \1498 );
not \U$42672 ( \43049 , \43047 );
and \U$42673 ( \43050 , \43049 , \1488 );
nor \U$42674 ( \43051 , \43048 , \43050 );
and \U$42675 ( \43052 , \43044 , \43051 );
and \U$42676 ( \43053 , \43036 , \43043 );
or \U$42677 ( \43054 , \43052 , \43053 );
and \U$42678 ( \43055 , \43029 , \43054 );
and \U$42679 ( \43056 , \43001 , \43028 );
or \U$42680 ( \43057 , \43055 , \43056 );
xor \U$42681 ( \43058 , \42975 , \43057 );
and \U$42682 ( \43059 , \7633 , RIae76190_36);
and \U$42683 ( \43060 , RIae760a0_34, \7631 );
nor \U$42684 ( \43061 , \43059 , \43060 );
and \U$42685 ( \43062 , \43061 , \7206 );
not \U$42686 ( \43063 , \43061 );
and \U$42687 ( \43064 , \43063 , \7205 );
nor \U$42688 ( \43065 , \43062 , \43064 );
and \U$42689 ( \43066 , \6172 , RIae76460_42);
and \U$42690 ( \43067 , RIae76550_44, \6170 );
nor \U$42691 ( \43068 , \43066 , \43067 );
and \U$42692 ( \43069 , \43068 , \6176 );
not \U$42693 ( \43070 , \43068 );
and \U$42694 ( \43071 , \43070 , \6175 );
nor \U$42695 ( \43072 , \43069 , \43071 );
xor \U$42696 ( \43073 , \43065 , \43072 );
and \U$42697 ( \43074 , \6941 , RIae76730_48);
and \U$42698 ( \43075 , RIae76640_46, \6939 );
nor \U$42699 ( \43076 , \43074 , \43075 );
and \U$42700 ( \43077 , \43076 , \6314 );
not \U$42701 ( \43078 , \43076 );
and \U$42702 ( \43079 , \43078 , \6945 );
nor \U$42703 ( \43080 , \43077 , \43079 );
and \U$42704 ( \43081 , \43073 , \43080 );
and \U$42705 ( \43082 , \43065 , \43072 );
or \U$42706 ( \43083 , \43081 , \43082 );
and \U$42707 ( \43084 , \10548 , RIae76be0_58);
and \U$42708 ( \43085 , RIae78ad0_124, \10546 );
nor \U$42709 ( \43086 , \43084 , \43085 );
and \U$42710 ( \43087 , \43086 , \10421 );
not \U$42711 ( \43088 , \43086 );
and \U$42712 ( \43089 , \43088 , \10118 );
nor \U$42713 ( \43090 , \43087 , \43089 );
xor \U$42714 ( \43091 , \43090 , \12184 );
and \U$42715 ( \43092 , \11470 , RIae78d28_129);
and \U$42716 ( \43093 , RIae78e18_131, \11468 );
nor \U$42717 ( \43094 , \43092 , \43093 );
and \U$42718 ( \43095 , \43094 , \10936 );
not \U$42719 ( \43096 , \43094 );
and \U$42720 ( \43097 , \43096 , \11474 );
nor \U$42721 ( \43098 , \43095 , \43097 );
and \U$42722 ( \43099 , \43091 , \43098 );
and \U$42723 ( \43100 , \43090 , \12184 );
or \U$42724 ( \43101 , \43099 , \43100 );
xor \U$42725 ( \43102 , \43083 , \43101 );
and \U$42726 ( \43103 , \8371 , RIae76370_40);
and \U$42727 ( \43104 , RIae76280_38, \8369 );
nor \U$42728 ( \43105 , \43103 , \43104 );
and \U$42729 ( \43106 , \43105 , \8020 );
not \U$42730 ( \43107 , \43105 );
and \U$42731 ( \43108 , \43107 , \8019 );
nor \U$42732 ( \43109 , \43106 , \43108 );
and \U$42733 ( \43110 , \8966 , RIae76af0_56);
and \U$42734 ( \43111 , RIae76a00_54, \8964 );
nor \U$42735 ( \43112 , \43110 , \43111 );
and \U$42736 ( \43113 , \43112 , \8799 );
not \U$42737 ( \43114 , \43112 );
and \U$42738 ( \43115 , \43114 , \8789 );
nor \U$42739 ( \43116 , \43113 , \43115 );
xor \U$42740 ( \43117 , \43109 , \43116 );
and \U$42741 ( \43118 , \9760 , RIae76820_50);
and \U$42742 ( \43119 , RIae76910_52, \9758 );
nor \U$42743 ( \43120 , \43118 , \43119 );
and \U$42744 ( \43121 , \43120 , \9273 );
not \U$42745 ( \43122 , \43120 );
and \U$42746 ( \43123 , \43122 , \9272 );
nor \U$42747 ( \43124 , \43121 , \43123 );
and \U$42748 ( \43125 , \43117 , \43124 );
and \U$42749 ( \43126 , \43109 , \43116 );
or \U$42750 ( \43127 , \43125 , \43126 );
and \U$42751 ( \43128 , \43102 , \43127 );
and \U$42752 ( \43129 , \43083 , \43101 );
or \U$42753 ( \43130 , \43128 , \43129 );
and \U$42754 ( \43131 , \43058 , \43130 );
and \U$42755 ( \43132 , \42975 , \43057 );
or \U$42756 ( \43133 , \43131 , \43132 );
xor \U$42757 ( \43134 , \42894 , \43133 );
xor \U$42758 ( \43135 , \42170 , \10936 );
xor \U$42759 ( \43136 , \43135 , \42178 );
xor \U$42760 ( \43137 , \42483 , \42485 );
xor \U$42761 ( \43138 , \43137 , \42488 );
and \U$42762 ( \43139 , \43136 , \43138 );
xor \U$42763 ( \43140 , \42189 , \42196 );
xor \U$42764 ( \43141 , \43140 , \42204 );
xor \U$42765 ( \43142 , \42458 , \42463 );
xor \U$42766 ( \43143 , \43141 , \43142 );
xor \U$42767 ( \43144 , \42483 , \42485 );
xor \U$42768 ( \43145 , \43144 , \42488 );
and \U$42769 ( \43146 , \43143 , \43145 );
and \U$42770 ( \43147 , \43136 , \43143 );
or \U$42771 ( \43148 , \43139 , \43146 , \43147 );
and \U$42772 ( \43149 , \43134 , \43148 );
and \U$42773 ( \43150 , \42894 , \43133 );
or \U$42774 ( \43151 , \43149 , \43150 );
xor \U$42775 ( \43152 , \42856 , \43151 );
xor \U$42776 ( \43153 , \42579 , \42656 );
xor \U$42777 ( \43154 , \43153 , \42738 );
xor \U$42778 ( \43155 , \42468 , \42480 );
xor \U$42779 ( \43156 , \43155 , \42491 );
and \U$42780 ( \43157 , \43154 , \43156 );
xor \U$42781 ( \43158 , \42321 , \42323 );
xor \U$42782 ( \43159 , \43158 , \42326 );
xor \U$42783 ( \43160 , \42748 , \42755 );
xor \U$42784 ( \43161 , \43159 , \43160 );
xor \U$42785 ( \43162 , \42468 , \42480 );
xor \U$42786 ( \43163 , \43162 , \42491 );
and \U$42787 ( \43164 , \43161 , \43163 );
and \U$42788 ( \43165 , \43154 , \43161 );
or \U$42789 ( \43166 , \43157 , \43164 , \43165 );
and \U$42790 ( \43167 , \43152 , \43166 );
and \U$42791 ( \43168 , \42856 , \43151 );
nor \U$42792 ( \43169 , \43167 , \43168 );
xor \U$42793 ( \43170 , \42834 , \43169 );
xor \U$42794 ( \43171 , \42445 , \42450 );
xor \U$42795 ( \43172 , \43171 , \42453 );
and \U$42796 ( \43173 , \43170 , \43172 );
and \U$42797 ( \43174 , \42834 , \43169 );
or \U$42798 ( \43175 , \43173 , \43174 );
not \U$42799 ( \43176 , \42038 );
not \U$42800 ( \43177 , \42358 );
and \U$42801 ( \43178 , \43176 , \43177 );
and \U$42802 ( \43179 , \42038 , \42358 );
nor \U$42803 ( \43180 , \43178 , \43179 );
not \U$42804 ( \43181 , \43180 );
not \U$42805 ( \43182 , \42052 );
and \U$42806 ( \43183 , \43181 , \43182 );
and \U$42807 ( \43184 , \43180 , \42052 );
nor \U$42808 ( \43185 , \43183 , \43184 );
xor \U$42809 ( \43186 , \43175 , \43185 );
xor \U$42810 ( \43187 , \42456 , \42797 );
xor \U$42811 ( \43188 , \43187 , \42804 );
and \U$42812 ( \43189 , \43186 , \43188 );
and \U$42813 ( \43190 , \43175 , \43185 );
or \U$42814 ( \43191 , \43189 , \43190 );
not \U$42815 ( \43192 , \43191 );
not \U$42816 ( \43193 , \42437 );
not \U$42817 ( \43194 , \42807 );
not \U$42818 ( \43195 , \42439 );
and \U$42819 ( \43196 , \43194 , \43195 );
and \U$42820 ( \43197 , \42807 , \42439 );
nor \U$42821 ( \43198 , \43196 , \43197 );
not \U$42822 ( \43199 , \43198 );
or \U$42823 ( \43200 , \43193 , \43199 );
or \U$42824 ( \43201 , \43198 , \42437 );
nand \U$42825 ( \43202 , \43200 , \43201 );
nand \U$42826 ( \43203 , \43192 , \43202 );
or \U$42827 ( \43204 , \42817 , \43203 );
xnor \U$42828 ( \43205 , \43203 , \42817 );
not \U$42829 ( \43206 , \43202 );
not \U$42830 ( \43207 , \43191 );
or \U$42831 ( \43208 , \43206 , \43207 );
or \U$42832 ( \43209 , \43202 , \43191 );
nand \U$42833 ( \43210 , \43208 , \43209 );
xor \U$42834 ( \43211 , \42834 , \43169 );
xor \U$42835 ( \43212 , \43211 , \43172 );
xor \U$42836 ( \43213 , \42763 , \42769 );
xor \U$42837 ( \43214 , \43213 , \42794 );
or \U$42838 ( \43215 , \43212 , \43214 );
not \U$42839 ( \43216 , \43214 );
not \U$42840 ( \43217 , \43212 );
or \U$42841 ( \43218 , \43216 , \43217 );
xor \U$42842 ( \43219 , \43083 , \43101 );
xor \U$42843 ( \43220 , \43219 , \43127 );
xor \U$42844 ( \43221 , \43001 , \43028 );
xor \U$42845 ( \43222 , \43221 , \43054 );
xor \U$42846 ( \43223 , \43220 , \43222 );
xor \U$42847 ( \43224 , \42919 , \42945 );
xor \U$42848 ( \43225 , \43224 , \42972 );
and \U$42849 ( \43226 , \43223 , \43225 );
and \U$42850 ( \43227 , \43220 , \43222 );
or \U$42851 ( \43228 , \43226 , \43227 );
xor \U$42852 ( \43229 , \42604 , \42627 );
xor \U$42853 ( \43230 , \43229 , \42653 );
xor \U$42854 ( \43231 , \43228 , \43230 );
or \U$42855 ( \43232 , \42877 , \42867 );
nand \U$42856 ( \43233 , \43232 , \42878 );
xor \U$42857 ( \43234 , \42858 , \42860 );
xor \U$42858 ( \43235 , \43234 , \42863 );
and \U$42859 ( \43236 , \43233 , \43235 );
xor \U$42860 ( \43237 , \42635 , \42642 );
xor \U$42861 ( \43238 , \43237 , \42650 );
xor \U$42862 ( \43239 , \42881 , \42886 );
xor \U$42863 ( \43240 , \43238 , \43239 );
xor \U$42864 ( \43241 , \42858 , \42860 );
xor \U$42865 ( \43242 , \43241 , \42863 );
and \U$42866 ( \43243 , \43240 , \43242 );
and \U$42867 ( \43244 , \43233 , \43240 );
or \U$42868 ( \43245 , \43236 , \43243 , \43244 );
and \U$42869 ( \43246 , \43231 , \43245 );
and \U$42870 ( \43247 , \43228 , \43230 );
or \U$42871 ( \43248 , \43246 , \43247 );
and \U$42872 ( \43249 , \4247 , RIae75dd0_28);
and \U$42873 ( \43250 , RIae75650_12, \4245 );
nor \U$42874 ( \43251 , \43249 , \43250 );
and \U$42875 ( \43252 , \43251 , \3989 );
not \U$42876 ( \43253 , \43251 );
and \U$42877 ( \43254 , \43253 , \4251 );
nor \U$42878 ( \43255 , \43252 , \43254 );
not \U$42879 ( \43256 , \3218 );
and \U$42880 ( \43257 , \3214 , RIae75920_18);
and \U$42881 ( \43258 , RIae75fb0_32, \3212 );
nor \U$42882 ( \43259 , \43257 , \43258 );
not \U$42883 ( \43260 , \43259 );
or \U$42884 ( \43261 , \43256 , \43260 );
or \U$42885 ( \43262 , \43259 , \2774 );
nand \U$42886 ( \43263 , \43261 , \43262 );
xor \U$42887 ( \43264 , \43255 , \43263 );
and \U$42888 ( \43265 , \3730 , RIae75ec0_30);
and \U$42889 ( \43266 , RIae75ce0_26, \3728 );
nor \U$42890 ( \43267 , \43265 , \43266 );
and \U$42891 ( \43268 , \43267 , \3732 );
not \U$42892 ( \43269 , \43267 );
and \U$42893 ( \43270 , \43269 , \3422 );
nor \U$42894 ( \43271 , \43268 , \43270 );
and \U$42895 ( \43272 , \43264 , \43271 );
and \U$42896 ( \43273 , \43255 , \43263 );
or \U$42897 ( \43274 , \43272 , \43273 );
and \U$42898 ( \43275 , \2607 , RIae78710_116);
and \U$42899 ( \43276 , RIae75bf0_24, \2605 );
nor \U$42900 ( \43277 , \43275 , \43276 );
and \U$42901 ( \43278 , \43277 , \2611 );
not \U$42902 ( \43279 , \43277 );
and \U$42903 ( \43280 , \43279 , \2397 );
nor \U$42904 ( \43281 , \43278 , \43280 );
and \U$42905 ( \43282 , \2224 , RIae788f0_120);
and \U$42906 ( \43283 , RIae78800_118, \2222 );
nor \U$42907 ( \43284 , \43282 , \43283 );
and \U$42908 ( \43285 , \43284 , \2061 );
not \U$42909 ( \43286 , \43284 );
and \U$42910 ( \43287 , \43286 , \2060 );
nor \U$42911 ( \43288 , \43285 , \43287 );
xor \U$42912 ( \43289 , \43281 , \43288 );
not \U$42913 ( \43290 , \3089 );
and \U$42914 ( \43291 , \2783 , RIae75b00_22);
and \U$42915 ( \43292 , RIae75a10_20, \2781 );
nor \U$42916 ( \43293 , \43291 , \43292 );
not \U$42917 ( \43294 , \43293 );
or \U$42918 ( \43295 , \43290 , \43294 );
or \U$42919 ( \43296 , \43293 , \2789 );
nand \U$42920 ( \43297 , \43295 , \43296 );
and \U$42921 ( \43298 , \43289 , \43297 );
and \U$42922 ( \43299 , \43281 , \43288 );
or \U$42923 ( \43300 , \43298 , \43299 );
xor \U$42924 ( \43301 , \43274 , \43300 );
and \U$42925 ( \43302 , \5399 , RIae75740_14);
and \U$42926 ( \43303 , RIae75290_4, \5397 );
nor \U$42927 ( \43304 , \43302 , \43303 );
and \U$42928 ( \43305 , \43304 , \5016 );
not \U$42929 ( \43306 , \43304 );
and \U$42930 ( \43307 , \43306 , \5403 );
nor \U$42931 ( \43308 , \43305 , \43307 );
and \U$42932 ( \43309 , \4688 , RIae75560_10);
and \U$42933 ( \43310 , RIae75830_16, \4686 );
nor \U$42934 ( \43311 , \43309 , \43310 );
and \U$42935 ( \43312 , \43311 , \4481 );
not \U$42936 ( \43313 , \43311 );
and \U$42937 ( \43314 , \43313 , \4482 );
nor \U$42938 ( \43315 , \43312 , \43314 );
xor \U$42939 ( \43316 , \43308 , \43315 );
and \U$42940 ( \43317 , \5896 , RIae751a0_2);
and \U$42941 ( \43318 , RIae75380_6, \5894 );
nor \U$42942 ( \43319 , \43317 , \43318 );
and \U$42943 ( \43320 , \43319 , \5590 );
not \U$42944 ( \43321 , \43319 );
and \U$42945 ( \43322 , \43321 , \5589 );
nor \U$42946 ( \43323 , \43320 , \43322 );
and \U$42947 ( \43324 , \43316 , \43323 );
and \U$42948 ( \43325 , \43308 , \43315 );
or \U$42949 ( \43326 , \43324 , \43325 );
and \U$42950 ( \43327 , \43301 , \43326 );
and \U$42951 ( \43328 , \43274 , \43300 );
or \U$42952 ( \43329 , \43327 , \43328 );
and \U$42953 ( \43330 , \1376 , RIae784b8_111);
and \U$42954 ( \43331 , RIae77cc0_94, \1374 );
nor \U$42955 ( \43332 , \43330 , \43331 );
and \U$42956 ( \43333 , \43332 , \1380 );
not \U$42957 ( \43334 , \43332 );
and \U$42958 ( \43335 , \43334 , \1261 );
nor \U$42959 ( \43336 , \43333 , \43335 );
and \U$42960 ( \43337 , \1593 , RIae77bd0_92);
and \U$42961 ( \43338 , RIae77db0_96, \1591 );
nor \U$42962 ( \43339 , \43337 , \43338 );
and \U$42963 ( \43340 , \43339 , \1498 );
not \U$42964 ( \43341 , \43339 );
and \U$42965 ( \43342 , \43341 , \1488 );
nor \U$42966 ( \43343 , \43340 , \43342 );
xor \U$42967 ( \43344 , \43336 , \43343 );
and \U$42968 ( \43345 , \1939 , RIae77ea0_98);
and \U$42969 ( \43346 , RIae789e0_122, \1937 );
nor \U$42970 ( \43347 , \43345 , \43346 );
and \U$42971 ( \43348 , \43347 , \1735 );
not \U$42972 ( \43349 , \43347 );
and \U$42973 ( \43350 , \43349 , \1734 );
nor \U$42974 ( \43351 , \43348 , \43350 );
and \U$42975 ( \43352 , \43344 , \43351 );
and \U$42976 ( \43353 , \43336 , \43343 );
or \U$42977 ( \43354 , \43352 , \43353 );
and \U$42978 ( \43355 , \672 , RIae78170_104);
and \U$42979 ( \43356 , RIae77f90_100, \670 );
nor \U$42980 ( \43357 , \43355 , \43356 );
and \U$42981 ( \43358 , \43357 , \588 );
not \U$42982 ( \43359 , \43357 );
and \U$42983 ( \43360 , \43359 , \587 );
nor \U$42984 ( \43361 , \43358 , \43360 );
not \U$42985 ( \43362 , \787 );
and \U$42986 ( \43363 , \883 , RIae78080_102);
and \U$42987 ( \43364 , RIae78260_106, \881 );
nor \U$42988 ( \43365 , \43363 , \43364 );
not \U$42989 ( \43366 , \43365 );
or \U$42990 ( \43367 , \43362 , \43366 );
or \U$42991 ( \43368 , \43365 , \787 );
nand \U$42992 ( \43369 , \43367 , \43368 );
xor \U$42993 ( \43370 , \43361 , \43369 );
and \U$42994 ( \43371 , \1138 , RIae78620_114);
and \U$42995 ( \43372 , RIae78440_110, \1136 );
nor \U$42996 ( \43373 , \43371 , \43372 );
and \U$42997 ( \43374 , \43373 , \1012 );
not \U$42998 ( \43375 , \43373 );
and \U$42999 ( \43376 , \43375 , \1142 );
nor \U$43000 ( \43377 , \43374 , \43376 );
and \U$43001 ( \43378 , \43370 , \43377 );
and \U$43002 ( \43379 , \43361 , \43369 );
or \U$43003 ( \43380 , \43378 , \43379 );
xor \U$43004 ( \43381 , \43354 , \43380 );
not \U$43005 ( \43382 , \400 );
and \U$43006 ( \43383 , \436 , RIae76cd0_60);
and \U$43007 ( \43384 , RIae77108_69, \434 );
nor \U$43008 ( \43385 , \43383 , \43384 );
not \U$43009 ( \43386 , \43385 );
or \U$43010 ( \43387 , \43382 , \43386 );
or \U$43011 ( \43388 , \43385 , \400 );
nand \U$43012 ( \43389 , \43387 , \43388 );
not \U$43013 ( \43390 , \469 );
and \U$43014 ( \43391 , \514 , RIae77090_68);
and \U$43015 ( \43392 , RIae77270_72, \512 );
nor \U$43016 ( \43393 , \43391 , \43392 );
not \U$43017 ( \43394 , \43393 );
or \U$43018 ( \43395 , \43390 , \43394 );
or \U$43019 ( \43396 , \43393 , \471 );
nand \U$43020 ( \43397 , \43395 , \43396 );
xor \U$43021 ( \43398 , \43389 , \43397 );
and \U$43022 ( \43399 , \558 , RIae77360_74);
and \U$43023 ( \43400 , RIae78350_108, \556 );
nor \U$43024 ( \43401 , \43399 , \43400 );
and \U$43025 ( \43402 , \43401 , \504 );
not \U$43026 ( \43403 , \43401 );
and \U$43027 ( \43404 , \43403 , \562 );
nor \U$43028 ( \43405 , \43402 , \43404 );
and \U$43029 ( \43406 , \43398 , \43405 );
and \U$43030 ( \43407 , \43389 , \43397 );
or \U$43031 ( \43408 , \43406 , \43407 );
and \U$43032 ( \43409 , \43381 , \43408 );
and \U$43033 ( \43410 , \43354 , \43380 );
or \U$43034 ( \43411 , \43409 , \43410 );
xor \U$43035 ( \43412 , \43329 , \43411 );
and \U$43036 ( \43413 , \6941 , RIae76550_44);
and \U$43037 ( \43414 , RIae76730_48, \6939 );
nor \U$43038 ( \43415 , \43413 , \43414 );
and \U$43039 ( \43416 , \43415 , \6314 );
not \U$43040 ( \43417 , \43415 );
and \U$43041 ( \43418 , \43417 , \6945 );
nor \U$43042 ( \43419 , \43416 , \43418 );
and \U$43043 ( \43420 , \6172 , RIae75470_8);
and \U$43044 ( \43421 , RIae76460_42, \6170 );
nor \U$43045 ( \43422 , \43420 , \43421 );
and \U$43046 ( \43423 , \43422 , \6176 );
not \U$43047 ( \43424 , \43422 );
and \U$43048 ( \43425 , \43424 , \6175 );
nor \U$43049 ( \43426 , \43423 , \43425 );
xor \U$43050 ( \43427 , \43419 , \43426 );
and \U$43051 ( \43428 , \7633 , RIae76640_46);
and \U$43052 ( \43429 , RIae76190_36, \7631 );
nor \U$43053 ( \43430 , \43428 , \43429 );
and \U$43054 ( \43431 , \43430 , \7206 );
not \U$43055 ( \43432 , \43430 );
and \U$43056 ( \43433 , \43432 , \7205 );
nor \U$43057 ( \43434 , \43431 , \43433 );
and \U$43058 ( \43435 , \43427 , \43434 );
and \U$43059 ( \43436 , \43419 , \43426 );
or \U$43060 ( \43437 , \43435 , \43436 );
and \U$43061 ( \43438 , \10548 , RIae76910_52);
and \U$43062 ( \43439 , RIae76be0_58, \10546 );
nor \U$43063 ( \43440 , \43438 , \43439 );
and \U$43064 ( \43441 , \43440 , \10421 );
not \U$43065 ( \43442 , \43440 );
and \U$43066 ( \43443 , \43442 , \10118 );
nor \U$43067 ( \43444 , \43441 , \43443 );
nand \U$43068 ( \43445 , RIae78e18_131, \12180 );
and \U$43069 ( \43446 , \43445 , \12184 );
not \U$43070 ( \43447 , \43445 );
and \U$43071 ( \43448 , \43447 , \11827 );
nor \U$43072 ( \43449 , \43446 , \43448 );
xor \U$43073 ( \43450 , \43444 , \43449 );
and \U$43074 ( \43451 , \11470 , RIae78ad0_124);
and \U$43075 ( \43452 , RIae78d28_129, \11468 );
nor \U$43076 ( \43453 , \43451 , \43452 );
and \U$43077 ( \43454 , \43453 , \10936 );
not \U$43078 ( \43455 , \43453 );
and \U$43079 ( \43456 , \43455 , \11474 );
nor \U$43080 ( \43457 , \43454 , \43456 );
and \U$43081 ( \43458 , \43450 , \43457 );
and \U$43082 ( \43459 , \43444 , \43449 );
or \U$43083 ( \43460 , \43458 , \43459 );
xor \U$43084 ( \43461 , \43437 , \43460 );
and \U$43085 ( \43462 , \8371 , RIae760a0_34);
and \U$43086 ( \43463 , RIae76370_40, \8369 );
nor \U$43087 ( \43464 , \43462 , \43463 );
and \U$43088 ( \43465 , \43464 , \8020 );
not \U$43089 ( \43466 , \43464 );
and \U$43090 ( \43467 , \43466 , \8019 );
nor \U$43091 ( \43468 , \43465 , \43467 );
and \U$43092 ( \43469 , \8966 , RIae76280_38);
and \U$43093 ( \43470 , RIae76af0_56, \8964 );
nor \U$43094 ( \43471 , \43469 , \43470 );
and \U$43095 ( \43472 , \43471 , \8799 );
not \U$43096 ( \43473 , \43471 );
and \U$43097 ( \43474 , \43473 , \8789 );
nor \U$43098 ( \43475 , \43472 , \43474 );
xor \U$43099 ( \43476 , \43468 , \43475 );
and \U$43100 ( \43477 , \9760 , RIae76a00_54);
and \U$43101 ( \43478 , RIae76820_50, \9758 );
nor \U$43102 ( \43479 , \43477 , \43478 );
and \U$43103 ( \43480 , \43479 , \9273 );
not \U$43104 ( \43481 , \43479 );
and \U$43105 ( \43482 , \43481 , \9764 );
nor \U$43106 ( \43483 , \43480 , \43482 );
and \U$43107 ( \43484 , \43476 , \43483 );
and \U$43108 ( \43485 , \43468 , \43475 );
or \U$43109 ( \43486 , \43484 , \43485 );
and \U$43110 ( \43487 , \43461 , \43486 );
and \U$43111 ( \43488 , \43437 , \43460 );
or \U$43112 ( \43489 , \43487 , \43488 );
and \U$43113 ( \43490 , \43412 , \43489 );
and \U$43114 ( \43491 , \43329 , \43411 );
or \U$43115 ( \43492 , \43490 , \43491 );
xor \U$43116 ( \43493 , \42611 , \42616 );
xor \U$43117 ( \43494 , \43493 , \42624 );
xor \U$43118 ( \43495 , \42586 , \42593 );
xor \U$43119 ( \43496 , \43495 , \42601 );
and \U$43120 ( \43497 , \43494 , \43496 );
xor \U$43121 ( \43498 , \43090 , \12184 );
xor \U$43122 ( \43499 , \43498 , \43098 );
xor \U$43123 ( \43500 , \43065 , \43072 );
xor \U$43124 ( \43501 , \43500 , \43080 );
and \U$43125 ( \43502 , \43499 , \43501 );
xor \U$43126 ( \43503 , \43109 , \43116 );
xor \U$43127 ( \43504 , \43503 , \43124 );
xor \U$43128 ( \43505 , \43065 , \43072 );
xor \U$43129 ( \43506 , \43505 , \43080 );
and \U$43130 ( \43507 , \43504 , \43506 );
and \U$43131 ( \43508 , \43499 , \43504 );
or \U$43132 ( \43509 , \43502 , \43507 , \43508 );
xor \U$43133 ( \43510 , \42586 , \42593 );
xor \U$43134 ( \43511 , \43510 , \42601 );
and \U$43135 ( \43512 , \43509 , \43511 );
and \U$43136 ( \43513 , \43494 , \43509 );
or \U$43137 ( \43514 , \43497 , \43512 , \43513 );
xor \U$43138 ( \43515 , \43492 , \43514 );
xor \U$43139 ( \43516 , \42927 , \42934 );
xor \U$43140 ( \43517 , \43516 , \42942 );
xor \U$43141 ( \43518 , \42901 , \42908 );
xor \U$43142 ( \43519 , \43518 , \42916 );
and \U$43143 ( \43520 , \43517 , \43519 );
xor \U$43144 ( \43521 , \42953 , \42961 );
xor \U$43145 ( \43522 , \43521 , \42969 );
xor \U$43146 ( \43523 , \42901 , \42908 );
xor \U$43147 ( \43524 , \43523 , \42916 );
and \U$43148 ( \43525 , \43522 , \43524 );
and \U$43149 ( \43526 , \43517 , \43522 );
or \U$43150 ( \43527 , \43520 , \43525 , \43526 );
not \U$43151 ( \43528 , \388 );
and \U$43152 ( \43529 , \384 , RIae76dc0_62);
and \U$43153 ( \43530 , RIae76cd0_60, \382 );
nor \U$43154 ( \43531 , \43529 , \43530 );
not \U$43155 ( \43532 , \43531 );
or \U$43156 ( \43533 , \43528 , \43532 );
or \U$43157 ( \43534 , \43531 , \392 );
nand \U$43158 ( \43535 , \43533 , \43534 );
not \U$43159 ( \43536 , RIae76eb0_64);
nor \U$43160 ( \43537 , \43536 , \491 );
xor \U$43161 ( \43538 , \43535 , \43537 );
nand \U$43162 ( \43539 , RIae76fa0_66, RIae78b48_125);
and \U$43163 ( \43540 , \384 , RIae76eb0_64);
and \U$43164 ( \43541 , RIae76dc0_62, \382 );
nor \U$43165 ( \43542 , \43540 , \43541 );
not \U$43166 ( \43543 , \43542 );
not \U$43167 ( \43544 , \392 );
and \U$43168 ( \43545 , \43543 , \43544 );
and \U$43169 ( \43546 , \43542 , \388 );
nor \U$43170 ( \43547 , \43545 , \43546 );
nand \U$43171 ( \43548 , \43539 , \43547 );
and \U$43172 ( \43549 , \43538 , \43548 );
and \U$43173 ( \43550 , \43535 , \43537 );
or \U$43174 ( \43551 , \43549 , \43550 );
xor \U$43175 ( \43552 , \43527 , \43551 );
xor \U$43176 ( \43553 , \42982 , \42989 );
xor \U$43177 ( \43554 , \43553 , \42998 );
xor \U$43178 ( \43555 , \43008 , \43016 );
xor \U$43179 ( \43556 , \43555 , \43025 );
xor \U$43180 ( \43557 , \43554 , \43556 );
xor \U$43181 ( \43558 , \43036 , \43043 );
xor \U$43182 ( \43559 , \43558 , \43051 );
and \U$43183 ( \43560 , \43557 , \43559 );
and \U$43184 ( \43561 , \43554 , \43556 );
or \U$43185 ( \43562 , \43560 , \43561 );
and \U$43186 ( \43563 , \43552 , \43562 );
and \U$43187 ( \43564 , \43527 , \43551 );
or \U$43188 ( \43565 , \43563 , \43564 );
and \U$43189 ( \43566 , \43515 , \43565 );
and \U$43190 ( \43567 , \43492 , \43514 );
or \U$43191 ( \43568 , \43566 , \43567 );
xor \U$43192 ( \43569 , \43248 , \43568 );
xor \U$43193 ( \43570 , \42682 , \42707 );
xor \U$43194 ( \43571 , \43570 , \42735 );
xor \U$43195 ( \43572 , \42836 , \42843 );
xor \U$43196 ( \43573 , \43571 , \43572 );
xor \U$43197 ( \43574 , \42866 , \42878 );
xor \U$43198 ( \43575 , \43574 , \42891 );
and \U$43199 ( \43576 , \43573 , \43575 );
xor \U$43200 ( \43577 , \42483 , \42485 );
xor \U$43201 ( \43578 , \43577 , \42488 );
xor \U$43202 ( \43579 , \43136 , \43143 );
xor \U$43203 ( \43580 , \43578 , \43579 );
xor \U$43204 ( \43581 , \42866 , \42878 );
xor \U$43205 ( \43582 , \43581 , \42891 );
and \U$43206 ( \43583 , \43580 , \43582 );
and \U$43207 ( \43584 , \43573 , \43580 );
or \U$43208 ( \43585 , \43576 , \43583 , \43584 );
and \U$43209 ( \43586 , \43569 , \43585 );
and \U$43210 ( \43587 , \43248 , \43568 );
or \U$43211 ( \43588 , \43586 , \43587 );
xor \U$43212 ( \43589 , \42894 , \43133 );
xor \U$43213 ( \43590 , \43589 , \43148 );
xor \U$43214 ( \43591 , \42848 , \42850 );
xor \U$43215 ( \43592 , \43591 , \42853 );
and \U$43216 ( \43593 , \43590 , \43592 );
xor \U$43217 ( \43594 , \42468 , \42480 );
xor \U$43218 ( \43595 , \43594 , \42491 );
xor \U$43219 ( \43596 , \43154 , \43161 );
xor \U$43220 ( \43597 , \43595 , \43596 );
xor \U$43221 ( \43598 , \42848 , \42850 );
xor \U$43222 ( \43599 , \43598 , \42853 );
and \U$43223 ( \43600 , \43597 , \43599 );
and \U$43224 ( \43601 , \43590 , \43597 );
or \U$43225 ( \43602 , \43593 , \43600 , \43601 );
xor \U$43226 ( \43603 , \43588 , \43602 );
xor \U$43227 ( \43604 , \42822 , \42824 );
xor \U$43228 ( \43605 , \43604 , \42831 );
and \U$43229 ( \43606 , \43603 , \43605 );
and \U$43230 ( \43607 , \43588 , \43602 );
or \U$43231 ( \43608 , \43606 , \43607 );
nand \U$43232 ( \43609 , \43218 , \43608 );
nand \U$43233 ( \43610 , \43215 , \43609 );
not \U$43234 ( \43611 , \43610 );
xor \U$43235 ( \43612 , \43175 , \43185 );
xor \U$43236 ( \43613 , \43612 , \43188 );
nor \U$43237 ( \43614 , \43611 , \43613 );
and \U$43238 ( \43615 , \43210 , \43614 );
xor \U$43239 ( \43616 , \43614 , \43210 );
xor \U$43240 ( \43617 , \42856 , \43151 );
xor \U$43241 ( \43618 , \43617 , \43166 );
xor \U$43242 ( \43619 , \43588 , \43602 );
xor \U$43243 ( \43620 , \43619 , \43605 );
and \U$43244 ( \43621 , \43618 , \43620 );
xor \U$43245 ( \43622 , \42975 , \43057 );
xor \U$43246 ( \43623 , \43622 , \43130 );
xor \U$43247 ( \43624 , \43228 , \43230 );
xor \U$43248 ( \43625 , \43624 , \43245 );
and \U$43249 ( \43626 , \43623 , \43625 );
xor \U$43250 ( \43627 , \42866 , \42878 );
xor \U$43251 ( \43628 , \43627 , \42891 );
xor \U$43252 ( \43629 , \43573 , \43580 );
xor \U$43253 ( \43630 , \43628 , \43629 );
xor \U$43254 ( \43631 , \43228 , \43230 );
xor \U$43255 ( \43632 , \43631 , \43245 );
and \U$43256 ( \43633 , \43630 , \43632 );
and \U$43257 ( \43634 , \43623 , \43630 );
or \U$43258 ( \43635 , \43626 , \43633 , \43634 );
xor \U$43259 ( \43636 , \42586 , \42593 );
xor \U$43260 ( \43637 , \43636 , \42601 );
xor \U$43261 ( \43638 , \43494 , \43509 );
xor \U$43262 ( \43639 , \43637 , \43638 );
xor \U$43263 ( \43640 , \43329 , \43411 );
xor \U$43264 ( \43641 , \43640 , \43489 );
xor \U$43265 ( \43642 , \43639 , \43641 );
xor \U$43266 ( \43643 , \43527 , \43551 );
xor \U$43267 ( \43644 , \43643 , \43562 );
and \U$43268 ( \43645 , \43642 , \43644 );
and \U$43269 ( \43646 , \43639 , \43641 );
or \U$43270 ( \43647 , \43645 , \43646 );
xor \U$43271 ( \43648 , \43336 , \43343 );
xor \U$43272 ( \43649 , \43648 , \43351 );
xor \U$43273 ( \43650 , \43361 , \43369 );
xor \U$43274 ( \43651 , \43650 , \43377 );
and \U$43275 ( \43652 , \43649 , \43651 );
xor \U$43276 ( \43653 , \43281 , \43288 );
xor \U$43277 ( \43654 , \43653 , \43297 );
xor \U$43278 ( \43655 , \43361 , \43369 );
xor \U$43279 ( \43656 , \43655 , \43377 );
and \U$43280 ( \43657 , \43654 , \43656 );
and \U$43281 ( \43658 , \43649 , \43654 );
or \U$43282 ( \43659 , \43652 , \43657 , \43658 );
not \U$43283 ( \43660 , \392 );
and \U$43284 ( \43661 , \384 , RIae76fa0_66);
and \U$43285 ( \43662 , RIae76eb0_64, \382 );
nor \U$43286 ( \43663 , \43661 , \43662 );
not \U$43287 ( \43664 , \43663 );
or \U$43288 ( \43665 , \43660 , \43664 );
or \U$43289 ( \43666 , \43663 , \392 );
nand \U$43290 ( \43667 , \43665 , \43666 );
not \U$43291 ( \43668 , RIae77900_86);
nor \U$43292 ( \43669 , \43668 , \491 );
xor \U$43293 ( \43670 , \43667 , \43669 );
not \U$43294 ( \43671 , \400 );
and \U$43295 ( \43672 , \436 , RIae76dc0_62);
and \U$43296 ( \43673 , RIae76cd0_60, \434 );
nor \U$43297 ( \43674 , \43672 , \43673 );
not \U$43298 ( \43675 , \43674 );
or \U$43299 ( \43676 , \43671 , \43675 );
or \U$43300 ( \43677 , \43674 , \400 );
nand \U$43301 ( \43678 , \43676 , \43677 );
and \U$43302 ( \43679 , \43670 , \43678 );
and \U$43303 ( \43680 , \43667 , \43669 );
or \U$43304 ( \43681 , \43679 , \43680 );
or \U$43305 ( \43682 , \43547 , \43539 );
nand \U$43306 ( \43683 , \43682 , \43548 );
xor \U$43307 ( \43684 , \43681 , \43683 );
xor \U$43308 ( \43685 , \43389 , \43397 );
xor \U$43309 ( \43686 , \43685 , \43405 );
and \U$43310 ( \43687 , \43684 , \43686 );
and \U$43311 ( \43688 , \43681 , \43683 );
or \U$43312 ( \43689 , \43687 , \43688 );
xor \U$43313 ( \43690 , \43659 , \43689 );
xor \U$43314 ( \43691 , \43308 , \43315 );
xor \U$43315 ( \43692 , \43691 , \43323 );
xor \U$43316 ( \43693 , \43255 , \43263 );
xor \U$43317 ( \43694 , \43693 , \43271 );
and \U$43318 ( \43695 , \43692 , \43694 );
xor \U$43319 ( \43696 , \43419 , \43426 );
xor \U$43320 ( \43697 , \43696 , \43434 );
xor \U$43321 ( \43698 , \43255 , \43263 );
xor \U$43322 ( \43699 , \43698 , \43271 );
and \U$43323 ( \43700 , \43697 , \43699 );
and \U$43324 ( \43701 , \43692 , \43697 );
or \U$43325 ( \43702 , \43695 , \43700 , \43701 );
and \U$43326 ( \43703 , \43690 , \43702 );
and \U$43327 ( \43704 , \43659 , \43689 );
or \U$43328 ( \43705 , \43703 , \43704 );
and \U$43329 ( \43706 , \1939 , RIae77db0_96);
and \U$43330 ( \43707 , RIae77ea0_98, \1937 );
nor \U$43331 ( \43708 , \43706 , \43707 );
and \U$43332 ( \43709 , \43708 , \1735 );
not \U$43333 ( \43710 , \43708 );
and \U$43334 ( \43711 , \43710 , \1734 );
nor \U$43335 ( \43712 , \43709 , \43711 );
and \U$43336 ( \43713 , \1593 , RIae77cc0_94);
and \U$43337 ( \43714 , RIae77bd0_92, \1591 );
nor \U$43338 ( \43715 , \43713 , \43714 );
and \U$43339 ( \43716 , \43715 , \1498 );
not \U$43340 ( \43717 , \43715 );
and \U$43341 ( \43718 , \43717 , \1488 );
nor \U$43342 ( \43719 , \43716 , \43718 );
xor \U$43343 ( \43720 , \43712 , \43719 );
and \U$43344 ( \43721 , \2224 , RIae789e0_122);
and \U$43345 ( \43722 , RIae788f0_120, \2222 );
nor \U$43346 ( \43723 , \43721 , \43722 );
and \U$43347 ( \43724 , \43723 , \2061 );
not \U$43348 ( \43725 , \43723 );
and \U$43349 ( \43726 , \43725 , \2060 );
nor \U$43350 ( \43727 , \43724 , \43726 );
and \U$43351 ( \43728 , \43720 , \43727 );
and \U$43352 ( \43729 , \43712 , \43719 );
or \U$43353 ( \43730 , \43728 , \43729 );
and \U$43354 ( \43731 , \1376 , RIae78440_110);
and \U$43355 ( \43732 , RIae784b8_111, \1374 );
nor \U$43356 ( \43733 , \43731 , \43732 );
and \U$43357 ( \43734 , \43733 , \1380 );
not \U$43358 ( \43735 , \43733 );
and \U$43359 ( \43736 , \43735 , \1261 );
nor \U$43360 ( \43737 , \43734 , \43736 );
not \U$43361 ( \43738 , \787 );
and \U$43362 ( \43739 , \883 , RIae77f90_100);
and \U$43363 ( \43740 , RIae78080_102, \881 );
nor \U$43364 ( \43741 , \43739 , \43740 );
not \U$43365 ( \43742 , \43741 );
or \U$43366 ( \43743 , \43738 , \43742 );
or \U$43367 ( \43744 , \43741 , \787 );
nand \U$43368 ( \43745 , \43743 , \43744 );
xor \U$43369 ( \43746 , \43737 , \43745 );
and \U$43370 ( \43747 , \1138 , RIae78260_106);
and \U$43371 ( \43748 , RIae78620_114, \1136 );
nor \U$43372 ( \43749 , \43747 , \43748 );
and \U$43373 ( \43750 , \43749 , \1012 );
not \U$43374 ( \43751 , \43749 );
and \U$43375 ( \43752 , \43751 , \1142 );
nor \U$43376 ( \43753 , \43750 , \43752 );
and \U$43377 ( \43754 , \43746 , \43753 );
and \U$43378 ( \43755 , \43737 , \43745 );
or \U$43379 ( \43756 , \43754 , \43755 );
xor \U$43380 ( \43757 , \43730 , \43756 );
and \U$43381 ( \43758 , \672 , RIae78350_108);
and \U$43382 ( \43759 , RIae78170_104, \670 );
nor \U$43383 ( \43760 , \43758 , \43759 );
and \U$43384 ( \43761 , \43760 , \588 );
not \U$43385 ( \43762 , \43760 );
and \U$43386 ( \43763 , \43762 , \587 );
nor \U$43387 ( \43764 , \43761 , \43763 );
not \U$43388 ( \43765 , \469 );
and \U$43389 ( \43766 , \514 , RIae77108_69);
and \U$43390 ( \43767 , RIae77090_68, \512 );
nor \U$43391 ( \43768 , \43766 , \43767 );
not \U$43392 ( \43769 , \43768 );
or \U$43393 ( \43770 , \43765 , \43769 );
or \U$43394 ( \43771 , \43768 , \469 );
nand \U$43395 ( \43772 , \43770 , \43771 );
xor \U$43396 ( \43773 , \43764 , \43772 );
and \U$43397 ( \43774 , \558 , RIae77270_72);
and \U$43398 ( \43775 , RIae77360_74, \556 );
nor \U$43399 ( \43776 , \43774 , \43775 );
and \U$43400 ( \43777 , \43776 , \504 );
not \U$43401 ( \43778 , \43776 );
and \U$43402 ( \43779 , \43778 , \562 );
nor \U$43403 ( \43780 , \43777 , \43779 );
and \U$43404 ( \43781 , \43773 , \43780 );
and \U$43405 ( \43782 , \43764 , \43772 );
or \U$43406 ( \43783 , \43781 , \43782 );
and \U$43407 ( \43784 , \43757 , \43783 );
and \U$43408 ( \43785 , \43730 , \43756 );
or \U$43409 ( \43786 , \43784 , \43785 );
and \U$43410 ( \43787 , \7633 , RIae76730_48);
and \U$43411 ( \43788 , RIae76640_46, \7631 );
nor \U$43412 ( \43789 , \43787 , \43788 );
and \U$43413 ( \43790 , \43789 , \7206 );
not \U$43414 ( \43791 , \43789 );
and \U$43415 ( \43792 , \43791 , \7205 );
nor \U$43416 ( \43793 , \43790 , \43792 );
and \U$43417 ( \43794 , \6941 , RIae76460_42);
and \U$43418 ( \43795 , RIae76550_44, \6939 );
nor \U$43419 ( \43796 , \43794 , \43795 );
and \U$43420 ( \43797 , \43796 , \6314 );
not \U$43421 ( \43798 , \43796 );
and \U$43422 ( \43799 , \43798 , \6945 );
nor \U$43423 ( \43800 , \43797 , \43799 );
xor \U$43424 ( \43801 , \43793 , \43800 );
and \U$43425 ( \43802 , \8371 , RIae76190_36);
and \U$43426 ( \43803 , RIae760a0_34, \8369 );
nor \U$43427 ( \43804 , \43802 , \43803 );
and \U$43428 ( \43805 , \43804 , \8020 );
not \U$43429 ( \43806 , \43804 );
and \U$43430 ( \43807 , \43806 , \8019 );
nor \U$43431 ( \43808 , \43805 , \43807 );
and \U$43432 ( \43809 , \43801 , \43808 );
and \U$43433 ( \43810 , \43793 , \43800 );
or \U$43434 ( \43811 , \43809 , \43810 );
and \U$43435 ( \43812 , \11470 , RIae76be0_58);
and \U$43436 ( \43813 , RIae78ad0_124, \11468 );
nor \U$43437 ( \43814 , \43812 , \43813 );
and \U$43438 ( \43815 , \43814 , \10936 );
not \U$43439 ( \43816 , \43814 );
and \U$43440 ( \43817 , \43816 , \11474 );
nor \U$43441 ( \43818 , \43815 , \43817 );
xor \U$43442 ( \43819 , \43818 , \13063 );
and \U$43443 ( \43820 , \12180 , RIae78d28_129);
and \U$43444 ( \43821 , RIae78e18_131, \12178 );
nor \U$43445 ( \43822 , \43820 , \43821 );
and \U$43446 ( \43823 , \43822 , \12184 );
not \U$43447 ( \43824 , \43822 );
and \U$43448 ( \43825 , \43824 , \11827 );
nor \U$43449 ( \43826 , \43823 , \43825 );
and \U$43450 ( \43827 , \43819 , \43826 );
and \U$43451 ( \43828 , \43818 , \13063 );
or \U$43452 ( \43829 , \43827 , \43828 );
xor \U$43453 ( \43830 , \43811 , \43829 );
and \U$43454 ( \43831 , \8966 , RIae76370_40);
and \U$43455 ( \43832 , RIae76280_38, \8964 );
nor \U$43456 ( \43833 , \43831 , \43832 );
and \U$43457 ( \43834 , \43833 , \8799 );
not \U$43458 ( \43835 , \43833 );
and \U$43459 ( \43836 , \43835 , \8789 );
nor \U$43460 ( \43837 , \43834 , \43836 );
and \U$43461 ( \43838 , \9760 , RIae76af0_56);
and \U$43462 ( \43839 , RIae76a00_54, \9758 );
nor \U$43463 ( \43840 , \43838 , \43839 );
and \U$43464 ( \43841 , \43840 , \9273 );
not \U$43465 ( \43842 , \43840 );
and \U$43466 ( \43843 , \43842 , \9272 );
nor \U$43467 ( \43844 , \43841 , \43843 );
xor \U$43468 ( \43845 , \43837 , \43844 );
and \U$43469 ( \43846 , \10548 , RIae76820_50);
and \U$43470 ( \43847 , RIae76910_52, \10546 );
nor \U$43471 ( \43848 , \43846 , \43847 );
and \U$43472 ( \43849 , \43848 , \10421 );
not \U$43473 ( \43850 , \43848 );
and \U$43474 ( \43851 , \43850 , \10118 );
nor \U$43475 ( \43852 , \43849 , \43851 );
and \U$43476 ( \43853 , \43845 , \43852 );
and \U$43477 ( \43854 , \43837 , \43844 );
or \U$43478 ( \43855 , \43853 , \43854 );
and \U$43479 ( \43856 , \43830 , \43855 );
and \U$43480 ( \43857 , \43811 , \43829 );
or \U$43481 ( \43858 , \43856 , \43857 );
xor \U$43482 ( \43859 , \43786 , \43858 );
and \U$43483 ( \43860 , \5896 , RIae75290_4);
and \U$43484 ( \43861 , RIae751a0_2, \5894 );
nor \U$43485 ( \43862 , \43860 , \43861 );
and \U$43486 ( \43863 , \43862 , \5590 );
not \U$43487 ( \43864 , \43862 );
and \U$43488 ( \43865 , \43864 , \5589 );
nor \U$43489 ( \43866 , \43863 , \43865 );
and \U$43490 ( \43867 , \5399 , RIae75830_16);
and \U$43491 ( \43868 , RIae75740_14, \5397 );
nor \U$43492 ( \43869 , \43867 , \43868 );
and \U$43493 ( \43870 , \43869 , \5016 );
not \U$43494 ( \43871 , \43869 );
and \U$43495 ( \43872 , \43871 , \5403 );
nor \U$43496 ( \43873 , \43870 , \43872 );
xor \U$43497 ( \43874 , \43866 , \43873 );
and \U$43498 ( \43875 , \6172 , RIae75380_6);
and \U$43499 ( \43876 , RIae75470_8, \6170 );
nor \U$43500 ( \43877 , \43875 , \43876 );
and \U$43501 ( \43878 , \43877 , \6176 );
not \U$43502 ( \43879 , \43877 );
and \U$43503 ( \43880 , \43879 , \6175 );
nor \U$43504 ( \43881 , \43878 , \43880 );
and \U$43505 ( \43882 , \43874 , \43881 );
and \U$43506 ( \43883 , \43866 , \43873 );
or \U$43507 ( \43884 , \43882 , \43883 );
and \U$43508 ( \43885 , \4247 , RIae75ce0_26);
and \U$43509 ( \43886 , RIae75dd0_28, \4245 );
nor \U$43510 ( \43887 , \43885 , \43886 );
and \U$43511 ( \43888 , \43887 , \3989 );
not \U$43512 ( \43889 , \43887 );
and \U$43513 ( \43890 , \43889 , \4251 );
nor \U$43514 ( \43891 , \43888 , \43890 );
and \U$43515 ( \43892 , \3730 , RIae75fb0_32);
and \U$43516 ( \43893 , RIae75ec0_30, \3728 );
nor \U$43517 ( \43894 , \43892 , \43893 );
and \U$43518 ( \43895 , \43894 , \3732 );
not \U$43519 ( \43896 , \43894 );
and \U$43520 ( \43897 , \43896 , \3422 );
nor \U$43521 ( \43898 , \43895 , \43897 );
xor \U$43522 ( \43899 , \43891 , \43898 );
and \U$43523 ( \43900 , \4688 , RIae75650_12);
and \U$43524 ( \43901 , RIae75560_10, \4686 );
nor \U$43525 ( \43902 , \43900 , \43901 );
and \U$43526 ( \43903 , \43902 , \4481 );
not \U$43527 ( \43904 , \43902 );
and \U$43528 ( \43905 , \43904 , \4482 );
nor \U$43529 ( \43906 , \43903 , \43905 );
and \U$43530 ( \43907 , \43899 , \43906 );
and \U$43531 ( \43908 , \43891 , \43898 );
or \U$43532 ( \43909 , \43907 , \43908 );
xor \U$43533 ( \43910 , \43884 , \43909 );
and \U$43534 ( \43911 , \2607 , RIae78800_118);
and \U$43535 ( \43912 , RIae78710_116, \2605 );
nor \U$43536 ( \43913 , \43911 , \43912 );
and \U$43537 ( \43914 , \43913 , \2611 );
not \U$43538 ( \43915 , \43913 );
and \U$43539 ( \43916 , \43915 , \2397 );
nor \U$43540 ( \43917 , \43914 , \43916 );
not \U$43541 ( \43918 , \2789 );
and \U$43542 ( \43919 , \2783 , RIae75bf0_24);
and \U$43543 ( \43920 , RIae75b00_22, \2781 );
nor \U$43544 ( \43921 , \43919 , \43920 );
not \U$43545 ( \43922 , \43921 );
or \U$43546 ( \43923 , \43918 , \43922 );
or \U$43547 ( \43924 , \43921 , \3089 );
nand \U$43548 ( \43925 , \43923 , \43924 );
xor \U$43549 ( \43926 , \43917 , \43925 );
not \U$43550 ( \43927 , \2774 );
and \U$43551 ( \43928 , \3214 , RIae75a10_20);
and \U$43552 ( \43929 , RIae75920_18, \3212 );
nor \U$43553 ( \43930 , \43928 , \43929 );
not \U$43554 ( \43931 , \43930 );
or \U$43555 ( \43932 , \43927 , \43931 );
or \U$43556 ( \43933 , \43930 , \2774 );
nand \U$43557 ( \43934 , \43932 , \43933 );
and \U$43558 ( \43935 , \43926 , \43934 );
and \U$43559 ( \43936 , \43917 , \43925 );
or \U$43560 ( \43937 , \43935 , \43936 );
and \U$43561 ( \43938 , \43910 , \43937 );
and \U$43562 ( \43939 , \43884 , \43909 );
or \U$43563 ( \43940 , \43938 , \43939 );
and \U$43564 ( \43941 , \43859 , \43940 );
and \U$43565 ( \43942 , \43786 , \43858 );
or \U$43566 ( \43943 , \43941 , \43942 );
xor \U$43567 ( \43944 , \43705 , \43943 );
xor \U$43568 ( \43945 , \43065 , \43072 );
xor \U$43569 ( \43946 , \43945 , \43080 );
xor \U$43570 ( \43947 , \43499 , \43504 );
xor \U$43571 ( \43948 , \43946 , \43947 );
xor \U$43572 ( \43949 , \43554 , \43556 );
xor \U$43573 ( \43950 , \43949 , \43559 );
and \U$43574 ( \43951 , \43948 , \43950 );
xor \U$43575 ( \43952 , \42901 , \42908 );
xor \U$43576 ( \43953 , \43952 , \42916 );
xor \U$43577 ( \43954 , \43517 , \43522 );
xor \U$43578 ( \43955 , \43953 , \43954 );
xor \U$43579 ( \43956 , \43554 , \43556 );
xor \U$43580 ( \43957 , \43956 , \43559 );
and \U$43581 ( \43958 , \43955 , \43957 );
and \U$43582 ( \43959 , \43948 , \43955 );
or \U$43583 ( \43960 , \43951 , \43958 , \43959 );
and \U$43584 ( \43961 , \43944 , \43960 );
and \U$43585 ( \43962 , \43705 , \43943 );
or \U$43586 ( \43963 , \43961 , \43962 );
xor \U$43587 ( \43964 , \43647 , \43963 );
xor \U$43588 ( \43965 , \43535 , \43537 );
xor \U$43589 ( \43966 , \43965 , \43548 );
xor \U$43590 ( \43967 , \43354 , \43380 );
xor \U$43591 ( \43968 , \43967 , \43408 );
and \U$43592 ( \43969 , \43966 , \43968 );
xor \U$43593 ( \43970 , \43274 , \43300 );
xor \U$43594 ( \43971 , \43970 , \43326 );
xor \U$43595 ( \43972 , \43354 , \43380 );
xor \U$43596 ( \43973 , \43972 , \43408 );
and \U$43597 ( \43974 , \43971 , \43973 );
and \U$43598 ( \43975 , \43966 , \43971 );
or \U$43599 ( \43976 , \43969 , \43974 , \43975 );
xor \U$43600 ( \43977 , \43220 , \43222 );
xor \U$43601 ( \43978 , \43977 , \43225 );
and \U$43602 ( \43979 , \43976 , \43978 );
xor \U$43603 ( \43980 , \42858 , \42860 );
xor \U$43604 ( \43981 , \43980 , \42863 );
xor \U$43605 ( \43982 , \43233 , \43240 );
xor \U$43606 ( \43983 , \43981 , \43982 );
xor \U$43607 ( \43984 , \43220 , \43222 );
xor \U$43608 ( \43985 , \43984 , \43225 );
and \U$43609 ( \43986 , \43983 , \43985 );
and \U$43610 ( \43987 , \43976 , \43983 );
or \U$43611 ( \43988 , \43979 , \43986 , \43987 );
and \U$43612 ( \43989 , \43964 , \43988 );
and \U$43613 ( \43990 , \43647 , \43963 );
or \U$43614 ( \43991 , \43989 , \43990 );
xor \U$43615 ( \43992 , \43635 , \43991 );
xor \U$43616 ( \43993 , \42848 , \42850 );
xor \U$43617 ( \43994 , \43993 , \42853 );
xor \U$43618 ( \43995 , \43590 , \43597 );
xor \U$43619 ( \43996 , \43994 , \43995 );
and \U$43620 ( \43997 , \43992 , \43996 );
and \U$43621 ( \43998 , \43635 , \43991 );
or \U$43622 ( \43999 , \43997 , \43998 );
xor \U$43623 ( \44000 , \43588 , \43602 );
xor \U$43624 ( \44001 , \44000 , \43605 );
and \U$43625 ( \44002 , \43999 , \44001 );
and \U$43626 ( \44003 , \43618 , \43999 );
or \U$43627 ( \44004 , \43621 , \44002 , \44003 );
not \U$43628 ( \44005 , \44004 );
not \U$43629 ( \44006 , \43214 );
not \U$43630 ( \44007 , \43608 );
or \U$43631 ( \44008 , \44006 , \44007 );
or \U$43632 ( \44009 , \43608 , \43214 );
nand \U$43633 ( \44010 , \44008 , \44009 );
not \U$43634 ( \44011 , \44010 );
not \U$43635 ( \44012 , \43212 );
and \U$43636 ( \44013 , \44011 , \44012 );
and \U$43637 ( \44014 , \44010 , \43212 );
nor \U$43638 ( \44015 , \44013 , \44014 );
not \U$43639 ( \44016 , \44015 );
or \U$43640 ( \44017 , \44005 , \44016 );
or \U$43641 ( \44018 , \44015 , \44004 );
nand \U$43642 ( \44019 , \44017 , \44018 );
xor \U$43643 ( \44020 , \43647 , \43963 );
xor \U$43644 ( \44021 , \44020 , \43988 );
xor \U$43645 ( \44022 , \43228 , \43230 );
xor \U$43646 ( \44023 , \44022 , \43245 );
xor \U$43647 ( \44024 , \43623 , \43630 );
xor \U$43648 ( \44025 , \44023 , \44024 );
and \U$43649 ( \44026 , \44021 , \44025 );
xor \U$43650 ( \44027 , \43248 , \43568 );
xor \U$43651 ( \44028 , \44027 , \43585 );
xor \U$43652 ( \44029 , \44026 , \44028 );
xor \U$43653 ( \44030 , \43786 , \43858 );
xor \U$43654 ( \44031 , \44030 , \43940 );
xor \U$43655 ( \44032 , \43659 , \43689 );
xor \U$43656 ( \44033 , \44032 , \43702 );
and \U$43657 ( \44034 , \44031 , \44033 );
xor \U$43658 ( \44035 , \43554 , \43556 );
xor \U$43659 ( \44036 , \44035 , \43559 );
xor \U$43660 ( \44037 , \43948 , \43955 );
xor \U$43661 ( \44038 , \44036 , \44037 );
xor \U$43662 ( \44039 , \43659 , \43689 );
xor \U$43663 ( \44040 , \44039 , \43702 );
and \U$43664 ( \44041 , \44038 , \44040 );
and \U$43665 ( \44042 , \44031 , \44038 );
or \U$43666 ( \44043 , \44034 , \44041 , \44042 );
and \U$43667 ( \44044 , \5399 , RIae75560_10);
and \U$43668 ( \44045 , RIae75830_16, \5397 );
nor \U$43669 ( \44046 , \44044 , \44045 );
and \U$43670 ( \44047 , \44046 , \5016 );
not \U$43671 ( \44048 , \44046 );
and \U$43672 ( \44049 , \44048 , \5403 );
nor \U$43673 ( \44050 , \44047 , \44049 );
and \U$43674 ( \44051 , \5896 , RIae75740_14);
and \U$43675 ( \44052 , RIae75290_4, \5894 );
nor \U$43676 ( \44053 , \44051 , \44052 );
and \U$43677 ( \44054 , \44053 , \5590 );
not \U$43678 ( \44055 , \44053 );
and \U$43679 ( \44056 , \44055 , \5589 );
nor \U$43680 ( \44057 , \44054 , \44056 );
xor \U$43681 ( \44058 , \44050 , \44057 );
and \U$43682 ( \44059 , \6172 , RIae751a0_2);
and \U$43683 ( \44060 , RIae75380_6, \6170 );
nor \U$43684 ( \44061 , \44059 , \44060 );
and \U$43685 ( \44062 , \44061 , \6176 );
not \U$43686 ( \44063 , \44061 );
and \U$43687 ( \44064 , \44063 , \6175 );
nor \U$43688 ( \44065 , \44062 , \44064 );
and \U$43689 ( \44066 , \44058 , \44065 );
and \U$43690 ( \44067 , \44050 , \44057 );
or \U$43691 ( \44068 , \44066 , \44067 );
not \U$43692 ( \44069 , \3218 );
and \U$43693 ( \44070 , \3214 , RIae75b00_22);
and \U$43694 ( \44071 , RIae75a10_20, \3212 );
nor \U$43695 ( \44072 , \44070 , \44071 );
not \U$43696 ( \44073 , \44072 );
or \U$43697 ( \44074 , \44069 , \44073 );
or \U$43698 ( \44075 , \44072 , \3218 );
nand \U$43699 ( \44076 , \44074 , \44075 );
and \U$43700 ( \44077 , \2607 , RIae788f0_120);
and \U$43701 ( \44078 , RIae78800_118, \2605 );
nor \U$43702 ( \44079 , \44077 , \44078 );
and \U$43703 ( \44080 , \44079 , \2611 );
not \U$43704 ( \44081 , \44079 );
and \U$43705 ( \44082 , \44081 , \2397 );
nor \U$43706 ( \44083 , \44080 , \44082 );
xor \U$43707 ( \44084 , \44076 , \44083 );
not \U$43708 ( \44085 , \2789 );
and \U$43709 ( \44086 , \2783 , RIae78710_116);
and \U$43710 ( \44087 , RIae75bf0_24, \2781 );
nor \U$43711 ( \44088 , \44086 , \44087 );
not \U$43712 ( \44089 , \44088 );
or \U$43713 ( \44090 , \44085 , \44089 );
or \U$43714 ( \44091 , \44088 , \3089 );
nand \U$43715 ( \44092 , \44090 , \44091 );
and \U$43716 ( \44093 , \44084 , \44092 );
and \U$43717 ( \44094 , \44076 , \44083 );
or \U$43718 ( \44095 , \44093 , \44094 );
xor \U$43719 ( \44096 , \44068 , \44095 );
and \U$43720 ( \44097 , \3730 , RIae75920_18);
and \U$43721 ( \44098 , RIae75fb0_32, \3728 );
nor \U$43722 ( \44099 , \44097 , \44098 );
and \U$43723 ( \44100 , \44099 , \3732 );
not \U$43724 ( \44101 , \44099 );
and \U$43725 ( \44102 , \44101 , \3422 );
nor \U$43726 ( \44103 , \44100 , \44102 );
and \U$43727 ( \44104 , \4247 , RIae75ec0_30);
and \U$43728 ( \44105 , RIae75ce0_26, \4245 );
nor \U$43729 ( \44106 , \44104 , \44105 );
and \U$43730 ( \44107 , \44106 , \3989 );
not \U$43731 ( \44108 , \44106 );
and \U$43732 ( \44109 , \44108 , \4251 );
nor \U$43733 ( \44110 , \44107 , \44109 );
xor \U$43734 ( \44111 , \44103 , \44110 );
and \U$43735 ( \44112 , \4688 , RIae75dd0_28);
and \U$43736 ( \44113 , RIae75650_12, \4686 );
nor \U$43737 ( \44114 , \44112 , \44113 );
and \U$43738 ( \44115 , \44114 , \4481 );
not \U$43739 ( \44116 , \44114 );
and \U$43740 ( \44117 , \44116 , \4482 );
nor \U$43741 ( \44118 , \44115 , \44117 );
and \U$43742 ( \44119 , \44111 , \44118 );
and \U$43743 ( \44120 , \44103 , \44110 );
or \U$43744 ( \44121 , \44119 , \44120 );
and \U$43745 ( \44122 , \44096 , \44121 );
and \U$43746 ( \44123 , \44068 , \44095 );
or \U$43747 ( \44124 , \44122 , \44123 );
not \U$43748 ( \44125 , \787 );
and \U$43749 ( \44126 , \883 , RIae78170_104);
and \U$43750 ( \44127 , RIae77f90_100, \881 );
nor \U$43751 ( \44128 , \44126 , \44127 );
not \U$43752 ( \44129 , \44128 );
or \U$43753 ( \44130 , \44125 , \44129 );
or \U$43754 ( \44131 , \44128 , \789 );
nand \U$43755 ( \44132 , \44130 , \44131 );
and \U$43756 ( \44133 , \1138 , RIae78080_102);
and \U$43757 ( \44134 , RIae78260_106, \1136 );
nor \U$43758 ( \44135 , \44133 , \44134 );
and \U$43759 ( \44136 , \44135 , \1012 );
not \U$43760 ( \44137 , \44135 );
and \U$43761 ( \44138 , \44137 , \1142 );
nor \U$43762 ( \44139 , \44136 , \44138 );
xor \U$43763 ( \44140 , \44132 , \44139 );
and \U$43764 ( \44141 , \1376 , RIae78620_114);
and \U$43765 ( \44142 , RIae78440_110, \1374 );
nor \U$43766 ( \44143 , \44141 , \44142 );
and \U$43767 ( \44144 , \44143 , \1380 );
not \U$43768 ( \44145 , \44143 );
and \U$43769 ( \44146 , \44145 , \1261 );
nor \U$43770 ( \44147 , \44144 , \44146 );
and \U$43771 ( \44148 , \44140 , \44147 );
and \U$43772 ( \44149 , \44132 , \44139 );
or \U$43773 ( \44150 , \44148 , \44149 );
and \U$43774 ( \44151 , \558 , RIae77090_68);
and \U$43775 ( \44152 , RIae77270_72, \556 );
nor \U$43776 ( \44153 , \44151 , \44152 );
and \U$43777 ( \44154 , \44153 , \504 );
not \U$43778 ( \44155 , \44153 );
and \U$43779 ( \44156 , \44155 , \562 );
nor \U$43780 ( \44157 , \44154 , \44156 );
not \U$43781 ( \44158 , \469 );
and \U$43782 ( \44159 , \514 , RIae76cd0_60);
and \U$43783 ( \44160 , RIae77108_69, \512 );
nor \U$43784 ( \44161 , \44159 , \44160 );
not \U$43785 ( \44162 , \44161 );
or \U$43786 ( \44163 , \44158 , \44162 );
or \U$43787 ( \44164 , \44161 , \469 );
nand \U$43788 ( \44165 , \44163 , \44164 );
xor \U$43789 ( \44166 , \44157 , \44165 );
and \U$43790 ( \44167 , \672 , RIae77360_74);
and \U$43791 ( \44168 , RIae78350_108, \670 );
nor \U$43792 ( \44169 , \44167 , \44168 );
and \U$43793 ( \44170 , \44169 , \588 );
not \U$43794 ( \44171 , \44169 );
and \U$43795 ( \44172 , \44171 , \587 );
nor \U$43796 ( \44173 , \44170 , \44172 );
and \U$43797 ( \44174 , \44166 , \44173 );
and \U$43798 ( \44175 , \44157 , \44165 );
or \U$43799 ( \44176 , \44174 , \44175 );
xor \U$43800 ( \44177 , \44150 , \44176 );
and \U$43801 ( \44178 , \1593 , RIae784b8_111);
and \U$43802 ( \44179 , RIae77cc0_94, \1591 );
nor \U$43803 ( \44180 , \44178 , \44179 );
and \U$43804 ( \44181 , \44180 , \1498 );
not \U$43805 ( \44182 , \44180 );
and \U$43806 ( \44183 , \44182 , \1488 );
nor \U$43807 ( \44184 , \44181 , \44183 );
and \U$43808 ( \44185 , \1939 , RIae77bd0_92);
and \U$43809 ( \44186 , RIae77db0_96, \1937 );
nor \U$43810 ( \44187 , \44185 , \44186 );
and \U$43811 ( \44188 , \44187 , \1735 );
not \U$43812 ( \44189 , \44187 );
and \U$43813 ( \44190 , \44189 , \1734 );
nor \U$43814 ( \44191 , \44188 , \44190 );
xor \U$43815 ( \44192 , \44184 , \44191 );
and \U$43816 ( \44193 , \2224 , RIae77ea0_98);
and \U$43817 ( \44194 , RIae789e0_122, \2222 );
nor \U$43818 ( \44195 , \44193 , \44194 );
and \U$43819 ( \44196 , \44195 , \2061 );
not \U$43820 ( \44197 , \44195 );
and \U$43821 ( \44198 , \44197 , \2060 );
nor \U$43822 ( \44199 , \44196 , \44198 );
and \U$43823 ( \44200 , \44192 , \44199 );
and \U$43824 ( \44201 , \44184 , \44191 );
or \U$43825 ( \44202 , \44200 , \44201 );
and \U$43826 ( \44203 , \44177 , \44202 );
and \U$43827 ( \44204 , \44150 , \44176 );
or \U$43828 ( \44205 , \44203 , \44204 );
xor \U$43829 ( \44206 , \44124 , \44205 );
and \U$43830 ( \44207 , \6941 , RIae75470_8);
and \U$43831 ( \44208 , RIae76460_42, \6939 );
nor \U$43832 ( \44209 , \44207 , \44208 );
and \U$43833 ( \44210 , \44209 , \6314 );
not \U$43834 ( \44211 , \44209 );
and \U$43835 ( \44212 , \44211 , \6945 );
nor \U$43836 ( \44213 , \44210 , \44212 );
and \U$43837 ( \44214 , \7633 , RIae76550_44);
and \U$43838 ( \44215 , RIae76730_48, \7631 );
nor \U$43839 ( \44216 , \44214 , \44215 );
and \U$43840 ( \44217 , \44216 , \7206 );
not \U$43841 ( \44218 , \44216 );
and \U$43842 ( \44219 , \44218 , \7205 );
nor \U$43843 ( \44220 , \44217 , \44219 );
xor \U$43844 ( \44221 , \44213 , \44220 );
and \U$43845 ( \44222 , \8371 , RIae76640_46);
and \U$43846 ( \44223 , RIae76190_36, \8369 );
nor \U$43847 ( \44224 , \44222 , \44223 );
and \U$43848 ( \44225 , \44224 , \8020 );
not \U$43849 ( \44226 , \44224 );
and \U$43850 ( \44227 , \44226 , \8019 );
nor \U$43851 ( \44228 , \44225 , \44227 );
and \U$43852 ( \44229 , \44221 , \44228 );
and \U$43853 ( \44230 , \44213 , \44220 );
or \U$43854 ( \44231 , \44229 , \44230 );
and \U$43855 ( \44232 , \11470 , RIae76910_52);
and \U$43856 ( \44233 , RIae76be0_58, \11468 );
nor \U$43857 ( \44234 , \44232 , \44233 );
and \U$43858 ( \44235 , \44234 , \10936 );
not \U$43859 ( \44236 , \44234 );
and \U$43860 ( \44237 , \44236 , \11474 );
nor \U$43861 ( \44238 , \44235 , \44237 );
nand \U$43862 ( \44239 , RIae78e18_131, \13059 );
and \U$43863 ( \44240 , \44239 , \13063 );
not \U$43864 ( \44241 , \44239 );
and \U$43865 ( \44242 , \44241 , \12718 );
nor \U$43866 ( \44243 , \44240 , \44242 );
xor \U$43867 ( \44244 , \44238 , \44243 );
and \U$43868 ( \44245 , \12180 , RIae78ad0_124);
and \U$43869 ( \44246 , RIae78d28_129, \12178 );
nor \U$43870 ( \44247 , \44245 , \44246 );
and \U$43871 ( \44248 , \44247 , \12184 );
not \U$43872 ( \44249 , \44247 );
and \U$43873 ( \44250 , \44249 , \11827 );
nor \U$43874 ( \44251 , \44248 , \44250 );
and \U$43875 ( \44252 , \44244 , \44251 );
and \U$43876 ( \44253 , \44238 , \44243 );
or \U$43877 ( \44254 , \44252 , \44253 );
xor \U$43878 ( \44255 , \44231 , \44254 );
and \U$43879 ( \44256 , \8966 , RIae760a0_34);
and \U$43880 ( \44257 , RIae76370_40, \8964 );
nor \U$43881 ( \44258 , \44256 , \44257 );
and \U$43882 ( \44259 , \44258 , \8799 );
not \U$43883 ( \44260 , \44258 );
and \U$43884 ( \44261 , \44260 , \8789 );
nor \U$43885 ( \44262 , \44259 , \44261 );
and \U$43886 ( \44263 , \9760 , RIae76280_38);
and \U$43887 ( \44264 , RIae76af0_56, \9758 );
nor \U$43888 ( \44265 , \44263 , \44264 );
and \U$43889 ( \44266 , \44265 , \9273 );
not \U$43890 ( \44267 , \44265 );
and \U$43891 ( \44268 , \44267 , \9764 );
nor \U$43892 ( \44269 , \44266 , \44268 );
xor \U$43893 ( \44270 , \44262 , \44269 );
and \U$43894 ( \44271 , \10548 , RIae76a00_54);
and \U$43895 ( \44272 , RIae76820_50, \10546 );
nor \U$43896 ( \44273 , \44271 , \44272 );
and \U$43897 ( \44274 , \44273 , \10421 );
not \U$43898 ( \44275 , \44273 );
and \U$43899 ( \44276 , \44275 , \10118 );
nor \U$43900 ( \44277 , \44274 , \44276 );
and \U$43901 ( \44278 , \44270 , \44277 );
and \U$43902 ( \44279 , \44262 , \44269 );
or \U$43903 ( \44280 , \44278 , \44279 );
and \U$43904 ( \44281 , \44255 , \44280 );
and \U$43905 ( \44282 , \44231 , \44254 );
or \U$43906 ( \44283 , \44281 , \44282 );
and \U$43907 ( \44284 , \44206 , \44283 );
and \U$43908 ( \44285 , \44124 , \44205 );
or \U$43909 ( \44286 , \44284 , \44285 );
xor \U$43910 ( \44287 , \43468 , \43475 );
xor \U$43911 ( \44288 , \44287 , \43483 );
xor \U$43912 ( \44289 , \43444 , \43449 );
xor \U$43913 ( \44290 , \44289 , \43457 );
xor \U$43914 ( \44291 , \44288 , \44290 );
xor \U$43915 ( \44292 , \43255 , \43263 );
xor \U$43916 ( \44293 , \44292 , \43271 );
xor \U$43917 ( \44294 , \43692 , \43697 );
xor \U$43918 ( \44295 , \44293 , \44294 );
and \U$43919 ( \44296 , \44291 , \44295 );
and \U$43920 ( \44297 , \44288 , \44290 );
or \U$43921 ( \44298 , \44296 , \44297 );
xor \U$43922 ( \44299 , \44286 , \44298 );
and \U$43923 ( \44300 , \384 , RIae77900_86);
and \U$43924 ( \44301 , RIae76fa0_66, \382 );
nor \U$43925 ( \44302 , \44300 , \44301 );
not \U$43926 ( \44303 , \44302 );
not \U$43927 ( \44304 , \388 );
and \U$43928 ( \44305 , \44303 , \44304 );
and \U$43929 ( \44306 , \44302 , \388 );
nor \U$43930 ( \44307 , \44305 , \44306 );
nand \U$43931 ( \44308 , RIae77810_84, RIae78b48_125);
or \U$43932 ( \44309 , \44307 , \44308 );
not \U$43933 ( \44310 , \44308 );
not \U$43934 ( \44311 , \44307 );
or \U$43935 ( \44312 , \44310 , \44311 );
not \U$43936 ( \44313 , \402 );
and \U$43937 ( \44314 , \436 , RIae76eb0_64);
and \U$43938 ( \44315 , RIae76dc0_62, \434 );
nor \U$43939 ( \44316 , \44314 , \44315 );
not \U$43940 ( \44317 , \44316 );
or \U$43941 ( \44318 , \44313 , \44317 );
or \U$43942 ( \44319 , \44316 , \400 );
nand \U$43943 ( \44320 , \44318 , \44319 );
nand \U$43944 ( \44321 , \44312 , \44320 );
nand \U$43945 ( \44322 , \44309 , \44321 );
xor \U$43946 ( \44323 , \43667 , \43669 );
xor \U$43947 ( \44324 , \44323 , \43678 );
and \U$43948 ( \44325 , \44322 , \44324 );
xor \U$43949 ( \44326 , \43764 , \43772 );
xor \U$43950 ( \44327 , \44326 , \43780 );
xor \U$43951 ( \44328 , \43667 , \43669 );
xor \U$43952 ( \44329 , \44328 , \43678 );
and \U$43953 ( \44330 , \44327 , \44329 );
and \U$43954 ( \44331 , \44322 , \44327 );
or \U$43955 ( \44332 , \44325 , \44330 , \44331 );
xor \U$43956 ( \44333 , \43712 , \43719 );
xor \U$43957 ( \44334 , \44333 , \43727 );
xor \U$43958 ( \44335 , \43737 , \43745 );
xor \U$43959 ( \44336 , \44335 , \43753 );
xor \U$43960 ( \44337 , \44334 , \44336 );
xor \U$43961 ( \44338 , \43917 , \43925 );
xor \U$43962 ( \44339 , \44338 , \43934 );
and \U$43963 ( \44340 , \44337 , \44339 );
and \U$43964 ( \44341 , \44334 , \44336 );
or \U$43965 ( \44342 , \44340 , \44341 );
xor \U$43966 ( \44343 , \44332 , \44342 );
xor \U$43967 ( \44344 , \43866 , \43873 );
xor \U$43968 ( \44345 , \44344 , \43881 );
xor \U$43969 ( \44346 , \43891 , \43898 );
xor \U$43970 ( \44347 , \44346 , \43906 );
and \U$43971 ( \44348 , \44345 , \44347 );
xor \U$43972 ( \44349 , \43793 , \43800 );
xor \U$43973 ( \44350 , \44349 , \43808 );
xor \U$43974 ( \44351 , \43891 , \43898 );
xor \U$43975 ( \44352 , \44351 , \43906 );
and \U$43976 ( \44353 , \44350 , \44352 );
and \U$43977 ( \44354 , \44345 , \44350 );
or \U$43978 ( \44355 , \44348 , \44353 , \44354 );
and \U$43979 ( \44356 , \44343 , \44355 );
and \U$43980 ( \44357 , \44332 , \44342 );
or \U$43981 ( \44358 , \44356 , \44357 );
and \U$43982 ( \44359 , \44299 , \44358 );
and \U$43983 ( \44360 , \44286 , \44298 );
or \U$43984 ( \44361 , \44359 , \44360 );
xor \U$43985 ( \44362 , \44043 , \44361 );
xor \U$43986 ( \44363 , \43730 , \43756 );
xor \U$43987 ( \44364 , \44363 , \43783 );
xor \U$43988 ( \44365 , \43681 , \43683 );
xor \U$43989 ( \44366 , \44365 , \43686 );
and \U$43990 ( \44367 , \44364 , \44366 );
xor \U$43991 ( \44368 , \43361 , \43369 );
xor \U$43992 ( \44369 , \44368 , \43377 );
xor \U$43993 ( \44370 , \43649 , \43654 );
xor \U$43994 ( \44371 , \44369 , \44370 );
xor \U$43995 ( \44372 , \43681 , \43683 );
xor \U$43996 ( \44373 , \44372 , \43686 );
and \U$43997 ( \44374 , \44371 , \44373 );
and \U$43998 ( \44375 , \44364 , \44371 );
or \U$43999 ( \44376 , \44367 , \44374 , \44375 );
xor \U$44000 ( \44377 , \43437 , \43460 );
xor \U$44001 ( \44378 , \44377 , \43486 );
xor \U$44002 ( \44379 , \44376 , \44378 );
xor \U$44003 ( \44380 , \43354 , \43380 );
xor \U$44004 ( \44381 , \44380 , \43408 );
xor \U$44005 ( \44382 , \43966 , \43971 );
xor \U$44006 ( \44383 , \44381 , \44382 );
and \U$44007 ( \44384 , \44379 , \44383 );
and \U$44008 ( \44385 , \44376 , \44378 );
or \U$44009 ( \44386 , \44384 , \44385 );
and \U$44010 ( \44387 , \44362 , \44386 );
and \U$44011 ( \44388 , \44043 , \44361 );
or \U$44012 ( \44389 , \44387 , \44388 );
xor \U$44013 ( \44390 , \43492 , \43514 );
xor \U$44014 ( \44391 , \44390 , \43565 );
xor \U$44015 ( \44392 , \44389 , \44391 );
xor \U$44016 ( \44393 , \43705 , \43943 );
xor \U$44017 ( \44394 , \44393 , \43960 );
xor \U$44018 ( \44395 , \43639 , \43641 );
xor \U$44019 ( \44396 , \44395 , \43644 );
and \U$44020 ( \44397 , \44394 , \44396 );
xor \U$44021 ( \44398 , \43220 , \43222 );
xor \U$44022 ( \44399 , \44398 , \43225 );
xor \U$44023 ( \44400 , \43976 , \43983 );
xor \U$44024 ( \44401 , \44399 , \44400 );
xor \U$44025 ( \44402 , \43639 , \43641 );
xor \U$44026 ( \44403 , \44402 , \43644 );
and \U$44027 ( \44404 , \44401 , \44403 );
and \U$44028 ( \44405 , \44394 , \44401 );
or \U$44029 ( \44406 , \44397 , \44404 , \44405 );
and \U$44030 ( \44407 , \44392 , \44406 );
and \U$44031 ( \44408 , \44389 , \44391 );
or \U$44032 ( \44409 , \44407 , \44408 );
and \U$44033 ( \44410 , \44029 , \44409 );
and \U$44034 ( \44411 , \44026 , \44028 );
or \U$44035 ( \44412 , \44410 , \44411 );
xor \U$44036 ( \44413 , \43588 , \43602 );
xor \U$44037 ( \44414 , \44413 , \43605 );
xor \U$44038 ( \44415 , \43618 , \43999 );
xor \U$44039 ( \44416 , \44414 , \44415 );
and \U$44040 ( \44417 , \44412 , \44416 );
and \U$44041 ( \44418 , \44019 , \44417 );
xor \U$44042 ( \44419 , \44417 , \44019 );
xor \U$44043 ( \44420 , \44412 , \44416 );
not \U$44044 ( \44421 , \44420 );
xor \U$44045 ( \44422 , \44286 , \44298 );
xor \U$44046 ( \44423 , \44422 , \44358 );
xor \U$44047 ( \44424 , \44376 , \44378 );
xor \U$44048 ( \44425 , \44424 , \44383 );
and \U$44049 ( \44426 , \44423 , \44425 );
xor \U$44050 ( \44427 , \43659 , \43689 );
xor \U$44051 ( \44428 , \44427 , \43702 );
xor \U$44052 ( \44429 , \44031 , \44038 );
xor \U$44053 ( \44430 , \44428 , \44429 );
xor \U$44054 ( \44431 , \44376 , \44378 );
xor \U$44055 ( \44432 , \44431 , \44383 );
and \U$44056 ( \44433 , \44430 , \44432 );
and \U$44057 ( \44434 , \44423 , \44430 );
or \U$44058 ( \44435 , \44426 , \44433 , \44434 );
xor \U$44059 ( \44436 , \43811 , \43829 );
xor \U$44060 ( \44437 , \44436 , \43855 );
xor \U$44061 ( \44438 , \44288 , \44290 );
xor \U$44062 ( \44439 , \44438 , \44295 );
and \U$44063 ( \44440 , \44437 , \44439 );
xor \U$44064 ( \44441 , \43681 , \43683 );
xor \U$44065 ( \44442 , \44441 , \43686 );
xor \U$44066 ( \44443 , \44364 , \44371 );
xor \U$44067 ( \44444 , \44442 , \44443 );
xor \U$44068 ( \44445 , \44288 , \44290 );
xor \U$44069 ( \44446 , \44445 , \44295 );
and \U$44070 ( \44447 , \44444 , \44446 );
and \U$44071 ( \44448 , \44437 , \44444 );
or \U$44072 ( \44449 , \44440 , \44447 , \44448 );
and \U$44073 ( \44450 , \5399 , RIae75650_12);
and \U$44074 ( \44451 , RIae75560_10, \5397 );
nor \U$44075 ( \44452 , \44450 , \44451 );
and \U$44076 ( \44453 , \44452 , \5016 );
not \U$44077 ( \44454 , \44452 );
and \U$44078 ( \44455 , \44454 , \5403 );
nor \U$44079 ( \44456 , \44453 , \44455 );
and \U$44080 ( \44457 , \4247 , RIae75fb0_32);
and \U$44081 ( \44458 , RIae75ec0_30, \4245 );
nor \U$44082 ( \44459 , \44457 , \44458 );
and \U$44083 ( \44460 , \44459 , \3989 );
not \U$44084 ( \44461 , \44459 );
and \U$44085 ( \44462 , \44461 , \4251 );
nor \U$44086 ( \44463 , \44460 , \44462 );
xor \U$44087 ( \44464 , \44456 , \44463 );
and \U$44088 ( \44465 , \4688 , RIae75ce0_26);
and \U$44089 ( \44466 , RIae75dd0_28, \4686 );
nor \U$44090 ( \44467 , \44465 , \44466 );
and \U$44091 ( \44468 , \44467 , \4481 );
not \U$44092 ( \44469 , \44467 );
and \U$44093 ( \44470 , \44469 , \4482 );
nor \U$44094 ( \44471 , \44468 , \44470 );
and \U$44095 ( \44472 , \44464 , \44471 );
and \U$44096 ( \44473 , \44456 , \44463 );
or \U$44097 ( \44474 , \44472 , \44473 );
and \U$44098 ( \44475 , \3730 , RIae75a10_20);
and \U$44099 ( \44476 , RIae75920_18, \3728 );
nor \U$44100 ( \44477 , \44475 , \44476 );
and \U$44101 ( \44478 , \44477 , \3732 );
not \U$44102 ( \44479 , \44477 );
and \U$44103 ( \44480 , \44479 , \3422 );
nor \U$44104 ( \44481 , \44478 , \44480 );
not \U$44105 ( \44482 , \2789 );
and \U$44106 ( \44483 , \2783 , RIae78800_118);
and \U$44107 ( \44484 , RIae78710_116, \2781 );
nor \U$44108 ( \44485 , \44483 , \44484 );
not \U$44109 ( \44486 , \44485 );
or \U$44110 ( \44487 , \44482 , \44486 );
or \U$44111 ( \44488 , \44485 , \3089 );
nand \U$44112 ( \44489 , \44487 , \44488 );
xor \U$44113 ( \44490 , \44481 , \44489 );
not \U$44114 ( \44491 , \3218 );
and \U$44115 ( \44492 , \3214 , RIae75bf0_24);
and \U$44116 ( \44493 , RIae75b00_22, \3212 );
nor \U$44117 ( \44494 , \44492 , \44493 );
not \U$44118 ( \44495 , \44494 );
or \U$44119 ( \44496 , \44491 , \44495 );
or \U$44120 ( \44497 , \44494 , \2774 );
nand \U$44121 ( \44498 , \44496 , \44497 );
and \U$44122 ( \44499 , \44490 , \44498 );
and \U$44123 ( \44500 , \44481 , \44489 );
or \U$44124 ( \44501 , \44499 , \44500 );
xor \U$44125 ( \44502 , \44474 , \44501 );
and \U$44126 ( \44503 , \5896 , RIae75830_16);
and \U$44127 ( \44504 , RIae75740_14, \5894 );
nor \U$44128 ( \44505 , \44503 , \44504 );
and \U$44129 ( \44506 , \44505 , \5590 );
not \U$44130 ( \44507 , \44505 );
and \U$44131 ( \44508 , \44507 , \5589 );
nor \U$44132 ( \44509 , \44506 , \44508 );
and \U$44133 ( \44510 , \6172 , RIae75290_4);
and \U$44134 ( \44511 , RIae751a0_2, \6170 );
nor \U$44135 ( \44512 , \44510 , \44511 );
and \U$44136 ( \44513 , \44512 , \6176 );
not \U$44137 ( \44514 , \44512 );
and \U$44138 ( \44515 , \44514 , \6175 );
nor \U$44139 ( \44516 , \44513 , \44515 );
xor \U$44140 ( \44517 , \44509 , \44516 );
and \U$44141 ( \44518 , \6941 , RIae75380_6);
and \U$44142 ( \44519 , RIae75470_8, \6939 );
nor \U$44143 ( \44520 , \44518 , \44519 );
and \U$44144 ( \44521 , \44520 , \6314 );
not \U$44145 ( \44522 , \44520 );
and \U$44146 ( \44523 , \44522 , \6945 );
nor \U$44147 ( \44524 , \44521 , \44523 );
and \U$44148 ( \44525 , \44517 , \44524 );
and \U$44149 ( \44526 , \44509 , \44516 );
or \U$44150 ( \44527 , \44525 , \44526 );
and \U$44151 ( \44528 , \44502 , \44527 );
and \U$44152 ( \44529 , \44474 , \44501 );
or \U$44153 ( \44530 , \44528 , \44529 );
and \U$44154 ( \44531 , \7633 , RIae76460_42);
and \U$44155 ( \44532 , RIae76550_44, \7631 );
nor \U$44156 ( \44533 , \44531 , \44532 );
and \U$44157 ( \44534 , \44533 , \7206 );
not \U$44158 ( \44535 , \44533 );
and \U$44159 ( \44536 , \44535 , \7205 );
nor \U$44160 ( \44537 , \44534 , \44536 );
and \U$44161 ( \44538 , \8371 , RIae76730_48);
and \U$44162 ( \44539 , RIae76640_46, \8369 );
nor \U$44163 ( \44540 , \44538 , \44539 );
and \U$44164 ( \44541 , \44540 , \8020 );
not \U$44165 ( \44542 , \44540 );
and \U$44166 ( \44543 , \44542 , \8019 );
nor \U$44167 ( \44544 , \44541 , \44543 );
xor \U$44168 ( \44545 , \44537 , \44544 );
and \U$44169 ( \44546 , \8966 , RIae76190_36);
and \U$44170 ( \44547 , RIae760a0_34, \8964 );
nor \U$44171 ( \44548 , \44546 , \44547 );
and \U$44172 ( \44549 , \44548 , \8799 );
not \U$44173 ( \44550 , \44548 );
and \U$44174 ( \44551 , \44550 , \8789 );
nor \U$44175 ( \44552 , \44549 , \44551 );
and \U$44176 ( \44553 , \44545 , \44552 );
and \U$44177 ( \44554 , \44537 , \44544 );
or \U$44178 ( \44555 , \44553 , \44554 );
and \U$44179 ( \44556 , \12180 , RIae76be0_58);
and \U$44180 ( \44557 , RIae78ad0_124, \12178 );
nor \U$44181 ( \44558 , \44556 , \44557 );
and \U$44182 ( \44559 , \44558 , \12184 );
not \U$44183 ( \44560 , \44558 );
and \U$44184 ( \44561 , \44560 , \11827 );
nor \U$44185 ( \44562 , \44559 , \44561 );
xor \U$44186 ( \44563 , \44562 , \13502 );
and \U$44187 ( \44564 , \13059 , RIae78d28_129);
and \U$44188 ( \44565 , RIae78e18_131, \13057 );
nor \U$44189 ( \44566 , \44564 , \44565 );
and \U$44190 ( \44567 , \44566 , \13063 );
not \U$44191 ( \44568 , \44566 );
and \U$44192 ( \44569 , \44568 , \12718 );
nor \U$44193 ( \44570 , \44567 , \44569 );
and \U$44194 ( \44571 , \44563 , \44570 );
and \U$44195 ( \44572 , \44562 , \13502 );
or \U$44196 ( \44573 , \44571 , \44572 );
xor \U$44197 ( \44574 , \44555 , \44573 );
and \U$44198 ( \44575 , \9760 , RIae76370_40);
and \U$44199 ( \44576 , RIae76280_38, \9758 );
nor \U$44200 ( \44577 , \44575 , \44576 );
and \U$44201 ( \44578 , \44577 , \9273 );
not \U$44202 ( \44579 , \44577 );
and \U$44203 ( \44580 , \44579 , \9764 );
nor \U$44204 ( \44581 , \44578 , \44580 );
and \U$44205 ( \44582 , \10548 , RIae76af0_56);
and \U$44206 ( \44583 , RIae76a00_54, \10546 );
nor \U$44207 ( \44584 , \44582 , \44583 );
and \U$44208 ( \44585 , \44584 , \10421 );
not \U$44209 ( \44586 , \44584 );
and \U$44210 ( \44587 , \44586 , \10118 );
nor \U$44211 ( \44588 , \44585 , \44587 );
xor \U$44212 ( \44589 , \44581 , \44588 );
and \U$44213 ( \44590 , \11470 , RIae76820_50);
and \U$44214 ( \44591 , RIae76910_52, \11468 );
nor \U$44215 ( \44592 , \44590 , \44591 );
and \U$44216 ( \44593 , \44592 , \10936 );
not \U$44217 ( \44594 , \44592 );
and \U$44218 ( \44595 , \44594 , \11474 );
nor \U$44219 ( \44596 , \44593 , \44595 );
and \U$44220 ( \44597 , \44589 , \44596 );
and \U$44221 ( \44598 , \44581 , \44588 );
or \U$44222 ( \44599 , \44597 , \44598 );
and \U$44223 ( \44600 , \44574 , \44599 );
and \U$44224 ( \44601 , \44555 , \44573 );
or \U$44225 ( \44602 , \44600 , \44601 );
xor \U$44226 ( \44603 , \44530 , \44602 );
and \U$44227 ( \44604 , \1138 , RIae77f90_100);
and \U$44228 ( \44605 , RIae78080_102, \1136 );
nor \U$44229 ( \44606 , \44604 , \44605 );
and \U$44230 ( \44607 , \44606 , \1012 );
not \U$44231 ( \44608 , \44606 );
and \U$44232 ( \44609 , \44608 , \1142 );
nor \U$44233 ( \44610 , \44607 , \44609 );
and \U$44234 ( \44611 , \1376 , RIae78260_106);
and \U$44235 ( \44612 , RIae78620_114, \1374 );
nor \U$44236 ( \44613 , \44611 , \44612 );
and \U$44237 ( \44614 , \44613 , \1380 );
not \U$44238 ( \44615 , \44613 );
and \U$44239 ( \44616 , \44615 , \1261 );
nor \U$44240 ( \44617 , \44614 , \44616 );
xor \U$44241 ( \44618 , \44610 , \44617 );
and \U$44242 ( \44619 , \1593 , RIae78440_110);
and \U$44243 ( \44620 , RIae784b8_111, \1591 );
nor \U$44244 ( \44621 , \44619 , \44620 );
and \U$44245 ( \44622 , \44621 , \1498 );
not \U$44246 ( \44623 , \44621 );
and \U$44247 ( \44624 , \44623 , \1488 );
nor \U$44248 ( \44625 , \44622 , \44624 );
and \U$44249 ( \44626 , \44618 , \44625 );
and \U$44250 ( \44627 , \44610 , \44617 );
or \U$44251 ( \44628 , \44626 , \44627 );
and \U$44252 ( \44629 , \558 , RIae77108_69);
and \U$44253 ( \44630 , RIae77090_68, \556 );
nor \U$44254 ( \44631 , \44629 , \44630 );
and \U$44255 ( \44632 , \44631 , \504 );
not \U$44256 ( \44633 , \44631 );
and \U$44257 ( \44634 , \44633 , \562 );
nor \U$44258 ( \44635 , \44632 , \44634 );
and \U$44259 ( \44636 , \672 , RIae77270_72);
and \U$44260 ( \44637 , RIae77360_74, \670 );
nor \U$44261 ( \44638 , \44636 , \44637 );
and \U$44262 ( \44639 , \44638 , \588 );
not \U$44263 ( \44640 , \44638 );
and \U$44264 ( \44641 , \44640 , \587 );
nor \U$44265 ( \44642 , \44639 , \44641 );
xor \U$44266 ( \44643 , \44635 , \44642 );
not \U$44267 ( \44644 , \787 );
and \U$44268 ( \44645 , \883 , RIae78350_108);
and \U$44269 ( \44646 , RIae78170_104, \881 );
nor \U$44270 ( \44647 , \44645 , \44646 );
not \U$44271 ( \44648 , \44647 );
or \U$44272 ( \44649 , \44644 , \44648 );
or \U$44273 ( \44650 , \44647 , \787 );
nand \U$44274 ( \44651 , \44649 , \44650 );
and \U$44275 ( \44652 , \44643 , \44651 );
and \U$44276 ( \44653 , \44635 , \44642 );
or \U$44277 ( \44654 , \44652 , \44653 );
xor \U$44278 ( \44655 , \44628 , \44654 );
and \U$44279 ( \44656 , \2224 , RIae77db0_96);
and \U$44280 ( \44657 , RIae77ea0_98, \2222 );
nor \U$44281 ( \44658 , \44656 , \44657 );
and \U$44282 ( \44659 , \44658 , \2061 );
not \U$44283 ( \44660 , \44658 );
and \U$44284 ( \44661 , \44660 , \2060 );
nor \U$44285 ( \44662 , \44659 , \44661 );
and \U$44286 ( \44663 , \1939 , RIae77cc0_94);
and \U$44287 ( \44664 , RIae77bd0_92, \1937 );
nor \U$44288 ( \44665 , \44663 , \44664 );
and \U$44289 ( \44666 , \44665 , \1735 );
not \U$44290 ( \44667 , \44665 );
and \U$44291 ( \44668 , \44667 , \1734 );
nor \U$44292 ( \44669 , \44666 , \44668 );
xor \U$44293 ( \44670 , \44662 , \44669 );
and \U$44294 ( \44671 , \2607 , RIae789e0_122);
and \U$44295 ( \44672 , RIae788f0_120, \2605 );
nor \U$44296 ( \44673 , \44671 , \44672 );
and \U$44297 ( \44674 , \44673 , \2611 );
not \U$44298 ( \44675 , \44673 );
and \U$44299 ( \44676 , \44675 , \2396 );
nor \U$44300 ( \44677 , \44674 , \44676 );
and \U$44301 ( \44678 , \44670 , \44677 );
and \U$44302 ( \44679 , \44662 , \44669 );
or \U$44303 ( \44680 , \44678 , \44679 );
and \U$44304 ( \44681 , \44655 , \44680 );
and \U$44305 ( \44682 , \44628 , \44654 );
or \U$44306 ( \44683 , \44681 , \44682 );
and \U$44307 ( \44684 , \44603 , \44683 );
and \U$44308 ( \44685 , \44530 , \44602 );
or \U$44309 ( \44686 , \44684 , \44685 );
xor \U$44310 ( \44687 , \43837 , \43844 );
xor \U$44311 ( \44688 , \44687 , \43852 );
xor \U$44312 ( \44689 , \43818 , \13063 );
xor \U$44313 ( \44690 , \44689 , \43826 );
xor \U$44314 ( \44691 , \44688 , \44690 );
xor \U$44315 ( \44692 , \44238 , \44243 );
xor \U$44316 ( \44693 , \44692 , \44251 );
xor \U$44317 ( \44694 , \44262 , \44269 );
xor \U$44318 ( \44695 , \44694 , \44277 );
and \U$44319 ( \44696 , \44693 , \44695 );
xor \U$44320 ( \44697 , \44213 , \44220 );
xor \U$44321 ( \44698 , \44697 , \44228 );
xor \U$44322 ( \44699 , \44262 , \44269 );
xor \U$44323 ( \44700 , \44699 , \44277 );
and \U$44324 ( \44701 , \44698 , \44700 );
and \U$44325 ( \44702 , \44693 , \44698 );
or \U$44326 ( \44703 , \44696 , \44701 , \44702 );
and \U$44327 ( \44704 , \44691 , \44703 );
and \U$44328 ( \44705 , \44688 , \44690 );
or \U$44329 ( \44706 , \44704 , \44705 );
xor \U$44330 ( \44707 , \44686 , \44706 );
xor \U$44331 ( \44708 , \44103 , \44110 );
xor \U$44332 ( \44709 , \44708 , \44118 );
xor \U$44333 ( \44710 , \44076 , \44083 );
xor \U$44334 ( \44711 , \44710 , \44092 );
xor \U$44335 ( \44712 , \44709 , \44711 );
xor \U$44336 ( \44713 , \44050 , \44057 );
xor \U$44337 ( \44714 , \44713 , \44065 );
and \U$44338 ( \44715 , \44712 , \44714 );
and \U$44339 ( \44716 , \44709 , \44711 );
or \U$44340 ( \44717 , \44715 , \44716 );
and \U$44341 ( \44718 , \384 , RIae77810_84);
and \U$44342 ( \44719 , RIae77900_86, \382 );
nor \U$44343 ( \44720 , \44718 , \44719 );
not \U$44344 ( \44721 , \44720 );
not \U$44345 ( \44722 , \388 );
and \U$44346 ( \44723 , \44721 , \44722 );
and \U$44347 ( \44724 , \44720 , \388 );
nor \U$44348 ( \44725 , \44723 , \44724 );
not \U$44349 ( \44726 , \44725 );
and \U$44350 ( \44727 , \436 , RIae76fa0_66);
and \U$44351 ( \44728 , RIae76eb0_64, \434 );
nor \U$44352 ( \44729 , \44727 , \44728 );
not \U$44353 ( \44730 , \44729 );
not \U$44354 ( \44731 , \402 );
and \U$44355 ( \44732 , \44730 , \44731 );
and \U$44356 ( \44733 , \44729 , \400 );
nor \U$44357 ( \44734 , \44732 , \44733 );
not \U$44358 ( \44735 , \44734 );
and \U$44359 ( \44736 , \44726 , \44735 );
and \U$44360 ( \44737 , \44734 , \44725 );
and \U$44361 ( \44738 , \514 , RIae76dc0_62);
and \U$44362 ( \44739 , RIae76cd0_60, \512 );
nor \U$44363 ( \44740 , \44738 , \44739 );
not \U$44364 ( \44741 , \44740 );
not \U$44365 ( \44742 , \471 );
and \U$44366 ( \44743 , \44741 , \44742 );
and \U$44367 ( \44744 , \44740 , \469 );
nor \U$44368 ( \44745 , \44743 , \44744 );
nor \U$44369 ( \44746 , \44737 , \44745 );
nor \U$44370 ( \44747 , \44736 , \44746 );
not \U$44371 ( \44748 , \44307 );
not \U$44372 ( \44749 , \44320 );
or \U$44373 ( \44750 , \44748 , \44749 );
or \U$44374 ( \44751 , \44307 , \44320 );
nand \U$44375 ( \44752 , \44750 , \44751 );
not \U$44376 ( \44753 , \44752 );
not \U$44377 ( \44754 , \44308 );
and \U$44378 ( \44755 , \44753 , \44754 );
and \U$44379 ( \44756 , \44752 , \44308 );
nor \U$44380 ( \44757 , \44755 , \44756 );
nand \U$44381 ( \44758 , \44747 , \44757 );
xor \U$44382 ( \44759 , \44717 , \44758 );
xor \U$44383 ( \44760 , \44132 , \44139 );
xor \U$44384 ( \44761 , \44760 , \44147 );
xor \U$44385 ( \44762 , \44157 , \44165 );
xor \U$44386 ( \44763 , \44762 , \44173 );
and \U$44387 ( \44764 , \44761 , \44763 );
xor \U$44388 ( \44765 , \44184 , \44191 );
xor \U$44389 ( \44766 , \44765 , \44199 );
xor \U$44390 ( \44767 , \44157 , \44165 );
xor \U$44391 ( \44768 , \44767 , \44173 );
and \U$44392 ( \44769 , \44766 , \44768 );
and \U$44393 ( \44770 , \44761 , \44766 );
or \U$44394 ( \44771 , \44764 , \44769 , \44770 );
and \U$44395 ( \44772 , \44759 , \44771 );
and \U$44396 ( \44773 , \44717 , \44758 );
or \U$44397 ( \44774 , \44772 , \44773 );
and \U$44398 ( \44775 , \44707 , \44774 );
and \U$44399 ( \44776 , \44686 , \44706 );
or \U$44400 ( \44777 , \44775 , \44776 );
xor \U$44401 ( \44778 , \44449 , \44777 );
xor \U$44402 ( \44779 , \44231 , \44254 );
xor \U$44403 ( \44780 , \44779 , \44280 );
xor \U$44404 ( \44781 , \44150 , \44176 );
xor \U$44405 ( \44782 , \44781 , \44202 );
and \U$44406 ( \44783 , \44780 , \44782 );
xor \U$44407 ( \44784 , \44068 , \44095 );
xor \U$44408 ( \44785 , \44784 , \44121 );
xor \U$44409 ( \44786 , \44150 , \44176 );
xor \U$44410 ( \44787 , \44786 , \44202 );
and \U$44411 ( \44788 , \44785 , \44787 );
and \U$44412 ( \44789 , \44780 , \44785 );
or \U$44413 ( \44790 , \44783 , \44788 , \44789 );
xor \U$44414 ( \44791 , \43884 , \43909 );
xor \U$44415 ( \44792 , \44791 , \43937 );
xor \U$44416 ( \44793 , \44790 , \44792 );
xor \U$44417 ( \44794 , \43667 , \43669 );
xor \U$44418 ( \44795 , \44794 , \43678 );
xor \U$44419 ( \44796 , \44322 , \44327 );
xor \U$44420 ( \44797 , \44795 , \44796 );
xor \U$44421 ( \44798 , \44334 , \44336 );
xor \U$44422 ( \44799 , \44798 , \44339 );
and \U$44423 ( \44800 , \44797 , \44799 );
xor \U$44424 ( \44801 , \43891 , \43898 );
xor \U$44425 ( \44802 , \44801 , \43906 );
xor \U$44426 ( \44803 , \44345 , \44350 );
xor \U$44427 ( \44804 , \44802 , \44803 );
xor \U$44428 ( \44805 , \44334 , \44336 );
xor \U$44429 ( \44806 , \44805 , \44339 );
and \U$44430 ( \44807 , \44804 , \44806 );
and \U$44431 ( \44808 , \44797 , \44804 );
or \U$44432 ( \44809 , \44800 , \44807 , \44808 );
and \U$44433 ( \44810 , \44793 , \44809 );
and \U$44434 ( \44811 , \44790 , \44792 );
or \U$44435 ( \44812 , \44810 , \44811 );
and \U$44436 ( \44813 , \44778 , \44812 );
and \U$44437 ( \44814 , \44449 , \44777 );
or \U$44438 ( \44815 , \44813 , \44814 );
xor \U$44439 ( \44816 , \44435 , \44815 );
xor \U$44440 ( \44817 , \43639 , \43641 );
xor \U$44441 ( \44818 , \44817 , \43644 );
xor \U$44442 ( \44819 , \44394 , \44401 );
xor \U$44443 ( \44820 , \44818 , \44819 );
and \U$44444 ( \44821 , \44816 , \44820 );
and \U$44445 ( \44822 , \44435 , \44815 );
or \U$44446 ( \44823 , \44821 , \44822 );
xor \U$44447 ( \44824 , \44021 , \44025 );
xor \U$44448 ( \44825 , \44823 , \44824 );
xor \U$44449 ( \44826 , \44389 , \44391 );
xor \U$44450 ( \44827 , \44826 , \44406 );
and \U$44451 ( \44828 , \44825 , \44827 );
and \U$44452 ( \44829 , \44823 , \44824 );
or \U$44453 ( \44830 , \44828 , \44829 );
xor \U$44454 ( \44831 , \43635 , \43991 );
xor \U$44455 ( \44832 , \44831 , \43996 );
xor \U$44456 ( \44833 , \44830 , \44832 );
xor \U$44457 ( \44834 , \44026 , \44028 );
xor \U$44458 ( \44835 , \44834 , \44409 );
and \U$44459 ( \44836 , \44833 , \44835 );
and \U$44460 ( \44837 , \44830 , \44832 );
or \U$44461 ( \44838 , \44836 , \44837 );
not \U$44462 ( \44839 , \44838 );
or \U$44463 ( \44840 , \44421 , \44839 );
xor \U$44464 ( \44841 , \44830 , \44832 );
xor \U$44465 ( \44842 , \44841 , \44835 );
xor \U$44466 ( \44843 , \44530 , \44602 );
xor \U$44467 ( \44844 , \44843 , \44683 );
xor \U$44468 ( \44845 , \44688 , \44690 );
xor \U$44469 ( \44846 , \44845 , \44703 );
and \U$44470 ( \44847 , \44844 , \44846 );
xor \U$44471 ( \44848 , \44717 , \44758 );
xor \U$44472 ( \44849 , \44848 , \44771 );
xor \U$44473 ( \44850 , \44688 , \44690 );
xor \U$44474 ( \44851 , \44850 , \44703 );
and \U$44475 ( \44852 , \44849 , \44851 );
and \U$44476 ( \44853 , \44844 , \44849 );
or \U$44477 ( \44854 , \44847 , \44852 , \44853 );
xor \U$44478 ( \44855 , \44456 , \44463 );
xor \U$44479 ( \44856 , \44855 , \44471 );
xor \U$44480 ( \44857 , \44662 , \44669 );
xor \U$44481 ( \44858 , \44857 , \44677 );
xor \U$44482 ( \44859 , \44856 , \44858 );
xor \U$44483 ( \44860 , \44481 , \44489 );
xor \U$44484 ( \44861 , \44860 , \44498 );
and \U$44485 ( \44862 , \44859 , \44861 );
and \U$44486 ( \44863 , \44856 , \44858 );
or \U$44487 ( \44864 , \44862 , \44863 );
nand \U$44488 ( \44865 , RIae77ae0_90, RIae78b48_125);
not \U$44489 ( \44866 , \44865 );
not \U$44490 ( \44867 , RIae779f0_88);
nor \U$44491 ( \44868 , \44867 , \491 );
xor \U$44492 ( \44869 , \44866 , \44868 );
not \U$44493 ( \44870 , \402 );
and \U$44494 ( \44871 , \436 , RIae77900_86);
and \U$44495 ( \44872 , RIae76fa0_66, \434 );
nor \U$44496 ( \44873 , \44871 , \44872 );
not \U$44497 ( \44874 , \44873 );
or \U$44498 ( \44875 , \44870 , \44874 );
or \U$44499 ( \44876 , \44873 , \402 );
nand \U$44500 ( \44877 , \44875 , \44876 );
not \U$44501 ( \44878 , \388 );
and \U$44502 ( \44879 , \384 , RIae779f0_88);
and \U$44503 ( \44880 , RIae77810_84, \382 );
nor \U$44504 ( \44881 , \44879 , \44880 );
not \U$44505 ( \44882 , \44881 );
or \U$44506 ( \44883 , \44878 , \44882 );
or \U$44507 ( \44884 , \44881 , \392 );
nand \U$44508 ( \44885 , \44883 , \44884 );
xor \U$44509 ( \44886 , \44877 , \44885 );
not \U$44510 ( \44887 , \471 );
and \U$44511 ( \44888 , \514 , RIae76eb0_64);
and \U$44512 ( \44889 , RIae76dc0_62, \512 );
nor \U$44513 ( \44890 , \44888 , \44889 );
not \U$44514 ( \44891 , \44890 );
or \U$44515 ( \44892 , \44887 , \44891 );
or \U$44516 ( \44893 , \44890 , \469 );
nand \U$44517 ( \44894 , \44892 , \44893 );
and \U$44518 ( \44895 , \44886 , \44894 );
and \U$44519 ( \44896 , \44877 , \44885 );
or \U$44520 ( \44897 , \44895 , \44896 );
and \U$44521 ( \44898 , \44869 , \44897 );
and \U$44522 ( \44899 , \44866 , \44868 );
or \U$44523 ( \44900 , \44898 , \44899 );
xor \U$44524 ( \44901 , \44864 , \44900 );
not \U$44525 ( \44902 , \44725 );
xor \U$44526 ( \44903 , \44734 , \44745 );
not \U$44527 ( \44904 , \44903 );
or \U$44528 ( \44905 , \44902 , \44904 );
or \U$44529 ( \44906 , \44903 , \44725 );
nand \U$44530 ( \44907 , \44905 , \44906 );
xor \U$44531 ( \44908 , \44635 , \44642 );
xor \U$44532 ( \44909 , \44908 , \44651 );
and \U$44533 ( \44910 , \44907 , \44909 );
xor \U$44534 ( \44911 , \44610 , \44617 );
xor \U$44535 ( \44912 , \44911 , \44625 );
xor \U$44536 ( \44913 , \44635 , \44642 );
xor \U$44537 ( \44914 , \44913 , \44651 );
and \U$44538 ( \44915 , \44912 , \44914 );
and \U$44539 ( \44916 , \44907 , \44912 );
or \U$44540 ( \44917 , \44910 , \44915 , \44916 );
and \U$44541 ( \44918 , \44901 , \44917 );
and \U$44542 ( \44919 , \44864 , \44900 );
or \U$44543 ( \44920 , \44918 , \44919 );
and \U$44544 ( \44921 , \2224 , RIae77bd0_92);
and \U$44545 ( \44922 , RIae77db0_96, \2222 );
nor \U$44546 ( \44923 , \44921 , \44922 );
and \U$44547 ( \44924 , \44923 , \2061 );
not \U$44548 ( \44925 , \44923 );
and \U$44549 ( \44926 , \44925 , \2060 );
nor \U$44550 ( \44927 , \44924 , \44926 );
and \U$44551 ( \44928 , \1939 , RIae784b8_111);
and \U$44552 ( \44929 , RIae77cc0_94, \1937 );
nor \U$44553 ( \44930 , \44928 , \44929 );
and \U$44554 ( \44931 , \44930 , \1735 );
not \U$44555 ( \44932 , \44930 );
and \U$44556 ( \44933 , \44932 , \1734 );
nor \U$44557 ( \44934 , \44931 , \44933 );
xor \U$44558 ( \44935 , \44927 , \44934 );
and \U$44559 ( \44936 , \2607 , RIae77ea0_98);
and \U$44560 ( \44937 , RIae789e0_122, \2605 );
nor \U$44561 ( \44938 , \44936 , \44937 );
and \U$44562 ( \44939 , \44938 , \2611 );
not \U$44563 ( \44940 , \44938 );
and \U$44564 ( \44941 , \44940 , \2397 );
nor \U$44565 ( \44942 , \44939 , \44941 );
and \U$44566 ( \44943 , \44935 , \44942 );
and \U$44567 ( \44944 , \44927 , \44934 );
or \U$44568 ( \44945 , \44943 , \44944 );
and \U$44569 ( \44946 , \1138 , RIae78170_104);
and \U$44570 ( \44947 , RIae77f90_100, \1136 );
nor \U$44571 ( \44948 , \44946 , \44947 );
and \U$44572 ( \44949 , \44948 , \1012 );
not \U$44573 ( \44950 , \44948 );
and \U$44574 ( \44951 , \44950 , \1142 );
nor \U$44575 ( \44952 , \44949 , \44951 );
and \U$44576 ( \44953 , \1376 , RIae78080_102);
and \U$44577 ( \44954 , RIae78260_106, \1374 );
nor \U$44578 ( \44955 , \44953 , \44954 );
and \U$44579 ( \44956 , \44955 , \1380 );
not \U$44580 ( \44957 , \44955 );
and \U$44581 ( \44958 , \44957 , \1261 );
nor \U$44582 ( \44959 , \44956 , \44958 );
xor \U$44583 ( \44960 , \44952 , \44959 );
and \U$44584 ( \44961 , \1593 , RIae78620_114);
and \U$44585 ( \44962 , RIae78440_110, \1591 );
nor \U$44586 ( \44963 , \44961 , \44962 );
and \U$44587 ( \44964 , \44963 , \1498 );
not \U$44588 ( \44965 , \44963 );
and \U$44589 ( \44966 , \44965 , \1488 );
nor \U$44590 ( \44967 , \44964 , \44966 );
and \U$44591 ( \44968 , \44960 , \44967 );
and \U$44592 ( \44969 , \44952 , \44959 );
or \U$44593 ( \44970 , \44968 , \44969 );
xor \U$44594 ( \44971 , \44945 , \44970 );
and \U$44595 ( \44972 , \672 , RIae77090_68);
and \U$44596 ( \44973 , RIae77270_72, \670 );
nor \U$44597 ( \44974 , \44972 , \44973 );
and \U$44598 ( \44975 , \44974 , \588 );
not \U$44599 ( \44976 , \44974 );
and \U$44600 ( \44977 , \44976 , \587 );
nor \U$44601 ( \44978 , \44975 , \44977 );
and \U$44602 ( \44979 , \558 , RIae76cd0_60);
and \U$44603 ( \44980 , RIae77108_69, \556 );
nor \U$44604 ( \44981 , \44979 , \44980 );
and \U$44605 ( \44982 , \44981 , \504 );
not \U$44606 ( \44983 , \44981 );
and \U$44607 ( \44984 , \44983 , \562 );
nor \U$44608 ( \44985 , \44982 , \44984 );
xor \U$44609 ( \44986 , \44978 , \44985 );
not \U$44610 ( \44987 , \789 );
and \U$44611 ( \44988 , \883 , RIae77360_74);
and \U$44612 ( \44989 , RIae78350_108, \881 );
nor \U$44613 ( \44990 , \44988 , \44989 );
not \U$44614 ( \44991 , \44990 );
or \U$44615 ( \44992 , \44987 , \44991 );
or \U$44616 ( \44993 , \44990 , \787 );
nand \U$44617 ( \44994 , \44992 , \44993 );
and \U$44618 ( \44995 , \44986 , \44994 );
and \U$44619 ( \44996 , \44978 , \44985 );
or \U$44620 ( \44997 , \44995 , \44996 );
and \U$44621 ( \44998 , \44971 , \44997 );
and \U$44622 ( \44999 , \44945 , \44970 );
or \U$44623 ( \45000 , \44998 , \44999 );
and \U$44624 ( \45001 , \9760 , RIae760a0_34);
and \U$44625 ( \45002 , RIae76370_40, \9758 );
nor \U$44626 ( \45003 , \45001 , \45002 );
and \U$44627 ( \45004 , \45003 , \9273 );
not \U$44628 ( \45005 , \45003 );
and \U$44629 ( \45006 , \45005 , \9272 );
nor \U$44630 ( \45007 , \45004 , \45006 );
and \U$44631 ( \45008 , \10548 , RIae76280_38);
and \U$44632 ( \45009 , RIae76af0_56, \10546 );
nor \U$44633 ( \45010 , \45008 , \45009 );
and \U$44634 ( \45011 , \45010 , \10421 );
not \U$44635 ( \45012 , \45010 );
and \U$44636 ( \45013 , \45012 , \10118 );
nor \U$44637 ( \45014 , \45011 , \45013 );
xor \U$44638 ( \45015 , \45007 , \45014 );
and \U$44639 ( \45016 , \11470 , RIae76a00_54);
and \U$44640 ( \45017 , RIae76820_50, \11468 );
nor \U$44641 ( \45018 , \45016 , \45017 );
and \U$44642 ( \45019 , \45018 , \10936 );
not \U$44643 ( \45020 , \45018 );
and \U$44644 ( \45021 , \45020 , \11474 );
nor \U$44645 ( \45022 , \45019 , \45021 );
and \U$44646 ( \45023 , \45015 , \45022 );
and \U$44647 ( \45024 , \45007 , \45014 );
or \U$44648 ( \45025 , \45023 , \45024 );
and \U$44649 ( \45026 , \12180 , RIae76910_52);
and \U$44650 ( \45027 , RIae76be0_58, \12178 );
nor \U$44651 ( \45028 , \45026 , \45027 );
and \U$44652 ( \45029 , \45028 , \12184 );
not \U$44653 ( \45030 , \45028 );
and \U$44654 ( \45031 , \45030 , \11827 );
nor \U$44655 ( \45032 , \45029 , \45031 );
nand \U$44656 ( \45033 , RIae78e18_131, \14059 );
and \U$44657 ( \45034 , \45033 , \13502 );
not \U$44658 ( \45035 , \45033 );
and \U$44659 ( \45036 , \45035 , \14063 );
nor \U$44660 ( \45037 , \45034 , \45036 );
xor \U$44661 ( \45038 , \45032 , \45037 );
and \U$44662 ( \45039 , \13059 , RIae78ad0_124);
and \U$44663 ( \45040 , RIae78d28_129, \13057 );
nor \U$44664 ( \45041 , \45039 , \45040 );
and \U$44665 ( \45042 , \45041 , \13063 );
not \U$44666 ( \45043 , \45041 );
and \U$44667 ( \45044 , \45043 , \12718 );
nor \U$44668 ( \45045 , \45042 , \45044 );
and \U$44669 ( \45046 , \45038 , \45045 );
and \U$44670 ( \45047 , \45032 , \45037 );
or \U$44671 ( \45048 , \45046 , \45047 );
xor \U$44672 ( \45049 , \45025 , \45048 );
and \U$44673 ( \45050 , \8371 , RIae76550_44);
and \U$44674 ( \45051 , RIae76730_48, \8369 );
nor \U$44675 ( \45052 , \45050 , \45051 );
and \U$44676 ( \45053 , \45052 , \8020 );
not \U$44677 ( \45054 , \45052 );
and \U$44678 ( \45055 , \45054 , \8019 );
nor \U$44679 ( \45056 , \45053 , \45055 );
and \U$44680 ( \45057 , \7633 , RIae75470_8);
and \U$44681 ( \45058 , RIae76460_42, \7631 );
nor \U$44682 ( \45059 , \45057 , \45058 );
and \U$44683 ( \45060 , \45059 , \7206 );
not \U$44684 ( \45061 , \45059 );
and \U$44685 ( \45062 , \45061 , \7205 );
nor \U$44686 ( \45063 , \45060 , \45062 );
xor \U$44687 ( \45064 , \45056 , \45063 );
and \U$44688 ( \45065 , \8966 , RIae76640_46);
and \U$44689 ( \45066 , RIae76190_36, \8964 );
nor \U$44690 ( \45067 , \45065 , \45066 );
and \U$44691 ( \45068 , \45067 , \8799 );
not \U$44692 ( \45069 , \45067 );
and \U$44693 ( \45070 , \45069 , \8789 );
nor \U$44694 ( \45071 , \45068 , \45070 );
and \U$44695 ( \45072 , \45064 , \45071 );
and \U$44696 ( \45073 , \45056 , \45063 );
or \U$44697 ( \45074 , \45072 , \45073 );
and \U$44698 ( \45075 , \45049 , \45074 );
and \U$44699 ( \45076 , \45025 , \45048 );
or \U$44700 ( \45077 , \45075 , \45076 );
xor \U$44701 ( \45078 , \45000 , \45077 );
and \U$44702 ( \45079 , \4247 , RIae75920_18);
and \U$44703 ( \45080 , RIae75fb0_32, \4245 );
nor \U$44704 ( \45081 , \45079 , \45080 );
and \U$44705 ( \45082 , \45081 , \3989 );
not \U$44706 ( \45083 , \45081 );
and \U$44707 ( \45084 , \45083 , \4251 );
nor \U$44708 ( \45085 , \45082 , \45084 );
and \U$44709 ( \45086 , \4688 , RIae75ec0_30);
and \U$44710 ( \45087 , RIae75ce0_26, \4686 );
nor \U$44711 ( \45088 , \45086 , \45087 );
and \U$44712 ( \45089 , \45088 , \4481 );
not \U$44713 ( \45090 , \45088 );
and \U$44714 ( \45091 , \45090 , \4482 );
nor \U$44715 ( \45092 , \45089 , \45091 );
xor \U$44716 ( \45093 , \45085 , \45092 );
and \U$44717 ( \45094 , \5399 , RIae75dd0_28);
and \U$44718 ( \45095 , RIae75650_12, \5397 );
nor \U$44719 ( \45096 , \45094 , \45095 );
and \U$44720 ( \45097 , \45096 , \5016 );
not \U$44721 ( \45098 , \45096 );
and \U$44722 ( \45099 , \45098 , \5403 );
nor \U$44723 ( \45100 , \45097 , \45099 );
and \U$44724 ( \45101 , \45093 , \45100 );
and \U$44725 ( \45102 , \45085 , \45092 );
or \U$44726 ( \45103 , \45101 , \45102 );
not \U$44727 ( \45104 , \3089 );
and \U$44728 ( \45105 , \2783 , RIae788f0_120);
and \U$44729 ( \45106 , RIae78800_118, \2781 );
nor \U$44730 ( \45107 , \45105 , \45106 );
not \U$44731 ( \45108 , \45107 );
or \U$44732 ( \45109 , \45104 , \45108 );
or \U$44733 ( \45110 , \45107 , \3089 );
nand \U$44734 ( \45111 , \45109 , \45110 );
not \U$44735 ( \45112 , \3218 );
and \U$44736 ( \45113 , \3214 , RIae78710_116);
and \U$44737 ( \45114 , RIae75bf0_24, \3212 );
nor \U$44738 ( \45115 , \45113 , \45114 );
not \U$44739 ( \45116 , \45115 );
or \U$44740 ( \45117 , \45112 , \45116 );
or \U$44741 ( \45118 , \45115 , \3218 );
nand \U$44742 ( \45119 , \45117 , \45118 );
xor \U$44743 ( \45120 , \45111 , \45119 );
and \U$44744 ( \45121 , \3730 , RIae75b00_22);
and \U$44745 ( \45122 , RIae75a10_20, \3728 );
nor \U$44746 ( \45123 , \45121 , \45122 );
and \U$44747 ( \45124 , \45123 , \3732 );
not \U$44748 ( \45125 , \45123 );
and \U$44749 ( \45126 , \45125 , \3422 );
nor \U$44750 ( \45127 , \45124 , \45126 );
and \U$44751 ( \45128 , \45120 , \45127 );
and \U$44752 ( \45129 , \45111 , \45119 );
or \U$44753 ( \45130 , \45128 , \45129 );
xor \U$44754 ( \45131 , \45103 , \45130 );
and \U$44755 ( \45132 , \6172 , RIae75740_14);
and \U$44756 ( \45133 , RIae75290_4, \6170 );
nor \U$44757 ( \45134 , \45132 , \45133 );
and \U$44758 ( \45135 , \45134 , \6176 );
not \U$44759 ( \45136 , \45134 );
and \U$44760 ( \45137 , \45136 , \6175 );
nor \U$44761 ( \45138 , \45135 , \45137 );
and \U$44762 ( \45139 , \5896 , RIae75560_10);
and \U$44763 ( \45140 , RIae75830_16, \5894 );
nor \U$44764 ( \45141 , \45139 , \45140 );
and \U$44765 ( \45142 , \45141 , \5590 );
not \U$44766 ( \45143 , \45141 );
and \U$44767 ( \45144 , \45143 , \5589 );
nor \U$44768 ( \45145 , \45142 , \45144 );
xor \U$44769 ( \45146 , \45138 , \45145 );
and \U$44770 ( \45147 , \6941 , RIae751a0_2);
and \U$44771 ( \45148 , RIae75380_6, \6939 );
nor \U$44772 ( \45149 , \45147 , \45148 );
and \U$44773 ( \45150 , \45149 , \6314 );
not \U$44774 ( \45151 , \45149 );
and \U$44775 ( \45152 , \45151 , \6945 );
nor \U$44776 ( \45153 , \45150 , \45152 );
and \U$44777 ( \45154 , \45146 , \45153 );
and \U$44778 ( \45155 , \45138 , \45145 );
or \U$44779 ( \45156 , \45154 , \45155 );
and \U$44780 ( \45157 , \45131 , \45156 );
and \U$44781 ( \45158 , \45103 , \45130 );
or \U$44782 ( \45159 , \45157 , \45158 );
and \U$44783 ( \45160 , \45078 , \45159 );
and \U$44784 ( \45161 , \45000 , \45077 );
or \U$44785 ( \45162 , \45160 , \45161 );
xor \U$44786 ( \45163 , \44920 , \45162 );
xor \U$44787 ( \45164 , \44537 , \44544 );
xor \U$44788 ( \45165 , \45164 , \44552 );
xor \U$44789 ( \45166 , \44509 , \44516 );
xor \U$44790 ( \45167 , \45166 , \44524 );
and \U$44791 ( \45168 , \45165 , \45167 );
xor \U$44792 ( \45169 , \44581 , \44588 );
xor \U$44793 ( \45170 , \45169 , \44596 );
xor \U$44794 ( \45171 , \44509 , \44516 );
xor \U$44795 ( \45172 , \45171 , \44524 );
and \U$44796 ( \45173 , \45170 , \45172 );
and \U$44797 ( \45174 , \45165 , \45170 );
or \U$44798 ( \45175 , \45168 , \45173 , \45174 );
xor \U$44799 ( \45176 , \44709 , \44711 );
xor \U$44800 ( \45177 , \45176 , \44714 );
and \U$44801 ( \45178 , \45175 , \45177 );
xor \U$44802 ( \45179 , \44262 , \44269 );
xor \U$44803 ( \45180 , \45179 , \44277 );
xor \U$44804 ( \45181 , \44693 , \44698 );
xor \U$44805 ( \45182 , \45180 , \45181 );
xor \U$44806 ( \45183 , \44709 , \44711 );
xor \U$44807 ( \45184 , \45183 , \44714 );
and \U$44808 ( \45185 , \45182 , \45184 );
and \U$44809 ( \45186 , \45175 , \45182 );
or \U$44810 ( \45187 , \45178 , \45185 , \45186 );
and \U$44811 ( \45188 , \45163 , \45187 );
and \U$44812 ( \45189 , \44920 , \45162 );
or \U$44813 ( \45190 , \45188 , \45189 );
xor \U$44814 ( \45191 , \44854 , \45190 );
xor \U$44815 ( \45192 , \44150 , \44176 );
xor \U$44816 ( \45193 , \45192 , \44202 );
xor \U$44817 ( \45194 , \44780 , \44785 );
xor \U$44818 ( \45195 , \45193 , \45194 );
xor \U$44819 ( \45196 , \44628 , \44654 );
xor \U$44820 ( \45197 , \45196 , \44680 );
or \U$44821 ( \45198 , \44757 , \44747 );
nand \U$44822 ( \45199 , \45198 , \44758 );
xor \U$44823 ( \45200 , \45197 , \45199 );
xor \U$44824 ( \45201 , \44157 , \44165 );
xor \U$44825 ( \45202 , \45201 , \44173 );
xor \U$44826 ( \45203 , \44761 , \44766 );
xor \U$44827 ( \45204 , \45202 , \45203 );
and \U$44828 ( \45205 , \45200 , \45204 );
and \U$44829 ( \45206 , \45197 , \45199 );
or \U$44830 ( \45207 , \45205 , \45206 );
xor \U$44831 ( \45208 , \45195 , \45207 );
xor \U$44832 ( \45209 , \44334 , \44336 );
xor \U$44833 ( \45210 , \45209 , \44339 );
xor \U$44834 ( \45211 , \44797 , \44804 );
xor \U$44835 ( \45212 , \45210 , \45211 );
and \U$44836 ( \45213 , \45208 , \45212 );
and \U$44837 ( \45214 , \45195 , \45207 );
or \U$44838 ( \45215 , \45213 , \45214 );
and \U$44839 ( \45216 , \45191 , \45215 );
and \U$44840 ( \45217 , \44854 , \45190 );
or \U$44841 ( \45218 , \45216 , \45217 );
xor \U$44842 ( \45219 , \44332 , \44342 );
xor \U$44843 ( \45220 , \45219 , \44355 );
xor \U$44844 ( \45221 , \44124 , \44205 );
xor \U$44845 ( \45222 , \45221 , \44283 );
xor \U$44846 ( \45223 , \45220 , \45222 );
xor \U$44847 ( \45224 , \44288 , \44290 );
xor \U$44848 ( \45225 , \45224 , \44295 );
xor \U$44849 ( \45226 , \44437 , \44444 );
xor \U$44850 ( \45227 , \45225 , \45226 );
and \U$44851 ( \45228 , \45223 , \45227 );
and \U$44852 ( \45229 , \45220 , \45222 );
or \U$44853 ( \45230 , \45228 , \45229 );
xor \U$44854 ( \45231 , \45218 , \45230 );
xor \U$44855 ( \45232 , \44376 , \44378 );
xor \U$44856 ( \45233 , \45232 , \44383 );
xor \U$44857 ( \45234 , \44423 , \44430 );
xor \U$44858 ( \45235 , \45233 , \45234 );
and \U$44859 ( \45236 , \45231 , \45235 );
and \U$44860 ( \45237 , \45218 , \45230 );
or \U$44861 ( \45238 , \45236 , \45237 );
xor \U$44862 ( \45239 , \44043 , \44361 );
xor \U$44863 ( \45240 , \45239 , \44386 );
xor \U$44864 ( \45241 , \45238 , \45240 );
xor \U$44865 ( \45242 , \44435 , \44815 );
xor \U$44866 ( \45243 , \45242 , \44820 );
and \U$44867 ( \45244 , \45241 , \45243 );
and \U$44868 ( \45245 , \45238 , \45240 );
or \U$44869 ( \45246 , \45244 , \45245 );
xor \U$44870 ( \45247 , \44823 , \44824 );
xor \U$44871 ( \45248 , \45247 , \44827 );
and \U$44872 ( \45249 , \45246 , \45248 );
and \U$44873 ( \45250 , \44842 , \45249 );
xor \U$44874 ( \45251 , \45249 , \44842 );
xor \U$44875 ( \45252 , \45246 , \45248 );
not \U$44876 ( \45253 , \45252 );
xor \U$44877 ( \45254 , \44449 , \44777 );
xor \U$44878 ( \45255 , \45254 , \44812 );
xor \U$44879 ( \45256 , \44686 , \44706 );
xor \U$44880 ( \45257 , \45256 , \44774 );
xor \U$44881 ( \45258 , \45220 , \45222 );
xor \U$44882 ( \45259 , \45258 , \45227 );
and \U$44883 ( \45260 , \45257 , \45259 );
xor \U$44884 ( \45261 , \44854 , \45190 );
xor \U$44885 ( \45262 , \45261 , \45215 );
xor \U$44886 ( \45263 , \45220 , \45222 );
xor \U$44887 ( \45264 , \45263 , \45227 );
and \U$44888 ( \45265 , \45262 , \45264 );
and \U$44889 ( \45266 , \45257 , \45262 );
or \U$44890 ( \45267 , \45260 , \45265 , \45266 );
xor \U$44891 ( \45268 , \45255 , \45267 );
xor \U$44892 ( \45269 , \45025 , \45048 );
xor \U$44893 ( \45270 , \45269 , \45074 );
xor \U$44894 ( \45271 , \44945 , \44970 );
xor \U$44895 ( \45272 , \45271 , \44997 );
and \U$44896 ( \45273 , \45270 , \45272 );
xor \U$44897 ( \45274 , \45103 , \45130 );
xor \U$44898 ( \45275 , \45274 , \45156 );
xor \U$44899 ( \45276 , \44945 , \44970 );
xor \U$44900 ( \45277 , \45276 , \44997 );
and \U$44901 ( \45278 , \45275 , \45277 );
and \U$44902 ( \45279 , \45270 , \45275 );
or \U$44903 ( \45280 , \45273 , \45278 , \45279 );
xor \U$44904 ( \45281 , \44474 , \44501 );
xor \U$44905 ( \45282 , \45281 , \44527 );
xor \U$44906 ( \45283 , \45280 , \45282 );
xor \U$44907 ( \45284 , \44866 , \44868 );
xor \U$44908 ( \45285 , \45284 , \44897 );
xor \U$44909 ( \45286 , \44856 , \44858 );
xor \U$44910 ( \45287 , \45286 , \44861 );
and \U$44911 ( \45288 , \45285 , \45287 );
xor \U$44912 ( \45289 , \44635 , \44642 );
xor \U$44913 ( \45290 , \45289 , \44651 );
xor \U$44914 ( \45291 , \44907 , \44912 );
xor \U$44915 ( \45292 , \45290 , \45291 );
xor \U$44916 ( \45293 , \44856 , \44858 );
xor \U$44917 ( \45294 , \45293 , \44861 );
and \U$44918 ( \45295 , \45292 , \45294 );
and \U$44919 ( \45296 , \45285 , \45292 );
or \U$44920 ( \45297 , \45288 , \45295 , \45296 );
and \U$44921 ( \45298 , \45283 , \45297 );
and \U$44922 ( \45299 , \45280 , \45282 );
or \U$44923 ( \45300 , \45298 , \45299 );
xor \U$44924 ( \45301 , \45111 , \45119 );
xor \U$44925 ( \45302 , \45301 , \45127 );
xor \U$44926 ( \45303 , \45138 , \45145 );
xor \U$44927 ( \45304 , \45303 , \45153 );
and \U$44928 ( \45305 , \45302 , \45304 );
xor \U$44929 ( \45306 , \45085 , \45092 );
xor \U$44930 ( \45307 , \45306 , \45100 );
xor \U$44931 ( \45308 , \45138 , \45145 );
xor \U$44932 ( \45309 , \45308 , \45153 );
and \U$44933 ( \45310 , \45307 , \45309 );
and \U$44934 ( \45311 , \45302 , \45307 );
or \U$44935 ( \45312 , \45305 , \45310 , \45311 );
not \U$44936 ( \45313 , \400 );
and \U$44937 ( \45314 , \436 , RIae77810_84);
and \U$44938 ( \45315 , RIae77900_86, \434 );
nor \U$44939 ( \45316 , \45314 , \45315 );
not \U$44940 ( \45317 , \45316 );
or \U$44941 ( \45318 , \45313 , \45317 );
or \U$44942 ( \45319 , \45316 , \402 );
nand \U$44943 ( \45320 , \45318 , \45319 );
not \U$44944 ( \45321 , \471 );
and \U$44945 ( \45322 , \514 , RIae76fa0_66);
and \U$44946 ( \45323 , RIae76eb0_64, \512 );
nor \U$44947 ( \45324 , \45322 , \45323 );
not \U$44948 ( \45325 , \45324 );
or \U$44949 ( \45326 , \45321 , \45325 );
or \U$44950 ( \45327 , \45324 , \471 );
nand \U$44951 ( \45328 , \45326 , \45327 );
xor \U$44952 ( \45329 , \45320 , \45328 );
and \U$44953 ( \45330 , \558 , RIae76dc0_62);
and \U$44954 ( \45331 , RIae76cd0_60, \556 );
nor \U$44955 ( \45332 , \45330 , \45331 );
and \U$44956 ( \45333 , \45332 , \504 );
not \U$44957 ( \45334 , \45332 );
and \U$44958 ( \45335 , \45334 , \562 );
nor \U$44959 ( \45336 , \45333 , \45335 );
and \U$44960 ( \45337 , \45329 , \45336 );
and \U$44961 ( \45338 , \45320 , \45328 );
or \U$44962 ( \45339 , \45337 , \45338 );
xor \U$44963 ( \45340 , \45339 , \44865 );
xor \U$44964 ( \45341 , \44877 , \44885 );
xor \U$44965 ( \45342 , \45341 , \44894 );
and \U$44966 ( \45343 , \45340 , \45342 );
and \U$44967 ( \45344 , \45339 , \44865 );
or \U$44968 ( \45345 , \45343 , \45344 );
xor \U$44969 ( \45346 , \45312 , \45345 );
xor \U$44970 ( \45347 , \44952 , \44959 );
xor \U$44971 ( \45348 , \45347 , \44967 );
xor \U$44972 ( \45349 , \44978 , \44985 );
xor \U$44973 ( \45350 , \45349 , \44994 );
xor \U$44974 ( \45351 , \45348 , \45350 );
xor \U$44975 ( \45352 , \44927 , \44934 );
xor \U$44976 ( \45353 , \45352 , \44942 );
and \U$44977 ( \45354 , \45351 , \45353 );
and \U$44978 ( \45355 , \45348 , \45350 );
or \U$44979 ( \45356 , \45354 , \45355 );
and \U$44980 ( \45357 , \45346 , \45356 );
and \U$44981 ( \45358 , \45312 , \45345 );
or \U$44982 ( \45359 , \45357 , \45358 );
not \U$44983 ( \45360 , \2789 );
and \U$44984 ( \45361 , \2783 , RIae789e0_122);
and \U$44985 ( \45362 , RIae788f0_120, \2781 );
nor \U$44986 ( \45363 , \45361 , \45362 );
not \U$44987 ( \45364 , \45363 );
or \U$44988 ( \45365 , \45360 , \45364 );
or \U$44989 ( \45366 , \45363 , \3089 );
nand \U$44990 ( \45367 , \45365 , \45366 );
and \U$44991 ( \45368 , \2224 , RIae77cc0_94);
and \U$44992 ( \45369 , RIae77bd0_92, \2222 );
nor \U$44993 ( \45370 , \45368 , \45369 );
and \U$44994 ( \45371 , \45370 , \2061 );
not \U$44995 ( \45372 , \45370 );
and \U$44996 ( \45373 , \45372 , \2060 );
nor \U$44997 ( \45374 , \45371 , \45373 );
xor \U$44998 ( \45375 , \45367 , \45374 );
and \U$44999 ( \45376 , \2607 , RIae77db0_96);
and \U$45000 ( \45377 , RIae77ea0_98, \2605 );
nor \U$45001 ( \45378 , \45376 , \45377 );
and \U$45002 ( \45379 , \45378 , \2611 );
not \U$45003 ( \45380 , \45378 );
and \U$45004 ( \45381 , \45380 , \2397 );
nor \U$45005 ( \45382 , \45379 , \45381 );
and \U$45006 ( \45383 , \45375 , \45382 );
and \U$45007 ( \45384 , \45367 , \45374 );
or \U$45008 ( \45385 , \45383 , \45384 );
and \U$45009 ( \45386 , \1939 , RIae78440_110);
and \U$45010 ( \45387 , RIae784b8_111, \1937 );
nor \U$45011 ( \45388 , \45386 , \45387 );
and \U$45012 ( \45389 , \45388 , \1735 );
not \U$45013 ( \45390 , \45388 );
and \U$45014 ( \45391 , \45390 , \1734 );
nor \U$45015 ( \45392 , \45389 , \45391 );
and \U$45016 ( \45393 , \1376 , RIae77f90_100);
and \U$45017 ( \45394 , RIae78080_102, \1374 );
nor \U$45018 ( \45395 , \45393 , \45394 );
and \U$45019 ( \45396 , \45395 , \1380 );
not \U$45020 ( \45397 , \45395 );
and \U$45021 ( \45398 , \45397 , \1261 );
nor \U$45022 ( \45399 , \45396 , \45398 );
xor \U$45023 ( \45400 , \45392 , \45399 );
and \U$45024 ( \45401 , \1593 , RIae78260_106);
and \U$45025 ( \45402 , RIae78620_114, \1591 );
nor \U$45026 ( \45403 , \45401 , \45402 );
and \U$45027 ( \45404 , \45403 , \1498 );
not \U$45028 ( \45405 , \45403 );
and \U$45029 ( \45406 , \45405 , \1488 );
nor \U$45030 ( \45407 , \45404 , \45406 );
and \U$45031 ( \45408 , \45400 , \45407 );
and \U$45032 ( \45409 , \45392 , \45399 );
or \U$45033 ( \45410 , \45408 , \45409 );
xor \U$45034 ( \45411 , \45385 , \45410 );
and \U$45035 ( \45412 , \1138 , RIae78350_108);
and \U$45036 ( \45413 , RIae78170_104, \1136 );
nor \U$45037 ( \45414 , \45412 , \45413 );
and \U$45038 ( \45415 , \45414 , \1012 );
not \U$45039 ( \45416 , \45414 );
and \U$45040 ( \45417 , \45416 , \1142 );
nor \U$45041 ( \45418 , \45415 , \45417 );
and \U$45042 ( \45419 , \672 , RIae77108_69);
and \U$45043 ( \45420 , RIae77090_68, \670 );
nor \U$45044 ( \45421 , \45419 , \45420 );
and \U$45045 ( \45422 , \45421 , \588 );
not \U$45046 ( \45423 , \45421 );
and \U$45047 ( \45424 , \45423 , \587 );
nor \U$45048 ( \45425 , \45422 , \45424 );
xor \U$45049 ( \45426 , \45418 , \45425 );
not \U$45050 ( \45427 , \787 );
and \U$45051 ( \45428 , \883 , RIae77270_72);
and \U$45052 ( \45429 , RIae77360_74, \881 );
nor \U$45053 ( \45430 , \45428 , \45429 );
not \U$45054 ( \45431 , \45430 );
or \U$45055 ( \45432 , \45427 , \45431 );
or \U$45056 ( \45433 , \45430 , \787 );
nand \U$45057 ( \45434 , \45432 , \45433 );
and \U$45058 ( \45435 , \45426 , \45434 );
and \U$45059 ( \45436 , \45418 , \45425 );
or \U$45060 ( \45437 , \45435 , \45436 );
and \U$45061 ( \45438 , \45411 , \45437 );
and \U$45062 ( \45439 , \45385 , \45410 );
or \U$45063 ( \45440 , \45438 , \45439 );
and \U$45064 ( \45441 , \8371 , RIae76460_42);
and \U$45065 ( \45442 , RIae76550_44, \8369 );
nor \U$45066 ( \45443 , \45441 , \45442 );
and \U$45067 ( \45444 , \45443 , \8020 );
not \U$45068 ( \45445 , \45443 );
and \U$45069 ( \45446 , \45445 , \8019 );
nor \U$45070 ( \45447 , \45444 , \45446 );
and \U$45071 ( \45448 , \8966 , RIae76730_48);
and \U$45072 ( \45449 , RIae76640_46, \8964 );
nor \U$45073 ( \45450 , \45448 , \45449 );
and \U$45074 ( \45451 , \45450 , \8799 );
not \U$45075 ( \45452 , \45450 );
and \U$45076 ( \45453 , \45452 , \8789 );
nor \U$45077 ( \45454 , \45451 , \45453 );
xor \U$45078 ( \45455 , \45447 , \45454 );
and \U$45079 ( \45456 , \9760 , RIae76190_36);
and \U$45080 ( \45457 , RIae760a0_34, \9758 );
nor \U$45081 ( \45458 , \45456 , \45457 );
and \U$45082 ( \45459 , \45458 , \9273 );
not \U$45083 ( \45460 , \45458 );
and \U$45084 ( \45461 , \45460 , \9764 );
nor \U$45085 ( \45462 , \45459 , \45461 );
and \U$45086 ( \45463 , \45455 , \45462 );
and \U$45087 ( \45464 , \45447 , \45454 );
or \U$45088 ( \45465 , \45463 , \45464 );
and \U$45089 ( \45466 , \13059 , RIae76be0_58);
and \U$45090 ( \45467 , RIae78ad0_124, \13057 );
nor \U$45091 ( \45468 , \45466 , \45467 );
and \U$45092 ( \45469 , \45468 , \13063 );
not \U$45093 ( \45470 , \45468 );
and \U$45094 ( \45471 , \45470 , \12718 );
nor \U$45095 ( \45472 , \45469 , \45471 );
xor \U$45096 ( \45473 , \45472 , \14463 );
and \U$45097 ( \45474 , \14059 , RIae78d28_129);
and \U$45098 ( \45475 , RIae78e18_131, \14057 );
nor \U$45099 ( \45476 , \45474 , \45475 );
and \U$45100 ( \45477 , \45476 , \13502 );
not \U$45101 ( \45478 , \45476 );
and \U$45102 ( \45479 , \45478 , \14063 );
nor \U$45103 ( \45480 , \45477 , \45479 );
and \U$45104 ( \45481 , \45473 , \45480 );
and \U$45105 ( \45482 , \45472 , \14463 );
or \U$45106 ( \45483 , \45481 , \45482 );
xor \U$45107 ( \45484 , \45465 , \45483 );
and \U$45108 ( \45485 , \12180 , RIae76820_50);
and \U$45109 ( \45486 , RIae76910_52, \12178 );
nor \U$45110 ( \45487 , \45485 , \45486 );
and \U$45111 ( \45488 , \45487 , \12184 );
not \U$45112 ( \45489 , \45487 );
and \U$45113 ( \45490 , \45489 , \11827 );
nor \U$45114 ( \45491 , \45488 , \45490 );
and \U$45115 ( \45492 , \10548 , RIae76370_40);
and \U$45116 ( \45493 , RIae76280_38, \10546 );
nor \U$45117 ( \45494 , \45492 , \45493 );
and \U$45118 ( \45495 , \45494 , \10421 );
not \U$45119 ( \45496 , \45494 );
and \U$45120 ( \45497 , \45496 , \10118 );
nor \U$45121 ( \45498 , \45495 , \45497 );
xor \U$45122 ( \45499 , \45491 , \45498 );
and \U$45123 ( \45500 , \11470 , RIae76af0_56);
and \U$45124 ( \45501 , RIae76a00_54, \11468 );
nor \U$45125 ( \45502 , \45500 , \45501 );
and \U$45126 ( \45503 , \45502 , \10936 );
not \U$45127 ( \45504 , \45502 );
and \U$45128 ( \45505 , \45504 , \11474 );
nor \U$45129 ( \45506 , \45503 , \45505 );
and \U$45130 ( \45507 , \45499 , \45506 );
and \U$45131 ( \45508 , \45491 , \45498 );
or \U$45132 ( \45509 , \45507 , \45508 );
and \U$45133 ( \45510 , \45484 , \45509 );
and \U$45134 ( \45511 , \45465 , \45483 );
or \U$45135 ( \45512 , \45510 , \45511 );
xor \U$45136 ( \45513 , \45440 , \45512 );
and \U$45137 ( \45514 , \6941 , RIae75290_4);
and \U$45138 ( \45515 , RIae751a0_2, \6939 );
nor \U$45139 ( \45516 , \45514 , \45515 );
and \U$45140 ( \45517 , \45516 , \6314 );
not \U$45141 ( \45518 , \45516 );
and \U$45142 ( \45519 , \45518 , \6945 );
nor \U$45143 ( \45520 , \45517 , \45519 );
and \U$45144 ( \45521 , \6172 , RIae75830_16);
and \U$45145 ( \45522 , RIae75740_14, \6170 );
nor \U$45146 ( \45523 , \45521 , \45522 );
and \U$45147 ( \45524 , \45523 , \6176 );
not \U$45148 ( \45525 , \45523 );
and \U$45149 ( \45526 , \45525 , \6175 );
nor \U$45150 ( \45527 , \45524 , \45526 );
xor \U$45151 ( \45528 , \45520 , \45527 );
and \U$45152 ( \45529 , \7633 , RIae75380_6);
and \U$45153 ( \45530 , RIae75470_8, \7631 );
nor \U$45154 ( \45531 , \45529 , \45530 );
and \U$45155 ( \45532 , \45531 , \7206 );
not \U$45156 ( \45533 , \45531 );
and \U$45157 ( \45534 , \45533 , \7205 );
nor \U$45158 ( \45535 , \45532 , \45534 );
and \U$45159 ( \45536 , \45528 , \45535 );
and \U$45160 ( \45537 , \45520 , \45527 );
or \U$45161 ( \45538 , \45536 , \45537 );
and \U$45162 ( \45539 , \5896 , RIae75650_12);
and \U$45163 ( \45540 , RIae75560_10, \5894 );
nor \U$45164 ( \45541 , \45539 , \45540 );
and \U$45165 ( \45542 , \45541 , \5590 );
not \U$45166 ( \45543 , \45541 );
and \U$45167 ( \45544 , \45543 , \5589 );
nor \U$45168 ( \45545 , \45542 , \45544 );
and \U$45169 ( \45546 , \4688 , RIae75fb0_32);
and \U$45170 ( \45547 , RIae75ec0_30, \4686 );
nor \U$45171 ( \45548 , \45546 , \45547 );
and \U$45172 ( \45549 , \45548 , \4481 );
not \U$45173 ( \45550 , \45548 );
and \U$45174 ( \45551 , \45550 , \4482 );
nor \U$45175 ( \45552 , \45549 , \45551 );
xor \U$45176 ( \45553 , \45545 , \45552 );
and \U$45177 ( \45554 , \5399 , RIae75ce0_26);
and \U$45178 ( \45555 , RIae75dd0_28, \5397 );
nor \U$45179 ( \45556 , \45554 , \45555 );
and \U$45180 ( \45557 , \45556 , \5016 );
not \U$45181 ( \45558 , \45556 );
and \U$45182 ( \45559 , \45558 , \5403 );
nor \U$45183 ( \45560 , \45557 , \45559 );
and \U$45184 ( \45561 , \45553 , \45560 );
and \U$45185 ( \45562 , \45545 , \45552 );
or \U$45186 ( \45563 , \45561 , \45562 );
xor \U$45187 ( \45564 , \45538 , \45563 );
and \U$45188 ( \45565 , \4247 , RIae75a10_20);
and \U$45189 ( \45566 , RIae75920_18, \4245 );
nor \U$45190 ( \45567 , \45565 , \45566 );
and \U$45191 ( \45568 , \45567 , \3989 );
not \U$45192 ( \45569 , \45567 );
and \U$45193 ( \45570 , \45569 , \4251 );
nor \U$45194 ( \45571 , \45568 , \45570 );
not \U$45195 ( \45572 , \2774 );
and \U$45196 ( \45573 , \3214 , RIae78800_118);
and \U$45197 ( \45574 , RIae78710_116, \3212 );
nor \U$45198 ( \45575 , \45573 , \45574 );
not \U$45199 ( \45576 , \45575 );
or \U$45200 ( \45577 , \45572 , \45576 );
or \U$45201 ( \45578 , \45575 , \3218 );
nand \U$45202 ( \45579 , \45577 , \45578 );
xor \U$45203 ( \45580 , \45571 , \45579 );
and \U$45204 ( \45581 , \3730 , RIae75bf0_24);
and \U$45205 ( \45582 , RIae75b00_22, \3728 );
nor \U$45206 ( \45583 , \45581 , \45582 );
and \U$45207 ( \45584 , \45583 , \3732 );
not \U$45208 ( \45585 , \45583 );
and \U$45209 ( \45586 , \45585 , \3422 );
nor \U$45210 ( \45587 , \45584 , \45586 );
and \U$45211 ( \45588 , \45580 , \45587 );
and \U$45212 ( \45589 , \45571 , \45579 );
or \U$45213 ( \45590 , \45588 , \45589 );
and \U$45214 ( \45591 , \45564 , \45590 );
and \U$45215 ( \45592 , \45538 , \45563 );
or \U$45216 ( \45593 , \45591 , \45592 );
and \U$45217 ( \45594 , \45513 , \45593 );
and \U$45218 ( \45595 , \45440 , \45512 );
or \U$45219 ( \45596 , \45594 , \45595 );
xor \U$45220 ( \45597 , \45359 , \45596 );
xor \U$45221 ( \45598 , \45032 , \45037 );
xor \U$45222 ( \45599 , \45598 , \45045 );
xor \U$45223 ( \45600 , \45007 , \45014 );
xor \U$45224 ( \45601 , \45600 , \45022 );
and \U$45225 ( \45602 , \45599 , \45601 );
xor \U$45226 ( \45603 , \45056 , \45063 );
xor \U$45227 ( \45604 , \45603 , \45071 );
xor \U$45228 ( \45605 , \45007 , \45014 );
xor \U$45229 ( \45606 , \45605 , \45022 );
and \U$45230 ( \45607 , \45604 , \45606 );
and \U$45231 ( \45608 , \45599 , \45604 );
or \U$45232 ( \45609 , \45602 , \45607 , \45608 );
xor \U$45233 ( \45610 , \44562 , \13502 );
xor \U$45234 ( \45611 , \45610 , \44570 );
xor \U$45235 ( \45612 , \45609 , \45611 );
xor \U$45236 ( \45613 , \44509 , \44516 );
xor \U$45237 ( \45614 , \45613 , \44524 );
xor \U$45238 ( \45615 , \45165 , \45170 );
xor \U$45239 ( \45616 , \45614 , \45615 );
and \U$45240 ( \45617 , \45612 , \45616 );
and \U$45241 ( \45618 , \45609 , \45611 );
or \U$45242 ( \45619 , \45617 , \45618 );
and \U$45243 ( \45620 , \45597 , \45619 );
and \U$45244 ( \45621 , \45359 , \45596 );
or \U$45245 ( \45622 , \45620 , \45621 );
xor \U$45246 ( \45623 , \45300 , \45622 );
xor \U$45247 ( \45624 , \44555 , \44573 );
xor \U$45248 ( \45625 , \45624 , \44599 );
xor \U$45249 ( \45626 , \45197 , \45199 );
xor \U$45250 ( \45627 , \45626 , \45204 );
and \U$45251 ( \45628 , \45625 , \45627 );
xor \U$45252 ( \45629 , \44709 , \44711 );
xor \U$45253 ( \45630 , \45629 , \44714 );
xor \U$45254 ( \45631 , \45175 , \45182 );
xor \U$45255 ( \45632 , \45630 , \45631 );
xor \U$45256 ( \45633 , \45197 , \45199 );
xor \U$45257 ( \45634 , \45633 , \45204 );
and \U$45258 ( \45635 , \45632 , \45634 );
and \U$45259 ( \45636 , \45625 , \45632 );
or \U$45260 ( \45637 , \45628 , \45635 , \45636 );
and \U$45261 ( \45638 , \45623 , \45637 );
and \U$45262 ( \45639 , \45300 , \45622 );
or \U$45263 ( \45640 , \45638 , \45639 );
xor \U$45264 ( \45641 , \44790 , \44792 );
xor \U$45265 ( \45642 , \45641 , \44809 );
xor \U$45266 ( \45643 , \45640 , \45642 );
xor \U$45267 ( \45644 , \44920 , \45162 );
xor \U$45268 ( \45645 , \45644 , \45187 );
xor \U$45269 ( \45646 , \45195 , \45207 );
xor \U$45270 ( \45647 , \45646 , \45212 );
and \U$45271 ( \45648 , \45645 , \45647 );
xor \U$45272 ( \45649 , \44688 , \44690 );
xor \U$45273 ( \45650 , \45649 , \44703 );
xor \U$45274 ( \45651 , \44844 , \44849 );
xor \U$45275 ( \45652 , \45650 , \45651 );
xor \U$45276 ( \45653 , \45195 , \45207 );
xor \U$45277 ( \45654 , \45653 , \45212 );
and \U$45278 ( \45655 , \45652 , \45654 );
and \U$45279 ( \45656 , \45645 , \45652 );
or \U$45280 ( \45657 , \45648 , \45655 , \45656 );
and \U$45281 ( \45658 , \45643 , \45657 );
and \U$45282 ( \45659 , \45640 , \45642 );
or \U$45283 ( \45660 , \45658 , \45659 );
and \U$45284 ( \45661 , \45268 , \45660 );
and \U$45285 ( \45662 , \45255 , \45267 );
nor \U$45286 ( \45663 , \45661 , \45662 );
not \U$45287 ( \45664 , \45663 );
xor \U$45288 ( \45665 , \45238 , \45240 );
xor \U$45289 ( \45666 , \45665 , \45243 );
nand \U$45290 ( \45667 , \45664 , \45666 );
or \U$45291 ( \45668 , \45253 , \45667 );
not \U$45292 ( \45669 , \45252 );
not \U$45293 ( \45670 , \45667 );
and \U$45294 ( \45671 , \45669 , \45670 );
and \U$45295 ( \45672 , \45252 , \45667 );
nor \U$45296 ( \45673 , \45671 , \45672 );
not \U$45297 ( \45674 , RIae77450_76);
nor \U$45298 ( \45675 , \45674 , \491 );
xor \U$45299 ( \45676 , \45320 , \45328 );
xor \U$45300 ( \45677 , \45676 , \45336 );
and \U$45301 ( \45678 , \45675 , \45677 );
xor \U$45302 ( \45679 , \45418 , \45425 );
xor \U$45303 ( \45680 , \45679 , \45434 );
xor \U$45304 ( \45681 , \45320 , \45328 );
xor \U$45305 ( \45682 , \45681 , \45336 );
and \U$45306 ( \45683 , \45680 , \45682 );
and \U$45307 ( \45684 , \45675 , \45680 );
or \U$45308 ( \45685 , \45678 , \45683 , \45684 );
nand \U$45309 ( \45686 , RIae776a8_81, RIae78b48_125);
and \U$45310 ( \45687 , \384 , RIae77450_76);
and \U$45311 ( \45688 , RIae77ae0_90, \382 );
nor \U$45312 ( \45689 , \45687 , \45688 );
not \U$45313 ( \45690 , \45689 );
not \U$45314 ( \45691 , \388 );
and \U$45315 ( \45692 , \45690 , \45691 );
and \U$45316 ( \45693 , \45689 , \392 );
nor \U$45317 ( \45694 , \45692 , \45693 );
nand \U$45318 ( \45695 , \45686 , \45694 );
not \U$45319 ( \45696 , \388 );
and \U$45320 ( \45697 , \384 , RIae77ae0_90);
and \U$45321 ( \45698 , RIae779f0_88, \382 );
nor \U$45322 ( \45699 , \45697 , \45698 );
not \U$45323 ( \45700 , \45699 );
or \U$45324 ( \45701 , \45696 , \45700 );
or \U$45325 ( \45702 , \45699 , \392 );
nand \U$45326 ( \45703 , \45701 , \45702 );
xor \U$45327 ( \45704 , \45695 , \45703 );
and \U$45328 ( \45705 , \558 , RIae76eb0_64);
and \U$45329 ( \45706 , RIae76dc0_62, \556 );
nor \U$45330 ( \45707 , \45705 , \45706 );
and \U$45331 ( \45708 , \45707 , \504 );
not \U$45332 ( \45709 , \45707 );
and \U$45333 ( \45710 , \45709 , \562 );
nor \U$45334 ( \45711 , \45708 , \45710 );
not \U$45335 ( \45712 , \400 );
and \U$45336 ( \45713 , \436 , RIae779f0_88);
and \U$45337 ( \45714 , RIae77810_84, \434 );
nor \U$45338 ( \45715 , \45713 , \45714 );
not \U$45339 ( \45716 , \45715 );
or \U$45340 ( \45717 , \45712 , \45716 );
or \U$45341 ( \45718 , \45715 , \400 );
nand \U$45342 ( \45719 , \45717 , \45718 );
xor \U$45343 ( \45720 , \45711 , \45719 );
not \U$45344 ( \45721 , \471 );
and \U$45345 ( \45722 , \514 , RIae77900_86);
and \U$45346 ( \45723 , RIae76fa0_66, \512 );
nor \U$45347 ( \45724 , \45722 , \45723 );
not \U$45348 ( \45725 , \45724 );
or \U$45349 ( \45726 , \45721 , \45725 );
or \U$45350 ( \45727 , \45724 , \471 );
nand \U$45351 ( \45728 , \45726 , \45727 );
and \U$45352 ( \45729 , \45720 , \45728 );
and \U$45353 ( \45730 , \45711 , \45719 );
or \U$45354 ( \45731 , \45729 , \45730 );
and \U$45355 ( \45732 , \45704 , \45731 );
and \U$45356 ( \45733 , \45695 , \45703 );
or \U$45357 ( \45734 , \45732 , \45733 );
xor \U$45358 ( \45735 , \45685 , \45734 );
xor \U$45359 ( \45736 , \45367 , \45374 );
xor \U$45360 ( \45737 , \45736 , \45382 );
xor \U$45361 ( \45738 , \45392 , \45399 );
xor \U$45362 ( \45739 , \45738 , \45407 );
xor \U$45363 ( \45740 , \45737 , \45739 );
xor \U$45364 ( \45741 , \45571 , \45579 );
xor \U$45365 ( \45742 , \45741 , \45587 );
and \U$45366 ( \45743 , \45740 , \45742 );
and \U$45367 ( \45744 , \45737 , \45739 );
or \U$45368 ( \45745 , \45743 , \45744 );
xor \U$45369 ( \45746 , \45735 , \45745 );
xor \U$45370 ( \45747 , \45545 , \45552 );
xor \U$45371 ( \45748 , \45747 , \45560 );
xor \U$45372 ( \45749 , \45520 , \45527 );
xor \U$45373 ( \45750 , \45749 , \45535 );
and \U$45374 ( \45751 , \45748 , \45750 );
xor \U$45375 ( \45752 , \45447 , \45454 );
xor \U$45376 ( \45753 , \45752 , \45462 );
xor \U$45377 ( \45754 , \45520 , \45527 );
xor \U$45378 ( \45755 , \45754 , \45535 );
and \U$45379 ( \45756 , \45753 , \45755 );
and \U$45380 ( \45757 , \45748 , \45753 );
or \U$45381 ( \45758 , \45751 , \45756 , \45757 );
xor \U$45382 ( \45759 , \45491 , \45498 );
xor \U$45383 ( \45760 , \45759 , \45506 );
xor \U$45384 ( \45761 , \45472 , \14463 );
xor \U$45385 ( \45762 , \45761 , \45480 );
and \U$45386 ( \45763 , \45760 , \45762 );
xor \U$45387 ( \45764 , \45758 , \45763 );
xor \U$45388 ( \45765 , \45007 , \45014 );
xor \U$45389 ( \45766 , \45765 , \45022 );
xor \U$45390 ( \45767 , \45599 , \45604 );
xor \U$45391 ( \45768 , \45766 , \45767 );
xor \U$45392 ( \45769 , \45764 , \45768 );
and \U$45393 ( \45770 , \45746 , \45769 );
xor \U$45394 ( \45771 , \45348 , \45350 );
xor \U$45395 ( \45772 , \45771 , \45353 );
xor \U$45396 ( \45773 , \45339 , \44865 );
xor \U$45397 ( \45774 , \45773 , \45342 );
xor \U$45398 ( \45775 , \45138 , \45145 );
xor \U$45399 ( \45776 , \45775 , \45153 );
xor \U$45400 ( \45777 , \45302 , \45307 );
xor \U$45401 ( \45778 , \45776 , \45777 );
xor \U$45402 ( \45779 , \45774 , \45778 );
xor \U$45403 ( \45780 , \45772 , \45779 );
xor \U$45404 ( \45781 , \45758 , \45763 );
xor \U$45405 ( \45782 , \45781 , \45768 );
and \U$45406 ( \45783 , \45780 , \45782 );
and \U$45407 ( \45784 , \45746 , \45780 );
or \U$45408 ( \45785 , \45770 , \45783 , \45784 );
not \U$45409 ( \45786 , \2789 );
and \U$45410 ( \45787 , \2783 , RIae77ea0_98);
and \U$45411 ( \45788 , RIae789e0_122, \2781 );
nor \U$45412 ( \45789 , \45787 , \45788 );
not \U$45413 ( \45790 , \45789 );
or \U$45414 ( \45791 , \45786 , \45790 );
or \U$45415 ( \45792 , \45789 , \3089 );
nand \U$45416 ( \45793 , \45791 , \45792 );
and \U$45417 ( \45794 , \2224 , RIae784b8_111);
and \U$45418 ( \45795 , RIae77cc0_94, \2222 );
nor \U$45419 ( \45796 , \45794 , \45795 );
and \U$45420 ( \45797 , \45796 , \2061 );
not \U$45421 ( \45798 , \45796 );
and \U$45422 ( \45799 , \45798 , \2060 );
nor \U$45423 ( \45800 , \45797 , \45799 );
xor \U$45424 ( \45801 , \45793 , \45800 );
and \U$45425 ( \45802 , \2607 , RIae77bd0_92);
and \U$45426 ( \45803 , RIae77db0_96, \2605 );
nor \U$45427 ( \45804 , \45802 , \45803 );
and \U$45428 ( \45805 , \45804 , \2611 );
not \U$45429 ( \45806 , \45804 );
and \U$45430 ( \45807 , \45806 , \2397 );
nor \U$45431 ( \45808 , \45805 , \45807 );
xor \U$45432 ( \45809 , \45801 , \45808 );
and \U$45433 ( \45810 , \3730 , RIae78710_116);
and \U$45434 ( \45811 , RIae75bf0_24, \3728 );
nor \U$45435 ( \45812 , \45810 , \45811 );
and \U$45436 ( \45813 , \45812 , \3732 );
not \U$45437 ( \45814 , \45812 );
and \U$45438 ( \45815 , \45814 , \3422 );
nor \U$45439 ( \45816 , \45813 , \45815 );
not \U$45440 ( \45817 , \2774 );
and \U$45441 ( \45818 , \3214 , RIae788f0_120);
and \U$45442 ( \45819 , RIae78800_118, \3212 );
nor \U$45443 ( \45820 , \45818 , \45819 );
not \U$45444 ( \45821 , \45820 );
or \U$45445 ( \45822 , \45817 , \45821 );
or \U$45446 ( \45823 , \45820 , \3218 );
nand \U$45447 ( \45824 , \45822 , \45823 );
xor \U$45448 ( \45825 , \45816 , \45824 );
and \U$45449 ( \45826 , \4247 , RIae75b00_22);
and \U$45450 ( \45827 , RIae75a10_20, \4245 );
nor \U$45451 ( \45828 , \45826 , \45827 );
and \U$45452 ( \45829 , \45828 , \3989 );
not \U$45453 ( \45830 , \45828 );
and \U$45454 ( \45831 , \45830 , \4251 );
nor \U$45455 ( \45832 , \45829 , \45831 );
xor \U$45456 ( \45833 , \45825 , \45832 );
xor \U$45457 ( \45834 , \45809 , \45833 );
and \U$45458 ( \45835 , \5399 , RIae75ec0_30);
and \U$45459 ( \45836 , RIae75ce0_26, \5397 );
nor \U$45460 ( \45837 , \45835 , \45836 );
and \U$45461 ( \45838 , \45837 , \5016 );
not \U$45462 ( \45839 , \45837 );
and \U$45463 ( \45840 , \45839 , \5403 );
nor \U$45464 ( \45841 , \45838 , \45840 );
and \U$45465 ( \45842 , \4688 , RIae75920_18);
and \U$45466 ( \45843 , RIae75fb0_32, \4686 );
nor \U$45467 ( \45844 , \45842 , \45843 );
and \U$45468 ( \45845 , \45844 , \4481 );
not \U$45469 ( \45846 , \45844 );
and \U$45470 ( \45847 , \45846 , \4482 );
nor \U$45471 ( \45848 , \45845 , \45847 );
xor \U$45472 ( \45849 , \45841 , \45848 );
and \U$45473 ( \45850 , \5896 , RIae75dd0_28);
and \U$45474 ( \45851 , RIae75650_12, \5894 );
nor \U$45475 ( \45852 , \45850 , \45851 );
and \U$45476 ( \45853 , \45852 , \5590 );
not \U$45477 ( \45854 , \45852 );
and \U$45478 ( \45855 , \45854 , \5589 );
nor \U$45479 ( \45856 , \45853 , \45855 );
xor \U$45480 ( \45857 , \45849 , \45856 );
and \U$45481 ( \45858 , \45834 , \45857 );
and \U$45482 ( \45859 , \45809 , \45833 );
or \U$45483 ( \45860 , \45858 , \45859 );
not \U$45484 ( \45861 , \388 );
and \U$45485 ( \45862 , \384 , RIae776a8_81);
and \U$45486 ( \45863 , RIae77450_76, \382 );
nor \U$45487 ( \45864 , \45862 , \45863 );
not \U$45488 ( \45865 , \45864 );
or \U$45489 ( \45866 , \45861 , \45865 );
or \U$45490 ( \45867 , \45864 , \392 );
nand \U$45491 ( \45868 , \45866 , \45867 );
not \U$45492 ( \45869 , RIae77540_78);
nor \U$45493 ( \45870 , \45869 , \491 );
xor \U$45494 ( \45871 , \45868 , \45870 );
not \U$45495 ( \45872 , \402 );
and \U$45496 ( \45873 , \436 , RIae77ae0_90);
and \U$45497 ( \45874 , RIae779f0_88, \434 );
nor \U$45498 ( \45875 , \45873 , \45874 );
not \U$45499 ( \45876 , \45875 );
or \U$45500 ( \45877 , \45872 , \45876 );
or \U$45501 ( \45878 , \45875 , \400 );
nand \U$45502 ( \45879 , \45877 , \45878 );
and \U$45503 ( \45880 , \45871 , \45879 );
and \U$45504 ( \45881 , \45868 , \45870 );
or \U$45505 ( \45882 , \45880 , \45881 );
or \U$45506 ( \45883 , \45694 , \45686 );
nand \U$45507 ( \45884 , \45883 , \45695 );
xor \U$45508 ( \45885 , \45882 , \45884 );
and \U$45509 ( \45886 , \672 , RIae76dc0_62);
and \U$45510 ( \45887 , RIae76cd0_60, \670 );
nor \U$45511 ( \45888 , \45886 , \45887 );
and \U$45512 ( \45889 , \45888 , \588 );
not \U$45513 ( \45890 , \45888 );
and \U$45514 ( \45891 , \45890 , \587 );
nor \U$45515 ( \45892 , \45889 , \45891 );
not \U$45516 ( \45893 , \471 );
and \U$45517 ( \45894 , \514 , RIae77810_84);
and \U$45518 ( \45895 , RIae77900_86, \512 );
nor \U$45519 ( \45896 , \45894 , \45895 );
not \U$45520 ( \45897 , \45896 );
or \U$45521 ( \45898 , \45893 , \45897 );
or \U$45522 ( \45899 , \45896 , \471 );
nand \U$45523 ( \45900 , \45898 , \45899 );
xor \U$45524 ( \45901 , \45892 , \45900 );
and \U$45525 ( \45902 , \558 , RIae76fa0_66);
and \U$45526 ( \45903 , RIae76eb0_64, \556 );
nor \U$45527 ( \45904 , \45902 , \45903 );
and \U$45528 ( \45905 , \45904 , \504 );
not \U$45529 ( \45906 , \45904 );
and \U$45530 ( \45907 , \45906 , \562 );
nor \U$45531 ( \45908 , \45905 , \45907 );
and \U$45532 ( \45909 , \45901 , \45908 );
and \U$45533 ( \45910 , \45892 , \45900 );
or \U$45534 ( \45911 , \45909 , \45910 );
and \U$45535 ( \45912 , \45885 , \45911 );
and \U$45536 ( \45913 , \45882 , \45884 );
or \U$45537 ( \45914 , \45912 , \45913 );
xor \U$45538 ( \45915 , \45860 , \45914 );
and \U$45539 ( \45916 , \1138 , RIae77360_74);
and \U$45540 ( \45917 , RIae78350_108, \1136 );
nor \U$45541 ( \45918 , \45916 , \45917 );
and \U$45542 ( \45919 , \45918 , \1012 );
not \U$45543 ( \45920 , \45918 );
and \U$45544 ( \45921 , \45920 , \1142 );
nor \U$45545 ( \45922 , \45919 , \45921 );
and \U$45546 ( \45923 , \672 , RIae76cd0_60);
and \U$45547 ( \45924 , RIae77108_69, \670 );
nor \U$45548 ( \45925 , \45923 , \45924 );
and \U$45549 ( \45926 , \45925 , \588 );
not \U$45550 ( \45927 , \45925 );
and \U$45551 ( \45928 , \45927 , \587 );
nor \U$45552 ( \45929 , \45926 , \45928 );
xor \U$45553 ( \45930 , \45922 , \45929 );
not \U$45554 ( \45931 , \789 );
and \U$45555 ( \45932 , \883 , RIae77090_68);
and \U$45556 ( \45933 , RIae77270_72, \881 );
nor \U$45557 ( \45934 , \45932 , \45933 );
not \U$45558 ( \45935 , \45934 );
or \U$45559 ( \45936 , \45931 , \45935 );
or \U$45560 ( \45937 , \45934 , \787 );
nand \U$45561 ( \45938 , \45936 , \45937 );
xor \U$45562 ( \45939 , \45930 , \45938 );
xor \U$45563 ( \45940 , \45711 , \45719 );
xor \U$45564 ( \45941 , \45940 , \45728 );
and \U$45565 ( \45942 , \45939 , \45941 );
and \U$45566 ( \45943 , \1939 , RIae78620_114);
and \U$45567 ( \45944 , RIae78440_110, \1937 );
nor \U$45568 ( \45945 , \45943 , \45944 );
and \U$45569 ( \45946 , \45945 , \1735 );
not \U$45570 ( \45947 , \45945 );
and \U$45571 ( \45948 , \45947 , \1734 );
nor \U$45572 ( \45949 , \45946 , \45948 );
and \U$45573 ( \45950 , \1376 , RIae78170_104);
and \U$45574 ( \45951 , RIae77f90_100, \1374 );
nor \U$45575 ( \45952 , \45950 , \45951 );
and \U$45576 ( \45953 , \45952 , \1380 );
not \U$45577 ( \45954 , \45952 );
and \U$45578 ( \45955 , \45954 , \1261 );
nor \U$45579 ( \45956 , \45953 , \45955 );
xor \U$45580 ( \45957 , \45949 , \45956 );
and \U$45581 ( \45958 , \1593 , RIae78080_102);
and \U$45582 ( \45959 , RIae78260_106, \1591 );
nor \U$45583 ( \45960 , \45958 , \45959 );
and \U$45584 ( \45961 , \45960 , \1498 );
not \U$45585 ( \45962 , \45960 );
and \U$45586 ( \45963 , \45962 , \1488 );
nor \U$45587 ( \45964 , \45961 , \45963 );
xor \U$45588 ( \45965 , \45957 , \45964 );
xor \U$45589 ( \45966 , \45711 , \45719 );
xor \U$45590 ( \45967 , \45966 , \45728 );
and \U$45591 ( \45968 , \45965 , \45967 );
and \U$45592 ( \45969 , \45939 , \45965 );
or \U$45593 ( \45970 , \45942 , \45968 , \45969 );
and \U$45594 ( \45971 , \45915 , \45970 );
and \U$45595 ( \45972 , \45860 , \45914 );
or \U$45596 ( \45973 , \45971 , \45972 );
and \U$45597 ( \45974 , \6941 , RIae75830_16);
and \U$45598 ( \45975 , RIae75740_14, \6939 );
nor \U$45599 ( \45976 , \45974 , \45975 );
and \U$45600 ( \45977 , \45976 , \6945 );
not \U$45601 ( \45978 , \45976 );
and \U$45602 ( \45979 , \45978 , \6314 );
nor \U$45603 ( \45980 , \45977 , \45979 );
and \U$45604 ( \45981 , \8371 , RIae75380_6);
and \U$45605 ( \45982 , RIae75470_8, \8369 );
nor \U$45606 ( \45983 , \45981 , \45982 );
and \U$45607 ( \45984 , \45983 , \8019 );
not \U$45608 ( \45985 , \45983 );
and \U$45609 ( \45986 , \45985 , \8020 );
nor \U$45610 ( \45987 , \45984 , \45986 );
or \U$45611 ( \45988 , \45980 , \45987 );
not \U$45612 ( \45989 , \45987 );
not \U$45613 ( \45990 , \45980 );
or \U$45614 ( \45991 , \45989 , \45990 );
and \U$45615 ( \45992 , \7633 , RIae75290_4);
and \U$45616 ( \45993 , RIae751a0_2, \7631 );
nor \U$45617 ( \45994 , \45992 , \45993 );
and \U$45618 ( \45995 , \45994 , \7206 );
not \U$45619 ( \45996 , \45994 );
and \U$45620 ( \45997 , \45996 , \7205 );
nor \U$45621 ( \45998 , \45995 , \45997 );
nand \U$45622 ( \45999 , \45991 , \45998 );
nand \U$45623 ( \46000 , \45988 , \45999 );
and \U$45624 ( \46001 , \5399 , RIae75fb0_32);
and \U$45625 ( \46002 , RIae75ec0_30, \5397 );
nor \U$45626 ( \46003 , \46001 , \46002 );
and \U$45627 ( \46004 , \46003 , \5403 );
not \U$45628 ( \46005 , \46003 );
and \U$45629 ( \46006 , \46005 , \5016 );
nor \U$45630 ( \46007 , \46004 , \46006 );
and \U$45631 ( \46008 , \5896 , RIae75ce0_26);
and \U$45632 ( \46009 , RIae75dd0_28, \5894 );
nor \U$45633 ( \46010 , \46008 , \46009 );
and \U$45634 ( \46011 , \46010 , \5589 );
not \U$45635 ( \46012 , \46010 );
and \U$45636 ( \46013 , \46012 , \5590 );
nor \U$45637 ( \46014 , \46011 , \46013 );
or \U$45638 ( \46015 , \46007 , \46014 );
not \U$45639 ( \46016 , \46014 );
not \U$45640 ( \46017 , \46007 );
or \U$45641 ( \46018 , \46016 , \46017 );
and \U$45642 ( \46019 , \6172 , RIae75650_12);
and \U$45643 ( \46020 , RIae75560_10, \6170 );
nor \U$45644 ( \46021 , \46019 , \46020 );
and \U$45645 ( \46022 , \46021 , \6176 );
not \U$45646 ( \46023 , \46021 );
and \U$45647 ( \46024 , \46023 , \6175 );
nor \U$45648 ( \46025 , \46022 , \46024 );
nand \U$45649 ( \46026 , \46018 , \46025 );
nand \U$45650 ( \46027 , \46015 , \46026 );
xor \U$45651 ( \46028 , \46000 , \46027 );
and \U$45652 ( \46029 , \3730 , RIae78800_118);
and \U$45653 ( \46030 , RIae78710_116, \3728 );
nor \U$45654 ( \46031 , \46029 , \46030 );
and \U$45655 ( \46032 , \46031 , \3422 );
not \U$45656 ( \46033 , \46031 );
and \U$45657 ( \46034 , \46033 , \3732 );
nor \U$45658 ( \46035 , \46032 , \46034 );
and \U$45659 ( \46036 , \4247 , RIae75bf0_24);
and \U$45660 ( \46037 , RIae75b00_22, \4245 );
nor \U$45661 ( \46038 , \46036 , \46037 );
and \U$45662 ( \46039 , \46038 , \4251 );
not \U$45663 ( \46040 , \46038 );
and \U$45664 ( \46041 , \46040 , \3989 );
nor \U$45665 ( \46042 , \46039 , \46041 );
or \U$45666 ( \46043 , \46035 , \46042 );
not \U$45667 ( \46044 , \46042 );
not \U$45668 ( \46045 , \46035 );
or \U$45669 ( \46046 , \46044 , \46045 );
and \U$45670 ( \46047 , \4688 , RIae75a10_20);
and \U$45671 ( \46048 , RIae75920_18, \4686 );
nor \U$45672 ( \46049 , \46047 , \46048 );
and \U$45673 ( \46050 , \46049 , \4481 );
not \U$45674 ( \46051 , \46049 );
and \U$45675 ( \46052 , \46051 , \4482 );
nor \U$45676 ( \46053 , \46050 , \46052 );
nand \U$45677 ( \46054 , \46046 , \46053 );
nand \U$45678 ( \46055 , \46043 , \46054 );
and \U$45679 ( \46056 , \46028 , \46055 );
and \U$45680 ( \46057 , \46000 , \46027 );
or \U$45681 ( \46058 , \46056 , \46057 );
and \U$45682 ( \46059 , \2607 , RIae77cc0_94);
and \U$45683 ( \46060 , RIae77bd0_92, \2605 );
nor \U$45684 ( \46061 , \46059 , \46060 );
and \U$45685 ( \46062 , \46061 , \2397 );
not \U$45686 ( \46063 , \46061 );
and \U$45687 ( \46064 , \46063 , \2611 );
nor \U$45688 ( \46065 , \46062 , \46064 );
and \U$45689 ( \46066 , \2783 , RIae77db0_96);
and \U$45690 ( \46067 , RIae77ea0_98, \2781 );
nor \U$45691 ( \46068 , \46066 , \46067 );
not \U$45692 ( \46069 , \46068 );
not \U$45693 ( \46070 , \2789 );
and \U$45694 ( \46071 , \46069 , \46070 );
and \U$45695 ( \46072 , \46068 , \3089 );
nor \U$45696 ( \46073 , \46071 , \46072 );
or \U$45697 ( \46074 , \46065 , \46073 );
not \U$45698 ( \46075 , \46073 );
not \U$45699 ( \46076 , \46065 );
or \U$45700 ( \46077 , \46075 , \46076 );
not \U$45701 ( \46078 , \2774 );
and \U$45702 ( \46079 , \3214 , RIae789e0_122);
and \U$45703 ( \46080 , RIae788f0_120, \3212 );
nor \U$45704 ( \46081 , \46079 , \46080 );
not \U$45705 ( \46082 , \46081 );
or \U$45706 ( \46083 , \46078 , \46082 );
or \U$45707 ( \46084 , \46081 , \2774 );
nand \U$45708 ( \46085 , \46083 , \46084 );
nand \U$45709 ( \46086 , \46077 , \46085 );
nand \U$45710 ( \46087 , \46074 , \46086 );
and \U$45711 ( \46088 , \1939 , RIae78260_106);
and \U$45712 ( \46089 , RIae78620_114, \1937 );
nor \U$45713 ( \46090 , \46088 , \46089 );
and \U$45714 ( \46091 , \46090 , \1734 );
not \U$45715 ( \46092 , \46090 );
and \U$45716 ( \46093 , \46092 , \1735 );
nor \U$45717 ( \46094 , \46091 , \46093 );
and \U$45718 ( \46095 , \2224 , RIae78440_110);
and \U$45719 ( \46096 , RIae784b8_111, \2222 );
nor \U$45720 ( \46097 , \46095 , \46096 );
and \U$45721 ( \46098 , \46097 , \2060 );
not \U$45722 ( \46099 , \46097 );
and \U$45723 ( \46100 , \46099 , \2061 );
nor \U$45724 ( \46101 , \46098 , \46100 );
xor \U$45725 ( \46102 , \46094 , \46101 );
and \U$45726 ( \46103 , \1593 , RIae77f90_100);
and \U$45727 ( \46104 , RIae78080_102, \1591 );
nor \U$45728 ( \46105 , \46103 , \46104 );
and \U$45729 ( \46106 , \46105 , \1488 );
not \U$45730 ( \46107 , \46105 );
and \U$45731 ( \46108 , \46107 , \1498 );
nor \U$45732 ( \46109 , \46106 , \46108 );
and \U$45733 ( \46110 , \46102 , \46109 );
and \U$45734 ( \46111 , \46094 , \46101 );
nor \U$45735 ( \46112 , \46110 , \46111 );
xor \U$45736 ( \46113 , \46087 , \46112 );
and \U$45737 ( \46114 , \1138 , RIae77270_72);
and \U$45738 ( \46115 , RIae77360_74, \1136 );
nor \U$45739 ( \46116 , \46114 , \46115 );
and \U$45740 ( \46117 , \46116 , \1012 );
not \U$45741 ( \46118 , \46116 );
and \U$45742 ( \46119 , \46118 , \1142 );
nor \U$45743 ( \46120 , \46117 , \46119 );
not \U$45744 ( \46121 , \787 );
and \U$45745 ( \46122 , \883 , RIae77108_69);
and \U$45746 ( \46123 , RIae77090_68, \881 );
nor \U$45747 ( \46124 , \46122 , \46123 );
not \U$45748 ( \46125 , \46124 );
or \U$45749 ( \46126 , \46121 , \46125 );
or \U$45750 ( \46127 , \46124 , \789 );
nand \U$45751 ( \46128 , \46126 , \46127 );
xor \U$45752 ( \46129 , \46120 , \46128 );
and \U$45753 ( \46130 , \1376 , RIae78350_108);
and \U$45754 ( \46131 , RIae78170_104, \1374 );
nor \U$45755 ( \46132 , \46130 , \46131 );
and \U$45756 ( \46133 , \46132 , \1380 );
not \U$45757 ( \46134 , \46132 );
and \U$45758 ( \46135 , \46134 , \1261 );
nor \U$45759 ( \46136 , \46133 , \46135 );
and \U$45760 ( \46137 , \46129 , \46136 );
and \U$45761 ( \46138 , \46120 , \46128 );
or \U$45762 ( \46139 , \46137 , \46138 );
and \U$45763 ( \46140 , \46113 , \46139 );
and \U$45764 ( \46141 , \46087 , \46112 );
or \U$45765 ( \46142 , \46140 , \46141 );
xor \U$45766 ( \46143 , \46058 , \46142 );
and \U$45767 ( \46144 , \8966 , RIae76460_42);
and \U$45768 ( \46145 , RIae76550_44, \8964 );
nor \U$45769 ( \46146 , \46144 , \46145 );
and \U$45770 ( \46147 , \46146 , \8789 );
not \U$45771 ( \46148 , \46146 );
and \U$45772 ( \46149 , \46148 , \8799 );
nor \U$45773 ( \46150 , \46147 , \46149 );
and \U$45774 ( \46151 , \9760 , RIae76730_48);
and \U$45775 ( \46152 , RIae76640_46, \9758 );
nor \U$45776 ( \46153 , \46151 , \46152 );
and \U$45777 ( \46154 , \46153 , \9272 );
not \U$45778 ( \46155 , \46153 );
and \U$45779 ( \46156 , \46155 , \9273 );
nor \U$45780 ( \46157 , \46154 , \46156 );
xor \U$45781 ( \46158 , \46150 , \46157 );
and \U$45782 ( \46159 , \10548 , RIae76190_36);
and \U$45783 ( \46160 , RIae760a0_34, \10546 );
nor \U$45784 ( \46161 , \46159 , \46160 );
and \U$45785 ( \46162 , \46161 , \10118 );
not \U$45786 ( \46163 , \46161 );
and \U$45787 ( \46164 , \46163 , \10421 );
nor \U$45788 ( \46165 , \46162 , \46164 );
and \U$45789 ( \46166 , \46158 , \46165 );
and \U$45790 ( \46167 , \46150 , \46157 );
or \U$45791 ( \46168 , \46166 , \46167 );
and \U$45792 ( \46169 , \11470 , RIae76370_40);
and \U$45793 ( \46170 , RIae76280_38, \11468 );
nor \U$45794 ( \46171 , \46169 , \46170 );
and \U$45795 ( \46172 , \46171 , \11474 );
not \U$45796 ( \46173 , \46171 );
and \U$45797 ( \46174 , \46173 , \10936 );
nor \U$45798 ( \46175 , \46172 , \46174 );
not \U$45799 ( \46176 , \46175 );
and \U$45800 ( \46177 , \13059 , RIae76820_50);
and \U$45801 ( \46178 , RIae76910_52, \13057 );
nor \U$45802 ( \46179 , \46177 , \46178 );
and \U$45803 ( \46180 , \46179 , \12718 );
not \U$45804 ( \46181 , \46179 );
and \U$45805 ( \46182 , \46181 , \13063 );
nor \U$45806 ( \46183 , \46180 , \46182 );
not \U$45807 ( \46184 , \46183 );
and \U$45808 ( \46185 , \46176 , \46184 );
and \U$45809 ( \46186 , \46183 , \46175 );
and \U$45810 ( \46187 , \12180 , RIae76af0_56);
and \U$45811 ( \46188 , RIae76a00_54, \12178 );
nor \U$45812 ( \46189 , \46187 , \46188 );
and \U$45813 ( \46190 , \46189 , \11827 );
not \U$45814 ( \46191 , \46189 );
and \U$45815 ( \46192 , \46191 , \12184 );
nor \U$45816 ( \46193 , \46190 , \46192 );
nor \U$45817 ( \46194 , \46186 , \46193 );
nor \U$45818 ( \46195 , \46185 , \46194 );
or \U$45819 ( \46196 , \46168 , \46195 );
not \U$45820 ( \46197 , \46168 );
not \U$45821 ( \46198 , \46195 );
or \U$45822 ( \46199 , \46197 , \46198 );
and \U$45823 ( \46200 , \14059 , RIae76be0_58);
and \U$45824 ( \46201 , RIae78ad0_124, \14057 );
nor \U$45825 ( \46202 , \46200 , \46201 );
and \U$45826 ( \46203 , \46202 , \14063 );
not \U$45827 ( \46204 , \46202 );
and \U$45828 ( \46205 , \46204 , \13502 );
nor \U$45829 ( \46206 , \46203 , \46205 );
or \U$45830 ( \46207 , \46206 , RIae7aa38_191);
not \U$45831 ( \46208 , RIae7aa38_191);
not \U$45832 ( \46209 , \46206 );
or \U$45833 ( \46210 , \46208 , \46209 );
and \U$45834 ( \46211 , \14964 , RIae78d28_129);
and \U$45835 ( \46212 , RIae78e18_131, \14962 );
nor \U$45836 ( \46213 , \46211 , \46212 );
and \U$45837 ( \46214 , \46213 , \14463 );
not \U$45838 ( \46215 , \46213 );
and \U$45839 ( \46216 , \46215 , \14462 );
nor \U$45840 ( \46217 , \46214 , \46216 );
nand \U$45841 ( \46218 , \46210 , \46217 );
nand \U$45842 ( \46219 , \46207 , \46218 );
nand \U$45843 ( \46220 , \46199 , \46219 );
nand \U$45844 ( \46221 , \46196 , \46220 );
and \U$45845 ( \46222 , \46143 , \46221 );
and \U$45846 ( \46223 , \46058 , \46142 );
or \U$45847 ( \46224 , \46222 , \46223 );
xor \U$45848 ( \46225 , \45973 , \46224 );
and \U$45849 ( \46226 , \7633 , RIae751a0_2);
and \U$45850 ( \46227 , RIae75380_6, \7631 );
nor \U$45851 ( \46228 , \46226 , \46227 );
and \U$45852 ( \46229 , \46228 , \7206 );
not \U$45853 ( \46230 , \46228 );
and \U$45854 ( \46231 , \46230 , \7205 );
nor \U$45855 ( \46232 , \46229 , \46231 );
and \U$45856 ( \46233 , \6172 , RIae75560_10);
and \U$45857 ( \46234 , RIae75830_16, \6170 );
nor \U$45858 ( \46235 , \46233 , \46234 );
and \U$45859 ( \46236 , \46235 , \6176 );
not \U$45860 ( \46237 , \46235 );
and \U$45861 ( \46238 , \46237 , \6175 );
nor \U$45862 ( \46239 , \46236 , \46238 );
xor \U$45863 ( \46240 , \46232 , \46239 );
and \U$45864 ( \46241 , \6941 , RIae75740_14);
and \U$45865 ( \46242 , RIae75290_4, \6939 );
nor \U$45866 ( \46243 , \46241 , \46242 );
and \U$45867 ( \46244 , \46243 , \6314 );
not \U$45868 ( \46245 , \46243 );
and \U$45869 ( \46246 , \46245 , \6945 );
nor \U$45870 ( \46247 , \46244 , \46246 );
xor \U$45871 ( \46248 , \46240 , \46247 );
and \U$45872 ( \46249 , \10548 , RIae760a0_34);
and \U$45873 ( \46250 , RIae76370_40, \10546 );
nor \U$45874 ( \46251 , \46249 , \46250 );
and \U$45875 ( \46252 , \46251 , \10421 );
not \U$45876 ( \46253 , \46251 );
and \U$45877 ( \46254 , \46253 , \10118 );
nor \U$45878 ( \46255 , \46252 , \46254 );
and \U$45879 ( \46256 , \11470 , RIae76280_38);
and \U$45880 ( \46257 , RIae76af0_56, \11468 );
nor \U$45881 ( \46258 , \46256 , \46257 );
and \U$45882 ( \46259 , \46258 , \10936 );
not \U$45883 ( \46260 , \46258 );
and \U$45884 ( \46261 , \46260 , \11474 );
nor \U$45885 ( \46262 , \46259 , \46261 );
xor \U$45886 ( \46263 , \46255 , \46262 );
and \U$45887 ( \46264 , \12180 , RIae76a00_54);
and \U$45888 ( \46265 , RIae76820_50, \12178 );
nor \U$45889 ( \46266 , \46264 , \46265 );
and \U$45890 ( \46267 , \46266 , \12184 );
not \U$45891 ( \46268 , \46266 );
and \U$45892 ( \46269 , \46268 , \11827 );
nor \U$45893 ( \46270 , \46267 , \46269 );
xor \U$45894 ( \46271 , \46263 , \46270 );
and \U$45895 ( \46272 , \46248 , \46271 );
and \U$45896 ( \46273 , \8966 , RIae76550_44);
and \U$45897 ( \46274 , RIae76730_48, \8964 );
nor \U$45898 ( \46275 , \46273 , \46274 );
and \U$45899 ( \46276 , \46275 , \8799 );
not \U$45900 ( \46277 , \46275 );
and \U$45901 ( \46278 , \46277 , \8789 );
nor \U$45902 ( \46279 , \46276 , \46278 );
and \U$45903 ( \46280 , \8371 , RIae75470_8);
and \U$45904 ( \46281 , RIae76460_42, \8369 );
nor \U$45905 ( \46282 , \46280 , \46281 );
and \U$45906 ( \46283 , \46282 , \8020 );
not \U$45907 ( \46284 , \46282 );
and \U$45908 ( \46285 , \46284 , \8019 );
nor \U$45909 ( \46286 , \46283 , \46285 );
xor \U$45910 ( \46287 , \46279 , \46286 );
and \U$45911 ( \46288 , \9760 , RIae76640_46);
and \U$45912 ( \46289 , RIae76190_36, \9758 );
nor \U$45913 ( \46290 , \46288 , \46289 );
and \U$45914 ( \46291 , \46290 , \9273 );
not \U$45915 ( \46292 , \46290 );
and \U$45916 ( \46293 , \46292 , \9272 );
nor \U$45917 ( \46294 , \46291 , \46293 );
xor \U$45918 ( \46295 , \46287 , \46294 );
xor \U$45919 ( \46296 , \46255 , \46262 );
xor \U$45920 ( \46297 , \46296 , \46270 );
and \U$45921 ( \46298 , \46295 , \46297 );
and \U$45922 ( \46299 , \46248 , \46295 );
or \U$45923 ( \46300 , \46272 , \46298 , \46299 );
xor \U$45924 ( \46301 , \45760 , \45762 );
xor \U$45925 ( \46302 , \46300 , \46301 );
xor \U$45926 ( \46303 , \45520 , \45527 );
xor \U$45927 ( \46304 , \46303 , \45535 );
xor \U$45928 ( \46305 , \45748 , \45753 );
xor \U$45929 ( \46306 , \46304 , \46305 );
and \U$45930 ( \46307 , \46302 , \46306 );
and \U$45931 ( \46308 , \46300 , \46301 );
or \U$45932 ( \46309 , \46307 , \46308 );
and \U$45933 ( \46310 , \46225 , \46309 );
and \U$45934 ( \46311 , \45973 , \46224 );
or \U$45935 ( \46312 , \46310 , \46311 );
xor \U$45936 ( \46313 , \45785 , \46312 );
xor \U$45937 ( \46314 , \45695 , \45703 );
xor \U$45938 ( \46315 , \46314 , \45731 );
xor \U$45939 ( \46316 , \45737 , \45739 );
xor \U$45940 ( \46317 , \46316 , \45742 );
and \U$45941 ( \46318 , \46315 , \46317 );
xor \U$45942 ( \46319 , \45320 , \45328 );
xor \U$45943 ( \46320 , \46319 , \45336 );
xor \U$45944 ( \46321 , \45675 , \45680 );
xor \U$45945 ( \46322 , \46320 , \46321 );
xor \U$45946 ( \46323 , \45737 , \45739 );
xor \U$45947 ( \46324 , \46323 , \45742 );
and \U$45948 ( \46325 , \46322 , \46324 );
and \U$45949 ( \46326 , \46315 , \46322 );
or \U$45950 ( \46327 , \46318 , \46325 , \46326 );
xor \U$45951 ( \46328 , \46255 , \46262 );
and \U$45952 ( \46329 , \46328 , \46270 );
and \U$45953 ( \46330 , \46255 , \46262 );
or \U$45954 ( \46331 , \46329 , \46330 );
and \U$45955 ( \46332 , \13059 , RIae76910_52);
and \U$45956 ( \46333 , RIae76be0_58, \13057 );
nor \U$45957 ( \46334 , \46332 , \46333 );
and \U$45958 ( \46335 , \46334 , \13063 );
not \U$45959 ( \46336 , \46334 );
and \U$45960 ( \46337 , \46336 , \12718 );
nor \U$45961 ( \46338 , \46335 , \46337 );
nand \U$45962 ( \46339 , RIae78e18_131, \14964 );
and \U$45963 ( \46340 , \46339 , \14463 );
not \U$45964 ( \46341 , \46339 );
and \U$45965 ( \46342 , \46341 , \14462 );
nor \U$45966 ( \46343 , \46340 , \46342 );
xor \U$45967 ( \46344 , \46338 , \46343 );
and \U$45968 ( \46345 , \14059 , RIae78ad0_124);
and \U$45969 ( \46346 , RIae78d28_129, \14057 );
nor \U$45970 ( \46347 , \46345 , \46346 );
and \U$45971 ( \46348 , \46347 , \13502 );
not \U$45972 ( \46349 , \46347 );
and \U$45973 ( \46350 , \46349 , \14063 );
nor \U$45974 ( \46351 , \46348 , \46350 );
and \U$45975 ( \46352 , \46344 , \46351 );
and \U$45976 ( \46353 , \46338 , \46343 );
or \U$45977 ( \46354 , \46352 , \46353 );
xor \U$45978 ( \46355 , \46331 , \46354 );
xor \U$45979 ( \46356 , \46279 , \46286 );
and \U$45980 ( \46357 , \46356 , \46294 );
and \U$45981 ( \46358 , \46279 , \46286 );
or \U$45982 ( \46359 , \46357 , \46358 );
xor \U$45983 ( \46360 , \46355 , \46359 );
xor \U$45984 ( \46361 , \45841 , \45848 );
and \U$45985 ( \46362 , \46361 , \45856 );
and \U$45986 ( \46363 , \45841 , \45848 );
or \U$45987 ( \46364 , \46362 , \46363 );
xor \U$45988 ( \46365 , \45816 , \45824 );
and \U$45989 ( \46366 , \46365 , \45832 );
and \U$45990 ( \46367 , \45816 , \45824 );
or \U$45991 ( \46368 , \46366 , \46367 );
xor \U$45992 ( \46369 , \46364 , \46368 );
xor \U$45993 ( \46370 , \46232 , \46239 );
and \U$45994 ( \46371 , \46370 , \46247 );
and \U$45995 ( \46372 , \46232 , \46239 );
or \U$45996 ( \46373 , \46371 , \46372 );
xor \U$45997 ( \46374 , \46369 , \46373 );
and \U$45998 ( \46375 , \46360 , \46374 );
xor \U$45999 ( \46376 , \45949 , \45956 );
and \U$46000 ( \46377 , \46376 , \45964 );
and \U$46001 ( \46378 , \45949 , \45956 );
or \U$46002 ( \46379 , \46377 , \46378 );
xor \U$46003 ( \46380 , \45922 , \45929 );
and \U$46004 ( \46381 , \46380 , \45938 );
and \U$46005 ( \46382 , \45922 , \45929 );
or \U$46006 ( \46383 , \46381 , \46382 );
xor \U$46007 ( \46384 , \46379 , \46383 );
xor \U$46008 ( \46385 , \45793 , \45800 );
and \U$46009 ( \46386 , \46385 , \45808 );
and \U$46010 ( \46387 , \45793 , \45800 );
or \U$46011 ( \46388 , \46386 , \46387 );
xor \U$46012 ( \46389 , \46384 , \46388 );
xor \U$46013 ( \46390 , \46364 , \46368 );
xor \U$46014 ( \46391 , \46390 , \46373 );
and \U$46015 ( \46392 , \46389 , \46391 );
and \U$46016 ( \46393 , \46360 , \46389 );
or \U$46017 ( \46394 , \46375 , \46392 , \46393 );
xor \U$46018 ( \46395 , \46327 , \46394 );
xor \U$46019 ( \46396 , \45385 , \45410 );
xor \U$46020 ( \46397 , \46396 , \45437 );
xor \U$46021 ( \46398 , \45465 , \45483 );
xor \U$46022 ( \46399 , \46398 , \45509 );
xor \U$46023 ( \46400 , \45538 , \45563 );
xor \U$46024 ( \46401 , \46400 , \45590 );
xor \U$46025 ( \46402 , \46399 , \46401 );
xor \U$46026 ( \46403 , \46397 , \46402 );
and \U$46027 ( \46404 , \46395 , \46403 );
and \U$46028 ( \46405 , \46327 , \46394 );
or \U$46029 ( \46406 , \46404 , \46405 );
and \U$46030 ( \46407 , \46313 , \46406 );
and \U$46031 ( \46408 , \45785 , \46312 );
or \U$46032 ( \46409 , \46407 , \46408 );
xor \U$46033 ( \46410 , \45280 , \45282 );
xor \U$46034 ( \46411 , \46410 , \45297 );
xor \U$46035 ( \46412 , \46409 , \46411 );
xor \U$46036 ( \46413 , \45440 , \45512 );
xor \U$46037 ( \46414 , \46413 , \45593 );
xor \U$46038 ( \46415 , \45348 , \45350 );
xor \U$46039 ( \46416 , \46415 , \45353 );
and \U$46040 ( \46417 , \45774 , \46416 );
xor \U$46041 ( \46418 , \45348 , \45350 );
xor \U$46042 ( \46419 , \46418 , \45353 );
and \U$46043 ( \46420 , \45778 , \46419 );
and \U$46044 ( \46421 , \45774 , \45778 );
or \U$46045 ( \46422 , \46417 , \46420 , \46421 );
xor \U$46046 ( \46423 , \45385 , \45410 );
xor \U$46047 ( \46424 , \46423 , \45437 );
and \U$46048 ( \46425 , \46399 , \46424 );
xor \U$46049 ( \46426 , \45385 , \45410 );
xor \U$46050 ( \46427 , \46426 , \45437 );
and \U$46051 ( \46428 , \46401 , \46427 );
and \U$46052 ( \46429 , \46399 , \46401 );
or \U$46053 ( \46430 , \46425 , \46428 , \46429 );
xor \U$46054 ( \46431 , \46422 , \46430 );
xor \U$46055 ( \46432 , \44945 , \44970 );
xor \U$46056 ( \46433 , \46432 , \44997 );
xor \U$46057 ( \46434 , \45270 , \45275 );
xor \U$46058 ( \46435 , \46433 , \46434 );
xor \U$46059 ( \46436 , \46431 , \46435 );
and \U$46060 ( \46437 , \46414 , \46436 );
xor \U$46061 ( \46438 , \45312 , \45345 );
xor \U$46062 ( \46439 , \46438 , \45356 );
xor \U$46063 ( \46440 , \45609 , \45611 );
xor \U$46064 ( \46441 , \46440 , \45616 );
xor \U$46065 ( \46442 , \44856 , \44858 );
xor \U$46066 ( \46443 , \46442 , \44861 );
xor \U$46067 ( \46444 , \45285 , \45292 );
xor \U$46068 ( \46445 , \46443 , \46444 );
xor \U$46069 ( \46446 , \46441 , \46445 );
xor \U$46070 ( \46447 , \46439 , \46446 );
xor \U$46071 ( \46448 , \46422 , \46430 );
xor \U$46072 ( \46449 , \46448 , \46435 );
and \U$46073 ( \46450 , \46447 , \46449 );
and \U$46074 ( \46451 , \46414 , \46447 );
or \U$46075 ( \46452 , \46437 , \46450 , \46451 );
and \U$46076 ( \46453 , \46412 , \46452 );
and \U$46077 ( \46454 , \46409 , \46411 );
or \U$46078 ( \46455 , \46453 , \46454 );
xor \U$46079 ( \46456 , \45300 , \45622 );
xor \U$46080 ( \46457 , \46456 , \45637 );
xor \U$46081 ( \46458 , \46455 , \46457 );
xor \U$46082 ( \46459 , \44864 , \44900 );
xor \U$46083 ( \46460 , \46459 , \44917 );
xor \U$46084 ( \46461 , \45000 , \45077 );
xor \U$46085 ( \46462 , \46461 , \45159 );
xor \U$46086 ( \46463 , \45197 , \45199 );
xor \U$46087 ( \46464 , \46463 , \45204 );
xor \U$46088 ( \46465 , \45625 , \45632 );
xor \U$46089 ( \46466 , \46464 , \46465 );
xor \U$46090 ( \46467 , \46462 , \46466 );
xor \U$46091 ( \46468 , \46460 , \46467 );
xor \U$46092 ( \46469 , \45359 , \45596 );
xor \U$46093 ( \46470 , \46469 , \45619 );
xor \U$46094 ( \46471 , \46468 , \46470 );
xor \U$46095 ( \46472 , \46422 , \46430 );
and \U$46096 ( \46473 , \46472 , \46435 );
and \U$46097 ( \46474 , \46422 , \46430 );
or \U$46098 ( \46475 , \46473 , \46474 );
xor \U$46099 ( \46476 , \45685 , \45734 );
and \U$46100 ( \46477 , \46476 , \45745 );
and \U$46101 ( \46478 , \45685 , \45734 );
or \U$46102 ( \46479 , \46477 , \46478 );
xor \U$46103 ( \46480 , \46364 , \46368 );
and \U$46104 ( \46481 , \46480 , \46373 );
and \U$46105 ( \46482 , \46364 , \46368 );
or \U$46106 ( \46483 , \46481 , \46482 );
xor \U$46107 ( \46484 , \46379 , \46383 );
and \U$46108 ( \46485 , \46484 , \46388 );
and \U$46109 ( \46486 , \46379 , \46383 );
or \U$46110 ( \46487 , \46485 , \46486 );
xor \U$46111 ( \46488 , \46483 , \46487 );
xor \U$46112 ( \46489 , \46331 , \46354 );
and \U$46113 ( \46490 , \46489 , \46359 );
and \U$46114 ( \46491 , \46331 , \46354 );
or \U$46115 ( \46492 , \46490 , \46491 );
and \U$46116 ( \46493 , \46488 , \46492 );
and \U$46117 ( \46494 , \46483 , \46487 );
or \U$46118 ( \46495 , \46493 , \46494 );
xor \U$46119 ( \46496 , \46479 , \46495 );
xor \U$46120 ( \46497 , \45758 , \45763 );
and \U$46121 ( \46498 , \46497 , \45768 );
and \U$46122 ( \46499 , \45758 , \45763 );
or \U$46123 ( \46500 , \46498 , \46499 );
and \U$46124 ( \46501 , \46496 , \46500 );
and \U$46125 ( \46502 , \46479 , \46495 );
or \U$46126 ( \46503 , \46501 , \46502 );
xor \U$46127 ( \46504 , \46475 , \46503 );
xor \U$46128 ( \46505 , \45312 , \45345 );
xor \U$46129 ( \46506 , \46505 , \45356 );
and \U$46130 ( \46507 , \46441 , \46506 );
xor \U$46131 ( \46508 , \45312 , \45345 );
xor \U$46132 ( \46509 , \46508 , \45356 );
and \U$46133 ( \46510 , \46445 , \46509 );
and \U$46134 ( \46511 , \46441 , \46445 );
or \U$46135 ( \46512 , \46507 , \46510 , \46511 );
xor \U$46136 ( \46513 , \46504 , \46512 );
and \U$46137 ( \46514 , \46471 , \46513 );
and \U$46138 ( \46515 , \46468 , \46470 );
or \U$46139 ( \46516 , \46514 , \46515 );
and \U$46140 ( \46517 , \46458 , \46516 );
and \U$46141 ( \46518 , \46455 , \46457 );
or \U$46142 ( \46519 , \46517 , \46518 );
xor \U$46143 ( \46520 , \45640 , \45642 );
xor \U$46144 ( \46521 , \46520 , \45657 );
xor \U$46145 ( \46522 , \46475 , \46503 );
and \U$46146 ( \46523 , \46522 , \46512 );
and \U$46147 ( \46524 , \46475 , \46503 );
or \U$46148 ( \46525 , \46523 , \46524 );
xor \U$46149 ( \46526 , \44864 , \44900 );
xor \U$46150 ( \46527 , \46526 , \44917 );
and \U$46151 ( \46528 , \46462 , \46527 );
xor \U$46152 ( \46529 , \44864 , \44900 );
xor \U$46153 ( \46530 , \46529 , \44917 );
and \U$46154 ( \46531 , \46466 , \46530 );
and \U$46155 ( \46532 , \46462 , \46466 );
or \U$46156 ( \46533 , \46528 , \46531 , \46532 );
xor \U$46157 ( \46534 , \46525 , \46533 );
xor \U$46158 ( \46535 , \45195 , \45207 );
xor \U$46159 ( \46536 , \46535 , \45212 );
xor \U$46160 ( \46537 , \45645 , \45652 );
xor \U$46161 ( \46538 , \46536 , \46537 );
and \U$46162 ( \46539 , \46534 , \46538 );
and \U$46163 ( \46540 , \46525 , \46533 );
or \U$46164 ( \46541 , \46539 , \46540 );
xor \U$46165 ( \46542 , \45220 , \45222 );
xor \U$46166 ( \46543 , \46542 , \45227 );
xor \U$46167 ( \46544 , \45257 , \45262 );
xor \U$46168 ( \46545 , \46543 , \46544 );
xor \U$46169 ( \46546 , \46541 , \46545 );
xor \U$46170 ( \46547 , \46521 , \46546 );
and \U$46171 ( \46548 , \46519 , \46547 );
not \U$46172 ( \46549 , \46548 );
xor \U$46173 ( \46550 , \45640 , \45642 );
xor \U$46174 ( \46551 , \46550 , \45657 );
and \U$46175 ( \46552 , \46541 , \46551 );
xor \U$46176 ( \46553 , \45640 , \45642 );
xor \U$46177 ( \46554 , \46553 , \45657 );
and \U$46178 ( \46555 , \46545 , \46554 );
and \U$46179 ( \46556 , \46541 , \46545 );
or \U$46180 ( \46557 , \46552 , \46555 , \46556 );
xor \U$46181 ( \46558 , \45218 , \45230 );
xor \U$46182 ( \46559 , \46558 , \45235 );
xor \U$46183 ( \46560 , \46557 , \46559 );
xor \U$46184 ( \46561 , \45255 , \45267 );
xor \U$46185 ( \46562 , \46561 , \45660 );
xor \U$46186 ( \46563 , \46560 , \46562 );
not \U$46187 ( \46564 , \46563 );
or \U$46188 ( \46565 , \46549 , \46564 );
xor \U$46189 ( \46566 , \45711 , \45719 );
xor \U$46190 ( \46567 , \46566 , \45728 );
xor \U$46191 ( \46568 , \45939 , \45965 );
xor \U$46192 ( \46569 , \46567 , \46568 );
xor \U$46193 ( \46570 , \45809 , \45833 );
xor \U$46194 ( \46571 , \46570 , \45857 );
and \U$46195 ( \46572 , \46569 , \46571 );
xor \U$46196 ( \46573 , \46255 , \46262 );
xor \U$46197 ( \46574 , \46573 , \46270 );
xor \U$46198 ( \46575 , \46248 , \46295 );
xor \U$46199 ( \46576 , \46574 , \46575 );
xor \U$46200 ( \46577 , \45809 , \45833 );
xor \U$46201 ( \46578 , \46577 , \45857 );
and \U$46202 ( \46579 , \46576 , \46578 );
and \U$46203 ( \46580 , \46569 , \46576 );
or \U$46204 ( \46581 , \46572 , \46579 , \46580 );
xor \U$46205 ( \46582 , \46000 , \46027 );
xor \U$46206 ( \46583 , \46582 , \46055 );
xor \U$46207 ( \46584 , \46087 , \46112 );
xor \U$46208 ( \46585 , \46584 , \46139 );
xor \U$46209 ( \46586 , \46583 , \46585 );
xor \U$46210 ( \46587 , \45882 , \45884 );
xor \U$46211 ( \46588 , \46587 , \45911 );
and \U$46212 ( \46589 , \46586 , \46588 );
and \U$46213 ( \46590 , \46583 , \46585 );
or \U$46214 ( \46591 , \46589 , \46590 );
xor \U$46215 ( \46592 , \46581 , \46591 );
xor \U$46216 ( \46593 , \46364 , \46368 );
xor \U$46217 ( \46594 , \46593 , \46373 );
xor \U$46218 ( \46595 , \46360 , \46389 );
xor \U$46219 ( \46596 , \46594 , \46595 );
and \U$46220 ( \46597 , \46592 , \46596 );
and \U$46221 ( \46598 , \46581 , \46591 );
or \U$46222 ( \46599 , \46597 , \46598 );
and \U$46223 ( \46600 , \1593 , RIae78170_104);
and \U$46224 ( \46601 , RIae77f90_100, \1591 );
nor \U$46225 ( \46602 , \46600 , \46601 );
and \U$46226 ( \46603 , \46602 , \1488 );
not \U$46227 ( \46604 , \46602 );
and \U$46228 ( \46605 , \46604 , \1498 );
nor \U$46229 ( \46606 , \46603 , \46605 );
and \U$46230 ( \46607 , \1138 , RIae77090_68);
and \U$46231 ( \46608 , RIae77270_72, \1136 );
nor \U$46232 ( \46609 , \46607 , \46608 );
and \U$46233 ( \46610 , \46609 , \1142 );
not \U$46234 ( \46611 , \46609 );
and \U$46235 ( \46612 , \46611 , \1012 );
nor \U$46236 ( \46613 , \46610 , \46612 );
xor \U$46237 ( \46614 , \46606 , \46613 );
and \U$46238 ( \46615 , \1376 , RIae77360_74);
and \U$46239 ( \46616 , RIae78350_108, \1374 );
nor \U$46240 ( \46617 , \46615 , \46616 );
and \U$46241 ( \46618 , \46617 , \1261 );
not \U$46242 ( \46619 , \46617 );
and \U$46243 ( \46620 , \46619 , \1380 );
nor \U$46244 ( \46621 , \46618 , \46620 );
and \U$46245 ( \46622 , \46614 , \46621 );
and \U$46246 ( \46623 , \46606 , \46613 );
or \U$46247 ( \46624 , \46622 , \46623 );
and \U$46248 ( \46625 , \2607 , RIae784b8_111);
and \U$46249 ( \46626 , RIae77cc0_94, \2605 );
nor \U$46250 ( \46627 , \46625 , \46626 );
and \U$46251 ( \46628 , \46627 , \2397 );
not \U$46252 ( \46629 , \46627 );
and \U$46253 ( \46630 , \46629 , \2611 );
nor \U$46254 ( \46631 , \46628 , \46630 );
and \U$46255 ( \46632 , \1939 , RIae78080_102);
and \U$46256 ( \46633 , RIae78260_106, \1937 );
nor \U$46257 ( \46634 , \46632 , \46633 );
and \U$46258 ( \46635 , \46634 , \1734 );
not \U$46259 ( \46636 , \46634 );
and \U$46260 ( \46637 , \46636 , \1735 );
nor \U$46261 ( \46638 , \46635 , \46637 );
xor \U$46262 ( \46639 , \46631 , \46638 );
and \U$46263 ( \46640 , \2224 , RIae78620_114);
and \U$46264 ( \46641 , RIae78440_110, \2222 );
nor \U$46265 ( \46642 , \46640 , \46641 );
and \U$46266 ( \46643 , \46642 , \2060 );
not \U$46267 ( \46644 , \46642 );
and \U$46268 ( \46645 , \46644 , \2061 );
nor \U$46269 ( \46646 , \46643 , \46645 );
and \U$46270 ( \46647 , \46639 , \46646 );
and \U$46271 ( \46648 , \46631 , \46638 );
or \U$46272 ( \46649 , \46647 , \46648 );
xor \U$46273 ( \46650 , \46624 , \46649 );
and \U$46274 ( \46651 , \3214 , RIae77ea0_98);
and \U$46275 ( \46652 , RIae789e0_122, \3212 );
nor \U$46276 ( \46653 , \46651 , \46652 );
not \U$46277 ( \46654 , \46653 );
not \U$46278 ( \46655 , \3218 );
and \U$46279 ( \46656 , \46654 , \46655 );
and \U$46280 ( \46657 , \46653 , \3218 );
nor \U$46281 ( \46658 , \46656 , \46657 );
and \U$46282 ( \46659 , \2783 , RIae77bd0_92);
and \U$46283 ( \46660 , RIae77db0_96, \2781 );
nor \U$46284 ( \46661 , \46659 , \46660 );
not \U$46285 ( \46662 , \46661 );
not \U$46286 ( \46663 , \3089 );
and \U$46287 ( \46664 , \46662 , \46663 );
and \U$46288 ( \46665 , \46661 , \2789 );
nor \U$46289 ( \46666 , \46664 , \46665 );
xor \U$46290 ( \46667 , \46658 , \46666 );
and \U$46291 ( \46668 , \3730 , RIae788f0_120);
and \U$46292 ( \46669 , RIae78800_118, \3728 );
nor \U$46293 ( \46670 , \46668 , \46669 );
and \U$46294 ( \46671 , \46670 , \3422 );
not \U$46295 ( \46672 , \46670 );
and \U$46296 ( \46673 , \46672 , \3732 );
nor \U$46297 ( \46674 , \46671 , \46673 );
and \U$46298 ( \46675 , \46667 , \46674 );
and \U$46299 ( \46676 , \46658 , \46666 );
or \U$46300 ( \46677 , \46675 , \46676 );
and \U$46301 ( \46678 , \46650 , \46677 );
and \U$46302 ( \46679 , \46624 , \46649 );
nor \U$46303 ( \46680 , \46678 , \46679 );
and \U$46304 ( \46681 , \14059 , RIae76910_52);
and \U$46305 ( \46682 , RIae76be0_58, \14057 );
nor \U$46306 ( \46683 , \46681 , \46682 );
and \U$46307 ( \46684 , \46683 , \14063 );
not \U$46308 ( \46685 , \46683 );
and \U$46309 ( \46686 , \46685 , \13502 );
nor \U$46310 ( \46687 , \46684 , \46686 );
and \U$46311 ( \46688 , \12180 , RIae76280_38);
and \U$46312 ( \46689 , RIae76af0_56, \12178 );
nor \U$46313 ( \46690 , \46688 , \46689 );
and \U$46314 ( \46691 , \46690 , \11827 );
not \U$46315 ( \46692 , \46690 );
and \U$46316 ( \46693 , \46692 , \12184 );
nor \U$46317 ( \46694 , \46691 , \46693 );
xor \U$46318 ( \46695 , \46687 , \46694 );
and \U$46319 ( \46696 , \13059 , RIae76a00_54);
and \U$46320 ( \46697 , RIae76820_50, \13057 );
nor \U$46321 ( \46698 , \46696 , \46697 );
and \U$46322 ( \46699 , \46698 , \12718 );
not \U$46323 ( \46700 , \46698 );
and \U$46324 ( \46701 , \46700 , \13063 );
nor \U$46325 ( \46702 , \46699 , \46701 );
and \U$46326 ( \46703 , \46695 , \46702 );
and \U$46327 ( \46704 , \46687 , \46694 );
or \U$46328 ( \46705 , \46703 , \46704 );
and \U$46329 ( \46706 , \14964 , RIae78ad0_124);
and \U$46330 ( \46707 , RIae78d28_129, \14962 );
nor \U$46331 ( \46708 , \46706 , \46707 );
and \U$46332 ( \46709 , \46708 , \14462 );
not \U$46333 ( \46710 , \46708 );
and \U$46334 ( \46711 , \46710 , \14463 );
nor \U$46335 ( \46712 , \46709 , \46711 );
not \U$46336 ( \46713 , \46712 );
and \U$46337 ( \46714 , \15726 , RIae78e18_131);
nor \U$46338 ( \46715 , \46714 , \14959 );
nand \U$46339 ( \46716 , \46713 , \46715 );
or \U$46340 ( \46717 , \46705 , \46716 );
not \U$46341 ( \46718 , \46716 );
not \U$46342 ( \46719 , \46705 );
or \U$46343 ( \46720 , \46718 , \46719 );
and \U$46344 ( \46721 , \9760 , RIae76550_44);
and \U$46345 ( \46722 , RIae76730_48, \9758 );
nor \U$46346 ( \46723 , \46721 , \46722 );
and \U$46347 ( \46724 , \46723 , \9272 );
not \U$46348 ( \46725 , \46723 );
and \U$46349 ( \46726 , \46725 , \9273 );
nor \U$46350 ( \46727 , \46724 , \46726 );
and \U$46351 ( \46728 , \11470 , RIae760a0_34);
and \U$46352 ( \46729 , RIae76370_40, \11468 );
nor \U$46353 ( \46730 , \46728 , \46729 );
and \U$46354 ( \46731 , \46730 , \11474 );
not \U$46355 ( \46732 , \46730 );
and \U$46356 ( \46733 , \46732 , \10936 );
nor \U$46357 ( \46734 , \46731 , \46733 );
or \U$46358 ( \46735 , \46727 , \46734 );
not \U$46359 ( \46736 , \46734 );
not \U$46360 ( \46737 , \46727 );
or \U$46361 ( \46738 , \46736 , \46737 );
and \U$46362 ( \46739 , \10548 , RIae76640_46);
and \U$46363 ( \46740 , RIae76190_36, \10546 );
nor \U$46364 ( \46741 , \46739 , \46740 );
and \U$46365 ( \46742 , \46741 , \10421 );
not \U$46366 ( \46743 , \46741 );
and \U$46367 ( \46744 , \46743 , \10118 );
nor \U$46368 ( \46745 , \46742 , \46744 );
nand \U$46369 ( \46746 , \46738 , \46745 );
nand \U$46370 ( \46747 , \46735 , \46746 );
nand \U$46371 ( \46748 , \46720 , \46747 );
nand \U$46372 ( \46749 , \46717 , \46748 );
xor \U$46373 ( \46750 , \46680 , \46749 );
and \U$46374 ( \46751 , \4688 , RIae75b00_22);
and \U$46375 ( \46752 , RIae75a10_20, \4686 );
nor \U$46376 ( \46753 , \46751 , \46752 );
and \U$46377 ( \46754 , \46753 , \4482 );
not \U$46378 ( \46755 , \46753 );
and \U$46379 ( \46756 , \46755 , \4481 );
nor \U$46380 ( \46757 , \46754 , \46756 );
and \U$46381 ( \46758 , \4247 , RIae78710_116);
and \U$46382 ( \46759 , RIae75bf0_24, \4245 );
nor \U$46383 ( \46760 , \46758 , \46759 );
and \U$46384 ( \46761 , \46760 , \4251 );
not \U$46385 ( \46762 , \46760 );
and \U$46386 ( \46763 , \46762 , \3989 );
nor \U$46387 ( \46764 , \46761 , \46763 );
xor \U$46388 ( \46765 , \46757 , \46764 );
and \U$46389 ( \46766 , \5399 , RIae75920_18);
and \U$46390 ( \46767 , RIae75fb0_32, \5397 );
nor \U$46391 ( \46768 , \46766 , \46767 );
and \U$46392 ( \46769 , \46768 , \5403 );
not \U$46393 ( \46770 , \46768 );
and \U$46394 ( \46771 , \46770 , \5016 );
nor \U$46395 ( \46772 , \46769 , \46771 );
and \U$46396 ( \46773 , \46765 , \46772 );
and \U$46397 ( \46774 , \46757 , \46764 );
or \U$46398 ( \46775 , \46773 , \46774 );
and \U$46399 ( \46776 , \6941 , RIae75560_10);
and \U$46400 ( \46777 , RIae75830_16, \6939 );
nor \U$46401 ( \46778 , \46776 , \46777 );
and \U$46402 ( \46779 , \46778 , \6945 );
not \U$46403 ( \46780 , \46778 );
and \U$46404 ( \46781 , \46780 , \6314 );
nor \U$46405 ( \46782 , \46779 , \46781 );
and \U$46406 ( \46783 , \5896 , RIae75ec0_30);
and \U$46407 ( \46784 , RIae75ce0_26, \5894 );
nor \U$46408 ( \46785 , \46783 , \46784 );
and \U$46409 ( \46786 , \46785 , \5589 );
not \U$46410 ( \46787 , \46785 );
and \U$46411 ( \46788 , \46787 , \5590 );
nor \U$46412 ( \46789 , \46786 , \46788 );
xor \U$46413 ( \46790 , \46782 , \46789 );
and \U$46414 ( \46791 , \6172 , RIae75dd0_28);
and \U$46415 ( \46792 , RIae75650_12, \6170 );
nor \U$46416 ( \46793 , \46791 , \46792 );
and \U$46417 ( \46794 , \46793 , \6175 );
not \U$46418 ( \46795 , \46793 );
and \U$46419 ( \46796 , \46795 , \6176 );
nor \U$46420 ( \46797 , \46794 , \46796 );
and \U$46421 ( \46798 , \46790 , \46797 );
and \U$46422 ( \46799 , \46782 , \46789 );
or \U$46423 ( \46800 , \46798 , \46799 );
xor \U$46424 ( \46801 , \46775 , \46800 );
and \U$46425 ( \46802 , \8371 , RIae751a0_2);
and \U$46426 ( \46803 , RIae75380_6, \8369 );
nor \U$46427 ( \46804 , \46802 , \46803 );
and \U$46428 ( \46805 , \46804 , \8019 );
not \U$46429 ( \46806 , \46804 );
and \U$46430 ( \46807 , \46806 , \8020 );
nor \U$46431 ( \46808 , \46805 , \46807 );
and \U$46432 ( \46809 , \7633 , RIae75740_14);
and \U$46433 ( \46810 , RIae75290_4, \7631 );
nor \U$46434 ( \46811 , \46809 , \46810 );
and \U$46435 ( \46812 , \46811 , \7205 );
not \U$46436 ( \46813 , \46811 );
and \U$46437 ( \46814 , \46813 , \7206 );
nor \U$46438 ( \46815 , \46812 , \46814 );
xor \U$46439 ( \46816 , \46808 , \46815 );
and \U$46440 ( \46817 , \8966 , RIae75470_8);
and \U$46441 ( \46818 , RIae76460_42, \8964 );
nor \U$46442 ( \46819 , \46817 , \46818 );
and \U$46443 ( \46820 , \46819 , \8789 );
not \U$46444 ( \46821 , \46819 );
and \U$46445 ( \46822 , \46821 , \8799 );
nor \U$46446 ( \46823 , \46820 , \46822 );
and \U$46447 ( \46824 , \46816 , \46823 );
and \U$46448 ( \46825 , \46808 , \46815 );
or \U$46449 ( \46826 , \46824 , \46825 );
and \U$46450 ( \46827 , \46801 , \46826 );
and \U$46451 ( \46828 , \46775 , \46800 );
nor \U$46452 ( \46829 , \46827 , \46828 );
and \U$46453 ( \46830 , \46750 , \46829 );
and \U$46454 ( \46831 , \46680 , \46749 );
or \U$46455 ( \46832 , \46830 , \46831 );
not \U$46456 ( \46833 , \46175 );
xor \U$46457 ( \46834 , \46193 , \46183 );
not \U$46458 ( \46835 , \46834 );
or \U$46459 ( \46836 , \46833 , \46835 );
or \U$46460 ( \46837 , \46834 , \46175 );
nand \U$46461 ( \46838 , \46836 , \46837 );
not \U$46462 ( \46839 , \46838 );
and \U$46463 ( \46840 , \46217 , \14959 );
not \U$46464 ( \46841 , \46217 );
and \U$46465 ( \46842 , \46841 , RIae7aa38_191);
nor \U$46466 ( \46843 , \46840 , \46842 );
not \U$46467 ( \46844 , \46843 );
not \U$46468 ( \46845 , \46206 );
and \U$46469 ( \46846 , \46844 , \46845 );
and \U$46470 ( \46847 , \46843 , \46206 );
nor \U$46471 ( \46848 , \46846 , \46847 );
nor \U$46472 ( \46849 , \46839 , \46848 );
xor \U$46473 ( \46850 , \46338 , \46343 );
xor \U$46474 ( \46851 , \46850 , \46351 );
xor \U$46475 ( \46852 , \46849 , \46851 );
not \U$46476 ( \46853 , \46014 );
not \U$46477 ( \46854 , \46025 );
or \U$46478 ( \46855 , \46853 , \46854 );
or \U$46479 ( \46856 , \46014 , \46025 );
nand \U$46480 ( \46857 , \46855 , \46856 );
not \U$46481 ( \46858 , \46857 );
not \U$46482 ( \46859 , \46007 );
and \U$46483 ( \46860 , \46858 , \46859 );
and \U$46484 ( \46861 , \46857 , \46007 );
nor \U$46485 ( \46862 , \46860 , \46861 );
xor \U$46486 ( \46863 , \46150 , \46157 );
xor \U$46487 ( \46864 , \46863 , \46165 );
xor \U$46488 ( \46865 , \46862 , \46864 );
not \U$46489 ( \46866 , \45987 );
not \U$46490 ( \46867 , \45998 );
or \U$46491 ( \46868 , \46866 , \46867 );
or \U$46492 ( \46869 , \45987 , \45998 );
nand \U$46493 ( \46870 , \46868 , \46869 );
not \U$46494 ( \46871 , \46870 );
not \U$46495 ( \46872 , \45980 );
and \U$46496 ( \46873 , \46871 , \46872 );
and \U$46497 ( \46874 , \46870 , \45980 );
nor \U$46498 ( \46875 , \46873 , \46874 );
and \U$46499 ( \46876 , \46865 , \46875 );
and \U$46500 ( \46877 , \46862 , \46864 );
nor \U$46501 ( \46878 , \46876 , \46877 );
and \U$46502 ( \46879 , \46852 , \46878 );
and \U$46503 ( \46880 , \46849 , \46851 );
or \U$46504 ( \46881 , \46879 , \46880 );
xor \U$46505 ( \46882 , \46832 , \46881 );
xor \U$46506 ( \46883 , \45868 , \45870 );
xor \U$46507 ( \46884 , \46883 , \45879 );
xor \U$46508 ( \46885 , \45892 , \45900 );
xor \U$46509 ( \46886 , \46885 , \45908 );
and \U$46510 ( \46887 , \46884 , \46886 );
xor \U$46511 ( \46888 , \46120 , \46128 );
xor \U$46512 ( \46889 , \46888 , \46136 );
xor \U$46513 ( \46890 , \45892 , \45900 );
xor \U$46514 ( \46891 , \46890 , \45908 );
and \U$46515 ( \46892 , \46889 , \46891 );
and \U$46516 ( \46893 , \46884 , \46889 );
or \U$46517 ( \46894 , \46887 , \46892 , \46893 );
and \U$46518 ( \46895 , \436 , RIae77450_76);
and \U$46519 ( \46896 , RIae77ae0_90, \434 );
nor \U$46520 ( \46897 , \46895 , \46896 );
not \U$46521 ( \46898 , \46897 );
not \U$46522 ( \46899 , \400 );
and \U$46523 ( \46900 , \46898 , \46899 );
and \U$46524 ( \46901 , \46897 , \400 );
nor \U$46525 ( \46902 , \46900 , \46901 );
and \U$46526 ( \46903 , \514 , RIae779f0_88);
and \U$46527 ( \46904 , RIae77810_84, \512 );
nor \U$46528 ( \46905 , \46903 , \46904 );
not \U$46529 ( \46906 , \46905 );
not \U$46530 ( \46907 , \469 );
and \U$46531 ( \46908 , \46906 , \46907 );
and \U$46532 ( \46909 , \46905 , \469 );
nor \U$46533 ( \46910 , \46908 , \46909 );
xor \U$46534 ( \46911 , \46902 , \46910 );
and \U$46535 ( \46912 , \384 , RIae77540_78);
and \U$46536 ( \46913 , RIae776a8_81, \382 );
nor \U$46537 ( \46914 , \46912 , \46913 );
not \U$46538 ( \46915 , \46914 );
not \U$46539 ( \46916 , \392 );
and \U$46540 ( \46917 , \46915 , \46916 );
and \U$46541 ( \46918 , \46914 , \388 );
nor \U$46542 ( \46919 , \46917 , \46918 );
and \U$46543 ( \46920 , \46911 , \46919 );
and \U$46544 ( \46921 , \46902 , \46910 );
nor \U$46545 ( \46922 , \46920 , \46921 );
and \U$46546 ( \46923 , \558 , RIae77900_86);
and \U$46547 ( \46924 , RIae76fa0_66, \556 );
nor \U$46548 ( \46925 , \46923 , \46924 );
and \U$46549 ( \46926 , \46925 , \562 );
not \U$46550 ( \46927 , \46925 );
and \U$46551 ( \46928 , \46927 , \504 );
nor \U$46552 ( \46929 , \46926 , \46928 );
and \U$46553 ( \46930 , \672 , RIae76eb0_64);
and \U$46554 ( \46931 , RIae76dc0_62, \670 );
nor \U$46555 ( \46932 , \46930 , \46931 );
and \U$46556 ( \46933 , \46932 , \587 );
not \U$46557 ( \46934 , \46932 );
and \U$46558 ( \46935 , \46934 , \588 );
nor \U$46559 ( \46936 , \46933 , \46935 );
or \U$46560 ( \46937 , \46929 , \46936 );
not \U$46561 ( \46938 , \46936 );
not \U$46562 ( \46939 , \46929 );
or \U$46563 ( \46940 , \46938 , \46939 );
not \U$46564 ( \46941 , \787 );
and \U$46565 ( \46942 , \883 , RIae76cd0_60);
and \U$46566 ( \46943 , RIae77108_69, \881 );
nor \U$46567 ( \46944 , \46942 , \46943 );
not \U$46568 ( \46945 , \46944 );
or \U$46569 ( \46946 , \46941 , \46945 );
or \U$46570 ( \46947 , \46944 , \789 );
nand \U$46571 ( \46948 , \46946 , \46947 );
nand \U$46572 ( \46949 , \46940 , \46948 );
nand \U$46573 ( \46950 , \46937 , \46949 );
nor \U$46574 ( \46951 , \46922 , \46950 );
not \U$46575 ( \46952 , \46951 );
xor \U$46576 ( \46953 , \46894 , \46952 );
xor \U$46577 ( \46954 , \46094 , \46101 );
xor \U$46578 ( \46955 , \46954 , \46109 );
not \U$46579 ( \46956 , \46073 );
not \U$46580 ( \46957 , \46085 );
or \U$46581 ( \46958 , \46956 , \46957 );
or \U$46582 ( \46959 , \46073 , \46085 );
nand \U$46583 ( \46960 , \46958 , \46959 );
not \U$46584 ( \46961 , \46960 );
not \U$46585 ( \46962 , \46065 );
and \U$46586 ( \46963 , \46961 , \46962 );
and \U$46587 ( \46964 , \46960 , \46065 );
nor \U$46588 ( \46965 , \46963 , \46964 );
xor \U$46589 ( \46966 , \46955 , \46965 );
not \U$46590 ( \46967 , \46042 );
not \U$46591 ( \46968 , \46053 );
or \U$46592 ( \46969 , \46967 , \46968 );
or \U$46593 ( \46970 , \46042 , \46053 );
nand \U$46594 ( \46971 , \46969 , \46970 );
not \U$46595 ( \46972 , \46971 );
not \U$46596 ( \46973 , \46035 );
and \U$46597 ( \46974 , \46972 , \46973 );
and \U$46598 ( \46975 , \46971 , \46035 );
nor \U$46599 ( \46976 , \46974 , \46975 );
and \U$46600 ( \46977 , \46966 , \46976 );
and \U$46601 ( \46978 , \46955 , \46965 );
nor \U$46602 ( \46979 , \46977 , \46978 );
and \U$46603 ( \46980 , \46953 , \46979 );
and \U$46604 ( \46981 , \46894 , \46952 );
or \U$46605 ( \46982 , \46980 , \46981 );
and \U$46606 ( \46983 , \46882 , \46982 );
and \U$46607 ( \46984 , \46832 , \46881 );
or \U$46608 ( \46985 , \46983 , \46984 );
xor \U$46609 ( \46986 , \46599 , \46985 );
xor \U$46610 ( \46987 , \45860 , \45914 );
xor \U$46611 ( \46988 , \46987 , \45970 );
xor \U$46612 ( \46989 , \46300 , \46301 );
xor \U$46613 ( \46990 , \46989 , \46306 );
and \U$46614 ( \46991 , \46988 , \46990 );
xor \U$46615 ( \46992 , \45737 , \45739 );
xor \U$46616 ( \46993 , \46992 , \45742 );
xor \U$46617 ( \46994 , \46315 , \46322 );
xor \U$46618 ( \46995 , \46993 , \46994 );
xor \U$46619 ( \46996 , \46300 , \46301 );
xor \U$46620 ( \46997 , \46996 , \46306 );
and \U$46621 ( \46998 , \46995 , \46997 );
and \U$46622 ( \46999 , \46988 , \46995 );
or \U$46623 ( \47000 , \46991 , \46998 , \46999 );
and \U$46624 ( \47001 , \46986 , \47000 );
and \U$46625 ( \47002 , \46599 , \46985 );
or \U$46626 ( \47003 , \47001 , \47002 );
xor \U$46627 ( \47004 , \46479 , \46495 );
xor \U$46628 ( \47005 , \47004 , \46500 );
xor \U$46629 ( \47006 , \47003 , \47005 );
xor \U$46630 ( \47007 , \46483 , \46487 );
xor \U$46631 ( \47008 , \47007 , \46492 );
xor \U$46632 ( \47009 , \46327 , \46394 );
xor \U$46633 ( \47010 , \47009 , \46403 );
and \U$46634 ( \47011 , \47008 , \47010 );
xor \U$46635 ( \47012 , \45758 , \45763 );
xor \U$46636 ( \47013 , \47012 , \45768 );
xor \U$46637 ( \47014 , \45746 , \45780 );
xor \U$46638 ( \47015 , \47013 , \47014 );
xor \U$46639 ( \47016 , \46327 , \46394 );
xor \U$46640 ( \47017 , \47016 , \46403 );
and \U$46641 ( \47018 , \47015 , \47017 );
and \U$46642 ( \47019 , \47008 , \47015 );
or \U$46643 ( \47020 , \47011 , \47018 , \47019 );
and \U$46644 ( \47021 , \47006 , \47020 );
and \U$46645 ( \47022 , \47003 , \47005 );
or \U$46646 ( \47023 , \47021 , \47022 );
xor \U$46647 ( \47024 , \46468 , \46470 );
xor \U$46648 ( \47025 , \47024 , \46513 );
and \U$46649 ( \47026 , \47023 , \47025 );
xor \U$46650 ( \47027 , \46409 , \46411 );
xor \U$46651 ( \47028 , \47027 , \46452 );
xor \U$46652 ( \47029 , \46468 , \46470 );
xor \U$46653 ( \47030 , \47029 , \46513 );
and \U$46654 ( \47031 , \47028 , \47030 );
and \U$46655 ( \47032 , \47023 , \47028 );
or \U$46656 ( \47033 , \47026 , \47031 , \47032 );
xor \U$46657 ( \47034 , \46525 , \46533 );
xor \U$46658 ( \47035 , \47034 , \46538 );
xor \U$46659 ( \47036 , \47033 , \47035 );
xor \U$46660 ( \47037 , \46455 , \46457 );
xor \U$46661 ( \47038 , \47037 , \46516 );
and \U$46662 ( \47039 , \47036 , \47038 );
and \U$46663 ( \47040 , \47033 , \47035 );
or \U$46664 ( \47041 , \47039 , \47040 );
xor \U$46665 ( \47042 , \46519 , \46547 );
and \U$46666 ( \47043 , \47041 , \47042 );
xor \U$46667 ( \47044 , \47042 , \47041 );
xor \U$46668 ( \47045 , \45785 , \46312 );
xor \U$46669 ( \47046 , \47045 , \46406 );
xor \U$46670 ( \47047 , \47003 , \47005 );
xor \U$46671 ( \47048 , \47047 , \47020 );
and \U$46672 ( \47049 , \47046 , \47048 );
xor \U$46673 ( \47050 , \46599 , \46985 );
xor \U$46674 ( \47051 , \47050 , \47000 );
xor \U$46675 ( \47052 , \46327 , \46394 );
xor \U$46676 ( \47053 , \47052 , \46403 );
xor \U$46677 ( \47054 , \47008 , \47015 );
xor \U$46678 ( \47055 , \47053 , \47054 );
and \U$46679 ( \47056 , \47051 , \47055 );
xor \U$46680 ( \47057 , \46422 , \46430 );
xor \U$46681 ( \47058 , \47057 , \46435 );
xor \U$46682 ( \47059 , \46414 , \46447 );
xor \U$46683 ( \47060 , \47058 , \47059 );
xor \U$46684 ( \47061 , \47056 , \47060 );
xor \U$46685 ( \47062 , \46775 , \46800 );
xor \U$46686 ( \47063 , \47062 , \46826 );
not \U$46687 ( \47064 , \46747 );
not \U$46688 ( \47065 , \46705 );
or \U$46689 ( \47066 , \47064 , \47065 );
or \U$46690 ( \47067 , \46705 , \46747 );
nand \U$46691 ( \47068 , \47066 , \47067 );
not \U$46692 ( \47069 , \47068 );
not \U$46693 ( \47070 , \46716 );
and \U$46694 ( \47071 , \47069 , \47070 );
and \U$46695 ( \47072 , \47068 , \46716 );
nor \U$46696 ( \47073 , \47071 , \47072 );
xor \U$46697 ( \47074 , \47063 , \47073 );
xor \U$46698 ( \47075 , \46624 , \46649 );
xor \U$46699 ( \47076 , \47075 , \46677 );
and \U$46700 ( \47077 , \47074 , \47076 );
and \U$46701 ( \47078 , \47063 , \47073 );
or \U$46702 ( \47079 , \47077 , \47078 );
not \U$46703 ( \47080 , \46219 );
not \U$46704 ( \47081 , \46195 );
or \U$46705 ( \47082 , \47080 , \47081 );
or \U$46706 ( \47083 , \46195 , \46219 );
nand \U$46707 ( \47084 , \47082 , \47083 );
not \U$46708 ( \47085 , \47084 );
not \U$46709 ( \47086 , \46168 );
and \U$46710 ( \47087 , \47085 , \47086 );
and \U$46711 ( \47088 , \47084 , \46168 );
nor \U$46712 ( \47089 , \47087 , \47088 );
or \U$46713 ( \47090 , \47079 , \47089 );
not \U$46714 ( \47091 , \47089 );
not \U$46715 ( \47092 , \47079 );
or \U$46716 ( \47093 , \47091 , \47092 );
xor \U$46717 ( \47094 , \46955 , \46965 );
xor \U$46718 ( \47095 , \47094 , \46976 );
and \U$46719 ( \47096 , \46922 , \46950 );
nor \U$46720 ( \47097 , \47096 , \46951 );
or \U$46721 ( \47098 , \47095 , \47097 );
not \U$46722 ( \47099 , \47097 );
not \U$46723 ( \47100 , \47095 );
or \U$46724 ( \47101 , \47099 , \47100 );
xor \U$46725 ( \47102 , \45892 , \45900 );
xor \U$46726 ( \47103 , \47102 , \45908 );
xor \U$46727 ( \47104 , \46884 , \46889 );
xor \U$46728 ( \47105 , \47103 , \47104 );
nand \U$46729 ( \47106 , \47101 , \47105 );
nand \U$46730 ( \47107 , \47098 , \47106 );
nand \U$46731 ( \47108 , \47093 , \47107 );
nand \U$46732 ( \47109 , \47090 , \47108 );
and \U$46733 ( \47110 , \2607 , RIae78440_110);
and \U$46734 ( \47111 , RIae784b8_111, \2605 );
nor \U$46735 ( \47112 , \47110 , \47111 );
and \U$46736 ( \47113 , \47112 , \2397 );
not \U$46737 ( \47114 , \47112 );
and \U$46738 ( \47115 , \47114 , \2611 );
nor \U$46739 ( \47116 , \47113 , \47115 );
not \U$46740 ( \47117 , \47116 );
and \U$46741 ( \47118 , \2783 , RIae77cc0_94);
and \U$46742 ( \47119 , RIae77bd0_92, \2781 );
nor \U$46743 ( \47120 , \47118 , \47119 );
not \U$46744 ( \47121 , \47120 );
not \U$46745 ( \47122 , \3089 );
and \U$46746 ( \47123 , \47121 , \47122 );
and \U$46747 ( \47124 , \47120 , \2789 );
nor \U$46748 ( \47125 , \47123 , \47124 );
not \U$46749 ( \47126 , \47125 );
and \U$46750 ( \47127 , \47117 , \47126 );
and \U$46751 ( \47128 , \47125 , \47116 );
and \U$46752 ( \47129 , \3214 , RIae77db0_96);
and \U$46753 ( \47130 , RIae77ea0_98, \3212 );
nor \U$46754 ( \47131 , \47129 , \47130 );
not \U$46755 ( \47132 , \47131 );
not \U$46756 ( \47133 , \2774 );
and \U$46757 ( \47134 , \47132 , \47133 );
and \U$46758 ( \47135 , \47131 , \2774 );
nor \U$46759 ( \47136 , \47134 , \47135 );
nor \U$46760 ( \47137 , \47128 , \47136 );
nor \U$46761 ( \47138 , \47127 , \47137 );
and \U$46762 ( \47139 , \1593 , RIae78350_108);
and \U$46763 ( \47140 , RIae78170_104, \1591 );
nor \U$46764 ( \47141 , \47139 , \47140 );
and \U$46765 ( \47142 , \47141 , \1488 );
not \U$46766 ( \47143 , \47141 );
and \U$46767 ( \47144 , \47143 , \1498 );
nor \U$46768 ( \47145 , \47142 , \47144 );
not \U$46769 ( \47146 , \47145 );
and \U$46770 ( \47147 , \2224 , RIae78260_106);
and \U$46771 ( \47148 , RIae78620_114, \2222 );
nor \U$46772 ( \47149 , \47147 , \47148 );
and \U$46773 ( \47150 , \47149 , \2060 );
not \U$46774 ( \47151 , \47149 );
and \U$46775 ( \47152 , \47151 , \2061 );
nor \U$46776 ( \47153 , \47150 , \47152 );
not \U$46777 ( \47154 , \47153 );
and \U$46778 ( \47155 , \47146 , \47154 );
and \U$46779 ( \47156 , \47153 , \47145 );
and \U$46780 ( \47157 , \1939 , RIae77f90_100);
and \U$46781 ( \47158 , RIae78080_102, \1937 );
nor \U$46782 ( \47159 , \47157 , \47158 );
and \U$46783 ( \47160 , \47159 , \1734 );
not \U$46784 ( \47161 , \47159 );
and \U$46785 ( \47162 , \47161 , \1735 );
nor \U$46786 ( \47163 , \47160 , \47162 );
nor \U$46787 ( \47164 , \47156 , \47163 );
nor \U$46788 ( \47165 , \47155 , \47164 );
xor \U$46789 ( \47166 , \47138 , \47165 );
and \U$46790 ( \47167 , \883 , RIae76dc0_62);
and \U$46791 ( \47168 , RIae76cd0_60, \881 );
nor \U$46792 ( \47169 , \47167 , \47168 );
not \U$46793 ( \47170 , \47169 );
not \U$46794 ( \47171 , \787 );
and \U$46795 ( \47172 , \47170 , \47171 );
and \U$46796 ( \47173 , \47169 , \787 );
nor \U$46797 ( \47174 , \47172 , \47173 );
not \U$46798 ( \47175 , \47174 );
and \U$46799 ( \47176 , \1138 , RIae77108_69);
and \U$46800 ( \47177 , RIae77090_68, \1136 );
nor \U$46801 ( \47178 , \47176 , \47177 );
and \U$46802 ( \47179 , \47178 , \1142 );
not \U$46803 ( \47180 , \47178 );
and \U$46804 ( \47181 , \47180 , \1012 );
nor \U$46805 ( \47182 , \47179 , \47181 );
not \U$46806 ( \47183 , \47182 );
and \U$46807 ( \47184 , \47175 , \47183 );
and \U$46808 ( \47185 , \47182 , \47174 );
and \U$46809 ( \47186 , \1376 , RIae77270_72);
and \U$46810 ( \47187 , RIae77360_74, \1374 );
nor \U$46811 ( \47188 , \47186 , \47187 );
and \U$46812 ( \47189 , \47188 , \1261 );
not \U$46813 ( \47190 , \47188 );
and \U$46814 ( \47191 , \47190 , \1380 );
nor \U$46815 ( \47192 , \47189 , \47191 );
nor \U$46816 ( \47193 , \47185 , \47192 );
nor \U$46817 ( \47194 , \47184 , \47193 );
and \U$46818 ( \47195 , \47166 , \47194 );
and \U$46819 ( \47196 , \47138 , \47165 );
or \U$46820 ( \47197 , \47195 , \47196 );
and \U$46821 ( \47198 , \8966 , RIae75380_6);
and \U$46822 ( \47199 , RIae75470_8, \8964 );
nor \U$46823 ( \47200 , \47198 , \47199 );
and \U$46824 ( \47201 , \47200 , \8789 );
not \U$46825 ( \47202 , \47200 );
and \U$46826 ( \47203 , \47202 , \8799 );
nor \U$46827 ( \47204 , \47201 , \47203 );
not \U$46828 ( \47205 , \47204 );
and \U$46829 ( \47206 , \10548 , RIae76730_48);
and \U$46830 ( \47207 , RIae76640_46, \10546 );
nor \U$46831 ( \47208 , \47206 , \47207 );
and \U$46832 ( \47209 , \47208 , \10118 );
not \U$46833 ( \47210 , \47208 );
and \U$46834 ( \47211 , \47210 , \10421 );
nor \U$46835 ( \47212 , \47209 , \47211 );
not \U$46836 ( \47213 , \47212 );
and \U$46837 ( \47214 , \47205 , \47213 );
and \U$46838 ( \47215 , \47212 , \47204 );
and \U$46839 ( \47216 , \9760 , RIae76460_42);
and \U$46840 ( \47217 , RIae76550_44, \9758 );
nor \U$46841 ( \47218 , \47216 , \47217 );
and \U$46842 ( \47219 , \47218 , \9272 );
not \U$46843 ( \47220 , \47218 );
and \U$46844 ( \47221 , \47220 , \9273 );
nor \U$46845 ( \47222 , \47219 , \47221 );
nor \U$46846 ( \47223 , \47215 , \47222 );
nor \U$46847 ( \47224 , \47214 , \47223 );
and \U$46848 ( \47225 , \14964 , RIae76be0_58);
and \U$46849 ( \47226 , RIae78ad0_124, \14962 );
nor \U$46850 ( \47227 , \47225 , \47226 );
and \U$46851 ( \47228 , \47227 , \14462 );
not \U$46852 ( \47229 , \47227 );
and \U$46853 ( \47230 , \47229 , \14463 );
nor \U$46854 ( \47231 , \47228 , \47230 );
and \U$46855 ( \47232 , \15726 , RIae78d28_129);
and \U$46856 ( \47233 , RIae78e18_131, RIae7aab0_192);
nor \U$46857 ( \47234 , \47232 , \47233 );
and \U$46858 ( \47235 , \47234 , RIae7aa38_191);
not \U$46859 ( \47236 , \47234 );
and \U$46860 ( \47237 , \47236 , \14959 );
nor \U$46861 ( \47238 , \47235 , \47237 );
xor \U$46862 ( \47239 , \47231 , \47238 );
and \U$46863 ( \47240 , \14059 , RIae76820_50);
and \U$46864 ( \47241 , RIae76910_52, \14057 );
nor \U$46865 ( \47242 , \47240 , \47241 );
and \U$46866 ( \47243 , \47242 , \14063 );
not \U$46867 ( \47244 , \47242 );
and \U$46868 ( \47245 , \47244 , \13502 );
nor \U$46869 ( \47246 , \47243 , \47245 );
and \U$46870 ( \47247 , \47239 , \47246 );
and \U$46871 ( \47248 , \47231 , \47238 );
or \U$46872 ( \47249 , \47247 , \47248 );
xor \U$46873 ( \47250 , \47224 , \47249 );
and \U$46874 ( \47251 , \11470 , RIae76190_36);
and \U$46875 ( \47252 , RIae760a0_34, \11468 );
nor \U$46876 ( \47253 , \47251 , \47252 );
and \U$46877 ( \47254 , \47253 , \11474 );
not \U$46878 ( \47255 , \47253 );
and \U$46879 ( \47256 , \47255 , \10936 );
nor \U$46880 ( \47257 , \47254 , \47256 );
not \U$46881 ( \47258 , \47257 );
and \U$46882 ( \47259 , \12180 , RIae76370_40);
and \U$46883 ( \47260 , RIae76280_38, \12178 );
nor \U$46884 ( \47261 , \47259 , \47260 );
and \U$46885 ( \47262 , \47261 , \11827 );
not \U$46886 ( \47263 , \47261 );
and \U$46887 ( \47264 , \47263 , \12184 );
nor \U$46888 ( \47265 , \47262 , \47264 );
not \U$46889 ( \47266 , \47265 );
and \U$46890 ( \47267 , \47258 , \47266 );
and \U$46891 ( \47268 , \47265 , \47257 );
and \U$46892 ( \47269 , \13059 , RIae76af0_56);
and \U$46893 ( \47270 , RIae76a00_54, \13057 );
nor \U$46894 ( \47271 , \47269 , \47270 );
and \U$46895 ( \47272 , \47271 , \12718 );
not \U$46896 ( \47273 , \47271 );
and \U$46897 ( \47274 , \47273 , \13063 );
nor \U$46898 ( \47275 , \47272 , \47274 );
nor \U$46899 ( \47276 , \47268 , \47275 );
nor \U$46900 ( \47277 , \47267 , \47276 );
and \U$46901 ( \47278 , \47250 , \47277 );
and \U$46902 ( \47279 , \47224 , \47249 );
or \U$46903 ( \47280 , \47278 , \47279 );
xor \U$46904 ( \47281 , \47197 , \47280 );
and \U$46905 ( \47282 , \5399 , RIae75a10_20);
and \U$46906 ( \47283 , RIae75920_18, \5397 );
nor \U$46907 ( \47284 , \47282 , \47283 );
and \U$46908 ( \47285 , \47284 , \5403 );
not \U$46909 ( \47286 , \47284 );
and \U$46910 ( \47287 , \47286 , \5016 );
nor \U$46911 ( \47288 , \47285 , \47287 );
not \U$46912 ( \47289 , \47288 );
and \U$46913 ( \47290 , \5896 , RIae75fb0_32);
and \U$46914 ( \47291 , RIae75ec0_30, \5894 );
nor \U$46915 ( \47292 , \47290 , \47291 );
and \U$46916 ( \47293 , \47292 , \5589 );
not \U$46917 ( \47294 , \47292 );
and \U$46918 ( \47295 , \47294 , \5590 );
nor \U$46919 ( \47296 , \47293 , \47295 );
not \U$46920 ( \47297 , \47296 );
and \U$46921 ( \47298 , \47289 , \47297 );
and \U$46922 ( \47299 , \47296 , \47288 );
and \U$46923 ( \47300 , \6172 , RIae75ce0_26);
and \U$46924 ( \47301 , RIae75dd0_28, \6170 );
nor \U$46925 ( \47302 , \47300 , \47301 );
and \U$46926 ( \47303 , \47302 , \6175 );
not \U$46927 ( \47304 , \47302 );
and \U$46928 ( \47305 , \47304 , \6176 );
nor \U$46929 ( \47306 , \47303 , \47305 );
nor \U$46930 ( \47307 , \47299 , \47306 );
nor \U$46931 ( \47308 , \47298 , \47307 );
and \U$46932 ( \47309 , \4247 , RIae78800_118);
and \U$46933 ( \47310 , RIae78710_116, \4245 );
nor \U$46934 ( \47311 , \47309 , \47310 );
and \U$46935 ( \47312 , \47311 , \3989 );
not \U$46936 ( \47313 , \47311 );
and \U$46937 ( \47314 , \47313 , \4251 );
nor \U$46938 ( \47315 , \47312 , \47314 );
and \U$46939 ( \47316 , \4688 , RIae75bf0_24);
and \U$46940 ( \47317 , RIae75b00_22, \4686 );
nor \U$46941 ( \47318 , \47316 , \47317 );
and \U$46942 ( \47319 , \47318 , \4481 );
not \U$46943 ( \47320 , \47318 );
and \U$46944 ( \47321 , \47320 , \4482 );
nor \U$46945 ( \47322 , \47319 , \47321 );
xor \U$46946 ( \47323 , \47315 , \47322 );
and \U$46947 ( \47324 , \3730 , RIae789e0_122);
and \U$46948 ( \47325 , RIae788f0_120, \3728 );
nor \U$46949 ( \47326 , \47324 , \47325 );
and \U$46950 ( \47327 , \47326 , \3732 );
not \U$46951 ( \47328 , \47326 );
and \U$46952 ( \47329 , \47328 , \3422 );
nor \U$46953 ( \47330 , \47327 , \47329 );
and \U$46954 ( \47331 , \47323 , \47330 );
and \U$46955 ( \47332 , \47315 , \47322 );
nor \U$46956 ( \47333 , \47331 , \47332 );
xor \U$46957 ( \47334 , \47308 , \47333 );
and \U$46958 ( \47335 , \6941 , RIae75650_12);
and \U$46959 ( \47336 , RIae75560_10, \6939 );
nor \U$46960 ( \47337 , \47335 , \47336 );
and \U$46961 ( \47338 , \47337 , \6945 );
not \U$46962 ( \47339 , \47337 );
and \U$46963 ( \47340 , \47339 , \6314 );
nor \U$46964 ( \47341 , \47338 , \47340 );
not \U$46965 ( \47342 , \47341 );
and \U$46966 ( \47343 , \7633 , RIae75830_16);
and \U$46967 ( \47344 , RIae75740_14, \7631 );
nor \U$46968 ( \47345 , \47343 , \47344 );
and \U$46969 ( \47346 , \47345 , \7205 );
not \U$46970 ( \47347 , \47345 );
and \U$46971 ( \47348 , \47347 , \7206 );
nor \U$46972 ( \47349 , \47346 , \47348 );
not \U$46973 ( \47350 , \47349 );
and \U$46974 ( \47351 , \47342 , \47350 );
and \U$46975 ( \47352 , \47349 , \47341 );
and \U$46976 ( \47353 , \8371 , RIae75290_4);
and \U$46977 ( \47354 , RIae751a0_2, \8369 );
nor \U$46978 ( \47355 , \47353 , \47354 );
and \U$46979 ( \47356 , \47355 , \8019 );
not \U$46980 ( \47357 , \47355 );
and \U$46981 ( \47358 , \47357 , \8020 );
nor \U$46982 ( \47359 , \47356 , \47358 );
nor \U$46983 ( \47360 , \47352 , \47359 );
nor \U$46984 ( \47361 , \47351 , \47360 );
and \U$46985 ( \47362 , \47334 , \47361 );
and \U$46986 ( \47363 , \47308 , \47333 );
or \U$46987 ( \47364 , \47362 , \47363 );
and \U$46988 ( \47365 , \47281 , \47364 );
and \U$46989 ( \47366 , \47197 , \47280 );
or \U$46990 ( \47367 , \47365 , \47366 );
not \U$46991 ( \47368 , \46936 );
not \U$46992 ( \47369 , \46948 );
or \U$46993 ( \47370 , \47368 , \47369 );
or \U$46994 ( \47371 , \46936 , \46948 );
nand \U$46995 ( \47372 , \47370 , \47371 );
not \U$46996 ( \47373 , \47372 );
not \U$46997 ( \47374 , \46929 );
and \U$46998 ( \47375 , \47373 , \47374 );
and \U$46999 ( \47376 , \47372 , \46929 );
nor \U$47000 ( \47377 , \47375 , \47376 );
xor \U$47001 ( \47378 , \46606 , \46613 );
xor \U$47002 ( \47379 , \47378 , \46621 );
xor \U$47003 ( \47380 , \47377 , \47379 );
xor \U$47004 ( \47381 , \46631 , \46638 );
xor \U$47005 ( \47382 , \47381 , \46646 );
and \U$47006 ( \47383 , \47380 , \47382 );
and \U$47007 ( \47384 , \47377 , \47379 );
or \U$47008 ( \47385 , \47383 , \47384 );
and \U$47009 ( \47386 , \514 , RIae77ae0_90);
and \U$47010 ( \47387 , RIae779f0_88, \512 );
nor \U$47011 ( \47388 , \47386 , \47387 );
not \U$47012 ( \47389 , \47388 );
not \U$47013 ( \47390 , \471 );
and \U$47014 ( \47391 , \47389 , \47390 );
and \U$47015 ( \47392 , \47388 , \469 );
nor \U$47016 ( \47393 , \47391 , \47392 );
not \U$47017 ( \47394 , \47393 );
and \U$47018 ( \47395 , \672 , RIae76fa0_66);
and \U$47019 ( \47396 , RIae76eb0_64, \670 );
nor \U$47020 ( \47397 , \47395 , \47396 );
and \U$47021 ( \47398 , \47397 , \587 );
not \U$47022 ( \47399 , \47397 );
and \U$47023 ( \47400 , \47399 , \588 );
nor \U$47024 ( \47401 , \47398 , \47400 );
not \U$47025 ( \47402 , \47401 );
and \U$47026 ( \47403 , \47394 , \47402 );
and \U$47027 ( \47404 , \47401 , \47393 );
and \U$47028 ( \47405 , \558 , RIae77810_84);
and \U$47029 ( \47406 , RIae77900_86, \556 );
nor \U$47030 ( \47407 , \47405 , \47406 );
and \U$47031 ( \47408 , \47407 , \562 );
not \U$47032 ( \47409 , \47407 );
and \U$47033 ( \47410 , \47409 , \504 );
nor \U$47034 ( \47411 , \47408 , \47410 );
nor \U$47035 ( \47412 , \47404 , \47411 );
nor \U$47036 ( \47413 , \47403 , \47412 );
nand \U$47037 ( \47414 , RIae77630_80, RIae78b48_125);
xor \U$47038 ( \47415 , \47413 , \47414 );
xor \U$47039 ( \47416 , \46902 , \46910 );
xor \U$47040 ( \47417 , \47416 , \46919 );
and \U$47041 ( \47418 , \47415 , \47417 );
and \U$47042 ( \47419 , \47413 , \47414 );
or \U$47043 ( \47420 , \47418 , \47419 );
xor \U$47044 ( \47421 , \47385 , \47420 );
xor \U$47045 ( \47422 , \46757 , \46764 );
xor \U$47046 ( \47423 , \47422 , \46772 );
xor \U$47047 ( \47424 , \46658 , \46666 );
xor \U$47048 ( \47425 , \47424 , \46674 );
and \U$47049 ( \47426 , \47423 , \47425 );
xor \U$47050 ( \47427 , \46782 , \46789 );
xor \U$47051 ( \47428 , \47427 , \46797 );
xor \U$47052 ( \47429 , \46658 , \46666 );
xor \U$47053 ( \47430 , \47429 , \46674 );
and \U$47054 ( \47431 , \47428 , \47430 );
and \U$47055 ( \47432 , \47423 , \47428 );
or \U$47056 ( \47433 , \47426 , \47431 , \47432 );
and \U$47057 ( \47434 , \47421 , \47433 );
and \U$47058 ( \47435 , \47385 , \47420 );
or \U$47059 ( \47436 , \47434 , \47435 );
xor \U$47060 ( \47437 , \47367 , \47436 );
xor \U$47061 ( \47438 , \46808 , \46815 );
xor \U$47062 ( \47439 , \47438 , \46823 );
not \U$47063 ( \47440 , \46734 );
not \U$47064 ( \47441 , \46745 );
or \U$47065 ( \47442 , \47440 , \47441 );
or \U$47066 ( \47443 , \46734 , \46745 );
nand \U$47067 ( \47444 , \47442 , \47443 );
not \U$47068 ( \47445 , \47444 );
not \U$47069 ( \47446 , \46727 );
and \U$47070 ( \47447 , \47445 , \47446 );
and \U$47071 ( \47448 , \47444 , \46727 );
nor \U$47072 ( \47449 , \47447 , \47448 );
xor \U$47073 ( \47450 , \47439 , \47449 );
xor \U$47074 ( \47451 , \46687 , \46694 );
xor \U$47075 ( \47452 , \47451 , \46702 );
and \U$47076 ( \47453 , \47450 , \47452 );
and \U$47077 ( \47454 , \47439 , \47449 );
or \U$47078 ( \47455 , \47453 , \47454 );
not \U$47079 ( \47456 , \46848 );
not \U$47080 ( \47457 , \46838 );
and \U$47081 ( \47458 , \47456 , \47457 );
and \U$47082 ( \47459 , \46848 , \46838 );
nor \U$47083 ( \47460 , \47458 , \47459 );
xor \U$47084 ( \47461 , \47455 , \47460 );
xor \U$47085 ( \47462 , \46862 , \46864 );
xor \U$47086 ( \47463 , \47462 , \46875 );
and \U$47087 ( \47464 , \47461 , \47463 );
and \U$47088 ( \47465 , \47455 , \47460 );
or \U$47089 ( \47466 , \47464 , \47465 );
and \U$47090 ( \47467 , \47437 , \47466 );
and \U$47091 ( \47468 , \47367 , \47436 );
nor \U$47092 ( \47469 , \47467 , \47468 );
xor \U$47093 ( \47470 , \47109 , \47469 );
xor \U$47094 ( \47471 , \46849 , \46851 );
xor \U$47095 ( \47472 , \47471 , \46878 );
xor \U$47096 ( \47473 , \46583 , \46585 );
xor \U$47097 ( \47474 , \47473 , \46588 );
and \U$47098 ( \47475 , \47472 , \47474 );
xor \U$47099 ( \47476 , \45809 , \45833 );
xor \U$47100 ( \47477 , \47476 , \45857 );
xor \U$47101 ( \47478 , \46569 , \46576 );
xor \U$47102 ( \47479 , \47477 , \47478 );
xor \U$47103 ( \47480 , \46583 , \46585 );
xor \U$47104 ( \47481 , \47480 , \46588 );
and \U$47105 ( \47482 , \47479 , \47481 );
and \U$47106 ( \47483 , \47472 , \47479 );
or \U$47107 ( \47484 , \47475 , \47482 , \47483 );
and \U$47108 ( \47485 , \47470 , \47484 );
and \U$47109 ( \47486 , \47109 , \47469 );
or \U$47110 ( \47487 , \47485 , \47486 );
xor \U$47111 ( \47488 , \45973 , \46224 );
xor \U$47112 ( \47489 , \47488 , \46309 );
xor \U$47113 ( \47490 , \47487 , \47489 );
xor \U$47114 ( \47491 , \46058 , \46142 );
xor \U$47115 ( \47492 , \47491 , \46221 );
xor \U$47116 ( \47493 , \46581 , \46591 );
xor \U$47117 ( \47494 , \47493 , \46596 );
and \U$47118 ( \47495 , \47492 , \47494 );
xor \U$47119 ( \47496 , \46300 , \46301 );
xor \U$47120 ( \47497 , \47496 , \46306 );
xor \U$47121 ( \47498 , \46988 , \46995 );
xor \U$47122 ( \47499 , \47497 , \47498 );
xor \U$47123 ( \47500 , \46581 , \46591 );
xor \U$47124 ( \47501 , \47500 , \46596 );
and \U$47125 ( \47502 , \47499 , \47501 );
and \U$47126 ( \47503 , \47492 , \47499 );
or \U$47127 ( \47504 , \47495 , \47502 , \47503 );
and \U$47128 ( \47505 , \47490 , \47504 );
and \U$47129 ( \47506 , \47487 , \47489 );
or \U$47130 ( \47507 , \47505 , \47506 );
and \U$47131 ( \47508 , \47061 , \47507 );
and \U$47132 ( \47509 , \47056 , \47060 );
or \U$47133 ( \47510 , \47508 , \47509 );
xor \U$47134 ( \47511 , \47049 , \47510 );
xor \U$47135 ( \47512 , \46468 , \46470 );
xor \U$47136 ( \47513 , \47512 , \46513 );
xor \U$47137 ( \47514 , \47023 , \47028 );
xor \U$47138 ( \47515 , \47513 , \47514 );
and \U$47139 ( \47516 , \47511 , \47515 );
and \U$47140 ( \47517 , \47049 , \47510 );
or \U$47141 ( \47518 , \47516 , \47517 );
not \U$47142 ( \47519 , \47518 );
xor \U$47143 ( \47520 , \47033 , \47035 );
xor \U$47144 ( \47521 , \47520 , \47038 );
not \U$47145 ( \47522 , \47521 );
or \U$47146 ( \47523 , \47519 , \47522 );
xor \U$47147 ( \47524 , \47049 , \47510 );
xor \U$47148 ( \47525 , \47524 , \47515 );
xor \U$47149 ( \47526 , \47046 , \47048 );
not \U$47150 ( \47527 , \47526 );
xor \U$47151 ( \47528 , \47056 , \47060 );
xor \U$47152 ( \47529 , \47528 , \47507 );
not \U$47153 ( \47530 , \47529 );
or \U$47154 ( \47531 , \47527 , \47530 );
or \U$47155 ( \47532 , \47529 , \47526 );
xor \U$47156 ( \47533 , \47051 , \47055 );
not \U$47157 ( \47534 , \47533 );
xor \U$47158 ( \47535 , \47487 , \47489 );
xor \U$47159 ( \47536 , \47535 , \47504 );
not \U$47160 ( \47537 , \47536 );
or \U$47161 ( \47538 , \47534 , \47537 );
or \U$47162 ( \47539 , \47536 , \47533 );
xor \U$47163 ( \47540 , \46680 , \46749 );
xor \U$47164 ( \47541 , \47540 , \46829 );
xor \U$47165 ( \47542 , \46894 , \46952 );
xor \U$47166 ( \47543 , \47542 , \46979 );
and \U$47167 ( \47544 , \47541 , \47543 );
xor \U$47168 ( \47545 , \46583 , \46585 );
xor \U$47169 ( \47546 , \47545 , \46588 );
xor \U$47170 ( \47547 , \47472 , \47479 );
xor \U$47171 ( \47548 , \47546 , \47547 );
xor \U$47172 ( \47549 , \46894 , \46952 );
xor \U$47173 ( \47550 , \47549 , \46979 );
and \U$47174 ( \47551 , \47548 , \47550 );
and \U$47175 ( \47552 , \47541 , \47548 );
or \U$47176 ( \47553 , \47544 , \47551 , \47552 );
xor \U$47177 ( \47554 , \46832 , \46881 );
xor \U$47178 ( \47555 , \47554 , \46982 );
xor \U$47179 ( \47556 , \47553 , \47555 );
not \U$47180 ( \47557 , \3218 );
and \U$47181 ( \47558 , \3214 , RIae77bd0_92);
and \U$47182 ( \47559 , RIae77db0_96, \3212 );
nor \U$47183 ( \47560 , \47558 , \47559 );
not \U$47184 ( \47561 , \47560 );
or \U$47185 ( \47562 , \47557 , \47561 );
or \U$47186 ( \47563 , \47560 , \2774 );
nand \U$47187 ( \47564 , \47562 , \47563 );
not \U$47188 ( \47565 , \3089 );
and \U$47189 ( \47566 , \2783 , RIae784b8_111);
and \U$47190 ( \47567 , RIae77cc0_94, \2781 );
nor \U$47191 ( \47568 , \47566 , \47567 );
not \U$47192 ( \47569 , \47568 );
or \U$47193 ( \47570 , \47565 , \47569 );
or \U$47194 ( \47571 , \47568 , \2789 );
nand \U$47195 ( \47572 , \47570 , \47571 );
xor \U$47196 ( \47573 , \47564 , \47572 );
and \U$47197 ( \47574 , \3730 , RIae77ea0_98);
and \U$47198 ( \47575 , RIae789e0_122, \3728 );
nor \U$47199 ( \47576 , \47574 , \47575 );
and \U$47200 ( \47577 , \47576 , \3732 );
not \U$47201 ( \47578 , \47576 );
and \U$47202 ( \47579 , \47578 , \3422 );
nor \U$47203 ( \47580 , \47577 , \47579 );
and \U$47204 ( \47581 , \47573 , \47580 );
and \U$47205 ( \47582 , \47564 , \47572 );
or \U$47206 ( \47583 , \47581 , \47582 );
and \U$47207 ( \47584 , \2607 , RIae78620_114);
and \U$47208 ( \47585 , RIae78440_110, \2605 );
nor \U$47209 ( \47586 , \47584 , \47585 );
and \U$47210 ( \47587 , \47586 , \2611 );
not \U$47211 ( \47588 , \47586 );
and \U$47212 ( \47589 , \47588 , \2397 );
nor \U$47213 ( \47590 , \47587 , \47589 );
and \U$47214 ( \47591 , \1939 , RIae78170_104);
and \U$47215 ( \47592 , RIae77f90_100, \1937 );
nor \U$47216 ( \47593 , \47591 , \47592 );
and \U$47217 ( \47594 , \47593 , \1735 );
not \U$47218 ( \47595 , \47593 );
and \U$47219 ( \47596 , \47595 , \1734 );
nor \U$47220 ( \47597 , \47594 , \47596 );
xor \U$47221 ( \47598 , \47590 , \47597 );
and \U$47222 ( \47599 , \2224 , RIae78080_102);
and \U$47223 ( \47600 , RIae78260_106, \2222 );
nor \U$47224 ( \47601 , \47599 , \47600 );
and \U$47225 ( \47602 , \47601 , \2061 );
not \U$47226 ( \47603 , \47601 );
and \U$47227 ( \47604 , \47603 , \2060 );
nor \U$47228 ( \47605 , \47602 , \47604 );
and \U$47229 ( \47606 , \47598 , \47605 );
and \U$47230 ( \47607 , \47590 , \47597 );
or \U$47231 ( \47608 , \47606 , \47607 );
xor \U$47232 ( \47609 , \47583 , \47608 );
and \U$47233 ( \47610 , \1376 , RIae77090_68);
and \U$47234 ( \47611 , RIae77270_72, \1374 );
nor \U$47235 ( \47612 , \47610 , \47611 );
and \U$47236 ( \47613 , \47612 , \1380 );
not \U$47237 ( \47614 , \47612 );
and \U$47238 ( \47615 , \47614 , \1261 );
nor \U$47239 ( \47616 , \47613 , \47615 );
and \U$47240 ( \47617 , \1138 , RIae76cd0_60);
and \U$47241 ( \47618 , RIae77108_69, \1136 );
nor \U$47242 ( \47619 , \47617 , \47618 );
and \U$47243 ( \47620 , \47619 , \1012 );
not \U$47244 ( \47621 , \47619 );
and \U$47245 ( \47622 , \47621 , \1142 );
nor \U$47246 ( \47623 , \47620 , \47622 );
xor \U$47247 ( \47624 , \47616 , \47623 );
and \U$47248 ( \47625 , \1593 , RIae77360_74);
and \U$47249 ( \47626 , RIae78350_108, \1591 );
nor \U$47250 ( \47627 , \47625 , \47626 );
and \U$47251 ( \47628 , \47627 , \1498 );
not \U$47252 ( \47629 , \47627 );
and \U$47253 ( \47630 , \47629 , \1488 );
nor \U$47254 ( \47631 , \47628 , \47630 );
and \U$47255 ( \47632 , \47624 , \47631 );
and \U$47256 ( \47633 , \47616 , \47623 );
or \U$47257 ( \47634 , \47632 , \47633 );
and \U$47258 ( \47635 , \47609 , \47634 );
and \U$47259 ( \47636 , \47583 , \47608 );
or \U$47260 ( \47637 , \47635 , \47636 );
and \U$47261 ( \47638 , \11470 , RIae76640_46);
and \U$47262 ( \47639 , RIae76190_36, \11468 );
nor \U$47263 ( \47640 , \47638 , \47639 );
and \U$47264 ( \47641 , \47640 , \10936 );
not \U$47265 ( \47642 , \47640 );
and \U$47266 ( \47643 , \47642 , \11474 );
nor \U$47267 ( \47644 , \47641 , \47643 );
and \U$47268 ( \47645 , \9760 , RIae75470_8);
and \U$47269 ( \47646 , RIae76460_42, \9758 );
nor \U$47270 ( \47647 , \47645 , \47646 );
and \U$47271 ( \47648 , \47647 , \9273 );
not \U$47272 ( \47649 , \47647 );
and \U$47273 ( \47650 , \47649 , \9764 );
nor \U$47274 ( \47651 , \47648 , \47650 );
xor \U$47275 ( \47652 , \47644 , \47651 );
and \U$47276 ( \47653 , \10548 , RIae76550_44);
and \U$47277 ( \47654 , RIae76730_48, \10546 );
nor \U$47278 ( \47655 , \47653 , \47654 );
and \U$47279 ( \47656 , \47655 , \10421 );
not \U$47280 ( \47657 , \47655 );
and \U$47281 ( \47658 , \47657 , \10118 );
nor \U$47282 ( \47659 , \47656 , \47658 );
and \U$47283 ( \47660 , \47652 , \47659 );
and \U$47284 ( \47661 , \47644 , \47651 );
or \U$47285 ( \47662 , \47660 , \47661 );
and \U$47286 ( \47663 , \15726 , RIae78ad0_124);
and \U$47287 ( \47664 , RIae78d28_129, RIae7aab0_192);
nor \U$47288 ( \47665 , \47663 , \47664 );
and \U$47289 ( \47666 , \47665 , \14959 );
not \U$47290 ( \47667 , \47665 );
and \U$47291 ( \47668 , \47667 , RIae7aa38_191);
nor \U$47292 ( \47669 , \47666 , \47668 );
xor \U$47293 ( \47670 , \47669 , \392 );
and \U$47294 ( \47671 , \14964 , RIae76910_52);
and \U$47295 ( \47672 , RIae76be0_58, \14962 );
nor \U$47296 ( \47673 , \47671 , \47672 );
and \U$47297 ( \47674 , \47673 , \14463 );
not \U$47298 ( \47675 , \47673 );
and \U$47299 ( \47676 , \47675 , \14462 );
nor \U$47300 ( \47677 , \47674 , \47676 );
and \U$47301 ( \47678 , \47670 , \47677 );
and \U$47302 ( \47679 , \47669 , \392 );
or \U$47303 ( \47680 , \47678 , \47679 );
xor \U$47304 ( \47681 , \47662 , \47680 );
and \U$47305 ( \47682 , \14059 , RIae76a00_54);
and \U$47306 ( \47683 , RIae76820_50, \14057 );
nor \U$47307 ( \47684 , \47682 , \47683 );
and \U$47308 ( \47685 , \47684 , \13502 );
not \U$47309 ( \47686 , \47684 );
and \U$47310 ( \47687 , \47686 , \14063 );
nor \U$47311 ( \47688 , \47685 , \47687 );
and \U$47312 ( \47689 , \12180 , RIae760a0_34);
and \U$47313 ( \47690 , RIae76370_40, \12178 );
nor \U$47314 ( \47691 , \47689 , \47690 );
and \U$47315 ( \47692 , \47691 , \12184 );
not \U$47316 ( \47693 , \47691 );
and \U$47317 ( \47694 , \47693 , \11827 );
nor \U$47318 ( \47695 , \47692 , \47694 );
xor \U$47319 ( \47696 , \47688 , \47695 );
and \U$47320 ( \47697 , \13059 , RIae76280_38);
and \U$47321 ( \47698 , RIae76af0_56, \13057 );
nor \U$47322 ( \47699 , \47697 , \47698 );
and \U$47323 ( \47700 , \47699 , \13063 );
not \U$47324 ( \47701 , \47699 );
and \U$47325 ( \47702 , \47701 , \12718 );
nor \U$47326 ( \47703 , \47700 , \47702 );
and \U$47327 ( \47704 , \47696 , \47703 );
and \U$47328 ( \47705 , \47688 , \47695 );
or \U$47329 ( \47706 , \47704 , \47705 );
and \U$47330 ( \47707 , \47681 , \47706 );
and \U$47331 ( \47708 , \47662 , \47680 );
or \U$47332 ( \47709 , \47707 , \47708 );
xor \U$47333 ( \47710 , \47637 , \47709 );
and \U$47334 ( \47711 , \6172 , RIae75ec0_30);
and \U$47335 ( \47712 , RIae75ce0_26, \6170 );
nor \U$47336 ( \47713 , \47711 , \47712 );
and \U$47337 ( \47714 , \47713 , \6176 );
not \U$47338 ( \47715 , \47713 );
and \U$47339 ( \47716 , \47715 , \6175 );
nor \U$47340 ( \47717 , \47714 , \47716 );
and \U$47341 ( \47718 , \5896 , RIae75920_18);
and \U$47342 ( \47719 , RIae75fb0_32, \5894 );
nor \U$47343 ( \47720 , \47718 , \47719 );
and \U$47344 ( \47721 , \47720 , \5590 );
not \U$47345 ( \47722 , \47720 );
and \U$47346 ( \47723 , \47722 , \5589 );
nor \U$47347 ( \47724 , \47721 , \47723 );
xor \U$47348 ( \47725 , \47717 , \47724 );
and \U$47349 ( \47726 , \6941 , RIae75dd0_28);
and \U$47350 ( \47727 , RIae75650_12, \6939 );
nor \U$47351 ( \47728 , \47726 , \47727 );
and \U$47352 ( \47729 , \47728 , \6314 );
not \U$47353 ( \47730 , \47728 );
and \U$47354 ( \47731 , \47730 , \6945 );
nor \U$47355 ( \47732 , \47729 , \47731 );
and \U$47356 ( \47733 , \47725 , \47732 );
and \U$47357 ( \47734 , \47717 , \47724 );
or \U$47358 ( \47735 , \47733 , \47734 );
and \U$47359 ( \47736 , \4247 , RIae788f0_120);
and \U$47360 ( \47737 , RIae78800_118, \4245 );
nor \U$47361 ( \47738 , \47736 , \47737 );
and \U$47362 ( \47739 , \47738 , \3989 );
not \U$47363 ( \47740 , \47738 );
and \U$47364 ( \47741 , \47740 , \4251 );
nor \U$47365 ( \47742 , \47739 , \47741 );
and \U$47366 ( \47743 , \4688 , RIae78710_116);
and \U$47367 ( \47744 , RIae75bf0_24, \4686 );
nor \U$47368 ( \47745 , \47743 , \47744 );
and \U$47369 ( \47746 , \47745 , \4481 );
not \U$47370 ( \47747 , \47745 );
and \U$47371 ( \47748 , \47747 , \4482 );
nor \U$47372 ( \47749 , \47746 , \47748 );
xor \U$47373 ( \47750 , \47742 , \47749 );
and \U$47374 ( \47751 , \5399 , RIae75b00_22);
and \U$47375 ( \47752 , RIae75a10_20, \5397 );
nor \U$47376 ( \47753 , \47751 , \47752 );
and \U$47377 ( \47754 , \47753 , \5016 );
not \U$47378 ( \47755 , \47753 );
and \U$47379 ( \47756 , \47755 , \5403 );
nor \U$47380 ( \47757 , \47754 , \47756 );
and \U$47381 ( \47758 , \47750 , \47757 );
and \U$47382 ( \47759 , \47742 , \47749 );
or \U$47383 ( \47760 , \47758 , \47759 );
xor \U$47384 ( \47761 , \47735 , \47760 );
and \U$47385 ( \47762 , \8966 , RIae751a0_2);
and \U$47386 ( \47763 , RIae75380_6, \8964 );
nor \U$47387 ( \47764 , \47762 , \47763 );
and \U$47388 ( \47765 , \47764 , \8799 );
not \U$47389 ( \47766 , \47764 );
and \U$47390 ( \47767 , \47766 , \8789 );
nor \U$47391 ( \47768 , \47765 , \47767 );
and \U$47392 ( \47769 , \7633 , RIae75560_10);
and \U$47393 ( \47770 , RIae75830_16, \7631 );
nor \U$47394 ( \47771 , \47769 , \47770 );
and \U$47395 ( \47772 , \47771 , \7206 );
not \U$47396 ( \47773 , \47771 );
and \U$47397 ( \47774 , \47773 , \7205 );
nor \U$47398 ( \47775 , \47772 , \47774 );
xor \U$47399 ( \47776 , \47768 , \47775 );
and \U$47400 ( \47777 , \8371 , RIae75740_14);
and \U$47401 ( \47778 , RIae75290_4, \8369 );
nor \U$47402 ( \47779 , \47777 , \47778 );
and \U$47403 ( \47780 , \47779 , \8020 );
not \U$47404 ( \47781 , \47779 );
and \U$47405 ( \47782 , \47781 , \8019 );
nor \U$47406 ( \47783 , \47780 , \47782 );
and \U$47407 ( \47784 , \47776 , \47783 );
and \U$47408 ( \47785 , \47768 , \47775 );
or \U$47409 ( \47786 , \47784 , \47785 );
and \U$47410 ( \47787 , \47761 , \47786 );
and \U$47411 ( \47788 , \47735 , \47760 );
or \U$47412 ( \47789 , \47787 , \47788 );
and \U$47413 ( \47790 , \47710 , \47789 );
and \U$47414 ( \47791 , \47637 , \47709 );
nor \U$47415 ( \47792 , \47790 , \47791 );
not \U$47416 ( \47793 , \47792 );
xor \U$47417 ( \47794 , \47231 , \47238 );
xor \U$47418 ( \47795 , \47794 , \47246 );
not \U$47419 ( \47796 , \47795 );
not \U$47420 ( \47797 , \47257 );
xor \U$47421 ( \47798 , \47265 , \47275 );
not \U$47422 ( \47799 , \47798 );
or \U$47423 ( \47800 , \47797 , \47799 );
or \U$47424 ( \47801 , \47798 , \47257 );
nand \U$47425 ( \47802 , \47800 , \47801 );
nand \U$47426 ( \47803 , \47796 , \47802 );
not \U$47427 ( \47804 , \46712 );
not \U$47428 ( \47805 , \46715 );
and \U$47429 ( \47806 , \47804 , \47805 );
and \U$47430 ( \47807 , \46712 , \46715 );
nor \U$47431 ( \47808 , \47806 , \47807 );
xor \U$47432 ( \47809 , \47803 , \47808 );
not \U$47433 ( \47810 , \47288 );
xor \U$47434 ( \47811 , \47296 , \47306 );
not \U$47435 ( \47812 , \47811 );
or \U$47436 ( \47813 , \47810 , \47812 );
or \U$47437 ( \47814 , \47811 , \47288 );
nand \U$47438 ( \47815 , \47813 , \47814 );
not \U$47439 ( \47816 , \47341 );
xor \U$47440 ( \47817 , \47349 , \47359 );
not \U$47441 ( \47818 , \47817 );
or \U$47442 ( \47819 , \47816 , \47818 );
or \U$47443 ( \47820 , \47817 , \47341 );
nand \U$47444 ( \47821 , \47819 , \47820 );
xor \U$47445 ( \47822 , \47815 , \47821 );
not \U$47446 ( \47823 , \47204 );
xor \U$47447 ( \47824 , \47222 , \47212 );
not \U$47448 ( \47825 , \47824 );
or \U$47449 ( \47826 , \47823 , \47825 );
or \U$47450 ( \47827 , \47824 , \47204 );
nand \U$47451 ( \47828 , \47826 , \47827 );
and \U$47452 ( \47829 , \47822 , \47828 );
and \U$47453 ( \47830 , \47815 , \47821 );
nor \U$47454 ( \47831 , \47829 , \47830 );
and \U$47455 ( \47832 , \47809 , \47831 );
and \U$47456 ( \47833 , \47803 , \47808 );
or \U$47457 ( \47834 , \47832 , \47833 );
not \U$47458 ( \47835 , \47834 );
and \U$47459 ( \47836 , \47793 , \47835 );
and \U$47460 ( \47837 , \47792 , \47834 );
not \U$47461 ( \47838 , \47116 );
xor \U$47462 ( \47839 , \47125 , \47136 );
not \U$47463 ( \47840 , \47839 );
or \U$47464 ( \47841 , \47838 , \47840 );
or \U$47465 ( \47842 , \47839 , \47116 );
nand \U$47466 ( \47843 , \47841 , \47842 );
xor \U$47467 ( \47844 , \47315 , \47322 );
xor \U$47468 ( \47845 , \47844 , \47330 );
xor \U$47469 ( \47846 , \47843 , \47845 );
not \U$47470 ( \47847 , \47145 );
xor \U$47471 ( \47848 , \47163 , \47153 );
not \U$47472 ( \47849 , \47848 );
or \U$47473 ( \47850 , \47847 , \47849 );
or \U$47474 ( \47851 , \47848 , \47145 );
nand \U$47475 ( \47852 , \47850 , \47851 );
and \U$47476 ( \47853 , \47846 , \47852 );
and \U$47477 ( \47854 , \47843 , \47845 );
nor \U$47478 ( \47855 , \47853 , \47854 );
not \U$47479 ( \47856 , \47855 );
and \U$47480 ( \47857 , \514 , RIae77450_76);
and \U$47481 ( \47858 , RIae77ae0_90, \512 );
nor \U$47482 ( \47859 , \47857 , \47858 );
not \U$47483 ( \47860 , \47859 );
not \U$47484 ( \47861 , \471 );
and \U$47485 ( \47862 , \47860 , \47861 );
and \U$47486 ( \47863 , \47859 , \469 );
nor \U$47487 ( \47864 , \47862 , \47863 );
not \U$47488 ( \47865 , \47864 );
not \U$47489 ( \47866 , \388 );
nand \U$47490 ( \47867 , RIae77630_80, \382 );
not \U$47491 ( \47868 , \47867 );
and \U$47492 ( \47869 , \47866 , \47868 );
and \U$47493 ( \47870 , \388 , \47867 );
nor \U$47494 ( \47871 , \47869 , \47870 );
not \U$47495 ( \47872 , \47871 );
and \U$47496 ( \47873 , \47865 , \47872 );
and \U$47497 ( \47874 , \47864 , \47871 );
and \U$47498 ( \47875 , \436 , RIae77540_78);
and \U$47499 ( \47876 , RIae776a8_81, \434 );
nor \U$47500 ( \47877 , \47875 , \47876 );
not \U$47501 ( \47878 , \47877 );
not \U$47502 ( \47879 , \400 );
and \U$47503 ( \47880 , \47878 , \47879 );
and \U$47504 ( \47881 , \47877 , \400 );
nor \U$47505 ( \47882 , \47880 , \47881 );
nor \U$47506 ( \47883 , \47874 , \47882 );
nor \U$47507 ( \47884 , \47873 , \47883 );
not \U$47508 ( \47885 , \47884 );
and \U$47509 ( \47886 , \436 , RIae776a8_81);
and \U$47510 ( \47887 , RIae77450_76, \434 );
nor \U$47511 ( \47888 , \47886 , \47887 );
not \U$47512 ( \47889 , \47888 );
not \U$47513 ( \47890 , \400 );
and \U$47514 ( \47891 , \47889 , \47890 );
and \U$47515 ( \47892 , \47888 , \400 );
nor \U$47516 ( \47893 , \47891 , \47892 );
not \U$47517 ( \47894 , \47893 );
and \U$47518 ( \47895 , \47885 , \47894 );
and \U$47519 ( \47896 , \47884 , \47893 );
and \U$47520 ( \47897 , \558 , RIae779f0_88);
and \U$47521 ( \47898 , RIae77810_84, \556 );
nor \U$47522 ( \47899 , \47897 , \47898 );
and \U$47523 ( \47900 , \47899 , \562 );
not \U$47524 ( \47901 , \47899 );
and \U$47525 ( \47902 , \47901 , \504 );
nor \U$47526 ( \47903 , \47900 , \47902 );
not \U$47527 ( \47904 , \47903 );
and \U$47528 ( \47905 , \883 , RIae76eb0_64);
and \U$47529 ( \47906 , RIae76dc0_62, \881 );
nor \U$47530 ( \47907 , \47905 , \47906 );
not \U$47531 ( \47908 , \47907 );
not \U$47532 ( \47909 , \789 );
and \U$47533 ( \47910 , \47908 , \47909 );
and \U$47534 ( \47911 , \47907 , \787 );
nor \U$47535 ( \47912 , \47910 , \47911 );
not \U$47536 ( \47913 , \47912 );
and \U$47537 ( \47914 , \47904 , \47913 );
and \U$47538 ( \47915 , \47912 , \47903 );
and \U$47539 ( \47916 , \672 , RIae77900_86);
and \U$47540 ( \47917 , RIae76fa0_66, \670 );
nor \U$47541 ( \47918 , \47916 , \47917 );
and \U$47542 ( \47919 , \47918 , \587 );
not \U$47543 ( \47920 , \47918 );
and \U$47544 ( \47921 , \47920 , \588 );
nor \U$47545 ( \47922 , \47919 , \47921 );
nor \U$47546 ( \47923 , \47915 , \47922 );
nor \U$47547 ( \47924 , \47914 , \47923 );
nor \U$47548 ( \47925 , \47896 , \47924 );
nor \U$47549 ( \47926 , \47895 , \47925 );
not \U$47550 ( \47927 , \47926 );
and \U$47551 ( \47928 , \47856 , \47927 );
and \U$47552 ( \47929 , \47855 , \47926 );
not \U$47553 ( \47930 , \47393 );
xor \U$47554 ( \47931 , \47411 , \47401 );
not \U$47555 ( \47932 , \47931 );
or \U$47556 ( \47933 , \47930 , \47932 );
or \U$47557 ( \47934 , \47931 , \47393 );
nand \U$47558 ( \47935 , \47933 , \47934 );
not \U$47559 ( \47936 , \392 );
and \U$47560 ( \47937 , \384 , RIae77630_80);
and \U$47561 ( \47938 , RIae77540_78, \382 );
nor \U$47562 ( \47939 , \47937 , \47938 );
not \U$47563 ( \47940 , \47939 );
or \U$47564 ( \47941 , \47936 , \47940 );
or \U$47565 ( \47942 , \47939 , \392 );
nand \U$47566 ( \47943 , \47941 , \47942 );
xor \U$47567 ( \47944 , \47935 , \47943 );
not \U$47568 ( \47945 , \47174 );
xor \U$47569 ( \47946 , \47182 , \47192 );
not \U$47570 ( \47947 , \47946 );
or \U$47571 ( \47948 , \47945 , \47947 );
or \U$47572 ( \47949 , \47946 , \47174 );
nand \U$47573 ( \47950 , \47948 , \47949 );
and \U$47574 ( \47951 , \47944 , \47950 );
and \U$47575 ( \47952 , \47935 , \47943 );
or \U$47576 ( \47953 , \47951 , \47952 );
not \U$47577 ( \47954 , \47953 );
nor \U$47578 ( \47955 , \47929 , \47954 );
nor \U$47579 ( \47956 , \47928 , \47955 );
nor \U$47580 ( \47957 , \47837 , \47956 );
nor \U$47581 ( \47958 , \47836 , \47957 );
xor \U$47582 ( \47959 , \47377 , \47379 );
xor \U$47583 ( \47960 , \47959 , \47382 );
xor \U$47584 ( \47961 , \47439 , \47449 );
xor \U$47585 ( \47962 , \47961 , \47452 );
and \U$47586 ( \47963 , \47960 , \47962 );
xor \U$47587 ( \47964 , \46658 , \46666 );
xor \U$47588 ( \47965 , \47964 , \46674 );
xor \U$47589 ( \47966 , \47423 , \47428 );
xor \U$47590 ( \47967 , \47965 , \47966 );
xor \U$47591 ( \47968 , \47439 , \47449 );
xor \U$47592 ( \47969 , \47968 , \47452 );
and \U$47593 ( \47970 , \47967 , \47969 );
and \U$47594 ( \47971 , \47960 , \47967 );
or \U$47595 ( \47972 , \47963 , \47970 , \47971 );
xor \U$47596 ( \47973 , \47413 , \47414 );
xor \U$47597 ( \47974 , \47973 , \47417 );
xor \U$47598 ( \47975 , \47308 , \47333 );
xor \U$47599 ( \47976 , \47975 , \47361 );
and \U$47600 ( \47977 , \47974 , \47976 );
xor \U$47601 ( \47978 , \47138 , \47165 );
xor \U$47602 ( \47979 , \47978 , \47194 );
xor \U$47603 ( \47980 , \47308 , \47333 );
xor \U$47604 ( \47981 , \47980 , \47361 );
and \U$47605 ( \47982 , \47979 , \47981 );
and \U$47606 ( \47983 , \47974 , \47979 );
or \U$47607 ( \47984 , \47977 , \47982 , \47983 );
xor \U$47608 ( \47985 , \47972 , \47984 );
xor \U$47609 ( \47986 , \47063 , \47073 );
xor \U$47610 ( \47987 , \47986 , \47076 );
and \U$47611 ( \47988 , \47985 , \47987 );
and \U$47612 ( \47989 , \47972 , \47984 );
or \U$47613 ( \47990 , \47988 , \47989 );
xor \U$47614 ( \47991 , \47958 , \47990 );
not \U$47615 ( \47992 , \47095 );
not \U$47616 ( \47993 , \47105 );
or \U$47617 ( \47994 , \47992 , \47993 );
or \U$47618 ( \47995 , \47105 , \47095 );
nand \U$47619 ( \47996 , \47994 , \47995 );
not \U$47620 ( \47997 , \47996 );
not \U$47621 ( \47998 , \47097 );
and \U$47622 ( \47999 , \47997 , \47998 );
and \U$47623 ( \48000 , \47996 , \47097 );
nor \U$47624 ( \48001 , \47999 , \48000 );
xor \U$47625 ( \48002 , \47385 , \47420 );
xor \U$47626 ( \48003 , \48002 , \47433 );
xor \U$47627 ( \48004 , \48001 , \48003 );
xor \U$47628 ( \48005 , \47455 , \47460 );
xor \U$47629 ( \48006 , \48005 , \47463 );
and \U$47630 ( \48007 , \48004 , \48006 );
and \U$47631 ( \48008 , \48001 , \48003 );
or \U$47632 ( \48009 , \48007 , \48008 );
and \U$47633 ( \48010 , \47991 , \48009 );
and \U$47634 ( \48011 , \47958 , \47990 );
nor \U$47635 ( \48012 , \48010 , \48011 );
and \U$47636 ( \48013 , \47556 , \48012 );
and \U$47637 ( \48014 , \47553 , \47555 );
or \U$47638 ( \48015 , \48013 , \48014 );
nand \U$47639 ( \48016 , \47539 , \48015 );
nand \U$47640 ( \48017 , \47538 , \48016 );
nand \U$47641 ( \48018 , \47532 , \48017 );
nand \U$47642 ( \48019 , \47531 , \48018 );
and \U$47643 ( \48020 , \47525 , \48019 );
xor \U$47644 ( \48021 , \48019 , \47525 );
not \U$47645 ( \48022 , \47855 );
not \U$47646 ( \48023 , \47926 );
not \U$47647 ( \48024 , \47953 );
or \U$47648 ( \48025 , \48023 , \48024 );
or \U$47649 ( \48026 , \47953 , \47926 );
nand \U$47650 ( \48027 , \48025 , \48026 );
not \U$47651 ( \48028 , \48027 );
or \U$47652 ( \48029 , \48022 , \48028 );
or \U$47653 ( \48030 , \48027 , \47855 );
nand \U$47654 ( \48031 , \48029 , \48030 );
xor \U$47655 ( \48032 , \47637 , \47709 );
xor \U$47656 ( \48033 , \48032 , \47789 );
xor \U$47657 ( \48034 , \48031 , \48033 );
xor \U$47658 ( \48035 , \47803 , \47808 );
xor \U$47659 ( \48036 , \48035 , \47831 );
not \U$47660 ( \48037 , \48036 );
xor \U$47661 ( \48038 , \47308 , \47333 );
xor \U$47662 ( \48039 , \48038 , \47361 );
xor \U$47663 ( \48040 , \47974 , \47979 );
xor \U$47664 ( \48041 , \48039 , \48040 );
xor \U$47665 ( \48042 , \47439 , \47449 );
xor \U$47666 ( \48043 , \48042 , \47452 );
xor \U$47667 ( \48044 , \47960 , \47967 );
xor \U$47668 ( \48045 , \48043 , \48044 );
xor \U$47669 ( \48046 , \48041 , \48045 );
not \U$47670 ( \48047 , \48046 );
or \U$47671 ( \48048 , \48037 , \48047 );
or \U$47672 ( \48049 , \48046 , \48036 );
nand \U$47673 ( \48050 , \48048 , \48049 );
and \U$47674 ( \48051 , \48034 , \48050 );
and \U$47675 ( \48052 , \48031 , \48033 );
or \U$47676 ( \48053 , \48051 , \48052 );
not \U$47677 ( \48054 , \47834 );
xor \U$47678 ( \48055 , \47792 , \47956 );
not \U$47679 ( \48056 , \48055 );
or \U$47680 ( \48057 , \48054 , \48056 );
or \U$47681 ( \48058 , \48055 , \47834 );
nand \U$47682 ( \48059 , \48057 , \48058 );
xor \U$47683 ( \48060 , \48053 , \48059 );
xor \U$47684 ( \48061 , \47742 , \47749 );
xor \U$47685 ( \48062 , \48061 , \47757 );
xor \U$47686 ( \48063 , \47717 , \47724 );
xor \U$47687 ( \48064 , \48063 , \47732 );
and \U$47688 ( \48065 , \48062 , \48064 );
xor \U$47689 ( \48066 , \47768 , \47775 );
xor \U$47690 ( \48067 , \48066 , \47783 );
xor \U$47691 ( \48068 , \47717 , \47724 );
xor \U$47692 ( \48069 , \48068 , \47732 );
and \U$47693 ( \48070 , \48067 , \48069 );
and \U$47694 ( \48071 , \48062 , \48067 );
or \U$47695 ( \48072 , \48065 , \48070 , \48071 );
not \U$47696 ( \48073 , \47871 );
xor \U$47697 ( \48074 , \47882 , \47864 );
not \U$47698 ( \48075 , \48074 );
or \U$47699 ( \48076 , \48073 , \48075 );
or \U$47700 ( \48077 , \48074 , \47871 );
nand \U$47701 ( \48078 , \48076 , \48077 );
not \U$47702 ( \48079 , \469 );
and \U$47703 ( \48080 , \514 , RIae776a8_81);
and \U$47704 ( \48081 , RIae77450_76, \512 );
nor \U$47705 ( \48082 , \48080 , \48081 );
not \U$47706 ( \48083 , \48082 );
or \U$47707 ( \48084 , \48079 , \48083 );
or \U$47708 ( \48085 , \48082 , \471 );
nand \U$47709 ( \48086 , \48084 , \48085 );
and \U$47710 ( \48087 , \558 , RIae77ae0_90);
and \U$47711 ( \48088 , RIae779f0_88, \556 );
nor \U$47712 ( \48089 , \48087 , \48088 );
and \U$47713 ( \48090 , \48089 , \504 );
not \U$47714 ( \48091 , \48089 );
and \U$47715 ( \48092 , \48091 , \562 );
nor \U$47716 ( \48093 , \48090 , \48092 );
xor \U$47717 ( \48094 , \48086 , \48093 );
and \U$47718 ( \48095 , \672 , RIae77810_84);
and \U$47719 ( \48096 , RIae77900_86, \670 );
nor \U$47720 ( \48097 , \48095 , \48096 );
and \U$47721 ( \48098 , \48097 , \588 );
not \U$47722 ( \48099 , \48097 );
and \U$47723 ( \48100 , \48099 , \587 );
nor \U$47724 ( \48101 , \48098 , \48100 );
and \U$47725 ( \48102 , \48094 , \48101 );
and \U$47726 ( \48103 , \48086 , \48093 );
or \U$47727 ( \48104 , \48102 , \48103 );
xor \U$47728 ( \48105 , \48078 , \48104 );
not \U$47729 ( \48106 , \47903 );
xor \U$47730 ( \48107 , \47922 , \47912 );
not \U$47731 ( \48108 , \48107 );
or \U$47732 ( \48109 , \48106 , \48108 );
or \U$47733 ( \48110 , \48107 , \47903 );
nand \U$47734 ( \48111 , \48109 , \48110 );
and \U$47735 ( \48112 , \48105 , \48111 );
and \U$47736 ( \48113 , \48078 , \48104 );
or \U$47737 ( \48114 , \48112 , \48113 );
xor \U$47738 ( \48115 , \48072 , \48114 );
xor \U$47739 ( \48116 , \47616 , \47623 );
xor \U$47740 ( \48117 , \48116 , \47631 );
xor \U$47741 ( \48118 , \47590 , \47597 );
xor \U$47742 ( \48119 , \48118 , \47605 );
and \U$47743 ( \48120 , \48117 , \48119 );
xor \U$47744 ( \48121 , \47564 , \47572 );
xor \U$47745 ( \48122 , \48121 , \47580 );
xor \U$47746 ( \48123 , \47590 , \47597 );
xor \U$47747 ( \48124 , \48123 , \47605 );
and \U$47748 ( \48125 , \48122 , \48124 );
and \U$47749 ( \48126 , \48117 , \48122 );
or \U$47750 ( \48127 , \48120 , \48125 , \48126 );
xor \U$47751 ( \48128 , \48115 , \48127 );
and \U$47752 ( \48129 , \2224 , RIae77f90_100);
and \U$47753 ( \48130 , RIae78080_102, \2222 );
nor \U$47754 ( \48131 , \48129 , \48130 );
and \U$47755 ( \48132 , \48131 , \2061 );
not \U$47756 ( \48133 , \48131 );
and \U$47757 ( \48134 , \48133 , \2060 );
nor \U$47758 ( \48135 , \48132 , \48134 );
and \U$47759 ( \48136 , \1593 , RIae77270_72);
and \U$47760 ( \48137 , RIae77360_74, \1591 );
nor \U$47761 ( \48138 , \48136 , \48137 );
and \U$47762 ( \48139 , \48138 , \1498 );
not \U$47763 ( \48140 , \48138 );
and \U$47764 ( \48141 , \48140 , \1488 );
nor \U$47765 ( \48142 , \48139 , \48141 );
xor \U$47766 ( \48143 , \48135 , \48142 );
and \U$47767 ( \48144 , \1939 , RIae78350_108);
and \U$47768 ( \48145 , RIae78170_104, \1937 );
nor \U$47769 ( \48146 , \48144 , \48145 );
and \U$47770 ( \48147 , \48146 , \1735 );
not \U$47771 ( \48148 , \48146 );
and \U$47772 ( \48149 , \48148 , \1734 );
nor \U$47773 ( \48150 , \48147 , \48149 );
and \U$47774 ( \48151 , \48143 , \48150 );
and \U$47775 ( \48152 , \48135 , \48142 );
or \U$47776 ( \48153 , \48151 , \48152 );
not \U$47777 ( \48154 , \787 );
and \U$47778 ( \48155 , \883 , RIae76fa0_66);
and \U$47779 ( \48156 , RIae76eb0_64, \881 );
nor \U$47780 ( \48157 , \48155 , \48156 );
not \U$47781 ( \48158 , \48157 );
or \U$47782 ( \48159 , \48154 , \48158 );
or \U$47783 ( \48160 , \48157 , \789 );
nand \U$47784 ( \48161 , \48159 , \48160 );
and \U$47785 ( \48162 , \1138 , RIae76dc0_62);
and \U$47786 ( \48163 , RIae76cd0_60, \1136 );
nor \U$47787 ( \48164 , \48162 , \48163 );
and \U$47788 ( \48165 , \48164 , \1012 );
not \U$47789 ( \48166 , \48164 );
and \U$47790 ( \48167 , \48166 , \1142 );
nor \U$47791 ( \48168 , \48165 , \48167 );
xor \U$47792 ( \48169 , \48161 , \48168 );
and \U$47793 ( \48170 , \1376 , RIae77108_69);
and \U$47794 ( \48171 , RIae77090_68, \1374 );
nor \U$47795 ( \48172 , \48170 , \48171 );
and \U$47796 ( \48173 , \48172 , \1380 );
not \U$47797 ( \48174 , \48172 );
and \U$47798 ( \48175 , \48174 , \1261 );
nor \U$47799 ( \48176 , \48173 , \48175 );
and \U$47800 ( \48177 , \48169 , \48176 );
and \U$47801 ( \48178 , \48161 , \48168 );
or \U$47802 ( \48179 , \48177 , \48178 );
xor \U$47803 ( \48180 , \48153 , \48179 );
not \U$47804 ( \48181 , \3218 );
and \U$47805 ( \48182 , \3214 , RIae77cc0_94);
and \U$47806 ( \48183 , RIae77bd0_92, \3212 );
nor \U$47807 ( \48184 , \48182 , \48183 );
not \U$47808 ( \48185 , \48184 );
or \U$47809 ( \48186 , \48181 , \48185 );
or \U$47810 ( \48187 , \48184 , \2774 );
nand \U$47811 ( \48188 , \48186 , \48187 );
and \U$47812 ( \48189 , \2607 , RIae78260_106);
and \U$47813 ( \48190 , RIae78620_114, \2605 );
nor \U$47814 ( \48191 , \48189 , \48190 );
and \U$47815 ( \48192 , \48191 , \2611 );
not \U$47816 ( \48193 , \48191 );
and \U$47817 ( \48194 , \48193 , \2397 );
nor \U$47818 ( \48195 , \48192 , \48194 );
xor \U$47819 ( \48196 , \48188 , \48195 );
not \U$47820 ( \48197 , \2789 );
and \U$47821 ( \48198 , \2783 , RIae78440_110);
and \U$47822 ( \48199 , RIae784b8_111, \2781 );
nor \U$47823 ( \48200 , \48198 , \48199 );
not \U$47824 ( \48201 , \48200 );
or \U$47825 ( \48202 , \48197 , \48201 );
or \U$47826 ( \48203 , \48200 , \3089 );
nand \U$47827 ( \48204 , \48202 , \48203 );
and \U$47828 ( \48205 , \48196 , \48204 );
and \U$47829 ( \48206 , \48188 , \48195 );
or \U$47830 ( \48207 , \48205 , \48206 );
and \U$47831 ( \48208 , \48180 , \48207 );
and \U$47832 ( \48209 , \48153 , \48179 );
or \U$47833 ( \48210 , \48208 , \48209 );
and \U$47834 ( \48211 , \11470 , RIae76730_48);
and \U$47835 ( \48212 , RIae76640_46, \11468 );
nor \U$47836 ( \48213 , \48211 , \48212 );
and \U$47837 ( \48214 , \48213 , \10936 );
not \U$47838 ( \48215 , \48213 );
and \U$47839 ( \48216 , \48215 , \11474 );
nor \U$47840 ( \48217 , \48214 , \48216 );
and \U$47841 ( \48218 , \12180 , RIae76190_36);
and \U$47842 ( \48219 , RIae760a0_34, \12178 );
nor \U$47843 ( \48220 , \48218 , \48219 );
and \U$47844 ( \48221 , \48220 , \12184 );
not \U$47845 ( \48222 , \48220 );
and \U$47846 ( \48223 , \48222 , \11827 );
nor \U$47847 ( \48224 , \48221 , \48223 );
xor \U$47848 ( \48225 , \48217 , \48224 );
and \U$47849 ( \48226 , \13059 , RIae76370_40);
and \U$47850 ( \48227 , RIae76280_38, \13057 );
nor \U$47851 ( \48228 , \48226 , \48227 );
and \U$47852 ( \48229 , \48228 , \13063 );
not \U$47853 ( \48230 , \48228 );
and \U$47854 ( \48231 , \48230 , \12718 );
nor \U$47855 ( \48232 , \48229 , \48231 );
and \U$47856 ( \48233 , \48225 , \48232 );
and \U$47857 ( \48234 , \48217 , \48224 );
or \U$47858 ( \48235 , \48233 , \48234 );
and \U$47859 ( \48236 , \14964 , RIae76820_50);
and \U$47860 ( \48237 , RIae76910_52, \14962 );
nor \U$47861 ( \48238 , \48236 , \48237 );
and \U$47862 ( \48239 , \48238 , \14463 );
not \U$47863 ( \48240 , \48238 );
and \U$47864 ( \48241 , \48240 , \14462 );
nor \U$47865 ( \48242 , \48239 , \48241 );
and \U$47866 ( \48243 , \15726 , RIae76be0_58);
and \U$47867 ( \48244 , RIae78ad0_124, RIae7aab0_192);
nor \U$47868 ( \48245 , \48243 , \48244 );
and \U$47869 ( \48246 , \48245 , \14959 );
not \U$47870 ( \48247 , \48245 );
and \U$47871 ( \48248 , \48247 , RIae7aa38_191);
nor \U$47872 ( \48249 , \48246 , \48248 );
xor \U$47873 ( \48250 , \48242 , \48249 );
and \U$47874 ( \48251 , \14059 , RIae76af0_56);
and \U$47875 ( \48252 , RIae76a00_54, \14057 );
nor \U$47876 ( \48253 , \48251 , \48252 );
and \U$47877 ( \48254 , \48253 , \13502 );
not \U$47878 ( \48255 , \48253 );
and \U$47879 ( \48256 , \48255 , \14063 );
nor \U$47880 ( \48257 , \48254 , \48256 );
and \U$47881 ( \48258 , \48250 , \48257 );
and \U$47882 ( \48259 , \48242 , \48249 );
or \U$47883 ( \48260 , \48258 , \48259 );
xor \U$47884 ( \48261 , \48235 , \48260 );
and \U$47885 ( \48262 , \10548 , RIae76460_42);
and \U$47886 ( \48263 , RIae76550_44, \10546 );
nor \U$47887 ( \48264 , \48262 , \48263 );
and \U$47888 ( \48265 , \48264 , \10421 );
not \U$47889 ( \48266 , \48264 );
and \U$47890 ( \48267 , \48266 , \10118 );
nor \U$47891 ( \48268 , \48265 , \48267 );
and \U$47892 ( \48269 , \8966 , RIae75290_4);
and \U$47893 ( \48270 , RIae751a0_2, \8964 );
nor \U$47894 ( \48271 , \48269 , \48270 );
and \U$47895 ( \48272 , \48271 , \8799 );
not \U$47896 ( \48273 , \48271 );
and \U$47897 ( \48274 , \48273 , \8789 );
nor \U$47898 ( \48275 , \48272 , \48274 );
xor \U$47899 ( \48276 , \48268 , \48275 );
and \U$47900 ( \48277 , \9760 , RIae75380_6);
and \U$47901 ( \48278 , RIae75470_8, \9758 );
nor \U$47902 ( \48279 , \48277 , \48278 );
and \U$47903 ( \48280 , \48279 , \9273 );
not \U$47904 ( \48281 , \48279 );
and \U$47905 ( \48282 , \48281 , \9272 );
nor \U$47906 ( \48283 , \48280 , \48282 );
and \U$47907 ( \48284 , \48276 , \48283 );
and \U$47908 ( \48285 , \48268 , \48275 );
or \U$47909 ( \48286 , \48284 , \48285 );
and \U$47910 ( \48287 , \48261 , \48286 );
and \U$47911 ( \48288 , \48235 , \48260 );
or \U$47912 ( \48289 , \48287 , \48288 );
xor \U$47913 ( \48290 , \48210 , \48289 );
and \U$47914 ( \48291 , \8371 , RIae75830_16);
and \U$47915 ( \48292 , RIae75740_14, \8369 );
nor \U$47916 ( \48293 , \48291 , \48292 );
and \U$47917 ( \48294 , \48293 , \8020 );
not \U$47918 ( \48295 , \48293 );
and \U$47919 ( \48296 , \48295 , \8019 );
nor \U$47920 ( \48297 , \48294 , \48296 );
and \U$47921 ( \48298 , \6941 , RIae75ce0_26);
and \U$47922 ( \48299 , RIae75dd0_28, \6939 );
nor \U$47923 ( \48300 , \48298 , \48299 );
and \U$47924 ( \48301 , \48300 , \6314 );
not \U$47925 ( \48302 , \48300 );
and \U$47926 ( \48303 , \48302 , \6945 );
nor \U$47927 ( \48304 , \48301 , \48303 );
xor \U$47928 ( \48305 , \48297 , \48304 );
and \U$47929 ( \48306 , \7633 , RIae75650_12);
and \U$47930 ( \48307 , RIae75560_10, \7631 );
nor \U$47931 ( \48308 , \48306 , \48307 );
and \U$47932 ( \48309 , \48308 , \7206 );
not \U$47933 ( \48310 , \48308 );
and \U$47934 ( \48311 , \48310 , \7205 );
nor \U$47935 ( \48312 , \48309 , \48311 );
and \U$47936 ( \48313 , \48305 , \48312 );
and \U$47937 ( \48314 , \48297 , \48304 );
or \U$47938 ( \48315 , \48313 , \48314 );
and \U$47939 ( \48316 , \5896 , RIae75a10_20);
and \U$47940 ( \48317 , RIae75920_18, \5894 );
nor \U$47941 ( \48318 , \48316 , \48317 );
and \U$47942 ( \48319 , \48318 , \5590 );
not \U$47943 ( \48320 , \48318 );
and \U$47944 ( \48321 , \48320 , \5589 );
nor \U$47945 ( \48322 , \48319 , \48321 );
and \U$47946 ( \48323 , \5399 , RIae75bf0_24);
and \U$47947 ( \48324 , RIae75b00_22, \5397 );
nor \U$47948 ( \48325 , \48323 , \48324 );
and \U$47949 ( \48326 , \48325 , \5016 );
not \U$47950 ( \48327 , \48325 );
and \U$47951 ( \48328 , \48327 , \5403 );
nor \U$47952 ( \48329 , \48326 , \48328 );
xor \U$47953 ( \48330 , \48322 , \48329 );
and \U$47954 ( \48331 , \6172 , RIae75fb0_32);
and \U$47955 ( \48332 , RIae75ec0_30, \6170 );
nor \U$47956 ( \48333 , \48331 , \48332 );
and \U$47957 ( \48334 , \48333 , \6176 );
not \U$47958 ( \48335 , \48333 );
and \U$47959 ( \48336 , \48335 , \6175 );
nor \U$47960 ( \48337 , \48334 , \48336 );
and \U$47961 ( \48338 , \48330 , \48337 );
and \U$47962 ( \48339 , \48322 , \48329 );
or \U$47963 ( \48340 , \48338 , \48339 );
xor \U$47964 ( \48341 , \48315 , \48340 );
and \U$47965 ( \48342 , \4247 , RIae789e0_122);
and \U$47966 ( \48343 , RIae788f0_120, \4245 );
nor \U$47967 ( \48344 , \48342 , \48343 );
and \U$47968 ( \48345 , \48344 , \3989 );
not \U$47969 ( \48346 , \48344 );
and \U$47970 ( \48347 , \48346 , \4251 );
nor \U$47971 ( \48348 , \48345 , \48347 );
and \U$47972 ( \48349 , \3730 , RIae77db0_96);
and \U$47973 ( \48350 , RIae77ea0_98, \3728 );
nor \U$47974 ( \48351 , \48349 , \48350 );
and \U$47975 ( \48352 , \48351 , \3732 );
not \U$47976 ( \48353 , \48351 );
and \U$47977 ( \48354 , \48353 , \3422 );
nor \U$47978 ( \48355 , \48352 , \48354 );
xor \U$47979 ( \48356 , \48348 , \48355 );
and \U$47980 ( \48357 , \4688 , RIae78800_118);
and \U$47981 ( \48358 , RIae78710_116, \4686 );
nor \U$47982 ( \48359 , \48357 , \48358 );
and \U$47983 ( \48360 , \48359 , \4481 );
not \U$47984 ( \48361 , \48359 );
and \U$47985 ( \48362 , \48361 , \4482 );
nor \U$47986 ( \48363 , \48360 , \48362 );
and \U$47987 ( \48364 , \48356 , \48363 );
and \U$47988 ( \48365 , \48348 , \48355 );
or \U$47989 ( \48366 , \48364 , \48365 );
and \U$47990 ( \48367 , \48341 , \48366 );
and \U$47991 ( \48368 , \48315 , \48340 );
or \U$47992 ( \48369 , \48367 , \48368 );
xor \U$47993 ( \48370 , \48290 , \48369 );
xor \U$47994 ( \48371 , \48128 , \48370 );
xor \U$47995 ( \48372 , \47644 , \47651 );
xor \U$47996 ( \48373 , \48372 , \47659 );
xor \U$47997 ( \48374 , \47688 , \47695 );
xor \U$47998 ( \48375 , \48374 , \47703 );
xor \U$47999 ( \48376 , \48373 , \48375 );
xor \U$48000 ( \48377 , \47669 , \392 );
xor \U$48001 ( \48378 , \48377 , \47677 );
and \U$48002 ( \48379 , \48376 , \48378 );
and \U$48003 ( \48380 , \48373 , \48375 );
or \U$48004 ( \48381 , \48379 , \48380 );
not \U$48005 ( \48382 , \47802 );
not \U$48006 ( \48383 , \47795 );
or \U$48007 ( \48384 , \48382 , \48383 );
or \U$48008 ( \48385 , \47795 , \47802 );
nand \U$48009 ( \48386 , \48384 , \48385 );
xor \U$48010 ( \48387 , \48381 , \48386 );
xor \U$48011 ( \48388 , \47815 , \47821 );
xor \U$48012 ( \48389 , \48388 , \47828 );
xor \U$48013 ( \48390 , \48387 , \48389 );
and \U$48014 ( \48391 , \48371 , \48390 );
and \U$48015 ( \48392 , \48128 , \48370 );
or \U$48016 ( \48393 , \48391 , \48392 );
xor \U$48017 ( \48394 , \48086 , \48093 );
xor \U$48018 ( \48395 , \48394 , \48101 );
xor \U$48019 ( \48396 , \48161 , \48168 );
xor \U$48020 ( \48397 , \48396 , \48176 );
xor \U$48021 ( \48398 , \48395 , \48397 );
xor \U$48022 ( \48399 , \48135 , \48142 );
xor \U$48023 ( \48400 , \48399 , \48150 );
and \U$48024 ( \48401 , \48398 , \48400 );
and \U$48025 ( \48402 , \48395 , \48397 );
or \U$48026 ( \48403 , \48401 , \48402 );
nand \U$48027 ( \48404 , RIae77630_80, \434 );
not \U$48028 ( \48405 , \48404 );
not \U$48029 ( \48406 , \400 );
or \U$48030 ( \48407 , \48405 , \48406 );
or \U$48031 ( \48408 , \400 , \48404 );
nand \U$48032 ( \48409 , \48407 , \48408 );
not \U$48033 ( \48410 , \469 );
and \U$48034 ( \48411 , \514 , RIae77540_78);
and \U$48035 ( \48412 , RIae776a8_81, \512 );
nor \U$48036 ( \48413 , \48411 , \48412 );
not \U$48037 ( \48414 , \48413 );
or \U$48038 ( \48415 , \48410 , \48414 );
or \U$48039 ( \48416 , \48413 , \469 );
nand \U$48040 ( \48417 , \48415 , \48416 );
and \U$48041 ( \48418 , \48409 , \48417 );
not \U$48042 ( \48419 , \400 );
and \U$48043 ( \48420 , \436 , RIae77630_80);
and \U$48044 ( \48421 , RIae77540_78, \434 );
nor \U$48045 ( \48422 , \48420 , \48421 );
not \U$48046 ( \48423 , \48422 );
or \U$48047 ( \48424 , \48419 , \48423 );
or \U$48048 ( \48425 , \48422 , \402 );
nand \U$48049 ( \48426 , \48424 , \48425 );
xor \U$48050 ( \48427 , \48418 , \48426 );
not \U$48051 ( \48428 , \789 );
and \U$48052 ( \48429 , \883 , RIae77900_86);
and \U$48053 ( \48430 , RIae76fa0_66, \881 );
nor \U$48054 ( \48431 , \48429 , \48430 );
not \U$48055 ( \48432 , \48431 );
or \U$48056 ( \48433 , \48428 , \48432 );
or \U$48057 ( \48434 , \48431 , \789 );
nand \U$48058 ( \48435 , \48433 , \48434 );
and \U$48059 ( \48436 , \558 , RIae77450_76);
and \U$48060 ( \48437 , RIae77ae0_90, \556 );
nor \U$48061 ( \48438 , \48436 , \48437 );
and \U$48062 ( \48439 , \48438 , \504 );
not \U$48063 ( \48440 , \48438 );
and \U$48064 ( \48441 , \48440 , \562 );
nor \U$48065 ( \48442 , \48439 , \48441 );
xor \U$48066 ( \48443 , \48435 , \48442 );
and \U$48067 ( \48444 , \672 , RIae779f0_88);
and \U$48068 ( \48445 , RIae77810_84, \670 );
nor \U$48069 ( \48446 , \48444 , \48445 );
and \U$48070 ( \48447 , \48446 , \588 );
not \U$48071 ( \48448 , \48446 );
and \U$48072 ( \48449 , \48448 , \587 );
nor \U$48073 ( \48450 , \48447 , \48449 );
and \U$48074 ( \48451 , \48443 , \48450 );
and \U$48075 ( \48452 , \48435 , \48442 );
or \U$48076 ( \48453 , \48451 , \48452 );
and \U$48077 ( \48454 , \48427 , \48453 );
and \U$48078 ( \48455 , \48418 , \48426 );
or \U$48079 ( \48456 , \48454 , \48455 );
xor \U$48080 ( \48457 , \48403 , \48456 );
xor \U$48081 ( \48458 , \48188 , \48195 );
xor \U$48082 ( \48459 , \48458 , \48204 );
xor \U$48083 ( \48460 , \48322 , \48329 );
xor \U$48084 ( \48461 , \48460 , \48337 );
and \U$48085 ( \48462 , \48459 , \48461 );
xor \U$48086 ( \48463 , \48348 , \48355 );
xor \U$48087 ( \48464 , \48463 , \48363 );
xor \U$48088 ( \48465 , \48322 , \48329 );
xor \U$48089 ( \48466 , \48465 , \48337 );
and \U$48090 ( \48467 , \48464 , \48466 );
and \U$48091 ( \48468 , \48459 , \48464 );
or \U$48092 ( \48469 , \48462 , \48467 , \48468 );
and \U$48093 ( \48470 , \48457 , \48469 );
and \U$48094 ( \48471 , \48403 , \48456 );
or \U$48095 ( \48472 , \48470 , \48471 );
not \U$48096 ( \48473 , \3089 );
and \U$48097 ( \48474 , \2783 , RIae78620_114);
and \U$48098 ( \48475 , RIae78440_110, \2781 );
nor \U$48099 ( \48476 , \48474 , \48475 );
not \U$48100 ( \48477 , \48476 );
or \U$48101 ( \48478 , \48473 , \48477 );
or \U$48102 ( \48479 , \48476 , \2789 );
nand \U$48103 ( \48480 , \48478 , \48479 );
not \U$48104 ( \48481 , \2774 );
and \U$48105 ( \48482 , \3214 , RIae784b8_111);
and \U$48106 ( \48483 , RIae77cc0_94, \3212 );
nor \U$48107 ( \48484 , \48482 , \48483 );
not \U$48108 ( \48485 , \48484 );
or \U$48109 ( \48486 , \48481 , \48485 );
or \U$48110 ( \48487 , \48484 , \2774 );
nand \U$48111 ( \48488 , \48486 , \48487 );
xor \U$48112 ( \48489 , \48480 , \48488 );
and \U$48113 ( \48490 , \3730 , RIae77bd0_92);
and \U$48114 ( \48491 , RIae77db0_96, \3728 );
nor \U$48115 ( \48492 , \48490 , \48491 );
and \U$48116 ( \48493 , \48492 , \3732 );
not \U$48117 ( \48494 , \48492 );
and \U$48118 ( \48495 , \48494 , \3421 );
nor \U$48119 ( \48496 , \48493 , \48495 );
and \U$48120 ( \48497 , \48489 , \48496 );
and \U$48121 ( \48498 , \48480 , \48488 );
or \U$48122 ( \48499 , \48497 , \48498 );
and \U$48123 ( \48500 , \1138 , RIae76eb0_64);
and \U$48124 ( \48501 , RIae76dc0_62, \1136 );
nor \U$48125 ( \48502 , \48500 , \48501 );
and \U$48126 ( \48503 , \48502 , \1012 );
not \U$48127 ( \48504 , \48502 );
and \U$48128 ( \48505 , \48504 , \1142 );
nor \U$48129 ( \48506 , \48503 , \48505 );
and \U$48130 ( \48507 , \1376 , RIae76cd0_60);
and \U$48131 ( \48508 , RIae77108_69, \1374 );
nor \U$48132 ( \48509 , \48507 , \48508 );
and \U$48133 ( \48510 , \48509 , \1380 );
not \U$48134 ( \48511 , \48509 );
and \U$48135 ( \48512 , \48511 , \1261 );
nor \U$48136 ( \48513 , \48510 , \48512 );
xor \U$48137 ( \48514 , \48506 , \48513 );
and \U$48138 ( \48515 , \1593 , RIae77090_68);
and \U$48139 ( \48516 , RIae77270_72, \1591 );
nor \U$48140 ( \48517 , \48515 , \48516 );
and \U$48141 ( \48518 , \48517 , \1498 );
not \U$48142 ( \48519 , \48517 );
and \U$48143 ( \48520 , \48519 , \1488 );
nor \U$48144 ( \48521 , \48518 , \48520 );
and \U$48145 ( \48522 , \48514 , \48521 );
and \U$48146 ( \48523 , \48506 , \48513 );
or \U$48147 ( \48524 , \48522 , \48523 );
xor \U$48148 ( \48525 , \48499 , \48524 );
and \U$48149 ( \48526 , \2607 , RIae78080_102);
and \U$48150 ( \48527 , RIae78260_106, \2605 );
nor \U$48151 ( \48528 , \48526 , \48527 );
and \U$48152 ( \48529 , \48528 , \2611 );
not \U$48153 ( \48530 , \48528 );
and \U$48154 ( \48531 , \48530 , \2397 );
nor \U$48155 ( \48532 , \48529 , \48531 );
and \U$48156 ( \48533 , \1939 , RIae77360_74);
and \U$48157 ( \48534 , RIae78350_108, \1937 );
nor \U$48158 ( \48535 , \48533 , \48534 );
and \U$48159 ( \48536 , \48535 , \1735 );
not \U$48160 ( \48537 , \48535 );
and \U$48161 ( \48538 , \48537 , \1734 );
nor \U$48162 ( \48539 , \48536 , \48538 );
xor \U$48163 ( \48540 , \48532 , \48539 );
and \U$48164 ( \48541 , \2224 , RIae78170_104);
and \U$48165 ( \48542 , RIae77f90_100, \2222 );
nor \U$48166 ( \48543 , \48541 , \48542 );
and \U$48167 ( \48544 , \48543 , \2061 );
not \U$48168 ( \48545 , \48543 );
and \U$48169 ( \48546 , \48545 , \2060 );
nor \U$48170 ( \48547 , \48544 , \48546 );
and \U$48171 ( \48548 , \48540 , \48547 );
and \U$48172 ( \48549 , \48532 , \48539 );
or \U$48173 ( \48550 , \48548 , \48549 );
and \U$48174 ( \48551 , \48525 , \48550 );
and \U$48175 ( \48552 , \48499 , \48524 );
or \U$48176 ( \48553 , \48551 , \48552 );
and \U$48177 ( \48554 , \10548 , RIae75470_8);
and \U$48178 ( \48555 , RIae76460_42, \10546 );
nor \U$48179 ( \48556 , \48554 , \48555 );
and \U$48180 ( \48557 , \48556 , \10421 );
not \U$48181 ( \48558 , \48556 );
and \U$48182 ( \48559 , \48558 , \10118 );
nor \U$48183 ( \48560 , \48557 , \48559 );
and \U$48184 ( \48561 , \9760 , RIae751a0_2);
and \U$48185 ( \48562 , RIae75380_6, \9758 );
nor \U$48186 ( \48563 , \48561 , \48562 );
and \U$48187 ( \48564 , \48563 , \9273 );
not \U$48188 ( \48565 , \48563 );
and \U$48189 ( \48566 , \48565 , \9764 );
nor \U$48190 ( \48567 , \48564 , \48566 );
xor \U$48191 ( \48568 , \48560 , \48567 );
and \U$48192 ( \48569 , \11470 , RIae76550_44);
and \U$48193 ( \48570 , RIae76730_48, \11468 );
nor \U$48194 ( \48571 , \48569 , \48570 );
and \U$48195 ( \48572 , \48571 , \10936 );
not \U$48196 ( \48573 , \48571 );
and \U$48197 ( \48574 , \48573 , \11474 );
nor \U$48198 ( \48575 , \48572 , \48574 );
and \U$48199 ( \48576 , \48568 , \48575 );
and \U$48200 ( \48577 , \48560 , \48567 );
or \U$48201 ( \48578 , \48576 , \48577 );
and \U$48202 ( \48579 , \15726 , RIae76910_52);
and \U$48203 ( \48580 , RIae76be0_58, RIae7aab0_192);
nor \U$48204 ( \48581 , \48579 , \48580 );
and \U$48205 ( \48582 , \48581 , \14959 );
not \U$48206 ( \48583 , \48581 );
and \U$48207 ( \48584 , \48583 , RIae7aa38_191);
nor \U$48208 ( \48585 , \48582 , \48584 );
xor \U$48209 ( \48586 , \48585 , \400 );
and \U$48210 ( \48587 , \14964 , RIae76a00_54);
and \U$48211 ( \48588 , RIae76820_50, \14962 );
nor \U$48212 ( \48589 , \48587 , \48588 );
and \U$48213 ( \48590 , \48589 , \14463 );
not \U$48214 ( \48591 , \48589 );
and \U$48215 ( \48592 , \48591 , \14462 );
nor \U$48216 ( \48593 , \48590 , \48592 );
and \U$48217 ( \48594 , \48586 , \48593 );
and \U$48218 ( \48595 , \48585 , \400 );
or \U$48219 ( \48596 , \48594 , \48595 );
xor \U$48220 ( \48597 , \48578 , \48596 );
and \U$48221 ( \48598 , \12180 , RIae76640_46);
and \U$48222 ( \48599 , RIae76190_36, \12178 );
nor \U$48223 ( \48600 , \48598 , \48599 );
and \U$48224 ( \48601 , \48600 , \12184 );
not \U$48225 ( \48602 , \48600 );
and \U$48226 ( \48603 , \48602 , \11827 );
nor \U$48227 ( \48604 , \48601 , \48603 );
and \U$48228 ( \48605 , \13059 , RIae760a0_34);
and \U$48229 ( \48606 , RIae76370_40, \13057 );
nor \U$48230 ( \48607 , \48605 , \48606 );
and \U$48231 ( \48608 , \48607 , \13063 );
not \U$48232 ( \48609 , \48607 );
and \U$48233 ( \48610 , \48609 , \12718 );
nor \U$48234 ( \48611 , \48608 , \48610 );
xor \U$48235 ( \48612 , \48604 , \48611 );
and \U$48236 ( \48613 , \14059 , RIae76280_38);
and \U$48237 ( \48614 , RIae76af0_56, \14057 );
nor \U$48238 ( \48615 , \48613 , \48614 );
and \U$48239 ( \48616 , \48615 , \13502 );
not \U$48240 ( \48617 , \48615 );
and \U$48241 ( \48618 , \48617 , \14063 );
nor \U$48242 ( \48619 , \48616 , \48618 );
and \U$48243 ( \48620 , \48612 , \48619 );
and \U$48244 ( \48621 , \48604 , \48611 );
or \U$48245 ( \48622 , \48620 , \48621 );
and \U$48246 ( \48623 , \48597 , \48622 );
and \U$48247 ( \48624 , \48578 , \48596 );
or \U$48248 ( \48625 , \48623 , \48624 );
xor \U$48249 ( \48626 , \48553 , \48625 );
and \U$48250 ( \48627 , \8371 , RIae75560_10);
and \U$48251 ( \48628 , RIae75830_16, \8369 );
nor \U$48252 ( \48629 , \48627 , \48628 );
and \U$48253 ( \48630 , \48629 , \8020 );
not \U$48254 ( \48631 , \48629 );
and \U$48255 ( \48632 , \48631 , \8019 );
nor \U$48256 ( \48633 , \48630 , \48632 );
and \U$48257 ( \48634 , \7633 , RIae75dd0_28);
and \U$48258 ( \48635 , RIae75650_12, \7631 );
nor \U$48259 ( \48636 , \48634 , \48635 );
and \U$48260 ( \48637 , \48636 , \7206 );
not \U$48261 ( \48638 , \48636 );
and \U$48262 ( \48639 , \48638 , \7205 );
nor \U$48263 ( \48640 , \48637 , \48639 );
xor \U$48264 ( \48641 , \48633 , \48640 );
and \U$48265 ( \48642 , \8966 , RIae75740_14);
and \U$48266 ( \48643 , RIae75290_4, \8964 );
nor \U$48267 ( \48644 , \48642 , \48643 );
and \U$48268 ( \48645 , \48644 , \8799 );
not \U$48269 ( \48646 , \48644 );
and \U$48270 ( \48647 , \48646 , \8789 );
nor \U$48271 ( \48648 , \48645 , \48647 );
and \U$48272 ( \48649 , \48641 , \48648 );
and \U$48273 ( \48650 , \48633 , \48640 );
or \U$48274 ( \48651 , \48649 , \48650 );
and \U$48275 ( \48652 , \5896 , RIae75b00_22);
and \U$48276 ( \48653 , RIae75a10_20, \5894 );
nor \U$48277 ( \48654 , \48652 , \48653 );
and \U$48278 ( \48655 , \48654 , \5590 );
not \U$48279 ( \48656 , \48654 );
and \U$48280 ( \48657 , \48656 , \5589 );
nor \U$48281 ( \48658 , \48655 , \48657 );
and \U$48282 ( \48659 , \6172 , RIae75920_18);
and \U$48283 ( \48660 , RIae75fb0_32, \6170 );
nor \U$48284 ( \48661 , \48659 , \48660 );
and \U$48285 ( \48662 , \48661 , \6176 );
not \U$48286 ( \48663 , \48661 );
and \U$48287 ( \48664 , \48663 , \6175 );
nor \U$48288 ( \48665 , \48662 , \48664 );
xor \U$48289 ( \48666 , \48658 , \48665 );
and \U$48290 ( \48667 , \6941 , RIae75ec0_30);
and \U$48291 ( \48668 , RIae75ce0_26, \6939 );
nor \U$48292 ( \48669 , \48667 , \48668 );
and \U$48293 ( \48670 , \48669 , \6314 );
not \U$48294 ( \48671 , \48669 );
and \U$48295 ( \48672 , \48671 , \6945 );
nor \U$48296 ( \48673 , \48670 , \48672 );
and \U$48297 ( \48674 , \48666 , \48673 );
and \U$48298 ( \48675 , \48658 , \48665 );
or \U$48299 ( \48676 , \48674 , \48675 );
xor \U$48300 ( \48677 , \48651 , \48676 );
and \U$48301 ( \48678 , \5399 , RIae78710_116);
and \U$48302 ( \48679 , RIae75bf0_24, \5397 );
nor \U$48303 ( \48680 , \48678 , \48679 );
and \U$48304 ( \48681 , \48680 , \5016 );
not \U$48305 ( \48682 , \48680 );
and \U$48306 ( \48683 , \48682 , \5403 );
nor \U$48307 ( \48684 , \48681 , \48683 );
and \U$48308 ( \48685 , \4247 , RIae77ea0_98);
and \U$48309 ( \48686 , RIae789e0_122, \4245 );
nor \U$48310 ( \48687 , \48685 , \48686 );
and \U$48311 ( \48688 , \48687 , \3989 );
not \U$48312 ( \48689 , \48687 );
and \U$48313 ( \48690 , \48689 , \4251 );
nor \U$48314 ( \48691 , \48688 , \48690 );
xor \U$48315 ( \48692 , \48684 , \48691 );
and \U$48316 ( \48693 , \4688 , RIae788f0_120);
and \U$48317 ( \48694 , RIae78800_118, \4686 );
nor \U$48318 ( \48695 , \48693 , \48694 );
and \U$48319 ( \48696 , \48695 , \4481 );
not \U$48320 ( \48697 , \48695 );
and \U$48321 ( \48698 , \48697 , \4482 );
nor \U$48322 ( \48699 , \48696 , \48698 );
and \U$48323 ( \48700 , \48692 , \48699 );
and \U$48324 ( \48701 , \48684 , \48691 );
or \U$48325 ( \48702 , \48700 , \48701 );
and \U$48326 ( \48703 , \48677 , \48702 );
and \U$48327 ( \48704 , \48651 , \48676 );
or \U$48328 ( \48705 , \48703 , \48704 );
and \U$48329 ( \48706 , \48626 , \48705 );
and \U$48330 ( \48707 , \48553 , \48625 );
or \U$48331 ( \48708 , \48706 , \48707 );
xor \U$48332 ( \48709 , \48472 , \48708 );
xor \U$48333 ( \48710 , \48297 , \48304 );
xor \U$48334 ( \48711 , \48710 , \48312 );
xor \U$48335 ( \48712 , \48217 , \48224 );
xor \U$48336 ( \48713 , \48712 , \48232 );
and \U$48337 ( \48714 , \48711 , \48713 );
xor \U$48338 ( \48715 , \48268 , \48275 );
xor \U$48339 ( \48716 , \48715 , \48283 );
xor \U$48340 ( \48717 , \48217 , \48224 );
xor \U$48341 ( \48718 , \48717 , \48232 );
and \U$48342 ( \48719 , \48716 , \48718 );
and \U$48343 ( \48720 , \48711 , \48716 );
or \U$48344 ( \48721 , \48714 , \48719 , \48720 );
xor \U$48345 ( \48722 , \48373 , \48375 );
xor \U$48346 ( \48723 , \48722 , \48378 );
and \U$48347 ( \48724 , \48721 , \48723 );
xor \U$48348 ( \48725 , \47717 , \47724 );
xor \U$48349 ( \48726 , \48725 , \47732 );
xor \U$48350 ( \48727 , \48062 , \48067 );
xor \U$48351 ( \48728 , \48726 , \48727 );
xor \U$48352 ( \48729 , \48373 , \48375 );
xor \U$48353 ( \48730 , \48729 , \48378 );
and \U$48354 ( \48731 , \48728 , \48730 );
and \U$48355 ( \48732 , \48721 , \48728 );
or \U$48356 ( \48733 , \48724 , \48731 , \48732 );
and \U$48357 ( \48734 , \48709 , \48733 );
and \U$48358 ( \48735 , \48472 , \48708 );
or \U$48359 ( \48736 , \48734 , \48735 );
xor \U$48360 ( \48737 , \48393 , \48736 );
xor \U$48361 ( \48738 , \47583 , \47608 );
xor \U$48362 ( \48739 , \48738 , \47634 );
xor \U$48363 ( \48740 , \47662 , \47680 );
xor \U$48364 ( \48741 , \48740 , \47706 );
xor \U$48365 ( \48742 , \48739 , \48741 );
xor \U$48366 ( \48743 , \47735 , \47760 );
xor \U$48367 ( \48744 , \48743 , \47786 );
xor \U$48368 ( \48745 , \48742 , \48744 );
xor \U$48369 ( \48746 , \47590 , \47597 );
xor \U$48370 ( \48747 , \48746 , \47605 );
xor \U$48371 ( \48748 , \48117 , \48122 );
xor \U$48372 ( \48749 , \48747 , \48748 );
xor \U$48373 ( \48750 , \48153 , \48179 );
xor \U$48374 ( \48751 , \48750 , \48207 );
xor \U$48375 ( \48752 , \48749 , \48751 );
xor \U$48376 ( \48753 , \48078 , \48104 );
xor \U$48377 ( \48754 , \48753 , \48111 );
and \U$48378 ( \48755 , \48752 , \48754 );
and \U$48379 ( \48756 , \48749 , \48751 );
or \U$48380 ( \48757 , \48755 , \48756 );
xor \U$48381 ( \48758 , \48745 , \48757 );
xor \U$48382 ( \48759 , \47935 , \47943 );
xor \U$48383 ( \48760 , \48759 , \47950 );
not \U$48384 ( \48761 , \47893 );
xor \U$48385 ( \48762 , \47884 , \47924 );
not \U$48386 ( \48763 , \48762 );
or \U$48387 ( \48764 , \48761 , \48763 );
or \U$48388 ( \48765 , \48762 , \47893 );
nand \U$48389 ( \48766 , \48764 , \48765 );
xor \U$48390 ( \48767 , \48760 , \48766 );
xor \U$48391 ( \48768 , \47843 , \47845 );
xor \U$48392 ( \48769 , \48768 , \47852 );
xor \U$48393 ( \48770 , \48767 , \48769 );
and \U$48394 ( \48771 , \48758 , \48770 );
and \U$48395 ( \48772 , \48745 , \48757 );
or \U$48396 ( \48773 , \48771 , \48772 );
and \U$48397 ( \48774 , \48737 , \48773 );
and \U$48398 ( \48775 , \48393 , \48736 );
or \U$48399 ( \48776 , \48774 , \48775 );
and \U$48400 ( \48777 , \48060 , \48776 );
and \U$48401 ( \48778 , \48053 , \48059 );
or \U$48402 ( \48779 , \48777 , \48778 );
not \U$48403 ( \48780 , \48779 );
not \U$48404 ( \48781 , \48041 );
not \U$48405 ( \48782 , \48036 );
and \U$48406 ( \48783 , \48781 , \48782 );
and \U$48407 ( \48784 , \48041 , \48036 );
nor \U$48408 ( \48785 , \48784 , \48045 );
nor \U$48409 ( \48786 , \48783 , \48785 );
xor \U$48410 ( \48787 , \48739 , \48741 );
and \U$48411 ( \48788 , \48787 , \48744 );
and \U$48412 ( \48789 , \48739 , \48741 );
nor \U$48413 ( \48790 , \48788 , \48789 );
not \U$48414 ( \48791 , \48790 );
xor \U$48415 ( \48792 , \47224 , \47249 );
xor \U$48416 ( \48793 , \48792 , \47277 );
not \U$48417 ( \48794 , \48793 );
and \U$48418 ( \48795 , \48791 , \48794 );
and \U$48419 ( \48796 , \48790 , \48793 );
xor \U$48420 ( \48797 , \48760 , \48766 );
and \U$48421 ( \48798 , \48797 , \48769 );
and \U$48422 ( \48799 , \48760 , \48766 );
nor \U$48423 ( \48800 , \48798 , \48799 );
nor \U$48424 ( \48801 , \48796 , \48800 );
nor \U$48425 ( \48802 , \48795 , \48801 );
or \U$48426 ( \48803 , \48786 , \48802 );
not \U$48427 ( \48804 , \48802 );
not \U$48428 ( \48805 , \48786 );
or \U$48429 ( \48806 , \48804 , \48805 );
xor \U$48430 ( \48807 , \48072 , \48114 );
and \U$48431 ( \48808 , \48807 , \48127 );
and \U$48432 ( \48809 , \48072 , \48114 );
or \U$48433 ( \48810 , \48808 , \48809 );
xor \U$48434 ( \48811 , \48210 , \48289 );
and \U$48435 ( \48812 , \48811 , \48369 );
and \U$48436 ( \48813 , \48210 , \48289 );
or \U$48437 ( \48814 , \48812 , \48813 );
xor \U$48438 ( \48815 , \48810 , \48814 );
xor \U$48439 ( \48816 , \48381 , \48386 );
and \U$48440 ( \48817 , \48816 , \48389 );
and \U$48441 ( \48818 , \48381 , \48386 );
or \U$48442 ( \48819 , \48817 , \48818 );
and \U$48443 ( \48820 , \48815 , \48819 );
and \U$48444 ( \48821 , \48810 , \48814 );
or \U$48445 ( \48822 , \48820 , \48821 );
nand \U$48446 ( \48823 , \48806 , \48822 );
nand \U$48447 ( \48824 , \48803 , \48823 );
not \U$48448 ( \48825 , \48824 );
xor \U$48449 ( \48826 , \47197 , \47280 );
xor \U$48450 ( \48827 , \48826 , \47364 );
xor \U$48451 ( \48828 , \47972 , \47984 );
xor \U$48452 ( \48829 , \48828 , \47987 );
and \U$48453 ( \48830 , \48827 , \48829 );
xor \U$48454 ( \48831 , \48001 , \48003 );
xor \U$48455 ( \48832 , \48831 , \48006 );
xor \U$48456 ( \48833 , \47972 , \47984 );
xor \U$48457 ( \48834 , \48833 , \47987 );
and \U$48458 ( \48835 , \48832 , \48834 );
and \U$48459 ( \48836 , \48827 , \48832 );
or \U$48460 ( \48837 , \48830 , \48835 , \48836 );
not \U$48461 ( \48838 , \48837 );
or \U$48462 ( \48839 , \48825 , \48838 );
or \U$48463 ( \48840 , \48837 , \48824 );
nand \U$48464 ( \48841 , \48839 , \48840 );
not \U$48465 ( \48842 , \48841 );
not \U$48466 ( \48843 , \47107 );
not \U$48467 ( \48844 , \47079 );
or \U$48468 ( \48845 , \48843 , \48844 );
or \U$48469 ( \48846 , \47079 , \47107 );
nand \U$48470 ( \48847 , \48845 , \48846 );
not \U$48471 ( \48848 , \48847 );
not \U$48472 ( \48849 , \47089 );
and \U$48473 ( \48850 , \48848 , \48849 );
and \U$48474 ( \48851 , \48847 , \47089 );
nor \U$48475 ( \48852 , \48850 , \48851 );
not \U$48476 ( \48853 , \48852 );
and \U$48477 ( \48854 , \48842 , \48853 );
and \U$48478 ( \48855 , \48841 , \48852 );
nor \U$48479 ( \48856 , \48854 , \48855 );
not \U$48480 ( \48857 , \48856 );
or \U$48481 ( \48858 , \48780 , \48857 );
or \U$48482 ( \48859 , \48856 , \48779 );
nand \U$48483 ( \48860 , \48858 , \48859 );
not \U$48484 ( \48861 , \48860 );
xor \U$48485 ( \48862 , \47367 , \47436 );
xor \U$48486 ( \48863 , \48862 , \47466 );
xor \U$48487 ( \48864 , \47958 , \47990 );
xor \U$48488 ( \48865 , \48864 , \48009 );
xnor \U$48489 ( \48866 , \48863 , \48865 );
not \U$48490 ( \48867 , \48866 );
xor \U$48491 ( \48868 , \46894 , \46952 );
xor \U$48492 ( \48869 , \48868 , \46979 );
xor \U$48493 ( \48870 , \47541 , \47548 );
xor \U$48494 ( \48871 , \48869 , \48870 );
not \U$48495 ( \48872 , \48871 );
and \U$48496 ( \48873 , \48867 , \48872 );
and \U$48497 ( \48874 , \48866 , \48871 );
nor \U$48498 ( \48875 , \48873 , \48874 );
not \U$48499 ( \48876 , \48875 );
and \U$48500 ( \48877 , \48861 , \48876 );
and \U$48501 ( \48878 , \48860 , \48875 );
nor \U$48502 ( \48879 , \48877 , \48878 );
not \U$48503 ( \48880 , \48879 );
not \U$48504 ( \48881 , \48822 );
not \U$48505 ( \48882 , \48802 );
or \U$48506 ( \48883 , \48881 , \48882 );
or \U$48507 ( \48884 , \48802 , \48822 );
nand \U$48508 ( \48885 , \48883 , \48884 );
not \U$48509 ( \48886 , \48885 );
not \U$48510 ( \48887 , \48786 );
and \U$48511 ( \48888 , \48886 , \48887 );
and \U$48512 ( \48889 , \48885 , \48786 );
nor \U$48513 ( \48890 , \48888 , \48889 );
not \U$48514 ( \48891 , \48890 );
xor \U$48515 ( \48892 , \48053 , \48059 );
xor \U$48516 ( \48893 , \48892 , \48776 );
nand \U$48517 ( \48894 , \48891 , \48893 );
xor \U$48518 ( \48895 , \48472 , \48708 );
xor \U$48519 ( \48896 , \48895 , \48733 );
xor \U$48520 ( \48897 , \48128 , \48370 );
xor \U$48521 ( \48898 , \48897 , \48390 );
and \U$48522 ( \48899 , \48896 , \48898 );
xor \U$48523 ( \48900 , \48745 , \48757 );
xor \U$48524 ( \48901 , \48900 , \48770 );
xor \U$48525 ( \48902 , \48128 , \48370 );
xor \U$48526 ( \48903 , \48902 , \48390 );
and \U$48527 ( \48904 , \48901 , \48903 );
and \U$48528 ( \48905 , \48896 , \48901 );
or \U$48529 ( \48906 , \48899 , \48904 , \48905 );
not \U$48530 ( \48907 , \48793 );
xor \U$48531 ( \48908 , \48790 , \48800 );
not \U$48532 ( \48909 , \48908 );
or \U$48533 ( \48910 , \48907 , \48909 );
or \U$48534 ( \48911 , \48908 , \48793 );
nand \U$48535 ( \48912 , \48910 , \48911 );
and \U$48536 ( \48913 , \48906 , \48912 );
not \U$48537 ( \48914 , \48906 );
not \U$48538 ( \48915 , \48912 );
and \U$48539 ( \48916 , \48914 , \48915 );
xor \U$48540 ( \48917 , \48235 , \48260 );
xor \U$48541 ( \48918 , \48917 , \48286 );
xor \U$48542 ( \48919 , \48749 , \48751 );
xor \U$48543 ( \48920 , \48919 , \48754 );
and \U$48544 ( \48921 , \48918 , \48920 );
xor \U$48545 ( \48922 , \48373 , \48375 );
xor \U$48546 ( \48923 , \48922 , \48378 );
xor \U$48547 ( \48924 , \48721 , \48728 );
xor \U$48548 ( \48925 , \48923 , \48924 );
xor \U$48549 ( \48926 , \48749 , \48751 );
xor \U$48550 ( \48927 , \48926 , \48754 );
and \U$48551 ( \48928 , \48925 , \48927 );
and \U$48552 ( \48929 , \48918 , \48925 );
or \U$48553 ( \48930 , \48921 , \48928 , \48929 );
xor \U$48554 ( \48931 , \48506 , \48513 );
xor \U$48555 ( \48932 , \48931 , \48521 );
xor \U$48556 ( \48933 , \48532 , \48539 );
xor \U$48557 ( \48934 , \48933 , \48547 );
xor \U$48558 ( \48935 , \48932 , \48934 );
xor \U$48559 ( \48936 , \48480 , \48488 );
xor \U$48560 ( \48937 , \48936 , \48496 );
and \U$48561 ( \48938 , \48935 , \48937 );
and \U$48562 ( \48939 , \48932 , \48934 );
or \U$48563 ( \48940 , \48938 , \48939 );
and \U$48564 ( \48941 , \672 , RIae77ae0_90);
and \U$48565 ( \48942 , RIae779f0_88, \670 );
nor \U$48566 ( \48943 , \48941 , \48942 );
and \U$48567 ( \48944 , \48943 , \588 );
not \U$48568 ( \48945 , \48943 );
and \U$48569 ( \48946 , \48945 , \587 );
nor \U$48570 ( \48947 , \48944 , \48946 );
not \U$48571 ( \48948 , \469 );
and \U$48572 ( \48949 , \514 , RIae77630_80);
and \U$48573 ( \48950 , RIae77540_78, \512 );
nor \U$48574 ( \48951 , \48949 , \48950 );
not \U$48575 ( \48952 , \48951 );
or \U$48576 ( \48953 , \48948 , \48952 );
or \U$48577 ( \48954 , \48951 , \469 );
nand \U$48578 ( \48955 , \48953 , \48954 );
xor \U$48579 ( \48956 , \48947 , \48955 );
and \U$48580 ( \48957 , \558 , RIae776a8_81);
and \U$48581 ( \48958 , RIae77450_76, \556 );
nor \U$48582 ( \48959 , \48957 , \48958 );
and \U$48583 ( \48960 , \48959 , \504 );
not \U$48584 ( \48961 , \48959 );
and \U$48585 ( \48962 , \48961 , \562 );
nor \U$48586 ( \48963 , \48960 , \48962 );
and \U$48587 ( \48964 , \48956 , \48963 );
and \U$48588 ( \48965 , \48947 , \48955 );
or \U$48589 ( \48966 , \48964 , \48965 );
xor \U$48590 ( \48967 , \48409 , \48417 );
xor \U$48591 ( \48968 , \48966 , \48967 );
xor \U$48592 ( \48969 , \48435 , \48442 );
xor \U$48593 ( \48970 , \48969 , \48450 );
and \U$48594 ( \48971 , \48968 , \48970 );
and \U$48595 ( \48972 , \48966 , \48967 );
or \U$48596 ( \48973 , \48971 , \48972 );
xor \U$48597 ( \48974 , \48940 , \48973 );
xor \U$48598 ( \48975 , \48658 , \48665 );
xor \U$48599 ( \48976 , \48975 , \48673 );
xor \U$48600 ( \48977 , \48684 , \48691 );
xor \U$48601 ( \48978 , \48977 , \48699 );
and \U$48602 ( \48979 , \48976 , \48978 );
xor \U$48603 ( \48980 , \48633 , \48640 );
xor \U$48604 ( \48981 , \48980 , \48648 );
xor \U$48605 ( \48982 , \48684 , \48691 );
xor \U$48606 ( \48983 , \48982 , \48699 );
and \U$48607 ( \48984 , \48981 , \48983 );
and \U$48608 ( \48985 , \48976 , \48981 );
or \U$48609 ( \48986 , \48979 , \48984 , \48985 );
and \U$48610 ( \48987 , \48974 , \48986 );
and \U$48611 ( \48988 , \48940 , \48973 );
or \U$48612 ( \48989 , \48987 , \48988 );
and \U$48613 ( \48990 , \6941 , RIae75fb0_32);
and \U$48614 ( \48991 , RIae75ec0_30, \6939 );
nor \U$48615 ( \48992 , \48990 , \48991 );
and \U$48616 ( \48993 , \48992 , \6314 );
not \U$48617 ( \48994 , \48992 );
and \U$48618 ( \48995 , \48994 , \6945 );
nor \U$48619 ( \48996 , \48993 , \48995 );
and \U$48620 ( \48997 , \7633 , RIae75ce0_26);
and \U$48621 ( \48998 , RIae75dd0_28, \7631 );
nor \U$48622 ( \48999 , \48997 , \48998 );
and \U$48623 ( \49000 , \48999 , \7206 );
not \U$48624 ( \49001 , \48999 );
and \U$48625 ( \49002 , \49001 , \7205 );
nor \U$48626 ( \49003 , \49000 , \49002 );
xor \U$48627 ( \49004 , \48996 , \49003 );
and \U$48628 ( \49005 , \8371 , RIae75650_12);
and \U$48629 ( \49006 , RIae75560_10, \8369 );
nor \U$48630 ( \49007 , \49005 , \49006 );
and \U$48631 ( \49008 , \49007 , \8020 );
not \U$48632 ( \49009 , \49007 );
and \U$48633 ( \49010 , \49009 , \8019 );
nor \U$48634 ( \49011 , \49008 , \49010 );
and \U$48635 ( \49012 , \49004 , \49011 );
and \U$48636 ( \49013 , \48996 , \49003 );
or \U$48637 ( \49014 , \49012 , \49013 );
and \U$48638 ( \49015 , \4688 , RIae789e0_122);
and \U$48639 ( \49016 , RIae788f0_120, \4686 );
nor \U$48640 ( \49017 , \49015 , \49016 );
and \U$48641 ( \49018 , \49017 , \4481 );
not \U$48642 ( \49019 , \49017 );
and \U$48643 ( \49020 , \49019 , \4482 );
nor \U$48644 ( \49021 , \49018 , \49020 );
and \U$48645 ( \49022 , \3730 , RIae77cc0_94);
and \U$48646 ( \49023 , RIae77bd0_92, \3728 );
nor \U$48647 ( \49024 , \49022 , \49023 );
and \U$48648 ( \49025 , \49024 , \3732 );
not \U$48649 ( \49026 , \49024 );
and \U$48650 ( \49027 , \49026 , \3422 );
nor \U$48651 ( \49028 , \49025 , \49027 );
xor \U$48652 ( \49029 , \49021 , \49028 );
and \U$48653 ( \49030 , \4247 , RIae77db0_96);
and \U$48654 ( \49031 , RIae77ea0_98, \4245 );
nor \U$48655 ( \49032 , \49030 , \49031 );
and \U$48656 ( \49033 , \49032 , \3989 );
not \U$48657 ( \49034 , \49032 );
and \U$48658 ( \49035 , \49034 , \4251 );
nor \U$48659 ( \49036 , \49033 , \49035 );
and \U$48660 ( \49037 , \49029 , \49036 );
and \U$48661 ( \49038 , \49021 , \49028 );
or \U$48662 ( \49039 , \49037 , \49038 );
xor \U$48663 ( \49040 , \49014 , \49039 );
and \U$48664 ( \49041 , \5399 , RIae78800_118);
and \U$48665 ( \49042 , RIae78710_116, \5397 );
nor \U$48666 ( \49043 , \49041 , \49042 );
and \U$48667 ( \49044 , \49043 , \5016 );
not \U$48668 ( \49045 , \49043 );
and \U$48669 ( \49046 , \49045 , \5403 );
nor \U$48670 ( \49047 , \49044 , \49046 );
and \U$48671 ( \49048 , \5896 , RIae75bf0_24);
and \U$48672 ( \49049 , RIae75b00_22, \5894 );
nor \U$48673 ( \49050 , \49048 , \49049 );
and \U$48674 ( \49051 , \49050 , \5590 );
not \U$48675 ( \49052 , \49050 );
and \U$48676 ( \49053 , \49052 , \5589 );
nor \U$48677 ( \49054 , \49051 , \49053 );
xor \U$48678 ( \49055 , \49047 , \49054 );
and \U$48679 ( \49056 , \6172 , RIae75a10_20);
and \U$48680 ( \49057 , RIae75920_18, \6170 );
nor \U$48681 ( \49058 , \49056 , \49057 );
and \U$48682 ( \49059 , \49058 , \6176 );
not \U$48683 ( \49060 , \49058 );
and \U$48684 ( \49061 , \49060 , \6175 );
nor \U$48685 ( \49062 , \49059 , \49061 );
and \U$48686 ( \49063 , \49055 , \49062 );
and \U$48687 ( \49064 , \49047 , \49054 );
or \U$48688 ( \49065 , \49063 , \49064 );
and \U$48689 ( \49066 , \49040 , \49065 );
and \U$48690 ( \49067 , \49014 , \49039 );
or \U$48691 ( \49068 , \49066 , \49067 );
and \U$48692 ( \49069 , \10548 , RIae75380_6);
and \U$48693 ( \49070 , RIae75470_8, \10546 );
nor \U$48694 ( \49071 , \49069 , \49070 );
and \U$48695 ( \49072 , \49071 , \10421 );
not \U$48696 ( \49073 , \49071 );
and \U$48697 ( \49074 , \49073 , \10118 );
nor \U$48698 ( \49075 , \49072 , \49074 );
and \U$48699 ( \49076 , \8966 , RIae75830_16);
and \U$48700 ( \49077 , RIae75740_14, \8964 );
nor \U$48701 ( \49078 , \49076 , \49077 );
and \U$48702 ( \49079 , \49078 , \8799 );
not \U$48703 ( \49080 , \49078 );
and \U$48704 ( \49081 , \49080 , \8789 );
nor \U$48705 ( \49082 , \49079 , \49081 );
xor \U$48706 ( \49083 , \49075 , \49082 );
and \U$48707 ( \49084 , \9760 , RIae75290_4);
and \U$48708 ( \49085 , RIae751a0_2, \9758 );
nor \U$48709 ( \49086 , \49084 , \49085 );
and \U$48710 ( \49087 , \49086 , \9273 );
not \U$48711 ( \49088 , \49086 );
and \U$48712 ( \49089 , \49088 , \9272 );
nor \U$48713 ( \49090 , \49087 , \49089 );
and \U$48714 ( \49091 , \49083 , \49090 );
and \U$48715 ( \49092 , \49075 , \49082 );
or \U$48716 ( \49093 , \49091 , \49092 );
and \U$48717 ( \49094 , \14964 , RIae76af0_56);
and \U$48718 ( \49095 , RIae76a00_54, \14962 );
nor \U$48719 ( \49096 , \49094 , \49095 );
and \U$48720 ( \49097 , \49096 , \14463 );
not \U$48721 ( \49098 , \49096 );
and \U$48722 ( \49099 , \49098 , \14462 );
nor \U$48723 ( \49100 , \49097 , \49099 );
and \U$48724 ( \49101 , \15726 , RIae76820_50);
and \U$48725 ( \49102 , RIae76910_52, RIae7aab0_192);
nor \U$48726 ( \49103 , \49101 , \49102 );
and \U$48727 ( \49104 , \49103 , \14959 );
not \U$48728 ( \49105 , \49103 );
and \U$48729 ( \49106 , \49105 , RIae7aa38_191);
nor \U$48730 ( \49107 , \49104 , \49106 );
xor \U$48731 ( \49108 , \49100 , \49107 );
and \U$48732 ( \49109 , \14059 , RIae76370_40);
and \U$48733 ( \49110 , RIae76280_38, \14057 );
nor \U$48734 ( \49111 , \49109 , \49110 );
and \U$48735 ( \49112 , \49111 , \13502 );
not \U$48736 ( \49113 , \49111 );
and \U$48737 ( \49114 , \49113 , \14063 );
nor \U$48738 ( \49115 , \49112 , \49114 );
and \U$48739 ( \49116 , \49108 , \49115 );
and \U$48740 ( \49117 , \49100 , \49107 );
or \U$48741 ( \49118 , \49116 , \49117 );
xor \U$48742 ( \49119 , \49093 , \49118 );
and \U$48743 ( \49120 , \12180 , RIae76730_48);
and \U$48744 ( \49121 , RIae76640_46, \12178 );
nor \U$48745 ( \49122 , \49120 , \49121 );
and \U$48746 ( \49123 , \49122 , \12184 );
not \U$48747 ( \49124 , \49122 );
and \U$48748 ( \49125 , \49124 , \11827 );
nor \U$48749 ( \49126 , \49123 , \49125 );
and \U$48750 ( \49127 , \11470 , RIae76460_42);
and \U$48751 ( \49128 , RIae76550_44, \11468 );
nor \U$48752 ( \49129 , \49127 , \49128 );
and \U$48753 ( \49130 , \49129 , \10936 );
not \U$48754 ( \49131 , \49129 );
and \U$48755 ( \49132 , \49131 , \11474 );
nor \U$48756 ( \49133 , \49130 , \49132 );
xor \U$48757 ( \49134 , \49126 , \49133 );
and \U$48758 ( \49135 , \13059 , RIae76190_36);
and \U$48759 ( \49136 , RIae760a0_34, \13057 );
nor \U$48760 ( \49137 , \49135 , \49136 );
and \U$48761 ( \49138 , \49137 , \13063 );
not \U$48762 ( \49139 , \49137 );
and \U$48763 ( \49140 , \49139 , \12718 );
nor \U$48764 ( \49141 , \49138 , \49140 );
and \U$48765 ( \49142 , \49134 , \49141 );
and \U$48766 ( \49143 , \49126 , \49133 );
or \U$48767 ( \49144 , \49142 , \49143 );
and \U$48768 ( \49145 , \49119 , \49144 );
and \U$48769 ( \49146 , \49093 , \49118 );
or \U$48770 ( \49147 , \49145 , \49146 );
xor \U$48771 ( \49148 , \49068 , \49147 );
and \U$48772 ( \49149 , \1939 , RIae77270_72);
and \U$48773 ( \49150 , RIae77360_74, \1937 );
nor \U$48774 ( \49151 , \49149 , \49150 );
and \U$48775 ( \49152 , \49151 , \1735 );
not \U$48776 ( \49153 , \49151 );
and \U$48777 ( \49154 , \49153 , \1734 );
nor \U$48778 ( \49155 , \49152 , \49154 );
and \U$48779 ( \49156 , \1593 , RIae77108_69);
and \U$48780 ( \49157 , RIae77090_68, \1591 );
nor \U$48781 ( \49158 , \49156 , \49157 );
and \U$48782 ( \49159 , \49158 , \1498 );
not \U$48783 ( \49160 , \49158 );
and \U$48784 ( \49161 , \49160 , \1488 );
nor \U$48785 ( \49162 , \49159 , \49161 );
xor \U$48786 ( \49163 , \49155 , \49162 );
and \U$48787 ( \49164 , \2224 , RIae78350_108);
and \U$48788 ( \49165 , RIae78170_104, \2222 );
nor \U$48789 ( \49166 , \49164 , \49165 );
and \U$48790 ( \49167 , \49166 , \2061 );
not \U$48791 ( \49168 , \49166 );
and \U$48792 ( \49169 , \49168 , \2060 );
nor \U$48793 ( \49170 , \49167 , \49169 );
and \U$48794 ( \49171 , \49163 , \49170 );
and \U$48795 ( \49172 , \49155 , \49162 );
or \U$48796 ( \49173 , \49171 , \49172 );
not \U$48797 ( \49174 , \789 );
and \U$48798 ( \49175 , \883 , RIae77810_84);
and \U$48799 ( \49176 , RIae77900_86, \881 );
nor \U$48800 ( \49177 , \49175 , \49176 );
not \U$48801 ( \49178 , \49177 );
or \U$48802 ( \49179 , \49174 , \49178 );
or \U$48803 ( \49180 , \49177 , \789 );
nand \U$48804 ( \49181 , \49179 , \49180 );
and \U$48805 ( \49182 , \1138 , RIae76fa0_66);
and \U$48806 ( \49183 , RIae76eb0_64, \1136 );
nor \U$48807 ( \49184 , \49182 , \49183 );
and \U$48808 ( \49185 , \49184 , \1012 );
not \U$48809 ( \49186 , \49184 );
and \U$48810 ( \49187 , \49186 , \1142 );
nor \U$48811 ( \49188 , \49185 , \49187 );
xor \U$48812 ( \49189 , \49181 , \49188 );
and \U$48813 ( \49190 , \1376 , RIae76dc0_62);
and \U$48814 ( \49191 , RIae76cd0_60, \1374 );
nor \U$48815 ( \49192 , \49190 , \49191 );
and \U$48816 ( \49193 , \49192 , \1380 );
not \U$48817 ( \49194 , \49192 );
and \U$48818 ( \49195 , \49194 , \1261 );
nor \U$48819 ( \49196 , \49193 , \49195 );
and \U$48820 ( \49197 , \49189 , \49196 );
and \U$48821 ( \49198 , \49181 , \49188 );
or \U$48822 ( \49199 , \49197 , \49198 );
xor \U$48823 ( \49200 , \49173 , \49199 );
not \U$48824 ( \49201 , \3218 );
and \U$48825 ( \49202 , \3214 , RIae78440_110);
and \U$48826 ( \49203 , RIae784b8_111, \3212 );
nor \U$48827 ( \49204 , \49202 , \49203 );
not \U$48828 ( \49205 , \49204 );
or \U$48829 ( \49206 , \49201 , \49205 );
or \U$48830 ( \49207 , \49204 , \2774 );
nand \U$48831 ( \49208 , \49206 , \49207 );
and \U$48832 ( \49209 , \2607 , RIae77f90_100);
and \U$48833 ( \49210 , RIae78080_102, \2605 );
nor \U$48834 ( \49211 , \49209 , \49210 );
and \U$48835 ( \49212 , \49211 , \2611 );
not \U$48836 ( \49213 , \49211 );
and \U$48837 ( \49214 , \49213 , \2397 );
nor \U$48838 ( \49215 , \49212 , \49214 );
xor \U$48839 ( \49216 , \49208 , \49215 );
not \U$48840 ( \49217 , \2789 );
and \U$48841 ( \49218 , \2783 , RIae78260_106);
and \U$48842 ( \49219 , RIae78620_114, \2781 );
nor \U$48843 ( \49220 , \49218 , \49219 );
not \U$48844 ( \49221 , \49220 );
or \U$48845 ( \49222 , \49217 , \49221 );
or \U$48846 ( \49223 , \49220 , \2789 );
nand \U$48847 ( \49224 , \49222 , \49223 );
and \U$48848 ( \49225 , \49216 , \49224 );
and \U$48849 ( \49226 , \49208 , \49215 );
or \U$48850 ( \49227 , \49225 , \49226 );
and \U$48851 ( \49228 , \49200 , \49227 );
and \U$48852 ( \49229 , \49173 , \49199 );
or \U$48853 ( \49230 , \49228 , \49229 );
and \U$48854 ( \49231 , \49148 , \49230 );
and \U$48855 ( \49232 , \49068 , \49147 );
or \U$48856 ( \49233 , \49231 , \49232 );
xor \U$48857 ( \49234 , \48989 , \49233 );
xor \U$48858 ( \49235 , \48560 , \48567 );
xor \U$48859 ( \49236 , \49235 , \48575 );
xor \U$48860 ( \49237 , \48585 , \400 );
xor \U$48861 ( \49238 , \49237 , \48593 );
and \U$48862 ( \49239 , \49236 , \49238 );
xor \U$48863 ( \49240 , \48604 , \48611 );
xor \U$48864 ( \49241 , \49240 , \48619 );
xor \U$48865 ( \49242 , \48585 , \400 );
xor \U$48866 ( \49243 , \49242 , \48593 );
and \U$48867 ( \49244 , \49241 , \49243 );
and \U$48868 ( \49245 , \49236 , \49241 );
or \U$48869 ( \49246 , \49239 , \49244 , \49245 );
xor \U$48870 ( \49247 , \48242 , \48249 );
xor \U$48871 ( \49248 , \49247 , \48257 );
xor \U$48872 ( \49249 , \49246 , \49248 );
xor \U$48873 ( \49250 , \48217 , \48224 );
xor \U$48874 ( \49251 , \49250 , \48232 );
xor \U$48875 ( \49252 , \48711 , \48716 );
xor \U$48876 ( \49253 , \49251 , \49252 );
and \U$48877 ( \49254 , \49249 , \49253 );
and \U$48878 ( \49255 , \49246 , \49248 );
or \U$48879 ( \49256 , \49254 , \49255 );
and \U$48880 ( \49257 , \49234 , \49256 );
and \U$48881 ( \49258 , \48989 , \49233 );
or \U$48882 ( \49259 , \49257 , \49258 );
xor \U$48883 ( \49260 , \48930 , \49259 );
xor \U$48884 ( \49261 , \48499 , \48524 );
xor \U$48885 ( \49262 , \49261 , \48550 );
xor \U$48886 ( \49263 , \48578 , \48596 );
xor \U$48887 ( \49264 , \49263 , \48622 );
and \U$48888 ( \49265 , \49262 , \49264 );
xor \U$48889 ( \49266 , \48651 , \48676 );
xor \U$48890 ( \49267 , \49266 , \48702 );
xor \U$48891 ( \49268 , \48578 , \48596 );
xor \U$48892 ( \49269 , \49268 , \48622 );
and \U$48893 ( \49270 , \49267 , \49269 );
and \U$48894 ( \49271 , \49262 , \49267 );
or \U$48895 ( \49272 , \49265 , \49270 , \49271 );
xor \U$48896 ( \49273 , \48315 , \48340 );
xor \U$48897 ( \49274 , \49273 , \48366 );
xor \U$48898 ( \49275 , \49272 , \49274 );
xor \U$48899 ( \49276 , \48418 , \48426 );
xor \U$48900 ( \49277 , \49276 , \48453 );
xor \U$48901 ( \49278 , \48395 , \48397 );
xor \U$48902 ( \49279 , \49278 , \48400 );
and \U$48903 ( \49280 , \49277 , \49279 );
xor \U$48904 ( \49281 , \48322 , \48329 );
xor \U$48905 ( \49282 , \49281 , \48337 );
xor \U$48906 ( \49283 , \48459 , \48464 );
xor \U$48907 ( \49284 , \49282 , \49283 );
xor \U$48908 ( \49285 , \48395 , \48397 );
xor \U$48909 ( \49286 , \49285 , \48400 );
and \U$48910 ( \49287 , \49284 , \49286 );
and \U$48911 ( \49288 , \49277 , \49284 );
or \U$48912 ( \49289 , \49280 , \49287 , \49288 );
and \U$48913 ( \49290 , \49275 , \49289 );
and \U$48914 ( \49291 , \49272 , \49274 );
or \U$48915 ( \49292 , \49290 , \49291 );
and \U$48916 ( \49293 , \49260 , \49292 );
and \U$48917 ( \49294 , \48930 , \49259 );
nor \U$48918 ( \49295 , \49293 , \49294 );
nor \U$48919 ( \49296 , \48916 , \49295 );
nor \U$48920 ( \49297 , \48913 , \49296 );
not \U$48921 ( \49298 , \49297 );
xor \U$48922 ( \49299 , \47972 , \47984 );
xor \U$48923 ( \49300 , \49299 , \47987 );
xor \U$48924 ( \49301 , \48827 , \48832 );
xor \U$48925 ( \49302 , \49300 , \49301 );
not \U$48926 ( \49303 , \49302 );
and \U$48927 ( \49304 , \49298 , \49303 );
and \U$48928 ( \49305 , \49297 , \49302 );
xor \U$48929 ( \49306 , \48031 , \48033 );
xor \U$48930 ( \49307 , \49306 , \48050 );
xor \U$48931 ( \49308 , \48393 , \48736 );
xor \U$48932 ( \49309 , \49308 , \48773 );
xor \U$48933 ( \49310 , \49307 , \49309 );
xor \U$48934 ( \49311 , \48810 , \48814 );
xor \U$48935 ( \49312 , \49311 , \48819 );
and \U$48936 ( \49313 , \49310 , \49312 );
and \U$48937 ( \49314 , \49307 , \49309 );
nor \U$48938 ( \49315 , \49313 , \49314 );
nor \U$48939 ( \49316 , \49305 , \49315 );
nor \U$48940 ( \49317 , \49304 , \49316 );
xor \U$48941 ( \49318 , \48894 , \49317 );
not \U$48942 ( \49319 , \49318 );
or \U$48943 ( \49320 , \48880 , \49319 );
or \U$48944 ( \49321 , \49318 , \48879 );
nand \U$48945 ( \49322 , \49320 , \49321 );
xor \U$48946 ( \49323 , \49307 , \49309 );
xor \U$48947 ( \49324 , \49323 , \49312 );
xor \U$48948 ( \49325 , \49208 , \49215 );
xor \U$48949 ( \49326 , \49325 , \49224 );
xor \U$48950 ( \49327 , \49155 , \49162 );
xor \U$48951 ( \49328 , \49327 , \49170 );
and \U$48952 ( \49329 , \49326 , \49328 );
xor \U$48953 ( \49330 , \49021 , \49028 );
xor \U$48954 ( \49331 , \49330 , \49036 );
xor \U$48955 ( \49332 , \49155 , \49162 );
xor \U$48956 ( \49333 , \49332 , \49170 );
and \U$48957 ( \49334 , \49331 , \49333 );
and \U$48958 ( \49335 , \49326 , \49331 );
or \U$48959 ( \49336 , \49329 , \49334 , \49335 );
xor \U$48960 ( \49337 , \48947 , \48955 );
xor \U$48961 ( \49338 , \49337 , \48963 );
and \U$48962 ( \49339 , \672 , RIae77450_76);
and \U$48963 ( \49340 , RIae77ae0_90, \670 );
nor \U$48964 ( \49341 , \49339 , \49340 );
and \U$48965 ( \49342 , \49341 , \588 );
not \U$48966 ( \49343 , \49341 );
and \U$48967 ( \49344 , \49343 , \587 );
nor \U$48968 ( \49345 , \49342 , \49344 );
and \U$48969 ( \49346 , \558 , RIae77540_78);
and \U$48970 ( \49347 , RIae776a8_81, \556 );
nor \U$48971 ( \49348 , \49346 , \49347 );
and \U$48972 ( \49349 , \49348 , \504 );
not \U$48973 ( \49350 , \49348 );
and \U$48974 ( \49351 , \49350 , \562 );
nor \U$48975 ( \49352 , \49349 , \49351 );
xor \U$48976 ( \49353 , \49345 , \49352 );
not \U$48977 ( \49354 , \789 );
and \U$48978 ( \49355 , \883 , RIae779f0_88);
and \U$48979 ( \49356 , RIae77810_84, \881 );
nor \U$48980 ( \49357 , \49355 , \49356 );
not \U$48981 ( \49358 , \49357 );
or \U$48982 ( \49359 , \49354 , \49358 );
or \U$48983 ( \49360 , \49357 , \789 );
nand \U$48984 ( \49361 , \49359 , \49360 );
and \U$48985 ( \49362 , \49353 , \49361 );
and \U$48986 ( \49363 , \49345 , \49352 );
or \U$48987 ( \49364 , \49362 , \49363 );
xor \U$48988 ( \49365 , \49338 , \49364 );
xor \U$48989 ( \49366 , \49181 , \49188 );
xor \U$48990 ( \49367 , \49366 , \49196 );
and \U$48991 ( \49368 , \49365 , \49367 );
and \U$48992 ( \49369 , \49338 , \49364 );
or \U$48993 ( \49370 , \49368 , \49369 );
xor \U$48994 ( \49371 , \49336 , \49370 );
xor \U$48995 ( \49372 , \49047 , \49054 );
xor \U$48996 ( \49373 , \49372 , \49062 );
xor \U$48997 ( \49374 , \49075 , \49082 );
xor \U$48998 ( \49375 , \49374 , \49090 );
and \U$48999 ( \49376 , \49373 , \49375 );
xor \U$49000 ( \49377 , \48996 , \49003 );
xor \U$49001 ( \49378 , \49377 , \49011 );
xor \U$49002 ( \49379 , \49075 , \49082 );
xor \U$49003 ( \49380 , \49379 , \49090 );
and \U$49004 ( \49381 , \49378 , \49380 );
and \U$49005 ( \49382 , \49373 , \49378 );
or \U$49006 ( \49383 , \49376 , \49381 , \49382 );
and \U$49007 ( \49384 , \49371 , \49383 );
and \U$49008 ( \49385 , \49336 , \49370 );
or \U$49009 ( \49386 , \49384 , \49385 );
and \U$49010 ( \49387 , \4247 , RIae77bd0_92);
and \U$49011 ( \49388 , RIae77db0_96, \4245 );
nor \U$49012 ( \49389 , \49387 , \49388 );
and \U$49013 ( \49390 , \49389 , \4251 );
not \U$49014 ( \49391 , \49389 );
and \U$49015 ( \49392 , \49391 , \3989 );
nor \U$49016 ( \49393 , \49390 , \49392 );
not \U$49017 ( \49394 , \49393 );
and \U$49018 ( \49395 , \4688 , RIae77ea0_98);
and \U$49019 ( \49396 , RIae789e0_122, \4686 );
nor \U$49020 ( \49397 , \49395 , \49396 );
and \U$49021 ( \49398 , \49397 , \4482 );
not \U$49022 ( \49399 , \49397 );
and \U$49023 ( \49400 , \49399 , \4481 );
nor \U$49024 ( \49401 , \49398 , \49400 );
not \U$49025 ( \49402 , \49401 );
and \U$49026 ( \49403 , \49394 , \49402 );
and \U$49027 ( \49404 , \49401 , \49393 );
and \U$49028 ( \49405 , \5399 , RIae788f0_120);
and \U$49029 ( \49406 , RIae78800_118, \5397 );
nor \U$49030 ( \49407 , \49405 , \49406 );
and \U$49031 ( \49408 , \49407 , \5403 );
not \U$49032 ( \49409 , \49407 );
and \U$49033 ( \49410 , \49409 , \5016 );
nor \U$49034 ( \49411 , \49408 , \49410 );
nor \U$49035 ( \49412 , \49404 , \49411 );
nor \U$49036 ( \49413 , \49403 , \49412 );
and \U$49037 ( \49414 , \5896 , RIae78710_116);
and \U$49038 ( \49415 , RIae75bf0_24, \5894 );
nor \U$49039 ( \49416 , \49414 , \49415 );
and \U$49040 ( \49417 , \49416 , \5589 );
not \U$49041 ( \49418 , \49416 );
and \U$49042 ( \49419 , \49418 , \5590 );
nor \U$49043 ( \49420 , \49417 , \49419 );
not \U$49044 ( \49421 , \49420 );
and \U$49045 ( \49422 , \6172 , RIae75b00_22);
and \U$49046 ( \49423 , RIae75a10_20, \6170 );
nor \U$49047 ( \49424 , \49422 , \49423 );
and \U$49048 ( \49425 , \49424 , \6175 );
not \U$49049 ( \49426 , \49424 );
and \U$49050 ( \49427 , \49426 , \6176 );
nor \U$49051 ( \49428 , \49425 , \49427 );
not \U$49052 ( \49429 , \49428 );
and \U$49053 ( \49430 , \49421 , \49429 );
and \U$49054 ( \49431 , \49428 , \49420 );
and \U$49055 ( \49432 , \6941 , RIae75920_18);
and \U$49056 ( \49433 , RIae75fb0_32, \6939 );
nor \U$49057 ( \49434 , \49432 , \49433 );
and \U$49058 ( \49435 , \49434 , \6945 );
not \U$49059 ( \49436 , \49434 );
and \U$49060 ( \49437 , \49436 , \6314 );
nor \U$49061 ( \49438 , \49435 , \49437 );
nor \U$49062 ( \49439 , \49431 , \49438 );
nor \U$49063 ( \49440 , \49430 , \49439 );
xor \U$49064 ( \49441 , \49413 , \49440 );
and \U$49065 ( \49442 , \7633 , RIae75ec0_30);
and \U$49066 ( \49443 , RIae75ce0_26, \7631 );
nor \U$49067 ( \49444 , \49442 , \49443 );
and \U$49068 ( \49445 , \49444 , \7205 );
not \U$49069 ( \49446 , \49444 );
and \U$49070 ( \49447 , \49446 , \7206 );
nor \U$49071 ( \49448 , \49445 , \49447 );
not \U$49072 ( \49449 , \49448 );
and \U$49073 ( \49450 , \8371 , RIae75dd0_28);
and \U$49074 ( \49451 , RIae75650_12, \8369 );
nor \U$49075 ( \49452 , \49450 , \49451 );
and \U$49076 ( \49453 , \49452 , \8019 );
not \U$49077 ( \49454 , \49452 );
and \U$49078 ( \49455 , \49454 , \8020 );
nor \U$49079 ( \49456 , \49453 , \49455 );
not \U$49080 ( \49457 , \49456 );
and \U$49081 ( \49458 , \49449 , \49457 );
and \U$49082 ( \49459 , \49456 , \49448 );
and \U$49083 ( \49460 , \8966 , RIae75560_10);
and \U$49084 ( \49461 , RIae75830_16, \8964 );
nor \U$49085 ( \49462 , \49460 , \49461 );
and \U$49086 ( \49463 , \49462 , \8789 );
not \U$49087 ( \49464 , \49462 );
and \U$49088 ( \49465 , \49464 , \8799 );
nor \U$49089 ( \49466 , \49463 , \49465 );
nor \U$49090 ( \49467 , \49459 , \49466 );
nor \U$49091 ( \49468 , \49458 , \49467 );
and \U$49092 ( \49469 , \49441 , \49468 );
and \U$49093 ( \49470 , \49413 , \49440 );
nor \U$49094 ( \49471 , \49469 , \49470 );
and \U$49095 ( \49472 , \10548 , RIae751a0_2);
and \U$49096 ( \49473 , RIae75380_6, \10546 );
nor \U$49097 ( \49474 , \49472 , \49473 );
and \U$49098 ( \49475 , \49474 , \10421 );
not \U$49099 ( \49476 , \49474 );
and \U$49100 ( \49477 , \49476 , \10118 );
nor \U$49101 ( \49478 , \49475 , \49477 );
and \U$49102 ( \49479 , \9760 , RIae75740_14);
and \U$49103 ( \49480 , RIae75290_4, \9758 );
nor \U$49104 ( \49481 , \49479 , \49480 );
and \U$49105 ( \49482 , \49481 , \9273 );
not \U$49106 ( \49483 , \49481 );
and \U$49107 ( \49484 , \49483 , \9272 );
nor \U$49108 ( \49485 , \49482 , \49484 );
xor \U$49109 ( \49486 , \49478 , \49485 );
and \U$49110 ( \49487 , \11470 , RIae75470_8);
and \U$49111 ( \49488 , RIae76460_42, \11468 );
nor \U$49112 ( \49489 , \49487 , \49488 );
and \U$49113 ( \49490 , \49489 , \10936 );
not \U$49114 ( \49491 , \49489 );
and \U$49115 ( \49492 , \49491 , \11474 );
nor \U$49116 ( \49493 , \49490 , \49492 );
and \U$49117 ( \49494 , \49486 , \49493 );
and \U$49118 ( \49495 , \49478 , \49485 );
or \U$49119 ( \49496 , \49494 , \49495 );
and \U$49120 ( \49497 , \15726 , RIae76a00_54);
and \U$49121 ( \49498 , RIae76820_50, RIae7aab0_192);
nor \U$49122 ( \49499 , \49497 , \49498 );
and \U$49123 ( \49500 , \49499 , \14959 );
not \U$49124 ( \49501 , \49499 );
and \U$49125 ( \49502 , \49501 , RIae7aa38_191);
nor \U$49126 ( \49503 , \49500 , \49502 );
xor \U$49127 ( \49504 , \49503 , \469 );
and \U$49128 ( \49505 , \14964 , RIae76280_38);
and \U$49129 ( \49506 , RIae76af0_56, \14962 );
nor \U$49130 ( \49507 , \49505 , \49506 );
and \U$49131 ( \49508 , \49507 , \14463 );
not \U$49132 ( \49509 , \49507 );
and \U$49133 ( \49510 , \49509 , \14462 );
nor \U$49134 ( \49511 , \49508 , \49510 );
and \U$49135 ( \49512 , \49504 , \49511 );
and \U$49136 ( \49513 , \49503 , \469 );
or \U$49137 ( \49514 , \49512 , \49513 );
xor \U$49138 ( \49515 , \49496 , \49514 );
and \U$49139 ( \49516 , \12180 , RIae76550_44);
and \U$49140 ( \49517 , RIae76730_48, \12178 );
nor \U$49141 ( \49518 , \49516 , \49517 );
and \U$49142 ( \49519 , \49518 , \12184 );
not \U$49143 ( \49520 , \49518 );
and \U$49144 ( \49521 , \49520 , \11827 );
nor \U$49145 ( \49522 , \49519 , \49521 );
and \U$49146 ( \49523 , \13059 , RIae76640_46);
and \U$49147 ( \49524 , RIae76190_36, \13057 );
nor \U$49148 ( \49525 , \49523 , \49524 );
and \U$49149 ( \49526 , \49525 , \13063 );
not \U$49150 ( \49527 , \49525 );
and \U$49151 ( \49528 , \49527 , \12718 );
nor \U$49152 ( \49529 , \49526 , \49528 );
xor \U$49153 ( \49530 , \49522 , \49529 );
and \U$49154 ( \49531 , \14059 , RIae760a0_34);
and \U$49155 ( \49532 , RIae76370_40, \14057 );
nor \U$49156 ( \49533 , \49531 , \49532 );
and \U$49157 ( \49534 , \49533 , \13502 );
not \U$49158 ( \49535 , \49533 );
and \U$49159 ( \49536 , \49535 , \14063 );
nor \U$49160 ( \49537 , \49534 , \49536 );
and \U$49161 ( \49538 , \49530 , \49537 );
and \U$49162 ( \49539 , \49522 , \49529 );
or \U$49163 ( \49540 , \49538 , \49539 );
and \U$49164 ( \49541 , \49515 , \49540 );
and \U$49165 ( \49542 , \49496 , \49514 );
or \U$49166 ( \49543 , \49541 , \49542 );
xor \U$49167 ( \49544 , \49471 , \49543 );
and \U$49168 ( \49545 , \3730 , RIae784b8_111);
and \U$49169 ( \49546 , RIae77cc0_94, \3728 );
nor \U$49170 ( \49547 , \49545 , \49546 );
and \U$49171 ( \49548 , \49547 , \3732 );
not \U$49172 ( \49549 , \49547 );
and \U$49173 ( \49550 , \49549 , \3422 );
nor \U$49174 ( \49551 , \49548 , \49550 );
not \U$49175 ( \49552 , \3089 );
and \U$49176 ( \49553 , \2783 , RIae78080_102);
and \U$49177 ( \49554 , RIae78260_106, \2781 );
nor \U$49178 ( \49555 , \49553 , \49554 );
not \U$49179 ( \49556 , \49555 );
or \U$49180 ( \49557 , \49552 , \49556 );
or \U$49181 ( \49558 , \49555 , \2789 );
nand \U$49182 ( \49559 , \49557 , \49558 );
xor \U$49183 ( \49560 , \49551 , \49559 );
not \U$49184 ( \49561 , \2774 );
and \U$49185 ( \49562 , \3214 , RIae78620_114);
and \U$49186 ( \49563 , RIae78440_110, \3212 );
nor \U$49187 ( \49564 , \49562 , \49563 );
not \U$49188 ( \49565 , \49564 );
or \U$49189 ( \49566 , \49561 , \49565 );
or \U$49190 ( \49567 , \49564 , \3218 );
nand \U$49191 ( \49568 , \49566 , \49567 );
and \U$49192 ( \49569 , \49560 , \49568 );
and \U$49193 ( \49570 , \49551 , \49559 );
or \U$49194 ( \49571 , \49569 , \49570 );
and \U$49195 ( \49572 , \1939 , RIae77090_68);
and \U$49196 ( \49573 , RIae77270_72, \1937 );
nor \U$49197 ( \49574 , \49572 , \49573 );
and \U$49198 ( \49575 , \49574 , \1735 );
not \U$49199 ( \49576 , \49574 );
and \U$49200 ( \49577 , \49576 , \1734 );
nor \U$49201 ( \49578 , \49575 , \49577 );
and \U$49202 ( \49579 , \2224 , RIae77360_74);
and \U$49203 ( \49580 , RIae78350_108, \2222 );
nor \U$49204 ( \49581 , \49579 , \49580 );
and \U$49205 ( \49582 , \49581 , \2061 );
not \U$49206 ( \49583 , \49581 );
and \U$49207 ( \49584 , \49583 , \2060 );
nor \U$49208 ( \49585 , \49582 , \49584 );
xor \U$49209 ( \49586 , \49578 , \49585 );
and \U$49210 ( \49587 , \2607 , RIae78170_104);
and \U$49211 ( \49588 , RIae77f90_100, \2605 );
nor \U$49212 ( \49589 , \49587 , \49588 );
and \U$49213 ( \49590 , \49589 , \2611 );
not \U$49214 ( \49591 , \49589 );
and \U$49215 ( \49592 , \49591 , \2397 );
nor \U$49216 ( \49593 , \49590 , \49592 );
and \U$49217 ( \49594 , \49586 , \49593 );
and \U$49218 ( \49595 , \49578 , \49585 );
or \U$49219 ( \49596 , \49594 , \49595 );
xor \U$49220 ( \49597 , \49571 , \49596 );
and \U$49221 ( \49598 , \1593 , RIae76cd0_60);
and \U$49222 ( \49599 , RIae77108_69, \1591 );
nor \U$49223 ( \49600 , \49598 , \49599 );
and \U$49224 ( \49601 , \49600 , \1498 );
not \U$49225 ( \49602 , \49600 );
and \U$49226 ( \49603 , \49602 , \1488 );
nor \U$49227 ( \49604 , \49601 , \49603 );
and \U$49228 ( \49605 , \1138 , RIae77900_86);
and \U$49229 ( \49606 , RIae76fa0_66, \1136 );
nor \U$49230 ( \49607 , \49605 , \49606 );
and \U$49231 ( \49608 , \49607 , \1012 );
not \U$49232 ( \49609 , \49607 );
and \U$49233 ( \49610 , \49609 , \1142 );
nor \U$49234 ( \49611 , \49608 , \49610 );
xor \U$49235 ( \49612 , \49604 , \49611 );
and \U$49236 ( \49613 , \1376 , RIae76eb0_64);
and \U$49237 ( \49614 , RIae76dc0_62, \1374 );
nor \U$49238 ( \49615 , \49613 , \49614 );
and \U$49239 ( \49616 , \49615 , \1380 );
not \U$49240 ( \49617 , \49615 );
and \U$49241 ( \49618 , \49617 , \1261 );
nor \U$49242 ( \49619 , \49616 , \49618 );
and \U$49243 ( \49620 , \49612 , \49619 );
and \U$49244 ( \49621 , \49604 , \49611 );
or \U$49245 ( \49622 , \49620 , \49621 );
and \U$49246 ( \49623 , \49597 , \49622 );
and \U$49247 ( \49624 , \49571 , \49596 );
or \U$49248 ( \49625 , \49623 , \49624 );
and \U$49249 ( \49626 , \49544 , \49625 );
and \U$49250 ( \49627 , \49471 , \49543 );
or \U$49251 ( \49628 , \49626 , \49627 );
xor \U$49252 ( \49629 , \49386 , \49628 );
xor \U$49253 ( \49630 , \48684 , \48691 );
xor \U$49254 ( \49631 , \49630 , \48699 );
xor \U$49255 ( \49632 , \48976 , \48981 );
xor \U$49256 ( \49633 , \49631 , \49632 );
xor \U$49257 ( \49634 , \48932 , \48934 );
xor \U$49258 ( \49635 , \49634 , \48937 );
and \U$49259 ( \49636 , \49633 , \49635 );
xor \U$49260 ( \49637 , \48585 , \400 );
xor \U$49261 ( \49638 , \49637 , \48593 );
xor \U$49262 ( \49639 , \49236 , \49241 );
xor \U$49263 ( \49640 , \49638 , \49639 );
xor \U$49264 ( \49641 , \48932 , \48934 );
xor \U$49265 ( \49642 , \49641 , \48937 );
and \U$49266 ( \49643 , \49640 , \49642 );
and \U$49267 ( \49644 , \49633 , \49640 );
or \U$49268 ( \49645 , \49636 , \49643 , \49644 );
and \U$49269 ( \49646 , \49629 , \49645 );
and \U$49270 ( \49647 , \49386 , \49628 );
or \U$49271 ( \49648 , \49646 , \49647 );
xor \U$49272 ( \49649 , \48578 , \48596 );
xor \U$49273 ( \49650 , \49649 , \48622 );
xor \U$49274 ( \49651 , \49262 , \49267 );
xor \U$49275 ( \49652 , \49650 , \49651 );
xor \U$49276 ( \49653 , \49173 , \49199 );
xor \U$49277 ( \49654 , \49653 , \49227 );
xor \U$49278 ( \49655 , \49014 , \49039 );
xor \U$49279 ( \49656 , \49655 , \49065 );
and \U$49280 ( \49657 , \49654 , \49656 );
xor \U$49281 ( \49658 , \48966 , \48967 );
xor \U$49282 ( \49659 , \49658 , \48970 );
xor \U$49283 ( \49660 , \49014 , \49039 );
xor \U$49284 ( \49661 , \49660 , \49065 );
and \U$49285 ( \49662 , \49659 , \49661 );
and \U$49286 ( \49663 , \49654 , \49659 );
or \U$49287 ( \49664 , \49657 , \49662 , \49663 );
xor \U$49288 ( \49665 , \49652 , \49664 );
xor \U$49289 ( \49666 , \48395 , \48397 );
xor \U$49290 ( \49667 , \49666 , \48400 );
xor \U$49291 ( \49668 , \49277 , \49284 );
xor \U$49292 ( \49669 , \49667 , \49668 );
and \U$49293 ( \49670 , \49665 , \49669 );
and \U$49294 ( \49671 , \49652 , \49664 );
or \U$49295 ( \49672 , \49670 , \49671 );
xor \U$49296 ( \49673 , \49648 , \49672 );
xor \U$49297 ( \49674 , \49068 , \49147 );
xor \U$49298 ( \49675 , \49674 , \49230 );
xor \U$49299 ( \49676 , \49246 , \49248 );
xor \U$49300 ( \49677 , \49676 , \49253 );
and \U$49301 ( \49678 , \49675 , \49677 );
xor \U$49302 ( \49679 , \48940 , \48973 );
xor \U$49303 ( \49680 , \49679 , \48986 );
xor \U$49304 ( \49681 , \49246 , \49248 );
xor \U$49305 ( \49682 , \49681 , \49253 );
and \U$49306 ( \49683 , \49680 , \49682 );
and \U$49307 ( \49684 , \49675 , \49680 );
or \U$49308 ( \49685 , \49678 , \49683 , \49684 );
and \U$49309 ( \49686 , \49673 , \49685 );
and \U$49310 ( \49687 , \49648 , \49672 );
or \U$49311 ( \49688 , \49686 , \49687 );
xor \U$49312 ( \49689 , \48553 , \48625 );
xor \U$49313 ( \49690 , \49689 , \48705 );
xor \U$49314 ( \49691 , \48403 , \48456 );
xor \U$49315 ( \49692 , \49691 , \48469 );
and \U$49316 ( \49693 , \49690 , \49692 );
xor \U$49317 ( \49694 , \48749 , \48751 );
xor \U$49318 ( \49695 , \49694 , \48754 );
xor \U$49319 ( \49696 , \48918 , \48925 );
xor \U$49320 ( \49697 , \49695 , \49696 );
xor \U$49321 ( \49698 , \48403 , \48456 );
xor \U$49322 ( \49699 , \49698 , \48469 );
and \U$49323 ( \49700 , \49697 , \49699 );
and \U$49324 ( \49701 , \49690 , \49697 );
or \U$49325 ( \49702 , \49693 , \49700 , \49701 );
xor \U$49326 ( \49703 , \49688 , \49702 );
xor \U$49327 ( \49704 , \48128 , \48370 );
xor \U$49328 ( \49705 , \49704 , \48390 );
xor \U$49329 ( \49706 , \48896 , \48901 );
xor \U$49330 ( \49707 , \49705 , \49706 );
and \U$49331 ( \49708 , \49703 , \49707 );
and \U$49332 ( \49709 , \49688 , \49702 );
or \U$49333 ( \49710 , \49708 , \49709 );
xor \U$49334 ( \49711 , \49324 , \49710 );
not \U$49335 ( \49712 , \48912 );
not \U$49336 ( \49713 , \48906 );
not \U$49337 ( \49714 , \49295 );
and \U$49338 ( \49715 , \49713 , \49714 );
and \U$49339 ( \49716 , \48906 , \49295 );
nor \U$49340 ( \49717 , \49715 , \49716 );
not \U$49341 ( \49718 , \49717 );
or \U$49342 ( \49719 , \49712 , \49718 );
or \U$49343 ( \49720 , \49717 , \48912 );
nand \U$49344 ( \49721 , \49719 , \49720 );
and \U$49345 ( \49722 , \49711 , \49721 );
and \U$49346 ( \49723 , \49324 , \49710 );
or \U$49347 ( \49724 , \49722 , \49723 );
not \U$49348 ( \49725 , \48890 );
not \U$49349 ( \49726 , \48893 );
or \U$49350 ( \49727 , \49725 , \49726 );
or \U$49351 ( \49728 , \48893 , \48890 );
nand \U$49352 ( \49729 , \49727 , \49728 );
xor \U$49353 ( \49730 , \49724 , \49729 );
not \U$49354 ( \49731 , \49302 );
xor \U$49355 ( \49732 , \49315 , \49297 );
not \U$49356 ( \49733 , \49732 );
or \U$49357 ( \49734 , \49731 , \49733 );
or \U$49358 ( \49735 , \49732 , \49302 );
nand \U$49359 ( \49736 , \49734 , \49735 );
and \U$49360 ( \49737 , \49730 , \49736 );
and \U$49361 ( \49738 , \49724 , \49729 );
or \U$49362 ( \49739 , \49737 , \49738 );
and \U$49363 ( \49740 , \49322 , \49739 );
xor \U$49364 ( \49741 , \49739 , \49322 );
xor \U$49365 ( \49742 , \49688 , \49702 );
xor \U$49366 ( \49743 , \49742 , \49707 );
not \U$49367 ( \49744 , \49743 );
xor \U$49368 ( \49745 , \48930 , \49259 );
xor \U$49369 ( \49746 , \49745 , \49292 );
xor \U$49370 ( \49747 , \49471 , \49543 );
xor \U$49371 ( \49748 , \49747 , \49625 );
xor \U$49372 ( \49749 , \49336 , \49370 );
xor \U$49373 ( \49750 , \49749 , \49383 );
and \U$49374 ( \49751 , \49748 , \49750 );
xor \U$49375 ( \49752 , \48932 , \48934 );
xor \U$49376 ( \49753 , \49752 , \48937 );
xor \U$49377 ( \49754 , \49633 , \49640 );
xor \U$49378 ( \49755 , \49753 , \49754 );
xor \U$49379 ( \49756 , \49336 , \49370 );
xor \U$49380 ( \49757 , \49756 , \49383 );
and \U$49381 ( \49758 , \49755 , \49757 );
and \U$49382 ( \49759 , \49748 , \49755 );
or \U$49383 ( \49760 , \49751 , \49758 , \49759 );
xor \U$49384 ( \49761 , \49126 , \49133 );
xor \U$49385 ( \49762 , \49761 , \49141 );
xor \U$49386 ( \49763 , \49100 , \49107 );
xor \U$49387 ( \49764 , \49763 , \49115 );
xor \U$49388 ( \49765 , \49762 , \49764 );
xor \U$49389 ( \49766 , \49075 , \49082 );
xor \U$49390 ( \49767 , \49766 , \49090 );
xor \U$49391 ( \49768 , \49373 , \49378 );
xor \U$49392 ( \49769 , \49767 , \49768 );
and \U$49393 ( \49770 , \49765 , \49769 );
and \U$49394 ( \49771 , \49762 , \49764 );
or \U$49395 ( \49772 , \49770 , \49771 );
and \U$49396 ( \49773 , \3730 , RIae78440_110);
and \U$49397 ( \49774 , RIae784b8_111, \3728 );
nor \U$49398 ( \49775 , \49773 , \49774 );
and \U$49399 ( \49776 , \49775 , \3422 );
not \U$49400 ( \49777 , \49775 );
and \U$49401 ( \49778 , \49777 , \3732 );
nor \U$49402 ( \49779 , \49776 , \49778 );
not \U$49403 ( \49780 , \49779 );
and \U$49404 ( \49781 , \4247 , RIae77cc0_94);
and \U$49405 ( \49782 , RIae77bd0_92, \4245 );
nor \U$49406 ( \49783 , \49781 , \49782 );
and \U$49407 ( \49784 , \49783 , \4251 );
not \U$49408 ( \49785 , \49783 );
and \U$49409 ( \49786 , \49785 , \3989 );
nor \U$49410 ( \49787 , \49784 , \49786 );
not \U$49411 ( \49788 , \49787 );
and \U$49412 ( \49789 , \49780 , \49788 );
and \U$49413 ( \49790 , \49787 , \49779 );
and \U$49414 ( \49791 , \4688 , RIae77db0_96);
and \U$49415 ( \49792 , RIae77ea0_98, \4686 );
nor \U$49416 ( \49793 , \49791 , \49792 );
and \U$49417 ( \49794 , \49793 , \4482 );
not \U$49418 ( \49795 , \49793 );
and \U$49419 ( \49796 , \49795 , \4481 );
nor \U$49420 ( \49797 , \49794 , \49796 );
nor \U$49421 ( \49798 , \49790 , \49797 );
nor \U$49422 ( \49799 , \49789 , \49798 );
and \U$49423 ( \49800 , \5896 , RIae78800_118);
and \U$49424 ( \49801 , RIae78710_116, \5894 );
nor \U$49425 ( \49802 , \49800 , \49801 );
and \U$49426 ( \49803 , \49802 , \5590 );
not \U$49427 ( \49804 , \49802 );
and \U$49428 ( \49805 , \49804 , \5589 );
nor \U$49429 ( \49806 , \49803 , \49805 );
and \U$49430 ( \49807 , \6172 , RIae75bf0_24);
and \U$49431 ( \49808 , RIae75b00_22, \6170 );
nor \U$49432 ( \49809 , \49807 , \49808 );
and \U$49433 ( \49810 , \49809 , \6176 );
not \U$49434 ( \49811 , \49809 );
and \U$49435 ( \49812 , \49811 , \6175 );
nor \U$49436 ( \49813 , \49810 , \49812 );
xor \U$49437 ( \49814 , \49806 , \49813 );
and \U$49438 ( \49815 , \5399 , RIae789e0_122);
and \U$49439 ( \49816 , RIae788f0_120, \5397 );
nor \U$49440 ( \49817 , \49815 , \49816 );
and \U$49441 ( \49818 , \49817 , \5016 );
not \U$49442 ( \49819 , \49817 );
and \U$49443 ( \49820 , \49819 , \5403 );
nor \U$49444 ( \49821 , \49818 , \49820 );
and \U$49445 ( \49822 , \49814 , \49821 );
and \U$49446 ( \49823 , \49806 , \49813 );
nor \U$49447 ( \49824 , \49822 , \49823 );
xor \U$49448 ( \49825 , \49799 , \49824 );
and \U$49449 ( \49826 , \6941 , RIae75a10_20);
and \U$49450 ( \49827 , RIae75920_18, \6939 );
nor \U$49451 ( \49828 , \49826 , \49827 );
and \U$49452 ( \49829 , \49828 , \6945 );
not \U$49453 ( \49830 , \49828 );
and \U$49454 ( \49831 , \49830 , \6314 );
nor \U$49455 ( \49832 , \49829 , \49831 );
not \U$49456 ( \49833 , \49832 );
and \U$49457 ( \49834 , \7633 , RIae75fb0_32);
and \U$49458 ( \49835 , RIae75ec0_30, \7631 );
nor \U$49459 ( \49836 , \49834 , \49835 );
and \U$49460 ( \49837 , \49836 , \7205 );
not \U$49461 ( \49838 , \49836 );
and \U$49462 ( \49839 , \49838 , \7206 );
nor \U$49463 ( \49840 , \49837 , \49839 );
not \U$49464 ( \49841 , \49840 );
and \U$49465 ( \49842 , \49833 , \49841 );
and \U$49466 ( \49843 , \49840 , \49832 );
and \U$49467 ( \49844 , \8371 , RIae75ce0_26);
and \U$49468 ( \49845 , RIae75dd0_28, \8369 );
nor \U$49469 ( \49846 , \49844 , \49845 );
and \U$49470 ( \49847 , \49846 , \8019 );
not \U$49471 ( \49848 , \49846 );
and \U$49472 ( \49849 , \49848 , \8020 );
nor \U$49473 ( \49850 , \49847 , \49849 );
nor \U$49474 ( \49851 , \49843 , \49850 );
nor \U$49475 ( \49852 , \49842 , \49851 );
and \U$49476 ( \49853 , \49825 , \49852 );
and \U$49477 ( \49854 , \49799 , \49824 );
nor \U$49478 ( \49855 , \49853 , \49854 );
and \U$49479 ( \49856 , \1138 , RIae77810_84);
and \U$49480 ( \49857 , RIae77900_86, \1136 );
nor \U$49481 ( \49858 , \49856 , \49857 );
and \U$49482 ( \49859 , \49858 , \1012 );
not \U$49483 ( \49860 , \49858 );
and \U$49484 ( \49861 , \49860 , \1142 );
nor \U$49485 ( \49862 , \49859 , \49861 );
and \U$49486 ( \49863 , \1376 , RIae76fa0_66);
and \U$49487 ( \49864 , RIae76eb0_64, \1374 );
nor \U$49488 ( \49865 , \49863 , \49864 );
and \U$49489 ( \49866 , \49865 , \1380 );
not \U$49490 ( \49867 , \49865 );
and \U$49491 ( \49868 , \49867 , \1261 );
nor \U$49492 ( \49869 , \49866 , \49868 );
xor \U$49493 ( \49870 , \49862 , \49869 );
not \U$49494 ( \49871 , \787 );
and \U$49495 ( \49872 , \883 , RIae77ae0_90);
and \U$49496 ( \49873 , RIae779f0_88, \881 );
nor \U$49497 ( \49874 , \49872 , \49873 );
not \U$49498 ( \49875 , \49874 );
or \U$49499 ( \49876 , \49871 , \49875 );
or \U$49500 ( \49877 , \49874 , \787 );
nand \U$49501 ( \49878 , \49876 , \49877 );
and \U$49502 ( \49879 , \49870 , \49878 );
and \U$49503 ( \49880 , \49862 , \49869 );
nor \U$49504 ( \49881 , \49879 , \49880 );
and \U$49505 ( \49882 , \1939 , RIae77108_69);
and \U$49506 ( \49883 , RIae77090_68, \1937 );
nor \U$49507 ( \49884 , \49882 , \49883 );
and \U$49508 ( \49885 , \49884 , \1735 );
not \U$49509 ( \49886 , \49884 );
and \U$49510 ( \49887 , \49886 , \1734 );
nor \U$49511 ( \49888 , \49885 , \49887 );
and \U$49512 ( \49889 , \2224 , RIae77270_72);
and \U$49513 ( \49890 , RIae77360_74, \2222 );
nor \U$49514 ( \49891 , \49889 , \49890 );
and \U$49515 ( \49892 , \49891 , \2061 );
not \U$49516 ( \49893 , \49891 );
and \U$49517 ( \49894 , \49893 , \2060 );
nor \U$49518 ( \49895 , \49892 , \49894 );
xor \U$49519 ( \49896 , \49888 , \49895 );
and \U$49520 ( \49897 , \1593 , RIae76dc0_62);
and \U$49521 ( \49898 , RIae76cd0_60, \1591 );
nor \U$49522 ( \49899 , \49897 , \49898 );
and \U$49523 ( \49900 , \49899 , \1498 );
not \U$49524 ( \49901 , \49899 );
and \U$49525 ( \49902 , \49901 , \1488 );
nor \U$49526 ( \49903 , \49900 , \49902 );
and \U$49527 ( \49904 , \49896 , \49903 );
and \U$49528 ( \49905 , \49888 , \49895 );
nor \U$49529 ( \49906 , \49904 , \49905 );
xor \U$49530 ( \49907 , \49881 , \49906 );
and \U$49531 ( \49908 , \2607 , RIae78350_108);
and \U$49532 ( \49909 , RIae78170_104, \2605 );
nor \U$49533 ( \49910 , \49908 , \49909 );
and \U$49534 ( \49911 , \49910 , \2397 );
not \U$49535 ( \49912 , \49910 );
and \U$49536 ( \49913 , \49912 , \2611 );
nor \U$49537 ( \49914 , \49911 , \49913 );
not \U$49538 ( \49915 , \49914 );
and \U$49539 ( \49916 , \2783 , RIae77f90_100);
and \U$49540 ( \49917 , RIae78080_102, \2781 );
nor \U$49541 ( \49918 , \49916 , \49917 );
not \U$49542 ( \49919 , \49918 );
not \U$49543 ( \49920 , \2789 );
and \U$49544 ( \49921 , \49919 , \49920 );
and \U$49545 ( \49922 , \49918 , \3089 );
nor \U$49546 ( \49923 , \49921 , \49922 );
not \U$49547 ( \49924 , \49923 );
and \U$49548 ( \49925 , \49915 , \49924 );
and \U$49549 ( \49926 , \49923 , \49914 );
and \U$49550 ( \49927 , \3214 , RIae78260_106);
and \U$49551 ( \49928 , RIae78620_114, \3212 );
nor \U$49552 ( \49929 , \49927 , \49928 );
not \U$49553 ( \49930 , \49929 );
not \U$49554 ( \49931 , \3218 );
and \U$49555 ( \49932 , \49930 , \49931 );
and \U$49556 ( \49933 , \49929 , \3218 );
nor \U$49557 ( \49934 , \49932 , \49933 );
nor \U$49558 ( \49935 , \49926 , \49934 );
nor \U$49559 ( \49936 , \49925 , \49935 );
and \U$49560 ( \49937 , \49907 , \49936 );
and \U$49561 ( \49938 , \49881 , \49906 );
nor \U$49562 ( \49939 , \49937 , \49938 );
xor \U$49563 ( \49940 , \49855 , \49939 );
and \U$49564 ( \49941 , \9760 , RIae75830_16);
and \U$49565 ( \49942 , RIae75740_14, \9758 );
nor \U$49566 ( \49943 , \49941 , \49942 );
and \U$49567 ( \49944 , \49943 , \9273 );
not \U$49568 ( \49945 , \49943 );
and \U$49569 ( \49946 , \49945 , \9764 );
nor \U$49570 ( \49947 , \49944 , \49946 );
and \U$49571 ( \49948 , \10548 , RIae75290_4);
and \U$49572 ( \49949 , RIae751a0_2, \10546 );
nor \U$49573 ( \49950 , \49948 , \49949 );
and \U$49574 ( \49951 , \49950 , \10421 );
not \U$49575 ( \49952 , \49950 );
and \U$49576 ( \49953 , \49952 , \10118 );
nor \U$49577 ( \49954 , \49951 , \49953 );
xor \U$49578 ( \49955 , \49947 , \49954 );
and \U$49579 ( \49956 , \8966 , RIae75650_12);
and \U$49580 ( \49957 , RIae75560_10, \8964 );
nor \U$49581 ( \49958 , \49956 , \49957 );
and \U$49582 ( \49959 , \49958 , \8799 );
not \U$49583 ( \49960 , \49958 );
and \U$49584 ( \49961 , \49960 , \8789 );
nor \U$49585 ( \49962 , \49959 , \49961 );
and \U$49586 ( \49963 , \49955 , \49962 );
and \U$49587 ( \49964 , \49947 , \49954 );
nor \U$49588 ( \49965 , \49963 , \49964 );
and \U$49589 ( \49966 , \11470 , RIae75380_6);
and \U$49590 ( \49967 , RIae75470_8, \11468 );
nor \U$49591 ( \49968 , \49966 , \49967 );
and \U$49592 ( \49969 , \49968 , \11474 );
not \U$49593 ( \49970 , \49968 );
and \U$49594 ( \49971 , \49970 , \10936 );
nor \U$49595 ( \49972 , \49969 , \49971 );
not \U$49596 ( \49973 , \49972 );
and \U$49597 ( \49974 , \13059 , RIae76730_48);
and \U$49598 ( \49975 , RIae76640_46, \13057 );
nor \U$49599 ( \49976 , \49974 , \49975 );
and \U$49600 ( \49977 , \49976 , \12718 );
not \U$49601 ( \49978 , \49976 );
and \U$49602 ( \49979 , \49978 , \13063 );
nor \U$49603 ( \49980 , \49977 , \49979 );
not \U$49604 ( \49981 , \49980 );
and \U$49605 ( \49982 , \49973 , \49981 );
and \U$49606 ( \49983 , \49980 , \49972 );
and \U$49607 ( \49984 , \12180 , RIae76460_42);
and \U$49608 ( \49985 , RIae76550_44, \12178 );
nor \U$49609 ( \49986 , \49984 , \49985 );
and \U$49610 ( \49987 , \49986 , \11827 );
not \U$49611 ( \49988 , \49986 );
and \U$49612 ( \49989 , \49988 , \12184 );
nor \U$49613 ( \49990 , \49987 , \49989 );
nor \U$49614 ( \49991 , \49983 , \49990 );
nor \U$49615 ( \49992 , \49982 , \49991 );
or \U$49616 ( \49993 , \49965 , \49992 );
not \U$49617 ( \49994 , \49965 );
not \U$49618 ( \49995 , \49992 );
or \U$49619 ( \49996 , \49994 , \49995 );
and \U$49620 ( \49997 , \14059 , RIae76190_36);
and \U$49621 ( \49998 , RIae760a0_34, \14057 );
nor \U$49622 ( \49999 , \49997 , \49998 );
and \U$49623 ( \50000 , \49999 , \13502 );
not \U$49624 ( \50001 , \49999 );
and \U$49625 ( \50002 , \50001 , \14063 );
nor \U$49626 ( \50003 , \50000 , \50002 );
and \U$49627 ( \50004 , \15726 , RIae76af0_56);
and \U$49628 ( \50005 , RIae76a00_54, RIae7aab0_192);
nor \U$49629 ( \50006 , \50004 , \50005 );
and \U$49630 ( \50007 , \50006 , \14959 );
not \U$49631 ( \50008 , \50006 );
and \U$49632 ( \50009 , \50008 , RIae7aa38_191);
nor \U$49633 ( \50010 , \50007 , \50009 );
xor \U$49634 ( \50011 , \50003 , \50010 );
and \U$49635 ( \50012 , \14964 , RIae76370_40);
and \U$49636 ( \50013 , RIae76280_38, \14962 );
nor \U$49637 ( \50014 , \50012 , \50013 );
and \U$49638 ( \50015 , \50014 , \14463 );
not \U$49639 ( \50016 , \50014 );
and \U$49640 ( \50017 , \50016 , \14462 );
nor \U$49641 ( \50018 , \50015 , \50017 );
and \U$49642 ( \50019 , \50011 , \50018 );
and \U$49643 ( \50020 , \50003 , \50010 );
or \U$49644 ( \50021 , \50019 , \50020 );
nand \U$49645 ( \50022 , \49996 , \50021 );
nand \U$49646 ( \50023 , \49993 , \50022 );
and \U$49647 ( \50024 , \49940 , \50023 );
and \U$49648 ( \50025 , \49855 , \49939 );
or \U$49649 ( \50026 , \50024 , \50025 );
xor \U$49650 ( \50027 , \49772 , \50026 );
xor \U$49651 ( \50028 , \49578 , \49585 );
xor \U$49652 ( \50029 , \50028 , \49593 );
xor \U$49653 ( \50030 , \49551 , \49559 );
xor \U$49654 ( \50031 , \50030 , \49568 );
xor \U$49655 ( \50032 , \50029 , \50031 );
not \U$49656 ( \50033 , \49393 );
xor \U$49657 ( \50034 , \49401 , \49411 );
not \U$49658 ( \50035 , \50034 );
or \U$49659 ( \50036 , \50033 , \50035 );
or \U$49660 ( \50037 , \50034 , \49393 );
nand \U$49661 ( \50038 , \50036 , \50037 );
and \U$49662 ( \50039 , \50032 , \50038 );
and \U$49663 ( \50040 , \50029 , \50031 );
or \U$49664 ( \50041 , \50039 , \50040 );
nand \U$49665 ( \50042 , RIae77630_80, \512 );
not \U$49666 ( \50043 , \50042 );
not \U$49667 ( \50044 , \469 );
or \U$49668 ( \50045 , \50043 , \50044 );
or \U$49669 ( \50046 , \469 , \50042 );
nand \U$49670 ( \50047 , \50045 , \50046 );
xor \U$49671 ( \50048 , \49604 , \49611 );
xor \U$49672 ( \50049 , \50048 , \49619 );
and \U$49673 ( \50050 , \50047 , \50049 );
xor \U$49674 ( \50051 , \49345 , \49352 );
xor \U$49675 ( \50052 , \50051 , \49361 );
xor \U$49676 ( \50053 , \49604 , \49611 );
xor \U$49677 ( \50054 , \50053 , \49619 );
and \U$49678 ( \50055 , \50052 , \50054 );
and \U$49679 ( \50056 , \50047 , \50052 );
or \U$49680 ( \50057 , \50050 , \50055 , \50056 );
xor \U$49681 ( \50058 , \50041 , \50057 );
not \U$49682 ( \50059 , \49448 );
xor \U$49683 ( \50060 , \49456 , \49466 );
not \U$49684 ( \50061 , \50060 );
or \U$49685 ( \50062 , \50059 , \50061 );
or \U$49686 ( \50063 , \50060 , \49448 );
nand \U$49687 ( \50064 , \50062 , \50063 );
not \U$49688 ( \50065 , \49420 );
xor \U$49689 ( \50066 , \49428 , \49438 );
not \U$49690 ( \50067 , \50066 );
or \U$49691 ( \50068 , \50065 , \50067 );
or \U$49692 ( \50069 , \50066 , \49420 );
nand \U$49693 ( \50070 , \50068 , \50069 );
xor \U$49694 ( \50071 , \50064 , \50070 );
xor \U$49695 ( \50072 , \49478 , \49485 );
xor \U$49696 ( \50073 , \50072 , \49493 );
and \U$49697 ( \50074 , \50071 , \50073 );
and \U$49698 ( \50075 , \50064 , \50070 );
or \U$49699 ( \50076 , \50074 , \50075 );
and \U$49700 ( \50077 , \50058 , \50076 );
and \U$49701 ( \50078 , \50041 , \50057 );
or \U$49702 ( \50079 , \50077 , \50078 );
and \U$49703 ( \50080 , \50027 , \50079 );
and \U$49704 ( \50081 , \49772 , \50026 );
or \U$49705 ( \50082 , \50080 , \50081 );
xor \U$49706 ( \50083 , \49760 , \50082 );
xor \U$49707 ( \50084 , \49571 , \49596 );
xor \U$49708 ( \50085 , \50084 , \49622 );
xor \U$49709 ( \50086 , \49338 , \49364 );
xor \U$49710 ( \50087 , \50086 , \49367 );
and \U$49711 ( \50088 , \50085 , \50087 );
xor \U$49712 ( \50089 , \49155 , \49162 );
xor \U$49713 ( \50090 , \50089 , \49170 );
xor \U$49714 ( \50091 , \49326 , \49331 );
xor \U$49715 ( \50092 , \50090 , \50091 );
xor \U$49716 ( \50093 , \49338 , \49364 );
xor \U$49717 ( \50094 , \50093 , \49367 );
and \U$49718 ( \50095 , \50092 , \50094 );
and \U$49719 ( \50096 , \50085 , \50092 );
or \U$49720 ( \50097 , \50088 , \50095 , \50096 );
xor \U$49721 ( \50098 , \49093 , \49118 );
xor \U$49722 ( \50099 , \50098 , \49144 );
xor \U$49723 ( \50100 , \50097 , \50099 );
xor \U$49724 ( \50101 , \49014 , \49039 );
xor \U$49725 ( \50102 , \50101 , \49065 );
xor \U$49726 ( \50103 , \49654 , \49659 );
xor \U$49727 ( \50104 , \50102 , \50103 );
and \U$49728 ( \50105 , \50100 , \50104 );
and \U$49729 ( \50106 , \50097 , \50099 );
or \U$49730 ( \50107 , \50105 , \50106 );
and \U$49731 ( \50108 , \50083 , \50107 );
and \U$49732 ( \50109 , \49760 , \50082 );
or \U$49733 ( \50110 , \50108 , \50109 );
xor \U$49734 ( \50111 , \49272 , \49274 );
xor \U$49735 ( \50112 , \50111 , \49289 );
xor \U$49736 ( \50113 , \50110 , \50112 );
xor \U$49737 ( \50114 , \49386 , \49628 );
xor \U$49738 ( \50115 , \50114 , \49645 );
xor \U$49739 ( \50116 , \49652 , \49664 );
xor \U$49740 ( \50117 , \50116 , \49669 );
and \U$49741 ( \50118 , \50115 , \50117 );
xor \U$49742 ( \50119 , \49246 , \49248 );
xor \U$49743 ( \50120 , \50119 , \49253 );
xor \U$49744 ( \50121 , \49675 , \49680 );
xor \U$49745 ( \50122 , \50120 , \50121 );
xor \U$49746 ( \50123 , \49652 , \49664 );
xor \U$49747 ( \50124 , \50123 , \49669 );
and \U$49748 ( \50125 , \50122 , \50124 );
and \U$49749 ( \50126 , \50115 , \50122 );
or \U$49750 ( \50127 , \50118 , \50125 , \50126 );
and \U$49751 ( \50128 , \50113 , \50127 );
and \U$49752 ( \50129 , \50110 , \50112 );
or \U$49753 ( \50130 , \50128 , \50129 );
xor \U$49754 ( \50131 , \49746 , \50130 );
xor \U$49755 ( \50132 , \48403 , \48456 );
xor \U$49756 ( \50133 , \50132 , \48469 );
xor \U$49757 ( \50134 , \49690 , \49697 );
xor \U$49758 ( \50135 , \50133 , \50134 );
xor \U$49759 ( \50136 , \48989 , \49233 );
xor \U$49760 ( \50137 , \50136 , \49256 );
xor \U$49761 ( \50138 , \50135 , \50137 );
xor \U$49762 ( \50139 , \49648 , \49672 );
xor \U$49763 ( \50140 , \50139 , \49685 );
and \U$49764 ( \50141 , \50138 , \50140 );
and \U$49765 ( \50142 , \50135 , \50137 );
or \U$49766 ( \50143 , \50141 , \50142 );
xor \U$49767 ( \50144 , \50131 , \50143 );
not \U$49768 ( \50145 , \50144 );
or \U$49769 ( \50146 , \49744 , \50145 );
or \U$49770 ( \50147 , \50144 , \49743 );
xor \U$49771 ( \50148 , \49772 , \50026 );
xor \U$49772 ( \50149 , \50148 , \50079 );
xor \U$49773 ( \50150 , \50097 , \50099 );
xor \U$49774 ( \50151 , \50150 , \50104 );
and \U$49775 ( \50152 , \50149 , \50151 );
xor \U$49776 ( \50153 , \49336 , \49370 );
xor \U$49777 ( \50154 , \50153 , \49383 );
xor \U$49778 ( \50155 , \49748 , \49755 );
xor \U$49779 ( \50156 , \50154 , \50155 );
xor \U$49780 ( \50157 , \50097 , \50099 );
xor \U$49781 ( \50158 , \50157 , \50104 );
and \U$49782 ( \50159 , \50156 , \50158 );
and \U$49783 ( \50160 , \50149 , \50156 );
or \U$49784 ( \50161 , \50152 , \50159 , \50160 );
xor \U$49785 ( \50162 , \49496 , \49514 );
xor \U$49786 ( \50163 , \50162 , \49540 );
xor \U$49787 ( \50164 , \49762 , \49764 );
xor \U$49788 ( \50165 , \50164 , \49769 );
and \U$49789 ( \50166 , \50163 , \50165 );
xor \U$49790 ( \50167 , \49338 , \49364 );
xor \U$49791 ( \50168 , \50167 , \49367 );
xor \U$49792 ( \50169 , \50085 , \50092 );
xor \U$49793 ( \50170 , \50168 , \50169 );
xor \U$49794 ( \50171 , \49762 , \49764 );
xor \U$49795 ( \50172 , \50171 , \49769 );
and \U$49796 ( \50173 , \50170 , \50172 );
and \U$49797 ( \50174 , \50163 , \50170 );
or \U$49798 ( \50175 , \50166 , \50173 , \50174 );
and \U$49799 ( \50176 , \8966 , RIae75dd0_28);
and \U$49800 ( \50177 , RIae75650_12, \8964 );
nor \U$49801 ( \50178 , \50176 , \50177 );
and \U$49802 ( \50179 , \50178 , \8799 );
not \U$49803 ( \50180 , \50178 );
and \U$49804 ( \50181 , \50180 , \8789 );
nor \U$49805 ( \50182 , \50179 , \50181 );
and \U$49806 ( \50183 , \7633 , RIae75920_18);
and \U$49807 ( \50184 , RIae75fb0_32, \7631 );
nor \U$49808 ( \50185 , \50183 , \50184 );
and \U$49809 ( \50186 , \50185 , \7206 );
not \U$49810 ( \50187 , \50185 );
and \U$49811 ( \50188 , \50187 , \7205 );
nor \U$49812 ( \50189 , \50186 , \50188 );
xor \U$49813 ( \50190 , \50182 , \50189 );
and \U$49814 ( \50191 , \8371 , RIae75ec0_30);
and \U$49815 ( \50192 , RIae75ce0_26, \8369 );
nor \U$49816 ( \50193 , \50191 , \50192 );
and \U$49817 ( \50194 , \50193 , \8020 );
not \U$49818 ( \50195 , \50193 );
and \U$49819 ( \50196 , \50195 , \8019 );
nor \U$49820 ( \50197 , \50194 , \50196 );
and \U$49821 ( \50198 , \50190 , \50197 );
and \U$49822 ( \50199 , \50182 , \50189 );
or \U$49823 ( \50200 , \50198 , \50199 );
and \U$49824 ( \50201 , \4688 , RIae77bd0_92);
and \U$49825 ( \50202 , RIae77db0_96, \4686 );
nor \U$49826 ( \50203 , \50201 , \50202 );
and \U$49827 ( \50204 , \50203 , \4481 );
not \U$49828 ( \50205 , \50203 );
and \U$49829 ( \50206 , \50205 , \4482 );
nor \U$49830 ( \50207 , \50204 , \50206 );
and \U$49831 ( \50208 , \4247 , RIae784b8_111);
and \U$49832 ( \50209 , RIae77cc0_94, \4245 );
nor \U$49833 ( \50210 , \50208 , \50209 );
and \U$49834 ( \50211 , \50210 , \3989 );
not \U$49835 ( \50212 , \50210 );
and \U$49836 ( \50213 , \50212 , \4251 );
nor \U$49837 ( \50214 , \50211 , \50213 );
xor \U$49838 ( \50215 , \50207 , \50214 );
and \U$49839 ( \50216 , \5399 , RIae77ea0_98);
and \U$49840 ( \50217 , RIae789e0_122, \5397 );
nor \U$49841 ( \50218 , \50216 , \50217 );
and \U$49842 ( \50219 , \50218 , \5016 );
not \U$49843 ( \50220 , \50218 );
and \U$49844 ( \50221 , \50220 , \5403 );
nor \U$49845 ( \50222 , \50219 , \50221 );
and \U$49846 ( \50223 , \50215 , \50222 );
and \U$49847 ( \50224 , \50207 , \50214 );
or \U$49848 ( \50225 , \50223 , \50224 );
xor \U$49849 ( \50226 , \50200 , \50225 );
and \U$49850 ( \50227 , \5896 , RIae788f0_120);
and \U$49851 ( \50228 , RIae78800_118, \5894 );
nor \U$49852 ( \50229 , \50227 , \50228 );
and \U$49853 ( \50230 , \50229 , \5590 );
not \U$49854 ( \50231 , \50229 );
and \U$49855 ( \50232 , \50231 , \5589 );
nor \U$49856 ( \50233 , \50230 , \50232 );
and \U$49857 ( \50234 , \6172 , RIae78710_116);
and \U$49858 ( \50235 , RIae75bf0_24, \6170 );
nor \U$49859 ( \50236 , \50234 , \50235 );
and \U$49860 ( \50237 , \50236 , \6176 );
not \U$49861 ( \50238 , \50236 );
and \U$49862 ( \50239 , \50238 , \6175 );
nor \U$49863 ( \50240 , \50237 , \50239 );
xor \U$49864 ( \50241 , \50233 , \50240 );
and \U$49865 ( \50242 , \6941 , RIae75b00_22);
and \U$49866 ( \50243 , RIae75a10_20, \6939 );
nor \U$49867 ( \50244 , \50242 , \50243 );
and \U$49868 ( \50245 , \50244 , \6314 );
not \U$49869 ( \50246 , \50244 );
and \U$49870 ( \50247 , \50246 , \6945 );
nor \U$49871 ( \50248 , \50245 , \50247 );
and \U$49872 ( \50249 , \50241 , \50248 );
and \U$49873 ( \50250 , \50233 , \50240 );
or \U$49874 ( \50251 , \50249 , \50250 );
and \U$49875 ( \50252 , \50226 , \50251 );
and \U$49876 ( \50253 , \50200 , \50225 );
or \U$49877 ( \50254 , \50252 , \50253 );
and \U$49878 ( \50255 , \10548 , RIae75740_14);
and \U$49879 ( \50256 , RIae75290_4, \10546 );
nor \U$49880 ( \50257 , \50255 , \50256 );
and \U$49881 ( \50258 , \50257 , \10421 );
not \U$49882 ( \50259 , \50257 );
and \U$49883 ( \50260 , \50259 , \10118 );
nor \U$49884 ( \50261 , \50258 , \50260 );
and \U$49885 ( \50262 , \9760 , RIae75560_10);
and \U$49886 ( \50263 , RIae75830_16, \9758 );
nor \U$49887 ( \50264 , \50262 , \50263 );
and \U$49888 ( \50265 , \50264 , \9273 );
not \U$49889 ( \50266 , \50264 );
and \U$49890 ( \50267 , \50266 , \9272 );
nor \U$49891 ( \50268 , \50265 , \50267 );
xor \U$49892 ( \50269 , \50261 , \50268 );
and \U$49893 ( \50270 , \11470 , RIae751a0_2);
and \U$49894 ( \50271 , RIae75380_6, \11468 );
nor \U$49895 ( \50272 , \50270 , \50271 );
and \U$49896 ( \50273 , \50272 , \10936 );
not \U$49897 ( \50274 , \50272 );
and \U$49898 ( \50275 , \50274 , \11474 );
nor \U$49899 ( \50276 , \50273 , \50275 );
and \U$49900 ( \50277 , \50269 , \50276 );
and \U$49901 ( \50278 , \50261 , \50268 );
or \U$49902 ( \50279 , \50277 , \50278 );
and \U$49903 ( \50280 , \15726 , RIae76280_38);
and \U$49904 ( \50281 , RIae76af0_56, RIae7aab0_192);
nor \U$49905 ( \50282 , \50280 , \50281 );
and \U$49906 ( \50283 , \50282 , \14959 );
not \U$49907 ( \50284 , \50282 );
and \U$49908 ( \50285 , \50284 , RIae7aa38_191);
nor \U$49909 ( \50286 , \50283 , \50285 );
xor \U$49910 ( \50287 , \50286 , \562 );
and \U$49911 ( \50288 , \14964 , RIae760a0_34);
and \U$49912 ( \50289 , RIae76370_40, \14962 );
nor \U$49913 ( \50290 , \50288 , \50289 );
and \U$49914 ( \50291 , \50290 , \14463 );
not \U$49915 ( \50292 , \50290 );
and \U$49916 ( \50293 , \50292 , \14462 );
nor \U$49917 ( \50294 , \50291 , \50293 );
and \U$49918 ( \50295 , \50287 , \50294 );
and \U$49919 ( \50296 , \50286 , \562 );
or \U$49920 ( \50297 , \50295 , \50296 );
xor \U$49921 ( \50298 , \50279 , \50297 );
and \U$49922 ( \50299 , \14059 , RIae76640_46);
and \U$49923 ( \50300 , RIae76190_36, \14057 );
nor \U$49924 ( \50301 , \50299 , \50300 );
and \U$49925 ( \50302 , \50301 , \13502 );
not \U$49926 ( \50303 , \50301 );
and \U$49927 ( \50304 , \50303 , \14063 );
nor \U$49928 ( \50305 , \50302 , \50304 );
and \U$49929 ( \50306 , \12180 , RIae75470_8);
and \U$49930 ( \50307 , RIae76460_42, \12178 );
nor \U$49931 ( \50308 , \50306 , \50307 );
and \U$49932 ( \50309 , \50308 , \12184 );
not \U$49933 ( \50310 , \50308 );
and \U$49934 ( \50311 , \50310 , \11827 );
nor \U$49935 ( \50312 , \50309 , \50311 );
xor \U$49936 ( \50313 , \50305 , \50312 );
and \U$49937 ( \50314 , \13059 , RIae76550_44);
and \U$49938 ( \50315 , RIae76730_48, \13057 );
nor \U$49939 ( \50316 , \50314 , \50315 );
and \U$49940 ( \50317 , \50316 , \13063 );
not \U$49941 ( \50318 , \50316 );
and \U$49942 ( \50319 , \50318 , \12718 );
nor \U$49943 ( \50320 , \50317 , \50319 );
and \U$49944 ( \50321 , \50313 , \50320 );
and \U$49945 ( \50322 , \50305 , \50312 );
or \U$49946 ( \50323 , \50321 , \50322 );
and \U$49947 ( \50324 , \50298 , \50323 );
and \U$49948 ( \50325 , \50279 , \50297 );
or \U$49949 ( \50326 , \50324 , \50325 );
xor \U$49950 ( \50327 , \50254 , \50326 );
and \U$49951 ( \50328 , \2607 , RIae77360_74);
and \U$49952 ( \50329 , RIae78350_108, \2605 );
nor \U$49953 ( \50330 , \50328 , \50329 );
and \U$49954 ( \50331 , \50330 , \2611 );
not \U$49955 ( \50332 , \50330 );
and \U$49956 ( \50333 , \50332 , \2397 );
nor \U$49957 ( \50334 , \50331 , \50333 );
and \U$49958 ( \50335 , \1939 , RIae76cd0_60);
and \U$49959 ( \50336 , RIae77108_69, \1937 );
nor \U$49960 ( \50337 , \50335 , \50336 );
and \U$49961 ( \50338 , \50337 , \1735 );
not \U$49962 ( \50339 , \50337 );
and \U$49963 ( \50340 , \50339 , \1734 );
nor \U$49964 ( \50341 , \50338 , \50340 );
xor \U$49965 ( \50342 , \50334 , \50341 );
and \U$49966 ( \50343 , \2224 , RIae77090_68);
and \U$49967 ( \50344 , RIae77270_72, \2222 );
nor \U$49968 ( \50345 , \50343 , \50344 );
and \U$49969 ( \50346 , \50345 , \2061 );
not \U$49970 ( \50347 , \50345 );
and \U$49971 ( \50348 , \50347 , \2060 );
nor \U$49972 ( \50349 , \50346 , \50348 );
and \U$49973 ( \50350 , \50342 , \50349 );
and \U$49974 ( \50351 , \50334 , \50341 );
or \U$49975 ( \50352 , \50350 , \50351 );
and \U$49976 ( \50353 , \1138 , RIae779f0_88);
and \U$49977 ( \50354 , RIae77810_84, \1136 );
nor \U$49978 ( \50355 , \50353 , \50354 );
and \U$49979 ( \50356 , \50355 , \1142 );
not \U$49980 ( \50357 , \50355 );
and \U$49981 ( \50358 , \50357 , \1012 );
nor \U$49982 ( \50359 , \50356 , \50358 );
and \U$49983 ( \50360 , \1376 , RIae77900_86);
and \U$49984 ( \50361 , RIae76fa0_66, \1374 );
nor \U$49985 ( \50362 , \50360 , \50361 );
and \U$49986 ( \50363 , \50362 , \1261 );
not \U$49987 ( \50364 , \50362 );
and \U$49988 ( \50365 , \50364 , \1380 );
nor \U$49989 ( \50366 , \50363 , \50365 );
or \U$49990 ( \50367 , \50359 , \50366 );
not \U$49991 ( \50368 , \50366 );
not \U$49992 ( \50369 , \50359 );
or \U$49993 ( \50370 , \50368 , \50369 );
and \U$49994 ( \50371 , \1593 , RIae76eb0_64);
and \U$49995 ( \50372 , RIae76dc0_62, \1591 );
nor \U$49996 ( \50373 , \50371 , \50372 );
and \U$49997 ( \50374 , \50373 , \1498 );
not \U$49998 ( \50375 , \50373 );
and \U$49999 ( \50376 , \50375 , \1488 );
nor \U$50000 ( \50377 , \50374 , \50376 );
nand \U$50001 ( \50378 , \50370 , \50377 );
nand \U$50002 ( \50379 , \50367 , \50378 );
xor \U$50003 ( \50380 , \50352 , \50379 );
and \U$50004 ( \50381 , \3730 , RIae78620_114);
and \U$50005 ( \50382 , RIae78440_110, \3728 );
nor \U$50006 ( \50383 , \50381 , \50382 );
and \U$50007 ( \50384 , \50383 , \3732 );
not \U$50008 ( \50385 , \50383 );
and \U$50009 ( \50386 , \50385 , \3422 );
nor \U$50010 ( \50387 , \50384 , \50386 );
not \U$50011 ( \50388 , \2789 );
and \U$50012 ( \50389 , \2783 , RIae78170_104);
and \U$50013 ( \50390 , RIae77f90_100, \2781 );
nor \U$50014 ( \50391 , \50389 , \50390 );
not \U$50015 ( \50392 , \50391 );
or \U$50016 ( \50393 , \50388 , \50392 );
or \U$50017 ( \50394 , \50391 , \2789 );
nand \U$50018 ( \50395 , \50393 , \50394 );
xor \U$50019 ( \50396 , \50387 , \50395 );
not \U$50020 ( \50397 , \3218 );
and \U$50021 ( \50398 , \3214 , RIae78080_102);
and \U$50022 ( \50399 , RIae78260_106, \3212 );
nor \U$50023 ( \50400 , \50398 , \50399 );
not \U$50024 ( \50401 , \50400 );
or \U$50025 ( \50402 , \50397 , \50401 );
or \U$50026 ( \50403 , \50400 , \2774 );
nand \U$50027 ( \50404 , \50402 , \50403 );
and \U$50028 ( \50405 , \50396 , \50404 );
and \U$50029 ( \50406 , \50387 , \50395 );
or \U$50030 ( \50407 , \50405 , \50406 );
and \U$50031 ( \50408 , \50380 , \50407 );
and \U$50032 ( \50409 , \50352 , \50379 );
or \U$50033 ( \50410 , \50408 , \50409 );
and \U$50034 ( \50411 , \50327 , \50410 );
and \U$50035 ( \50412 , \50254 , \50326 );
or \U$50036 ( \50413 , \50411 , \50412 );
xor \U$50037 ( \50414 , \49503 , \469 );
xor \U$50038 ( \50415 , \50414 , \49511 );
xor \U$50039 ( \50416 , \49522 , \49529 );
xor \U$50040 ( \50417 , \50416 , \49537 );
and \U$50041 ( \50418 , \50415 , \50417 );
xor \U$50042 ( \50419 , \49947 , \49954 );
xor \U$50043 ( \50420 , \50419 , \49962 );
xor \U$50044 ( \50421 , \50003 , \50010 );
xor \U$50045 ( \50422 , \50421 , \50018 );
and \U$50046 ( \50423 , \50420 , \50422 );
not \U$50047 ( \50424 , \49972 );
xor \U$50048 ( \50425 , \49990 , \49980 );
not \U$50049 ( \50426 , \50425 );
or \U$50050 ( \50427 , \50424 , \50426 );
or \U$50051 ( \50428 , \50425 , \49972 );
nand \U$50052 ( \50429 , \50427 , \50428 );
xor \U$50053 ( \50430 , \50003 , \50010 );
xor \U$50054 ( \50431 , \50430 , \50018 );
and \U$50055 ( \50432 , \50429 , \50431 );
and \U$50056 ( \50433 , \50420 , \50429 );
or \U$50057 ( \50434 , \50423 , \50432 , \50433 );
xor \U$50058 ( \50435 , \49522 , \49529 );
xor \U$50059 ( \50436 , \50435 , \49537 );
and \U$50060 ( \50437 , \50434 , \50436 );
and \U$50061 ( \50438 , \50415 , \50434 );
or \U$50062 ( \50439 , \50418 , \50437 , \50438 );
xor \U$50063 ( \50440 , \50413 , \50439 );
xor \U$50064 ( \50441 , \49888 , \49895 );
xor \U$50065 ( \50442 , \50441 , \49903 );
xor \U$50066 ( \50443 , \49862 , \49869 );
xor \U$50067 ( \50444 , \50443 , \49878 );
xor \U$50068 ( \50445 , \50442 , \50444 );
not \U$50069 ( \50446 , \49914 );
xor \U$50070 ( \50447 , \49923 , \49934 );
not \U$50071 ( \50448 , \50447 );
or \U$50072 ( \50449 , \50446 , \50448 );
or \U$50073 ( \50450 , \50447 , \49914 );
nand \U$50074 ( \50451 , \50449 , \50450 );
and \U$50075 ( \50452 , \50445 , \50451 );
and \U$50076 ( \50453 , \50442 , \50444 );
or \U$50077 ( \50454 , \50452 , \50453 );
and \U$50078 ( \50455 , \672 , RIae776a8_81);
and \U$50079 ( \50456 , RIae77450_76, \670 );
nor \U$50080 ( \50457 , \50455 , \50456 );
and \U$50081 ( \50458 , \50457 , \588 );
not \U$50082 ( \50459 , \50457 );
and \U$50083 ( \50460 , \50459 , \587 );
nor \U$50084 ( \50461 , \50458 , \50460 );
and \U$50085 ( \50462 , \558 , RIae77630_80);
and \U$50086 ( \50463 , RIae77540_78, \556 );
nor \U$50087 ( \50464 , \50462 , \50463 );
and \U$50088 ( \50465 , \50464 , \504 );
not \U$50089 ( \50466 , \50464 );
and \U$50090 ( \50467 , \50466 , \562 );
nor \U$50091 ( \50468 , \50465 , \50467 );
xor \U$50092 ( \50469 , \50461 , \50468 );
nand \U$50093 ( \50470 , RIae77630_80, \556 );
and \U$50094 ( \50471 , \50470 , \504 );
not \U$50095 ( \50472 , \50470 );
and \U$50096 ( \50473 , \50472 , \562 );
nor \U$50097 ( \50474 , \50471 , \50473 );
not \U$50098 ( \50475 , \50474 );
and \U$50099 ( \50476 , \672 , RIae77540_78);
and \U$50100 ( \50477 , RIae776a8_81, \670 );
nor \U$50101 ( \50478 , \50476 , \50477 );
and \U$50102 ( \50479 , \50478 , \588 );
not \U$50103 ( \50480 , \50478 );
and \U$50104 ( \50481 , \50480 , \587 );
nor \U$50105 ( \50482 , \50479 , \50481 );
not \U$50106 ( \50483 , \50482 );
or \U$50107 ( \50484 , \50475 , \50483 );
or \U$50108 ( \50485 , \50482 , \50474 );
not \U$50109 ( \50486 , \787 );
and \U$50110 ( \50487 , \883 , RIae77450_76);
and \U$50111 ( \50488 , RIae77ae0_90, \881 );
nor \U$50112 ( \50489 , \50487 , \50488 );
not \U$50113 ( \50490 , \50489 );
or \U$50114 ( \50491 , \50486 , \50490 );
or \U$50115 ( \50492 , \50489 , \787 );
nand \U$50116 ( \50493 , \50491 , \50492 );
nand \U$50117 ( \50494 , \50485 , \50493 );
nand \U$50118 ( \50495 , \50484 , \50494 );
and \U$50119 ( \50496 , \50469 , \50495 );
and \U$50120 ( \50497 , \50461 , \50468 );
or \U$50121 ( \50498 , \50496 , \50497 );
xor \U$50122 ( \50499 , \50454 , \50498 );
xor \U$50123 ( \50500 , \49806 , \49813 );
xor \U$50124 ( \50501 , \50500 , \49821 );
not \U$50125 ( \50502 , \49779 );
xor \U$50126 ( \50503 , \49787 , \49797 );
not \U$50127 ( \50504 , \50503 );
or \U$50128 ( \50505 , \50502 , \50504 );
or \U$50129 ( \50506 , \50503 , \49779 );
nand \U$50130 ( \50507 , \50505 , \50506 );
xor \U$50131 ( \50508 , \50501 , \50507 );
not \U$50132 ( \50509 , \49832 );
xor \U$50133 ( \50510 , \49840 , \49850 );
not \U$50134 ( \50511 , \50510 );
or \U$50135 ( \50512 , \50509 , \50511 );
or \U$50136 ( \50513 , \50510 , \49832 );
nand \U$50137 ( \50514 , \50512 , \50513 );
and \U$50138 ( \50515 , \50508 , \50514 );
and \U$50139 ( \50516 , \50501 , \50507 );
or \U$50140 ( \50517 , \50515 , \50516 );
and \U$50141 ( \50518 , \50499 , \50517 );
and \U$50142 ( \50519 , \50454 , \50498 );
or \U$50143 ( \50520 , \50518 , \50519 );
and \U$50144 ( \50521 , \50440 , \50520 );
and \U$50145 ( \50522 , \50413 , \50439 );
or \U$50146 ( \50523 , \50521 , \50522 );
xor \U$50147 ( \50524 , \50175 , \50523 );
not \U$50148 ( \50525 , \50021 );
not \U$50149 ( \50526 , \49992 );
or \U$50150 ( \50527 , \50525 , \50526 );
or \U$50151 ( \50528 , \49992 , \50021 );
nand \U$50152 ( \50529 , \50527 , \50528 );
not \U$50153 ( \50530 , \50529 );
not \U$50154 ( \50531 , \49965 );
and \U$50155 ( \50532 , \50530 , \50531 );
and \U$50156 ( \50533 , \50529 , \49965 );
nor \U$50157 ( \50534 , \50532 , \50533 );
not \U$50158 ( \50535 , \50534 );
xor \U$50159 ( \50536 , \49881 , \49906 );
xor \U$50160 ( \50537 , \50536 , \49936 );
not \U$50161 ( \50538 , \50537 );
and \U$50162 ( \50539 , \50535 , \50538 );
and \U$50163 ( \50540 , \50534 , \50537 );
xor \U$50164 ( \50541 , \49799 , \49824 );
xor \U$50165 ( \50542 , \50541 , \49852 );
nor \U$50166 ( \50543 , \50540 , \50542 );
nor \U$50167 ( \50544 , \50539 , \50543 );
xor \U$50168 ( \50545 , \49413 , \49440 );
xor \U$50169 ( \50546 , \50545 , \49468 );
or \U$50170 ( \50547 , \50544 , \50546 );
not \U$50171 ( \50548 , \50546 );
not \U$50172 ( \50549 , \50544 );
or \U$50173 ( \50550 , \50548 , \50549 );
xor \U$50174 ( \50551 , \49604 , \49611 );
xor \U$50175 ( \50552 , \50551 , \49619 );
xor \U$50176 ( \50553 , \50047 , \50052 );
xor \U$50177 ( \50554 , \50552 , \50553 );
xor \U$50178 ( \50555 , \50029 , \50031 );
xor \U$50179 ( \50556 , \50555 , \50038 );
and \U$50180 ( \50557 , \50554 , \50556 );
xor \U$50181 ( \50558 , \50064 , \50070 );
xor \U$50182 ( \50559 , \50558 , \50073 );
xor \U$50183 ( \50560 , \50029 , \50031 );
xor \U$50184 ( \50561 , \50560 , \50038 );
and \U$50185 ( \50562 , \50559 , \50561 );
and \U$50186 ( \50563 , \50554 , \50559 );
or \U$50187 ( \50564 , \50557 , \50562 , \50563 );
nand \U$50188 ( \50565 , \50550 , \50564 );
nand \U$50189 ( \50566 , \50547 , \50565 );
and \U$50190 ( \50567 , \50524 , \50566 );
and \U$50191 ( \50568 , \50175 , \50523 );
or \U$50192 ( \50569 , \50567 , \50568 );
xor \U$50193 ( \50570 , \50161 , \50569 );
xor \U$50194 ( \50571 , \49652 , \49664 );
xor \U$50195 ( \50572 , \50571 , \49669 );
xor \U$50196 ( \50573 , \50115 , \50122 );
xor \U$50197 ( \50574 , \50572 , \50573 );
and \U$50198 ( \50575 , \50570 , \50574 );
and \U$50199 ( \50576 , \50161 , \50569 );
or \U$50200 ( \50577 , \50575 , \50576 );
xor \U$50201 ( \50578 , \50135 , \50137 );
xor \U$50202 ( \50579 , \50578 , \50140 );
and \U$50203 ( \50580 , \50577 , \50579 );
xor \U$50204 ( \50581 , \50110 , \50112 );
xor \U$50205 ( \50582 , \50581 , \50127 );
xor \U$50206 ( \50583 , \50135 , \50137 );
xor \U$50207 ( \50584 , \50583 , \50140 );
and \U$50208 ( \50585 , \50582 , \50584 );
and \U$50209 ( \50586 , \50577 , \50582 );
or \U$50210 ( \50587 , \50580 , \50585 , \50586 );
nand \U$50211 ( \50588 , \50147 , \50587 );
nand \U$50212 ( \50589 , \50146 , \50588 );
xor \U$50213 ( \50590 , \49746 , \50130 );
and \U$50214 ( \50591 , \50590 , \50143 );
and \U$50215 ( \50592 , \49746 , \50130 );
nor \U$50216 ( \50593 , \50591 , \50592 );
not \U$50217 ( \50594 , \50593 );
xor \U$50218 ( \50595 , \49324 , \49710 );
xor \U$50219 ( \50596 , \50595 , \49721 );
not \U$50220 ( \50597 , \50596 );
or \U$50221 ( \50598 , \50594 , \50597 );
or \U$50222 ( \50599 , \50596 , \50593 );
nand \U$50223 ( \50600 , \50598 , \50599 );
and \U$50224 ( \50601 , \50589 , \50600 );
xor \U$50225 ( \50602 , \50600 , \50589 );
xnor \U$50226 ( \50603 , \50587 , \50144 );
not \U$50227 ( \50604 , \50603 );
not \U$50228 ( \50605 , \49743 );
and \U$50229 ( \50606 , \50604 , \50605 );
and \U$50230 ( \50607 , \50603 , \49743 );
nor \U$50231 ( \50608 , \50606 , \50607 );
xor \U$50232 ( \50609 , \50161 , \50569 );
xor \U$50233 ( \50610 , \50609 , \50574 );
xor \U$50234 ( \50611 , \50254 , \50326 );
xor \U$50235 ( \50612 , \50611 , \50410 );
xor \U$50236 ( \50613 , \50454 , \50498 );
xor \U$50237 ( \50614 , \50613 , \50517 );
and \U$50238 ( \50615 , \50612 , \50614 );
xor \U$50239 ( \50616 , \49522 , \49529 );
xor \U$50240 ( \50617 , \50616 , \49537 );
xor \U$50241 ( \50618 , \50415 , \50434 );
xor \U$50242 ( \50619 , \50617 , \50618 );
xor \U$50243 ( \50620 , \50454 , \50498 );
xor \U$50244 ( \50621 , \50620 , \50517 );
and \U$50245 ( \50622 , \50619 , \50621 );
and \U$50246 ( \50623 , \50612 , \50619 );
or \U$50247 ( \50624 , \50615 , \50622 , \50623 );
xnor \U$50248 ( \50625 , \50493 , \50482 );
not \U$50249 ( \50626 , \50625 );
not \U$50250 ( \50627 , \50474 );
and \U$50251 ( \50628 , \50626 , \50627 );
and \U$50252 ( \50629 , \50625 , \50474 );
nor \U$50253 ( \50630 , \50628 , \50629 );
not \U$50254 ( \50631 , \50366 );
not \U$50255 ( \50632 , \50377 );
or \U$50256 ( \50633 , \50631 , \50632 );
or \U$50257 ( \50634 , \50366 , \50377 );
nand \U$50258 ( \50635 , \50633 , \50634 );
not \U$50259 ( \50636 , \50635 );
not \U$50260 ( \50637 , \50359 );
and \U$50261 ( \50638 , \50636 , \50637 );
and \U$50262 ( \50639 , \50635 , \50359 );
nor \U$50263 ( \50640 , \50638 , \50639 );
or \U$50264 ( \50641 , \50630 , \50640 );
not \U$50265 ( \50642 , \50640 );
not \U$50266 ( \50643 , \50630 );
or \U$50267 ( \50644 , \50642 , \50643 );
xor \U$50268 ( \50645 , \50334 , \50341 );
xor \U$50269 ( \50646 , \50645 , \50349 );
nand \U$50270 ( \50647 , \50644 , \50646 );
nand \U$50271 ( \50648 , \50641 , \50647 );
xor \U$50272 ( \50649 , \50387 , \50395 );
xor \U$50273 ( \50650 , \50649 , \50404 );
xor \U$50274 ( \50651 , \50233 , \50240 );
xor \U$50275 ( \50652 , \50651 , \50248 );
and \U$50276 ( \50653 , \50650 , \50652 );
xor \U$50277 ( \50654 , \50207 , \50214 );
xor \U$50278 ( \50655 , \50654 , \50222 );
xor \U$50279 ( \50656 , \50233 , \50240 );
xor \U$50280 ( \50657 , \50656 , \50248 );
and \U$50281 ( \50658 , \50655 , \50657 );
and \U$50282 ( \50659 , \50650 , \50655 );
or \U$50283 ( \50660 , \50653 , \50658 , \50659 );
xor \U$50284 ( \50661 , \50648 , \50660 );
xor \U$50285 ( \50662 , \50261 , \50268 );
xor \U$50286 ( \50663 , \50662 , \50276 );
xor \U$50287 ( \50664 , \50182 , \50189 );
xor \U$50288 ( \50665 , \50664 , \50197 );
xor \U$50289 ( \50666 , \50663 , \50665 );
xor \U$50290 ( \50667 , \50305 , \50312 );
xor \U$50291 ( \50668 , \50667 , \50320 );
and \U$50292 ( \50669 , \50666 , \50668 );
and \U$50293 ( \50670 , \50663 , \50665 );
or \U$50294 ( \50671 , \50669 , \50670 );
and \U$50295 ( \50672 , \50661 , \50671 );
and \U$50296 ( \50673 , \50648 , \50660 );
or \U$50297 ( \50674 , \50672 , \50673 );
and \U$50298 ( \50675 , \4688 , RIae77cc0_94);
and \U$50299 ( \50676 , RIae77bd0_92, \4686 );
nor \U$50300 ( \50677 , \50675 , \50676 );
and \U$50301 ( \50678 , \50677 , \4482 );
not \U$50302 ( \50679 , \50677 );
and \U$50303 ( \50680 , \50679 , \4481 );
nor \U$50304 ( \50681 , \50678 , \50680 );
and \U$50305 ( \50682 , \3730 , RIae78260_106);
and \U$50306 ( \50683 , RIae78620_114, \3728 );
nor \U$50307 ( \50684 , \50682 , \50683 );
and \U$50308 ( \50685 , \50684 , \3422 );
not \U$50309 ( \50686 , \50684 );
and \U$50310 ( \50687 , \50686 , \3732 );
nor \U$50311 ( \50688 , \50685 , \50687 );
xor \U$50312 ( \50689 , \50681 , \50688 );
and \U$50313 ( \50690 , \4247 , RIae78440_110);
and \U$50314 ( \50691 , RIae784b8_111, \4245 );
nor \U$50315 ( \50692 , \50690 , \50691 );
and \U$50316 ( \50693 , \50692 , \4251 );
not \U$50317 ( \50694 , \50692 );
and \U$50318 ( \50695 , \50694 , \3989 );
nor \U$50319 ( \50696 , \50693 , \50695 );
and \U$50320 ( \50697 , \50689 , \50696 );
and \U$50321 ( \50698 , \50681 , \50688 );
or \U$50322 ( \50699 , \50697 , \50698 );
and \U$50323 ( \50700 , \8371 , RIae75fb0_32);
and \U$50324 ( \50701 , RIae75ec0_30, \8369 );
nor \U$50325 ( \50702 , \50700 , \50701 );
and \U$50326 ( \50703 , \50702 , \8019 );
not \U$50327 ( \50704 , \50702 );
and \U$50328 ( \50705 , \50704 , \8020 );
nor \U$50329 ( \50706 , \50703 , \50705 );
and \U$50330 ( \50707 , \6941 , RIae75bf0_24);
and \U$50331 ( \50708 , RIae75b00_22, \6939 );
nor \U$50332 ( \50709 , \50707 , \50708 );
and \U$50333 ( \50710 , \50709 , \6945 );
not \U$50334 ( \50711 , \50709 );
and \U$50335 ( \50712 , \50711 , \6314 );
nor \U$50336 ( \50713 , \50710 , \50712 );
xor \U$50337 ( \50714 , \50706 , \50713 );
and \U$50338 ( \50715 , \7633 , RIae75a10_20);
and \U$50339 ( \50716 , RIae75920_18, \7631 );
nor \U$50340 ( \50717 , \50715 , \50716 );
and \U$50341 ( \50718 , \50717 , \7205 );
not \U$50342 ( \50719 , \50717 );
and \U$50343 ( \50720 , \50719 , \7206 );
nor \U$50344 ( \50721 , \50718 , \50720 );
and \U$50345 ( \50722 , \50714 , \50721 );
and \U$50346 ( \50723 , \50706 , \50713 );
or \U$50347 ( \50724 , \50722 , \50723 );
xor \U$50348 ( \50725 , \50699 , \50724 );
and \U$50349 ( \50726 , \5896 , RIae789e0_122);
and \U$50350 ( \50727 , RIae788f0_120, \5894 );
nor \U$50351 ( \50728 , \50726 , \50727 );
and \U$50352 ( \50729 , \50728 , \5590 );
not \U$50353 ( \50730 , \50728 );
and \U$50354 ( \50731 , \50730 , \5589 );
nor \U$50355 ( \50732 , \50729 , \50731 );
and \U$50356 ( \50733 , \6172 , RIae78800_118);
and \U$50357 ( \50734 , RIae78710_116, \6170 );
nor \U$50358 ( \50735 , \50733 , \50734 );
and \U$50359 ( \50736 , \50735 , \6176 );
not \U$50360 ( \50737 , \50735 );
and \U$50361 ( \50738 , \50737 , \6175 );
nor \U$50362 ( \50739 , \50736 , \50738 );
xor \U$50363 ( \50740 , \50732 , \50739 );
and \U$50364 ( \50741 , \5399 , RIae77db0_96);
and \U$50365 ( \50742 , RIae77ea0_98, \5397 );
nor \U$50366 ( \50743 , \50741 , \50742 );
and \U$50367 ( \50744 , \50743 , \5016 );
not \U$50368 ( \50745 , \50743 );
and \U$50369 ( \50746 , \50745 , \5403 );
nor \U$50370 ( \50747 , \50744 , \50746 );
and \U$50371 ( \50748 , \50740 , \50747 );
and \U$50372 ( \50749 , \50732 , \50739 );
nor \U$50373 ( \50750 , \50748 , \50749 );
and \U$50374 ( \50751 , \50725 , \50750 );
and \U$50375 ( \50752 , \50699 , \50724 );
nor \U$50376 ( \50753 , \50751 , \50752 );
and \U$50377 ( \50754 , \14964 , RIae76190_36);
and \U$50378 ( \50755 , RIae760a0_34, \14962 );
nor \U$50379 ( \50756 , \50754 , \50755 );
and \U$50380 ( \50757 , \50756 , \14462 );
not \U$50381 ( \50758 , \50756 );
and \U$50382 ( \50759 , \50758 , \14463 );
nor \U$50383 ( \50760 , \50757 , \50759 );
and \U$50384 ( \50761 , \15726 , RIae76370_40);
and \U$50385 ( \50762 , RIae76280_38, RIae7aab0_192);
nor \U$50386 ( \50763 , \50761 , \50762 );
and \U$50387 ( \50764 , \50763 , RIae7aa38_191);
not \U$50388 ( \50765 , \50763 );
and \U$50389 ( \50766 , \50765 , \14959 );
nor \U$50390 ( \50767 , \50764 , \50766 );
xor \U$50391 ( \50768 , \50760 , \50767 );
and \U$50392 ( \50769 , \14059 , RIae76730_48);
and \U$50393 ( \50770 , RIae76640_46, \14057 );
nor \U$50394 ( \50771 , \50769 , \50770 );
and \U$50395 ( \50772 , \50771 , \14063 );
not \U$50396 ( \50773 , \50771 );
and \U$50397 ( \50774 , \50773 , \13502 );
nor \U$50398 ( \50775 , \50772 , \50774 );
and \U$50399 ( \50776 , \50768 , \50775 );
and \U$50400 ( \50777 , \50760 , \50767 );
or \U$50401 ( \50778 , \50776 , \50777 );
and \U$50402 ( \50779 , \8966 , RIae75ce0_26);
and \U$50403 ( \50780 , RIae75dd0_28, \8964 );
nor \U$50404 ( \50781 , \50779 , \50780 );
and \U$50405 ( \50782 , \50781 , \8789 );
not \U$50406 ( \50783 , \50781 );
and \U$50407 ( \50784 , \50783 , \8799 );
nor \U$50408 ( \50785 , \50782 , \50784 );
not \U$50409 ( \50786 , \50785 );
and \U$50410 ( \50787 , \10548 , RIae75830_16);
and \U$50411 ( \50788 , RIae75740_14, \10546 );
nor \U$50412 ( \50789 , \50787 , \50788 );
and \U$50413 ( \50790 , \50789 , \10118 );
not \U$50414 ( \50791 , \50789 );
and \U$50415 ( \50792 , \50791 , \10421 );
nor \U$50416 ( \50793 , \50790 , \50792 );
not \U$50417 ( \50794 , \50793 );
and \U$50418 ( \50795 , \50786 , \50794 );
and \U$50419 ( \50796 , \50793 , \50785 );
and \U$50420 ( \50797 , \9760 , RIae75650_12);
and \U$50421 ( \50798 , RIae75560_10, \9758 );
nor \U$50422 ( \50799 , \50797 , \50798 );
and \U$50423 ( \50800 , \50799 , \9272 );
not \U$50424 ( \50801 , \50799 );
and \U$50425 ( \50802 , \50801 , \9273 );
nor \U$50426 ( \50803 , \50800 , \50802 );
nor \U$50427 ( \50804 , \50796 , \50803 );
nor \U$50428 ( \50805 , \50795 , \50804 );
xor \U$50429 ( \50806 , \50778 , \50805 );
and \U$50430 ( \50807 , \11470 , RIae75290_4);
and \U$50431 ( \50808 , RIae751a0_2, \11468 );
nor \U$50432 ( \50809 , \50807 , \50808 );
and \U$50433 ( \50810 , \50809 , \11474 );
not \U$50434 ( \50811 , \50809 );
and \U$50435 ( \50812 , \50811 , \10936 );
nor \U$50436 ( \50813 , \50810 , \50812 );
and \U$50437 ( \50814 , \12180 , RIae75380_6);
and \U$50438 ( \50815 , RIae75470_8, \12178 );
nor \U$50439 ( \50816 , \50814 , \50815 );
and \U$50440 ( \50817 , \50816 , \11827 );
not \U$50441 ( \50818 , \50816 );
and \U$50442 ( \50819 , \50818 , \12184 );
nor \U$50443 ( \50820 , \50817 , \50819 );
xor \U$50444 ( \50821 , \50813 , \50820 );
and \U$50445 ( \50822 , \13059 , RIae76460_42);
and \U$50446 ( \50823 , RIae76550_44, \13057 );
nor \U$50447 ( \50824 , \50822 , \50823 );
and \U$50448 ( \50825 , \50824 , \12718 );
not \U$50449 ( \50826 , \50824 );
and \U$50450 ( \50827 , \50826 , \13063 );
nor \U$50451 ( \50828 , \50825 , \50827 );
and \U$50452 ( \50829 , \50821 , \50828 );
and \U$50453 ( \50830 , \50813 , \50820 );
or \U$50454 ( \50831 , \50829 , \50830 );
and \U$50455 ( \50832 , \50806 , \50831 );
and \U$50456 ( \50833 , \50778 , \50805 );
nor \U$50457 ( \50834 , \50832 , \50833 );
xor \U$50458 ( \50835 , \50753 , \50834 );
and \U$50459 ( \50836 , \883 , RIae776a8_81);
and \U$50460 ( \50837 , RIae77450_76, \881 );
nor \U$50461 ( \50838 , \50836 , \50837 );
not \U$50462 ( \50839 , \50838 );
not \U$50463 ( \50840 , \789 );
and \U$50464 ( \50841 , \50839 , \50840 );
and \U$50465 ( \50842 , \50838 , \789 );
nor \U$50466 ( \50843 , \50841 , \50842 );
and \U$50467 ( \50844 , \1138 , RIae77ae0_90);
and \U$50468 ( \50845 , RIae779f0_88, \1136 );
nor \U$50469 ( \50846 , \50844 , \50845 );
and \U$50470 ( \50847 , \50846 , \1142 );
not \U$50471 ( \50848 , \50846 );
and \U$50472 ( \50849 , \50848 , \1012 );
nor \U$50473 ( \50850 , \50847 , \50849 );
xor \U$50474 ( \50851 , \50843 , \50850 );
and \U$50475 ( \50852 , \1376 , RIae77810_84);
and \U$50476 ( \50853 , RIae77900_86, \1374 );
nor \U$50477 ( \50854 , \50852 , \50853 );
and \U$50478 ( \50855 , \50854 , \1261 );
not \U$50479 ( \50856 , \50854 );
and \U$50480 ( \50857 , \50856 , \1380 );
nor \U$50481 ( \50858 , \50855 , \50857 );
and \U$50482 ( \50859 , \50851 , \50858 );
and \U$50483 ( \50860 , \50843 , \50850 );
or \U$50484 ( \50861 , \50859 , \50860 );
and \U$50485 ( \50862 , \2783 , RIae78350_108);
and \U$50486 ( \50863 , RIae78170_104, \2781 );
nor \U$50487 ( \50864 , \50862 , \50863 );
not \U$50488 ( \50865 , \50864 );
not \U$50489 ( \50866 , \2789 );
and \U$50490 ( \50867 , \50865 , \50866 );
and \U$50491 ( \50868 , \50864 , \2789 );
nor \U$50492 ( \50869 , \50867 , \50868 );
and \U$50493 ( \50870 , \2607 , RIae77270_72);
and \U$50494 ( \50871 , RIae77360_74, \2605 );
nor \U$50495 ( \50872 , \50870 , \50871 );
and \U$50496 ( \50873 , \50872 , \2397 );
not \U$50497 ( \50874 , \50872 );
and \U$50498 ( \50875 , \50874 , \2611 );
nor \U$50499 ( \50876 , \50873 , \50875 );
xor \U$50500 ( \50877 , \50869 , \50876 );
and \U$50501 ( \50878 , \3214 , RIae77f90_100);
and \U$50502 ( \50879 , RIae78080_102, \3212 );
nor \U$50503 ( \50880 , \50878 , \50879 );
not \U$50504 ( \50881 , \50880 );
not \U$50505 ( \50882 , \2774 );
and \U$50506 ( \50883 , \50881 , \50882 );
and \U$50507 ( \50884 , \50880 , \3218 );
nor \U$50508 ( \50885 , \50883 , \50884 );
and \U$50509 ( \50886 , \50877 , \50885 );
and \U$50510 ( \50887 , \50869 , \50876 );
or \U$50511 ( \50888 , \50886 , \50887 );
or \U$50512 ( \50889 , \50861 , \50888 );
not \U$50513 ( \50890 , \50861 );
not \U$50514 ( \50891 , \50888 );
or \U$50515 ( \50892 , \50890 , \50891 );
and \U$50516 ( \50893 , \1593 , RIae76fa0_66);
and \U$50517 ( \50894 , RIae76eb0_64, \1591 );
nor \U$50518 ( \50895 , \50893 , \50894 );
and \U$50519 ( \50896 , \50895 , \1488 );
not \U$50520 ( \50897 , \50895 );
and \U$50521 ( \50898 , \50897 , \1498 );
nor \U$50522 ( \50899 , \50896 , \50898 );
and \U$50523 ( \50900 , \1939 , RIae76dc0_62);
and \U$50524 ( \50901 , RIae76cd0_60, \1937 );
nor \U$50525 ( \50902 , \50900 , \50901 );
and \U$50526 ( \50903 , \50902 , \1734 );
not \U$50527 ( \50904 , \50902 );
and \U$50528 ( \50905 , \50904 , \1735 );
nor \U$50529 ( \50906 , \50903 , \50905 );
or \U$50530 ( \50907 , \50899 , \50906 );
not \U$50531 ( \50908 , \50906 );
not \U$50532 ( \50909 , \50899 );
or \U$50533 ( \50910 , \50908 , \50909 );
and \U$50534 ( \50911 , \2224 , RIae77108_69);
and \U$50535 ( \50912 , RIae77090_68, \2222 );
nor \U$50536 ( \50913 , \50911 , \50912 );
and \U$50537 ( \50914 , \50913 , \2061 );
not \U$50538 ( \50915 , \50913 );
and \U$50539 ( \50916 , \50915 , \2060 );
nor \U$50540 ( \50917 , \50914 , \50916 );
nand \U$50541 ( \50918 , \50910 , \50917 );
nand \U$50542 ( \50919 , \50907 , \50918 );
nand \U$50543 ( \50920 , \50892 , \50919 );
nand \U$50544 ( \50921 , \50889 , \50920 );
and \U$50545 ( \50922 , \50835 , \50921 );
and \U$50546 ( \50923 , \50753 , \50834 );
or \U$50547 ( \50924 , \50922 , \50923 );
xor \U$50548 ( \50925 , \50674 , \50924 );
xor \U$50549 ( \50926 , \50442 , \50444 );
xor \U$50550 ( \50927 , \50926 , \50451 );
xor \U$50551 ( \50928 , \50501 , \50507 );
xor \U$50552 ( \50929 , \50928 , \50514 );
and \U$50553 ( \50930 , \50927 , \50929 );
xor \U$50554 ( \50931 , \50003 , \50010 );
xor \U$50555 ( \50932 , \50931 , \50018 );
xor \U$50556 ( \50933 , \50420 , \50429 );
xor \U$50557 ( \50934 , \50932 , \50933 );
xor \U$50558 ( \50935 , \50501 , \50507 );
xor \U$50559 ( \50936 , \50935 , \50514 );
and \U$50560 ( \50937 , \50934 , \50936 );
and \U$50561 ( \50938 , \50927 , \50934 );
or \U$50562 ( \50939 , \50930 , \50937 , \50938 );
and \U$50563 ( \50940 , \50925 , \50939 );
and \U$50564 ( \50941 , \50674 , \50924 );
or \U$50565 ( \50942 , \50940 , \50941 );
xor \U$50566 ( \50943 , \50624 , \50942 );
not \U$50567 ( \50944 , \50534 );
xor \U$50568 ( \50945 , \50537 , \50542 );
not \U$50569 ( \50946 , \50945 );
or \U$50570 ( \50947 , \50944 , \50946 );
or \U$50571 ( \50948 , \50945 , \50534 );
nand \U$50572 ( \50949 , \50947 , \50948 );
xor \U$50573 ( \50950 , \50461 , \50468 );
xor \U$50574 ( \50951 , \50950 , \50495 );
xor \U$50575 ( \50952 , \50352 , \50379 );
xor \U$50576 ( \50953 , \50952 , \50407 );
and \U$50577 ( \50954 , \50951 , \50953 );
xor \U$50578 ( \50955 , \50200 , \50225 );
xor \U$50579 ( \50956 , \50955 , \50251 );
xor \U$50580 ( \50957 , \50352 , \50379 );
xor \U$50581 ( \50958 , \50957 , \50407 );
and \U$50582 ( \50959 , \50956 , \50958 );
and \U$50583 ( \50960 , \50951 , \50956 );
or \U$50584 ( \50961 , \50954 , \50959 , \50960 );
xor \U$50585 ( \50962 , \50949 , \50961 );
xor \U$50586 ( \50963 , \50029 , \50031 );
xor \U$50587 ( \50964 , \50963 , \50038 );
xor \U$50588 ( \50965 , \50554 , \50559 );
xor \U$50589 ( \50966 , \50964 , \50965 );
and \U$50590 ( \50967 , \50962 , \50966 );
and \U$50591 ( \50968 , \50949 , \50961 );
or \U$50592 ( \50969 , \50967 , \50968 );
and \U$50593 ( \50970 , \50943 , \50969 );
and \U$50594 ( \50971 , \50624 , \50942 );
or \U$50595 ( \50972 , \50970 , \50971 );
xor \U$50596 ( \50973 , \50041 , \50057 );
xor \U$50597 ( \50974 , \50973 , \50076 );
xor \U$50598 ( \50975 , \49855 , \49939 );
xor \U$50599 ( \50976 , \50975 , \50023 );
xor \U$50600 ( \50977 , \50974 , \50976 );
xor \U$50601 ( \50978 , \49762 , \49764 );
xor \U$50602 ( \50979 , \50978 , \49769 );
xor \U$50603 ( \50980 , \50163 , \50170 );
xor \U$50604 ( \50981 , \50979 , \50980 );
and \U$50605 ( \50982 , \50977 , \50981 );
and \U$50606 ( \50983 , \50974 , \50976 );
or \U$50607 ( \50984 , \50982 , \50983 );
xor \U$50608 ( \50985 , \50972 , \50984 );
xor \U$50609 ( \50986 , \50097 , \50099 );
xor \U$50610 ( \50987 , \50986 , \50104 );
xor \U$50611 ( \50988 , \50149 , \50156 );
xor \U$50612 ( \50989 , \50987 , \50988 );
and \U$50613 ( \50990 , \50985 , \50989 );
and \U$50614 ( \50991 , \50972 , \50984 );
or \U$50615 ( \50992 , \50990 , \50991 );
xor \U$50616 ( \50993 , \50610 , \50992 );
xor \U$50617 ( \50994 , \49760 , \50082 );
xor \U$50618 ( \50995 , \50994 , \50107 );
and \U$50619 ( \50996 , \50993 , \50995 );
and \U$50620 ( \50997 , \50610 , \50992 );
nor \U$50621 ( \50998 , \50996 , \50997 );
not \U$50622 ( \50999 , \50998 );
xor \U$50623 ( \51000 , \50135 , \50137 );
xor \U$50624 ( \51001 , \51000 , \50140 );
xor \U$50625 ( \51002 , \50577 , \50582 );
xor \U$50626 ( \51003 , \51001 , \51002 );
nand \U$50627 ( \51004 , \50999 , \51003 );
or \U$50628 ( \51005 , \50608 , \51004 );
xnor \U$50629 ( \51006 , \51004 , \50608 );
xor \U$50630 ( \51007 , \50753 , \50834 );
xor \U$50631 ( \51008 , \51007 , \50921 );
xor \U$50632 ( \51009 , \50648 , \50660 );
xor \U$50633 ( \51010 , \51009 , \50671 );
and \U$50634 ( \51011 , \51008 , \51010 );
xor \U$50635 ( \51012 , \50501 , \50507 );
xor \U$50636 ( \51013 , \51012 , \50514 );
xor \U$50637 ( \51014 , \50927 , \50934 );
xor \U$50638 ( \51015 , \51013 , \51014 );
xor \U$50639 ( \51016 , \50648 , \50660 );
xor \U$50640 ( \51017 , \51016 , \50671 );
and \U$50641 ( \51018 , \51015 , \51017 );
and \U$50642 ( \51019 , \51008 , \51015 );
or \U$50643 ( \51020 , \51011 , \51018 , \51019 );
xor \U$50644 ( \51021 , \50869 , \50876 );
xor \U$50645 ( \51022 , \51021 , \50885 );
xor \U$50646 ( \51023 , \50681 , \50688 );
xor \U$50647 ( \51024 , \51023 , \50696 );
or \U$50648 ( \51025 , \51022 , \51024 );
not \U$50649 ( \51026 , \51024 );
not \U$50650 ( \51027 , \51022 );
or \U$50651 ( \51028 , \51026 , \51027 );
xor \U$50652 ( \51029 , \50732 , \50739 );
xor \U$50653 ( \51030 , \51029 , \50747 );
nand \U$50654 ( \51031 , \51028 , \51030 );
nand \U$50655 ( \51032 , \51025 , \51031 );
and \U$50656 ( \51033 , \672 , RIae77630_80);
and \U$50657 ( \51034 , RIae77540_78, \670 );
nor \U$50658 ( \51035 , \51033 , \51034 );
and \U$50659 ( \51036 , \51035 , \587 );
not \U$50660 ( \51037 , \51035 );
and \U$50661 ( \51038 , \51037 , \588 );
nor \U$50662 ( \51039 , \51036 , \51038 );
xor \U$50663 ( \51040 , \50843 , \50850 );
xor \U$50664 ( \51041 , \51040 , \50858 );
xor \U$50665 ( \51042 , \51039 , \51041 );
not \U$50666 ( \51043 , \50906 );
not \U$50667 ( \51044 , \50917 );
or \U$50668 ( \51045 , \51043 , \51044 );
or \U$50669 ( \51046 , \50906 , \50917 );
nand \U$50670 ( \51047 , \51045 , \51046 );
not \U$50671 ( \51048 , \51047 );
not \U$50672 ( \51049 , \50899 );
and \U$50673 ( \51050 , \51048 , \51049 );
and \U$50674 ( \51051 , \51047 , \50899 );
nor \U$50675 ( \51052 , \51050 , \51051 );
and \U$50676 ( \51053 , \51042 , \51052 );
and \U$50677 ( \51054 , \51039 , \51041 );
nor \U$50678 ( \51055 , \51053 , \51054 );
xor \U$50679 ( \51056 , \51032 , \51055 );
xor \U$50680 ( \51057 , \50706 , \50713 );
xor \U$50681 ( \51058 , \51057 , \50721 );
xor \U$50682 ( \51059 , \50813 , \50820 );
xor \U$50683 ( \51060 , \51059 , \50828 );
or \U$50684 ( \51061 , \51058 , \51060 );
not \U$50685 ( \51062 , \51060 );
not \U$50686 ( \51063 , \51058 );
or \U$50687 ( \51064 , \51062 , \51063 );
not \U$50688 ( \51065 , \50785 );
xor \U$50689 ( \51066 , \50803 , \50793 );
not \U$50690 ( \51067 , \51066 );
or \U$50691 ( \51068 , \51065 , \51067 );
or \U$50692 ( \51069 , \51066 , \50785 );
nand \U$50693 ( \51070 , \51068 , \51069 );
nand \U$50694 ( \51071 , \51064 , \51070 );
nand \U$50695 ( \51072 , \51061 , \51071 );
and \U$50696 ( \51073 , \51056 , \51072 );
and \U$50697 ( \51074 , \51032 , \51055 );
or \U$50698 ( \51075 , \51073 , \51074 );
and \U$50699 ( \51076 , \4247 , RIae78620_114);
and \U$50700 ( \51077 , RIae78440_110, \4245 );
nor \U$50701 ( \51078 , \51076 , \51077 );
and \U$50702 ( \51079 , \51078 , \4251 );
not \U$50703 ( \51080 , \51078 );
and \U$50704 ( \51081 , \51080 , \3989 );
nor \U$50705 ( \51082 , \51079 , \51081 );
and \U$50706 ( \51083 , \4688 , RIae784b8_111);
and \U$50707 ( \51084 , RIae77cc0_94, \4686 );
nor \U$50708 ( \51085 , \51083 , \51084 );
and \U$50709 ( \51086 , \51085 , \4482 );
not \U$50710 ( \51087 , \51085 );
and \U$50711 ( \51088 , \51087 , \4481 );
nor \U$50712 ( \51089 , \51086 , \51088 );
xor \U$50713 ( \51090 , \51082 , \51089 );
and \U$50714 ( \51091 , \5399 , RIae77bd0_92);
and \U$50715 ( \51092 , RIae77db0_96, \5397 );
nor \U$50716 ( \51093 , \51091 , \51092 );
and \U$50717 ( \51094 , \51093 , \5403 );
not \U$50718 ( \51095 , \51093 );
and \U$50719 ( \51096 , \51095 , \5016 );
nor \U$50720 ( \51097 , \51094 , \51096 );
and \U$50721 ( \51098 , \51090 , \51097 );
and \U$50722 ( \51099 , \51082 , \51089 );
or \U$50723 ( \51100 , \51098 , \51099 );
and \U$50724 ( \51101 , \7633 , RIae75b00_22);
and \U$50725 ( \51102 , RIae75a10_20, \7631 );
nor \U$50726 ( \51103 , \51101 , \51102 );
and \U$50727 ( \51104 , \51103 , \7205 );
not \U$50728 ( \51105 , \51103 );
and \U$50729 ( \51106 , \51105 , \7206 );
nor \U$50730 ( \51107 , \51104 , \51106 );
not \U$50731 ( \51108 , \51107 );
and \U$50732 ( \51109 , \8966 , RIae75ec0_30);
and \U$50733 ( \51110 , RIae75ce0_26, \8964 );
nor \U$50734 ( \51111 , \51109 , \51110 );
and \U$50735 ( \51112 , \51111 , \8789 );
not \U$50736 ( \51113 , \51111 );
and \U$50737 ( \51114 , \51113 , \8799 );
nor \U$50738 ( \51115 , \51112 , \51114 );
not \U$50739 ( \51116 , \51115 );
and \U$50740 ( \51117 , \51108 , \51116 );
and \U$50741 ( \51118 , \51115 , \51107 );
and \U$50742 ( \51119 , \8371 , RIae75920_18);
and \U$50743 ( \51120 , RIae75fb0_32, \8369 );
nor \U$50744 ( \51121 , \51119 , \51120 );
and \U$50745 ( \51122 , \51121 , \8019 );
not \U$50746 ( \51123 , \51121 );
and \U$50747 ( \51124 , \51123 , \8020 );
nor \U$50748 ( \51125 , \51122 , \51124 );
nor \U$50749 ( \51126 , \51118 , \51125 );
nor \U$50750 ( \51127 , \51117 , \51126 );
or \U$50751 ( \51128 , \51100 , \51127 );
not \U$50752 ( \51129 , \51100 );
not \U$50753 ( \51130 , \51127 );
or \U$50754 ( \51131 , \51129 , \51130 );
and \U$50755 ( \51132 , \5896 , RIae77ea0_98);
and \U$50756 ( \51133 , RIae789e0_122, \5894 );
nor \U$50757 ( \51134 , \51132 , \51133 );
and \U$50758 ( \51135 , \51134 , \5590 );
not \U$50759 ( \51136 , \51134 );
and \U$50760 ( \51137 , \51136 , \5589 );
nor \U$50761 ( \51138 , \51135 , \51137 );
and \U$50762 ( \51139 , \6172 , RIae788f0_120);
and \U$50763 ( \51140 , RIae78800_118, \6170 );
nor \U$50764 ( \51141 , \51139 , \51140 );
and \U$50765 ( \51142 , \51141 , \6176 );
not \U$50766 ( \51143 , \51141 );
and \U$50767 ( \51144 , \51143 , \6175 );
nor \U$50768 ( \51145 , \51142 , \51144 );
xor \U$50769 ( \51146 , \51138 , \51145 );
and \U$50770 ( \51147 , \6941 , RIae78710_116);
and \U$50771 ( \51148 , RIae75bf0_24, \6939 );
nor \U$50772 ( \51149 , \51147 , \51148 );
and \U$50773 ( \51150 , \51149 , \6314 );
not \U$50774 ( \51151 , \51149 );
and \U$50775 ( \51152 , \51151 , \6945 );
nor \U$50776 ( \51153 , \51150 , \51152 );
and \U$50777 ( \51154 , \51146 , \51153 );
and \U$50778 ( \51155 , \51138 , \51145 );
or \U$50779 ( \51156 , \51154 , \51155 );
nand \U$50780 ( \51157 , \51131 , \51156 );
nand \U$50781 ( \51158 , \51128 , \51157 );
and \U$50782 ( \51159 , \13059 , RIae75470_8);
and \U$50783 ( \51160 , RIae76460_42, \13057 );
nor \U$50784 ( \51161 , \51159 , \51160 );
and \U$50785 ( \51162 , \51161 , \13063 );
not \U$50786 ( \51163 , \51161 );
and \U$50787 ( \51164 , \51163 , \12718 );
nor \U$50788 ( \51165 , \51162 , \51164 );
and \U$50789 ( \51166 , \12180 , RIae751a0_2);
and \U$50790 ( \51167 , RIae75380_6, \12178 );
nor \U$50791 ( \51168 , \51166 , \51167 );
and \U$50792 ( \51169 , \51168 , \12184 );
not \U$50793 ( \51170 , \51168 );
and \U$50794 ( \51171 , \51170 , \11827 );
nor \U$50795 ( \51172 , \51169 , \51171 );
xor \U$50796 ( \51173 , \51165 , \51172 );
and \U$50797 ( \51174 , \14059 , RIae76550_44);
and \U$50798 ( \51175 , RIae76730_48, \14057 );
nor \U$50799 ( \51176 , \51174 , \51175 );
and \U$50800 ( \51177 , \51176 , \13502 );
not \U$50801 ( \51178 , \51176 );
and \U$50802 ( \51179 , \51178 , \14063 );
nor \U$50803 ( \51180 , \51177 , \51179 );
and \U$50804 ( \51181 , \51173 , \51180 );
and \U$50805 ( \51182 , \51165 , \51172 );
or \U$50806 ( \51183 , \51181 , \51182 );
and \U$50807 ( \51184 , \15726 , RIae760a0_34);
and \U$50808 ( \51185 , RIae76370_40, RIae7aab0_192);
nor \U$50809 ( \51186 , \51184 , \51185 );
and \U$50810 ( \51187 , \51186 , \14959 );
not \U$50811 ( \51188 , \51186 );
and \U$50812 ( \51189 , \51188 , RIae7aa38_191);
nor \U$50813 ( \51190 , \51187 , \51189 );
xor \U$50814 ( \51191 , \51190 , \587 );
and \U$50815 ( \51192 , \14964 , RIae76640_46);
and \U$50816 ( \51193 , RIae76190_36, \14962 );
nor \U$50817 ( \51194 , \51192 , \51193 );
and \U$50818 ( \51195 , \51194 , \14463 );
not \U$50819 ( \51196 , \51194 );
and \U$50820 ( \51197 , \51196 , \14462 );
nor \U$50821 ( \51198 , \51195 , \51197 );
and \U$50822 ( \51199 , \51191 , \51198 );
and \U$50823 ( \51200 , \51190 , \587 );
or \U$50824 ( \51201 , \51199 , \51200 );
xor \U$50825 ( \51202 , \51183 , \51201 );
and \U$50826 ( \51203 , \9760 , RIae75dd0_28);
and \U$50827 ( \51204 , RIae75650_12, \9758 );
nor \U$50828 ( \51205 , \51203 , \51204 );
and \U$50829 ( \51206 , \51205 , \9273 );
not \U$50830 ( \51207 , \51205 );
and \U$50831 ( \51208 , \51207 , \9272 );
nor \U$50832 ( \51209 , \51206 , \51208 );
and \U$50833 ( \51210 , \10548 , RIae75560_10);
and \U$50834 ( \51211 , RIae75830_16, \10546 );
nor \U$50835 ( \51212 , \51210 , \51211 );
and \U$50836 ( \51213 , \51212 , \10421 );
not \U$50837 ( \51214 , \51212 );
and \U$50838 ( \51215 , \51214 , \10118 );
nor \U$50839 ( \51216 , \51213 , \51215 );
xor \U$50840 ( \51217 , \51209 , \51216 );
and \U$50841 ( \51218 , \11470 , RIae75740_14);
and \U$50842 ( \51219 , RIae75290_4, \11468 );
nor \U$50843 ( \51220 , \51218 , \51219 );
and \U$50844 ( \51221 , \51220 , \10936 );
not \U$50845 ( \51222 , \51220 );
and \U$50846 ( \51223 , \51222 , \11474 );
nor \U$50847 ( \51224 , \51221 , \51223 );
and \U$50848 ( \51225 , \51217 , \51224 );
and \U$50849 ( \51226 , \51209 , \51216 );
or \U$50850 ( \51227 , \51225 , \51226 );
and \U$50851 ( \51228 , \51202 , \51227 );
and \U$50852 ( \51229 , \51183 , \51201 );
or \U$50853 ( \51230 , \51228 , \51229 );
xor \U$50854 ( \51231 , \51158 , \51230 );
and \U$50855 ( \51232 , \2224 , RIae76cd0_60);
and \U$50856 ( \51233 , RIae77108_69, \2222 );
nor \U$50857 ( \51234 , \51232 , \51233 );
and \U$50858 ( \51235 , \51234 , \2060 );
not \U$50859 ( \51236 , \51234 );
and \U$50860 ( \51237 , \51236 , \2061 );
nor \U$50861 ( \51238 , \51235 , \51237 );
and \U$50862 ( \51239 , \1939 , RIae76eb0_64);
and \U$50863 ( \51240 , RIae76dc0_62, \1937 );
nor \U$50864 ( \51241 , \51239 , \51240 );
and \U$50865 ( \51242 , \51241 , \1734 );
not \U$50866 ( \51243 , \51241 );
and \U$50867 ( \51244 , \51243 , \1735 );
nor \U$50868 ( \51245 , \51242 , \51244 );
xor \U$50869 ( \51246 , \51238 , \51245 );
and \U$50870 ( \51247 , \2607 , RIae77090_68);
and \U$50871 ( \51248 , RIae77270_72, \2605 );
nor \U$50872 ( \51249 , \51247 , \51248 );
and \U$50873 ( \51250 , \51249 , \2397 );
not \U$50874 ( \51251 , \51249 );
and \U$50875 ( \51252 , \51251 , \2611 );
nor \U$50876 ( \51253 , \51250 , \51252 );
and \U$50877 ( \51254 , \51246 , \51253 );
and \U$50878 ( \51255 , \51238 , \51245 );
or \U$50879 ( \51256 , \51254 , \51255 );
and \U$50880 ( \51257 , \3730 , RIae78080_102);
and \U$50881 ( \51258 , RIae78260_106, \3728 );
nor \U$50882 ( \51259 , \51257 , \51258 );
and \U$50883 ( \51260 , \51259 , \3422 );
not \U$50884 ( \51261 , \51259 );
and \U$50885 ( \51262 , \51261 , \3732 );
nor \U$50886 ( \51263 , \51260 , \51262 );
and \U$50887 ( \51264 , \2783 , RIae77360_74);
and \U$50888 ( \51265 , RIae78350_108, \2781 );
nor \U$50889 ( \51266 , \51264 , \51265 );
not \U$50890 ( \51267 , \51266 );
not \U$50891 ( \51268 , \2789 );
and \U$50892 ( \51269 , \51267 , \51268 );
and \U$50893 ( \51270 , \51266 , \3089 );
nor \U$50894 ( \51271 , \51269 , \51270 );
xor \U$50895 ( \51272 , \51263 , \51271 );
and \U$50896 ( \51273 , \3214 , RIae78170_104);
and \U$50897 ( \51274 , RIae77f90_100, \3212 );
nor \U$50898 ( \51275 , \51273 , \51274 );
not \U$50899 ( \51276 , \51275 );
not \U$50900 ( \51277 , \3218 );
and \U$50901 ( \51278 , \51276 , \51277 );
and \U$50902 ( \51279 , \51275 , \2774 );
nor \U$50903 ( \51280 , \51278 , \51279 );
and \U$50904 ( \51281 , \51272 , \51280 );
and \U$50905 ( \51282 , \51263 , \51271 );
or \U$50906 ( \51283 , \51281 , \51282 );
or \U$50907 ( \51284 , \51256 , \51283 );
not \U$50908 ( \51285 , \51256 );
not \U$50909 ( \51286 , \51283 );
or \U$50910 ( \51287 , \51285 , \51286 );
and \U$50911 ( \51288 , \1593 , RIae77900_86);
and \U$50912 ( \51289 , RIae76fa0_66, \1591 );
nor \U$50913 ( \51290 , \51288 , \51289 );
and \U$50914 ( \51291 , \51290 , \1498 );
not \U$50915 ( \51292 , \51290 );
and \U$50916 ( \51293 , \51292 , \1488 );
nor \U$50917 ( \51294 , \51291 , \51293 );
and \U$50918 ( \51295 , \1138 , RIae77450_76);
and \U$50919 ( \51296 , RIae77ae0_90, \1136 );
nor \U$50920 ( \51297 , \51295 , \51296 );
and \U$50921 ( \51298 , \51297 , \1012 );
not \U$50922 ( \51299 , \51297 );
and \U$50923 ( \51300 , \51299 , \1142 );
nor \U$50924 ( \51301 , \51298 , \51300 );
xor \U$50925 ( \51302 , \51294 , \51301 );
and \U$50926 ( \51303 , \1376 , RIae779f0_88);
and \U$50927 ( \51304 , RIae77810_84, \1374 );
nor \U$50928 ( \51305 , \51303 , \51304 );
and \U$50929 ( \51306 , \51305 , \1380 );
not \U$50930 ( \51307 , \51305 );
and \U$50931 ( \51308 , \51307 , \1261 );
nor \U$50932 ( \51309 , \51306 , \51308 );
and \U$50933 ( \51310 , \51302 , \51309 );
and \U$50934 ( \51311 , \51294 , \51301 );
or \U$50935 ( \51312 , \51310 , \51311 );
nand \U$50936 ( \51313 , \51287 , \51312 );
nand \U$50937 ( \51314 , \51284 , \51313 );
and \U$50938 ( \51315 , \51231 , \51314 );
and \U$50939 ( \51316 , \51158 , \51230 );
or \U$50940 ( \51317 , \51315 , \51316 );
xor \U$50941 ( \51318 , \51075 , \51317 );
xor \U$50942 ( \51319 , \50286 , \562 );
xor \U$50943 ( \51320 , \51319 , \50294 );
xor \U$50944 ( \51321 , \50663 , \50665 );
xor \U$50945 ( \51322 , \51321 , \50668 );
and \U$50946 ( \51323 , \51320 , \51322 );
xor \U$50947 ( \51324 , \50233 , \50240 );
xor \U$50948 ( \51325 , \51324 , \50248 );
xor \U$50949 ( \51326 , \50650 , \50655 );
xor \U$50950 ( \51327 , \51325 , \51326 );
xor \U$50951 ( \51328 , \50663 , \50665 );
xor \U$50952 ( \51329 , \51328 , \50668 );
and \U$50953 ( \51330 , \51327 , \51329 );
and \U$50954 ( \51331 , \51320 , \51327 );
or \U$50955 ( \51332 , \51323 , \51330 , \51331 );
and \U$50956 ( \51333 , \51318 , \51332 );
and \U$50957 ( \51334 , \51075 , \51317 );
or \U$50958 ( \51335 , \51333 , \51334 );
xor \U$50959 ( \51336 , \51020 , \51335 );
not \U$50960 ( \51337 , \50919 );
not \U$50961 ( \51338 , \50861 );
or \U$50962 ( \51339 , \51337 , \51338 );
or \U$50963 ( \51340 , \50861 , \50919 );
nand \U$50964 ( \51341 , \51339 , \51340 );
not \U$50965 ( \51342 , \51341 );
not \U$50966 ( \51343 , \50888 );
and \U$50967 ( \51344 , \51342 , \51343 );
and \U$50968 ( \51345 , \51341 , \50888 );
nor \U$50969 ( \51346 , \51344 , \51345 );
xor \U$50970 ( \51347 , \50699 , \50724 );
xor \U$50971 ( \51348 , \51347 , \50750 );
xor \U$50972 ( \51349 , \51346 , \51348 );
not \U$50973 ( \51350 , \50646 );
not \U$50974 ( \51351 , \50630 );
or \U$50975 ( \51352 , \51350 , \51351 );
or \U$50976 ( \51353 , \50630 , \50646 );
nand \U$50977 ( \51354 , \51352 , \51353 );
not \U$50978 ( \51355 , \51354 );
not \U$50979 ( \51356 , \50640 );
and \U$50980 ( \51357 , \51355 , \51356 );
and \U$50981 ( \51358 , \51354 , \50640 );
nor \U$50982 ( \51359 , \51357 , \51358 );
and \U$50983 ( \51360 , \51349 , \51359 );
and \U$50984 ( \51361 , \51346 , \51348 );
nor \U$50985 ( \51362 , \51360 , \51361 );
xor \U$50986 ( \51363 , \50279 , \50297 );
xor \U$50987 ( \51364 , \51363 , \50323 );
xor \U$50988 ( \51365 , \51362 , \51364 );
xor \U$50989 ( \51366 , \50352 , \50379 );
xor \U$50990 ( \51367 , \51366 , \50407 );
xor \U$50991 ( \51368 , \50951 , \50956 );
xor \U$50992 ( \51369 , \51367 , \51368 );
and \U$50993 ( \51370 , \51365 , \51369 );
and \U$50994 ( \51371 , \51362 , \51364 );
or \U$50995 ( \51372 , \51370 , \51371 );
and \U$50996 ( \51373 , \51336 , \51372 );
and \U$50997 ( \51374 , \51020 , \51335 );
or \U$50998 ( \51375 , \51373 , \51374 );
not \U$50999 ( \51376 , \51375 );
xor \U$51000 ( \51377 , \50454 , \50498 );
xor \U$51001 ( \51378 , \51377 , \50517 );
xor \U$51002 ( \51379 , \50612 , \50619 );
xor \U$51003 ( \51380 , \51378 , \51379 );
xor \U$51004 ( \51381 , \50674 , \50924 );
xor \U$51005 ( \51382 , \51381 , \50939 );
and \U$51006 ( \51383 , \51380 , \51382 );
xor \U$51007 ( \51384 , \50949 , \50961 );
xor \U$51008 ( \51385 , \51384 , \50966 );
or \U$51009 ( \51386 , \51380 , \51382 );
and \U$51010 ( \51387 , \51385 , \51386 );
nor \U$51011 ( \51388 , \51383 , \51387 );
not \U$51012 ( \51389 , \51388 );
or \U$51013 ( \51390 , \51376 , \51389 );
or \U$51014 ( \51391 , \51388 , \51375 );
nand \U$51015 ( \51392 , \51390 , \51391 );
not \U$51016 ( \51393 , \51392 );
not \U$51017 ( \51394 , \50564 );
not \U$51018 ( \51395 , \50544 );
or \U$51019 ( \51396 , \51394 , \51395 );
or \U$51020 ( \51397 , \50544 , \50564 );
nand \U$51021 ( \51398 , \51396 , \51397 );
not \U$51022 ( \51399 , \51398 );
not \U$51023 ( \51400 , \50546 );
and \U$51024 ( \51401 , \51399 , \51400 );
and \U$51025 ( \51402 , \51398 , \50546 );
nor \U$51026 ( \51403 , \51401 , \51402 );
not \U$51027 ( \51404 , \51403 );
and \U$51028 ( \51405 , \51393 , \51404 );
and \U$51029 ( \51406 , \51392 , \51403 );
nor \U$51030 ( \51407 , \51405 , \51406 );
not \U$51031 ( \51408 , \51407 );
xor \U$51032 ( \51409 , \51075 , \51317 );
xor \U$51033 ( \51410 , \51409 , \51332 );
xor \U$51034 ( \51411 , \51362 , \51364 );
xor \U$51035 ( \51412 , \51411 , \51369 );
and \U$51036 ( \51413 , \51410 , \51412 );
xor \U$51037 ( \51414 , \50648 , \50660 );
xor \U$51038 ( \51415 , \51414 , \50671 );
xor \U$51039 ( \51416 , \51008 , \51015 );
xor \U$51040 ( \51417 , \51415 , \51416 );
xor \U$51041 ( \51418 , \51362 , \51364 );
xor \U$51042 ( \51419 , \51418 , \51369 );
and \U$51043 ( \51420 , \51417 , \51419 );
and \U$51044 ( \51421 , \51410 , \51417 );
or \U$51045 ( \51422 , \51413 , \51420 , \51421 );
xor \U$51046 ( \51423 , \51346 , \51348 );
xor \U$51047 ( \51424 , \51423 , \51359 );
xor \U$51048 ( \51425 , \50778 , \50805 );
xor \U$51049 ( \51426 , \51425 , \50831 );
or \U$51050 ( \51427 , \51424 , \51426 );
not \U$51051 ( \51428 , \51426 );
not \U$51052 ( \51429 , \51424 );
or \U$51053 ( \51430 , \51428 , \51429 );
not \U$51054 ( \51431 , \51312 );
not \U$51055 ( \51432 , \51283 );
or \U$51056 ( \51433 , \51431 , \51432 );
or \U$51057 ( \51434 , \51283 , \51312 );
nand \U$51058 ( \51435 , \51433 , \51434 );
not \U$51059 ( \51436 , \51435 );
not \U$51060 ( \51437 , \51256 );
and \U$51061 ( \51438 , \51436 , \51437 );
and \U$51062 ( \51439 , \51435 , \51256 );
nor \U$51063 ( \51440 , \51438 , \51439 );
not \U$51064 ( \51441 , \51156 );
not \U$51065 ( \51442 , \51100 );
or \U$51066 ( \51443 , \51441 , \51442 );
or \U$51067 ( \51444 , \51100 , \51156 );
nand \U$51068 ( \51445 , \51443 , \51444 );
not \U$51069 ( \51446 , \51445 );
not \U$51070 ( \51447 , \51127 );
and \U$51071 ( \51448 , \51446 , \51447 );
and \U$51072 ( \51449 , \51445 , \51127 );
nor \U$51073 ( \51450 , \51448 , \51449 );
xor \U$51074 ( \51451 , \51440 , \51450 );
xor \U$51075 ( \51452 , \51039 , \51041 );
xor \U$51076 ( \51453 , \51452 , \51052 );
and \U$51077 ( \51454 , \51451 , \51453 );
and \U$51078 ( \51455 , \51440 , \51450 );
nor \U$51079 ( \51456 , \51454 , \51455 );
nand \U$51080 ( \51457 , \51430 , \51456 );
nand \U$51081 ( \51458 , \51427 , \51457 );
not \U$51082 ( \51459 , \2774 );
and \U$51083 ( \51460 , \3214 , RIae78350_108);
and \U$51084 ( \51461 , RIae78170_104, \3212 );
nor \U$51085 ( \51462 , \51460 , \51461 );
not \U$51086 ( \51463 , \51462 );
or \U$51087 ( \51464 , \51459 , \51463 );
or \U$51088 ( \51465 , \51462 , \3218 );
nand \U$51089 ( \51466 , \51464 , \51465 );
and \U$51090 ( \51467 , \2607 , RIae77108_69);
and \U$51091 ( \51468 , RIae77090_68, \2605 );
nor \U$51092 ( \51469 , \51467 , \51468 );
and \U$51093 ( \51470 , \51469 , \2611 );
not \U$51094 ( \51471 , \51469 );
and \U$51095 ( \51472 , \51471 , \2397 );
nor \U$51096 ( \51473 , \51470 , \51472 );
xor \U$51097 ( \51474 , \51466 , \51473 );
not \U$51098 ( \51475 , \2789 );
and \U$51099 ( \51476 , \2783 , RIae77270_72);
and \U$51100 ( \51477 , RIae77360_74, \2781 );
nor \U$51101 ( \51478 , \51476 , \51477 );
not \U$51102 ( \51479 , \51478 );
or \U$51103 ( \51480 , \51475 , \51479 );
or \U$51104 ( \51481 , \51478 , \3089 );
nand \U$51105 ( \51482 , \51480 , \51481 );
and \U$51106 ( \51483 , \51474 , \51482 );
and \U$51107 ( \51484 , \51466 , \51473 );
or \U$51108 ( \51485 , \51483 , \51484 );
and \U$51109 ( \51486 , \1376 , RIae77ae0_90);
and \U$51110 ( \51487 , RIae779f0_88, \1374 );
nor \U$51111 ( \51488 , \51486 , \51487 );
and \U$51112 ( \51489 , \51488 , \1380 );
not \U$51113 ( \51490 , \51488 );
and \U$51114 ( \51491 , \51490 , \1261 );
nor \U$51115 ( \51492 , \51489 , \51491 );
not \U$51116 ( \51493 , \789 );
and \U$51117 ( \51494 , \883 , RIae77630_80);
and \U$51118 ( \51495 , RIae77540_78, \881 );
nor \U$51119 ( \51496 , \51494 , \51495 );
not \U$51120 ( \51497 , \51496 );
or \U$51121 ( \51498 , \51493 , \51497 );
or \U$51122 ( \51499 , \51496 , \789 );
nand \U$51123 ( \51500 , \51498 , \51499 );
xor \U$51124 ( \51501 , \51492 , \51500 );
and \U$51125 ( \51502 , \1138 , RIae776a8_81);
and \U$51126 ( \51503 , RIae77450_76, \1136 );
nor \U$51127 ( \51504 , \51502 , \51503 );
and \U$51128 ( \51505 , \51504 , \1012 );
not \U$51129 ( \51506 , \51504 );
and \U$51130 ( \51507 , \51506 , \1142 );
nor \U$51131 ( \51508 , \51505 , \51507 );
and \U$51132 ( \51509 , \51501 , \51508 );
and \U$51133 ( \51510 , \51492 , \51500 );
or \U$51134 ( \51511 , \51509 , \51510 );
xor \U$51135 ( \51512 , \51485 , \51511 );
and \U$51136 ( \51513 , \2224 , RIae76dc0_62);
and \U$51137 ( \51514 , RIae76cd0_60, \2222 );
nor \U$51138 ( \51515 , \51513 , \51514 );
and \U$51139 ( \51516 , \51515 , \2061 );
not \U$51140 ( \51517 , \51515 );
and \U$51141 ( \51518 , \51517 , \2060 );
nor \U$51142 ( \51519 , \51516 , \51518 );
and \U$51143 ( \51520 , \1593 , RIae77810_84);
and \U$51144 ( \51521 , RIae77900_86, \1591 );
nor \U$51145 ( \51522 , \51520 , \51521 );
and \U$51146 ( \51523 , \51522 , \1498 );
not \U$51147 ( \51524 , \51522 );
and \U$51148 ( \51525 , \51524 , \1488 );
nor \U$51149 ( \51526 , \51523 , \51525 );
xor \U$51150 ( \51527 , \51519 , \51526 );
and \U$51151 ( \51528 , \1939 , RIae76fa0_66);
and \U$51152 ( \51529 , RIae76eb0_64, \1937 );
nor \U$51153 ( \51530 , \51528 , \51529 );
and \U$51154 ( \51531 , \51530 , \1735 );
not \U$51155 ( \51532 , \51530 );
and \U$51156 ( \51533 , \51532 , \1734 );
nor \U$51157 ( \51534 , \51531 , \51533 );
and \U$51158 ( \51535 , \51527 , \51534 );
and \U$51159 ( \51536 , \51519 , \51526 );
or \U$51160 ( \51537 , \51535 , \51536 );
and \U$51161 ( \51538 , \51512 , \51537 );
and \U$51162 ( \51539 , \51485 , \51511 );
nor \U$51163 ( \51540 , \51538 , \51539 );
and \U$51164 ( \51541 , \13059 , RIae75380_6);
and \U$51165 ( \51542 , RIae75470_8, \13057 );
nor \U$51166 ( \51543 , \51541 , \51542 );
and \U$51167 ( \51544 , \51543 , \13063 );
not \U$51168 ( \51545 , \51543 );
and \U$51169 ( \51546 , \51545 , \12718 );
nor \U$51170 ( \51547 , \51544 , \51546 );
and \U$51171 ( \51548 , \11470 , RIae75830_16);
and \U$51172 ( \51549 , RIae75740_14, \11468 );
nor \U$51173 ( \51550 , \51548 , \51549 );
and \U$51174 ( \51551 , \51550 , \10936 );
not \U$51175 ( \51552 , \51550 );
and \U$51176 ( \51553 , \51552 , \11474 );
nor \U$51177 ( \51554 , \51551 , \51553 );
xor \U$51178 ( \51555 , \51547 , \51554 );
and \U$51179 ( \51556 , \12180 , RIae75290_4);
and \U$51180 ( \51557 , RIae751a0_2, \12178 );
nor \U$51181 ( \51558 , \51556 , \51557 );
and \U$51182 ( \51559 , \51558 , \12184 );
not \U$51183 ( \51560 , \51558 );
and \U$51184 ( \51561 , \51560 , \11827 );
nor \U$51185 ( \51562 , \51559 , \51561 );
and \U$51186 ( \51563 , \51555 , \51562 );
and \U$51187 ( \51564 , \51547 , \51554 );
or \U$51188 ( \51565 , \51563 , \51564 );
and \U$51189 ( \51566 , \8966 , RIae75fb0_32);
and \U$51190 ( \51567 , RIae75ec0_30, \8964 );
nor \U$51191 ( \51568 , \51566 , \51567 );
and \U$51192 ( \51569 , \51568 , \8799 );
not \U$51193 ( \51570 , \51568 );
and \U$51194 ( \51571 , \51570 , \8789 );
nor \U$51195 ( \51572 , \51569 , \51571 );
and \U$51196 ( \51573 , \9760 , RIae75ce0_26);
and \U$51197 ( \51574 , RIae75dd0_28, \9758 );
nor \U$51198 ( \51575 , \51573 , \51574 );
and \U$51199 ( \51576 , \51575 , \9273 );
not \U$51200 ( \51577 , \51575 );
and \U$51201 ( \51578 , \51577 , \9764 );
nor \U$51202 ( \51579 , \51576 , \51578 );
xor \U$51203 ( \51580 , \51572 , \51579 );
and \U$51204 ( \51581 , \10548 , RIae75650_12);
and \U$51205 ( \51582 , RIae75560_10, \10546 );
nor \U$51206 ( \51583 , \51581 , \51582 );
and \U$51207 ( \51584 , \51583 , \10421 );
not \U$51208 ( \51585 , \51583 );
and \U$51209 ( \51586 , \51585 , \10118 );
nor \U$51210 ( \51587 , \51584 , \51586 );
and \U$51211 ( \51588 , \51580 , \51587 );
and \U$51212 ( \51589 , \51572 , \51579 );
or \U$51213 ( \51590 , \51588 , \51589 );
xor \U$51214 ( \51591 , \51565 , \51590 );
and \U$51215 ( \51592 , \14964 , RIae76730_48);
and \U$51216 ( \51593 , RIae76640_46, \14962 );
nor \U$51217 ( \51594 , \51592 , \51593 );
and \U$51218 ( \51595 , \51594 , \14463 );
not \U$51219 ( \51596 , \51594 );
and \U$51220 ( \51597 , \51596 , \14462 );
nor \U$51221 ( \51598 , \51595 , \51597 );
and \U$51222 ( \51599 , \15726 , RIae76190_36);
and \U$51223 ( \51600 , RIae760a0_34, RIae7aab0_192);
nor \U$51224 ( \51601 , \51599 , \51600 );
and \U$51225 ( \51602 , \51601 , \14959 );
not \U$51226 ( \51603 , \51601 );
and \U$51227 ( \51604 , \51603 , RIae7aa38_191);
nor \U$51228 ( \51605 , \51602 , \51604 );
xor \U$51229 ( \51606 , \51598 , \51605 );
and \U$51230 ( \51607 , \14059 , RIae76460_42);
and \U$51231 ( \51608 , RIae76550_44, \14057 );
nor \U$51232 ( \51609 , \51607 , \51608 );
and \U$51233 ( \51610 , \51609 , \13502 );
not \U$51234 ( \51611 , \51609 );
and \U$51235 ( \51612 , \51611 , \14063 );
nor \U$51236 ( \51613 , \51610 , \51612 );
and \U$51237 ( \51614 , \51606 , \51613 );
and \U$51238 ( \51615 , \51598 , \51605 );
or \U$51239 ( \51616 , \51614 , \51615 );
and \U$51240 ( \51617 , \51591 , \51616 );
and \U$51241 ( \51618 , \51565 , \51590 );
nor \U$51242 ( \51619 , \51617 , \51618 );
xor \U$51243 ( \51620 , \51540 , \51619 );
and \U$51244 ( \51621 , \5399 , RIae77cc0_94);
and \U$51245 ( \51622 , RIae77bd0_92, \5397 );
nor \U$51246 ( \51623 , \51621 , \51622 );
and \U$51247 ( \51624 , \51623 , \5016 );
not \U$51248 ( \51625 , \51623 );
and \U$51249 ( \51626 , \51625 , \5403 );
nor \U$51250 ( \51627 , \51624 , \51626 );
and \U$51251 ( \51628 , \5896 , RIae77db0_96);
and \U$51252 ( \51629 , RIae77ea0_98, \5894 );
nor \U$51253 ( \51630 , \51628 , \51629 );
and \U$51254 ( \51631 , \51630 , \5590 );
not \U$51255 ( \51632 , \51630 );
and \U$51256 ( \51633 , \51632 , \5589 );
nor \U$51257 ( \51634 , \51631 , \51633 );
xor \U$51258 ( \51635 , \51627 , \51634 );
and \U$51259 ( \51636 , \6172 , RIae789e0_122);
and \U$51260 ( \51637 , RIae788f0_120, \6170 );
nor \U$51261 ( \51638 , \51636 , \51637 );
and \U$51262 ( \51639 , \51638 , \6176 );
not \U$51263 ( \51640 , \51638 );
and \U$51264 ( \51641 , \51640 , \6175 );
nor \U$51265 ( \51642 , \51639 , \51641 );
and \U$51266 ( \51643 , \51635 , \51642 );
and \U$51267 ( \51644 , \51627 , \51634 );
or \U$51268 ( \51645 , \51643 , \51644 );
and \U$51269 ( \51646 , \4247 , RIae78260_106);
and \U$51270 ( \51647 , RIae78620_114, \4245 );
nor \U$51271 ( \51648 , \51646 , \51647 );
and \U$51272 ( \51649 , \51648 , \3989 );
not \U$51273 ( \51650 , \51648 );
and \U$51274 ( \51651 , \51650 , \4251 );
nor \U$51275 ( \51652 , \51649 , \51651 );
and \U$51276 ( \51653 , \3730 , RIae77f90_100);
and \U$51277 ( \51654 , RIae78080_102, \3728 );
nor \U$51278 ( \51655 , \51653 , \51654 );
and \U$51279 ( \51656 , \51655 , \3732 );
not \U$51280 ( \51657 , \51655 );
and \U$51281 ( \51658 , \51657 , \3422 );
nor \U$51282 ( \51659 , \51656 , \51658 );
xor \U$51283 ( \51660 , \51652 , \51659 );
and \U$51284 ( \51661 , \4688 , RIae78440_110);
and \U$51285 ( \51662 , RIae784b8_111, \4686 );
nor \U$51286 ( \51663 , \51661 , \51662 );
and \U$51287 ( \51664 , \51663 , \4481 );
not \U$51288 ( \51665 , \51663 );
and \U$51289 ( \51666 , \51665 , \4482 );
nor \U$51290 ( \51667 , \51664 , \51666 );
and \U$51291 ( \51668 , \51660 , \51667 );
and \U$51292 ( \51669 , \51652 , \51659 );
or \U$51293 ( \51670 , \51668 , \51669 );
xor \U$51294 ( \51671 , \51645 , \51670 );
and \U$51295 ( \51672 , \6941 , RIae78800_118);
and \U$51296 ( \51673 , RIae78710_116, \6939 );
nor \U$51297 ( \51674 , \51672 , \51673 );
and \U$51298 ( \51675 , \51674 , \6314 );
not \U$51299 ( \51676 , \51674 );
and \U$51300 ( \51677 , \51676 , \6945 );
nor \U$51301 ( \51678 , \51675 , \51677 );
and \U$51302 ( \51679 , \7633 , RIae75bf0_24);
and \U$51303 ( \51680 , RIae75b00_22, \7631 );
nor \U$51304 ( \51681 , \51679 , \51680 );
and \U$51305 ( \51682 , \51681 , \7206 );
not \U$51306 ( \51683 , \51681 );
and \U$51307 ( \51684 , \51683 , \7205 );
nor \U$51308 ( \51685 , \51682 , \51684 );
xor \U$51309 ( \51686 , \51678 , \51685 );
and \U$51310 ( \51687 , \8371 , RIae75a10_20);
and \U$51311 ( \51688 , RIae75920_18, \8369 );
nor \U$51312 ( \51689 , \51687 , \51688 );
and \U$51313 ( \51690 , \51689 , \8020 );
not \U$51314 ( \51691 , \51689 );
and \U$51315 ( \51692 , \51691 , \8019 );
nor \U$51316 ( \51693 , \51690 , \51692 );
and \U$51317 ( \51694 , \51686 , \51693 );
and \U$51318 ( \51695 , \51678 , \51685 );
or \U$51319 ( \51696 , \51694 , \51695 );
and \U$51320 ( \51697 , \51671 , \51696 );
and \U$51321 ( \51698 , \51645 , \51670 );
nor \U$51322 ( \51699 , \51697 , \51698 );
and \U$51323 ( \51700 , \51620 , \51699 );
and \U$51324 ( \51701 , \51540 , \51619 );
or \U$51325 ( \51702 , \51700 , \51701 );
xor \U$51326 ( \51703 , \51238 , \51245 );
xor \U$51327 ( \51704 , \51703 , \51253 );
not \U$51328 ( \51705 , \51704 );
xor \U$51329 ( \51706 , \51263 , \51271 );
xor \U$51330 ( \51707 , \51706 , \51280 );
not \U$51331 ( \51708 , \51707 );
and \U$51332 ( \51709 , \51705 , \51708 );
and \U$51333 ( \51710 , \51707 , \51704 );
xor \U$51334 ( \51711 , \51082 , \51089 );
xor \U$51335 ( \51712 , \51711 , \51097 );
nor \U$51336 ( \51713 , \51710 , \51712 );
nor \U$51337 ( \51714 , \51709 , \51713 );
nand \U$51338 ( \51715 , RIae77630_80, \670 );
and \U$51339 ( \51716 , \51715 , \588 );
not \U$51340 ( \51717 , \51715 );
and \U$51341 ( \51718 , \51717 , \587 );
nor \U$51342 ( \51719 , \51716 , \51718 );
not \U$51343 ( \51720 , \787 );
and \U$51344 ( \51721 , \883 , RIae77540_78);
and \U$51345 ( \51722 , RIae776a8_81, \881 );
nor \U$51346 ( \51723 , \51721 , \51722 );
not \U$51347 ( \51724 , \51723 );
or \U$51348 ( \51725 , \51720 , \51724 );
or \U$51349 ( \51726 , \51723 , \789 );
nand \U$51350 ( \51727 , \51725 , \51726 );
xor \U$51351 ( \51728 , \51719 , \51727 );
xor \U$51352 ( \51729 , \51294 , \51301 );
xor \U$51353 ( \51730 , \51729 , \51309 );
and \U$51354 ( \51731 , \51728 , \51730 );
and \U$51355 ( \51732 , \51719 , \51727 );
nor \U$51356 ( \51733 , \51731 , \51732 );
xor \U$51357 ( \51734 , \51714 , \51733 );
xor \U$51358 ( \51735 , \51209 , \51216 );
xor \U$51359 ( \51736 , \51735 , \51224 );
xor \U$51360 ( \51737 , \51138 , \51145 );
xor \U$51361 ( \51738 , \51737 , \51153 );
and \U$51362 ( \51739 , \51736 , \51738 );
not \U$51363 ( \51740 , \51107 );
xor \U$51364 ( \51741 , \51125 , \51115 );
not \U$51365 ( \51742 , \51741 );
or \U$51366 ( \51743 , \51740 , \51742 );
or \U$51367 ( \51744 , \51741 , \51107 );
nand \U$51368 ( \51745 , \51743 , \51744 );
xor \U$51369 ( \51746 , \51138 , \51145 );
xor \U$51370 ( \51747 , \51746 , \51153 );
and \U$51371 ( \51748 , \51745 , \51747 );
and \U$51372 ( \51749 , \51736 , \51745 );
or \U$51373 ( \51750 , \51739 , \51748 , \51749 );
not \U$51374 ( \51751 , \51750 );
and \U$51375 ( \51752 , \51734 , \51751 );
and \U$51376 ( \51753 , \51714 , \51733 );
or \U$51377 ( \51754 , \51752 , \51753 );
xor \U$51378 ( \51755 , \51702 , \51754 );
not \U$51379 ( \51756 , \51024 );
not \U$51380 ( \51757 , \51030 );
or \U$51381 ( \51758 , \51756 , \51757 );
or \U$51382 ( \51759 , \51024 , \51030 );
nand \U$51383 ( \51760 , \51758 , \51759 );
not \U$51384 ( \51761 , \51760 );
not \U$51385 ( \51762 , \51022 );
and \U$51386 ( \51763 , \51761 , \51762 );
and \U$51387 ( \51764 , \51760 , \51022 );
nor \U$51388 ( \51765 , \51763 , \51764 );
xor \U$51389 ( \51766 , \50760 , \50767 );
xor \U$51390 ( \51767 , \51766 , \50775 );
xor \U$51391 ( \51768 , \51765 , \51767 );
not \U$51392 ( \51769 , \51058 );
not \U$51393 ( \51770 , \51070 );
or \U$51394 ( \51771 , \51769 , \51770 );
or \U$51395 ( \51772 , \51058 , \51070 );
nand \U$51396 ( \51773 , \51771 , \51772 );
not \U$51397 ( \51774 , \51773 );
not \U$51398 ( \51775 , \51060 );
and \U$51399 ( \51776 , \51774 , \51775 );
and \U$51400 ( \51777 , \51773 , \51060 );
nor \U$51401 ( \51778 , \51776 , \51777 );
and \U$51402 ( \51779 , \51768 , \51778 );
and \U$51403 ( \51780 , \51765 , \51767 );
or \U$51404 ( \51781 , \51779 , \51780 );
and \U$51405 ( \51782 , \51755 , \51781 );
and \U$51406 ( \51783 , \51702 , \51754 );
nor \U$51407 ( \51784 , \51782 , \51783 );
xor \U$51408 ( \51785 , \51458 , \51784 );
xor \U$51409 ( \51786 , \51158 , \51230 );
xor \U$51410 ( \51787 , \51786 , \51314 );
xor \U$51411 ( \51788 , \51032 , \51055 );
xor \U$51412 ( \51789 , \51788 , \51072 );
and \U$51413 ( \51790 , \51787 , \51789 );
xor \U$51414 ( \51791 , \50663 , \50665 );
xor \U$51415 ( \51792 , \51791 , \50668 );
xor \U$51416 ( \51793 , \51320 , \51327 );
xor \U$51417 ( \51794 , \51792 , \51793 );
xor \U$51418 ( \51795 , \51032 , \51055 );
xor \U$51419 ( \51796 , \51795 , \51072 );
and \U$51420 ( \51797 , \51794 , \51796 );
and \U$51421 ( \51798 , \51787 , \51794 );
or \U$51422 ( \51799 , \51790 , \51797 , \51798 );
and \U$51423 ( \51800 , \51785 , \51799 );
and \U$51424 ( \51801 , \51458 , \51784 );
or \U$51425 ( \51802 , \51800 , \51801 );
xor \U$51426 ( \51803 , \51422 , \51802 );
not \U$51427 ( \51804 , \51385 );
xnor \U$51428 ( \51805 , \51382 , \51380 );
not \U$51429 ( \51806 , \51805 );
or \U$51430 ( \51807 , \51804 , \51806 );
or \U$51431 ( \51808 , \51805 , \51385 );
nand \U$51432 ( \51809 , \51807 , \51808 );
and \U$51433 ( \51810 , \51803 , \51809 );
and \U$51434 ( \51811 , \51422 , \51802 );
or \U$51435 ( \51812 , \51810 , \51811 );
not \U$51436 ( \51813 , \51812 );
and \U$51437 ( \51814 , \51408 , \51813 );
and \U$51438 ( \51815 , \51407 , \51812 );
nor \U$51439 ( \51816 , \51814 , \51815 );
not \U$51440 ( \51817 , \51816 );
xor \U$51441 ( \51818 , \50974 , \50976 );
xor \U$51442 ( \51819 , \51818 , \50981 );
xor \U$51443 ( \51820 , \50413 , \50439 );
xor \U$51444 ( \51821 , \51820 , \50520 );
xor \U$51445 ( \51822 , \50624 , \50942 );
xor \U$51446 ( \51823 , \51822 , \50969 );
xor \U$51447 ( \51824 , \51821 , \51823 );
xor \U$51448 ( \51825 , \51819 , \51824 );
not \U$51449 ( \51826 , \51825 );
and \U$51450 ( \51827 , \51817 , \51826 );
and \U$51451 ( \51828 , \51816 , \51825 );
nor \U$51452 ( \51829 , \51827 , \51828 );
not \U$51453 ( \51830 , \51829 );
not \U$51454 ( \51831 , \51426 );
not \U$51455 ( \51832 , \51456 );
or \U$51456 ( \51833 , \51831 , \51832 );
or \U$51457 ( \51834 , \51456 , \51426 );
nand \U$51458 ( \51835 , \51833 , \51834 );
not \U$51459 ( \51836 , \51835 );
not \U$51460 ( \51837 , \51424 );
and \U$51461 ( \51838 , \51836 , \51837 );
and \U$51462 ( \51839 , \51835 , \51424 );
nor \U$51463 ( \51840 , \51838 , \51839 );
xor \U$51464 ( \51841 , \51702 , \51754 );
xor \U$51465 ( \51842 , \51841 , \51781 );
or \U$51466 ( \51843 , \51840 , \51842 );
not \U$51467 ( \51844 , \51842 );
not \U$51468 ( \51845 , \51840 );
or \U$51469 ( \51846 , \51844 , \51845 );
xor \U$51470 ( \51847 , \51032 , \51055 );
xor \U$51471 ( \51848 , \51847 , \51072 );
xor \U$51472 ( \51849 , \51787 , \51794 );
xor \U$51473 ( \51850 , \51848 , \51849 );
nand \U$51474 ( \51851 , \51846 , \51850 );
nand \U$51475 ( \51852 , \51843 , \51851 );
xor \U$51476 ( \51853 , \51165 , \51172 );
xor \U$51477 ( \51854 , \51853 , \51180 );
xor \U$51478 ( \51855 , \51190 , \587 );
xor \U$51479 ( \51856 , \51855 , \51198 );
and \U$51480 ( \51857 , \51854 , \51856 );
xor \U$51481 ( \51858 , \51138 , \51145 );
xor \U$51482 ( \51859 , \51858 , \51153 );
xor \U$51483 ( \51860 , \51736 , \51745 );
xor \U$51484 ( \51861 , \51859 , \51860 );
xor \U$51485 ( \51862 , \51190 , \587 );
xor \U$51486 ( \51863 , \51862 , \51198 );
and \U$51487 ( \51864 , \51861 , \51863 );
and \U$51488 ( \51865 , \51854 , \51861 );
or \U$51489 ( \51866 , \51857 , \51864 , \51865 );
and \U$51490 ( \51867 , \3730 , RIae78170_104);
and \U$51491 ( \51868 , RIae77f90_100, \3728 );
nor \U$51492 ( \51869 , \51867 , \51868 );
and \U$51493 ( \51870 , \51869 , \3732 );
not \U$51494 ( \51871 , \51869 );
and \U$51495 ( \51872 , \51871 , \3422 );
nor \U$51496 ( \51873 , \51870 , \51872 );
not \U$51497 ( \51874 , \2789 );
and \U$51498 ( \51875 , \2783 , RIae77090_68);
and \U$51499 ( \51876 , RIae77270_72, \2781 );
nor \U$51500 ( \51877 , \51875 , \51876 );
not \U$51501 ( \51878 , \51877 );
or \U$51502 ( \51879 , \51874 , \51878 );
or \U$51503 ( \51880 , \51877 , \2789 );
nand \U$51504 ( \51881 , \51879 , \51880 );
xor \U$51505 ( \51882 , \51873 , \51881 );
not \U$51506 ( \51883 , \2774 );
and \U$51507 ( \51884 , \3214 , RIae77360_74);
and \U$51508 ( \51885 , RIae78350_108, \3212 );
nor \U$51509 ( \51886 , \51884 , \51885 );
not \U$51510 ( \51887 , \51886 );
or \U$51511 ( \51888 , \51883 , \51887 );
or \U$51512 ( \51889 , \51886 , \3218 );
nand \U$51513 ( \51890 , \51888 , \51889 );
and \U$51514 ( \51891 , \51882 , \51890 );
and \U$51515 ( \51892 , \51873 , \51881 );
or \U$51516 ( \51893 , \51891 , \51892 );
and \U$51517 ( \51894 , \2607 , RIae76cd0_60);
and \U$51518 ( \51895 , RIae77108_69, \2605 );
nor \U$51519 ( \51896 , \51894 , \51895 );
and \U$51520 ( \51897 , \51896 , \2611 );
not \U$51521 ( \51898 , \51896 );
and \U$51522 ( \51899 , \51898 , \2397 );
nor \U$51523 ( \51900 , \51897 , \51899 );
and \U$51524 ( \51901 , \1939 , RIae77900_86);
and \U$51525 ( \51902 , RIae76fa0_66, \1937 );
nor \U$51526 ( \51903 , \51901 , \51902 );
and \U$51527 ( \51904 , \51903 , \1735 );
not \U$51528 ( \51905 , \51903 );
and \U$51529 ( \51906 , \51905 , \1734 );
nor \U$51530 ( \51907 , \51904 , \51906 );
xor \U$51531 ( \51908 , \51900 , \51907 );
and \U$51532 ( \51909 , \2224 , RIae76eb0_64);
and \U$51533 ( \51910 , RIae76dc0_62, \2222 );
nor \U$51534 ( \51911 , \51909 , \51910 );
and \U$51535 ( \51912 , \51911 , \2061 );
not \U$51536 ( \51913 , \51911 );
and \U$51537 ( \51914 , \51913 , \2060 );
nor \U$51538 ( \51915 , \51912 , \51914 );
and \U$51539 ( \51916 , \51908 , \51915 );
and \U$51540 ( \51917 , \51900 , \51907 );
or \U$51541 ( \51918 , \51916 , \51917 );
xor \U$51542 ( \51919 , \51893 , \51918 );
and \U$51543 ( \51920 , \1593 , RIae779f0_88);
and \U$51544 ( \51921 , RIae77810_84, \1591 );
nor \U$51545 ( \51922 , \51920 , \51921 );
and \U$51546 ( \51923 , \51922 , \1498 );
not \U$51547 ( \51924 , \51922 );
and \U$51548 ( \51925 , \51924 , \1488 );
nor \U$51549 ( \51926 , \51923 , \51925 );
and \U$51550 ( \51927 , \1138 , RIae77540_78);
and \U$51551 ( \51928 , RIae776a8_81, \1136 );
nor \U$51552 ( \51929 , \51927 , \51928 );
and \U$51553 ( \51930 , \51929 , \1012 );
not \U$51554 ( \51931 , \51929 );
and \U$51555 ( \51932 , \51931 , \1142 );
nor \U$51556 ( \51933 , \51930 , \51932 );
xor \U$51557 ( \51934 , \51926 , \51933 );
and \U$51558 ( \51935 , \1376 , RIae77450_76);
and \U$51559 ( \51936 , RIae77ae0_90, \1374 );
nor \U$51560 ( \51937 , \51935 , \51936 );
and \U$51561 ( \51938 , \51937 , \1380 );
not \U$51562 ( \51939 , \51937 );
and \U$51563 ( \51940 , \51939 , \1261 );
nor \U$51564 ( \51941 , \51938 , \51940 );
and \U$51565 ( \51942 , \51934 , \51941 );
and \U$51566 ( \51943 , \51926 , \51933 );
or \U$51567 ( \51944 , \51942 , \51943 );
and \U$51568 ( \51945 , \51919 , \51944 );
and \U$51569 ( \51946 , \51893 , \51918 );
or \U$51570 ( \51947 , \51945 , \51946 );
and \U$51571 ( \51948 , \11470 , RIae75560_10);
and \U$51572 ( \51949 , RIae75830_16, \11468 );
nor \U$51573 ( \51950 , \51948 , \51949 );
and \U$51574 ( \51951 , \51950 , \10936 );
not \U$51575 ( \51952 , \51950 );
and \U$51576 ( \51953 , \51952 , \11474 );
nor \U$51577 ( \51954 , \51951 , \51953 );
and \U$51578 ( \51955 , \9760 , RIae75ec0_30);
and \U$51579 ( \51956 , RIae75ce0_26, \9758 );
nor \U$51580 ( \51957 , \51955 , \51956 );
and \U$51581 ( \51958 , \51957 , \9273 );
not \U$51582 ( \51959 , \51957 );
and \U$51583 ( \51960 , \51959 , \9272 );
nor \U$51584 ( \51961 , \51958 , \51960 );
xor \U$51585 ( \51962 , \51954 , \51961 );
and \U$51586 ( \51963 , \10548 , RIae75dd0_28);
and \U$51587 ( \51964 , RIae75650_12, \10546 );
nor \U$51588 ( \51965 , \51963 , \51964 );
and \U$51589 ( \51966 , \51965 , \10421 );
not \U$51590 ( \51967 , \51965 );
and \U$51591 ( \51968 , \51967 , \10118 );
nor \U$51592 ( \51969 , \51966 , \51968 );
and \U$51593 ( \51970 , \51962 , \51969 );
and \U$51594 ( \51971 , \51954 , \51961 );
or \U$51595 ( \51972 , \51970 , \51971 );
and \U$51596 ( \51973 , \15726 , RIae76640_46);
and \U$51597 ( \51974 , RIae76190_36, RIae7aab0_192);
nor \U$51598 ( \51975 , \51973 , \51974 );
and \U$51599 ( \51976 , \51975 , \14959 );
not \U$51600 ( \51977 , \51975 );
and \U$51601 ( \51978 , \51977 , RIae7aa38_191);
nor \U$51602 ( \51979 , \51976 , \51978 );
xor \U$51603 ( \51980 , \51979 , \789 );
and \U$51604 ( \51981 , \14964 , RIae76550_44);
and \U$51605 ( \51982 , RIae76730_48, \14962 );
nor \U$51606 ( \51983 , \51981 , \51982 );
and \U$51607 ( \51984 , \51983 , \14463 );
not \U$51608 ( \51985 , \51983 );
and \U$51609 ( \51986 , \51985 , \14462 );
nor \U$51610 ( \51987 , \51984 , \51986 );
and \U$51611 ( \51988 , \51980 , \51987 );
and \U$51612 ( \51989 , \51979 , \789 );
or \U$51613 ( \51990 , \51988 , \51989 );
xor \U$51614 ( \51991 , \51972 , \51990 );
and \U$51615 ( \51992 , \12180 , RIae75740_14);
and \U$51616 ( \51993 , RIae75290_4, \12178 );
nor \U$51617 ( \51994 , \51992 , \51993 );
and \U$51618 ( \51995 , \51994 , \12184 );
not \U$51619 ( \51996 , \51994 );
and \U$51620 ( \51997 , \51996 , \11827 );
nor \U$51621 ( \51998 , \51995 , \51997 );
and \U$51622 ( \51999 , \13059 , RIae751a0_2);
and \U$51623 ( \52000 , RIae75380_6, \13057 );
nor \U$51624 ( \52001 , \51999 , \52000 );
and \U$51625 ( \52002 , \52001 , \13063 );
not \U$51626 ( \52003 , \52001 );
and \U$51627 ( \52004 , \52003 , \12718 );
nor \U$51628 ( \52005 , \52002 , \52004 );
xor \U$51629 ( \52006 , \51998 , \52005 );
and \U$51630 ( \52007 , \14059 , RIae75470_8);
and \U$51631 ( \52008 , RIae76460_42, \14057 );
nor \U$51632 ( \52009 , \52007 , \52008 );
and \U$51633 ( \52010 , \52009 , \13502 );
not \U$51634 ( \52011 , \52009 );
and \U$51635 ( \52012 , \52011 , \14063 );
nor \U$51636 ( \52013 , \52010 , \52012 );
and \U$51637 ( \52014 , \52006 , \52013 );
and \U$51638 ( \52015 , \51998 , \52005 );
or \U$51639 ( \52016 , \52014 , \52015 );
and \U$51640 ( \52017 , \51991 , \52016 );
and \U$51641 ( \52018 , \51972 , \51990 );
or \U$51642 ( \52019 , \52017 , \52018 );
xor \U$51643 ( \52020 , \51947 , \52019 );
and \U$51644 ( \52021 , \5896 , RIae77bd0_92);
and \U$51645 ( \52022 , RIae77db0_96, \5894 );
nor \U$51646 ( \52023 , \52021 , \52022 );
and \U$51647 ( \52024 , \52023 , \5590 );
not \U$51648 ( \52025 , \52023 );
and \U$51649 ( \52026 , \52025 , \5589 );
nor \U$51650 ( \52027 , \52024 , \52026 );
and \U$51651 ( \52028 , \6172 , RIae77ea0_98);
and \U$51652 ( \52029 , RIae789e0_122, \6170 );
nor \U$51653 ( \52030 , \52028 , \52029 );
and \U$51654 ( \52031 , \52030 , \6176 );
not \U$51655 ( \52032 , \52030 );
and \U$51656 ( \52033 , \52032 , \6175 );
nor \U$51657 ( \52034 , \52031 , \52033 );
xor \U$51658 ( \52035 , \52027 , \52034 );
and \U$51659 ( \52036 , \6941 , RIae788f0_120);
and \U$51660 ( \52037 , RIae78800_118, \6939 );
nor \U$51661 ( \52038 , \52036 , \52037 );
and \U$51662 ( \52039 , \52038 , \6314 );
not \U$51663 ( \52040 , \52038 );
and \U$51664 ( \52041 , \52040 , \6945 );
nor \U$51665 ( \52042 , \52039 , \52041 );
and \U$51666 ( \52043 , \52035 , \52042 );
and \U$51667 ( \52044 , \52027 , \52034 );
or \U$51668 ( \52045 , \52043 , \52044 );
and \U$51669 ( \52046 , \5399 , RIae784b8_111);
and \U$51670 ( \52047 , RIae77cc0_94, \5397 );
nor \U$51671 ( \52048 , \52046 , \52047 );
and \U$51672 ( \52049 , \52048 , \5016 );
not \U$51673 ( \52050 , \52048 );
and \U$51674 ( \52051 , \52050 , \5403 );
nor \U$51675 ( \52052 , \52049 , \52051 );
and \U$51676 ( \52053 , \4247 , RIae78080_102);
and \U$51677 ( \52054 , RIae78260_106, \4245 );
nor \U$51678 ( \52055 , \52053 , \52054 );
and \U$51679 ( \52056 , \52055 , \3989 );
not \U$51680 ( \52057 , \52055 );
and \U$51681 ( \52058 , \52057 , \4251 );
nor \U$51682 ( \52059 , \52056 , \52058 );
xor \U$51683 ( \52060 , \52052 , \52059 );
and \U$51684 ( \52061 , \4688 , RIae78620_114);
and \U$51685 ( \52062 , RIae78440_110, \4686 );
nor \U$51686 ( \52063 , \52061 , \52062 );
and \U$51687 ( \52064 , \52063 , \4481 );
not \U$51688 ( \52065 , \52063 );
and \U$51689 ( \52066 , \52065 , \4482 );
nor \U$51690 ( \52067 , \52064 , \52066 );
and \U$51691 ( \52068 , \52060 , \52067 );
and \U$51692 ( \52069 , \52052 , \52059 );
or \U$51693 ( \52070 , \52068 , \52069 );
xor \U$51694 ( \52071 , \52045 , \52070 );
and \U$51695 ( \52072 , \8966 , RIae75920_18);
and \U$51696 ( \52073 , RIae75fb0_32, \8964 );
nor \U$51697 ( \52074 , \52072 , \52073 );
and \U$51698 ( \52075 , \52074 , \8799 );
not \U$51699 ( \52076 , \52074 );
and \U$51700 ( \52077 , \52076 , \8789 );
nor \U$51701 ( \52078 , \52075 , \52077 );
and \U$51702 ( \52079 , \7633 , RIae78710_116);
and \U$51703 ( \52080 , RIae75bf0_24, \7631 );
nor \U$51704 ( \52081 , \52079 , \52080 );
and \U$51705 ( \52082 , \52081 , \7206 );
not \U$51706 ( \52083 , \52081 );
and \U$51707 ( \52084 , \52083 , \7205 );
nor \U$51708 ( \52085 , \52082 , \52084 );
xor \U$51709 ( \52086 , \52078 , \52085 );
and \U$51710 ( \52087 , \8371 , RIae75b00_22);
and \U$51711 ( \52088 , RIae75a10_20, \8369 );
nor \U$51712 ( \52089 , \52087 , \52088 );
and \U$51713 ( \52090 , \52089 , \8020 );
not \U$51714 ( \52091 , \52089 );
and \U$51715 ( \52092 , \52091 , \8019 );
nor \U$51716 ( \52093 , \52090 , \52092 );
and \U$51717 ( \52094 , \52086 , \52093 );
and \U$51718 ( \52095 , \52078 , \52085 );
or \U$51719 ( \52096 , \52094 , \52095 );
and \U$51720 ( \52097 , \52071 , \52096 );
and \U$51721 ( \52098 , \52045 , \52070 );
or \U$51722 ( \52099 , \52097 , \52098 );
and \U$51723 ( \52100 , \52020 , \52099 );
and \U$51724 ( \52101 , \51947 , \52019 );
or \U$51725 ( \52102 , \52100 , \52101 );
xor \U$51726 ( \52103 , \51866 , \52102 );
xor \U$51727 ( \52104 , \51572 , \51579 );
xor \U$51728 ( \52105 , \52104 , \51587 );
xor \U$51729 ( \52106 , \51598 , \51605 );
xor \U$51730 ( \52107 , \52106 , \51613 );
xor \U$51731 ( \52108 , \52105 , \52107 );
xor \U$51732 ( \52109 , \51547 , \51554 );
xor \U$51733 ( \52110 , \52109 , \51562 );
and \U$51734 ( \52111 , \52108 , \52110 );
and \U$51735 ( \52112 , \52105 , \52107 );
or \U$51736 ( \52113 , \52111 , \52112 );
xor \U$51737 ( \52114 , \51492 , \51500 );
xor \U$51738 ( \52115 , \52114 , \51508 );
xor \U$51739 ( \52116 , \51466 , \51473 );
xor \U$51740 ( \52117 , \52116 , \51482 );
and \U$51741 ( \52118 , \52115 , \52117 );
xor \U$51742 ( \52119 , \51519 , \51526 );
xor \U$51743 ( \52120 , \52119 , \51534 );
xor \U$51744 ( \52121 , \51466 , \51473 );
xor \U$51745 ( \52122 , \52121 , \51482 );
and \U$51746 ( \52123 , \52120 , \52122 );
and \U$51747 ( \52124 , \52115 , \52120 );
or \U$51748 ( \52125 , \52118 , \52123 , \52124 );
xor \U$51749 ( \52126 , \52113 , \52125 );
xor \U$51750 ( \52127 , \51652 , \51659 );
xor \U$51751 ( \52128 , \52127 , \51667 );
xor \U$51752 ( \52129 , \51627 , \51634 );
xor \U$51753 ( \52130 , \52129 , \51642 );
and \U$51754 ( \52131 , \52128 , \52130 );
xor \U$51755 ( \52132 , \51678 , \51685 );
xor \U$51756 ( \52133 , \52132 , \51693 );
xor \U$51757 ( \52134 , \51627 , \51634 );
xor \U$51758 ( \52135 , \52134 , \51642 );
and \U$51759 ( \52136 , \52133 , \52135 );
and \U$51760 ( \52137 , \52128 , \52133 );
or \U$51761 ( \52138 , \52131 , \52136 , \52137 );
and \U$51762 ( \52139 , \52126 , \52138 );
and \U$51763 ( \52140 , \52113 , \52125 );
or \U$51764 ( \52141 , \52139 , \52140 );
and \U$51765 ( \52142 , \52103 , \52141 );
and \U$51766 ( \52143 , \51866 , \52102 );
or \U$51767 ( \52144 , \52142 , \52143 );
xor \U$51768 ( \52145 , \51183 , \51201 );
xor \U$51769 ( \52146 , \52145 , \51227 );
not \U$51770 ( \52147 , \52146 );
xor \U$51771 ( \52148 , \51645 , \51670 );
xor \U$51772 ( \52149 , \52148 , \51696 );
xor \U$51773 ( \52150 , \51565 , \51590 );
xor \U$51774 ( \52151 , \52150 , \51616 );
and \U$51775 ( \52152 , \52149 , \52151 );
not \U$51776 ( \52153 , \52152 );
or \U$51777 ( \52154 , \52147 , \52153 );
or \U$51778 ( \52155 , \52152 , \52146 );
xor \U$51779 ( \52156 , \51485 , \51511 );
xor \U$51780 ( \52157 , \52156 , \51537 );
xor \U$51781 ( \52158 , \51719 , \51727 );
xor \U$51782 ( \52159 , \52158 , \51730 );
xor \U$51783 ( \52160 , \52157 , \52159 );
not \U$51784 ( \52161 , \51704 );
xor \U$51785 ( \52162 , \51707 , \51712 );
not \U$51786 ( \52163 , \52162 );
or \U$51787 ( \52164 , \52161 , \52163 );
or \U$51788 ( \52165 , \52162 , \51704 );
nand \U$51789 ( \52166 , \52164 , \52165 );
and \U$51790 ( \52167 , \52160 , \52166 );
and \U$51791 ( \52168 , \52157 , \52159 );
or \U$51792 ( \52169 , \52167 , \52168 );
nand \U$51793 ( \52170 , \52155 , \52169 );
nand \U$51794 ( \52171 , \52154 , \52170 );
xor \U$51795 ( \52172 , \52144 , \52171 );
xor \U$51796 ( \52173 , \51714 , \51733 );
xor \U$51797 ( \52174 , \52173 , \51751 );
xor \U$51798 ( \52175 , \51440 , \51450 );
xor \U$51799 ( \52176 , \52175 , \51453 );
xor \U$51800 ( \52177 , \52174 , \52176 );
xor \U$51801 ( \52178 , \51765 , \51767 );
xor \U$51802 ( \52179 , \52178 , \51778 );
and \U$51803 ( \52180 , \52177 , \52179 );
and \U$51804 ( \52181 , \52174 , \52176 );
nor \U$51805 ( \52182 , \52180 , \52181 );
and \U$51806 ( \52183 , \52172 , \52182 );
and \U$51807 ( \52184 , \52144 , \52171 );
or \U$51808 ( \52185 , \52183 , \52184 );
xor \U$51809 ( \52186 , \51852 , \52185 );
xor \U$51810 ( \52187 , \51362 , \51364 );
xor \U$51811 ( \52188 , \52187 , \51369 );
xor \U$51812 ( \52189 , \51410 , \51417 );
xor \U$51813 ( \52190 , \52188 , \52189 );
and \U$51814 ( \52191 , \52186 , \52190 );
and \U$51815 ( \52192 , \51852 , \52185 );
or \U$51816 ( \52193 , \52191 , \52192 );
xor \U$51817 ( \52194 , \51020 , \51335 );
xor \U$51818 ( \52195 , \52194 , \51372 );
xor \U$51819 ( \52196 , \52193 , \52195 );
xor \U$51820 ( \52197 , \51422 , \51802 );
xor \U$51821 ( \52198 , \52197 , \51809 );
and \U$51822 ( \52199 , \52196 , \52198 );
and \U$51823 ( \52200 , \52193 , \52195 );
or \U$51824 ( \52201 , \52199 , \52200 );
not \U$51825 ( \52202 , \52201 );
and \U$51826 ( \52203 , \51830 , \52202 );
and \U$51827 ( \52204 , \51829 , \52201 );
nor \U$51828 ( \52205 , \52203 , \52204 );
xor \U$51829 ( \52206 , \51852 , \52185 );
xor \U$51830 ( \52207 , \52206 , \52190 );
xor \U$51831 ( \52208 , \51458 , \51784 );
xor \U$51832 ( \52209 , \52208 , \51799 );
xor \U$51833 ( \52210 , \52207 , \52209 );
xnor \U$51834 ( \52211 , \51842 , \51840 );
not \U$51835 ( \52212 , \52211 );
not \U$51836 ( \52213 , \51850 );
and \U$51837 ( \52214 , \52212 , \52213 );
and \U$51838 ( \52215 , \52211 , \51850 );
nor \U$51839 ( \52216 , \52214 , \52215 );
xor \U$51840 ( \52217 , \51947 , \52019 );
xor \U$51841 ( \52218 , \52217 , \52099 );
xor \U$51842 ( \52219 , \51190 , \587 );
xor \U$51843 ( \52220 , \52219 , \51198 );
xor \U$51844 ( \52221 , \51854 , \51861 );
xor \U$51845 ( \52222 , \52220 , \52221 );
xor \U$51846 ( \52223 , \52218 , \52222 );
xor \U$51847 ( \52224 , \52113 , \52125 );
xor \U$51848 ( \52225 , \52224 , \52138 );
and \U$51849 ( \52226 , \52223 , \52225 );
and \U$51850 ( \52227 , \52218 , \52222 );
or \U$51851 ( \52228 , \52226 , \52227 );
xor \U$51852 ( \52229 , \52052 , \52059 );
xor \U$51853 ( \52230 , \52229 , \52067 );
xor \U$51854 ( \52231 , \51873 , \51881 );
xor \U$51855 ( \52232 , \52231 , \51890 );
and \U$51856 ( \52233 , \52230 , \52232 );
xor \U$51857 ( \52234 , \52027 , \52034 );
xor \U$51858 ( \52235 , \52234 , \52042 );
xor \U$51859 ( \52236 , \51873 , \51881 );
xor \U$51860 ( \52237 , \52236 , \51890 );
and \U$51861 ( \52238 , \52235 , \52237 );
and \U$51862 ( \52239 , \52230 , \52235 );
or \U$51863 ( \52240 , \52233 , \52238 , \52239 );
nand \U$51864 ( \52241 , RIae77630_80, \881 );
not \U$51865 ( \52242 , \52241 );
not \U$51866 ( \52243 , \787 );
or \U$51867 ( \52244 , \52242 , \52243 );
or \U$51868 ( \52245 , \787 , \52241 );
nand \U$51869 ( \52246 , \52244 , \52245 );
xor \U$51870 ( \52247 , \51926 , \51933 );
xor \U$51871 ( \52248 , \52247 , \51941 );
and \U$51872 ( \52249 , \52246 , \52248 );
xor \U$51873 ( \52250 , \51900 , \51907 );
xor \U$51874 ( \52251 , \52250 , \51915 );
xor \U$51875 ( \52252 , \51926 , \51933 );
xor \U$51876 ( \52253 , \52252 , \51941 );
and \U$51877 ( \52254 , \52251 , \52253 );
and \U$51878 ( \52255 , \52246 , \52251 );
or \U$51879 ( \52256 , \52249 , \52254 , \52255 );
xor \U$51880 ( \52257 , \52240 , \52256 );
xor \U$51881 ( \52258 , \52078 , \52085 );
xor \U$51882 ( \52259 , \52258 , \52093 );
xor \U$51883 ( \52260 , \51954 , \51961 );
xor \U$51884 ( \52261 , \52260 , \51969 );
xor \U$51885 ( \52262 , \52259 , \52261 );
xor \U$51886 ( \52263 , \51998 , \52005 );
xor \U$51887 ( \52264 , \52263 , \52013 );
and \U$51888 ( \52265 , \52262 , \52264 );
and \U$51889 ( \52266 , \52259 , \52261 );
or \U$51890 ( \52267 , \52265 , \52266 );
and \U$51891 ( \52268 , \52257 , \52267 );
and \U$51892 ( \52269 , \52240 , \52256 );
or \U$51893 ( \52270 , \52268 , \52269 );
and \U$51894 ( \52271 , \1593 , RIae77ae0_90);
and \U$51895 ( \52272 , RIae779f0_88, \1591 );
nor \U$51896 ( \52273 , \52271 , \52272 );
and \U$51897 ( \52274 , \52273 , \1488 );
not \U$51898 ( \52275 , \52273 );
and \U$51899 ( \52276 , \52275 , \1498 );
nor \U$51900 ( \52277 , \52274 , \52276 );
and \U$51901 ( \52278 , \2224 , RIae76fa0_66);
and \U$51902 ( \52279 , RIae76eb0_64, \2222 );
nor \U$51903 ( \52280 , \52278 , \52279 );
and \U$51904 ( \52281 , \52280 , \2060 );
not \U$51905 ( \52282 , \52280 );
and \U$51906 ( \52283 , \52282 , \2061 );
nor \U$51907 ( \52284 , \52281 , \52283 );
or \U$51908 ( \52285 , \52277 , \52284 );
not \U$51909 ( \52286 , \52284 );
not \U$51910 ( \52287 , \52277 );
or \U$51911 ( \52288 , \52286 , \52287 );
and \U$51912 ( \52289 , \1939 , RIae77810_84);
and \U$51913 ( \52290 , RIae77900_86, \1937 );
nor \U$51914 ( \52291 , \52289 , \52290 );
and \U$51915 ( \52292 , \52291 , \1735 );
not \U$51916 ( \52293 , \52291 );
and \U$51917 ( \52294 , \52293 , \1734 );
nor \U$51918 ( \52295 , \52292 , \52294 );
nand \U$51919 ( \52296 , \52288 , \52295 );
nand \U$51920 ( \52297 , \52285 , \52296 );
and \U$51921 ( \52298 , \1376 , RIae776a8_81);
and \U$51922 ( \52299 , RIae77450_76, \1374 );
nor \U$51923 ( \52300 , \52298 , \52299 );
and \U$51924 ( \52301 , \52300 , \1380 );
not \U$51925 ( \52302 , \52300 );
and \U$51926 ( \52303 , \52302 , \1261 );
nor \U$51927 ( \52304 , \52301 , \52303 );
and \U$51928 ( \52305 , \1138 , RIae77630_80);
and \U$51929 ( \52306 , RIae77540_78, \1136 );
nor \U$51930 ( \52307 , \52305 , \52306 );
and \U$51931 ( \52308 , \52307 , \1012 );
not \U$51932 ( \52309 , \52307 );
and \U$51933 ( \52310 , \52309 , \1142 );
nor \U$51934 ( \52311 , \52308 , \52310 );
and \U$51935 ( \52312 , \52304 , \52311 );
xor \U$51936 ( \52313 , \52297 , \52312 );
and \U$51937 ( \52314 , \2607 , RIae76dc0_62);
and \U$51938 ( \52315 , RIae76cd0_60, \2605 );
nor \U$51939 ( \52316 , \52314 , \52315 );
and \U$51940 ( \52317 , \52316 , \2611 );
not \U$51941 ( \52318 , \52316 );
and \U$51942 ( \52319 , \52318 , \2397 );
nor \U$51943 ( \52320 , \52317 , \52319 );
not \U$51944 ( \52321 , \2789 );
and \U$51945 ( \52322 , \2783 , RIae77108_69);
and \U$51946 ( \52323 , RIae77090_68, \2781 );
nor \U$51947 ( \52324 , \52322 , \52323 );
not \U$51948 ( \52325 , \52324 );
or \U$51949 ( \52326 , \52321 , \52325 );
or \U$51950 ( \52327 , \52324 , \3089 );
nand \U$51951 ( \52328 , \52326 , \52327 );
xor \U$51952 ( \52329 , \52320 , \52328 );
not \U$51953 ( \52330 , \2774 );
and \U$51954 ( \52331 , \3214 , RIae77270_72);
and \U$51955 ( \52332 , RIae77360_74, \3212 );
nor \U$51956 ( \52333 , \52331 , \52332 );
not \U$51957 ( \52334 , \52333 );
or \U$51958 ( \52335 , \52330 , \52334 );
or \U$51959 ( \52336 , \52333 , \3218 );
nand \U$51960 ( \52337 , \52335 , \52336 );
and \U$51961 ( \52338 , \52329 , \52337 );
and \U$51962 ( \52339 , \52320 , \52328 );
or \U$51963 ( \52340 , \52338 , \52339 );
and \U$51964 ( \52341 , \52313 , \52340 );
and \U$51965 ( \52342 , \52297 , \52312 );
or \U$51966 ( \52343 , \52341 , \52342 );
and \U$51967 ( \52344 , \12180 , RIae75830_16);
and \U$51968 ( \52345 , RIae75740_14, \12178 );
nor \U$51969 ( \52346 , \52344 , \52345 );
and \U$51970 ( \52347 , \52346 , \11827 );
not \U$51971 ( \52348 , \52346 );
and \U$51972 ( \52349 , \52348 , \12184 );
nor \U$51973 ( \52350 , \52347 , \52349 );
and \U$51974 ( \52351 , \13059 , RIae75290_4);
and \U$51975 ( \52352 , RIae751a0_2, \13057 );
nor \U$51976 ( \52353 , \52351 , \52352 );
and \U$51977 ( \52354 , \52353 , \12718 );
not \U$51978 ( \52355 , \52353 );
and \U$51979 ( \52356 , \52355 , \13063 );
nor \U$51980 ( \52357 , \52354 , \52356 );
xor \U$51981 ( \52358 , \52350 , \52357 );
and \U$51982 ( \52359 , \11470 , RIae75650_12);
and \U$51983 ( \52360 , RIae75560_10, \11468 );
nor \U$51984 ( \52361 , \52359 , \52360 );
and \U$51985 ( \52362 , \52361 , \11474 );
not \U$51986 ( \52363 , \52361 );
and \U$51987 ( \52364 , \52363 , \10936 );
nor \U$51988 ( \52365 , \52362 , \52364 );
and \U$51989 ( \52366 , \52358 , \52365 );
and \U$51990 ( \52367 , \52350 , \52357 );
nor \U$51991 ( \52368 , \52366 , \52367 );
and \U$51992 ( \52369 , \14059 , RIae75380_6);
and \U$51993 ( \52370 , RIae75470_8, \14057 );
nor \U$51994 ( \52371 , \52369 , \52370 );
and \U$51995 ( \52372 , \52371 , \13502 );
not \U$51996 ( \52373 , \52371 );
and \U$51997 ( \52374 , \52373 , \14063 );
nor \U$51998 ( \52375 , \52372 , \52374 );
and \U$51999 ( \52376 , \15726 , RIae76730_48);
and \U$52000 ( \52377 , RIae76640_46, RIae7aab0_192);
nor \U$52001 ( \52378 , \52376 , \52377 );
and \U$52002 ( \52379 , \52378 , \14959 );
not \U$52003 ( \52380 , \52378 );
and \U$52004 ( \52381 , \52380 , RIae7aa38_191);
nor \U$52005 ( \52382 , \52379 , \52381 );
xor \U$52006 ( \52383 , \52375 , \52382 );
and \U$52007 ( \52384 , \14964 , RIae76460_42);
and \U$52008 ( \52385 , RIae76550_44, \14962 );
nor \U$52009 ( \52386 , \52384 , \52385 );
and \U$52010 ( \52387 , \52386 , \14463 );
not \U$52011 ( \52388 , \52386 );
and \U$52012 ( \52389 , \52388 , \14462 );
nor \U$52013 ( \52390 , \52387 , \52389 );
and \U$52014 ( \52391 , \52383 , \52390 );
and \U$52015 ( \52392 , \52375 , \52382 );
or \U$52016 ( \52393 , \52391 , \52392 );
xor \U$52017 ( \52394 , \52368 , \52393 );
and \U$52018 ( \52395 , \8966 , RIae75a10_20);
and \U$52019 ( \52396 , RIae75920_18, \8964 );
nor \U$52020 ( \52397 , \52395 , \52396 );
and \U$52021 ( \52398 , \52397 , \8789 );
not \U$52022 ( \52399 , \52397 );
and \U$52023 ( \52400 , \52399 , \8799 );
nor \U$52024 ( \52401 , \52398 , \52400 );
and \U$52025 ( \52402 , \9760 , RIae75fb0_32);
and \U$52026 ( \52403 , RIae75ec0_30, \9758 );
nor \U$52027 ( \52404 , \52402 , \52403 );
and \U$52028 ( \52405 , \52404 , \9272 );
not \U$52029 ( \52406 , \52404 );
and \U$52030 ( \52407 , \52406 , \9273 );
nor \U$52031 ( \52408 , \52405 , \52407 );
or \U$52032 ( \52409 , \52401 , \52408 );
not \U$52033 ( \52410 , \52408 );
not \U$52034 ( \52411 , \52401 );
or \U$52035 ( \52412 , \52410 , \52411 );
and \U$52036 ( \52413 , \10548 , RIae75ce0_26);
and \U$52037 ( \52414 , RIae75dd0_28, \10546 );
nor \U$52038 ( \52415 , \52413 , \52414 );
and \U$52039 ( \52416 , \52415 , \10421 );
not \U$52040 ( \52417 , \52415 );
and \U$52041 ( \52418 , \52417 , \10118 );
nor \U$52042 ( \52419 , \52416 , \52418 );
nand \U$52043 ( \52420 , \52412 , \52419 );
nand \U$52044 ( \52421 , \52409 , \52420 );
and \U$52045 ( \52422 , \52394 , \52421 );
and \U$52046 ( \52423 , \52368 , \52393 );
or \U$52047 ( \52424 , \52422 , \52423 );
xor \U$52048 ( \52425 , \52343 , \52424 );
and \U$52049 ( \52426 , \5399 , RIae78440_110);
and \U$52050 ( \52427 , RIae784b8_111, \5397 );
nor \U$52051 ( \52428 , \52426 , \52427 );
and \U$52052 ( \52429 , \52428 , \5403 );
not \U$52053 ( \52430 , \52428 );
and \U$52054 ( \52431 , \52430 , \5016 );
nor \U$52055 ( \52432 , \52429 , \52431 );
and \U$52056 ( \52433 , \6172 , RIae77db0_96);
and \U$52057 ( \52434 , RIae77ea0_98, \6170 );
nor \U$52058 ( \52435 , \52433 , \52434 );
and \U$52059 ( \52436 , \52435 , \6175 );
not \U$52060 ( \52437 , \52435 );
and \U$52061 ( \52438 , \52437 , \6176 );
nor \U$52062 ( \52439 , \52436 , \52438 );
or \U$52063 ( \52440 , \52432 , \52439 );
not \U$52064 ( \52441 , \52439 );
not \U$52065 ( \52442 , \52432 );
or \U$52066 ( \52443 , \52441 , \52442 );
and \U$52067 ( \52444 , \5896 , RIae77cc0_94);
and \U$52068 ( \52445 , RIae77bd0_92, \5894 );
nor \U$52069 ( \52446 , \52444 , \52445 );
and \U$52070 ( \52447 , \52446 , \5590 );
not \U$52071 ( \52448 , \52446 );
and \U$52072 ( \52449 , \52448 , \5589 );
nor \U$52073 ( \52450 , \52447 , \52449 );
nand \U$52074 ( \52451 , \52443 , \52450 );
nand \U$52075 ( \52452 , \52440 , \52451 );
and \U$52076 ( \52453 , \3730 , RIae78350_108);
and \U$52077 ( \52454 , RIae78170_104, \3728 );
nor \U$52078 ( \52455 , \52453 , \52454 );
and \U$52079 ( \52456 , \52455 , \3422 );
not \U$52080 ( \52457 , \52455 );
and \U$52081 ( \52458 , \52457 , \3732 );
nor \U$52082 ( \52459 , \52456 , \52458 );
and \U$52083 ( \52460 , \4688 , RIae78260_106);
and \U$52084 ( \52461 , RIae78620_114, \4686 );
nor \U$52085 ( \52462 , \52460 , \52461 );
and \U$52086 ( \52463 , \52462 , \4482 );
not \U$52087 ( \52464 , \52462 );
and \U$52088 ( \52465 , \52464 , \4481 );
nor \U$52089 ( \52466 , \52463 , \52465 );
or \U$52090 ( \52467 , \52459 , \52466 );
not \U$52091 ( \52468 , \52466 );
not \U$52092 ( \52469 , \52459 );
or \U$52093 ( \52470 , \52468 , \52469 );
and \U$52094 ( \52471 , \4247 , RIae77f90_100);
and \U$52095 ( \52472 , RIae78080_102, \4245 );
nor \U$52096 ( \52473 , \52471 , \52472 );
and \U$52097 ( \52474 , \52473 , \3989 );
not \U$52098 ( \52475 , \52473 );
and \U$52099 ( \52476 , \52475 , \4251 );
nor \U$52100 ( \52477 , \52474 , \52476 );
nand \U$52101 ( \52478 , \52470 , \52477 );
nand \U$52102 ( \52479 , \52467 , \52478 );
xor \U$52103 ( \52480 , \52452 , \52479 );
and \U$52104 ( \52481 , \6941 , RIae789e0_122);
and \U$52105 ( \52482 , RIae788f0_120, \6939 );
nor \U$52106 ( \52483 , \52481 , \52482 );
and \U$52107 ( \52484 , \52483 , \6314 );
not \U$52108 ( \52485 , \52483 );
and \U$52109 ( \52486 , \52485 , \6945 );
nor \U$52110 ( \52487 , \52484 , \52486 );
and \U$52111 ( \52488 , \7633 , RIae78800_118);
and \U$52112 ( \52489 , RIae78710_116, \7631 );
nor \U$52113 ( \52490 , \52488 , \52489 );
and \U$52114 ( \52491 , \52490 , \7206 );
not \U$52115 ( \52492 , \52490 );
and \U$52116 ( \52493 , \52492 , \7205 );
nor \U$52117 ( \52494 , \52491 , \52493 );
xor \U$52118 ( \52495 , \52487 , \52494 );
and \U$52119 ( \52496 , \8371 , RIae75bf0_24);
and \U$52120 ( \52497 , RIae75b00_22, \8369 );
nor \U$52121 ( \52498 , \52496 , \52497 );
and \U$52122 ( \52499 , \52498 , \8020 );
not \U$52123 ( \52500 , \52498 );
and \U$52124 ( \52501 , \52500 , \8019 );
nor \U$52125 ( \52502 , \52499 , \52501 );
and \U$52126 ( \52503 , \52495 , \52502 );
and \U$52127 ( \52504 , \52487 , \52494 );
or \U$52128 ( \52505 , \52503 , \52504 );
and \U$52129 ( \52506 , \52480 , \52505 );
and \U$52130 ( \52507 , \52452 , \52479 );
or \U$52131 ( \52508 , \52506 , \52507 );
and \U$52132 ( \52509 , \52425 , \52508 );
and \U$52133 ( \52510 , \52343 , \52424 );
or \U$52134 ( \52511 , \52509 , \52510 );
xor \U$52135 ( \52512 , \52270 , \52511 );
xor \U$52136 ( \52513 , \51466 , \51473 );
xor \U$52137 ( \52514 , \52513 , \51482 );
xor \U$52138 ( \52515 , \52115 , \52120 );
xor \U$52139 ( \52516 , \52514 , \52515 );
xor \U$52140 ( \52517 , \52105 , \52107 );
xor \U$52141 ( \52518 , \52517 , \52110 );
and \U$52142 ( \52519 , \52516 , \52518 );
xor \U$52143 ( \52520 , \51627 , \51634 );
xor \U$52144 ( \52521 , \52520 , \51642 );
xor \U$52145 ( \52522 , \52128 , \52133 );
xor \U$52146 ( \52523 , \52521 , \52522 );
xor \U$52147 ( \52524 , \52105 , \52107 );
xor \U$52148 ( \52525 , \52524 , \52110 );
and \U$52149 ( \52526 , \52523 , \52525 );
and \U$52150 ( \52527 , \52516 , \52523 );
or \U$52151 ( \52528 , \52519 , \52526 , \52527 );
and \U$52152 ( \52529 , \52512 , \52528 );
and \U$52153 ( \52530 , \52270 , \52511 );
or \U$52154 ( \52531 , \52529 , \52530 );
and \U$52155 ( \52532 , \52228 , \52531 );
xor \U$52156 ( \52533 , \52045 , \52070 );
xor \U$52157 ( \52534 , \52533 , \52096 );
xor \U$52158 ( \52535 , \51972 , \51990 );
xor \U$52159 ( \52536 , \52535 , \52016 );
xor \U$52160 ( \52537 , \52534 , \52536 );
xor \U$52161 ( \52538 , \51893 , \51918 );
xor \U$52162 ( \52539 , \52538 , \51944 );
and \U$52163 ( \52540 , \52537 , \52539 );
and \U$52164 ( \52541 , \52534 , \52536 );
or \U$52165 ( \52542 , \52540 , \52541 );
xor \U$52166 ( \52543 , \52149 , \52151 );
xor \U$52167 ( \52544 , \52542 , \52543 );
xor \U$52168 ( \52545 , \52157 , \52159 );
xor \U$52169 ( \52546 , \52545 , \52166 );
and \U$52170 ( \52547 , \52544 , \52546 );
and \U$52171 ( \52548 , \52542 , \52543 );
or \U$52172 ( \52549 , \52547 , \52548 );
or \U$52173 ( \52550 , \52228 , \52531 );
and \U$52174 ( \52551 , \52549 , \52550 );
nor \U$52175 ( \52552 , \52532 , \52551 );
or \U$52176 ( \52553 , \52216 , \52552 );
not \U$52177 ( \52554 , \52552 );
not \U$52178 ( \52555 , \52216 );
or \U$52179 ( \52556 , \52554 , \52555 );
xor \U$52180 ( \52557 , \51540 , \51619 );
xor \U$52181 ( \52558 , \52557 , \51699 );
xnor \U$52182 ( \52559 , \52169 , \52152 );
not \U$52183 ( \52560 , \52559 );
not \U$52184 ( \52561 , \52146 );
and \U$52185 ( \52562 , \52560 , \52561 );
and \U$52186 ( \52563 , \52559 , \52146 );
nor \U$52187 ( \52564 , \52562 , \52563 );
xor \U$52188 ( \52565 , \52558 , \52564 );
xor \U$52189 ( \52566 , \52174 , \52176 );
xor \U$52190 ( \52567 , \52566 , \52179 );
and \U$52191 ( \52568 , \52565 , \52567 );
and \U$52192 ( \52569 , \52558 , \52564 );
nor \U$52193 ( \52570 , \52568 , \52569 );
nand \U$52194 ( \52571 , \52556 , \52570 );
nand \U$52195 ( \52572 , \52553 , \52571 );
and \U$52196 ( \52573 , \52210 , \52572 );
and \U$52197 ( \52574 , \52207 , \52209 );
nor \U$52198 ( \52575 , \52573 , \52574 );
not \U$52199 ( \52576 , \52575 );
xor \U$52200 ( \52577 , \52193 , \52195 );
xor \U$52201 ( \52578 , \52577 , \52198 );
nand \U$52202 ( \52579 , \52576 , \52578 );
or \U$52203 ( \52580 , \52205 , \52579 );
xnor \U$52204 ( \52581 , \52579 , \52205 );
xor \U$52205 ( \52582 , \52207 , \52209 );
xor \U$52206 ( \52583 , \52582 , \52572 );
not \U$52207 ( \52584 , \52583 );
xor \U$52208 ( \52585 , \52558 , \52564 );
xor \U$52209 ( \52586 , \52585 , \52567 );
not \U$52210 ( \52587 , \52586 );
not \U$52211 ( \52588 , \52549 );
xnor \U$52212 ( \52589 , \52531 , \52228 );
not \U$52213 ( \52590 , \52589 );
or \U$52214 ( \52591 , \52588 , \52590 );
or \U$52215 ( \52592 , \52589 , \52549 );
nand \U$52216 ( \52593 , \52591 , \52592 );
nand \U$52217 ( \52594 , \52587 , \52593 );
not \U$52218 ( \52595 , \52594 );
xor \U$52219 ( \52596 , \52144 , \52171 );
xor \U$52220 ( \52597 , \52596 , \52182 );
and \U$52221 ( \52598 , \52595 , \52597 );
not \U$52222 ( \52599 , \52597 );
nand \U$52223 ( \52600 , \52599 , \52594 );
not \U$52224 ( \52601 , \52466 );
not \U$52225 ( \52602 , \52477 );
or \U$52226 ( \52603 , \52601 , \52602 );
or \U$52227 ( \52604 , \52466 , \52477 );
nand \U$52228 ( \52605 , \52603 , \52604 );
not \U$52229 ( \52606 , \52605 );
not \U$52230 ( \52607 , \52459 );
and \U$52231 ( \52608 , \52606 , \52607 );
and \U$52232 ( \52609 , \52605 , \52459 );
nor \U$52233 ( \52610 , \52608 , \52609 );
not \U$52234 ( \52611 , \52439 );
not \U$52235 ( \52612 , \52450 );
or \U$52236 ( \52613 , \52611 , \52612 );
or \U$52237 ( \52614 , \52439 , \52450 );
nand \U$52238 ( \52615 , \52613 , \52614 );
not \U$52239 ( \52616 , \52615 );
not \U$52240 ( \52617 , \52432 );
and \U$52241 ( \52618 , \52616 , \52617 );
and \U$52242 ( \52619 , \52615 , \52432 );
nor \U$52243 ( \52620 , \52618 , \52619 );
or \U$52244 ( \52621 , \52610 , \52620 );
not \U$52245 ( \52622 , \52620 );
not \U$52246 ( \52623 , \52610 );
or \U$52247 ( \52624 , \52622 , \52623 );
xor \U$52248 ( \52625 , \52487 , \52494 );
xor \U$52249 ( \52626 , \52625 , \52502 );
nand \U$52250 ( \52627 , \52624 , \52626 );
nand \U$52251 ( \52628 , \52621 , \52627 );
not \U$52252 ( \52629 , \52284 );
not \U$52253 ( \52630 , \52295 );
or \U$52254 ( \52631 , \52629 , \52630 );
or \U$52255 ( \52632 , \52284 , \52295 );
nand \U$52256 ( \52633 , \52631 , \52632 );
not \U$52257 ( \52634 , \52633 );
not \U$52258 ( \52635 , \52277 );
and \U$52259 ( \52636 , \52634 , \52635 );
and \U$52260 ( \52637 , \52633 , \52277 );
nor \U$52261 ( \52638 , \52636 , \52637 );
xor \U$52262 ( \52639 , \52304 , \52311 );
not \U$52263 ( \52640 , \52639 );
or \U$52264 ( \52641 , \52638 , \52640 );
not \U$52265 ( \52642 , \52640 );
not \U$52266 ( \52643 , \52638 );
or \U$52267 ( \52644 , \52642 , \52643 );
xor \U$52268 ( \52645 , \52320 , \52328 );
xor \U$52269 ( \52646 , \52645 , \52337 );
nand \U$52270 ( \52647 , \52644 , \52646 );
nand \U$52271 ( \52648 , \52641 , \52647 );
xor \U$52272 ( \52649 , \52628 , \52648 );
not \U$52273 ( \52650 , \52408 );
not \U$52274 ( \52651 , \52419 );
or \U$52275 ( \52652 , \52650 , \52651 );
or \U$52276 ( \52653 , \52408 , \52419 );
nand \U$52277 ( \52654 , \52652 , \52653 );
not \U$52278 ( \52655 , \52654 );
not \U$52279 ( \52656 , \52401 );
and \U$52280 ( \52657 , \52655 , \52656 );
and \U$52281 ( \52658 , \52654 , \52401 );
nor \U$52282 ( \52659 , \52657 , \52658 );
xor \U$52283 ( \52660 , \52350 , \52357 );
xor \U$52284 ( \52661 , \52660 , \52365 );
or \U$52285 ( \52662 , \52659 , \52661 );
not \U$52286 ( \52663 , \52661 );
not \U$52287 ( \52664 , \52659 );
or \U$52288 ( \52665 , \52663 , \52664 );
xor \U$52289 ( \52666 , \52375 , \52382 );
xor \U$52290 ( \52667 , \52666 , \52390 );
nand \U$52291 ( \52668 , \52665 , \52667 );
nand \U$52292 ( \52669 , \52662 , \52668 );
and \U$52293 ( \52670 , \52649 , \52669 );
and \U$52294 ( \52671 , \52628 , \52648 );
or \U$52295 ( \52672 , \52670 , \52671 );
and \U$52296 ( \52673 , \8371 , RIae78710_116);
and \U$52297 ( \52674 , RIae75bf0_24, \8369 );
nor \U$52298 ( \52675 , \52673 , \52674 );
and \U$52299 ( \52676 , \52675 , \8019 );
not \U$52300 ( \52677 , \52675 );
and \U$52301 ( \52678 , \52677 , \8020 );
nor \U$52302 ( \52679 , \52676 , \52678 );
and \U$52303 ( \52680 , \8966 , RIae75b00_22);
and \U$52304 ( \52681 , RIae75a10_20, \8964 );
nor \U$52305 ( \52682 , \52680 , \52681 );
and \U$52306 ( \52683 , \52682 , \8789 );
not \U$52307 ( \52684 , \52682 );
and \U$52308 ( \52685 , \52684 , \8799 );
nor \U$52309 ( \52686 , \52683 , \52685 );
xor \U$52310 ( \52687 , \52679 , \52686 );
and \U$52311 ( \52688 , \7633 , RIae788f0_120);
and \U$52312 ( \52689 , RIae78800_118, \7631 );
nor \U$52313 ( \52690 , \52688 , \52689 );
and \U$52314 ( \52691 , \52690 , \7205 );
not \U$52315 ( \52692 , \52690 );
and \U$52316 ( \52693 , \52692 , \7206 );
nor \U$52317 ( \52694 , \52691 , \52693 );
and \U$52318 ( \52695 , \52687 , \52694 );
and \U$52319 ( \52696 , \52679 , \52686 );
nor \U$52320 ( \52697 , \52695 , \52696 );
and \U$52321 ( \52698 , \4688 , RIae78080_102);
and \U$52322 ( \52699 , RIae78260_106, \4686 );
nor \U$52323 ( \52700 , \52698 , \52699 );
and \U$52324 ( \52701 , \52700 , \4482 );
not \U$52325 ( \52702 , \52700 );
and \U$52326 ( \52703 , \52702 , \4481 );
nor \U$52327 ( \52704 , \52701 , \52703 );
and \U$52328 ( \52705 , \5399 , RIae78620_114);
and \U$52329 ( \52706 , RIae78440_110, \5397 );
nor \U$52330 ( \52707 , \52705 , \52706 );
and \U$52331 ( \52708 , \52707 , \5403 );
not \U$52332 ( \52709 , \52707 );
and \U$52333 ( \52710 , \52709 , \5016 );
nor \U$52334 ( \52711 , \52708 , \52710 );
xor \U$52335 ( \52712 , \52704 , \52711 );
and \U$52336 ( \52713 , \4247 , RIae78170_104);
and \U$52337 ( \52714 , RIae77f90_100, \4245 );
nor \U$52338 ( \52715 , \52713 , \52714 );
and \U$52339 ( \52716 , \52715 , \4251 );
not \U$52340 ( \52717 , \52715 );
and \U$52341 ( \52718 , \52717 , \3989 );
nor \U$52342 ( \52719 , \52716 , \52718 );
and \U$52343 ( \52720 , \52712 , \52719 );
and \U$52344 ( \52721 , \52704 , \52711 );
nor \U$52345 ( \52722 , \52720 , \52721 );
xor \U$52346 ( \52723 , \52697 , \52722 );
and \U$52347 ( \52724 , \5896 , RIae784b8_111);
and \U$52348 ( \52725 , RIae77cc0_94, \5894 );
nor \U$52349 ( \52726 , \52724 , \52725 );
and \U$52350 ( \52727 , \52726 , \5589 );
not \U$52351 ( \52728 , \52726 );
and \U$52352 ( \52729 , \52728 , \5590 );
nor \U$52353 ( \52730 , \52727 , \52729 );
and \U$52354 ( \52731 , \6172 , RIae77bd0_92);
and \U$52355 ( \52732 , RIae77db0_96, \6170 );
nor \U$52356 ( \52733 , \52731 , \52732 );
and \U$52357 ( \52734 , \52733 , \6175 );
not \U$52358 ( \52735 , \52733 );
and \U$52359 ( \52736 , \52735 , \6176 );
nor \U$52360 ( \52737 , \52734 , \52736 );
or \U$52361 ( \52738 , \52730 , \52737 );
not \U$52362 ( \52739 , \52737 );
not \U$52363 ( \52740 , \52730 );
or \U$52364 ( \52741 , \52739 , \52740 );
and \U$52365 ( \52742 , \6941 , RIae77ea0_98);
and \U$52366 ( \52743 , RIae789e0_122, \6939 );
nor \U$52367 ( \52744 , \52742 , \52743 );
and \U$52368 ( \52745 , \52744 , \6314 );
not \U$52369 ( \52746 , \52744 );
and \U$52370 ( \52747 , \52746 , \6945 );
nor \U$52371 ( \52748 , \52745 , \52747 );
nand \U$52372 ( \52749 , \52741 , \52748 );
nand \U$52373 ( \52750 , \52738 , \52749 );
and \U$52374 ( \52751 , \52723 , \52750 );
and \U$52375 ( \52752 , \52697 , \52722 );
or \U$52376 ( \52753 , \52751 , \52752 );
and \U$52377 ( \52754 , \12180 , RIae75560_10);
and \U$52378 ( \52755 , RIae75830_16, \12178 );
nor \U$52379 ( \52756 , \52754 , \52755 );
and \U$52380 ( \52757 , \52756 , \11827 );
not \U$52381 ( \52758 , \52756 );
and \U$52382 ( \52759 , \52758 , \12184 );
nor \U$52383 ( \52760 , \52757 , \52759 );
and \U$52384 ( \52761 , \14059 , RIae751a0_2);
and \U$52385 ( \52762 , RIae75380_6, \14057 );
nor \U$52386 ( \52763 , \52761 , \52762 );
and \U$52387 ( \52764 , \52763 , \14063 );
not \U$52388 ( \52765 , \52763 );
and \U$52389 ( \52766 , \52765 , \13502 );
nor \U$52390 ( \52767 , \52764 , \52766 );
or \U$52391 ( \52768 , \52760 , \52767 );
not \U$52392 ( \52769 , \52767 );
not \U$52393 ( \52770 , \52760 );
or \U$52394 ( \52771 , \52769 , \52770 );
and \U$52395 ( \52772 , \13059 , RIae75740_14);
and \U$52396 ( \52773 , RIae75290_4, \13057 );
nor \U$52397 ( \52774 , \52772 , \52773 );
and \U$52398 ( \52775 , \52774 , \13063 );
not \U$52399 ( \52776 , \52774 );
and \U$52400 ( \52777 , \52776 , \12718 );
nor \U$52401 ( \52778 , \52775 , \52777 );
nand \U$52402 ( \52779 , \52771 , \52778 );
nand \U$52403 ( \52780 , \52768 , \52779 );
and \U$52404 ( \52781 , \15726 , RIae76550_44);
and \U$52405 ( \52782 , RIae76730_48, RIae7aab0_192);
nor \U$52406 ( \52783 , \52781 , \52782 );
and \U$52407 ( \52784 , \52783 , \14959 );
not \U$52408 ( \52785 , \52783 );
and \U$52409 ( \52786 , \52785 , RIae7aa38_191);
nor \U$52410 ( \52787 , \52784 , \52786 );
xor \U$52411 ( \52788 , \52787 , \1142 );
and \U$52412 ( \52789 , \14964 , RIae75470_8);
and \U$52413 ( \52790 , RIae76460_42, \14962 );
nor \U$52414 ( \52791 , \52789 , \52790 );
and \U$52415 ( \52792 , \52791 , \14463 );
not \U$52416 ( \52793 , \52791 );
and \U$52417 ( \52794 , \52793 , \14462 );
nor \U$52418 ( \52795 , \52792 , \52794 );
and \U$52419 ( \52796 , \52788 , \52795 );
and \U$52420 ( \52797 , \52787 , \1142 );
or \U$52421 ( \52798 , \52796 , \52797 );
xor \U$52422 ( \52799 , \52780 , \52798 );
and \U$52423 ( \52800 , \9760 , RIae75920_18);
and \U$52424 ( \52801 , RIae75fb0_32, \9758 );
nor \U$52425 ( \52802 , \52800 , \52801 );
and \U$52426 ( \52803 , \52802 , \9764 );
not \U$52427 ( \52804 , \52802 );
and \U$52428 ( \52805 , \52804 , \9273 );
nor \U$52429 ( \52806 , \52803 , \52805 );
and \U$52430 ( \52807 , \10548 , RIae75ec0_30);
and \U$52431 ( \52808 , RIae75ce0_26, \10546 );
nor \U$52432 ( \52809 , \52807 , \52808 );
and \U$52433 ( \52810 , \52809 , \10118 );
not \U$52434 ( \52811 , \52809 );
and \U$52435 ( \52812 , \52811 , \10421 );
nor \U$52436 ( \52813 , \52810 , \52812 );
or \U$52437 ( \52814 , \52806 , \52813 );
not \U$52438 ( \52815 , \52813 );
not \U$52439 ( \52816 , \52806 );
or \U$52440 ( \52817 , \52815 , \52816 );
and \U$52441 ( \52818 , \11470 , RIae75dd0_28);
and \U$52442 ( \52819 , RIae75650_12, \11468 );
nor \U$52443 ( \52820 , \52818 , \52819 );
and \U$52444 ( \52821 , \52820 , \10936 );
not \U$52445 ( \52822 , \52820 );
and \U$52446 ( \52823 , \52822 , \11474 );
nor \U$52447 ( \52824 , \52821 , \52823 );
nand \U$52448 ( \52825 , \52817 , \52824 );
nand \U$52449 ( \52826 , \52814 , \52825 );
and \U$52450 ( \52827 , \52799 , \52826 );
and \U$52451 ( \52828 , \52780 , \52798 );
or \U$52452 ( \52829 , \52827 , \52828 );
xor \U$52453 ( \52830 , \52753 , \52829 );
and \U$52454 ( \52831 , \1939 , RIae779f0_88);
and \U$52455 ( \52832 , RIae77810_84, \1937 );
nor \U$52456 ( \52833 , \52831 , \52832 );
and \U$52457 ( \52834 , \52833 , \1734 );
not \U$52458 ( \52835 , \52833 );
and \U$52459 ( \52836 , \52835 , \1735 );
nor \U$52460 ( \52837 , \52834 , \52836 );
and \U$52461 ( \52838 , \2607 , RIae76eb0_64);
and \U$52462 ( \52839 , RIae76dc0_62, \2605 );
nor \U$52463 ( \52840 , \52838 , \52839 );
and \U$52464 ( \52841 , \52840 , \2397 );
not \U$52465 ( \52842 , \52840 );
and \U$52466 ( \52843 , \52842 , \2611 );
nor \U$52467 ( \52844 , \52841 , \52843 );
or \U$52468 ( \52845 , \52837 , \52844 );
not \U$52469 ( \52846 , \52844 );
not \U$52470 ( \52847 , \52837 );
or \U$52471 ( \52848 , \52846 , \52847 );
and \U$52472 ( \52849 , \2224 , RIae77900_86);
and \U$52473 ( \52850 , RIae76fa0_66, \2222 );
nor \U$52474 ( \52851 , \52849 , \52850 );
and \U$52475 ( \52852 , \52851 , \2061 );
not \U$52476 ( \52853 , \52851 );
and \U$52477 ( \52854 , \52853 , \2060 );
nor \U$52478 ( \52855 , \52852 , \52854 );
nand \U$52479 ( \52856 , \52848 , \52855 );
nand \U$52480 ( \52857 , \52845 , \52856 );
and \U$52481 ( \52858 , \1376 , RIae77540_78);
and \U$52482 ( \52859 , RIae776a8_81, \1374 );
nor \U$52483 ( \52860 , \52858 , \52859 );
and \U$52484 ( \52861 , \52860 , \1380 );
not \U$52485 ( \52862 , \52860 );
and \U$52486 ( \52863 , \52862 , \1261 );
nor \U$52487 ( \52864 , \52861 , \52863 );
nand \U$52488 ( \52865 , RIae77630_80, \1136 );
and \U$52489 ( \52866 , \52865 , \1012 );
not \U$52490 ( \52867 , \52865 );
and \U$52491 ( \52868 , \52867 , \1142 );
nor \U$52492 ( \52869 , \52866 , \52868 );
xor \U$52493 ( \52870 , \52864 , \52869 );
and \U$52494 ( \52871 , \1593 , RIae77450_76);
and \U$52495 ( \52872 , RIae77ae0_90, \1591 );
nor \U$52496 ( \52873 , \52871 , \52872 );
and \U$52497 ( \52874 , \52873 , \1498 );
not \U$52498 ( \52875 , \52873 );
and \U$52499 ( \52876 , \52875 , \1488 );
nor \U$52500 ( \52877 , \52874 , \52876 );
and \U$52501 ( \52878 , \52870 , \52877 );
and \U$52502 ( \52879 , \52864 , \52869 );
or \U$52503 ( \52880 , \52878 , \52879 );
xor \U$52504 ( \52881 , \52857 , \52880 );
and \U$52505 ( \52882 , \3214 , RIae77090_68);
and \U$52506 ( \52883 , RIae77270_72, \3212 );
nor \U$52507 ( \52884 , \52882 , \52883 );
not \U$52508 ( \52885 , \52884 );
not \U$52509 ( \52886 , \3218 );
and \U$52510 ( \52887 , \52885 , \52886 );
and \U$52511 ( \52888 , \52884 , \2774 );
nor \U$52512 ( \52889 , \52887 , \52888 );
and \U$52513 ( \52890 , \3730 , RIae77360_74);
and \U$52514 ( \52891 , RIae78350_108, \3728 );
nor \U$52515 ( \52892 , \52890 , \52891 );
and \U$52516 ( \52893 , \52892 , \3422 );
not \U$52517 ( \52894 , \52892 );
and \U$52518 ( \52895 , \52894 , \3732 );
nor \U$52519 ( \52896 , \52893 , \52895 );
xor \U$52520 ( \52897 , \52889 , \52896 );
and \U$52521 ( \52898 , \2783 , RIae76cd0_60);
and \U$52522 ( \52899 , RIae77108_69, \2781 );
nor \U$52523 ( \52900 , \52898 , \52899 );
not \U$52524 ( \52901 , \52900 );
not \U$52525 ( \52902 , \3089 );
and \U$52526 ( \52903 , \52901 , \52902 );
and \U$52527 ( \52904 , \52900 , \2789 );
nor \U$52528 ( \52905 , \52903 , \52904 );
and \U$52529 ( \52906 , \52897 , \52905 );
and \U$52530 ( \52907 , \52889 , \52896 );
nor \U$52531 ( \52908 , \52906 , \52907 );
and \U$52532 ( \52909 , \52881 , \52908 );
and \U$52533 ( \52910 , \52857 , \52880 );
or \U$52534 ( \52911 , \52909 , \52910 );
and \U$52535 ( \52912 , \52830 , \52911 );
and \U$52536 ( \52913 , \52753 , \52829 );
or \U$52537 ( \52914 , \52912 , \52913 );
xor \U$52538 ( \52915 , \52672 , \52914 );
xor \U$52539 ( \52916 , \51979 , \789 );
xor \U$52540 ( \52917 , \52916 , \51987 );
xor \U$52541 ( \52918 , \52259 , \52261 );
xor \U$52542 ( \52919 , \52918 , \52264 );
and \U$52543 ( \52920 , \52917 , \52919 );
xor \U$52544 ( \52921 , \51873 , \51881 );
xor \U$52545 ( \52922 , \52921 , \51890 );
xor \U$52546 ( \52923 , \52230 , \52235 );
xor \U$52547 ( \52924 , \52922 , \52923 );
xor \U$52548 ( \52925 , \52259 , \52261 );
xor \U$52549 ( \52926 , \52925 , \52264 );
and \U$52550 ( \52927 , \52924 , \52926 );
and \U$52551 ( \52928 , \52917 , \52924 );
or \U$52552 ( \52929 , \52920 , \52927 , \52928 );
and \U$52553 ( \52930 , \52915 , \52929 );
and \U$52554 ( \52931 , \52672 , \52914 );
or \U$52555 ( \52932 , \52930 , \52931 );
xor \U$52556 ( \52933 , \52343 , \52424 );
xor \U$52557 ( \52934 , \52933 , \52508 );
xor \U$52558 ( \52935 , \52240 , \52256 );
xor \U$52559 ( \52936 , \52935 , \52267 );
and \U$52560 ( \52937 , \52934 , \52936 );
xor \U$52561 ( \52938 , \52932 , \52937 );
xor \U$52562 ( \52939 , \52297 , \52312 );
xor \U$52563 ( \52940 , \52939 , \52340 );
xor \U$52564 ( \52941 , \52452 , \52479 );
xor \U$52565 ( \52942 , \52941 , \52505 );
and \U$52566 ( \52943 , \52940 , \52942 );
xor \U$52567 ( \52944 , \51926 , \51933 );
xor \U$52568 ( \52945 , \52944 , \51941 );
xor \U$52569 ( \52946 , \52246 , \52251 );
xor \U$52570 ( \52947 , \52945 , \52946 );
xor \U$52571 ( \52948 , \52452 , \52479 );
xor \U$52572 ( \52949 , \52948 , \52505 );
and \U$52573 ( \52950 , \52947 , \52949 );
and \U$52574 ( \52951 , \52940 , \52947 );
or \U$52575 ( \52952 , \52943 , \52950 , \52951 );
xor \U$52576 ( \52953 , \52534 , \52536 );
xor \U$52577 ( \52954 , \52953 , \52539 );
and \U$52578 ( \52955 , \52952 , \52954 );
xor \U$52579 ( \52956 , \52105 , \52107 );
xor \U$52580 ( \52957 , \52956 , \52110 );
xor \U$52581 ( \52958 , \52516 , \52523 );
xor \U$52582 ( \52959 , \52957 , \52958 );
xor \U$52583 ( \52960 , \52534 , \52536 );
xor \U$52584 ( \52961 , \52960 , \52539 );
and \U$52585 ( \52962 , \52959 , \52961 );
and \U$52586 ( \52963 , \52952 , \52959 );
or \U$52587 ( \52964 , \52955 , \52962 , \52963 );
and \U$52588 ( \52965 , \52938 , \52964 );
and \U$52589 ( \52966 , \52932 , \52937 );
or \U$52590 ( \52967 , \52965 , \52966 );
xor \U$52591 ( \52968 , \51866 , \52102 );
xor \U$52592 ( \52969 , \52968 , \52141 );
xor \U$52593 ( \52970 , \52967 , \52969 );
xor \U$52594 ( \52971 , \52270 , \52511 );
xor \U$52595 ( \52972 , \52971 , \52528 );
xor \U$52596 ( \52973 , \52218 , \52222 );
xor \U$52597 ( \52974 , \52973 , \52225 );
and \U$52598 ( \52975 , \52972 , \52974 );
xor \U$52599 ( \52976 , \52542 , \52543 );
xor \U$52600 ( \52977 , \52976 , \52546 );
xor \U$52601 ( \52978 , \52218 , \52222 );
xor \U$52602 ( \52979 , \52978 , \52225 );
and \U$52603 ( \52980 , \52977 , \52979 );
and \U$52604 ( \52981 , \52972 , \52977 );
or \U$52605 ( \52982 , \52975 , \52980 , \52981 );
and \U$52606 ( \52983 , \52970 , \52982 );
and \U$52607 ( \52984 , \52967 , \52969 );
or \U$52608 ( \52985 , \52983 , \52984 );
and \U$52609 ( \52986 , \52600 , \52985 );
nor \U$52610 ( \52987 , \52598 , \52986 );
not \U$52611 ( \52988 , \52987 );
and \U$52612 ( \52989 , \52584 , \52988 );
and \U$52613 ( \52990 , \52583 , \52987 );
nor \U$52614 ( \52991 , \52989 , \52990 );
not \U$52615 ( \52992 , \52552 );
not \U$52616 ( \52993 , \52570 );
or \U$52617 ( \52994 , \52992 , \52993 );
or \U$52618 ( \52995 , \52570 , \52552 );
nand \U$52619 ( \52996 , \52994 , \52995 );
not \U$52620 ( \52997 , \52996 );
not \U$52621 ( \52998 , \52216 );
and \U$52622 ( \52999 , \52997 , \52998 );
and \U$52623 ( \53000 , \52996 , \52216 );
nor \U$52624 ( \53001 , \52999 , \53000 );
not \U$52625 ( \53002 , \53001 );
not \U$52626 ( \53003 , \52597 );
not \U$52627 ( \53004 , \52985 );
not \U$52628 ( \53005 , \52594 );
and \U$52629 ( \53006 , \53004 , \53005 );
and \U$52630 ( \53007 , \52985 , \52594 );
nor \U$52631 ( \53008 , \53006 , \53007 );
not \U$52632 ( \53009 , \53008 );
or \U$52633 ( \53010 , \53003 , \53009 );
or \U$52634 ( \53011 , \53008 , \52597 );
nand \U$52635 ( \53012 , \53010 , \53011 );
nand \U$52636 ( \53013 , \53002 , \53012 );
or \U$52637 ( \53014 , \52991 , \53013 );
xnor \U$52638 ( \53015 , \53013 , \52991 );
not \U$52639 ( \53016 , \53001 );
not \U$52640 ( \53017 , \53012 );
or \U$52641 ( \53018 , \53016 , \53017 );
or \U$52642 ( \53019 , \53012 , \53001 );
nand \U$52643 ( \53020 , \53018 , \53019 );
not \U$52644 ( \53021 , \52593 );
not \U$52645 ( \53022 , \52586 );
or \U$52646 ( \53023 , \53021 , \53022 );
or \U$52647 ( \53024 , \52586 , \52593 );
nand \U$52648 ( \53025 , \53023 , \53024 );
not \U$52649 ( \53026 , \53025 );
xor \U$52650 ( \53027 , \52967 , \52969 );
xor \U$52651 ( \53028 , \53027 , \52982 );
not \U$52652 ( \53029 , \53028 );
or \U$52653 ( \53030 , \53026 , \53029 );
or \U$52654 ( \53031 , \53028 , \53025 );
xor \U$52655 ( \53032 , \52780 , \52798 );
xor \U$52656 ( \53033 , \53032 , \52826 );
xor \U$52657 ( \53034 , \52697 , \52722 );
xor \U$52658 ( \53035 , \53034 , \52750 );
xor \U$52659 ( \53036 , \53033 , \53035 );
xor \U$52660 ( \53037 , \52857 , \52880 );
xor \U$52661 ( \53038 , \53037 , \52908 );
and \U$52662 ( \53039 , \53036 , \53038 );
and \U$52663 ( \53040 , \53033 , \53035 );
or \U$52664 ( \53041 , \53039 , \53040 );
xor \U$52665 ( \53042 , \52368 , \52393 );
xor \U$52666 ( \53043 , \53042 , \52421 );
xor \U$52667 ( \53044 , \53041 , \53043 );
xor \U$52668 ( \53045 , \52452 , \52479 );
xor \U$52669 ( \53046 , \53045 , \52505 );
xor \U$52670 ( \53047 , \52940 , \52947 );
xor \U$52671 ( \53048 , \53046 , \53047 );
and \U$52672 ( \53049 , \53044 , \53048 );
and \U$52673 ( \53050 , \53041 , \53043 );
or \U$52674 ( \53051 , \53049 , \53050 );
and \U$52675 ( \53052 , \8371 , RIae78800_118);
and \U$52676 ( \53053 , RIae78710_116, \8369 );
nor \U$52677 ( \53054 , \53052 , \53053 );
and \U$52678 ( \53055 , \53054 , \8020 );
not \U$52679 ( \53056 , \53054 );
and \U$52680 ( \53057 , \53056 , \8019 );
nor \U$52681 ( \53058 , \53055 , \53057 );
and \U$52682 ( \53059 , \6941 , RIae77db0_96);
and \U$52683 ( \53060 , RIae77ea0_98, \6939 );
nor \U$52684 ( \53061 , \53059 , \53060 );
and \U$52685 ( \53062 , \53061 , \6314 );
not \U$52686 ( \53063 , \53061 );
and \U$52687 ( \53064 , \53063 , \6945 );
nor \U$52688 ( \53065 , \53062 , \53064 );
xor \U$52689 ( \53066 , \53058 , \53065 );
and \U$52690 ( \53067 , \7633 , RIae789e0_122);
and \U$52691 ( \53068 , RIae788f0_120, \7631 );
nor \U$52692 ( \53069 , \53067 , \53068 );
and \U$52693 ( \53070 , \53069 , \7206 );
not \U$52694 ( \53071 , \53069 );
and \U$52695 ( \53072 , \53071 , \7205 );
nor \U$52696 ( \53073 , \53070 , \53072 );
and \U$52697 ( \53074 , \53066 , \53073 );
and \U$52698 ( \53075 , \53058 , \53065 );
or \U$52699 ( \53076 , \53074 , \53075 );
and \U$52700 ( \53077 , \4688 , RIae77f90_100);
and \U$52701 ( \53078 , RIae78080_102, \4686 );
nor \U$52702 ( \53079 , \53077 , \53078 );
and \U$52703 ( \53080 , \53079 , \4481 );
not \U$52704 ( \53081 , \53079 );
and \U$52705 ( \53082 , \53081 , \4482 );
nor \U$52706 ( \53083 , \53080 , \53082 );
and \U$52707 ( \53084 , \3730 , RIae77270_72);
and \U$52708 ( \53085 , RIae77360_74, \3728 );
nor \U$52709 ( \53086 , \53084 , \53085 );
and \U$52710 ( \53087 , \53086 , \3732 );
not \U$52711 ( \53088 , \53086 );
and \U$52712 ( \53089 , \53088 , \3422 );
nor \U$52713 ( \53090 , \53087 , \53089 );
xor \U$52714 ( \53091 , \53083 , \53090 );
and \U$52715 ( \53092 , \4247 , RIae78350_108);
and \U$52716 ( \53093 , RIae78170_104, \4245 );
nor \U$52717 ( \53094 , \53092 , \53093 );
and \U$52718 ( \53095 , \53094 , \3989 );
not \U$52719 ( \53096 , \53094 );
and \U$52720 ( \53097 , \53096 , \4251 );
nor \U$52721 ( \53098 , \53095 , \53097 );
and \U$52722 ( \53099 , \53091 , \53098 );
and \U$52723 ( \53100 , \53083 , \53090 );
or \U$52724 ( \53101 , \53099 , \53100 );
xor \U$52725 ( \53102 , \53076 , \53101 );
and \U$52726 ( \53103 , \5896 , RIae78440_110);
and \U$52727 ( \53104 , RIae784b8_111, \5894 );
nor \U$52728 ( \53105 , \53103 , \53104 );
and \U$52729 ( \53106 , \53105 , \5590 );
not \U$52730 ( \53107 , \53105 );
and \U$52731 ( \53108 , \53107 , \5589 );
nor \U$52732 ( \53109 , \53106 , \53108 );
and \U$52733 ( \53110 , \5399 , RIae78260_106);
and \U$52734 ( \53111 , RIae78620_114, \5397 );
nor \U$52735 ( \53112 , \53110 , \53111 );
and \U$52736 ( \53113 , \53112 , \5016 );
not \U$52737 ( \53114 , \53112 );
and \U$52738 ( \53115 , \53114 , \5403 );
nor \U$52739 ( \53116 , \53113 , \53115 );
xor \U$52740 ( \53117 , \53109 , \53116 );
and \U$52741 ( \53118 , \6172 , RIae77cc0_94);
and \U$52742 ( \53119 , RIae77bd0_92, \6170 );
nor \U$52743 ( \53120 , \53118 , \53119 );
and \U$52744 ( \53121 , \53120 , \6176 );
not \U$52745 ( \53122 , \53120 );
and \U$52746 ( \53123 , \53122 , \6175 );
nor \U$52747 ( \53124 , \53121 , \53123 );
and \U$52748 ( \53125 , \53117 , \53124 );
and \U$52749 ( \53126 , \53109 , \53116 );
or \U$52750 ( \53127 , \53125 , \53126 );
and \U$52751 ( \53128 , \53102 , \53127 );
and \U$52752 ( \53129 , \53076 , \53101 );
or \U$52753 ( \53130 , \53128 , \53129 );
and \U$52754 ( \53131 , \9760 , RIae75a10_20);
and \U$52755 ( \53132 , RIae75920_18, \9758 );
nor \U$52756 ( \53133 , \53131 , \53132 );
and \U$52757 ( \53134 , \53133 , \9273 );
not \U$52758 ( \53135 , \53133 );
and \U$52759 ( \53136 , \53135 , \9272 );
nor \U$52760 ( \53137 , \53134 , \53136 );
and \U$52761 ( \53138 , \8966 , RIae75bf0_24);
and \U$52762 ( \53139 , RIae75b00_22, \8964 );
nor \U$52763 ( \53140 , \53138 , \53139 );
and \U$52764 ( \53141 , \53140 , \8799 );
not \U$52765 ( \53142 , \53140 );
and \U$52766 ( \53143 , \53142 , \8789 );
nor \U$52767 ( \53144 , \53141 , \53143 );
xor \U$52768 ( \53145 , \53137 , \53144 );
and \U$52769 ( \53146 , \10548 , RIae75fb0_32);
and \U$52770 ( \53147 , RIae75ec0_30, \10546 );
nor \U$52771 ( \53148 , \53146 , \53147 );
and \U$52772 ( \53149 , \53148 , \10421 );
not \U$52773 ( \53150 , \53148 );
and \U$52774 ( \53151 , \53150 , \10118 );
nor \U$52775 ( \53152 , \53149 , \53151 );
and \U$52776 ( \53153 , \53145 , \53152 );
and \U$52777 ( \53154 , \53137 , \53144 );
or \U$52778 ( \53155 , \53153 , \53154 );
and \U$52779 ( \53156 , \14964 , RIae75380_6);
and \U$52780 ( \53157 , RIae75470_8, \14962 );
nor \U$52781 ( \53158 , \53156 , \53157 );
and \U$52782 ( \53159 , \53158 , \14463 );
not \U$52783 ( \53160 , \53158 );
and \U$52784 ( \53161 , \53160 , \14462 );
nor \U$52785 ( \53162 , \53159 , \53161 );
and \U$52786 ( \53163 , \15726 , RIae76460_42);
and \U$52787 ( \53164 , RIae76550_44, RIae7aab0_192);
nor \U$52788 ( \53165 , \53163 , \53164 );
and \U$52789 ( \53166 , \53165 , \14959 );
not \U$52790 ( \53167 , \53165 );
and \U$52791 ( \53168 , \53167 , RIae7aa38_191);
nor \U$52792 ( \53169 , \53166 , \53168 );
xor \U$52793 ( \53170 , \53162 , \53169 );
and \U$52794 ( \53171 , \14059 , RIae75290_4);
and \U$52795 ( \53172 , RIae751a0_2, \14057 );
nor \U$52796 ( \53173 , \53171 , \53172 );
and \U$52797 ( \53174 , \53173 , \13502 );
not \U$52798 ( \53175 , \53173 );
and \U$52799 ( \53176 , \53175 , \14063 );
nor \U$52800 ( \53177 , \53174 , \53176 );
and \U$52801 ( \53178 , \53170 , \53177 );
and \U$52802 ( \53179 , \53162 , \53169 );
or \U$52803 ( \53180 , \53178 , \53179 );
xor \U$52804 ( \53181 , \53155 , \53180 );
and \U$52805 ( \53182 , \12180 , RIae75650_12);
and \U$52806 ( \53183 , RIae75560_10, \12178 );
nor \U$52807 ( \53184 , \53182 , \53183 );
and \U$52808 ( \53185 , \53184 , \12184 );
not \U$52809 ( \53186 , \53184 );
and \U$52810 ( \53187 , \53186 , \11827 );
nor \U$52811 ( \53188 , \53185 , \53187 );
and \U$52812 ( \53189 , \11470 , RIae75ce0_26);
and \U$52813 ( \53190 , RIae75dd0_28, \11468 );
nor \U$52814 ( \53191 , \53189 , \53190 );
and \U$52815 ( \53192 , \53191 , \10936 );
not \U$52816 ( \53193 , \53191 );
and \U$52817 ( \53194 , \53193 , \11474 );
nor \U$52818 ( \53195 , \53192 , \53194 );
xor \U$52819 ( \53196 , \53188 , \53195 );
and \U$52820 ( \53197 , \13059 , RIae75830_16);
and \U$52821 ( \53198 , RIae75740_14, \13057 );
nor \U$52822 ( \53199 , \53197 , \53198 );
and \U$52823 ( \53200 , \53199 , \13063 );
not \U$52824 ( \53201 , \53199 );
and \U$52825 ( \53202 , \53201 , \12718 );
nor \U$52826 ( \53203 , \53200 , \53202 );
and \U$52827 ( \53204 , \53196 , \53203 );
and \U$52828 ( \53205 , \53188 , \53195 );
or \U$52829 ( \53206 , \53204 , \53205 );
and \U$52830 ( \53207 , \53181 , \53206 );
and \U$52831 ( \53208 , \53155 , \53180 );
or \U$52832 ( \53209 , \53207 , \53208 );
xor \U$52833 ( \53210 , \53130 , \53209 );
not \U$52834 ( \53211 , \2774 );
and \U$52835 ( \53212 , \3214 , RIae77108_69);
and \U$52836 ( \53213 , RIae77090_68, \3212 );
nor \U$52837 ( \53214 , \53212 , \53213 );
not \U$52838 ( \53215 , \53214 );
or \U$52839 ( \53216 , \53211 , \53215 );
or \U$52840 ( \53217 , \53214 , \3218 );
nand \U$52841 ( \53218 , \53216 , \53217 );
and \U$52842 ( \53219 , \2607 , RIae76fa0_66);
and \U$52843 ( \53220 , RIae76eb0_64, \2605 );
nor \U$52844 ( \53221 , \53219 , \53220 );
and \U$52845 ( \53222 , \53221 , \2611 );
not \U$52846 ( \53223 , \53221 );
and \U$52847 ( \53224 , \53223 , \2396 );
nor \U$52848 ( \53225 , \53222 , \53224 );
xor \U$52849 ( \53226 , \53218 , \53225 );
not \U$52850 ( \53227 , \3089 );
and \U$52851 ( \53228 , \2783 , RIae76dc0_62);
and \U$52852 ( \53229 , RIae76cd0_60, \2781 );
nor \U$52853 ( \53230 , \53228 , \53229 );
not \U$52854 ( \53231 , \53230 );
or \U$52855 ( \53232 , \53227 , \53231 );
or \U$52856 ( \53233 , \53230 , \3089 );
nand \U$52857 ( \53234 , \53232 , \53233 );
and \U$52858 ( \53235 , \53226 , \53234 );
and \U$52859 ( \53236 , \53218 , \53225 );
or \U$52860 ( \53237 , \53235 , \53236 );
and \U$52861 ( \53238 , \1593 , RIae776a8_81);
and \U$52862 ( \53239 , RIae77450_76, \1591 );
nor \U$52863 ( \53240 , \53238 , \53239 );
and \U$52864 ( \53241 , \53240 , \1498 );
not \U$52865 ( \53242 , \53240 );
and \U$52866 ( \53243 , \53242 , \1488 );
nor \U$52867 ( \53244 , \53241 , \53243 );
and \U$52868 ( \53245 , \1939 , RIae77ae0_90);
and \U$52869 ( \53246 , RIae779f0_88, \1937 );
nor \U$52870 ( \53247 , \53245 , \53246 );
and \U$52871 ( \53248 , \53247 , \1735 );
not \U$52872 ( \53249 , \53247 );
and \U$52873 ( \53250 , \53249 , \1734 );
nor \U$52874 ( \53251 , \53248 , \53250 );
xor \U$52875 ( \53252 , \53244 , \53251 );
and \U$52876 ( \53253 , \2224 , RIae77810_84);
and \U$52877 ( \53254 , RIae77900_86, \2222 );
nor \U$52878 ( \53255 , \53253 , \53254 );
and \U$52879 ( \53256 , \53255 , \2061 );
not \U$52880 ( \53257 , \53255 );
and \U$52881 ( \53258 , \53257 , \2060 );
nor \U$52882 ( \53259 , \53256 , \53258 );
and \U$52883 ( \53260 , \53252 , \53259 );
and \U$52884 ( \53261 , \53244 , \53251 );
or \U$52885 ( \53262 , \53260 , \53261 );
xor \U$52886 ( \53263 , \53237 , \53262 );
xor \U$52887 ( \53264 , \52864 , \52869 );
xor \U$52888 ( \53265 , \53264 , \52877 );
and \U$52889 ( \53266 , \53263 , \53265 );
and \U$52890 ( \53267 , \53237 , \53262 );
or \U$52891 ( \53268 , \53266 , \53267 );
and \U$52892 ( \53269 , \53210 , \53268 );
and \U$52893 ( \53270 , \53130 , \53209 );
nor \U$52894 ( \53271 , \53269 , \53270 );
xor \U$52895 ( \53272 , \52679 , \52686 );
xor \U$52896 ( \53273 , \53272 , \52694 );
not \U$52897 ( \53274 , \53273 );
not \U$52898 ( \53275 , \52813 );
not \U$52899 ( \53276 , \52824 );
or \U$52900 ( \53277 , \53275 , \53276 );
or \U$52901 ( \53278 , \52813 , \52824 );
nand \U$52902 ( \53279 , \53277 , \53278 );
not \U$52903 ( \53280 , \53279 );
not \U$52904 ( \53281 , \52806 );
and \U$52905 ( \53282 , \53280 , \53281 );
and \U$52906 ( \53283 , \53279 , \52806 );
nor \U$52907 ( \53284 , \53282 , \53283 );
not \U$52908 ( \53285 , \53284 );
and \U$52909 ( \53286 , \53274 , \53285 );
and \U$52910 ( \53287 , \53284 , \53273 );
not \U$52911 ( \53288 , \52737 );
not \U$52912 ( \53289 , \52748 );
or \U$52913 ( \53290 , \53288 , \53289 );
or \U$52914 ( \53291 , \52737 , \52748 );
nand \U$52915 ( \53292 , \53290 , \53291 );
not \U$52916 ( \53293 , \53292 );
not \U$52917 ( \53294 , \52730 );
and \U$52918 ( \53295 , \53293 , \53294 );
and \U$52919 ( \53296 , \53292 , \52730 );
nor \U$52920 ( \53297 , \53295 , \53296 );
nor \U$52921 ( \53298 , \53287 , \53297 );
nor \U$52922 ( \53299 , \53286 , \53298 );
not \U$52923 ( \53300 , \52767 );
not \U$52924 ( \53301 , \52778 );
or \U$52925 ( \53302 , \53300 , \53301 );
or \U$52926 ( \53303 , \52767 , \52778 );
nand \U$52927 ( \53304 , \53302 , \53303 );
not \U$52928 ( \53305 , \53304 );
not \U$52929 ( \53306 , \52760 );
and \U$52930 ( \53307 , \53305 , \53306 );
and \U$52931 ( \53308 , \53304 , \52760 );
nor \U$52932 ( \53309 , \53307 , \53308 );
not \U$52933 ( \53310 , \53309 );
xor \U$52934 ( \53311 , \52787 , \1142 );
xor \U$52935 ( \53312 , \53311 , \52795 );
nand \U$52936 ( \53313 , \53310 , \53312 );
xor \U$52937 ( \53314 , \53299 , \53313 );
not \U$52938 ( \53315 , \52844 );
not \U$52939 ( \53316 , \52855 );
or \U$52940 ( \53317 , \53315 , \53316 );
or \U$52941 ( \53318 , \52844 , \52855 );
nand \U$52942 ( \53319 , \53317 , \53318 );
not \U$52943 ( \53320 , \53319 );
not \U$52944 ( \53321 , \52837 );
and \U$52945 ( \53322 , \53320 , \53321 );
and \U$52946 ( \53323 , \53319 , \52837 );
nor \U$52947 ( \53324 , \53322 , \53323 );
not \U$52948 ( \53325 , \53324 );
xor \U$52949 ( \53326 , \52704 , \52711 );
xor \U$52950 ( \53327 , \53326 , \52719 );
not \U$52951 ( \53328 , \53327 );
and \U$52952 ( \53329 , \53325 , \53328 );
and \U$52953 ( \53330 , \53327 , \53324 );
xor \U$52954 ( \53331 , \52889 , \52896 );
xor \U$52955 ( \53332 , \53331 , \52905 );
nor \U$52956 ( \53333 , \53330 , \53332 );
nor \U$52957 ( \53334 , \53329 , \53333 );
and \U$52958 ( \53335 , \53314 , \53334 );
and \U$52959 ( \53336 , \53299 , \53313 );
or \U$52960 ( \53337 , \53335 , \53336 );
xor \U$52961 ( \53338 , \53271 , \53337 );
not \U$52962 ( \53339 , \52638 );
not \U$52963 ( \53340 , \52646 );
and \U$52964 ( \53341 , \53339 , \53340 );
and \U$52965 ( \53342 , \52638 , \52646 );
nor \U$52966 ( \53343 , \53341 , \53342 );
not \U$52967 ( \53344 , \53343 );
not \U$52968 ( \53345 , \52639 );
and \U$52969 ( \53346 , \53344 , \53345 );
and \U$52970 ( \53347 , \53343 , \52639 );
nor \U$52971 ( \53348 , \53346 , \53347 );
not \U$52972 ( \53349 , \53348 );
not \U$52973 ( \53350 , \52620 );
not \U$52974 ( \53351 , \52626 );
or \U$52975 ( \53352 , \53350 , \53351 );
or \U$52976 ( \53353 , \52620 , \52626 );
nand \U$52977 ( \53354 , \53352 , \53353 );
not \U$52978 ( \53355 , \53354 );
not \U$52979 ( \53356 , \52610 );
and \U$52980 ( \53357 , \53355 , \53356 );
and \U$52981 ( \53358 , \53354 , \52610 );
nor \U$52982 ( \53359 , \53357 , \53358 );
not \U$52983 ( \53360 , \53359 );
and \U$52984 ( \53361 , \53349 , \53360 );
and \U$52985 ( \53362 , \53359 , \53348 );
not \U$52986 ( \53363 , \52659 );
not \U$52987 ( \53364 , \52667 );
or \U$52988 ( \53365 , \53363 , \53364 );
or \U$52989 ( \53366 , \52667 , \52659 );
nand \U$52990 ( \53367 , \53365 , \53366 );
not \U$52991 ( \53368 , \53367 );
not \U$52992 ( \53369 , \52661 );
and \U$52993 ( \53370 , \53368 , \53369 );
and \U$52994 ( \53371 , \53367 , \52661 );
nor \U$52995 ( \53372 , \53370 , \53371 );
nor \U$52996 ( \53373 , \53362 , \53372 );
nor \U$52997 ( \53374 , \53361 , \53373 );
and \U$52998 ( \53375 , \53338 , \53374 );
and \U$52999 ( \53376 , \53271 , \53337 );
nor \U$53000 ( \53377 , \53375 , \53376 );
xor \U$53001 ( \53378 , \53051 , \53377 );
xor \U$53002 ( \53379 , \52753 , \52829 );
xor \U$53003 ( \53380 , \53379 , \52911 );
xor \U$53004 ( \53381 , \52628 , \52648 );
xor \U$53005 ( \53382 , \53381 , \52669 );
and \U$53006 ( \53383 , \53380 , \53382 );
xor \U$53007 ( \53384 , \52259 , \52261 );
xor \U$53008 ( \53385 , \53384 , \52264 );
xor \U$53009 ( \53386 , \52917 , \52924 );
xor \U$53010 ( \53387 , \53385 , \53386 );
xor \U$53011 ( \53388 , \52628 , \52648 );
xor \U$53012 ( \53389 , \53388 , \52669 );
and \U$53013 ( \53390 , \53387 , \53389 );
and \U$53014 ( \53391 , \53380 , \53387 );
or \U$53015 ( \53392 , \53383 , \53390 , \53391 );
and \U$53016 ( \53393 , \53378 , \53392 );
and \U$53017 ( \53394 , \53051 , \53377 );
or \U$53018 ( \53395 , \53393 , \53394 );
xor \U$53019 ( \53396 , \52934 , \52936 );
xor \U$53020 ( \53397 , \52672 , \52914 );
xor \U$53021 ( \53398 , \53397 , \52929 );
and \U$53022 ( \53399 , \53396 , \53398 );
xor \U$53023 ( \53400 , \52534 , \52536 );
xor \U$53024 ( \53401 , \53400 , \52539 );
xor \U$53025 ( \53402 , \52952 , \52959 );
xor \U$53026 ( \53403 , \53401 , \53402 );
xor \U$53027 ( \53404 , \52672 , \52914 );
xor \U$53028 ( \53405 , \53404 , \52929 );
and \U$53029 ( \53406 , \53403 , \53405 );
and \U$53030 ( \53407 , \53396 , \53403 );
or \U$53031 ( \53408 , \53399 , \53406 , \53407 );
xor \U$53032 ( \53409 , \53395 , \53408 );
xor \U$53033 ( \53410 , \52218 , \52222 );
xor \U$53034 ( \53411 , \53410 , \52225 );
xor \U$53035 ( \53412 , \52972 , \52977 );
xor \U$53036 ( \53413 , \53411 , \53412 );
and \U$53037 ( \53414 , \53409 , \53413 );
and \U$53038 ( \53415 , \53395 , \53408 );
or \U$53039 ( \53416 , \53414 , \53415 );
nand \U$53040 ( \53417 , \53031 , \53416 );
nand \U$53041 ( \53418 , \53030 , \53417 );
and \U$53042 ( \53419 , \53020 , \53418 );
xor \U$53043 ( \53420 , \53418 , \53020 );
and \U$53044 ( \53421 , \6172 , RIae78350_108);
and \U$53045 ( \53422 , RIae78170_104, \6170 );
nor \U$53046 ( \53423 , \53421 , \53422 );
and \U$53047 ( \53424 , \53423 , \6176 );
not \U$53048 ( \53425 , \53423 );
and \U$53049 ( \53426 , \53425 , \6175 );
nor \U$53050 ( \53427 , \53424 , \53426 );
and \U$53051 ( \53428 , \5399 , RIae77108_69);
and \U$53052 ( \53429 , RIae77090_68, \5397 );
nor \U$53053 ( \53430 , \53428 , \53429 );
and \U$53054 ( \53431 , \53430 , \5016 );
not \U$53055 ( \53432 , \53430 );
and \U$53056 ( \53433 , \53432 , \5403 );
nor \U$53057 ( \53434 , \53431 , \53433 );
xor \U$53058 ( \53435 , \53427 , \53434 );
and \U$53059 ( \53436 , \5896 , RIae77270_72);
and \U$53060 ( \53437 , RIae77360_74, \5894 );
nor \U$53061 ( \53438 , \53436 , \53437 );
and \U$53062 ( \53439 , \53438 , \5590 );
not \U$53063 ( \53440 , \53438 );
and \U$53064 ( \53441 , \53440 , \5589 );
nor \U$53065 ( \53442 , \53439 , \53441 );
and \U$53066 ( \53443 , \53435 , \53442 );
and \U$53067 ( \53444 , \53427 , \53434 );
or \U$53068 ( \53445 , \53443 , \53444 );
and \U$53069 ( \53446 , \3730 , RIae77810_84);
and \U$53070 ( \53447 , RIae77900_86, \3728 );
nor \U$53071 ( \53448 , \53446 , \53447 );
and \U$53072 ( \53449 , \53448 , \3732 );
not \U$53073 ( \53450 , \53448 );
and \U$53074 ( \53451 , \53450 , \3422 );
nor \U$53075 ( \53452 , \53449 , \53451 );
and \U$53076 ( \53453 , \4247 , RIae76fa0_66);
and \U$53077 ( \53454 , RIae76eb0_64, \4245 );
nor \U$53078 ( \53455 , \53453 , \53454 );
and \U$53079 ( \53456 , \53455 , \3989 );
not \U$53080 ( \53457 , \53455 );
and \U$53081 ( \53458 , \53457 , \4251 );
nor \U$53082 ( \53459 , \53456 , \53458 );
xor \U$53083 ( \53460 , \53452 , \53459 );
and \U$53084 ( \53461 , \4688 , RIae76dc0_62);
and \U$53085 ( \53462 , RIae76cd0_60, \4686 );
nor \U$53086 ( \53463 , \53461 , \53462 );
and \U$53087 ( \53464 , \53463 , \4481 );
not \U$53088 ( \53465 , \53463 );
and \U$53089 ( \53466 , \53465 , \4482 );
nor \U$53090 ( \53467 , \53464 , \53466 );
and \U$53091 ( \53468 , \53460 , \53467 );
and \U$53092 ( \53469 , \53452 , \53459 );
or \U$53093 ( \53470 , \53468 , \53469 );
xor \U$53094 ( \53471 , \53445 , \53470 );
and \U$53095 ( \53472 , \6941 , RIae77f90_100);
and \U$53096 ( \53473 , RIae78080_102, \6939 );
nor \U$53097 ( \53474 , \53472 , \53473 );
and \U$53098 ( \53475 , \53474 , \6314 );
not \U$53099 ( \53476 , \53474 );
and \U$53100 ( \53477 , \53476 , \6945 );
nor \U$53101 ( \53478 , \53475 , \53477 );
and \U$53102 ( \53479 , \7633 , RIae78260_106);
and \U$53103 ( \53480 , RIae78620_114, \7631 );
nor \U$53104 ( \53481 , \53479 , \53480 );
and \U$53105 ( \53482 , \53481 , \7206 );
not \U$53106 ( \53483 , \53481 );
and \U$53107 ( \53484 , \53483 , \7205 );
nor \U$53108 ( \53485 , \53482 , \53484 );
xor \U$53109 ( \53486 , \53478 , \53485 );
and \U$53110 ( \53487 , \8371 , RIae78440_110);
and \U$53111 ( \53488 , RIae784b8_111, \8369 );
nor \U$53112 ( \53489 , \53487 , \53488 );
and \U$53113 ( \53490 , \53489 , \8020 );
not \U$53114 ( \53491 , \53489 );
and \U$53115 ( \53492 , \53491 , \8019 );
nor \U$53116 ( \53493 , \53490 , \53492 );
and \U$53117 ( \53494 , \53486 , \53493 );
and \U$53118 ( \53495 , \53478 , \53485 );
or \U$53119 ( \53496 , \53494 , \53495 );
and \U$53120 ( \53497 , \53471 , \53496 );
and \U$53121 ( \53498 , \53445 , \53470 );
or \U$53122 ( \53499 , \53497 , \53498 );
and \U$53123 ( \53500 , \10548 , RIae789e0_122);
and \U$53124 ( \53501 , RIae788f0_120, \10546 );
nor \U$53125 ( \53502 , \53500 , \53501 );
and \U$53126 ( \53503 , \53502 , \10421 );
not \U$53127 ( \53504 , \53502 );
and \U$53128 ( \53505 , \53504 , \10118 );
nor \U$53129 ( \53506 , \53503 , \53505 );
and \U$53130 ( \53507 , \8966 , RIae77cc0_94);
and \U$53131 ( \53508 , RIae77bd0_92, \8964 );
nor \U$53132 ( \53509 , \53507 , \53508 );
and \U$53133 ( \53510 , \53509 , \8799 );
not \U$53134 ( \53511 , \53509 );
and \U$53135 ( \53512 , \53511 , \8789 );
nor \U$53136 ( \53513 , \53510 , \53512 );
xor \U$53137 ( \53514 , \53506 , \53513 );
and \U$53138 ( \53515 , \9760 , RIae77db0_96);
and \U$53139 ( \53516 , RIae77ea0_98, \9758 );
nor \U$53140 ( \53517 , \53515 , \53516 );
and \U$53141 ( \53518 , \53517 , \9273 );
not \U$53142 ( \53519 , \53517 );
and \U$53143 ( \53520 , \53519 , \9764 );
nor \U$53144 ( \53521 , \53518 , \53520 );
and \U$53145 ( \53522 , \53514 , \53521 );
and \U$53146 ( \53523 , \53506 , \53513 );
or \U$53147 ( \53524 , \53522 , \53523 );
and \U$53148 ( \53525 , \14964 , RIae75ce0_26);
and \U$53149 ( \53526 , RIae75dd0_28, \14962 );
nor \U$53150 ( \53527 , \53525 , \53526 );
and \U$53151 ( \53528 , \53527 , \14463 );
not \U$53152 ( \53529 , \53527 );
and \U$53153 ( \53530 , \53529 , \14462 );
nor \U$53154 ( \53531 , \53528 , \53530 );
and \U$53155 ( \53532 , \15726 , RIae75650_12);
and \U$53156 ( \53533 , RIae75560_10, RIae7aab0_192);
nor \U$53157 ( \53534 , \53532 , \53533 );
and \U$53158 ( \53535 , \53534 , \14959 );
not \U$53159 ( \53536 , \53534 );
and \U$53160 ( \53537 , \53536 , RIae7aa38_191);
nor \U$53161 ( \53538 , \53535 , \53537 );
xor \U$53162 ( \53539 , \53531 , \53538 );
and \U$53163 ( \53540 , \14059 , RIae75fb0_32);
and \U$53164 ( \53541 , RIae75ec0_30, \14057 );
nor \U$53165 ( \53542 , \53540 , \53541 );
and \U$53166 ( \53543 , \53542 , \13502 );
not \U$53167 ( \53544 , \53542 );
and \U$53168 ( \53545 , \53544 , \14063 );
nor \U$53169 ( \53546 , \53543 , \53545 );
and \U$53170 ( \53547 , \53539 , \53546 );
and \U$53171 ( \53548 , \53531 , \53538 );
or \U$53172 ( \53549 , \53547 , \53548 );
xor \U$53173 ( \53550 , \53524 , \53549 );
and \U$53174 ( \53551 , \11470 , RIae78800_118);
and \U$53175 ( \53552 , RIae78710_116, \11468 );
nor \U$53176 ( \53553 , \53551 , \53552 );
and \U$53177 ( \53554 , \53553 , \10936 );
not \U$53178 ( \53555 , \53553 );
and \U$53179 ( \53556 , \53555 , \11474 );
nor \U$53180 ( \53557 , \53554 , \53556 );
and \U$53181 ( \53558 , \12180 , RIae75bf0_24);
and \U$53182 ( \53559 , RIae75b00_22, \12178 );
nor \U$53183 ( \53560 , \53558 , \53559 );
and \U$53184 ( \53561 , \53560 , \12184 );
not \U$53185 ( \53562 , \53560 );
and \U$53186 ( \53563 , \53562 , \11827 );
nor \U$53187 ( \53564 , \53561 , \53563 );
xor \U$53188 ( \53565 , \53557 , \53564 );
and \U$53189 ( \53566 , \13059 , RIae75a10_20);
and \U$53190 ( \53567 , RIae75920_18, \13057 );
nor \U$53191 ( \53568 , \53566 , \53567 );
and \U$53192 ( \53569 , \53568 , \13063 );
not \U$53193 ( \53570 , \53568 );
and \U$53194 ( \53571 , \53570 , \12718 );
nor \U$53195 ( \53572 , \53569 , \53571 );
and \U$53196 ( \53573 , \53565 , \53572 );
and \U$53197 ( \53574 , \53557 , \53564 );
or \U$53198 ( \53575 , \53573 , \53574 );
and \U$53199 ( \53576 , \53550 , \53575 );
and \U$53200 ( \53577 , \53524 , \53549 );
or \U$53201 ( \53578 , \53576 , \53577 );
xor \U$53202 ( \53579 , \53499 , \53578 );
not \U$53203 ( \53580 , \2774 );
and \U$53204 ( \53581 , \3214 , RIae77ae0_90);
and \U$53205 ( \53582 , RIae779f0_88, \3212 );
nor \U$53206 ( \53583 , \53581 , \53582 );
not \U$53207 ( \53584 , \53583 );
or \U$53208 ( \53585 , \53580 , \53584 );
or \U$53209 ( \53586 , \53583 , \3218 );
nand \U$53210 ( \53587 , \53585 , \53586 );
and \U$53211 ( \53588 , \2607 , RIae77630_80);
and \U$53212 ( \53589 , RIae77540_78, \2605 );
nor \U$53213 ( \53590 , \53588 , \53589 );
and \U$53214 ( \53591 , \53590 , \2611 );
not \U$53215 ( \53592 , \53590 );
and \U$53216 ( \53593 , \53592 , \2396 );
nor \U$53217 ( \53594 , \53591 , \53593 );
xor \U$53218 ( \53595 , \53587 , \53594 );
not \U$53219 ( \53596 , \3089 );
and \U$53220 ( \53597 , \2783 , RIae776a8_81);
and \U$53221 ( \53598 , RIae77450_76, \2781 );
nor \U$53222 ( \53599 , \53597 , \53598 );
not \U$53223 ( \53600 , \53599 );
or \U$53224 ( \53601 , \53596 , \53600 );
or \U$53225 ( \53602 , \53599 , \3089 );
nand \U$53226 ( \53603 , \53601 , \53602 );
and \U$53227 ( \53604 , \53595 , \53603 );
and \U$53228 ( \53605 , \53587 , \53594 );
or \U$53229 ( \53606 , \53604 , \53605 );
nand \U$53230 ( \53607 , RIae77630_80, \2222 );
and \U$53231 ( \53608 , \53607 , \2061 );
not \U$53232 ( \53609 , \53607 );
and \U$53233 ( \53610 , \53609 , \2060 );
nor \U$53234 ( \53611 , \53608 , \53610 );
and \U$53235 ( \53612 , \2607 , RIae77540_78);
and \U$53236 ( \53613 , RIae776a8_81, \2605 );
nor \U$53237 ( \53614 , \53612 , \53613 );
and \U$53238 ( \53615 , \53614 , \2611 );
not \U$53239 ( \53616 , \53614 );
and \U$53240 ( \53617 , \53616 , \2397 );
nor \U$53241 ( \53618 , \53615 , \53617 );
xor \U$53242 ( \53619 , \53611 , \53618 );
xor \U$53243 ( \53620 , \53606 , \53619 );
not \U$53244 ( \53621 , \3089 );
and \U$53245 ( \53622 , \2783 , RIae77450_76);
and \U$53246 ( \53623 , RIae77ae0_90, \2781 );
nor \U$53247 ( \53624 , \53622 , \53623 );
not \U$53248 ( \53625 , \53624 );
or \U$53249 ( \53626 , \53621 , \53625 );
or \U$53250 ( \53627 , \53624 , \2789 );
nand \U$53251 ( \53628 , \53626 , \53627 );
not \U$53252 ( \53629 , \2774 );
and \U$53253 ( \53630 , \3214 , RIae779f0_88);
and \U$53254 ( \53631 , RIae77810_84, \3212 );
nor \U$53255 ( \53632 , \53630 , \53631 );
not \U$53256 ( \53633 , \53632 );
or \U$53257 ( \53634 , \53629 , \53633 );
or \U$53258 ( \53635 , \53632 , \2774 );
nand \U$53259 ( \53636 , \53634 , \53635 );
xor \U$53260 ( \53637 , \53628 , \53636 );
and \U$53261 ( \53638 , \3730 , RIae77900_86);
and \U$53262 ( \53639 , RIae76fa0_66, \3728 );
nor \U$53263 ( \53640 , \53638 , \53639 );
and \U$53264 ( \53641 , \53640 , \3732 );
not \U$53265 ( \53642 , \53640 );
and \U$53266 ( \53643 , \53642 , \3422 );
nor \U$53267 ( \53644 , \53641 , \53643 );
xor \U$53268 ( \53645 , \53637 , \53644 );
and \U$53269 ( \53646 , \53620 , \53645 );
and \U$53270 ( \53647 , \53606 , \53619 );
or \U$53271 ( \53648 , \53646 , \53647 );
and \U$53272 ( \53649 , \53579 , \53648 );
and \U$53273 ( \53650 , \53499 , \53578 );
nor \U$53274 ( \53651 , \53649 , \53650 );
and \U$53275 ( \53652 , \9760 , RIae77ea0_98);
and \U$53276 ( \53653 , RIae789e0_122, \9758 );
nor \U$53277 ( \53654 , \53652 , \53653 );
and \U$53278 ( \53655 , \53654 , \9273 );
not \U$53279 ( \53656 , \53654 );
and \U$53280 ( \53657 , \53656 , \9764 );
nor \U$53281 ( \53658 , \53655 , \53657 );
and \U$53282 ( \53659 , \10548 , RIae788f0_120);
and \U$53283 ( \53660 , RIae78800_118, \10546 );
nor \U$53284 ( \53661 , \53659 , \53660 );
and \U$53285 ( \53662 , \53661 , \10421 );
not \U$53286 ( \53663 , \53661 );
and \U$53287 ( \53664 , \53663 , \10118 );
nor \U$53288 ( \53665 , \53662 , \53664 );
xor \U$53289 ( \53666 , \53658 , \53665 );
and \U$53290 ( \53667 , \11470 , RIae78710_116);
and \U$53291 ( \53668 , RIae75bf0_24, \11468 );
nor \U$53292 ( \53669 , \53667 , \53668 );
and \U$53293 ( \53670 , \53669 , \10936 );
not \U$53294 ( \53671 , \53669 );
and \U$53295 ( \53672 , \53671 , \11474 );
nor \U$53296 ( \53673 , \53670 , \53672 );
xor \U$53297 ( \53674 , \53666 , \53673 );
and \U$53298 ( \53675 , \15726 , RIae75560_10);
and \U$53299 ( \53676 , RIae75830_16, RIae7aab0_192);
nor \U$53300 ( \53677 , \53675 , \53676 );
and \U$53301 ( \53678 , \53677 , \14959 );
not \U$53302 ( \53679 , \53677 );
and \U$53303 ( \53680 , \53679 , RIae7aa38_191);
nor \U$53304 ( \53681 , \53678 , \53680 );
xor \U$53305 ( \53682 , \53681 , \2060 );
and \U$53306 ( \53683 , \14964 , RIae75dd0_28);
and \U$53307 ( \53684 , RIae75650_12, \14962 );
nor \U$53308 ( \53685 , \53683 , \53684 );
and \U$53309 ( \53686 , \53685 , \14463 );
not \U$53310 ( \53687 , \53685 );
and \U$53311 ( \53688 , \53687 , \14462 );
nor \U$53312 ( \53689 , \53686 , \53688 );
xor \U$53313 ( \53690 , \53682 , \53689 );
and \U$53314 ( \53691 , \53674 , \53690 );
and \U$53315 ( \53692 , \12180 , RIae75b00_22);
and \U$53316 ( \53693 , RIae75a10_20, \12178 );
nor \U$53317 ( \53694 , \53692 , \53693 );
and \U$53318 ( \53695 , \53694 , \12184 );
not \U$53319 ( \53696 , \53694 );
and \U$53320 ( \53697 , \53696 , \11827 );
nor \U$53321 ( \53698 , \53695 , \53697 );
and \U$53322 ( \53699 , \13059 , RIae75920_18);
and \U$53323 ( \53700 , RIae75fb0_32, \13057 );
nor \U$53324 ( \53701 , \53699 , \53700 );
and \U$53325 ( \53702 , \53701 , \13063 );
not \U$53326 ( \53703 , \53701 );
and \U$53327 ( \53704 , \53703 , \12718 );
nor \U$53328 ( \53705 , \53702 , \53704 );
xor \U$53329 ( \53706 , \53698 , \53705 );
and \U$53330 ( \53707 , \14059 , RIae75ec0_30);
and \U$53331 ( \53708 , RIae75ce0_26, \14057 );
nor \U$53332 ( \53709 , \53707 , \53708 );
and \U$53333 ( \53710 , \53709 , \13502 );
not \U$53334 ( \53711 , \53709 );
and \U$53335 ( \53712 , \53711 , \14063 );
nor \U$53336 ( \53713 , \53710 , \53712 );
xor \U$53337 ( \53714 , \53706 , \53713 );
xor \U$53338 ( \53715 , \53681 , \2060 );
xor \U$53339 ( \53716 , \53715 , \53689 );
and \U$53340 ( \53717 , \53714 , \53716 );
and \U$53341 ( \53718 , \53674 , \53714 );
or \U$53342 ( \53719 , \53691 , \53717 , \53718 );
not \U$53343 ( \53720 , \53719 );
not \U$53344 ( \53721 , \53720 );
and \U$53345 ( \53722 , \15726 , RIae75830_16);
and \U$53346 ( \53723 , RIae75740_14, RIae7aab0_192);
nor \U$53347 ( \53724 , \53722 , \53723 );
and \U$53348 ( \53725 , \53724 , RIae7aa38_191);
not \U$53349 ( \53726 , \53724 );
and \U$53350 ( \53727 , \53726 , \14959 );
nor \U$53351 ( \53728 , \53725 , \53727 );
not \U$53352 ( \53729 , \53728 );
and \U$53353 ( \53730 , \14964 , RIae75650_12);
and \U$53354 ( \53731 , RIae75560_10, \14962 );
nor \U$53355 ( \53732 , \53730 , \53731 );
and \U$53356 ( \53733 , \53732 , \14463 );
not \U$53357 ( \53734 , \53732 );
and \U$53358 ( \53735 , \53734 , \14462 );
nor \U$53359 ( \53736 , \53733 , \53735 );
not \U$53360 ( \53737 , \53736 );
or \U$53361 ( \53738 , \53729 , \53737 );
or \U$53362 ( \53739 , \53736 , \53728 );
nand \U$53363 ( \53740 , \53738 , \53739 );
not \U$53364 ( \53741 , \53740 );
and \U$53365 ( \53742 , \14059 , RIae75ce0_26);
and \U$53366 ( \53743 , RIae75dd0_28, \14057 );
nor \U$53367 ( \53744 , \53742 , \53743 );
and \U$53368 ( \53745 , \53744 , \14063 );
not \U$53369 ( \53746 , \53744 );
and \U$53370 ( \53747 , \53746 , \13502 );
nor \U$53371 ( \53748 , \53745 , \53747 );
not \U$53372 ( \53749 , \53748 );
and \U$53373 ( \53750 , \53741 , \53749 );
and \U$53374 ( \53751 , \53740 , \53748 );
nor \U$53375 ( \53752 , \53750 , \53751 );
not \U$53376 ( \53753 , \53752 );
and \U$53377 ( \53754 , \53721 , \53753 );
and \U$53378 ( \53755 , \53720 , \53752 );
and \U$53379 ( \53756 , \6172 , RIae78170_104);
and \U$53380 ( \53757 , RIae77f90_100, \6170 );
nor \U$53381 ( \53758 , \53756 , \53757 );
and \U$53382 ( \53759 , \53758 , \6175 );
not \U$53383 ( \53760 , \53758 );
and \U$53384 ( \53761 , \53760 , \6176 );
nor \U$53385 ( \53762 , \53759 , \53761 );
not \U$53386 ( \53763 , \53762 );
and \U$53387 ( \53764 , \6941 , RIae78080_102);
and \U$53388 ( \53765 , RIae78260_106, \6939 );
nor \U$53389 ( \53766 , \53764 , \53765 );
and \U$53390 ( \53767 , \53766 , \6314 );
not \U$53391 ( \53768 , \53766 );
and \U$53392 ( \53769 , \53768 , \6945 );
nor \U$53393 ( \53770 , \53767 , \53769 );
not \U$53394 ( \53771 , \53770 );
or \U$53395 ( \53772 , \53763 , \53771 );
or \U$53396 ( \53773 , \53762 , \53770 );
nand \U$53397 ( \53774 , \53772 , \53773 );
not \U$53398 ( \53775 , \53774 );
and \U$53399 ( \53776 , \5896 , RIae77360_74);
and \U$53400 ( \53777 , RIae78350_108, \5894 );
nor \U$53401 ( \53778 , \53776 , \53777 );
and \U$53402 ( \53779 , \53778 , \5589 );
not \U$53403 ( \53780 , \53778 );
and \U$53404 ( \53781 , \53780 , \5590 );
nor \U$53405 ( \53782 , \53779 , \53781 );
not \U$53406 ( \53783 , \53782 );
and \U$53407 ( \53784 , \53775 , \53783 );
and \U$53408 ( \53785 , \53774 , \53782 );
nor \U$53409 ( \53786 , \53784 , \53785 );
not \U$53410 ( \53787 , \53786 );
and \U$53411 ( \53788 , \8966 , RIae77bd0_92);
and \U$53412 ( \53789 , RIae77db0_96, \8964 );
nor \U$53413 ( \53790 , \53788 , \53789 );
and \U$53414 ( \53791 , \53790 , \8789 );
not \U$53415 ( \53792 , \53790 );
and \U$53416 ( \53793 , \53792 , \8799 );
nor \U$53417 ( \53794 , \53791 , \53793 );
not \U$53418 ( \53795 , \53794 );
and \U$53419 ( \53796 , \8371 , RIae784b8_111);
and \U$53420 ( \53797 , RIae77cc0_94, \8369 );
nor \U$53421 ( \53798 , \53796 , \53797 );
and \U$53422 ( \53799 , \53798 , \8020 );
not \U$53423 ( \53800 , \53798 );
and \U$53424 ( \53801 , \53800 , \8019 );
nor \U$53425 ( \53802 , \53799 , \53801 );
not \U$53426 ( \53803 , \53802 );
or \U$53427 ( \53804 , \53795 , \53803 );
or \U$53428 ( \53805 , \53794 , \53802 );
nand \U$53429 ( \53806 , \53804 , \53805 );
not \U$53430 ( \53807 , \53806 );
and \U$53431 ( \53808 , \7633 , RIae78620_114);
and \U$53432 ( \53809 , RIae78440_110, \7631 );
nor \U$53433 ( \53810 , \53808 , \53809 );
and \U$53434 ( \53811 , \53810 , \7205 );
not \U$53435 ( \53812 , \53810 );
and \U$53436 ( \53813 , \53812 , \7206 );
nor \U$53437 ( \53814 , \53811 , \53813 );
not \U$53438 ( \53815 , \53814 );
and \U$53439 ( \53816 , \53807 , \53815 );
and \U$53440 ( \53817 , \53806 , \53814 );
nor \U$53441 ( \53818 , \53816 , \53817 );
not \U$53442 ( \53819 , \53818 );
and \U$53443 ( \53820 , \53787 , \53819 );
and \U$53444 ( \53821 , \53818 , \53786 );
and \U$53445 ( \53822 , \4688 , RIae76cd0_60);
and \U$53446 ( \53823 , RIae77108_69, \4686 );
nor \U$53447 ( \53824 , \53822 , \53823 );
and \U$53448 ( \53825 , \53824 , \4482 );
not \U$53449 ( \53826 , \53824 );
and \U$53450 ( \53827 , \53826 , \4481 );
nor \U$53451 ( \53828 , \53825 , \53827 );
not \U$53452 ( \53829 , \53828 );
and \U$53453 ( \53830 , \5399 , RIae77090_68);
and \U$53454 ( \53831 , RIae77270_72, \5397 );
nor \U$53455 ( \53832 , \53830 , \53831 );
and \U$53456 ( \53833 , \53832 , \5016 );
not \U$53457 ( \53834 , \53832 );
and \U$53458 ( \53835 , \53834 , \5403 );
nor \U$53459 ( \53836 , \53833 , \53835 );
not \U$53460 ( \53837 , \53836 );
or \U$53461 ( \53838 , \53829 , \53837 );
or \U$53462 ( \53839 , \53828 , \53836 );
nand \U$53463 ( \53840 , \53838 , \53839 );
not \U$53464 ( \53841 , \53840 );
and \U$53465 ( \53842 , \4247 , RIae76eb0_64);
and \U$53466 ( \53843 , RIae76dc0_62, \4245 );
nor \U$53467 ( \53844 , \53842 , \53843 );
and \U$53468 ( \53845 , \53844 , \4251 );
not \U$53469 ( \53846 , \53844 );
and \U$53470 ( \53847 , \53846 , \3989 );
nor \U$53471 ( \53848 , \53845 , \53847 );
not \U$53472 ( \53849 , \53848 );
and \U$53473 ( \53850 , \53841 , \53849 );
and \U$53474 ( \53851 , \53840 , \53848 );
nor \U$53475 ( \53852 , \53850 , \53851 );
nor \U$53476 ( \53853 , \53821 , \53852 );
nor \U$53477 ( \53854 , \53820 , \53853 );
nor \U$53478 ( \53855 , \53755 , \53854 );
nor \U$53479 ( \53856 , \53754 , \53855 );
xor \U$53480 ( \53857 , \53651 , \53856 );
and \U$53481 ( \53858 , \2783 , RIae77ae0_90);
and \U$53482 ( \53859 , RIae779f0_88, \2781 );
nor \U$53483 ( \53860 , \53858 , \53859 );
not \U$53484 ( \53861 , \53860 );
not \U$53485 ( \53862 , \3089 );
and \U$53486 ( \53863 , \53861 , \53862 );
and \U$53487 ( \53864 , \53860 , \3089 );
nor \U$53488 ( \53865 , \53863 , \53864 );
not \U$53489 ( \53866 , \53865 );
not \U$53490 ( \53867 , \2774 );
and \U$53491 ( \53868 , \3214 , RIae77810_84);
and \U$53492 ( \53869 , RIae77900_86, \3212 );
nor \U$53493 ( \53870 , \53868 , \53869 );
not \U$53494 ( \53871 , \53870 );
or \U$53495 ( \53872 , \53867 , \53871 );
or \U$53496 ( \53873 , \53870 , \3218 );
nand \U$53497 ( \53874 , \53872 , \53873 );
not \U$53498 ( \53875 , \53874 );
or \U$53499 ( \53876 , \53866 , \53875 );
or \U$53500 ( \53877 , \53865 , \53874 );
nand \U$53501 ( \53878 , \53876 , \53877 );
not \U$53502 ( \53879 , \53878 );
and \U$53503 ( \53880 , \2607 , RIae776a8_81);
and \U$53504 ( \53881 , RIae77450_76, \2605 );
nor \U$53505 ( \53882 , \53880 , \53881 );
and \U$53506 ( \53883 , \53882 , \2397 );
not \U$53507 ( \53884 , \53882 );
and \U$53508 ( \53885 , \53884 , \2611 );
nor \U$53509 ( \53886 , \53883 , \53885 );
not \U$53510 ( \53887 , \53886 );
and \U$53511 ( \53888 , \53879 , \53887 );
and \U$53512 ( \53889 , \53878 , \53886 );
nor \U$53513 ( \53890 , \53888 , \53889 );
not \U$53514 ( \53891 , \53890 );
and \U$53515 ( \53892 , \6172 , RIae77f90_100);
and \U$53516 ( \53893 , RIae78080_102, \6170 );
nor \U$53517 ( \53894 , \53892 , \53893 );
and \U$53518 ( \53895 , \53894 , \6176 );
not \U$53519 ( \53896 , \53894 );
and \U$53520 ( \53897 , \53896 , \6175 );
nor \U$53521 ( \53898 , \53895 , \53897 );
and \U$53522 ( \53899 , \5399 , RIae77270_72);
and \U$53523 ( \53900 , RIae77360_74, \5397 );
nor \U$53524 ( \53901 , \53899 , \53900 );
and \U$53525 ( \53902 , \53901 , \5016 );
not \U$53526 ( \53903 , \53901 );
and \U$53527 ( \53904 , \53903 , \5403 );
nor \U$53528 ( \53905 , \53902 , \53904 );
xor \U$53529 ( \53906 , \53898 , \53905 );
and \U$53530 ( \53907 , \5896 , RIae78350_108);
and \U$53531 ( \53908 , RIae78170_104, \5894 );
nor \U$53532 ( \53909 , \53907 , \53908 );
and \U$53533 ( \53910 , \53909 , \5590 );
not \U$53534 ( \53911 , \53909 );
and \U$53535 ( \53912 , \53911 , \5589 );
nor \U$53536 ( \53913 , \53910 , \53912 );
xor \U$53537 ( \53914 , \53906 , \53913 );
not \U$53538 ( \53915 , \53914 );
or \U$53539 ( \53916 , \53891 , \53915 );
or \U$53540 ( \53917 , \53890 , \53914 );
nand \U$53541 ( \53918 , \53916 , \53917 );
not \U$53542 ( \53919 , \53918 );
and \U$53543 ( \53920 , \4247 , RIae76dc0_62);
and \U$53544 ( \53921 , RIae76cd0_60, \4245 );
nor \U$53545 ( \53922 , \53920 , \53921 );
and \U$53546 ( \53923 , \53922 , \4251 );
not \U$53547 ( \53924 , \53922 );
and \U$53548 ( \53925 , \53924 , \3989 );
nor \U$53549 ( \53926 , \53923 , \53925 );
and \U$53550 ( \53927 , \4688 , RIae77108_69);
and \U$53551 ( \53928 , RIae77090_68, \4686 );
nor \U$53552 ( \53929 , \53927 , \53928 );
and \U$53553 ( \53930 , \53929 , \4482 );
not \U$53554 ( \53931 , \53929 );
and \U$53555 ( \53932 , \53931 , \4481 );
nor \U$53556 ( \53933 , \53930 , \53932 );
xor \U$53557 ( \53934 , \53926 , \53933 );
and \U$53558 ( \53935 , \3730 , RIae76fa0_66);
and \U$53559 ( \53936 , RIae76eb0_64, \3728 );
nor \U$53560 ( \53937 , \53935 , \53936 );
and \U$53561 ( \53938 , \53937 , \3422 );
not \U$53562 ( \53939 , \53937 );
and \U$53563 ( \53940 , \53939 , \3732 );
nor \U$53564 ( \53941 , \53938 , \53940 );
xor \U$53565 ( \53942 , \53934 , \53941 );
not \U$53566 ( \53943 , \53942 );
and \U$53567 ( \53944 , \53919 , \53943 );
and \U$53568 ( \53945 , \53918 , \53942 );
nor \U$53569 ( \53946 , \53944 , \53945 );
not \U$53570 ( \53947 , \53946 );
xor \U$53571 ( \53948 , \53628 , \53636 );
and \U$53572 ( \53949 , \53948 , \53644 );
and \U$53573 ( \53950 , \53628 , \53636 );
or \U$53574 ( \53951 , \53949 , \53950 );
and \U$53575 ( \53952 , \53611 , \53618 );
xnor \U$53576 ( \53953 , \53951 , \53952 );
not \U$53577 ( \53954 , \53953 );
and \U$53578 ( \53955 , \2224 , RIae77630_80);
and \U$53579 ( \53956 , RIae77540_78, \2222 );
nor \U$53580 ( \53957 , \53955 , \53956 );
and \U$53581 ( \53958 , \53957 , \2061 );
not \U$53582 ( \53959 , \53957 );
and \U$53583 ( \53960 , \53959 , \2060 );
nor \U$53584 ( \53961 , \53958 , \53960 );
not \U$53585 ( \53962 , \53961 );
and \U$53586 ( \53963 , \53954 , \53962 );
and \U$53587 ( \53964 , \53953 , \53961 );
nor \U$53588 ( \53965 , \53963 , \53964 );
not \U$53589 ( \53966 , \53965 );
and \U$53590 ( \53967 , \53947 , \53966 );
and \U$53591 ( \53968 , \53946 , \53965 );
and \U$53592 ( \53969 , \8371 , RIae77cc0_94);
and \U$53593 ( \53970 , RIae77bd0_92, \8369 );
nor \U$53594 ( \53971 , \53969 , \53970 );
and \U$53595 ( \53972 , \53971 , \8019 );
not \U$53596 ( \53973 , \53971 );
and \U$53597 ( \53974 , \53973 , \8020 );
nor \U$53598 ( \53975 , \53972 , \53974 );
not \U$53599 ( \53976 , \53975 );
and \U$53600 ( \53977 , \7633 , RIae78440_110);
and \U$53601 ( \53978 , RIae784b8_111, \7631 );
nor \U$53602 ( \53979 , \53977 , \53978 );
and \U$53603 ( \53980 , \53979 , \7206 );
not \U$53604 ( \53981 , \53979 );
and \U$53605 ( \53982 , \53981 , \7205 );
nor \U$53606 ( \53983 , \53980 , \53982 );
not \U$53607 ( \53984 , \53983 );
or \U$53608 ( \53985 , \53976 , \53984 );
or \U$53609 ( \53986 , \53975 , \53983 );
nand \U$53610 ( \53987 , \53985 , \53986 );
not \U$53611 ( \53988 , \53987 );
and \U$53612 ( \53989 , \6941 , RIae78260_106);
and \U$53613 ( \53990 , RIae78620_114, \6939 );
nor \U$53614 ( \53991 , \53989 , \53990 );
and \U$53615 ( \53992 , \53991 , \6945 );
not \U$53616 ( \53993 , \53991 );
and \U$53617 ( \53994 , \53993 , \6314 );
nor \U$53618 ( \53995 , \53992 , \53994 );
not \U$53619 ( \53996 , \53995 );
and \U$53620 ( \53997 , \53988 , \53996 );
and \U$53621 ( \53998 , \53987 , \53995 );
nor \U$53622 ( \53999 , \53997 , \53998 );
not \U$53623 ( \54000 , \53999 );
and \U$53624 ( \54001 , \11470 , RIae75bf0_24);
and \U$53625 ( \54002 , RIae75b00_22, \11468 );
nor \U$53626 ( \54003 , \54001 , \54002 );
and \U$53627 ( \54004 , \54003 , \10936 );
not \U$53628 ( \54005 , \54003 );
and \U$53629 ( \54006 , \54005 , \11474 );
nor \U$53630 ( \54007 , \54004 , \54006 );
and \U$53631 ( \54008 , \12180 , RIae75a10_20);
and \U$53632 ( \54009 , RIae75920_18, \12178 );
nor \U$53633 ( \54010 , \54008 , \54009 );
and \U$53634 ( \54011 , \54010 , \12184 );
not \U$53635 ( \54012 , \54010 );
and \U$53636 ( \54013 , \54012 , \11827 );
nor \U$53637 ( \54014 , \54011 , \54013 );
xor \U$53638 ( \54015 , \54007 , \54014 );
and \U$53639 ( \54016 , \13059 , RIae75fb0_32);
and \U$53640 ( \54017 , RIae75ec0_30, \13057 );
nor \U$53641 ( \54018 , \54016 , \54017 );
and \U$53642 ( \54019 , \54018 , \13063 );
not \U$53643 ( \54020 , \54018 );
and \U$53644 ( \54021 , \54020 , \12718 );
nor \U$53645 ( \54022 , \54019 , \54021 );
xor \U$53646 ( \54023 , \54015 , \54022 );
not \U$53647 ( \54024 , \54023 );
or \U$53648 ( \54025 , \54000 , \54024 );
or \U$53649 ( \54026 , \53999 , \54023 );
nand \U$53650 ( \54027 , \54025 , \54026 );
not \U$53651 ( \54028 , \54027 );
and \U$53652 ( \54029 , \9760 , RIae789e0_122);
and \U$53653 ( \54030 , RIae788f0_120, \9758 );
nor \U$53654 ( \54031 , \54029 , \54030 );
and \U$53655 ( \54032 , \54031 , \9272 );
not \U$53656 ( \54033 , \54031 );
and \U$53657 ( \54034 , \54033 , \9273 );
nor \U$53658 ( \54035 , \54032 , \54034 );
and \U$53659 ( \54036 , \10548 , RIae78800_118);
and \U$53660 ( \54037 , RIae78710_116, \10546 );
nor \U$53661 ( \54038 , \54036 , \54037 );
and \U$53662 ( \54039 , \54038 , \10118 );
not \U$53663 ( \54040 , \54038 );
and \U$53664 ( \54041 , \54040 , \10421 );
nor \U$53665 ( \54042 , \54039 , \54041 );
xor \U$53666 ( \54043 , \54035 , \54042 );
and \U$53667 ( \54044 , \8966 , RIae77db0_96);
and \U$53668 ( \54045 , RIae77ea0_98, \8964 );
nor \U$53669 ( \54046 , \54044 , \54045 );
and \U$53670 ( \54047 , \54046 , \8789 );
not \U$53671 ( \54048 , \54046 );
and \U$53672 ( \54049 , \54048 , \8799 );
nor \U$53673 ( \54050 , \54047 , \54049 );
xor \U$53674 ( \54051 , \54043 , \54050 );
not \U$53675 ( \54052 , \54051 );
and \U$53676 ( \54053 , \54028 , \54052 );
and \U$53677 ( \54054 , \54027 , \54051 );
nor \U$53678 ( \54055 , \54053 , \54054 );
nor \U$53679 ( \54056 , \53968 , \54055 );
nor \U$53680 ( \54057 , \53967 , \54056 );
xor \U$53681 ( \54058 , \53857 , \54057 );
not \U$53682 ( \54059 , \54058 );
or \U$53683 ( \54060 , \53814 , \53794 );
not \U$53684 ( \54061 , \53794 );
not \U$53685 ( \54062 , \53814 );
or \U$53686 ( \54063 , \54061 , \54062 );
nand \U$53687 ( \54064 , \54063 , \53802 );
nand \U$53688 ( \54065 , \54060 , \54064 );
or \U$53689 ( \54066 , \53848 , \53828 );
not \U$53690 ( \54067 , \53828 );
not \U$53691 ( \54068 , \53848 );
or \U$53692 ( \54069 , \54067 , \54068 );
nand \U$53693 ( \54070 , \54069 , \53836 );
nand \U$53694 ( \54071 , \54066 , \54070 );
xor \U$53695 ( \54072 , \54065 , \54071 );
or \U$53696 ( \54073 , \53782 , \53762 );
not \U$53697 ( \54074 , \53762 );
not \U$53698 ( \54075 , \53782 );
or \U$53699 ( \54076 , \54074 , \54075 );
nand \U$53700 ( \54077 , \54076 , \53770 );
nand \U$53701 ( \54078 , \54073 , \54077 );
xor \U$53702 ( \54079 , \54072 , \54078 );
xor \U$53703 ( \54080 , \53658 , \53665 );
and \U$53704 ( \54081 , \54080 , \53673 );
and \U$53705 ( \54082 , \53658 , \53665 );
or \U$53706 ( \54083 , \54081 , \54082 );
xor \U$53707 ( \54084 , \53681 , \2060 );
and \U$53708 ( \54085 , \54084 , \53689 );
and \U$53709 ( \54086 , \53681 , \2060 );
or \U$53710 ( \54087 , \54085 , \54086 );
xor \U$53711 ( \54088 , \54083 , \54087 );
xor \U$53712 ( \54089 , \53698 , \53705 );
and \U$53713 ( \54090 , \54089 , \53713 );
and \U$53714 ( \54091 , \53698 , \53705 );
or \U$53715 ( \54092 , \54090 , \54091 );
xor \U$53716 ( \54093 , \54088 , \54092 );
xor \U$53717 ( \54094 , \54079 , \54093 );
not \U$53718 ( \54095 , \53946 );
xor \U$53719 ( \54096 , \53965 , \54055 );
not \U$53720 ( \54097 , \54096 );
or \U$53721 ( \54098 , \54095 , \54097 );
or \U$53722 ( \54099 , \54096 , \53946 );
nand \U$53723 ( \54100 , \54098 , \54099 );
and \U$53724 ( \54101 , \54094 , \54100 );
and \U$53725 ( \54102 , \54079 , \54093 );
or \U$53726 ( \54103 , \54101 , \54102 );
xor \U$53727 ( \54104 , \54083 , \54087 );
and \U$53728 ( \54105 , \54104 , \54092 );
and \U$53729 ( \54106 , \54083 , \54087 );
or \U$53730 ( \54107 , \54105 , \54106 );
not \U$53731 ( \54108 , \53961 );
not \U$53732 ( \54109 , \53952 );
or \U$53733 ( \54110 , \54108 , \54109 );
or \U$53734 ( \54111 , \53952 , \53961 );
nand \U$53735 ( \54112 , \54111 , \53951 );
nand \U$53736 ( \54113 , \54110 , \54112 );
xor \U$53737 ( \54114 , \54107 , \54113 );
xor \U$53738 ( \54115 , \54065 , \54071 );
and \U$53739 ( \54116 , \54115 , \54078 );
and \U$53740 ( \54117 , \54065 , \54071 );
or \U$53741 ( \54118 , \54116 , \54117 );
xor \U$53742 ( \54119 , \54114 , \54118 );
xor \U$53743 ( \54120 , \54103 , \54119 );
xor \U$53744 ( \54121 , \53445 , \53470 );
xor \U$53745 ( \54122 , \54121 , \53496 );
xor \U$53746 ( \54123 , \53606 , \53619 );
xor \U$53747 ( \54124 , \54123 , \53645 );
and \U$53748 ( \54125 , \54122 , \54124 );
not \U$53749 ( \54126 , \53786 );
xor \U$53750 ( \54127 , \53852 , \53818 );
not \U$53751 ( \54128 , \54127 );
or \U$53752 ( \54129 , \54126 , \54128 );
or \U$53753 ( \54130 , \54127 , \53786 );
nand \U$53754 ( \54131 , \54129 , \54130 );
xor \U$53755 ( \54132 , \53606 , \53619 );
xor \U$53756 ( \54133 , \54132 , \53645 );
and \U$53757 ( \54134 , \54131 , \54133 );
and \U$53758 ( \54135 , \54122 , \54131 );
or \U$53759 ( \54136 , \54125 , \54134 , \54135 );
and \U$53760 ( \54137 , \5896 , RIae77090_68);
and \U$53761 ( \54138 , RIae77270_72, \5894 );
nor \U$53762 ( \54139 , \54137 , \54138 );
and \U$53763 ( \54140 , \54139 , \5590 );
not \U$53764 ( \54141 , \54139 );
and \U$53765 ( \54142 , \54141 , \5589 );
nor \U$53766 ( \54143 , \54140 , \54142 );
and \U$53767 ( \54144 , \6172 , RIae77360_74);
and \U$53768 ( \54145 , RIae78350_108, \6170 );
nor \U$53769 ( \54146 , \54144 , \54145 );
and \U$53770 ( \54147 , \54146 , \6176 );
not \U$53771 ( \54148 , \54146 );
and \U$53772 ( \54149 , \54148 , \6175 );
nor \U$53773 ( \54150 , \54147 , \54149 );
xor \U$53774 ( \54151 , \54143 , \54150 );
and \U$53775 ( \54152 , \6941 , RIae78170_104);
and \U$53776 ( \54153 , RIae77f90_100, \6939 );
nor \U$53777 ( \54154 , \54152 , \54153 );
and \U$53778 ( \54155 , \54154 , \6314 );
not \U$53779 ( \54156 , \54154 );
and \U$53780 ( \54157 , \54156 , \6945 );
nor \U$53781 ( \54158 , \54155 , \54157 );
and \U$53782 ( \54159 , \54151 , \54158 );
and \U$53783 ( \54160 , \54143 , \54150 );
or \U$53784 ( \54161 , \54159 , \54160 );
and \U$53785 ( \54162 , \4247 , RIae77900_86);
and \U$53786 ( \54163 , RIae76fa0_66, \4245 );
nor \U$53787 ( \54164 , \54162 , \54163 );
and \U$53788 ( \54165 , \54164 , \3989 );
not \U$53789 ( \54166 , \54164 );
and \U$53790 ( \54167 , \54166 , \4251 );
nor \U$53791 ( \54168 , \54165 , \54167 );
and \U$53792 ( \54169 , \4688 , RIae76eb0_64);
and \U$53793 ( \54170 , RIae76dc0_62, \4686 );
nor \U$53794 ( \54171 , \54169 , \54170 );
and \U$53795 ( \54172 , \54171 , \4481 );
not \U$53796 ( \54173 , \54171 );
and \U$53797 ( \54174 , \54173 , \4482 );
nor \U$53798 ( \54175 , \54172 , \54174 );
xor \U$53799 ( \54176 , \54168 , \54175 );
and \U$53800 ( \54177 , \5399 , RIae76cd0_60);
and \U$53801 ( \54178 , RIae77108_69, \5397 );
nor \U$53802 ( \54179 , \54177 , \54178 );
and \U$53803 ( \54180 , \54179 , \5016 );
not \U$53804 ( \54181 , \54179 );
and \U$53805 ( \54182 , \54181 , \5403 );
nor \U$53806 ( \54183 , \54180 , \54182 );
and \U$53807 ( \54184 , \54176 , \54183 );
and \U$53808 ( \54185 , \54168 , \54175 );
or \U$53809 ( \54186 , \54184 , \54185 );
xor \U$53810 ( \54187 , \54161 , \54186 );
and \U$53811 ( \54188 , \7633 , RIae78080_102);
and \U$53812 ( \54189 , RIae78260_106, \7631 );
nor \U$53813 ( \54190 , \54188 , \54189 );
and \U$53814 ( \54191 , \54190 , \7206 );
not \U$53815 ( \54192 , \54190 );
and \U$53816 ( \54193 , \54192 , \7205 );
nor \U$53817 ( \54194 , \54191 , \54193 );
and \U$53818 ( \54195 , \8371 , RIae78620_114);
and \U$53819 ( \54196 , RIae78440_110, \8369 );
nor \U$53820 ( \54197 , \54195 , \54196 );
and \U$53821 ( \54198 , \54197 , \8020 );
not \U$53822 ( \54199 , \54197 );
and \U$53823 ( \54200 , \54199 , \8019 );
nor \U$53824 ( \54201 , \54198 , \54200 );
xor \U$53825 ( \54202 , \54194 , \54201 );
and \U$53826 ( \54203 , \8966 , RIae784b8_111);
and \U$53827 ( \54204 , RIae77cc0_94, \8964 );
nor \U$53828 ( \54205 , \54203 , \54204 );
and \U$53829 ( \54206 , \54205 , \8799 );
not \U$53830 ( \54207 , \54205 );
and \U$53831 ( \54208 , \54207 , \8789 );
nor \U$53832 ( \54209 , \54206 , \54208 );
and \U$53833 ( \54210 , \54202 , \54209 );
and \U$53834 ( \54211 , \54194 , \54201 );
or \U$53835 ( \54212 , \54210 , \54211 );
and \U$53836 ( \54213 , \54187 , \54212 );
and \U$53837 ( \54214 , \54161 , \54186 );
or \U$53838 ( \54215 , \54213 , \54214 );
and \U$53839 ( \54216 , \9760 , RIae77bd0_92);
and \U$53840 ( \54217 , RIae77db0_96, \9758 );
nor \U$53841 ( \54218 , \54216 , \54217 );
and \U$53842 ( \54219 , \54218 , \9273 );
not \U$53843 ( \54220 , \54218 );
and \U$53844 ( \54221 , \54220 , \9764 );
nor \U$53845 ( \54222 , \54219 , \54221 );
and \U$53846 ( \54223 , \10548 , RIae77ea0_98);
and \U$53847 ( \54224 , RIae789e0_122, \10546 );
nor \U$53848 ( \54225 , \54223 , \54224 );
and \U$53849 ( \54226 , \54225 , \10421 );
not \U$53850 ( \54227 , \54225 );
and \U$53851 ( \54228 , \54227 , \10118 );
nor \U$53852 ( \54229 , \54226 , \54228 );
xor \U$53853 ( \54230 , \54222 , \54229 );
and \U$53854 ( \54231 , \11470 , RIae788f0_120);
and \U$53855 ( \54232 , RIae78800_118, \11468 );
nor \U$53856 ( \54233 , \54231 , \54232 );
and \U$53857 ( \54234 , \54233 , \10936 );
not \U$53858 ( \54235 , \54233 );
and \U$53859 ( \54236 , \54235 , \11474 );
nor \U$53860 ( \54237 , \54234 , \54236 );
and \U$53861 ( \54238 , \54230 , \54237 );
and \U$53862 ( \54239 , \54222 , \54229 );
or \U$53863 ( \54240 , \54238 , \54239 );
and \U$53864 ( \54241 , \15726 , RIae75dd0_28);
and \U$53865 ( \54242 , RIae75650_12, RIae7aab0_192);
nor \U$53866 ( \54243 , \54241 , \54242 );
and \U$53867 ( \54244 , \54243 , \14959 );
not \U$53868 ( \54245 , \54243 );
and \U$53869 ( \54246 , \54245 , RIae7aa38_191);
nor \U$53870 ( \54247 , \54244 , \54246 );
xor \U$53871 ( \54248 , \54247 , \2397 );
and \U$53872 ( \54249 , \14964 , RIae75ec0_30);
and \U$53873 ( \54250 , RIae75ce0_26, \14962 );
nor \U$53874 ( \54251 , \54249 , \54250 );
and \U$53875 ( \54252 , \54251 , \14463 );
not \U$53876 ( \54253 , \54251 );
and \U$53877 ( \54254 , \54253 , \14462 );
nor \U$53878 ( \54255 , \54252 , \54254 );
and \U$53879 ( \54256 , \54248 , \54255 );
and \U$53880 ( \54257 , \54247 , \2397 );
or \U$53881 ( \54258 , \54256 , \54257 );
xor \U$53882 ( \54259 , \54240 , \54258 );
and \U$53883 ( \54260 , \12180 , RIae78710_116);
and \U$53884 ( \54261 , RIae75bf0_24, \12178 );
nor \U$53885 ( \54262 , \54260 , \54261 );
and \U$53886 ( \54263 , \54262 , \12184 );
not \U$53887 ( \54264 , \54262 );
and \U$53888 ( \54265 , \54264 , \11827 );
nor \U$53889 ( \54266 , \54263 , \54265 );
and \U$53890 ( \54267 , \13059 , RIae75b00_22);
and \U$53891 ( \54268 , RIae75a10_20, \13057 );
nor \U$53892 ( \54269 , \54267 , \54268 );
and \U$53893 ( \54270 , \54269 , \13063 );
not \U$53894 ( \54271 , \54269 );
and \U$53895 ( \54272 , \54271 , \12718 );
nor \U$53896 ( \54273 , \54270 , \54272 );
xor \U$53897 ( \54274 , \54266 , \54273 );
and \U$53898 ( \54275 , \14059 , RIae75920_18);
and \U$53899 ( \54276 , RIae75fb0_32, \14057 );
nor \U$53900 ( \54277 , \54275 , \54276 );
and \U$53901 ( \54278 , \54277 , \13502 );
not \U$53902 ( \54279 , \54277 );
and \U$53903 ( \54280 , \54279 , \14063 );
nor \U$53904 ( \54281 , \54278 , \54280 );
and \U$53905 ( \54282 , \54274 , \54281 );
and \U$53906 ( \54283 , \54266 , \54273 );
or \U$53907 ( \54284 , \54282 , \54283 );
and \U$53908 ( \54285 , \54259 , \54284 );
and \U$53909 ( \54286 , \54240 , \54258 );
or \U$53910 ( \54287 , \54285 , \54286 );
xor \U$53911 ( \54288 , \54215 , \54287 );
and \U$53912 ( \54289 , \3730 , RIae779f0_88);
and \U$53913 ( \54290 , RIae77810_84, \3728 );
nor \U$53914 ( \54291 , \54289 , \54290 );
and \U$53915 ( \54292 , \54291 , \3732 );
not \U$53916 ( \54293 , \54291 );
and \U$53917 ( \54294 , \54293 , \3422 );
nor \U$53918 ( \54295 , \54292 , \54294 );
not \U$53919 ( \54296 , \3089 );
and \U$53920 ( \54297 , \2783 , RIae77540_78);
and \U$53921 ( \54298 , RIae776a8_81, \2781 );
nor \U$53922 ( \54299 , \54297 , \54298 );
not \U$53923 ( \54300 , \54299 );
or \U$53924 ( \54301 , \54296 , \54300 );
or \U$53925 ( \54302 , \54299 , \3089 );
nand \U$53926 ( \54303 , \54301 , \54302 );
xor \U$53927 ( \54304 , \54295 , \54303 );
not \U$53928 ( \54305 , \2774 );
and \U$53929 ( \54306 , \3214 , RIae77450_76);
and \U$53930 ( \54307 , RIae77ae0_90, \3212 );
nor \U$53931 ( \54308 , \54306 , \54307 );
not \U$53932 ( \54309 , \54308 );
or \U$53933 ( \54310 , \54305 , \54309 );
or \U$53934 ( \54311 , \54308 , \2774 );
nand \U$53935 ( \54312 , \54310 , \54311 );
and \U$53936 ( \54313 , \54304 , \54312 );
and \U$53937 ( \54314 , \54295 , \54303 );
or \U$53938 ( \54315 , \54313 , \54314 );
xor \U$53939 ( \54316 , \53587 , \53594 );
xor \U$53940 ( \54317 , \54316 , \53603 );
and \U$53941 ( \54318 , \54315 , \54317 );
xor \U$53942 ( \54319 , \53452 , \53459 );
xor \U$53943 ( \54320 , \54319 , \53467 );
xor \U$53944 ( \54321 , \53587 , \53594 );
xor \U$53945 ( \54322 , \54321 , \53603 );
and \U$53946 ( \54323 , \54320 , \54322 );
and \U$53947 ( \54324 , \54315 , \54320 );
or \U$53948 ( \54325 , \54318 , \54323 , \54324 );
and \U$53949 ( \54326 , \54288 , \54325 );
and \U$53950 ( \54327 , \54215 , \54287 );
or \U$53951 ( \54328 , \54326 , \54327 );
xor \U$53952 ( \54329 , \54136 , \54328 );
xor \U$53953 ( \54330 , \53427 , \53434 );
xor \U$53954 ( \54331 , \54330 , \53442 );
xor \U$53955 ( \54332 , \53506 , \53513 );
xor \U$53956 ( \54333 , \54332 , \53521 );
and \U$53957 ( \54334 , \54331 , \54333 );
xor \U$53958 ( \54335 , \53478 , \53485 );
xor \U$53959 ( \54336 , \54335 , \53493 );
xor \U$53960 ( \54337 , \53506 , \53513 );
xor \U$53961 ( \54338 , \54337 , \53521 );
and \U$53962 ( \54339 , \54336 , \54338 );
and \U$53963 ( \54340 , \54331 , \54336 );
or \U$53964 ( \54341 , \54334 , \54339 , \54340 );
xor \U$53965 ( \54342 , \53557 , \53564 );
xor \U$53966 ( \54343 , \54342 , \53572 );
xor \U$53967 ( \54344 , \53531 , \53538 );
xor \U$53968 ( \54345 , \54344 , \53546 );
and \U$53969 ( \54346 , \54343 , \54345 );
xor \U$53970 ( \54347 , \54341 , \54346 );
xor \U$53971 ( \54348 , \53681 , \2060 );
xor \U$53972 ( \54349 , \54348 , \53689 );
xor \U$53973 ( \54350 , \53674 , \53714 );
xor \U$53974 ( \54351 , \54349 , \54350 );
and \U$53975 ( \54352 , \54347 , \54351 );
and \U$53976 ( \54353 , \54341 , \54346 );
or \U$53977 ( \54354 , \54352 , \54353 );
and \U$53978 ( \54355 , \54329 , \54354 );
and \U$53979 ( \54356 , \54136 , \54328 );
or \U$53980 ( \54357 , \54355 , \54356 );
xor \U$53981 ( \54358 , \54120 , \54357 );
not \U$53982 ( \54359 , \54358 );
or \U$53983 ( \54360 , \54059 , \54359 );
or \U$53984 ( \54361 , \54358 , \54058 );
nand \U$53985 ( \54362 , \54360 , \54361 );
xor \U$53986 ( \54363 , \53499 , \53578 );
xor \U$53987 ( \54364 , \54363 , \53648 );
xor \U$53988 ( \54365 , \54079 , \54093 );
xor \U$53989 ( \54366 , \54365 , \54100 );
and \U$53990 ( \54367 , \54364 , \54366 );
xor \U$53991 ( \54368 , \54136 , \54328 );
xor \U$53992 ( \54369 , \54368 , \54354 );
xor \U$53993 ( \54370 , \54079 , \54093 );
xor \U$53994 ( \54371 , \54370 , \54100 );
and \U$53995 ( \54372 , \54369 , \54371 );
and \U$53996 ( \54373 , \54364 , \54369 );
or \U$53997 ( \54374 , \54367 , \54372 , \54373 );
or \U$53998 ( \54375 , \53999 , \54051 );
not \U$53999 ( \54376 , \54051 );
not \U$54000 ( \54377 , \53999 );
or \U$54001 ( \54378 , \54376 , \54377 );
nand \U$54002 ( \54379 , \54378 , \54023 );
nand \U$54003 ( \54380 , \54375 , \54379 );
or \U$54004 ( \54381 , \53890 , \53942 );
not \U$54005 ( \54382 , \53942 );
not \U$54006 ( \54383 , \53890 );
or \U$54007 ( \54384 , \54382 , \54383 );
nand \U$54008 ( \54385 , \54384 , \53914 );
nand \U$54009 ( \54386 , \54381 , \54385 );
xor \U$54010 ( \54387 , \54380 , \54386 );
and \U$54011 ( \54388 , \15726 , RIae75740_14);
and \U$54012 ( \54389 , RIae75290_4, RIae7aab0_192);
nor \U$54013 ( \54390 , \54388 , \54389 );
and \U$54014 ( \54391 , \54390 , \14959 );
not \U$54015 ( \54392 , \54390 );
and \U$54016 ( \54393 , \54392 , RIae7aa38_191);
nor \U$54017 ( \54394 , \54391 , \54393 );
xor \U$54018 ( \54395 , \54394 , \1734 );
and \U$54019 ( \54396 , \14964 , RIae75560_10);
and \U$54020 ( \54397 , RIae75830_16, \14962 );
nor \U$54021 ( \54398 , \54396 , \54397 );
and \U$54022 ( \54399 , \54398 , \14463 );
not \U$54023 ( \54400 , \54398 );
and \U$54024 ( \54401 , \54400 , \14462 );
nor \U$54025 ( \54402 , \54399 , \54401 );
xor \U$54026 ( \54403 , \54395 , \54402 );
and \U$54027 ( \54404 , \12180 , RIae75920_18);
and \U$54028 ( \54405 , RIae75fb0_32, \12178 );
nor \U$54029 ( \54406 , \54404 , \54405 );
and \U$54030 ( \54407 , \54406 , \12184 );
not \U$54031 ( \54408 , \54406 );
and \U$54032 ( \54409 , \54408 , \11827 );
nor \U$54033 ( \54410 , \54407 , \54409 );
and \U$54034 ( \54411 , \13059 , RIae75ec0_30);
and \U$54035 ( \54412 , RIae75ce0_26, \13057 );
nor \U$54036 ( \54413 , \54411 , \54412 );
and \U$54037 ( \54414 , \54413 , \13063 );
not \U$54038 ( \54415 , \54413 );
and \U$54039 ( \54416 , \54415 , \12718 );
nor \U$54040 ( \54417 , \54414 , \54416 );
xor \U$54041 ( \54418 , \54410 , \54417 );
and \U$54042 ( \54419 , \14059 , RIae75dd0_28);
and \U$54043 ( \54420 , RIae75650_12, \14057 );
nor \U$54044 ( \54421 , \54419 , \54420 );
and \U$54045 ( \54422 , \54421 , \13502 );
not \U$54046 ( \54423 , \54421 );
and \U$54047 ( \54424 , \54423 , \14063 );
nor \U$54048 ( \54425 , \54422 , \54424 );
xor \U$54049 ( \54426 , \54418 , \54425 );
and \U$54050 ( \54427 , \11470 , RIae75b00_22);
and \U$54051 ( \54428 , RIae75a10_20, \11468 );
nor \U$54052 ( \54429 , \54427 , \54428 );
and \U$54053 ( \54430 , \54429 , \10936 );
not \U$54054 ( \54431 , \54429 );
and \U$54055 ( \54432 , \54431 , \11474 );
nor \U$54056 ( \54433 , \54430 , \54432 );
and \U$54057 ( \54434 , \9760 , RIae788f0_120);
and \U$54058 ( \54435 , RIae78800_118, \9758 );
nor \U$54059 ( \54436 , \54434 , \54435 );
and \U$54060 ( \54437 , \54436 , \9273 );
not \U$54061 ( \54438 , \54436 );
and \U$54062 ( \54439 , \54438 , \9272 );
nor \U$54063 ( \54440 , \54437 , \54439 );
xor \U$54064 ( \54441 , \54433 , \54440 );
and \U$54065 ( \54442 , \10548 , RIae78710_116);
and \U$54066 ( \54443 , RIae75bf0_24, \10546 );
nor \U$54067 ( \54444 , \54442 , \54443 );
and \U$54068 ( \54445 , \54444 , \10421 );
not \U$54069 ( \54446 , \54444 );
and \U$54070 ( \54447 , \54446 , \10118 );
nor \U$54071 ( \54448 , \54445 , \54447 );
xor \U$54072 ( \54449 , \54441 , \54448 );
xor \U$54073 ( \54450 , \54426 , \54449 );
xor \U$54074 ( \54451 , \54403 , \54450 );
xor \U$54075 ( \54452 , \54387 , \54451 );
xor \U$54076 ( \54453 , \54035 , \54042 );
and \U$54077 ( \54454 , \54453 , \54050 );
and \U$54078 ( \54455 , \54035 , \54042 );
nor \U$54079 ( \54456 , \54454 , \54455 );
or \U$54080 ( \54457 , \53748 , \53728 );
not \U$54081 ( \54458 , \53728 );
not \U$54082 ( \54459 , \53748 );
or \U$54083 ( \54460 , \54458 , \54459 );
nand \U$54084 ( \54461 , \54460 , \53736 );
nand \U$54085 ( \54462 , \54457 , \54461 );
xor \U$54086 ( \54463 , \54456 , \54462 );
xor \U$54087 ( \54464 , \54007 , \54014 );
and \U$54088 ( \54465 , \54464 , \54022 );
and \U$54089 ( \54466 , \54007 , \54014 );
or \U$54090 ( \54467 , \54465 , \54466 );
xor \U$54091 ( \54468 , \54463 , \54467 );
and \U$54092 ( \54469 , \6941 , RIae78620_114);
and \U$54093 ( \54470 , RIae78440_110, \6939 );
nor \U$54094 ( \54471 , \54469 , \54470 );
and \U$54095 ( \54472 , \54471 , \6314 );
not \U$54096 ( \54473 , \54471 );
and \U$54097 ( \54474 , \54473 , \6945 );
nor \U$54098 ( \54475 , \54472 , \54474 );
and \U$54099 ( \54476 , \5896 , RIae78170_104);
and \U$54100 ( \54477 , RIae77f90_100, \5894 );
nor \U$54101 ( \54478 , \54476 , \54477 );
and \U$54102 ( \54479 , \54478 , \5590 );
not \U$54103 ( \54480 , \54478 );
and \U$54104 ( \54481 , \54480 , \5589 );
nor \U$54105 ( \54482 , \54479 , \54481 );
xor \U$54106 ( \54483 , \54475 , \54482 );
and \U$54107 ( \54484 , \6172 , RIae78080_102);
and \U$54108 ( \54485 , RIae78260_106, \6170 );
nor \U$54109 ( \54486 , \54484 , \54485 );
and \U$54110 ( \54487 , \54486 , \6176 );
not \U$54111 ( \54488 , \54486 );
and \U$54112 ( \54489 , \54488 , \6175 );
nor \U$54113 ( \54490 , \54487 , \54489 );
xor \U$54114 ( \54491 , \54483 , \54490 );
and \U$54115 ( \54492 , \8966 , RIae77ea0_98);
and \U$54116 ( \54493 , RIae789e0_122, \8964 );
nor \U$54117 ( \54494 , \54492 , \54493 );
and \U$54118 ( \54495 , \54494 , \8799 );
not \U$54119 ( \54496 , \54494 );
and \U$54120 ( \54497 , \54496 , \8789 );
nor \U$54121 ( \54498 , \54495 , \54497 );
and \U$54122 ( \54499 , \7633 , RIae784b8_111);
and \U$54123 ( \54500 , RIae77cc0_94, \7631 );
nor \U$54124 ( \54501 , \54499 , \54500 );
and \U$54125 ( \54502 , \54501 , \7206 );
not \U$54126 ( \54503 , \54501 );
and \U$54127 ( \54504 , \54503 , \7205 );
nor \U$54128 ( \54505 , \54502 , \54504 );
xor \U$54129 ( \54506 , \54498 , \54505 );
and \U$54130 ( \54507 , \8371 , RIae77bd0_92);
and \U$54131 ( \54508 , RIae77db0_96, \8369 );
nor \U$54132 ( \54509 , \54507 , \54508 );
and \U$54133 ( \54510 , \54509 , \8020 );
not \U$54134 ( \54511 , \54509 );
and \U$54135 ( \54512 , \54511 , \8019 );
nor \U$54136 ( \54513 , \54510 , \54512 );
xor \U$54137 ( \54514 , \54506 , \54513 );
and \U$54138 ( \54515 , \4247 , RIae76cd0_60);
and \U$54139 ( \54516 , RIae77108_69, \4245 );
nor \U$54140 ( \54517 , \54515 , \54516 );
and \U$54141 ( \54518 , \54517 , \3989 );
not \U$54142 ( \54519 , \54517 );
and \U$54143 ( \54520 , \54519 , \4251 );
nor \U$54144 ( \54521 , \54518 , \54520 );
and \U$54145 ( \54522 , \4688 , RIae77090_68);
and \U$54146 ( \54523 , RIae77270_72, \4686 );
nor \U$54147 ( \54524 , \54522 , \54523 );
and \U$54148 ( \54525 , \54524 , \4481 );
not \U$54149 ( \54526 , \54524 );
and \U$54150 ( \54527 , \54526 , \4482 );
nor \U$54151 ( \54528 , \54525 , \54527 );
xor \U$54152 ( \54529 , \54521 , \54528 );
and \U$54153 ( \54530 , \5399 , RIae77360_74);
and \U$54154 ( \54531 , RIae78350_108, \5397 );
nor \U$54155 ( \54532 , \54530 , \54531 );
and \U$54156 ( \54533 , \54532 , \5016 );
not \U$54157 ( \54534 , \54532 );
and \U$54158 ( \54535 , \54534 , \5403 );
nor \U$54159 ( \54536 , \54533 , \54535 );
xor \U$54160 ( \54537 , \54529 , \54536 );
xor \U$54161 ( \54538 , \54514 , \54537 );
xor \U$54162 ( \54539 , \54491 , \54538 );
or \U$54163 ( \54540 , \53995 , \53975 );
not \U$54164 ( \54541 , \53975 );
not \U$54165 ( \54542 , \53995 );
or \U$54166 ( \54543 , \54541 , \54542 );
nand \U$54167 ( \54544 , \54543 , \53983 );
nand \U$54168 ( \54545 , \54540 , \54544 );
xor \U$54169 ( \54546 , \53898 , \53905 );
and \U$54170 ( \54547 , \54546 , \53913 );
and \U$54171 ( \54548 , \53898 , \53905 );
or \U$54172 ( \54549 , \54547 , \54548 );
xor \U$54173 ( \54550 , \54545 , \54549 );
xor \U$54174 ( \54551 , \53926 , \53933 );
and \U$54175 ( \54552 , \54551 , \53941 );
and \U$54176 ( \54553 , \53926 , \53933 );
nor \U$54177 ( \54554 , \54552 , \54553 );
xor \U$54178 ( \54555 , \54550 , \54554 );
xor \U$54179 ( \54556 , \54539 , \54555 );
and \U$54180 ( \54557 , \2224 , RIae77540_78);
and \U$54181 ( \54558 , RIae776a8_81, \2222 );
nor \U$54182 ( \54559 , \54557 , \54558 );
and \U$54183 ( \54560 , \54559 , \2061 );
not \U$54184 ( \54561 , \54559 );
and \U$54185 ( \54562 , \54561 , \2060 );
nor \U$54186 ( \54563 , \54560 , \54562 );
nand \U$54187 ( \54564 , RIae77630_80, \1937 );
and \U$54188 ( \54565 , \54564 , \1735 );
not \U$54189 ( \54566 , \54564 );
and \U$54190 ( \54567 , \54566 , \1734 );
nor \U$54191 ( \54568 , \54565 , \54567 );
xor \U$54192 ( \54569 , \54563 , \54568 );
and \U$54193 ( \54570 , \2607 , RIae77450_76);
and \U$54194 ( \54571 , RIae77ae0_90, \2605 );
nor \U$54195 ( \54572 , \54570 , \54571 );
and \U$54196 ( \54573 , \54572 , \2611 );
not \U$54197 ( \54574 , \54572 );
and \U$54198 ( \54575 , \54574 , \2397 );
nor \U$54199 ( \54576 , \54573 , \54575 );
xor \U$54200 ( \54577 , \54569 , \54576 );
or \U$54201 ( \54578 , \53886 , \53865 );
not \U$54202 ( \54579 , \53865 );
not \U$54203 ( \54580 , \53886 );
or \U$54204 ( \54581 , \54579 , \54580 );
nand \U$54205 ( \54582 , \54581 , \53874 );
nand \U$54206 ( \54583 , \54578 , \54582 );
not \U$54207 ( \54584 , \2789 );
and \U$54208 ( \54585 , \2783 , RIae779f0_88);
and \U$54209 ( \54586 , RIae77810_84, \2781 );
nor \U$54210 ( \54587 , \54585 , \54586 );
not \U$54211 ( \54588 , \54587 );
or \U$54212 ( \54589 , \54584 , \54588 );
or \U$54213 ( \54590 , \54587 , \3089 );
nand \U$54214 ( \54591 , \54589 , \54590 );
not \U$54215 ( \54592 , \3218 );
and \U$54216 ( \54593 , \3214 , RIae77900_86);
and \U$54217 ( \54594 , RIae76fa0_66, \3212 );
nor \U$54218 ( \54595 , \54593 , \54594 );
not \U$54219 ( \54596 , \54595 );
or \U$54220 ( \54597 , \54592 , \54596 );
or \U$54221 ( \54598 , \54595 , \3218 );
nand \U$54222 ( \54599 , \54597 , \54598 );
xor \U$54223 ( \54600 , \54591 , \54599 );
and \U$54224 ( \54601 , \3730 , RIae76eb0_64);
and \U$54225 ( \54602 , RIae76dc0_62, \3728 );
nor \U$54226 ( \54603 , \54601 , \54602 );
and \U$54227 ( \54604 , \54603 , \3732 );
not \U$54228 ( \54605 , \54603 );
and \U$54229 ( \54606 , \54605 , \3422 );
nor \U$54230 ( \54607 , \54604 , \54606 );
xor \U$54231 ( \54608 , \54600 , \54607 );
xor \U$54232 ( \54609 , \54583 , \54608 );
xor \U$54233 ( \54610 , \54577 , \54609 );
xor \U$54234 ( \54611 , \54556 , \54610 );
xor \U$54235 ( \54612 , \54468 , \54611 );
xor \U$54236 ( \54613 , \54452 , \54612 );
xor \U$54237 ( \54614 , \54374 , \54613 );
xor \U$54238 ( \54615 , \54161 , \54186 );
xor \U$54239 ( \54616 , \54615 , \54212 );
xor \U$54240 ( \54617 , \54240 , \54258 );
xor \U$54241 ( \54618 , \54617 , \54284 );
xor \U$54242 ( \54619 , \54616 , \54618 );
xor \U$54243 ( \54620 , \53587 , \53594 );
xor \U$54244 ( \54621 , \54620 , \53603 );
xor \U$54245 ( \54622 , \54315 , \54320 );
xor \U$54246 ( \54623 , \54621 , \54622 );
and \U$54247 ( \54624 , \54619 , \54623 );
and \U$54248 ( \54625 , \54616 , \54618 );
or \U$54249 ( \54626 , \54624 , \54625 );
and \U$54250 ( \54627 , \7633 , RIae77f90_100);
and \U$54251 ( \54628 , RIae78080_102, \7631 );
nor \U$54252 ( \54629 , \54627 , \54628 );
and \U$54253 ( \54630 , \54629 , \7206 );
not \U$54254 ( \54631 , \54629 );
and \U$54255 ( \54632 , \54631 , \7205 );
nor \U$54256 ( \54633 , \54630 , \54632 );
and \U$54257 ( \54634 , \6941 , RIae78350_108);
and \U$54258 ( \54635 , RIae78170_104, \6939 );
nor \U$54259 ( \54636 , \54634 , \54635 );
and \U$54260 ( \54637 , \54636 , \6314 );
not \U$54261 ( \54638 , \54636 );
and \U$54262 ( \54639 , \54638 , \6945 );
nor \U$54263 ( \54640 , \54637 , \54639 );
xor \U$54264 ( \54641 , \54633 , \54640 );
and \U$54265 ( \54642 , \8371 , RIae78260_106);
and \U$54266 ( \54643 , RIae78620_114, \8369 );
nor \U$54267 ( \54644 , \54642 , \54643 );
and \U$54268 ( \54645 , \54644 , \8020 );
not \U$54269 ( \54646 , \54644 );
and \U$54270 ( \54647 , \54646 , \8019 );
nor \U$54271 ( \54648 , \54645 , \54647 );
and \U$54272 ( \54649 , \54641 , \54648 );
and \U$54273 ( \54650 , \54633 , \54640 );
or \U$54274 ( \54651 , \54649 , \54650 );
and \U$54275 ( \54652 , \5896 , RIae77108_69);
and \U$54276 ( \54653 , RIae77090_68, \5894 );
nor \U$54277 ( \54654 , \54652 , \54653 );
and \U$54278 ( \54655 , \54654 , \5590 );
not \U$54279 ( \54656 , \54654 );
and \U$54280 ( \54657 , \54656 , \5589 );
nor \U$54281 ( \54658 , \54655 , \54657 );
and \U$54282 ( \54659 , \5399 , RIae76dc0_62);
and \U$54283 ( \54660 , RIae76cd0_60, \5397 );
nor \U$54284 ( \54661 , \54659 , \54660 );
and \U$54285 ( \54662 , \54661 , \5016 );
not \U$54286 ( \54663 , \54661 );
and \U$54287 ( \54664 , \54663 , \5403 );
nor \U$54288 ( \54665 , \54662 , \54664 );
xor \U$54289 ( \54666 , \54658 , \54665 );
and \U$54290 ( \54667 , \6172 , RIae77270_72);
and \U$54291 ( \54668 , RIae77360_74, \6170 );
nor \U$54292 ( \54669 , \54667 , \54668 );
and \U$54293 ( \54670 , \54669 , \6176 );
not \U$54294 ( \54671 , \54669 );
and \U$54295 ( \54672 , \54671 , \6175 );
nor \U$54296 ( \54673 , \54670 , \54672 );
and \U$54297 ( \54674 , \54666 , \54673 );
and \U$54298 ( \54675 , \54658 , \54665 );
or \U$54299 ( \54676 , \54674 , \54675 );
xor \U$54300 ( \54677 , \54651 , \54676 );
and \U$54301 ( \54678 , \4688 , RIae76fa0_66);
and \U$54302 ( \54679 , RIae76eb0_64, \4686 );
nor \U$54303 ( \54680 , \54678 , \54679 );
and \U$54304 ( \54681 , \54680 , \4481 );
not \U$54305 ( \54682 , \54680 );
and \U$54306 ( \54683 , \54682 , \4482 );
nor \U$54307 ( \54684 , \54681 , \54683 );
and \U$54308 ( \54685 , \3730 , RIae77ae0_90);
and \U$54309 ( \54686 , RIae779f0_88, \3728 );
nor \U$54310 ( \54687 , \54685 , \54686 );
and \U$54311 ( \54688 , \54687 , \3732 );
not \U$54312 ( \54689 , \54687 );
and \U$54313 ( \54690 , \54689 , \3422 );
nor \U$54314 ( \54691 , \54688 , \54690 );
xor \U$54315 ( \54692 , \54684 , \54691 );
and \U$54316 ( \54693 , \4247 , RIae77810_84);
and \U$54317 ( \54694 , RIae77900_86, \4245 );
nor \U$54318 ( \54695 , \54693 , \54694 );
and \U$54319 ( \54696 , \54695 , \3989 );
not \U$54320 ( \54697 , \54695 );
and \U$54321 ( \54698 , \54697 , \4251 );
nor \U$54322 ( \54699 , \54696 , \54698 );
and \U$54323 ( \54700 , \54692 , \54699 );
and \U$54324 ( \54701 , \54684 , \54691 );
or \U$54325 ( \54702 , \54700 , \54701 );
and \U$54326 ( \54703 , \54677 , \54702 );
and \U$54327 ( \54704 , \54651 , \54676 );
or \U$54328 ( \54705 , \54703 , \54704 );
and \U$54329 ( \54706 , \13059 , RIae75bf0_24);
and \U$54330 ( \54707 , RIae75b00_22, \13057 );
nor \U$54331 ( \54708 , \54706 , \54707 );
and \U$54332 ( \54709 , \54708 , \13063 );
not \U$54333 ( \54710 , \54708 );
and \U$54334 ( \54711 , \54710 , \12718 );
nor \U$54335 ( \54712 , \54709 , \54711 );
and \U$54336 ( \54713 , \11470 , RIae789e0_122);
and \U$54337 ( \54714 , RIae788f0_120, \11468 );
nor \U$54338 ( \54715 , \54713 , \54714 );
and \U$54339 ( \54716 , \54715 , \10936 );
not \U$54340 ( \54717 , \54715 );
and \U$54341 ( \54718 , \54717 , \11474 );
nor \U$54342 ( \54719 , \54716 , \54718 );
xor \U$54343 ( \54720 , \54712 , \54719 );
and \U$54344 ( \54721 , \12180 , RIae78800_118);
and \U$54345 ( \54722 , RIae78710_116, \12178 );
nor \U$54346 ( \54723 , \54721 , \54722 );
and \U$54347 ( \54724 , \54723 , \12184 );
not \U$54348 ( \54725 , \54723 );
and \U$54349 ( \54726 , \54725 , \11827 );
nor \U$54350 ( \54727 , \54724 , \54726 );
and \U$54351 ( \54728 , \54720 , \54727 );
and \U$54352 ( \54729 , \54712 , \54719 );
or \U$54353 ( \54730 , \54728 , \54729 );
and \U$54354 ( \54731 , \14964 , RIae75fb0_32);
and \U$54355 ( \54732 , RIae75ec0_30, \14962 );
nor \U$54356 ( \54733 , \54731 , \54732 );
and \U$54357 ( \54734 , \54733 , \14463 );
not \U$54358 ( \54735 , \54733 );
and \U$54359 ( \54736 , \54735 , \14462 );
nor \U$54360 ( \54737 , \54734 , \54736 );
and \U$54361 ( \54738 , \15726 , RIae75ce0_26);
and \U$54362 ( \54739 , RIae75dd0_28, RIae7aab0_192);
nor \U$54363 ( \54740 , \54738 , \54739 );
and \U$54364 ( \54741 , \54740 , \14959 );
not \U$54365 ( \54742 , \54740 );
and \U$54366 ( \54743 , \54742 , RIae7aa38_191);
nor \U$54367 ( \54744 , \54741 , \54743 );
xor \U$54368 ( \54745 , \54737 , \54744 );
and \U$54369 ( \54746 , \14059 , RIae75a10_20);
and \U$54370 ( \54747 , RIae75920_18, \14057 );
nor \U$54371 ( \54748 , \54746 , \54747 );
and \U$54372 ( \54749 , \54748 , \13502 );
not \U$54373 ( \54750 , \54748 );
and \U$54374 ( \54751 , \54750 , \14063 );
nor \U$54375 ( \54752 , \54749 , \54751 );
and \U$54376 ( \54753 , \54745 , \54752 );
and \U$54377 ( \54754 , \54737 , \54744 );
or \U$54378 ( \54755 , \54753 , \54754 );
xor \U$54379 ( \54756 , \54730 , \54755 );
and \U$54380 ( \54757 , \8966 , RIae78440_110);
and \U$54381 ( \54758 , RIae784b8_111, \8964 );
nor \U$54382 ( \54759 , \54757 , \54758 );
and \U$54383 ( \54760 , \54759 , \8799 );
not \U$54384 ( \54761 , \54759 );
and \U$54385 ( \54762 , \54761 , \8789 );
nor \U$54386 ( \54763 , \54760 , \54762 );
and \U$54387 ( \54764 , \9760 , RIae77cc0_94);
and \U$54388 ( \54765 , RIae77bd0_92, \9758 );
nor \U$54389 ( \54766 , \54764 , \54765 );
and \U$54390 ( \54767 , \54766 , \9273 );
not \U$54391 ( \54768 , \54766 );
and \U$54392 ( \54769 , \54768 , \9272 );
nor \U$54393 ( \54770 , \54767 , \54769 );
xor \U$54394 ( \54771 , \54763 , \54770 );
and \U$54395 ( \54772 , \10548 , RIae77db0_96);
and \U$54396 ( \54773 , RIae77ea0_98, \10546 );
nor \U$54397 ( \54774 , \54772 , \54773 );
and \U$54398 ( \54775 , \54774 , \10421 );
not \U$54399 ( \54776 , \54774 );
and \U$54400 ( \54777 , \54776 , \10118 );
nor \U$54401 ( \54778 , \54775 , \54777 );
and \U$54402 ( \54779 , \54771 , \54778 );
and \U$54403 ( \54780 , \54763 , \54770 );
or \U$54404 ( \54781 , \54779 , \54780 );
and \U$54405 ( \54782 , \54756 , \54781 );
and \U$54406 ( \54783 , \54730 , \54755 );
or \U$54407 ( \54784 , \54782 , \54783 );
xor \U$54408 ( \54785 , \54705 , \54784 );
xor \U$54409 ( \54786 , \54295 , \54303 );
xor \U$54410 ( \54787 , \54786 , \54312 );
nand \U$54411 ( \54788 , RIae77630_80, \2605 );
and \U$54412 ( \54789 , \54788 , \2611 );
not \U$54413 ( \54790 , \54788 );
and \U$54414 ( \54791 , \54790 , \2397 );
nor \U$54415 ( \54792 , \54789 , \54791 );
xor \U$54416 ( \54793 , \54787 , \54792 );
xor \U$54417 ( \54794 , \54168 , \54175 );
xor \U$54418 ( \54795 , \54794 , \54183 );
and \U$54419 ( \54796 , \54793 , \54795 );
and \U$54420 ( \54797 , \54787 , \54792 );
or \U$54421 ( \54798 , \54796 , \54797 );
and \U$54422 ( \54799 , \54785 , \54798 );
and \U$54423 ( \54800 , \54705 , \54784 );
or \U$54424 ( \54801 , \54799 , \54800 );
xor \U$54425 ( \54802 , \54626 , \54801 );
xor \U$54426 ( \54803 , \54143 , \54150 );
xor \U$54427 ( \54804 , \54803 , \54158 );
xor \U$54428 ( \54805 , \54194 , \54201 );
xor \U$54429 ( \54806 , \54805 , \54209 );
and \U$54430 ( \54807 , \54804 , \54806 );
xor \U$54431 ( \54808 , \54222 , \54229 );
xor \U$54432 ( \54809 , \54808 , \54237 );
xor \U$54433 ( \54810 , \54194 , \54201 );
xor \U$54434 ( \54811 , \54810 , \54209 );
and \U$54435 ( \54812 , \54809 , \54811 );
and \U$54436 ( \54813 , \54804 , \54809 );
or \U$54437 ( \54814 , \54807 , \54812 , \54813 );
xor \U$54438 ( \54815 , \54343 , \54345 );
xor \U$54439 ( \54816 , \54814 , \54815 );
xor \U$54440 ( \54817 , \53506 , \53513 );
xor \U$54441 ( \54818 , \54817 , \53521 );
xor \U$54442 ( \54819 , \54331 , \54336 );
xor \U$54443 ( \54820 , \54818 , \54819 );
and \U$54444 ( \54821 , \54816 , \54820 );
and \U$54445 ( \54822 , \54814 , \54815 );
or \U$54446 ( \54823 , \54821 , \54822 );
and \U$54447 ( \54824 , \54802 , \54823 );
and \U$54448 ( \54825 , \54626 , \54801 );
or \U$54449 ( \54826 , \54824 , \54825 );
not \U$54450 ( \54827 , \53752 );
xor \U$54451 ( \54828 , \53854 , \53720 );
not \U$54452 ( \54829 , \54828 );
or \U$54453 ( \54830 , \54827 , \54829 );
or \U$54454 ( \54831 , \54828 , \53752 );
nand \U$54455 ( \54832 , \54830 , \54831 );
xor \U$54456 ( \54833 , \54826 , \54832 );
xor \U$54457 ( \54834 , \53524 , \53549 );
xor \U$54458 ( \54835 , \54834 , \53575 );
xor \U$54459 ( \54836 , \54341 , \54346 );
xor \U$54460 ( \54837 , \54836 , \54351 );
and \U$54461 ( \54838 , \54835 , \54837 );
xor \U$54462 ( \54839 , \53606 , \53619 );
xor \U$54463 ( \54840 , \54839 , \53645 );
xor \U$54464 ( \54841 , \54122 , \54131 );
xor \U$54465 ( \54842 , \54840 , \54841 );
xor \U$54466 ( \54843 , \54341 , \54346 );
xor \U$54467 ( \54844 , \54843 , \54351 );
and \U$54468 ( \54845 , \54842 , \54844 );
and \U$54469 ( \54846 , \54835 , \54842 );
or \U$54470 ( \54847 , \54838 , \54845 , \54846 );
and \U$54471 ( \54848 , \54833 , \54847 );
and \U$54472 ( \54849 , \54826 , \54832 );
or \U$54473 ( \54850 , \54848 , \54849 );
xor \U$54474 ( \54851 , \54614 , \54850 );
xor \U$54475 ( \54852 , \54362 , \54851 );
xor \U$54476 ( \54853 , \54712 , \54719 );
xor \U$54477 ( \54854 , \54853 , \54727 );
xor \U$54478 ( \54855 , \54737 , \54744 );
xor \U$54479 ( \54856 , \54855 , \54752 );
xor \U$54480 ( \54857 , \54854 , \54856 );
xor \U$54481 ( \54858 , \54763 , \54770 );
xor \U$54482 ( \54859 , \54858 , \54778 );
and \U$54483 ( \54860 , \54857 , \54859 );
and \U$54484 ( \54861 , \54854 , \54856 );
or \U$54485 ( \54862 , \54860 , \54861 );
xor \U$54486 ( \54863 , \54266 , \54273 );
xor \U$54487 ( \54864 , \54863 , \54281 );
xor \U$54488 ( \54865 , \54862 , \54864 );
xor \U$54489 ( \54866 , \54684 , \54691 );
xor \U$54490 ( \54867 , \54866 , \54699 );
xor \U$54491 ( \54868 , \54658 , \54665 );
xor \U$54492 ( \54869 , \54868 , \54673 );
and \U$54493 ( \54870 , \54867 , \54869 );
xor \U$54494 ( \54871 , \54633 , \54640 );
xor \U$54495 ( \54872 , \54871 , \54648 );
xor \U$54496 ( \54873 , \54658 , \54665 );
xor \U$54497 ( \54874 , \54873 , \54673 );
and \U$54498 ( \54875 , \54872 , \54874 );
and \U$54499 ( \54876 , \54867 , \54872 );
or \U$54500 ( \54877 , \54870 , \54875 , \54876 );
and \U$54501 ( \54878 , \54865 , \54877 );
and \U$54502 ( \54879 , \54862 , \54864 );
or \U$54503 ( \54880 , \54878 , \54879 );
and \U$54504 ( \54881 , \13059 , RIae78710_116);
and \U$54505 ( \54882 , RIae75bf0_24, \13057 );
nor \U$54506 ( \54883 , \54881 , \54882 );
and \U$54507 ( \54884 , \54883 , \13063 );
not \U$54508 ( \54885 , \54883 );
and \U$54509 ( \54886 , \54885 , \12718 );
nor \U$54510 ( \54887 , \54884 , \54886 );
and \U$54511 ( \54888 , \12180 , RIae788f0_120);
and \U$54512 ( \54889 , RIae78800_118, \12178 );
nor \U$54513 ( \54890 , \54888 , \54889 );
and \U$54514 ( \54891 , \54890 , \12184 );
not \U$54515 ( \54892 , \54890 );
and \U$54516 ( \54893 , \54892 , \11827 );
nor \U$54517 ( \54894 , \54891 , \54893 );
xor \U$54518 ( \54895 , \54887 , \54894 );
and \U$54519 ( \54896 , \14059 , RIae75b00_22);
and \U$54520 ( \54897 , RIae75a10_20, \14057 );
nor \U$54521 ( \54898 , \54896 , \54897 );
and \U$54522 ( \54899 , \54898 , \13502 );
not \U$54523 ( \54900 , \54898 );
and \U$54524 ( \54901 , \54900 , \14063 );
nor \U$54525 ( \54902 , \54899 , \54901 );
and \U$54526 ( \54903 , \54895 , \54902 );
and \U$54527 ( \54904 , \54887 , \54894 );
or \U$54528 ( \54905 , \54903 , \54904 );
and \U$54529 ( \54906 , \15726 , RIae75ec0_30);
and \U$54530 ( \54907 , RIae75ce0_26, RIae7aab0_192);
nor \U$54531 ( \54908 , \54906 , \54907 );
and \U$54532 ( \54909 , \54908 , \14959 );
not \U$54533 ( \54910 , \54908 );
and \U$54534 ( \54911 , \54910 , RIae7aa38_191);
nor \U$54535 ( \54912 , \54909 , \54911 );
xor \U$54536 ( \54913 , \54912 , \2789 );
and \U$54537 ( \54914 , \14964 , RIae75920_18);
and \U$54538 ( \54915 , RIae75fb0_32, \14962 );
nor \U$54539 ( \54916 , \54914 , \54915 );
and \U$54540 ( \54917 , \54916 , \14463 );
not \U$54541 ( \54918 , \54916 );
and \U$54542 ( \54919 , \54918 , \14462 );
nor \U$54543 ( \54920 , \54917 , \54919 );
and \U$54544 ( \54921 , \54913 , \54920 );
and \U$54545 ( \54922 , \54912 , \2789 );
or \U$54546 ( \54923 , \54921 , \54922 );
xor \U$54547 ( \54924 , \54905 , \54923 );
and \U$54548 ( \54925 , \11470 , RIae77ea0_98);
and \U$54549 ( \54926 , RIae789e0_122, \11468 );
nor \U$54550 ( \54927 , \54925 , \54926 );
and \U$54551 ( \54928 , \54927 , \10936 );
not \U$54552 ( \54929 , \54927 );
and \U$54553 ( \54930 , \54929 , \11474 );
nor \U$54554 ( \54931 , \54928 , \54930 );
and \U$54555 ( \54932 , \9760 , RIae784b8_111);
and \U$54556 ( \54933 , RIae77cc0_94, \9758 );
nor \U$54557 ( \54934 , \54932 , \54933 );
and \U$54558 ( \54935 , \54934 , \9273 );
not \U$54559 ( \54936 , \54934 );
and \U$54560 ( \54937 , \54936 , \9272 );
nor \U$54561 ( \54938 , \54935 , \54937 );
xor \U$54562 ( \54939 , \54931 , \54938 );
and \U$54563 ( \54940 , \10548 , RIae77bd0_92);
and \U$54564 ( \54941 , RIae77db0_96, \10546 );
nor \U$54565 ( \54942 , \54940 , \54941 );
and \U$54566 ( \54943 , \54942 , \10421 );
not \U$54567 ( \54944 , \54942 );
and \U$54568 ( \54945 , \54944 , \10118 );
nor \U$54569 ( \54946 , \54943 , \54945 );
and \U$54570 ( \54947 , \54939 , \54946 );
and \U$54571 ( \54948 , \54931 , \54938 );
or \U$54572 ( \54949 , \54947 , \54948 );
and \U$54573 ( \54950 , \54924 , \54949 );
and \U$54574 ( \54951 , \54905 , \54923 );
or \U$54575 ( \54952 , \54950 , \54951 );
not \U$54576 ( \54953 , \2774 );
and \U$54577 ( \54954 , \3214 , RIae776a8_81);
and \U$54578 ( \54955 , RIae77450_76, \3212 );
nor \U$54579 ( \54956 , \54954 , \54955 );
not \U$54580 ( \54957 , \54956 );
or \U$54581 ( \54958 , \54953 , \54957 );
or \U$54582 ( \54959 , \54956 , \3218 );
nand \U$54583 ( \54960 , \54958 , \54959 );
not \U$54584 ( \54961 , \3089 );
and \U$54585 ( \54962 , \2783 , RIae77630_80);
and \U$54586 ( \54963 , RIae77540_78, \2781 );
nor \U$54587 ( \54964 , \54962 , \54963 );
not \U$54588 ( \54965 , \54964 );
or \U$54589 ( \54966 , \54961 , \54965 );
or \U$54590 ( \54967 , \54964 , \3089 );
nand \U$54591 ( \54968 , \54966 , \54967 );
xor \U$54592 ( \54969 , \54960 , \54968 );
and \U$54593 ( \54970 , \3730 , RIae77450_76);
and \U$54594 ( \54971 , RIae77ae0_90, \3728 );
nor \U$54595 ( \54972 , \54970 , \54971 );
and \U$54596 ( \54973 , \54972 , \3732 );
not \U$54597 ( \54974 , \54972 );
and \U$54598 ( \54975 , \54974 , \3421 );
nor \U$54599 ( \54976 , \54973 , \54975 );
nand \U$54600 ( \54977 , RIae77630_80, \2781 );
not \U$54601 ( \54978 , \54977 );
not \U$54602 ( \54979 , \2789 );
or \U$54603 ( \54980 , \54978 , \54979 );
or \U$54604 ( \54981 , \2789 , \54977 );
nand \U$54605 ( \54982 , \54980 , \54981 );
xor \U$54606 ( \54983 , \54976 , \54982 );
not \U$54607 ( \54984 , \2774 );
and \U$54608 ( \54985 , \3214 , RIae77540_78);
and \U$54609 ( \54986 , RIae776a8_81, \3212 );
nor \U$54610 ( \54987 , \54985 , \54986 );
not \U$54611 ( \54988 , \54987 );
or \U$54612 ( \54989 , \54984 , \54988 );
or \U$54613 ( \54990 , \54987 , \3218 );
nand \U$54614 ( \54991 , \54989 , \54990 );
and \U$54615 ( \54992 , \54983 , \54991 );
and \U$54616 ( \54993 , \54976 , \54982 );
or \U$54617 ( \54994 , \54992 , \54993 );
and \U$54618 ( \54995 , \54969 , \54994 );
and \U$54619 ( \54996 , \54960 , \54968 );
or \U$54620 ( \54997 , \54995 , \54996 );
xor \U$54621 ( \54998 , \54952 , \54997 );
and \U$54622 ( \54999 , \5896 , RIae76cd0_60);
and \U$54623 ( \55000 , RIae77108_69, \5894 );
nor \U$54624 ( \55001 , \54999 , \55000 );
and \U$54625 ( \55002 , \55001 , \5590 );
not \U$54626 ( \55003 , \55001 );
and \U$54627 ( \55004 , \55003 , \5589 );
nor \U$54628 ( \55005 , \55002 , \55004 );
and \U$54629 ( \55006 , \6172 , RIae77090_68);
and \U$54630 ( \55007 , RIae77270_72, \6170 );
nor \U$54631 ( \55008 , \55006 , \55007 );
and \U$54632 ( \55009 , \55008 , \6176 );
not \U$54633 ( \55010 , \55008 );
and \U$54634 ( \55011 , \55010 , \6175 );
nor \U$54635 ( \55012 , \55009 , \55011 );
xor \U$54636 ( \55013 , \55005 , \55012 );
and \U$54637 ( \55014 , \6941 , RIae77360_74);
and \U$54638 ( \55015 , RIae78350_108, \6939 );
nor \U$54639 ( \55016 , \55014 , \55015 );
and \U$54640 ( \55017 , \55016 , \6314 );
not \U$54641 ( \55018 , \55016 );
and \U$54642 ( \55019 , \55018 , \6945 );
nor \U$54643 ( \55020 , \55017 , \55019 );
and \U$54644 ( \55021 , \55013 , \55020 );
and \U$54645 ( \55022 , \55005 , \55012 );
or \U$54646 ( \55023 , \55021 , \55022 );
and \U$54647 ( \55024 , \5399 , RIae76eb0_64);
and \U$54648 ( \55025 , RIae76dc0_62, \5397 );
nor \U$54649 ( \55026 , \55024 , \55025 );
and \U$54650 ( \55027 , \55026 , \5016 );
not \U$54651 ( \55028 , \55026 );
and \U$54652 ( \55029 , \55028 , \5403 );
nor \U$54653 ( \55030 , \55027 , \55029 );
and \U$54654 ( \55031 , \4247 , RIae779f0_88);
and \U$54655 ( \55032 , RIae77810_84, \4245 );
nor \U$54656 ( \55033 , \55031 , \55032 );
and \U$54657 ( \55034 , \55033 , \3989 );
not \U$54658 ( \55035 , \55033 );
and \U$54659 ( \55036 , \55035 , \4251 );
nor \U$54660 ( \55037 , \55034 , \55036 );
xor \U$54661 ( \55038 , \55030 , \55037 );
and \U$54662 ( \55039 , \4688 , RIae77900_86);
and \U$54663 ( \55040 , RIae76fa0_66, \4686 );
nor \U$54664 ( \55041 , \55039 , \55040 );
and \U$54665 ( \55042 , \55041 , \4481 );
not \U$54666 ( \55043 , \55041 );
and \U$54667 ( \55044 , \55043 , \4482 );
nor \U$54668 ( \55045 , \55042 , \55044 );
and \U$54669 ( \55046 , \55038 , \55045 );
and \U$54670 ( \55047 , \55030 , \55037 );
or \U$54671 ( \55048 , \55046 , \55047 );
xor \U$54672 ( \55049 , \55023 , \55048 );
and \U$54673 ( \55050 , \8371 , RIae78080_102);
and \U$54674 ( \55051 , RIae78260_106, \8369 );
nor \U$54675 ( \55052 , \55050 , \55051 );
and \U$54676 ( \55053 , \55052 , \8020 );
not \U$54677 ( \55054 , \55052 );
and \U$54678 ( \55055 , \55054 , \8019 );
nor \U$54679 ( \55056 , \55053 , \55055 );
and \U$54680 ( \55057 , \7633 , RIae78170_104);
and \U$54681 ( \55058 , RIae77f90_100, \7631 );
nor \U$54682 ( \55059 , \55057 , \55058 );
and \U$54683 ( \55060 , \55059 , \7206 );
not \U$54684 ( \55061 , \55059 );
and \U$54685 ( \55062 , \55061 , \7205 );
nor \U$54686 ( \55063 , \55060 , \55062 );
xor \U$54687 ( \55064 , \55056 , \55063 );
and \U$54688 ( \55065 , \8966 , RIae78620_114);
and \U$54689 ( \55066 , RIae78440_110, \8964 );
nor \U$54690 ( \55067 , \55065 , \55066 );
and \U$54691 ( \55068 , \55067 , \8799 );
not \U$54692 ( \55069 , \55067 );
and \U$54693 ( \55070 , \55069 , \8789 );
nor \U$54694 ( \55071 , \55068 , \55070 );
and \U$54695 ( \55072 , \55064 , \55071 );
and \U$54696 ( \55073 , \55056 , \55063 );
or \U$54697 ( \55074 , \55072 , \55073 );
and \U$54698 ( \55075 , \55049 , \55074 );
and \U$54699 ( \55076 , \55023 , \55048 );
or \U$54700 ( \55077 , \55075 , \55076 );
and \U$54701 ( \55078 , \54998 , \55077 );
and \U$54702 ( \55079 , \54952 , \54997 );
or \U$54703 ( \55080 , \55078 , \55079 );
xor \U$54704 ( \55081 , \54880 , \55080 );
xor \U$54705 ( \55082 , \54247 , \2397 );
xor \U$54706 ( \55083 , \55082 , \54255 );
xor \U$54707 ( \55084 , \54787 , \54792 );
xor \U$54708 ( \55085 , \55084 , \54795 );
and \U$54709 ( \55086 , \55083 , \55085 );
xor \U$54710 ( \55087 , \54194 , \54201 );
xor \U$54711 ( \55088 , \55087 , \54209 );
xor \U$54712 ( \55089 , \54804 , \54809 );
xor \U$54713 ( \55090 , \55088 , \55089 );
xor \U$54714 ( \55091 , \54787 , \54792 );
xor \U$54715 ( \55092 , \55091 , \54795 );
and \U$54716 ( \55093 , \55090 , \55092 );
and \U$54717 ( \55094 , \55083 , \55090 );
or \U$54718 ( \55095 , \55086 , \55093 , \55094 );
and \U$54719 ( \55096 , \55081 , \55095 );
and \U$54720 ( \55097 , \54880 , \55080 );
or \U$54721 ( \55098 , \55096 , \55097 );
xor \U$54722 ( \55099 , \54215 , \54287 );
xor \U$54723 ( \55100 , \55099 , \54325 );
xor \U$54724 ( \55101 , \55098 , \55100 );
xor \U$54725 ( \55102 , \54705 , \54784 );
xor \U$54726 ( \55103 , \55102 , \54798 );
xor \U$54727 ( \55104 , \54616 , \54618 );
xor \U$54728 ( \55105 , \55104 , \54623 );
and \U$54729 ( \55106 , \55103 , \55105 );
xor \U$54730 ( \55107 , \54814 , \54815 );
xor \U$54731 ( \55108 , \55107 , \54820 );
xor \U$54732 ( \55109 , \54616 , \54618 );
xor \U$54733 ( \55110 , \55109 , \54623 );
and \U$54734 ( \55111 , \55108 , \55110 );
and \U$54735 ( \55112 , \55103 , \55108 );
or \U$54736 ( \55113 , \55106 , \55111 , \55112 );
and \U$54737 ( \55114 , \55101 , \55113 );
and \U$54738 ( \55115 , \55098 , \55100 );
or \U$54739 ( \55116 , \55114 , \55115 );
xor \U$54740 ( \55117 , \54626 , \54801 );
xor \U$54741 ( \55118 , \55117 , \54823 );
xor \U$54742 ( \55119 , \54341 , \54346 );
xor \U$54743 ( \55120 , \55119 , \54351 );
xor \U$54744 ( \55121 , \54835 , \54842 );
xor \U$54745 ( \55122 , \55120 , \55121 );
and \U$54746 ( \55123 , \55118 , \55122 );
xor \U$54747 ( \55124 , \55116 , \55123 );
xor \U$54748 ( \55125 , \54079 , \54093 );
xor \U$54749 ( \55126 , \55125 , \54100 );
xor \U$54750 ( \55127 , \54364 , \54369 );
xor \U$54751 ( \55128 , \55126 , \55127 );
and \U$54752 ( \55129 , \55124 , \55128 );
and \U$54753 ( \55130 , \55116 , \55123 );
or \U$54754 ( \55131 , \55129 , \55130 );
and \U$54755 ( \55132 , \54852 , \55131 );
and \U$54756 ( \55133 , \54362 , \54851 );
nor \U$54757 ( \55134 , \55132 , \55133 );
not \U$54758 ( \55135 , \54058 );
nand \U$54759 ( \55136 , \55135 , \54358 );
not \U$54760 ( \55137 , \55136 );
xor \U$54761 ( \55138 , \54374 , \54613 );
and \U$54762 ( \55139 , \55138 , \54850 );
and \U$54763 ( \55140 , \54374 , \54613 );
or \U$54764 ( \55141 , \55139 , \55140 );
not \U$54765 ( \55142 , \55141 );
or \U$54766 ( \55143 , \55137 , \55142 );
or \U$54767 ( \55144 , \55141 , \55136 );
nand \U$54768 ( \55145 , \55143 , \55144 );
not \U$54769 ( \55146 , \55145 );
xor \U$54770 ( \55147 , \54103 , \54119 );
and \U$54771 ( \55148 , \55147 , \54357 );
and \U$54772 ( \55149 , \54103 , \54119 );
or \U$54773 ( \55150 , \55148 , \55149 );
xor \U$54774 ( \55151 , \53651 , \53856 );
and \U$54775 ( \55152 , \55151 , \54057 );
and \U$54776 ( \55153 , \53651 , \53856 );
nor \U$54777 ( \55154 , \55152 , \55153 );
xor \U$54778 ( \55155 , \54545 , \54549 );
and \U$54779 ( \55156 , \55155 , \54554 );
and \U$54780 ( \55157 , \54545 , \54549 );
or \U$54781 ( \55158 , \55156 , \55157 );
xor \U$54782 ( \55159 , \54456 , \54462 );
and \U$54783 ( \55160 , \55159 , \54467 );
and \U$54784 ( \55161 , \54456 , \54462 );
or \U$54785 ( \55162 , \55160 , \55161 );
xor \U$54786 ( \55163 , \55158 , \55162 );
xor \U$54787 ( \55164 , \54563 , \54568 );
xor \U$54788 ( \55165 , \55164 , \54576 );
and \U$54789 ( \55166 , \54583 , \55165 );
xor \U$54790 ( \55167 , \54563 , \54568 );
xor \U$54791 ( \55168 , \55167 , \54576 );
and \U$54792 ( \55169 , \54608 , \55168 );
and \U$54793 ( \55170 , \54583 , \54608 );
or \U$54794 ( \55171 , \55166 , \55169 , \55170 );
xor \U$54795 ( \55172 , \55163 , \55171 );
xor \U$54796 ( \55173 , \55154 , \55172 );
xor \U$54797 ( \55174 , \54380 , \54386 );
xor \U$54798 ( \55175 , \55174 , \54451 );
and \U$54799 ( \55176 , \54468 , \55175 );
xor \U$54800 ( \55177 , \54380 , \54386 );
xor \U$54801 ( \55178 , \55177 , \54451 );
and \U$54802 ( \55179 , \54611 , \55178 );
and \U$54803 ( \55180 , \54468 , \54611 );
or \U$54804 ( \55181 , \55176 , \55179 , \55180 );
xor \U$54805 ( \55182 , \55173 , \55181 );
xnor \U$54806 ( \55183 , \55150 , \55182 );
not \U$54807 ( \55184 , \55183 );
xor \U$54808 ( \55185 , \54539 , \54555 );
and \U$54809 ( \55186 , \55185 , \54610 );
and \U$54810 ( \55187 , \54539 , \54555 );
or \U$54811 ( \55188 , \55186 , \55187 );
xor \U$54812 ( \55189 , \54107 , \54113 );
and \U$54813 ( \55190 , \55189 , \54118 );
and \U$54814 ( \55191 , \54107 , \54113 );
or \U$54815 ( \55192 , \55190 , \55191 );
xor \U$54816 ( \55193 , \55188 , \55192 );
xor \U$54817 ( \55194 , \54380 , \54386 );
and \U$54818 ( \55195 , \55194 , \54451 );
and \U$54819 ( \55196 , \54380 , \54386 );
or \U$54820 ( \55197 , \55195 , \55196 );
xor \U$54821 ( \55198 , \55193 , \55197 );
xor \U$54822 ( \55199 , \54563 , \54568 );
and \U$54823 ( \55200 , \55199 , \54576 );
and \U$54824 ( \55201 , \54563 , \54568 );
or \U$54825 ( \55202 , \55200 , \55201 );
and \U$54826 ( \55203 , \2224 , RIae776a8_81);
and \U$54827 ( \55204 , RIae77450_76, \2222 );
nor \U$54828 ( \55205 , \55203 , \55204 );
and \U$54829 ( \55206 , \55205 , \2061 );
not \U$54830 ( \55207 , \55205 );
and \U$54831 ( \55208 , \55207 , \2060 );
nor \U$54832 ( \55209 , \55206 , \55208 );
xor \U$54833 ( \55210 , \55202 , \55209 );
xor \U$54834 ( \55211 , \54591 , \54599 );
and \U$54835 ( \55212 , \55211 , \54607 );
and \U$54836 ( \55213 , \54591 , \54599 );
or \U$54837 ( \55214 , \55212 , \55213 );
xor \U$54838 ( \55215 , \55210 , \55214 );
xor \U$54839 ( \55216 , \54433 , \54440 );
and \U$54840 ( \55217 , \55216 , \54448 );
and \U$54841 ( \55218 , \54433 , \54440 );
or \U$54842 ( \55219 , \55217 , \55218 );
xor \U$54843 ( \55220 , \54394 , \1734 );
and \U$54844 ( \55221 , \55220 , \54402 );
and \U$54845 ( \55222 , \54394 , \1734 );
or \U$54846 ( \55223 , \55221 , \55222 );
xor \U$54847 ( \55224 , \55219 , \55223 );
xor \U$54848 ( \55225 , \54410 , \54417 );
and \U$54849 ( \55226 , \55225 , \54425 );
and \U$54850 ( \55227 , \54410 , \54417 );
or \U$54851 ( \55228 , \55226 , \55227 );
xor \U$54852 ( \55229 , \55224 , \55228 );
xor \U$54853 ( \55230 , \55215 , \55229 );
xor \U$54854 ( \55231 , \54498 , \54505 );
and \U$54855 ( \55232 , \55231 , \54513 );
and \U$54856 ( \55233 , \54498 , \54505 );
or \U$54857 ( \55234 , \55232 , \55233 );
xor \U$54858 ( \55235 , \54521 , \54528 );
and \U$54859 ( \55236 , \55235 , \54536 );
and \U$54860 ( \55237 , \54521 , \54528 );
or \U$54861 ( \55238 , \55236 , \55237 );
xor \U$54862 ( \55239 , \55234 , \55238 );
xor \U$54863 ( \55240 , \54475 , \54482 );
and \U$54864 ( \55241 , \55240 , \54490 );
and \U$54865 ( \55242 , \54475 , \54482 );
or \U$54866 ( \55243 , \55241 , \55242 );
xor \U$54867 ( \55244 , \55239 , \55243 );
xor \U$54868 ( \55245 , \55230 , \55244 );
and \U$54869 ( \55246 , \12180 , RIae75fb0_32);
and \U$54870 ( \55247 , RIae75ec0_30, \12178 );
nor \U$54871 ( \55248 , \55246 , \55247 );
and \U$54872 ( \55249 , \55248 , \11827 );
not \U$54873 ( \55250 , \55248 );
and \U$54874 ( \55251 , \55250 , \12184 );
nor \U$54875 ( \55252 , \55249 , \55251 );
not \U$54876 ( \55253 , \55252 );
and \U$54877 ( \55254 , \13059 , RIae75ce0_26);
and \U$54878 ( \55255 , RIae75dd0_28, \13057 );
nor \U$54879 ( \55256 , \55254 , \55255 );
and \U$54880 ( \55257 , \55256 , \13063 );
not \U$54881 ( \55258 , \55256 );
and \U$54882 ( \55259 , \55258 , \12718 );
nor \U$54883 ( \55260 , \55257 , \55259 );
not \U$54884 ( \55261 , \55260 );
or \U$54885 ( \55262 , \55253 , \55261 );
or \U$54886 ( \55263 , \55252 , \55260 );
nand \U$54887 ( \55264 , \55262 , \55263 );
not \U$54888 ( \55265 , \55264 );
and \U$54889 ( \55266 , \11470 , RIae75a10_20);
and \U$54890 ( \55267 , RIae75920_18, \11468 );
nor \U$54891 ( \55268 , \55266 , \55267 );
and \U$54892 ( \55269 , \55268 , \11474 );
not \U$54893 ( \55270 , \55268 );
and \U$54894 ( \55271 , \55270 , \10936 );
nor \U$54895 ( \55272 , \55269 , \55271 );
not \U$54896 ( \55273 , \55272 );
and \U$54897 ( \55274 , \55265 , \55273 );
and \U$54898 ( \55275 , \55264 , \55272 );
nor \U$54899 ( \55276 , \55274 , \55275 );
not \U$54900 ( \55277 , \55276 );
xor \U$54901 ( \55278 , \54475 , \54482 );
xor \U$54902 ( \55279 , \55278 , \54490 );
and \U$54903 ( \55280 , \54514 , \55279 );
xor \U$54904 ( \55281 , \54475 , \54482 );
xor \U$54905 ( \55282 , \55281 , \54490 );
and \U$54906 ( \55283 , \54537 , \55282 );
and \U$54907 ( \55284 , \54514 , \54537 );
or \U$54908 ( \55285 , \55280 , \55283 , \55284 );
not \U$54909 ( \55286 , \55285 );
xor \U$54910 ( \55287 , \54394 , \1734 );
xor \U$54911 ( \55288 , \55287 , \54402 );
and \U$54912 ( \55289 , \54426 , \55288 );
xor \U$54913 ( \55290 , \54394 , \1734 );
xor \U$54914 ( \55291 , \55290 , \54402 );
and \U$54915 ( \55292 , \54449 , \55291 );
and \U$54916 ( \55293 , \54426 , \54449 );
or \U$54917 ( \55294 , \55289 , \55292 , \55293 );
not \U$54918 ( \55295 , \55294 );
xor \U$54919 ( \55296 , \55286 , \55295 );
not \U$54920 ( \55297 , \55296 );
or \U$54921 ( \55298 , \55277 , \55297 );
or \U$54922 ( \55299 , \55296 , \55276 );
nand \U$54923 ( \55300 , \55298 , \55299 );
and \U$54924 ( \55301 , \5896 , RIae77f90_100);
and \U$54925 ( \55302 , RIae78080_102, \5894 );
nor \U$54926 ( \55303 , \55301 , \55302 );
and \U$54927 ( \55304 , \55303 , \5589 );
not \U$54928 ( \55305 , \55303 );
and \U$54929 ( \55306 , \55305 , \5590 );
nor \U$54930 ( \55307 , \55304 , \55306 );
not \U$54931 ( \55308 , \55307 );
and \U$54932 ( \55309 , \6172 , RIae78260_106);
and \U$54933 ( \55310 , RIae78620_114, \6170 );
nor \U$54934 ( \55311 , \55309 , \55310 );
and \U$54935 ( \55312 , \55311 , \6176 );
not \U$54936 ( \55313 , \55311 );
and \U$54937 ( \55314 , \55313 , \6175 );
nor \U$54938 ( \55315 , \55312 , \55314 );
not \U$54939 ( \55316 , \55315 );
or \U$54940 ( \55317 , \55308 , \55316 );
or \U$54941 ( \55318 , \55307 , \55315 );
nand \U$54942 ( \55319 , \55317 , \55318 );
not \U$54943 ( \55320 , \55319 );
and \U$54944 ( \55321 , \5399 , RIae78350_108);
and \U$54945 ( \55322 , RIae78170_104, \5397 );
nor \U$54946 ( \55323 , \55321 , \55322 );
and \U$54947 ( \55324 , \55323 , \5403 );
not \U$54948 ( \55325 , \55323 );
and \U$54949 ( \55326 , \55325 , \5016 );
nor \U$54950 ( \55327 , \55324 , \55326 );
not \U$54951 ( \55328 , \55327 );
and \U$54952 ( \55329 , \55320 , \55328 );
and \U$54953 ( \55330 , \55319 , \55327 );
nor \U$54954 ( \55331 , \55329 , \55330 );
not \U$54955 ( \55332 , \55331 );
and \U$54956 ( \55333 , \8371 , RIae77db0_96);
and \U$54957 ( \55334 , RIae77ea0_98, \8369 );
nor \U$54958 ( \55335 , \55333 , \55334 );
and \U$54959 ( \55336 , \55335 , \8020 );
not \U$54960 ( \55337 , \55335 );
and \U$54961 ( \55338 , \55337 , \8019 );
nor \U$54962 ( \55339 , \55336 , \55338 );
and \U$54963 ( \55340 , \6941 , RIae78440_110);
and \U$54964 ( \55341 , RIae784b8_111, \6939 );
nor \U$54965 ( \55342 , \55340 , \55341 );
and \U$54966 ( \55343 , \55342 , \6314 );
not \U$54967 ( \55344 , \55342 );
and \U$54968 ( \55345 , \55344 , \6945 );
nor \U$54969 ( \55346 , \55343 , \55345 );
xor \U$54970 ( \55347 , \55339 , \55346 );
and \U$54971 ( \55348 , \7633 , RIae77cc0_94);
and \U$54972 ( \55349 , RIae77bd0_92, \7631 );
nor \U$54973 ( \55350 , \55348 , \55349 );
and \U$54974 ( \55351 , \55350 , \7206 );
not \U$54975 ( \55352 , \55350 );
and \U$54976 ( \55353 , \55352 , \7205 );
nor \U$54977 ( \55354 , \55351 , \55353 );
xor \U$54978 ( \55355 , \55347 , \55354 );
not \U$54979 ( \55356 , \55355 );
or \U$54980 ( \55357 , \55332 , \55356 );
or \U$54981 ( \55358 , \55331 , \55355 );
nand \U$54982 ( \55359 , \55357 , \55358 );
not \U$54983 ( \55360 , \55359 );
and \U$54984 ( \55361 , \9760 , RIae78800_118);
and \U$54985 ( \55362 , RIae78710_116, \9758 );
nor \U$54986 ( \55363 , \55361 , \55362 );
and \U$54987 ( \55364 , \55363 , \9272 );
not \U$54988 ( \55365 , \55363 );
and \U$54989 ( \55366 , \55365 , \9273 );
nor \U$54990 ( \55367 , \55364 , \55366 );
and \U$54991 ( \55368 , \10548 , RIae75bf0_24);
and \U$54992 ( \55369 , RIae75b00_22, \10546 );
nor \U$54993 ( \55370 , \55368 , \55369 );
and \U$54994 ( \55371 , \55370 , \10118 );
not \U$54995 ( \55372 , \55370 );
and \U$54996 ( \55373 , \55372 , \10421 );
nor \U$54997 ( \55374 , \55371 , \55373 );
xor \U$54998 ( \55375 , \55367 , \55374 );
and \U$54999 ( \55376 , \8966 , RIae789e0_122);
and \U$55000 ( \55377 , RIae788f0_120, \8964 );
nor \U$55001 ( \55378 , \55376 , \55377 );
and \U$55002 ( \55379 , \55378 , \8789 );
not \U$55003 ( \55380 , \55378 );
and \U$55004 ( \55381 , \55380 , \8799 );
nor \U$55005 ( \55382 , \55379 , \55381 );
xor \U$55006 ( \55383 , \55375 , \55382 );
not \U$55007 ( \55384 , \55383 );
and \U$55008 ( \55385 , \55360 , \55384 );
and \U$55009 ( \55386 , \55359 , \55383 );
nor \U$55010 ( \55387 , \55385 , \55386 );
not \U$55011 ( \55388 , \55387 );
and \U$55012 ( \55389 , \15726 , RIae75290_4);
and \U$55013 ( \55390 , RIae751a0_2, RIae7aab0_192);
nor \U$55014 ( \55391 , \55389 , \55390 );
and \U$55015 ( \55392 , \55391 , RIae7aa38_191);
not \U$55016 ( \55393 , \55391 );
and \U$55017 ( \55394 , \55393 , \14959 );
nor \U$55018 ( \55395 , \55392 , \55394 );
not \U$55019 ( \55396 , \55395 );
and \U$55020 ( \55397 , \14964 , RIae75830_16);
and \U$55021 ( \55398 , RIae75740_14, \14962 );
nor \U$55022 ( \55399 , \55397 , \55398 );
and \U$55023 ( \55400 , \55399 , \14463 );
not \U$55024 ( \55401 , \55399 );
and \U$55025 ( \55402 , \55401 , \14462 );
nor \U$55026 ( \55403 , \55400 , \55402 );
not \U$55027 ( \55404 , \55403 );
or \U$55028 ( \55405 , \55396 , \55404 );
or \U$55029 ( \55406 , \55403 , \55395 );
nand \U$55030 ( \55407 , \55405 , \55406 );
not \U$55031 ( \55408 , \55407 );
and \U$55032 ( \55409 , \14059 , RIae75650_12);
and \U$55033 ( \55410 , RIae75560_10, \14057 );
nor \U$55034 ( \55411 , \55409 , \55410 );
and \U$55035 ( \55412 , \55411 , \14063 );
not \U$55036 ( \55413 , \55411 );
and \U$55037 ( \55414 , \55413 , \13502 );
nor \U$55038 ( \55415 , \55412 , \55414 );
not \U$55039 ( \55416 , \55415 );
and \U$55040 ( \55417 , \55408 , \55416 );
and \U$55041 ( \55418 , \55407 , \55415 );
nor \U$55042 ( \55419 , \55417 , \55418 );
and \U$55043 ( \55420 , \1939 , RIae77630_80);
and \U$55044 ( \55421 , RIae77540_78, \1937 );
nor \U$55045 ( \55422 , \55420 , \55421 );
and \U$55046 ( \55423 , \55422 , \1734 );
not \U$55047 ( \55424 , \55422 );
and \U$55048 ( \55425 , \55424 , \1735 );
nor \U$55049 ( \55426 , \55423 , \55425 );
not \U$55050 ( \55427 , \55426 );
and \U$55051 ( \55428 , \4688 , RIae77270_72);
and \U$55052 ( \55429 , RIae77360_74, \4686 );
nor \U$55053 ( \55430 , \55428 , \55429 );
and \U$55054 ( \55431 , \55430 , \4481 );
not \U$55055 ( \55432 , \55430 );
and \U$55056 ( \55433 , \55432 , \4482 );
nor \U$55057 ( \55434 , \55431 , \55433 );
and \U$55058 ( \55435 , \3730 , RIae76dc0_62);
and \U$55059 ( \55436 , RIae76cd0_60, \3728 );
nor \U$55060 ( \55437 , \55435 , \55436 );
and \U$55061 ( \55438 , \55437 , \3732 );
not \U$55062 ( \55439 , \55437 );
and \U$55063 ( \55440 , \55439 , \3422 );
nor \U$55064 ( \55441 , \55438 , \55440 );
xor \U$55065 ( \55442 , \55434 , \55441 );
and \U$55066 ( \55443 , \4247 , RIae77108_69);
and \U$55067 ( \55444 , RIae77090_68, \4245 );
nor \U$55068 ( \55445 , \55443 , \55444 );
and \U$55069 ( \55446 , \55445 , \3989 );
not \U$55070 ( \55447 , \55445 );
and \U$55071 ( \55448 , \55447 , \4251 );
nor \U$55072 ( \55449 , \55446 , \55448 );
xor \U$55073 ( \55450 , \55442 , \55449 );
not \U$55074 ( \55451 , \55450 );
or \U$55075 ( \55452 , \55427 , \55451 );
or \U$55076 ( \55453 , \55450 , \55426 );
nand \U$55077 ( \55454 , \55452 , \55453 );
not \U$55078 ( \55455 , \55454 );
and \U$55079 ( \55456 , \2783 , RIae77810_84);
and \U$55080 ( \55457 , RIae77900_86, \2781 );
nor \U$55081 ( \55458 , \55456 , \55457 );
not \U$55082 ( \55459 , \55458 );
not \U$55083 ( \55460 , \3089 );
and \U$55084 ( \55461 , \55459 , \55460 );
and \U$55085 ( \55462 , \55458 , \3089 );
nor \U$55086 ( \55463 , \55461 , \55462 );
not \U$55087 ( \55464 , \55463 );
not \U$55088 ( \55465 , \2774 );
and \U$55089 ( \55466 , \3214 , RIae76fa0_66);
and \U$55090 ( \55467 , RIae76eb0_64, \3212 );
nor \U$55091 ( \55468 , \55466 , \55467 );
not \U$55092 ( \55469 , \55468 );
or \U$55093 ( \55470 , \55465 , \55469 );
or \U$55094 ( \55471 , \55468 , \2774 );
nand \U$55095 ( \55472 , \55470 , \55471 );
not \U$55096 ( \55473 , \55472 );
or \U$55097 ( \55474 , \55464 , \55473 );
or \U$55098 ( \55475 , \55463 , \55472 );
nand \U$55099 ( \55476 , \55474 , \55475 );
not \U$55100 ( \55477 , \55476 );
and \U$55101 ( \55478 , \2607 , RIae77ae0_90);
and \U$55102 ( \55479 , RIae779f0_88, \2605 );
nor \U$55103 ( \55480 , \55478 , \55479 );
and \U$55104 ( \55481 , \55480 , \2397 );
not \U$55105 ( \55482 , \55480 );
and \U$55106 ( \55483 , \55482 , \2611 );
nor \U$55107 ( \55484 , \55481 , \55483 );
not \U$55108 ( \55485 , \55484 );
and \U$55109 ( \55486 , \55477 , \55485 );
and \U$55110 ( \55487 , \55476 , \55484 );
nor \U$55111 ( \55488 , \55486 , \55487 );
not \U$55112 ( \55489 , \55488 );
and \U$55113 ( \55490 , \55455 , \55489 );
and \U$55114 ( \55491 , \55454 , \55488 );
nor \U$55115 ( \55492 , \55490 , \55491 );
xor \U$55116 ( \55493 , \55419 , \55492 );
not \U$55117 ( \55494 , \55493 );
or \U$55118 ( \55495 , \55388 , \55494 );
or \U$55119 ( \55496 , \55493 , \55387 );
nand \U$55120 ( \55497 , \55495 , \55496 );
xor \U$55121 ( \55498 , \55300 , \55497 );
xor \U$55122 ( \55499 , \55245 , \55498 );
xor \U$55123 ( \55500 , \55198 , \55499 );
not \U$55124 ( \55501 , \55500 );
and \U$55125 ( \55502 , \55184 , \55501 );
and \U$55126 ( \55503 , \55183 , \55500 );
nor \U$55127 ( \55504 , \55502 , \55503 );
not \U$55128 ( \55505 , \55504 );
and \U$55129 ( \55506 , \55146 , \55505 );
and \U$55130 ( \55507 , \55145 , \55504 );
nor \U$55131 ( \55508 , \55506 , \55507 );
or \U$55132 ( \55509 , \55134 , \55508 );
xnor \U$55133 ( \55510 , \55508 , \55134 );
xor \U$55134 ( \55511 , \54960 , \54968 );
xor \U$55135 ( \55512 , \55511 , \54994 );
xor \U$55136 ( \55513 , \54905 , \54923 );
xor \U$55137 ( \55514 , \55513 , \54949 );
and \U$55138 ( \55515 , \55512 , \55514 );
xor \U$55139 ( \55516 , \55023 , \55048 );
xor \U$55140 ( \55517 , \55516 , \55074 );
xor \U$55141 ( \55518 , \54905 , \54923 );
xor \U$55142 ( \55519 , \55518 , \54949 );
and \U$55143 ( \55520 , \55517 , \55519 );
and \U$55144 ( \55521 , \55512 , \55517 );
or \U$55145 ( \55522 , \55515 , \55520 , \55521 );
and \U$55146 ( \55523 , \5399 , RIae76fa0_66);
and \U$55147 ( \55524 , RIae76eb0_64, \5397 );
nor \U$55148 ( \55525 , \55523 , \55524 );
and \U$55149 ( \55526 , \55525 , \5403 );
not \U$55150 ( \55527 , \55525 );
and \U$55151 ( \55528 , \55527 , \5016 );
nor \U$55152 ( \55529 , \55526 , \55528 );
and \U$55153 ( \55530 , \5896 , RIae76dc0_62);
and \U$55154 ( \55531 , RIae76cd0_60, \5894 );
nor \U$55155 ( \55532 , \55530 , \55531 );
and \U$55156 ( \55533 , \55532 , \5589 );
not \U$55157 ( \55534 , \55532 );
and \U$55158 ( \55535 , \55534 , \5590 );
nor \U$55159 ( \55536 , \55533 , \55535 );
or \U$55160 ( \55537 , \55529 , \55536 );
not \U$55161 ( \55538 , \55536 );
not \U$55162 ( \55539 , \55529 );
or \U$55163 ( \55540 , \55538 , \55539 );
and \U$55164 ( \55541 , \6172 , RIae77108_69);
and \U$55165 ( \55542 , RIae77090_68, \6170 );
nor \U$55166 ( \55543 , \55541 , \55542 );
and \U$55167 ( \55544 , \55543 , \6176 );
not \U$55168 ( \55545 , \55543 );
and \U$55169 ( \55546 , \55545 , \6175 );
nor \U$55170 ( \55547 , \55544 , \55546 );
nand \U$55171 ( \55548 , \55540 , \55547 );
nand \U$55172 ( \55549 , \55537 , \55548 );
and \U$55173 ( \55550 , \4688 , RIae77810_84);
and \U$55174 ( \55551 , RIae77900_86, \4686 );
nor \U$55175 ( \55552 , \55550 , \55551 );
and \U$55176 ( \55553 , \55552 , \4481 );
not \U$55177 ( \55554 , \55552 );
and \U$55178 ( \55555 , \55554 , \4482 );
nor \U$55179 ( \55556 , \55553 , \55555 );
and \U$55180 ( \55557 , \3730 , RIae776a8_81);
and \U$55181 ( \55558 , RIae77450_76, \3728 );
nor \U$55182 ( \55559 , \55557 , \55558 );
and \U$55183 ( \55560 , \55559 , \3732 );
not \U$55184 ( \55561 , \55559 );
and \U$55185 ( \55562 , \55561 , \3421 );
nor \U$55186 ( \55563 , \55560 , \55562 );
xor \U$55187 ( \55564 , \55556 , \55563 );
and \U$55188 ( \55565 , \4247 , RIae77ae0_90);
and \U$55189 ( \55566 , RIae779f0_88, \4245 );
nor \U$55190 ( \55567 , \55565 , \55566 );
and \U$55191 ( \55568 , \55567 , \3989 );
not \U$55192 ( \55569 , \55567 );
and \U$55193 ( \55570 , \55569 , \4251 );
nor \U$55194 ( \55571 , \55568 , \55570 );
and \U$55195 ( \55572 , \55564 , \55571 );
and \U$55196 ( \55573 , \55556 , \55563 );
or \U$55197 ( \55574 , \55572 , \55573 );
xor \U$55198 ( \55575 , \55549 , \55574 );
and \U$55199 ( \55576 , \7633 , RIae78350_108);
and \U$55200 ( \55577 , RIae78170_104, \7631 );
nor \U$55201 ( \55578 , \55576 , \55577 );
and \U$55202 ( \55579 , \55578 , \7205 );
not \U$55203 ( \55580 , \55578 );
and \U$55204 ( \55581 , \55580 , \7206 );
nor \U$55205 ( \55582 , \55579 , \55581 );
and \U$55206 ( \55583 , \8371 , RIae77f90_100);
and \U$55207 ( \55584 , RIae78080_102, \8369 );
nor \U$55208 ( \55585 , \55583 , \55584 );
and \U$55209 ( \55586 , \55585 , \8019 );
not \U$55210 ( \55587 , \55585 );
and \U$55211 ( \55588 , \55587 , \8020 );
nor \U$55212 ( \55589 , \55586 , \55588 );
xor \U$55213 ( \55590 , \55582 , \55589 );
and \U$55214 ( \55591 , \6941 , RIae77270_72);
and \U$55215 ( \55592 , RIae77360_74, \6939 );
nor \U$55216 ( \55593 , \55591 , \55592 );
and \U$55217 ( \55594 , \55593 , \6945 );
not \U$55218 ( \55595 , \55593 );
and \U$55219 ( \55596 , \55595 , \6314 );
nor \U$55220 ( \55597 , \55594 , \55596 );
and \U$55221 ( \55598 , \55590 , \55597 );
and \U$55222 ( \55599 , \55582 , \55589 );
nor \U$55223 ( \55600 , \55598 , \55599 );
and \U$55224 ( \55601 , \55575 , \55600 );
and \U$55225 ( \55602 , \55549 , \55574 );
or \U$55226 ( \55603 , \55601 , \55602 );
and \U$55227 ( \55604 , \10548 , RIae77cc0_94);
and \U$55228 ( \55605 , RIae77bd0_92, \10546 );
nor \U$55229 ( \55606 , \55604 , \55605 );
and \U$55230 ( \55607 , \55606 , \10421 );
not \U$55231 ( \55608 , \55606 );
and \U$55232 ( \55609 , \55608 , \10118 );
nor \U$55233 ( \55610 , \55607 , \55609 );
and \U$55234 ( \55611 , \8966 , RIae78260_106);
and \U$55235 ( \55612 , RIae78620_114, \8964 );
nor \U$55236 ( \55613 , \55611 , \55612 );
and \U$55237 ( \55614 , \55613 , \8799 );
not \U$55238 ( \55615 , \55613 );
and \U$55239 ( \55616 , \55615 , \8789 );
nor \U$55240 ( \55617 , \55614 , \55616 );
xor \U$55241 ( \55618 , \55610 , \55617 );
and \U$55242 ( \55619 , \9760 , RIae78440_110);
and \U$55243 ( \55620 , RIae784b8_111, \9758 );
nor \U$55244 ( \55621 , \55619 , \55620 );
and \U$55245 ( \55622 , \55621 , \9273 );
not \U$55246 ( \55623 , \55621 );
and \U$55247 ( \55624 , \55623 , \9272 );
nor \U$55248 ( \55625 , \55622 , \55624 );
and \U$55249 ( \55626 , \55618 , \55625 );
and \U$55250 ( \55627 , \55610 , \55617 );
or \U$55251 ( \55628 , \55626 , \55627 );
and \U$55252 ( \55629 , \14059 , RIae75bf0_24);
and \U$55253 ( \55630 , RIae75b00_22, \14057 );
nor \U$55254 ( \55631 , \55629 , \55630 );
and \U$55255 ( \55632 , \55631 , \14063 );
not \U$55256 ( \55633 , \55631 );
and \U$55257 ( \55634 , \55633 , \13502 );
nor \U$55258 ( \55635 , \55632 , \55634 );
and \U$55259 ( \55636 , \15726 , RIae75fb0_32);
and \U$55260 ( \55637 , RIae75ec0_30, RIae7aab0_192);
nor \U$55261 ( \55638 , \55636 , \55637 );
and \U$55262 ( \55639 , \55638 , RIae7aa38_191);
not \U$55263 ( \55640 , \55638 );
and \U$55264 ( \55641 , \55640 , \14959 );
nor \U$55265 ( \55642 , \55639 , \55641 );
or \U$55266 ( \55643 , \55635 , \55642 );
not \U$55267 ( \55644 , \55642 );
not \U$55268 ( \55645 , \55635 );
or \U$55269 ( \55646 , \55644 , \55645 );
and \U$55270 ( \55647 , \14964 , RIae75a10_20);
and \U$55271 ( \55648 , RIae75920_18, \14962 );
nor \U$55272 ( \55649 , \55647 , \55648 );
and \U$55273 ( \55650 , \55649 , \14463 );
not \U$55274 ( \55651 , \55649 );
and \U$55275 ( \55652 , \55651 , \14462 );
nor \U$55276 ( \55653 , \55650 , \55652 );
nand \U$55277 ( \55654 , \55646 , \55653 );
nand \U$55278 ( \55655 , \55643 , \55654 );
xor \U$55279 ( \55656 , \55628 , \55655 );
and \U$55280 ( \55657 , \11470 , RIae77db0_96);
and \U$55281 ( \55658 , RIae77ea0_98, \11468 );
nor \U$55282 ( \55659 , \55657 , \55658 );
and \U$55283 ( \55660 , \55659 , \11474 );
not \U$55284 ( \55661 , \55659 );
and \U$55285 ( \55662 , \55661 , \10936 );
nor \U$55286 ( \55663 , \55660 , \55662 );
and \U$55287 ( \55664 , \12180 , RIae789e0_122);
and \U$55288 ( \55665 , RIae788f0_120, \12178 );
nor \U$55289 ( \55666 , \55664 , \55665 );
and \U$55290 ( \55667 , \55666 , \11827 );
not \U$55291 ( \55668 , \55666 );
and \U$55292 ( \55669 , \55668 , \12184 );
nor \U$55293 ( \55670 , \55667 , \55669 );
or \U$55294 ( \55671 , \55663 , \55670 );
not \U$55295 ( \55672 , \55670 );
not \U$55296 ( \55673 , \55663 );
or \U$55297 ( \55674 , \55672 , \55673 );
and \U$55298 ( \55675 , \13059 , RIae78800_118);
and \U$55299 ( \55676 , RIae78710_116, \13057 );
nor \U$55300 ( \55677 , \55675 , \55676 );
and \U$55301 ( \55678 , \55677 , \13063 );
not \U$55302 ( \55679 , \55677 );
and \U$55303 ( \55680 , \55679 , \12718 );
nor \U$55304 ( \55681 , \55678 , \55680 );
nand \U$55305 ( \55682 , \55674 , \55681 );
nand \U$55306 ( \55683 , \55671 , \55682 );
and \U$55307 ( \55684 , \55656 , \55683 );
and \U$55308 ( \55685 , \55628 , \55655 );
or \U$55309 ( \55686 , \55684 , \55685 );
xor \U$55310 ( \55687 , \55603 , \55686 );
xor \U$55311 ( \55688 , \54976 , \54982 );
xor \U$55312 ( \55689 , \55688 , \54991 );
xor \U$55313 ( \55690 , \55005 , \55012 );
xor \U$55314 ( \55691 , \55690 , \55020 );
and \U$55315 ( \55692 , \55689 , \55691 );
xor \U$55316 ( \55693 , \55030 , \55037 );
xor \U$55317 ( \55694 , \55693 , \55045 );
xor \U$55318 ( \55695 , \55005 , \55012 );
xor \U$55319 ( \55696 , \55695 , \55020 );
and \U$55320 ( \55697 , \55694 , \55696 );
and \U$55321 ( \55698 , \55689 , \55694 );
or \U$55322 ( \55699 , \55692 , \55697 , \55698 );
and \U$55323 ( \55700 , \55687 , \55699 );
and \U$55324 ( \55701 , \55603 , \55686 );
or \U$55325 ( \55702 , \55700 , \55701 );
xor \U$55326 ( \55703 , \55522 , \55702 );
xor \U$55327 ( \55704 , \55056 , \55063 );
xor \U$55328 ( \55705 , \55704 , \55071 );
xor \U$55329 ( \55706 , \54931 , \54938 );
xor \U$55330 ( \55707 , \55706 , \54946 );
and \U$55331 ( \55708 , \55705 , \55707 );
xor \U$55332 ( \55709 , \54887 , \54894 );
xor \U$55333 ( \55710 , \55709 , \54902 );
xor \U$55334 ( \55711 , \54931 , \54938 );
xor \U$55335 ( \55712 , \55711 , \54946 );
and \U$55336 ( \55713 , \55710 , \55712 );
and \U$55337 ( \55714 , \55705 , \55710 );
or \U$55338 ( \55715 , \55708 , \55713 , \55714 );
xor \U$55339 ( \55716 , \54854 , \54856 );
xor \U$55340 ( \55717 , \55716 , \54859 );
and \U$55341 ( \55718 , \55715 , \55717 );
xor \U$55342 ( \55719 , \54658 , \54665 );
xor \U$55343 ( \55720 , \55719 , \54673 );
xor \U$55344 ( \55721 , \54867 , \54872 );
xor \U$55345 ( \55722 , \55720 , \55721 );
xor \U$55346 ( \55723 , \54854 , \54856 );
xor \U$55347 ( \55724 , \55723 , \54859 );
and \U$55348 ( \55725 , \55722 , \55724 );
and \U$55349 ( \55726 , \55715 , \55722 );
or \U$55350 ( \55727 , \55718 , \55725 , \55726 );
and \U$55351 ( \55728 , \55703 , \55727 );
and \U$55352 ( \55729 , \55522 , \55702 );
or \U$55353 ( \55730 , \55728 , \55729 );
xor \U$55354 ( \55731 , \54730 , \54755 );
xor \U$55355 ( \55732 , \55731 , \54781 );
xor \U$55356 ( \55733 , \54651 , \54676 );
xor \U$55357 ( \55734 , \55733 , \54702 );
xor \U$55358 ( \55735 , \55732 , \55734 );
xor \U$55359 ( \55736 , \54787 , \54792 );
xor \U$55360 ( \55737 , \55736 , \54795 );
xor \U$55361 ( \55738 , \55083 , \55090 );
xor \U$55362 ( \55739 , \55737 , \55738 );
and \U$55363 ( \55740 , \55735 , \55739 );
and \U$55364 ( \55741 , \55732 , \55734 );
or \U$55365 ( \55742 , \55740 , \55741 );
xor \U$55366 ( \55743 , \55730 , \55742 );
xor \U$55367 ( \55744 , \54616 , \54618 );
xor \U$55368 ( \55745 , \55744 , \54623 );
xor \U$55369 ( \55746 , \55103 , \55108 );
xor \U$55370 ( \55747 , \55745 , \55746 );
xor \U$55371 ( \55748 , \55743 , \55747 );
not \U$55372 ( \55749 , \55748 );
xor \U$55373 ( \55750 , \54952 , \54997 );
xor \U$55374 ( \55751 , \55750 , \55077 );
xor \U$55375 ( \55752 , \55732 , \55734 );
xor \U$55376 ( \55753 , \55752 , \55739 );
and \U$55377 ( \55754 , \55751 , \55753 );
xor \U$55378 ( \55755 , \55522 , \55702 );
xor \U$55379 ( \55756 , \55755 , \55727 );
xor \U$55380 ( \55757 , \55732 , \55734 );
xor \U$55381 ( \55758 , \55757 , \55739 );
and \U$55382 ( \55759 , \55756 , \55758 );
and \U$55383 ( \55760 , \55751 , \55756 );
or \U$55384 ( \55761 , \55754 , \55759 , \55760 );
xor \U$55385 ( \55762 , \54880 , \55080 );
xor \U$55386 ( \55763 , \55762 , \55095 );
xor \U$55387 ( \55764 , \55761 , \55763 );
xor \U$55388 ( \55765 , \55582 , \55589 );
xor \U$55389 ( \55766 , \55765 , \55597 );
not \U$55390 ( \55767 , \55670 );
not \U$55391 ( \55768 , \55681 );
or \U$55392 ( \55769 , \55767 , \55768 );
or \U$55393 ( \55770 , \55670 , \55681 );
nand \U$55394 ( \55771 , \55769 , \55770 );
not \U$55395 ( \55772 , \55771 );
not \U$55396 ( \55773 , \55663 );
and \U$55397 ( \55774 , \55772 , \55773 );
and \U$55398 ( \55775 , \55771 , \55663 );
nor \U$55399 ( \55776 , \55774 , \55775 );
or \U$55400 ( \55777 , \55766 , \55776 );
not \U$55401 ( \55778 , \55776 );
not \U$55402 ( \55779 , \55766 );
or \U$55403 ( \55780 , \55778 , \55779 );
xor \U$55404 ( \55781 , \55610 , \55617 );
xor \U$55405 ( \55782 , \55781 , \55625 );
nand \U$55406 ( \55783 , \55780 , \55782 );
nand \U$55407 ( \55784 , \55777 , \55783 );
xor \U$55408 ( \55785 , \54912 , \2789 );
xor \U$55409 ( \55786 , \55785 , \54920 );
xor \U$55410 ( \55787 , \55784 , \55786 );
xor \U$55411 ( \55788 , \54931 , \54938 );
xor \U$55412 ( \55789 , \55788 , \54946 );
xor \U$55413 ( \55790 , \55705 , \55710 );
xor \U$55414 ( \55791 , \55789 , \55790 );
and \U$55415 ( \55792 , \55787 , \55791 );
and \U$55416 ( \55793 , \55784 , \55786 );
or \U$55417 ( \55794 , \55792 , \55793 );
and \U$55418 ( \55795 , \4688 , RIae779f0_88);
and \U$55419 ( \55796 , RIae77810_84, \4686 );
nor \U$55420 ( \55797 , \55795 , \55796 );
and \U$55421 ( \55798 , \55797 , \4481 );
not \U$55422 ( \55799 , \55797 );
and \U$55423 ( \55800 , \55799 , \4482 );
nor \U$55424 ( \55801 , \55798 , \55800 );
and \U$55425 ( \55802 , \5399 , RIae77900_86);
and \U$55426 ( \55803 , RIae76fa0_66, \5397 );
nor \U$55427 ( \55804 , \55802 , \55803 );
and \U$55428 ( \55805 , \55804 , \5016 );
not \U$55429 ( \55806 , \55804 );
and \U$55430 ( \55807 , \55806 , \5403 );
nor \U$55431 ( \55808 , \55805 , \55807 );
xor \U$55432 ( \55809 , \55801 , \55808 );
and \U$55433 ( \55810 , \4247 , RIae77450_76);
and \U$55434 ( \55811 , RIae77ae0_90, \4245 );
nor \U$55435 ( \55812 , \55810 , \55811 );
and \U$55436 ( \55813 , \55812 , \3989 );
not \U$55437 ( \55814 , \55812 );
and \U$55438 ( \55815 , \55814 , \4251 );
nor \U$55439 ( \55816 , \55813 , \55815 );
and \U$55440 ( \55817 , \55809 , \55816 );
and \U$55441 ( \55818 , \55801 , \55808 );
nor \U$55442 ( \55819 , \55817 , \55818 );
and \U$55443 ( \55820 , \8371 , RIae78170_104);
and \U$55444 ( \55821 , RIae77f90_100, \8369 );
nor \U$55445 ( \55822 , \55820 , \55821 );
and \U$55446 ( \55823 , \55822 , \8020 );
not \U$55447 ( \55824 , \55822 );
and \U$55448 ( \55825 , \55824 , \8019 );
nor \U$55449 ( \55826 , \55823 , \55825 );
and \U$55450 ( \55827 , \8966 , RIae78080_102);
and \U$55451 ( \55828 , RIae78260_106, \8964 );
nor \U$55452 ( \55829 , \55827 , \55828 );
and \U$55453 ( \55830 , \55829 , \8799 );
not \U$55454 ( \55831 , \55829 );
and \U$55455 ( \55832 , \55831 , \8789 );
nor \U$55456 ( \55833 , \55830 , \55832 );
xor \U$55457 ( \55834 , \55826 , \55833 );
and \U$55458 ( \55835 , \7633 , RIae77360_74);
and \U$55459 ( \55836 , RIae78350_108, \7631 );
nor \U$55460 ( \55837 , \55835 , \55836 );
and \U$55461 ( \55838 , \55837 , \7206 );
not \U$55462 ( \55839 , \55837 );
and \U$55463 ( \55840 , \55839 , \7205 );
nor \U$55464 ( \55841 , \55838 , \55840 );
and \U$55465 ( \55842 , \55834 , \55841 );
and \U$55466 ( \55843 , \55826 , \55833 );
nor \U$55467 ( \55844 , \55842 , \55843 );
xor \U$55468 ( \55845 , \55819 , \55844 );
and \U$55469 ( \55846 , \6172 , RIae76cd0_60);
and \U$55470 ( \55847 , RIae77108_69, \6170 );
nor \U$55471 ( \55848 , \55846 , \55847 );
and \U$55472 ( \55849 , \55848 , \6176 );
not \U$55473 ( \55850 , \55848 );
and \U$55474 ( \55851 , \55850 , \6175 );
nor \U$55475 ( \55852 , \55849 , \55851 );
and \U$55476 ( \55853 , \6941 , RIae77090_68);
and \U$55477 ( \55854 , RIae77270_72, \6939 );
nor \U$55478 ( \55855 , \55853 , \55854 );
and \U$55479 ( \55856 , \55855 , \6314 );
not \U$55480 ( \55857 , \55855 );
and \U$55481 ( \55858 , \55857 , \6945 );
nor \U$55482 ( \55859 , \55856 , \55858 );
xor \U$55483 ( \55860 , \55852 , \55859 );
and \U$55484 ( \55861 , \5896 , RIae76eb0_64);
and \U$55485 ( \55862 , RIae76dc0_62, \5894 );
nor \U$55486 ( \55863 , \55861 , \55862 );
and \U$55487 ( \55864 , \55863 , \5590 );
not \U$55488 ( \55865 , \55863 );
and \U$55489 ( \55866 , \55865 , \5589 );
nor \U$55490 ( \55867 , \55864 , \55866 );
and \U$55491 ( \55868 , \55860 , \55867 );
and \U$55492 ( \55869 , \55852 , \55859 );
nor \U$55493 ( \55870 , \55868 , \55869 );
and \U$55494 ( \55871 , \55845 , \55870 );
and \U$55495 ( \55872 , \55819 , \55844 );
nor \U$55496 ( \55873 , \55871 , \55872 );
and \U$55497 ( \55874 , \15726 , RIae75920_18);
and \U$55498 ( \55875 , RIae75fb0_32, RIae7aab0_192);
nor \U$55499 ( \55876 , \55874 , \55875 );
and \U$55500 ( \55877 , \55876 , \14959 );
not \U$55501 ( \55878 , \55876 );
and \U$55502 ( \55879 , \55878 , RIae7aa38_191);
nor \U$55503 ( \55880 , \55877 , \55879 );
xor \U$55504 ( \55881 , \55880 , \2774 );
and \U$55505 ( \55882 , \14964 , RIae75b00_22);
and \U$55506 ( \55883 , RIae75a10_20, \14962 );
nor \U$55507 ( \55884 , \55882 , \55883 );
and \U$55508 ( \55885 , \55884 , \14463 );
not \U$55509 ( \55886 , \55884 );
and \U$55510 ( \55887 , \55886 , \14462 );
nor \U$55511 ( \55888 , \55885 , \55887 );
and \U$55512 ( \55889 , \55881 , \55888 );
and \U$55513 ( \55890 , \55880 , \2774 );
or \U$55514 ( \55891 , \55889 , \55890 );
not \U$55515 ( \55892 , \55891 );
and \U$55516 ( \55893 , \9760 , RIae78620_114);
and \U$55517 ( \55894 , RIae78440_110, \9758 );
nor \U$55518 ( \55895 , \55893 , \55894 );
and \U$55519 ( \55896 , \55895 , \9273 );
not \U$55520 ( \55897 , \55895 );
and \U$55521 ( \55898 , \55897 , \9272 );
nor \U$55522 ( \55899 , \55896 , \55898 );
and \U$55523 ( \55900 , \10548 , RIae784b8_111);
and \U$55524 ( \55901 , RIae77cc0_94, \10546 );
nor \U$55525 ( \55902 , \55900 , \55901 );
and \U$55526 ( \55903 , \55902 , \10421 );
not \U$55527 ( \55904 , \55902 );
and \U$55528 ( \55905 , \55904 , \10118 );
nor \U$55529 ( \55906 , \55903 , \55905 );
xor \U$55530 ( \55907 , \55899 , \55906 );
and \U$55531 ( \55908 , \11470 , RIae77bd0_92);
and \U$55532 ( \55909 , RIae77db0_96, \11468 );
nor \U$55533 ( \55910 , \55908 , \55909 );
and \U$55534 ( \55911 , \55910 , \10936 );
not \U$55535 ( \55912 , \55910 );
and \U$55536 ( \55913 , \55912 , \11474 );
nor \U$55537 ( \55914 , \55911 , \55913 );
and \U$55538 ( \55915 , \55907 , \55914 );
and \U$55539 ( \55916 , \55899 , \55906 );
or \U$55540 ( \55917 , \55915 , \55916 );
not \U$55541 ( \55918 , \55917 );
or \U$55542 ( \55919 , \55892 , \55918 );
or \U$55543 ( \55920 , \55917 , \55891 );
and \U$55544 ( \55921 , \12180 , RIae77ea0_98);
and \U$55545 ( \55922 , RIae789e0_122, \12178 );
nor \U$55546 ( \55923 , \55921 , \55922 );
and \U$55547 ( \55924 , \55923 , \11827 );
not \U$55548 ( \55925 , \55923 );
and \U$55549 ( \55926 , \55925 , \12184 );
nor \U$55550 ( \55927 , \55924 , \55926 );
and \U$55551 ( \55928 , \13059 , RIae788f0_120);
and \U$55552 ( \55929 , RIae78800_118, \13057 );
nor \U$55553 ( \55930 , \55928 , \55929 );
and \U$55554 ( \55931 , \55930 , \12718 );
not \U$55555 ( \55932 , \55930 );
and \U$55556 ( \55933 , \55932 , \13063 );
nor \U$55557 ( \55934 , \55931 , \55933 );
or \U$55558 ( \55935 , \55927 , \55934 );
not \U$55559 ( \55936 , \55934 );
not \U$55560 ( \55937 , \55927 );
or \U$55561 ( \55938 , \55936 , \55937 );
and \U$55562 ( \55939 , \14059 , RIae78710_116);
and \U$55563 ( \55940 , RIae75bf0_24, \14057 );
nor \U$55564 ( \55941 , \55939 , \55940 );
and \U$55565 ( \55942 , \55941 , \13502 );
not \U$55566 ( \55943 , \55941 );
and \U$55567 ( \55944 , \55943 , \14063 );
nor \U$55568 ( \55945 , \55942 , \55944 );
nand \U$55569 ( \55946 , \55938 , \55945 );
nand \U$55570 ( \55947 , \55935 , \55946 );
nand \U$55571 ( \55948 , \55920 , \55947 );
nand \U$55572 ( \55949 , \55919 , \55948 );
xor \U$55573 ( \55950 , \55873 , \55949 );
not \U$55574 ( \55951 , \55536 );
not \U$55575 ( \55952 , \55547 );
or \U$55576 ( \55953 , \55951 , \55952 );
or \U$55577 ( \55954 , \55536 , \55547 );
nand \U$55578 ( \55955 , \55953 , \55954 );
not \U$55579 ( \55956 , \55955 );
not \U$55580 ( \55957 , \55529 );
and \U$55581 ( \55958 , \55956 , \55957 );
and \U$55582 ( \55959 , \55955 , \55529 );
nor \U$55583 ( \55960 , \55958 , \55959 );
and \U$55584 ( \55961 , \3214 , RIae77630_80);
and \U$55585 ( \55962 , RIae77540_78, \3212 );
nor \U$55586 ( \55963 , \55961 , \55962 );
not \U$55587 ( \55964 , \55963 );
not \U$55588 ( \55965 , \2774 );
and \U$55589 ( \55966 , \55964 , \55965 );
and \U$55590 ( \55967 , \55963 , \3218 );
nor \U$55591 ( \55968 , \55966 , \55967 );
or \U$55592 ( \55969 , \55960 , \55968 );
not \U$55593 ( \55970 , \55968 );
not \U$55594 ( \55971 , \55960 );
or \U$55595 ( \55972 , \55970 , \55971 );
xor \U$55596 ( \55973 , \55556 , \55563 );
xor \U$55597 ( \55974 , \55973 , \55571 );
nand \U$55598 ( \55975 , \55972 , \55974 );
nand \U$55599 ( \55976 , \55969 , \55975 );
and \U$55600 ( \55977 , \55950 , \55976 );
and \U$55601 ( \55978 , \55873 , \55949 );
or \U$55602 ( \55979 , \55977 , \55978 );
xor \U$55603 ( \55980 , \55794 , \55979 );
xor \U$55604 ( \55981 , \55628 , \55655 );
xor \U$55605 ( \55982 , \55981 , \55683 );
xor \U$55606 ( \55983 , \55549 , \55574 );
xor \U$55607 ( \55984 , \55983 , \55600 );
and \U$55608 ( \55985 , \55982 , \55984 );
xor \U$55609 ( \55986 , \55005 , \55012 );
xor \U$55610 ( \55987 , \55986 , \55020 );
xor \U$55611 ( \55988 , \55689 , \55694 );
xor \U$55612 ( \55989 , \55987 , \55988 );
xor \U$55613 ( \55990 , \55549 , \55574 );
xor \U$55614 ( \55991 , \55990 , \55600 );
and \U$55615 ( \55992 , \55989 , \55991 );
and \U$55616 ( \55993 , \55982 , \55989 );
or \U$55617 ( \55994 , \55985 , \55992 , \55993 );
and \U$55618 ( \55995 , \55980 , \55994 );
and \U$55619 ( \55996 , \55794 , \55979 );
or \U$55620 ( \55997 , \55995 , \55996 );
xor \U$55621 ( \55998 , \54862 , \54864 );
xor \U$55622 ( \55999 , \55998 , \54877 );
xor \U$55623 ( \56000 , \55997 , \55999 );
xor \U$55624 ( \56001 , \54905 , \54923 );
xor \U$55625 ( \56002 , \56001 , \54949 );
xor \U$55626 ( \56003 , \55512 , \55517 );
xor \U$55627 ( \56004 , \56002 , \56003 );
xor \U$55628 ( \56005 , \55603 , \55686 );
xor \U$55629 ( \56006 , \56005 , \55699 );
and \U$55630 ( \56007 , \56004 , \56006 );
xor \U$55631 ( \56008 , \54854 , \54856 );
xor \U$55632 ( \56009 , \56008 , \54859 );
xor \U$55633 ( \56010 , \55715 , \55722 );
xor \U$55634 ( \56011 , \56009 , \56010 );
xor \U$55635 ( \56012 , \55603 , \55686 );
xor \U$55636 ( \56013 , \56012 , \55699 );
and \U$55637 ( \56014 , \56011 , \56013 );
and \U$55638 ( \56015 , \56004 , \56011 );
or \U$55639 ( \56016 , \56007 , \56014 , \56015 );
and \U$55640 ( \56017 , \56000 , \56016 );
and \U$55641 ( \56018 , \55997 , \55999 );
or \U$55642 ( \56019 , \56017 , \56018 );
xor \U$55643 ( \56020 , \55764 , \56019 );
not \U$55644 ( \56021 , \56020 );
or \U$55645 ( \56022 , \55749 , \56021 );
or \U$55646 ( \56023 , \56020 , \55748 );
xor \U$55647 ( \56024 , \55997 , \55999 );
xor \U$55648 ( \56025 , \56024 , \56016 );
not \U$55649 ( \56026 , \56025 );
xor \U$55650 ( \56027 , \55732 , \55734 );
xor \U$55651 ( \56028 , \56027 , \55739 );
xor \U$55652 ( \56029 , \55751 , \55756 );
xor \U$55653 ( \56030 , \56028 , \56029 );
not \U$55654 ( \56031 , \56030 );
or \U$55655 ( \56032 , \56026 , \56031 );
or \U$55656 ( \56033 , \56030 , \56025 );
xor \U$55657 ( \56034 , \55873 , \55949 );
xor \U$55658 ( \56035 , \56034 , \55976 );
xor \U$55659 ( \56036 , \55784 , \55786 );
xor \U$55660 ( \56037 , \56036 , \55791 );
and \U$55661 ( \56038 , \56035 , \56037 );
xor \U$55662 ( \56039 , \55549 , \55574 );
xor \U$55663 ( \56040 , \56039 , \55600 );
xor \U$55664 ( \56041 , \55982 , \55989 );
xor \U$55665 ( \56042 , \56040 , \56041 );
xor \U$55666 ( \56043 , \55784 , \55786 );
xor \U$55667 ( \56044 , \56043 , \55791 );
and \U$55668 ( \56045 , \56042 , \56044 );
and \U$55669 ( \56046 , \56035 , \56042 );
or \U$55670 ( \56047 , \56038 , \56045 , \56046 );
not \U$55671 ( \56048 , \55934 );
not \U$55672 ( \56049 , \55945 );
or \U$55673 ( \56050 , \56048 , \56049 );
or \U$55674 ( \56051 , \55934 , \55945 );
nand \U$55675 ( \56052 , \56050 , \56051 );
not \U$55676 ( \56053 , \56052 );
not \U$55677 ( \56054 , \55927 );
and \U$55678 ( \56055 , \56053 , \56054 );
and \U$55679 ( \56056 , \56052 , \55927 );
nor \U$55680 ( \56057 , \56055 , \56056 );
not \U$55681 ( \56058 , \56057 );
xor \U$55682 ( \56059 , \55880 , \2774 );
xor \U$55683 ( \56060 , \56059 , \55888 );
nand \U$55684 ( \56061 , \56058 , \56060 );
not \U$55685 ( \56062 , \55642 );
not \U$55686 ( \56063 , \55653 );
or \U$55687 ( \56064 , \56062 , \56063 );
or \U$55688 ( \56065 , \55653 , \55642 );
nand \U$55689 ( \56066 , \56064 , \56065 );
not \U$55690 ( \56067 , \56066 );
not \U$55691 ( \56068 , \55635 );
and \U$55692 ( \56069 , \56067 , \56068 );
and \U$55693 ( \56070 , \56066 , \55635 );
nor \U$55694 ( \56071 , \56069 , \56070 );
xor \U$55695 ( \56072 , \56061 , \56071 );
xor \U$55696 ( \56073 , \55826 , \55833 );
xor \U$55697 ( \56074 , \56073 , \55841 );
xor \U$55698 ( \56075 , \55899 , \55906 );
xor \U$55699 ( \56076 , \56075 , \55914 );
xor \U$55700 ( \56077 , \56074 , \56076 );
xor \U$55701 ( \56078 , \55852 , \55859 );
xor \U$55702 ( \56079 , \56078 , \55867 );
and \U$55703 ( \56080 , \56077 , \56079 );
and \U$55704 ( \56081 , \56074 , \56076 );
nor \U$55705 ( \56082 , \56080 , \56081 );
and \U$55706 ( \56083 , \56072 , \56082 );
and \U$55707 ( \56084 , \56061 , \56071 );
or \U$55708 ( \56085 , \56083 , \56084 );
and \U$55709 ( \56086 , \13059 , RIae789e0_122);
and \U$55710 ( \56087 , RIae788f0_120, \13057 );
nor \U$55711 ( \56088 , \56086 , \56087 );
and \U$55712 ( \56089 , \56088 , \13063 );
not \U$55713 ( \56090 , \56088 );
and \U$55714 ( \56091 , \56090 , \12718 );
nor \U$55715 ( \56092 , \56089 , \56091 );
and \U$55716 ( \56093 , \11470 , RIae77cc0_94);
and \U$55717 ( \56094 , RIae77bd0_92, \11468 );
nor \U$55718 ( \56095 , \56093 , \56094 );
and \U$55719 ( \56096 , \56095 , \10936 );
not \U$55720 ( \56097 , \56095 );
and \U$55721 ( \56098 , \56097 , \11474 );
nor \U$55722 ( \56099 , \56096 , \56098 );
xor \U$55723 ( \56100 , \56092 , \56099 );
and \U$55724 ( \56101 , \12180 , RIae77db0_96);
and \U$55725 ( \56102 , RIae77ea0_98, \12178 );
nor \U$55726 ( \56103 , \56101 , \56102 );
and \U$55727 ( \56104 , \56103 , \12184 );
not \U$55728 ( \56105 , \56103 );
and \U$55729 ( \56106 , \56105 , \11827 );
nor \U$55730 ( \56107 , \56104 , \56106 );
and \U$55731 ( \56108 , \56100 , \56107 );
and \U$55732 ( \56109 , \56092 , \56099 );
or \U$55733 ( \56110 , \56108 , \56109 );
and \U$55734 ( \56111 , \14059 , RIae78800_118);
and \U$55735 ( \56112 , RIae78710_116, \14057 );
nor \U$55736 ( \56113 , \56111 , \56112 );
and \U$55737 ( \56114 , \56113 , \14063 );
not \U$55738 ( \56115 , \56113 );
and \U$55739 ( \56116 , \56115 , \13502 );
nor \U$55740 ( \56117 , \56114 , \56116 );
and \U$55741 ( \56118 , \15726 , RIae75a10_20);
and \U$55742 ( \56119 , RIae75920_18, RIae7aab0_192);
nor \U$55743 ( \56120 , \56118 , \56119 );
and \U$55744 ( \56121 , \56120 , RIae7aa38_191);
not \U$55745 ( \56122 , \56120 );
and \U$55746 ( \56123 , \56122 , \14959 );
nor \U$55747 ( \56124 , \56121 , \56123 );
or \U$55748 ( \56125 , \56117 , \56124 );
not \U$55749 ( \56126 , \56124 );
not \U$55750 ( \56127 , \56117 );
or \U$55751 ( \56128 , \56126 , \56127 );
and \U$55752 ( \56129 , \14964 , RIae75bf0_24);
and \U$55753 ( \56130 , RIae75b00_22, \14962 );
nor \U$55754 ( \56131 , \56129 , \56130 );
and \U$55755 ( \56132 , \56131 , \14463 );
not \U$55756 ( \56133 , \56131 );
and \U$55757 ( \56134 , \56133 , \14462 );
nor \U$55758 ( \56135 , \56132 , \56134 );
nand \U$55759 ( \56136 , \56128 , \56135 );
nand \U$55760 ( \56137 , \56125 , \56136 );
xor \U$55761 ( \56138 , \56110 , \56137 );
and \U$55762 ( \56139 , \8966 , RIae77f90_100);
and \U$55763 ( \56140 , RIae78080_102, \8964 );
nor \U$55764 ( \56141 , \56139 , \56140 );
and \U$55765 ( \56142 , \56141 , \8789 );
not \U$55766 ( \56143 , \56141 );
and \U$55767 ( \56144 , \56143 , \8799 );
nor \U$55768 ( \56145 , \56142 , \56144 );
and \U$55769 ( \56146 , \9760 , RIae78260_106);
and \U$55770 ( \56147 , RIae78620_114, \9758 );
nor \U$55771 ( \56148 , \56146 , \56147 );
and \U$55772 ( \56149 , \56148 , \9272 );
not \U$55773 ( \56150 , \56148 );
and \U$55774 ( \56151 , \56150 , \9273 );
nor \U$55775 ( \56152 , \56149 , \56151 );
or \U$55776 ( \56153 , \56145 , \56152 );
not \U$55777 ( \56154 , \56152 );
not \U$55778 ( \56155 , \56145 );
or \U$55779 ( \56156 , \56154 , \56155 );
and \U$55780 ( \56157 , \10548 , RIae78440_110);
and \U$55781 ( \56158 , RIae784b8_111, \10546 );
nor \U$55782 ( \56159 , \56157 , \56158 );
and \U$55783 ( \56160 , \56159 , \10421 );
not \U$55784 ( \56161 , \56159 );
and \U$55785 ( \56162 , \56161 , \10118 );
nor \U$55786 ( \56163 , \56160 , \56162 );
nand \U$55787 ( \56164 , \56156 , \56163 );
nand \U$55788 ( \56165 , \56153 , \56164 );
and \U$55789 ( \56166 , \56138 , \56165 );
and \U$55790 ( \56167 , \56110 , \56137 );
nor \U$55791 ( \56168 , \56166 , \56167 );
nand \U$55792 ( \56169 , RIae77630_80, \3212 );
not \U$55793 ( \56170 , \56169 );
not \U$55794 ( \56171 , \2774 );
or \U$55795 ( \56172 , \56170 , \56171 );
or \U$55796 ( \56173 , \2774 , \56169 );
nand \U$55797 ( \56174 , \56172 , \56173 );
and \U$55798 ( \56175 , \3730 , RIae77540_78);
and \U$55799 ( \56176 , RIae776a8_81, \3728 );
nor \U$55800 ( \56177 , \56175 , \56176 );
and \U$55801 ( \56178 , \56177 , \3732 );
not \U$55802 ( \56179 , \56177 );
and \U$55803 ( \56180 , \56179 , \3422 );
nor \U$55804 ( \56181 , \56178 , \56180 );
xor \U$55805 ( \56182 , \56174 , \56181 );
xor \U$55806 ( \56183 , \55801 , \55808 );
xor \U$55807 ( \56184 , \56183 , \55816 );
and \U$55808 ( \56185 , \56182 , \56184 );
and \U$55809 ( \56186 , \56174 , \56181 );
nor \U$55810 ( \56187 , \56185 , \56186 );
xor \U$55811 ( \56188 , \56168 , \56187 );
and \U$55812 ( \56189 , \4247 , RIae776a8_81);
and \U$55813 ( \56190 , RIae77450_76, \4245 );
nor \U$55814 ( \56191 , \56189 , \56190 );
and \U$55815 ( \56192 , \56191 , \4251 );
not \U$55816 ( \56193 , \56191 );
and \U$55817 ( \56194 , \56193 , \3989 );
nor \U$55818 ( \56195 , \56192 , \56194 );
and \U$55819 ( \56196 , \3730 , RIae77630_80);
and \U$55820 ( \56197 , RIae77540_78, \3728 );
nor \U$55821 ( \56198 , \56196 , \56197 );
and \U$55822 ( \56199 , \56198 , \3422 );
not \U$55823 ( \56200 , \56198 );
and \U$55824 ( \56201 , \56200 , \3732 );
nor \U$55825 ( \56202 , \56199 , \56201 );
xor \U$55826 ( \56203 , \56195 , \56202 );
and \U$55827 ( \56204 , \4688 , RIae77ae0_90);
and \U$55828 ( \56205 , RIae779f0_88, \4686 );
nor \U$55829 ( \56206 , \56204 , \56205 );
and \U$55830 ( \56207 , \56206 , \4482 );
not \U$55831 ( \56208 , \56206 );
and \U$55832 ( \56209 , \56208 , \4481 );
nor \U$55833 ( \56210 , \56207 , \56209 );
and \U$55834 ( \56211 , \56203 , \56210 );
and \U$55835 ( \56212 , \56195 , \56202 );
or \U$55836 ( \56213 , \56211 , \56212 );
not \U$55837 ( \56214 , \56213 );
and \U$55838 ( \56215 , \7633 , RIae77270_72);
and \U$55839 ( \56216 , RIae77360_74, \7631 );
nor \U$55840 ( \56217 , \56215 , \56216 );
and \U$55841 ( \56218 , \56217 , \7205 );
not \U$55842 ( \56219 , \56217 );
and \U$55843 ( \56220 , \56219 , \7206 );
nor \U$55844 ( \56221 , \56218 , \56220 );
and \U$55845 ( \56222 , \6941 , RIae77108_69);
and \U$55846 ( \56223 , RIae77090_68, \6939 );
nor \U$55847 ( \56224 , \56222 , \56223 );
and \U$55848 ( \56225 , \56224 , \6945 );
not \U$55849 ( \56226 , \56224 );
and \U$55850 ( \56227 , \56226 , \6314 );
nor \U$55851 ( \56228 , \56225 , \56227 );
xor \U$55852 ( \56229 , \56221 , \56228 );
and \U$55853 ( \56230 , \8371 , RIae78350_108);
and \U$55854 ( \56231 , RIae78170_104, \8369 );
nor \U$55855 ( \56232 , \56230 , \56231 );
and \U$55856 ( \56233 , \56232 , \8019 );
not \U$55857 ( \56234 , \56232 );
and \U$55858 ( \56235 , \56234 , \8020 );
nor \U$55859 ( \56236 , \56233 , \56235 );
and \U$55860 ( \56237 , \56229 , \56236 );
and \U$55861 ( \56238 , \56221 , \56228 );
or \U$55862 ( \56239 , \56237 , \56238 );
not \U$55863 ( \56240 , \56239 );
and \U$55864 ( \56241 , \56214 , \56240 );
and \U$55865 ( \56242 , \56213 , \56239 );
and \U$55866 ( \56243 , \6172 , RIae76dc0_62);
and \U$55867 ( \56244 , RIae76cd0_60, \6170 );
nor \U$55868 ( \56245 , \56243 , \56244 );
and \U$55869 ( \56246 , \56245 , \6175 );
not \U$55870 ( \56247 , \56245 );
and \U$55871 ( \56248 , \56247 , \6176 );
nor \U$55872 ( \56249 , \56246 , \56248 );
and \U$55873 ( \56250 , \5399 , RIae77810_84);
and \U$55874 ( \56251 , RIae77900_86, \5397 );
nor \U$55875 ( \56252 , \56250 , \56251 );
and \U$55876 ( \56253 , \56252 , \5403 );
not \U$55877 ( \56254 , \56252 );
and \U$55878 ( \56255 , \56254 , \5016 );
nor \U$55879 ( \56256 , \56253 , \56255 );
xor \U$55880 ( \56257 , \56249 , \56256 );
and \U$55881 ( \56258 , \5896 , RIae76fa0_66);
and \U$55882 ( \56259 , RIae76eb0_64, \5894 );
nor \U$55883 ( \56260 , \56258 , \56259 );
and \U$55884 ( \56261 , \56260 , \5589 );
not \U$55885 ( \56262 , \56260 );
and \U$55886 ( \56263 , \56262 , \5590 );
nor \U$55887 ( \56264 , \56261 , \56263 );
and \U$55888 ( \56265 , \56257 , \56264 );
and \U$55889 ( \56266 , \56249 , \56256 );
or \U$55890 ( \56267 , \56265 , \56266 );
nor \U$55891 ( \56268 , \56242 , \56267 );
nor \U$55892 ( \56269 , \56241 , \56268 );
and \U$55893 ( \56270 , \56188 , \56269 );
and \U$55894 ( \56271 , \56168 , \56187 );
or \U$55895 ( \56272 , \56270 , \56271 );
xor \U$55896 ( \56273 , \56085 , \56272 );
not \U$55897 ( \56274 , \55968 );
not \U$55898 ( \56275 , \55974 );
or \U$55899 ( \56276 , \56274 , \56275 );
or \U$55900 ( \56277 , \55974 , \55968 );
nand \U$55901 ( \56278 , \56276 , \56277 );
not \U$55902 ( \56279 , \56278 );
not \U$55903 ( \56280 , \55960 );
and \U$55904 ( \56281 , \56279 , \56280 );
and \U$55905 ( \56282 , \56278 , \55960 );
nor \U$55906 ( \56283 , \56281 , \56282 );
not \U$55907 ( \56284 , \56283 );
xor \U$55908 ( \56285 , \55819 , \55844 );
xor \U$55909 ( \56286 , \56285 , \55870 );
not \U$55910 ( \56287 , \56286 );
and \U$55911 ( \56288 , \56284 , \56287 );
and \U$55912 ( \56289 , \56283 , \56286 );
not \U$55913 ( \56290 , \55766 );
not \U$55914 ( \56291 , \55782 );
or \U$55915 ( \56292 , \56290 , \56291 );
or \U$55916 ( \56293 , \55766 , \55782 );
nand \U$55917 ( \56294 , \56292 , \56293 );
not \U$55918 ( \56295 , \56294 );
not \U$55919 ( \56296 , \55776 );
and \U$55920 ( \56297 , \56295 , \56296 );
and \U$55921 ( \56298 , \56294 , \55776 );
nor \U$55922 ( \56299 , \56297 , \56298 );
nor \U$55923 ( \56300 , \56289 , \56299 );
nor \U$55924 ( \56301 , \56288 , \56300 );
and \U$55925 ( \56302 , \56273 , \56301 );
and \U$55926 ( \56303 , \56085 , \56272 );
nor \U$55927 ( \56304 , \56302 , \56303 );
xor \U$55928 ( \56305 , \56047 , \56304 );
xor \U$55929 ( \56306 , \55603 , \55686 );
xor \U$55930 ( \56307 , \56306 , \55699 );
xor \U$55931 ( \56308 , \56004 , \56011 );
xor \U$55932 ( \56309 , \56307 , \56308 );
and \U$55933 ( \56310 , \56305 , \56309 );
and \U$55934 ( \56311 , \56047 , \56304 );
or \U$55935 ( \56312 , \56310 , \56311 );
nand \U$55936 ( \56313 , \56033 , \56312 );
nand \U$55937 ( \56314 , \56032 , \56313 );
nand \U$55938 ( \56315 , \56023 , \56314 );
nand \U$55939 ( \56316 , \56022 , \56315 );
xor \U$55940 ( \56317 , \55761 , \55763 );
and \U$55941 ( \56318 , \56317 , \56019 );
and \U$55942 ( \56319 , \55761 , \55763 );
or \U$55943 ( \56320 , \56318 , \56319 );
not \U$55944 ( \56321 , \56320 );
xor \U$55945 ( \56322 , \55730 , \55742 );
and \U$55946 ( \56323 , \56322 , \55747 );
and \U$55947 ( \56324 , \55730 , \55742 );
or \U$55948 ( \56325 , \56323 , \56324 );
xor \U$55949 ( \56326 , \55098 , \55100 );
xor \U$55950 ( \56327 , \56326 , \55113 );
xnor \U$55951 ( \56328 , \56325 , \56327 );
not \U$55952 ( \56329 , \56328 );
xor \U$55953 ( \56330 , \55118 , \55122 );
not \U$55954 ( \56331 , \56330 );
and \U$55955 ( \56332 , \56329 , \56331 );
and \U$55956 ( \56333 , \56328 , \56330 );
nor \U$55957 ( \56334 , \56332 , \56333 );
not \U$55958 ( \56335 , \56334 );
or \U$55959 ( \56336 , \56321 , \56335 );
or \U$55960 ( \56337 , \56334 , \56320 );
nand \U$55961 ( \56338 , \56336 , \56337 );
and \U$55962 ( \56339 , \56316 , \56338 );
xor \U$55963 ( \56340 , \56316 , \56338 );
xor \U$55964 ( \56341 , \56061 , \56071 );
xor \U$55965 ( \56342 , \56341 , \56082 );
xnor \U$55966 ( \56343 , \55947 , \55917 );
not \U$55967 ( \56344 , \56343 );
not \U$55968 ( \56345 , \55891 );
and \U$55969 ( \56346 , \56344 , \56345 );
and \U$55970 ( \56347 , \56343 , \55891 );
nor \U$55971 ( \56348 , \56346 , \56347 );
or \U$55972 ( \56349 , \56342 , \56348 );
not \U$55973 ( \56350 , \56348 );
not \U$55974 ( \56351 , \56342 );
or \U$55975 ( \56352 , \56350 , \56351 );
not \U$55976 ( \56353 , \56283 );
xor \U$55977 ( \56354 , \56286 , \56299 );
not \U$55978 ( \56355 , \56354 );
or \U$55979 ( \56356 , \56353 , \56355 );
or \U$55980 ( \56357 , \56354 , \56283 );
nand \U$55981 ( \56358 , \56356 , \56357 );
nand \U$55982 ( \56359 , \56352 , \56358 );
nand \U$55983 ( \56360 , \56349 , \56359 );
xor \U$55984 ( \56361 , \56110 , \56137 );
xor \U$55985 ( \56362 , \56361 , \56165 );
xor \U$55986 ( \56363 , \56174 , \56181 );
xor \U$55987 ( \56364 , \56363 , \56184 );
xor \U$55988 ( \56365 , \56362 , \56364 );
not \U$55989 ( \56366 , \56239 );
xor \U$55990 ( \56367 , \56213 , \56267 );
not \U$55991 ( \56368 , \56367 );
or \U$55992 ( \56369 , \56366 , \56368 );
or \U$55993 ( \56370 , \56367 , \56239 );
nand \U$55994 ( \56371 , \56369 , \56370 );
and \U$55995 ( \56372 , \56365 , \56371 );
and \U$55996 ( \56373 , \56362 , \56364 );
or \U$55997 ( \56374 , \56372 , \56373 );
and \U$55998 ( \56375 , \4688 , RIae77450_76);
and \U$55999 ( \56376 , RIae77ae0_90, \4686 );
nor \U$56000 ( \56377 , \56375 , \56376 );
and \U$56001 ( \56378 , \56377 , \4482 );
not \U$56002 ( \56379 , \56377 );
and \U$56003 ( \56380 , \56379 , \4481 );
nor \U$56004 ( \56381 , \56378 , \56380 );
and \U$56005 ( \56382 , \4247 , RIae77540_78);
and \U$56006 ( \56383 , RIae776a8_81, \4245 );
nor \U$56007 ( \56384 , \56382 , \56383 );
and \U$56008 ( \56385 , \56384 , \4251 );
not \U$56009 ( \56386 , \56384 );
and \U$56010 ( \56387 , \56386 , \3989 );
nor \U$56011 ( \56388 , \56385 , \56387 );
xor \U$56012 ( \56389 , \56381 , \56388 );
and \U$56013 ( \56390 , \5399 , RIae779f0_88);
and \U$56014 ( \56391 , RIae77810_84, \5397 );
nor \U$56015 ( \56392 , \56390 , \56391 );
and \U$56016 ( \56393 , \56392 , \5403 );
not \U$56017 ( \56394 , \56392 );
and \U$56018 ( \56395 , \56394 , \5016 );
nor \U$56019 ( \56396 , \56393 , \56395 );
and \U$56020 ( \56397 , \56389 , \56396 );
and \U$56021 ( \56398 , \56381 , \56388 );
or \U$56022 ( \56399 , \56397 , \56398 );
and \U$56023 ( \56400 , \5896 , RIae77900_86);
and \U$56024 ( \56401 , RIae76fa0_66, \5894 );
nor \U$56025 ( \56402 , \56400 , \56401 );
and \U$56026 ( \56403 , \56402 , \5589 );
not \U$56027 ( \56404 , \56402 );
and \U$56028 ( \56405 , \56404 , \5590 );
nor \U$56029 ( \56406 , \56403 , \56405 );
not \U$56030 ( \56407 , \56406 );
and \U$56031 ( \56408 , \6172 , RIae76eb0_64);
and \U$56032 ( \56409 , RIae76dc0_62, \6170 );
nor \U$56033 ( \56410 , \56408 , \56409 );
and \U$56034 ( \56411 , \56410 , \6175 );
not \U$56035 ( \56412 , \56410 );
and \U$56036 ( \56413 , \56412 , \6176 );
nor \U$56037 ( \56414 , \56411 , \56413 );
not \U$56038 ( \56415 , \56414 );
and \U$56039 ( \56416 , \56407 , \56415 );
and \U$56040 ( \56417 , \56414 , \56406 );
and \U$56041 ( \56418 , \6941 , RIae76cd0_60);
and \U$56042 ( \56419 , RIae77108_69, \6939 );
nor \U$56043 ( \56420 , \56418 , \56419 );
and \U$56044 ( \56421 , \56420 , \6945 );
not \U$56045 ( \56422 , \56420 );
and \U$56046 ( \56423 , \56422 , \6314 );
nor \U$56047 ( \56424 , \56421 , \56423 );
nor \U$56048 ( \56425 , \56417 , \56424 );
nor \U$56049 ( \56426 , \56416 , \56425 );
or \U$56050 ( \56427 , \56399 , \56426 );
not \U$56051 ( \56428 , \56399 );
not \U$56052 ( \56429 , \56426 );
or \U$56053 ( \56430 , \56428 , \56429 );
and \U$56054 ( \56431 , \8371 , RIae77360_74);
and \U$56055 ( \56432 , RIae78350_108, \8369 );
nor \U$56056 ( \56433 , \56431 , \56432 );
and \U$56057 ( \56434 , \56433 , \8019 );
not \U$56058 ( \56435 , \56433 );
and \U$56059 ( \56436 , \56435 , \8020 );
nor \U$56060 ( \56437 , \56434 , \56436 );
and \U$56061 ( \56438 , \8966 , RIae78170_104);
and \U$56062 ( \56439 , RIae77f90_100, \8964 );
nor \U$56063 ( \56440 , \56438 , \56439 );
and \U$56064 ( \56441 , \56440 , \8789 );
not \U$56065 ( \56442 , \56440 );
and \U$56066 ( \56443 , \56442 , \8799 );
nor \U$56067 ( \56444 , \56441 , \56443 );
xor \U$56068 ( \56445 , \56437 , \56444 );
and \U$56069 ( \56446 , \7633 , RIae77090_68);
and \U$56070 ( \56447 , RIae77270_72, \7631 );
nor \U$56071 ( \56448 , \56446 , \56447 );
and \U$56072 ( \56449 , \56448 , \7205 );
not \U$56073 ( \56450 , \56448 );
and \U$56074 ( \56451 , \56450 , \7206 );
nor \U$56075 ( \56452 , \56449 , \56451 );
and \U$56076 ( \56453 , \56445 , \56452 );
and \U$56077 ( \56454 , \56437 , \56444 );
nor \U$56078 ( \56455 , \56453 , \56454 );
nand \U$56079 ( \56456 , \56430 , \56455 );
nand \U$56080 ( \56457 , \56427 , \56456 );
and \U$56081 ( \56458 , \13059 , RIae77ea0_98);
and \U$56082 ( \56459 , RIae789e0_122, \13057 );
nor \U$56083 ( \56460 , \56458 , \56459 );
and \U$56084 ( \56461 , \56460 , \12718 );
not \U$56085 ( \56462 , \56460 );
and \U$56086 ( \56463 , \56462 , \13063 );
nor \U$56087 ( \56464 , \56461 , \56463 );
and \U$56088 ( \56465 , \14059 , RIae788f0_120);
and \U$56089 ( \56466 , RIae78800_118, \14057 );
nor \U$56090 ( \56467 , \56465 , \56466 );
and \U$56091 ( \56468 , \56467 , \14063 );
not \U$56092 ( \56469 , \56467 );
and \U$56093 ( \56470 , \56469 , \13502 );
nor \U$56094 ( \56471 , \56468 , \56470 );
xor \U$56095 ( \56472 , \56464 , \56471 );
and \U$56096 ( \56473 , \12180 , RIae77bd0_92);
and \U$56097 ( \56474 , RIae77db0_96, \12178 );
nor \U$56098 ( \56475 , \56473 , \56474 );
and \U$56099 ( \56476 , \56475 , \11827 );
not \U$56100 ( \56477 , \56475 );
and \U$56101 ( \56478 , \56477 , \12184 );
nor \U$56102 ( \56479 , \56476 , \56478 );
and \U$56103 ( \56480 , \56472 , \56479 );
and \U$56104 ( \56481 , \56464 , \56471 );
nor \U$56105 ( \56482 , \56480 , \56481 );
and \U$56106 ( \56483 , \15726 , RIae75b00_22);
and \U$56107 ( \56484 , RIae75a10_20, RIae7aab0_192);
nor \U$56108 ( \56485 , \56483 , \56484 );
and \U$56109 ( \56486 , \56485 , RIae7aa38_191);
not \U$56110 ( \56487 , \56485 );
and \U$56111 ( \56488 , \56487 , \14959 );
nor \U$56112 ( \56489 , \56486 , \56488 );
or \U$56113 ( \56490 , \56489 , \3732 );
not \U$56114 ( \56491 , \3732 );
not \U$56115 ( \56492 , \56489 );
or \U$56116 ( \56493 , \56491 , \56492 );
and \U$56117 ( \56494 , \14964 , RIae78710_116);
and \U$56118 ( \56495 , RIae75bf0_24, \14962 );
nor \U$56119 ( \56496 , \56494 , \56495 );
and \U$56120 ( \56497 , \56496 , \14463 );
not \U$56121 ( \56498 , \56496 );
and \U$56122 ( \56499 , \56498 , \14462 );
nor \U$56123 ( \56500 , \56497 , \56499 );
nand \U$56124 ( \56501 , \56493 , \56500 );
nand \U$56125 ( \56502 , \56490 , \56501 );
xor \U$56126 ( \56503 , \56482 , \56502 );
and \U$56127 ( \56504 , \9760 , RIae78080_102);
and \U$56128 ( \56505 , RIae78260_106, \9758 );
nor \U$56129 ( \56506 , \56504 , \56505 );
and \U$56130 ( \56507 , \56506 , \9272 );
not \U$56131 ( \56508 , \56506 );
and \U$56132 ( \56509 , \56508 , \9273 );
nor \U$56133 ( \56510 , \56507 , \56509 );
and \U$56134 ( \56511 , \11470 , RIae784b8_111);
and \U$56135 ( \56512 , RIae77cc0_94, \11468 );
nor \U$56136 ( \56513 , \56511 , \56512 );
and \U$56137 ( \56514 , \56513 , \11474 );
not \U$56138 ( \56515 , \56513 );
and \U$56139 ( \56516 , \56515 , \10936 );
nor \U$56140 ( \56517 , \56514 , \56516 );
or \U$56141 ( \56518 , \56510 , \56517 );
not \U$56142 ( \56519 , \56517 );
not \U$56143 ( \56520 , \56510 );
or \U$56144 ( \56521 , \56519 , \56520 );
and \U$56145 ( \56522 , \10548 , RIae78620_114);
and \U$56146 ( \56523 , RIae78440_110, \10546 );
nor \U$56147 ( \56524 , \56522 , \56523 );
and \U$56148 ( \56525 , \56524 , \10421 );
not \U$56149 ( \56526 , \56524 );
and \U$56150 ( \56527 , \56526 , \10118 );
nor \U$56151 ( \56528 , \56525 , \56527 );
nand \U$56152 ( \56529 , \56521 , \56528 );
nand \U$56153 ( \56530 , \56518 , \56529 );
and \U$56154 ( \56531 , \56503 , \56530 );
and \U$56155 ( \56532 , \56482 , \56502 );
or \U$56156 ( \56533 , \56531 , \56532 );
xor \U$56157 ( \56534 , \56457 , \56533 );
xor \U$56158 ( \56535 , \56195 , \56202 );
xor \U$56159 ( \56536 , \56535 , \56210 );
xor \U$56160 ( \56537 , \56249 , \56256 );
xor \U$56161 ( \56538 , \56537 , \56264 );
xor \U$56162 ( \56539 , \56536 , \56538 );
xor \U$56163 ( \56540 , \56221 , \56228 );
xor \U$56164 ( \56541 , \56540 , \56236 );
and \U$56165 ( \56542 , \56539 , \56541 );
and \U$56166 ( \56543 , \56536 , \56538 );
nor \U$56167 ( \56544 , \56542 , \56543 );
and \U$56168 ( \56545 , \56534 , \56544 );
and \U$56169 ( \56546 , \56457 , \56533 );
or \U$56170 ( \56547 , \56545 , \56546 );
xor \U$56171 ( \56548 , \56374 , \56547 );
not \U$56172 ( \56549 , \56124 );
not \U$56173 ( \56550 , \56135 );
or \U$56174 ( \56551 , \56549 , \56550 );
or \U$56175 ( \56552 , \56135 , \56124 );
nand \U$56176 ( \56553 , \56551 , \56552 );
not \U$56177 ( \56554 , \56553 );
not \U$56178 ( \56555 , \56117 );
and \U$56179 ( \56556 , \56554 , \56555 );
and \U$56180 ( \56557 , \56553 , \56117 );
nor \U$56181 ( \56558 , \56556 , \56557 );
not \U$56182 ( \56559 , \56152 );
not \U$56183 ( \56560 , \56163 );
or \U$56184 ( \56561 , \56559 , \56560 );
or \U$56185 ( \56562 , \56152 , \56163 );
nand \U$56186 ( \56563 , \56561 , \56562 );
not \U$56187 ( \56564 , \56563 );
not \U$56188 ( \56565 , \56145 );
and \U$56189 ( \56566 , \56564 , \56565 );
and \U$56190 ( \56567 , \56563 , \56145 );
nor \U$56191 ( \56568 , \56566 , \56567 );
or \U$56192 ( \56569 , \56558 , \56568 );
not \U$56193 ( \56570 , \56568 );
not \U$56194 ( \56571 , \56558 );
or \U$56195 ( \56572 , \56570 , \56571 );
xor \U$56196 ( \56573 , \56092 , \56099 );
xor \U$56197 ( \56574 , \56573 , \56107 );
nand \U$56198 ( \56575 , \56572 , \56574 );
nand \U$56199 ( \56576 , \56569 , \56575 );
not \U$56200 ( \56577 , \56057 );
not \U$56201 ( \56578 , \56060 );
or \U$56202 ( \56579 , \56577 , \56578 );
or \U$56203 ( \56580 , \56060 , \56057 );
nand \U$56204 ( \56581 , \56579 , \56580 );
xor \U$56205 ( \56582 , \56576 , \56581 );
xor \U$56206 ( \56583 , \56074 , \56076 );
xor \U$56207 ( \56584 , \56583 , \56079 );
and \U$56208 ( \56585 , \56582 , \56584 );
and \U$56209 ( \56586 , \56576 , \56581 );
or \U$56210 ( \56587 , \56585 , \56586 );
and \U$56211 ( \56588 , \56548 , \56587 );
and \U$56212 ( \56589 , \56374 , \56547 );
or \U$56213 ( \56590 , \56588 , \56589 );
xor \U$56214 ( \56591 , \56360 , \56590 );
xor \U$56215 ( \56592 , \55784 , \55786 );
xor \U$56216 ( \56593 , \56592 , \55791 );
xor \U$56217 ( \56594 , \56035 , \56042 );
xor \U$56218 ( \56595 , \56593 , \56594 );
and \U$56219 ( \56596 , \56591 , \56595 );
and \U$56220 ( \56597 , \56360 , \56590 );
or \U$56221 ( \56598 , \56596 , \56597 );
xor \U$56222 ( \56599 , \55794 , \55979 );
xor \U$56223 ( \56600 , \56599 , \55994 );
xor \U$56224 ( \56601 , \56598 , \56600 );
xor \U$56225 ( \56602 , \56047 , \56304 );
xor \U$56226 ( \56603 , \56602 , \56309 );
xor \U$56227 ( \56604 , \56601 , \56603 );
not \U$56228 ( \56605 , \56604 );
xnor \U$56229 ( \56606 , \56348 , \56342 );
not \U$56230 ( \56607 , \56606 );
not \U$56231 ( \56608 , \56358 );
and \U$56232 ( \56609 , \56607 , \56608 );
and \U$56233 ( \56610 , \56606 , \56358 );
nor \U$56234 ( \56611 , \56609 , \56610 );
not \U$56235 ( \56612 , \56611 );
xor \U$56236 ( \56613 , \56374 , \56547 );
xor \U$56237 ( \56614 , \56613 , \56587 );
nand \U$56238 ( \56615 , \56612 , \56614 );
xor \U$56239 ( \56616 , \56085 , \56272 );
xor \U$56240 ( \56617 , \56616 , \56301 );
xor \U$56241 ( \56618 , \56615 , \56617 );
and \U$56242 ( \56619 , \12180 , RIae77cc0_94);
and \U$56243 ( \56620 , RIae77bd0_92, \12178 );
nor \U$56244 ( \56621 , \56619 , \56620 );
and \U$56245 ( \56622 , \56621 , \11827 );
not \U$56246 ( \56623 , \56621 );
and \U$56247 ( \56624 , \56623 , \12184 );
nor \U$56248 ( \56625 , \56622 , \56624 );
and \U$56249 ( \56626 , \11470 , RIae78440_110);
and \U$56250 ( \56627 , RIae784b8_111, \11468 );
nor \U$56251 ( \56628 , \56626 , \56627 );
and \U$56252 ( \56629 , \56628 , \11474 );
not \U$56253 ( \56630 , \56628 );
and \U$56254 ( \56631 , \56630 , \10936 );
nor \U$56255 ( \56632 , \56629 , \56631 );
xor \U$56256 ( \56633 , \56625 , \56632 );
and \U$56257 ( \56634 , \13059 , RIae77db0_96);
and \U$56258 ( \56635 , RIae77ea0_98, \13057 );
nor \U$56259 ( \56636 , \56634 , \56635 );
and \U$56260 ( \56637 , \56636 , \12718 );
not \U$56261 ( \56638 , \56636 );
and \U$56262 ( \56639 , \56638 , \13063 );
nor \U$56263 ( \56640 , \56637 , \56639 );
and \U$56264 ( \56641 , \56633 , \56640 );
and \U$56265 ( \56642 , \56625 , \56632 );
or \U$56266 ( \56643 , \56641 , \56642 );
and \U$56267 ( \56644 , \14059 , RIae789e0_122);
and \U$56268 ( \56645 , RIae788f0_120, \14057 );
nor \U$56269 ( \56646 , \56644 , \56645 );
and \U$56270 ( \56647 , \56646 , \14063 );
not \U$56271 ( \56648 , \56646 );
and \U$56272 ( \56649 , \56648 , \13502 );
nor \U$56273 ( \56650 , \56647 , \56649 );
and \U$56274 ( \56651 , \15726 , RIae75bf0_24);
and \U$56275 ( \56652 , RIae75b00_22, RIae7aab0_192);
nor \U$56276 ( \56653 , \56651 , \56652 );
and \U$56277 ( \56654 , \56653 , RIae7aa38_191);
not \U$56278 ( \56655 , \56653 );
and \U$56279 ( \56656 , \56655 , \14959 );
nor \U$56280 ( \56657 , \56654 , \56656 );
xor \U$56281 ( \56658 , \56650 , \56657 );
and \U$56282 ( \56659 , \14964 , RIae78800_118);
and \U$56283 ( \56660 , RIae78710_116, \14962 );
nor \U$56284 ( \56661 , \56659 , \56660 );
and \U$56285 ( \56662 , \56661 , \14462 );
not \U$56286 ( \56663 , \56661 );
and \U$56287 ( \56664 , \56663 , \14463 );
nor \U$56288 ( \56665 , \56662 , \56664 );
and \U$56289 ( \56666 , \56658 , \56665 );
and \U$56290 ( \56667 , \56650 , \56657 );
or \U$56291 ( \56668 , \56666 , \56667 );
or \U$56292 ( \56669 , \56643 , \56668 );
not \U$56293 ( \56670 , \56668 );
not \U$56294 ( \56671 , \56643 );
or \U$56295 ( \56672 , \56670 , \56671 );
and \U$56296 ( \56673 , \9760 , RIae77f90_100);
and \U$56297 ( \56674 , RIae78080_102, \9758 );
nor \U$56298 ( \56675 , \56673 , \56674 );
and \U$56299 ( \56676 , \56675 , \9272 );
not \U$56300 ( \56677 , \56675 );
and \U$56301 ( \56678 , \56677 , \9273 );
nor \U$56302 ( \56679 , \56676 , \56678 );
and \U$56303 ( \56680 , \10548 , RIae78260_106);
and \U$56304 ( \56681 , RIae78620_114, \10546 );
nor \U$56305 ( \56682 , \56680 , \56681 );
and \U$56306 ( \56683 , \56682 , \10118 );
not \U$56307 ( \56684 , \56682 );
and \U$56308 ( \56685 , \56684 , \10421 );
nor \U$56309 ( \56686 , \56683 , \56685 );
xor \U$56310 ( \56687 , \56679 , \56686 );
and \U$56311 ( \56688 , \8966 , RIae78350_108);
and \U$56312 ( \56689 , RIae78170_104, \8964 );
nor \U$56313 ( \56690 , \56688 , \56689 );
and \U$56314 ( \56691 , \56690 , \8789 );
not \U$56315 ( \56692 , \56690 );
and \U$56316 ( \56693 , \56692 , \8799 );
nor \U$56317 ( \56694 , \56691 , \56693 );
and \U$56318 ( \56695 , \56687 , \56694 );
and \U$56319 ( \56696 , \56679 , \56686 );
nor \U$56320 ( \56697 , \56695 , \56696 );
nand \U$56321 ( \56698 , \56672 , \56697 );
nand \U$56322 ( \56699 , \56669 , \56698 );
and \U$56323 ( \56700 , \4688 , RIae776a8_81);
and \U$56324 ( \56701 , RIae77450_76, \4686 );
nor \U$56325 ( \56702 , \56700 , \56701 );
and \U$56326 ( \56703 , \56702 , \4481 );
not \U$56327 ( \56704 , \56702 );
and \U$56328 ( \56705 , \56704 , \4482 );
nor \U$56329 ( \56706 , \56703 , \56705 );
and \U$56330 ( \56707 , \4247 , RIae77630_80);
and \U$56331 ( \56708 , RIae77540_78, \4245 );
nor \U$56332 ( \56709 , \56707 , \56708 );
and \U$56333 ( \56710 , \56709 , \3989 );
not \U$56334 ( \56711 , \56709 );
and \U$56335 ( \56712 , \56711 , \4251 );
nor \U$56336 ( \56713 , \56710 , \56712 );
and \U$56337 ( \56714 , \56706 , \56713 );
not \U$56338 ( \56715 , \56714 );
and \U$56339 ( \56716 , \8371 , RIae77270_72);
and \U$56340 ( \56717 , RIae77360_74, \8369 );
nor \U$56341 ( \56718 , \56716 , \56717 );
and \U$56342 ( \56719 , \56718 , \8020 );
not \U$56343 ( \56720 , \56718 );
and \U$56344 ( \56721 , \56720 , \8019 );
nor \U$56345 ( \56722 , \56719 , \56721 );
and \U$56346 ( \56723 , \6941 , RIae76dc0_62);
and \U$56347 ( \56724 , RIae76cd0_60, \6939 );
nor \U$56348 ( \56725 , \56723 , \56724 );
and \U$56349 ( \56726 , \56725 , \6314 );
not \U$56350 ( \56727 , \56725 );
and \U$56351 ( \56728 , \56727 , \6945 );
nor \U$56352 ( \56729 , \56726 , \56728 );
xor \U$56353 ( \56730 , \56722 , \56729 );
and \U$56354 ( \56731 , \7633 , RIae77108_69);
and \U$56355 ( \56732 , RIae77090_68, \7631 );
nor \U$56356 ( \56733 , \56731 , \56732 );
and \U$56357 ( \56734 , \56733 , \7206 );
not \U$56358 ( \56735 , \56733 );
and \U$56359 ( \56736 , \56735 , \7205 );
nor \U$56360 ( \56737 , \56734 , \56736 );
and \U$56361 ( \56738 , \56730 , \56737 );
and \U$56362 ( \56739 , \56722 , \56729 );
or \U$56363 ( \56740 , \56738 , \56739 );
not \U$56364 ( \56741 , \56740 );
or \U$56365 ( \56742 , \56715 , \56741 );
or \U$56366 ( \56743 , \56740 , \56714 );
and \U$56367 ( \56744 , \5399 , RIae77ae0_90);
and \U$56368 ( \56745 , RIae779f0_88, \5397 );
nor \U$56369 ( \56746 , \56744 , \56745 );
and \U$56370 ( \56747 , \56746 , \5016 );
not \U$56371 ( \56748 , \56746 );
and \U$56372 ( \56749 , \56748 , \5403 );
nor \U$56373 ( \56750 , \56747 , \56749 );
and \U$56374 ( \56751 , \5896 , RIae77810_84);
and \U$56375 ( \56752 , RIae77900_86, \5894 );
nor \U$56376 ( \56753 , \56751 , \56752 );
and \U$56377 ( \56754 , \56753 , \5590 );
not \U$56378 ( \56755 , \56753 );
and \U$56379 ( \56756 , \56755 , \5589 );
nor \U$56380 ( \56757 , \56754 , \56756 );
xor \U$56381 ( \56758 , \56750 , \56757 );
and \U$56382 ( \56759 , \6172 , RIae76fa0_66);
and \U$56383 ( \56760 , RIae76eb0_64, \6170 );
nor \U$56384 ( \56761 , \56759 , \56760 );
and \U$56385 ( \56762 , \56761 , \6176 );
not \U$56386 ( \56763 , \56761 );
and \U$56387 ( \56764 , \56763 , \6175 );
nor \U$56388 ( \56765 , \56762 , \56764 );
and \U$56389 ( \56766 , \56758 , \56765 );
and \U$56390 ( \56767 , \56750 , \56757 );
or \U$56391 ( \56768 , \56766 , \56767 );
nand \U$56392 ( \56769 , \56743 , \56768 );
nand \U$56393 ( \56770 , \56742 , \56769 );
xor \U$56394 ( \56771 , \56699 , \56770 );
xor \U$56395 ( \56772 , \56381 , \56388 );
xor \U$56396 ( \56773 , \56772 , \56396 );
nand \U$56397 ( \56774 , RIae77630_80, \3728 );
and \U$56398 ( \56775 , \56774 , \3422 );
not \U$56399 ( \56776 , \56774 );
and \U$56400 ( \56777 , \56776 , \3732 );
nor \U$56401 ( \56778 , \56775 , \56777 );
or \U$56402 ( \56779 , \56773 , \56778 );
not \U$56403 ( \56780 , \56778 );
not \U$56404 ( \56781 , \56773 );
or \U$56405 ( \56782 , \56780 , \56781 );
not \U$56406 ( \56783 , \56406 );
xor \U$56407 ( \56784 , \56414 , \56424 );
not \U$56408 ( \56785 , \56784 );
or \U$56409 ( \56786 , \56783 , \56785 );
or \U$56410 ( \56787 , \56784 , \56406 );
nand \U$56411 ( \56788 , \56786 , \56787 );
nand \U$56412 ( \56789 , \56782 , \56788 );
nand \U$56413 ( \56790 , \56779 , \56789 );
and \U$56414 ( \56791 , \56771 , \56790 );
and \U$56415 ( \56792 , \56699 , \56770 );
nor \U$56416 ( \56793 , \56791 , \56792 );
not \U$56417 ( \56794 , \56455 );
not \U$56418 ( \56795 , \56426 );
or \U$56419 ( \56796 , \56794 , \56795 );
or \U$56420 ( \56797 , \56426 , \56455 );
nand \U$56421 ( \56798 , \56796 , \56797 );
not \U$56422 ( \56799 , \56798 );
not \U$56423 ( \56800 , \56399 );
and \U$56424 ( \56801 , \56799 , \56800 );
and \U$56425 ( \56802 , \56798 , \56399 );
nor \U$56426 ( \56803 , \56801 , \56802 );
not \U$56427 ( \56804 , \56803 );
xor \U$56428 ( \56805 , \56482 , \56502 );
xor \U$56429 ( \56806 , \56805 , \56530 );
nand \U$56430 ( \56807 , \56804 , \56806 );
xor \U$56431 ( \56808 , \56793 , \56807 );
not \U$56432 ( \56809 , \56574 );
not \U$56433 ( \56810 , \56558 );
or \U$56434 ( \56811 , \56809 , \56810 );
or \U$56435 ( \56812 , \56558 , \56574 );
nand \U$56436 ( \56813 , \56811 , \56812 );
not \U$56437 ( \56814 , \56813 );
not \U$56438 ( \56815 , \56568 );
and \U$56439 ( \56816 , \56814 , \56815 );
and \U$56440 ( \56817 , \56813 , \56568 );
nor \U$56441 ( \56818 , \56816 , \56817 );
not \U$56442 ( \56819 , \56818 );
xor \U$56443 ( \56820 , \56536 , \56538 );
xor \U$56444 ( \56821 , \56820 , \56541 );
not \U$56445 ( \56822 , \56821 );
and \U$56446 ( \56823 , \56819 , \56822 );
and \U$56447 ( \56824 , \56818 , \56821 );
xor \U$56448 ( \56825 , \56464 , \56471 );
xor \U$56449 ( \56826 , \56825 , \56479 );
xor \U$56450 ( \56827 , \56437 , \56444 );
xor \U$56451 ( \56828 , \56827 , \56452 );
xor \U$56452 ( \56829 , \56826 , \56828 );
not \U$56453 ( \56830 , \56517 );
not \U$56454 ( \56831 , \56528 );
or \U$56455 ( \56832 , \56830 , \56831 );
or \U$56456 ( \56833 , \56517 , \56528 );
nand \U$56457 ( \56834 , \56832 , \56833 );
not \U$56458 ( \56835 , \56834 );
not \U$56459 ( \56836 , \56510 );
and \U$56460 ( \56837 , \56835 , \56836 );
and \U$56461 ( \56838 , \56834 , \56510 );
nor \U$56462 ( \56839 , \56837 , \56838 );
and \U$56463 ( \56840 , \56829 , \56839 );
and \U$56464 ( \56841 , \56826 , \56828 );
or \U$56465 ( \56842 , \56840 , \56841 );
nor \U$56466 ( \56843 , \56824 , \56842 );
nor \U$56467 ( \56844 , \56823 , \56843 );
and \U$56468 ( \56845 , \56808 , \56844 );
and \U$56469 ( \56846 , \56793 , \56807 );
or \U$56470 ( \56847 , \56845 , \56846 );
xor \U$56471 ( \56848 , \56168 , \56187 );
xor \U$56472 ( \56849 , \56848 , \56269 );
xor \U$56473 ( \56850 , \56847 , \56849 );
xor \U$56474 ( \56851 , \56457 , \56533 );
xor \U$56475 ( \56852 , \56851 , \56544 );
xor \U$56476 ( \56853 , \56362 , \56364 );
xor \U$56477 ( \56854 , \56853 , \56371 );
and \U$56478 ( \56855 , \56852 , \56854 );
xor \U$56479 ( \56856 , \56576 , \56581 );
xor \U$56480 ( \56857 , \56856 , \56584 );
xor \U$56481 ( \56858 , \56362 , \56364 );
xor \U$56482 ( \56859 , \56858 , \56371 );
and \U$56483 ( \56860 , \56857 , \56859 );
and \U$56484 ( \56861 , \56852 , \56857 );
or \U$56485 ( \56862 , \56855 , \56860 , \56861 );
not \U$56486 ( \56863 , \56862 );
and \U$56487 ( \56864 , \56850 , \56863 );
and \U$56488 ( \56865 , \56847 , \56849 );
or \U$56489 ( \56866 , \56864 , \56865 );
and \U$56490 ( \56867 , \56618 , \56866 );
and \U$56491 ( \56868 , \56615 , \56617 );
or \U$56492 ( \56869 , \56867 , \56868 );
not \U$56493 ( \56870 , \56869 );
and \U$56494 ( \56871 , \56605 , \56870 );
and \U$56495 ( \56872 , \56604 , \56869 );
nor \U$56496 ( \56873 , \56871 , \56872 );
xor \U$56497 ( \56874 , \56615 , \56617 );
xor \U$56498 ( \56875 , \56874 , \56866 );
not \U$56499 ( \56876 , \56875 );
xor \U$56500 ( \56877 , \56360 , \56590 );
xor \U$56501 ( \56878 , \56877 , \56595 );
nand \U$56502 ( \56879 , \56876 , \56878 );
or \U$56503 ( \56880 , \56873 , \56879 );
xnor \U$56504 ( \56881 , \56879 , \56873 );
not \U$56505 ( \56882 , \56878 );
not \U$56506 ( \56883 , \56875 );
or \U$56507 ( \56884 , \56882 , \56883 );
or \U$56508 ( \56885 , \56875 , \56878 );
nand \U$56509 ( \56886 , \56884 , \56885 );
xor \U$56510 ( \56887 , \56847 , \56849 );
xor \U$56511 ( \56888 , \56887 , \56863 );
not \U$56512 ( \56889 , \56611 );
not \U$56513 ( \56890 , \56614 );
and \U$56514 ( \56891 , \56889 , \56890 );
and \U$56515 ( \56892 , \56611 , \56614 );
nor \U$56516 ( \56893 , \56891 , \56892 );
or \U$56517 ( \56894 , \56888 , \56893 );
not \U$56518 ( \56895 , \56893 );
not \U$56519 ( \56896 , \56888 );
or \U$56520 ( \56897 , \56895 , \56896 );
and \U$56521 ( \56898 , \5399 , RIae77450_76);
and \U$56522 ( \56899 , RIae77ae0_90, \5397 );
nor \U$56523 ( \56900 , \56898 , \56899 );
and \U$56524 ( \56901 , \56900 , \5403 );
not \U$56525 ( \56902 , \56900 );
and \U$56526 ( \56903 , \56902 , \5016 );
nor \U$56527 ( \56904 , \56901 , \56903 );
nand \U$56528 ( \56905 , RIae77630_80, \4245 );
and \U$56529 ( \56906 , \56905 , \4251 );
not \U$56530 ( \56907 , \56905 );
and \U$56531 ( \56908 , \56907 , \3989 );
nor \U$56532 ( \56909 , \56906 , \56908 );
xor \U$56533 ( \56910 , \56904 , \56909 );
and \U$56534 ( \56911 , \4688 , RIae77540_78);
and \U$56535 ( \56912 , RIae776a8_81, \4686 );
nor \U$56536 ( \56913 , \56911 , \56912 );
and \U$56537 ( \56914 , \56913 , \4482 );
not \U$56538 ( \56915 , \56913 );
and \U$56539 ( \56916 , \56915 , \4481 );
nor \U$56540 ( \56917 , \56914 , \56916 );
and \U$56541 ( \56918 , \56910 , \56917 );
and \U$56542 ( \56919 , \56904 , \56909 );
or \U$56543 ( \56920 , \56918 , \56919 );
and \U$56544 ( \56921 , \5896 , RIae779f0_88);
and \U$56545 ( \56922 , RIae77810_84, \5894 );
nor \U$56546 ( \56923 , \56921 , \56922 );
and \U$56547 ( \56924 , \56923 , \5589 );
not \U$56548 ( \56925 , \56923 );
and \U$56549 ( \56926 , \56925 , \5590 );
nor \U$56550 ( \56927 , \56924 , \56926 );
not \U$56551 ( \56928 , \56927 );
and \U$56552 ( \56929 , \6172 , RIae77900_86);
and \U$56553 ( \56930 , RIae76fa0_66, \6170 );
nor \U$56554 ( \56931 , \56929 , \56930 );
and \U$56555 ( \56932 , \56931 , \6175 );
not \U$56556 ( \56933 , \56931 );
and \U$56557 ( \56934 , \56933 , \6176 );
nor \U$56558 ( \56935 , \56932 , \56934 );
not \U$56559 ( \56936 , \56935 );
and \U$56560 ( \56937 , \56928 , \56936 );
and \U$56561 ( \56938 , \56935 , \56927 );
and \U$56562 ( \56939 , \6941 , RIae76eb0_64);
and \U$56563 ( \56940 , RIae76dc0_62, \6939 );
nor \U$56564 ( \56941 , \56939 , \56940 );
and \U$56565 ( \56942 , \56941 , \6945 );
not \U$56566 ( \56943 , \56941 );
and \U$56567 ( \56944 , \56943 , \6314 );
nor \U$56568 ( \56945 , \56942 , \56944 );
nor \U$56569 ( \56946 , \56938 , \56945 );
nor \U$56570 ( \56947 , \56937 , \56946 );
xor \U$56571 ( \56948 , \56920 , \56947 );
and \U$56572 ( \56949 , \7633 , RIae76cd0_60);
and \U$56573 ( \56950 , RIae77108_69, \7631 );
nor \U$56574 ( \56951 , \56949 , \56950 );
and \U$56575 ( \56952 , \56951 , \7205 );
not \U$56576 ( \56953 , \56951 );
and \U$56577 ( \56954 , \56953 , \7206 );
nor \U$56578 ( \56955 , \56952 , \56954 );
not \U$56579 ( \56956 , \56955 );
and \U$56580 ( \56957 , \8371 , RIae77090_68);
and \U$56581 ( \56958 , RIae77270_72, \8369 );
nor \U$56582 ( \56959 , \56957 , \56958 );
and \U$56583 ( \56960 , \56959 , \8019 );
not \U$56584 ( \56961 , \56959 );
and \U$56585 ( \56962 , \56961 , \8020 );
nor \U$56586 ( \56963 , \56960 , \56962 );
not \U$56587 ( \56964 , \56963 );
and \U$56588 ( \56965 , \56956 , \56964 );
and \U$56589 ( \56966 , \56963 , \56955 );
and \U$56590 ( \56967 , \8966 , RIae77360_74);
and \U$56591 ( \56968 , RIae78350_108, \8964 );
nor \U$56592 ( \56969 , \56967 , \56968 );
and \U$56593 ( \56970 , \56969 , \8789 );
not \U$56594 ( \56971 , \56969 );
and \U$56595 ( \56972 , \56971 , \8799 );
nor \U$56596 ( \56973 , \56970 , \56972 );
nor \U$56597 ( \56974 , \56966 , \56973 );
nor \U$56598 ( \56975 , \56965 , \56974 );
and \U$56599 ( \56976 , \56948 , \56975 );
and \U$56600 ( \56977 , \56920 , \56947 );
nor \U$56601 ( \56978 , \56976 , \56977 );
and \U$56602 ( \56979 , \9760 , RIae78170_104);
and \U$56603 ( \56980 , RIae77f90_100, \9758 );
nor \U$56604 ( \56981 , \56979 , \56980 );
and \U$56605 ( \56982 , \56981 , \9273 );
not \U$56606 ( \56983 , \56981 );
and \U$56607 ( \56984 , \56983 , \9764 );
nor \U$56608 ( \56985 , \56982 , \56984 );
and \U$56609 ( \56986 , \10548 , RIae78080_102);
and \U$56610 ( \56987 , RIae78260_106, \10546 );
nor \U$56611 ( \56988 , \56986 , \56987 );
and \U$56612 ( \56989 , \56988 , \10421 );
not \U$56613 ( \56990 , \56988 );
and \U$56614 ( \56991 , \56990 , \10118 );
nor \U$56615 ( \56992 , \56989 , \56991 );
xor \U$56616 ( \56993 , \56985 , \56992 );
and \U$56617 ( \56994 , \11470 , RIae78620_114);
and \U$56618 ( \56995 , RIae78440_110, \11468 );
nor \U$56619 ( \56996 , \56994 , \56995 );
and \U$56620 ( \56997 , \56996 , \10936 );
not \U$56621 ( \56998 , \56996 );
and \U$56622 ( \56999 , \56998 , \11474 );
nor \U$56623 ( \57000 , \56997 , \56999 );
and \U$56624 ( \57001 , \56993 , \57000 );
and \U$56625 ( \57002 , \56985 , \56992 );
or \U$56626 ( \57003 , \57001 , \57002 );
and \U$56627 ( \57004 , \15726 , RIae78710_116);
and \U$56628 ( \57005 , RIae75bf0_24, RIae7aab0_192);
nor \U$56629 ( \57006 , \57004 , \57005 );
and \U$56630 ( \57007 , \57006 , \14959 );
not \U$56631 ( \57008 , \57006 );
and \U$56632 ( \57009 , \57008 , RIae7aa38_191);
nor \U$56633 ( \57010 , \57007 , \57009 );
xor \U$56634 ( \57011 , \57010 , \4251 );
and \U$56635 ( \57012 , \14964 , RIae788f0_120);
and \U$56636 ( \57013 , RIae78800_118, \14962 );
nor \U$56637 ( \57014 , \57012 , \57013 );
and \U$56638 ( \57015 , \57014 , \14463 );
not \U$56639 ( \57016 , \57014 );
and \U$56640 ( \57017 , \57016 , \14462 );
nor \U$56641 ( \57018 , \57015 , \57017 );
and \U$56642 ( \57019 , \57011 , \57018 );
and \U$56643 ( \57020 , \57010 , \4251 );
or \U$56644 ( \57021 , \57019 , \57020 );
xor \U$56645 ( \57022 , \57003 , \57021 );
and \U$56646 ( \57023 , \14059 , RIae77ea0_98);
and \U$56647 ( \57024 , RIae789e0_122, \14057 );
nor \U$56648 ( \57025 , \57023 , \57024 );
and \U$56649 ( \57026 , \57025 , \13502 );
not \U$56650 ( \57027 , \57025 );
and \U$56651 ( \57028 , \57027 , \14063 );
nor \U$56652 ( \57029 , \57026 , \57028 );
and \U$56653 ( \57030 , \12180 , RIae784b8_111);
and \U$56654 ( \57031 , RIae77cc0_94, \12178 );
nor \U$56655 ( \57032 , \57030 , \57031 );
and \U$56656 ( \57033 , \57032 , \12184 );
not \U$56657 ( \57034 , \57032 );
and \U$56658 ( \57035 , \57034 , \11827 );
nor \U$56659 ( \57036 , \57033 , \57035 );
xor \U$56660 ( \57037 , \57029 , \57036 );
and \U$56661 ( \57038 , \13059 , RIae77bd0_92);
and \U$56662 ( \57039 , RIae77db0_96, \13057 );
nor \U$56663 ( \57040 , \57038 , \57039 );
and \U$56664 ( \57041 , \57040 , \13063 );
not \U$56665 ( \57042 , \57040 );
and \U$56666 ( \57043 , \57042 , \12718 );
nor \U$56667 ( \57044 , \57041 , \57043 );
and \U$56668 ( \57045 , \57037 , \57044 );
and \U$56669 ( \57046 , \57029 , \57036 );
or \U$56670 ( \57047 , \57045 , \57046 );
and \U$56671 ( \57048 , \57022 , \57047 );
and \U$56672 ( \57049 , \57003 , \57021 );
or \U$56673 ( \57050 , \57048 , \57049 );
xor \U$56674 ( \57051 , \56978 , \57050 );
xor \U$56675 ( \57052 , \56706 , \56713 );
not \U$56676 ( \57053 , \57052 );
xor \U$56677 ( \57054 , \56750 , \56757 );
xor \U$56678 ( \57055 , \57054 , \56765 );
not \U$56679 ( \57056 , \57055 );
or \U$56680 ( \57057 , \57053 , \57056 );
or \U$56681 ( \57058 , \57055 , \57052 );
xor \U$56682 ( \57059 , \56722 , \56729 );
xor \U$56683 ( \57060 , \57059 , \56737 );
nand \U$56684 ( \57061 , \57058 , \57060 );
nand \U$56685 ( \57062 , \57057 , \57061 );
and \U$56686 ( \57063 , \57051 , \57062 );
and \U$56687 ( \57064 , \56978 , \57050 );
nor \U$56688 ( \57065 , \57063 , \57064 );
xor \U$56689 ( \57066 , \56826 , \56828 );
xor \U$56690 ( \57067 , \57066 , \56839 );
not \U$56691 ( \57068 , \57067 );
not \U$56692 ( \57069 , \56500 );
not \U$56693 ( \57070 , \56489 );
and \U$56694 ( \57071 , \57069 , \57070 );
and \U$56695 ( \57072 , \56500 , \56489 );
nor \U$56696 ( \57073 , \57071 , \57072 );
not \U$56697 ( \57074 , \57073 );
not \U$56698 ( \57075 , \3422 );
and \U$56699 ( \57076 , \57074 , \57075 );
and \U$56700 ( \57077 , \57073 , \3422 );
nor \U$56701 ( \57078 , \57076 , \57077 );
not \U$56702 ( \57079 , \57078 );
and \U$56703 ( \57080 , \57068 , \57079 );
and \U$56704 ( \57081 , \57067 , \57078 );
xor \U$56705 ( \57082 , \56679 , \56686 );
xor \U$56706 ( \57083 , \57082 , \56694 );
xor \U$56707 ( \57084 , \56650 , \56657 );
xor \U$56708 ( \57085 , \57084 , \56665 );
xor \U$56709 ( \57086 , \57083 , \57085 );
xor \U$56710 ( \57087 , \56625 , \56632 );
xor \U$56711 ( \57088 , \57087 , \56640 );
and \U$56712 ( \57089 , \57086 , \57088 );
and \U$56713 ( \57090 , \57083 , \57085 );
or \U$56714 ( \57091 , \57089 , \57090 );
nor \U$56715 ( \57092 , \57081 , \57091 );
nor \U$56716 ( \57093 , \57080 , \57092 );
xor \U$56717 ( \57094 , \57065 , \57093 );
not \U$56718 ( \57095 , \56697 );
not \U$56719 ( \57096 , \56668 );
or \U$56720 ( \57097 , \57095 , \57096 );
or \U$56721 ( \57098 , \56668 , \56697 );
nand \U$56722 ( \57099 , \57097 , \57098 );
not \U$56723 ( \57100 , \57099 );
not \U$56724 ( \57101 , \56643 );
and \U$56725 ( \57102 , \57100 , \57101 );
and \U$56726 ( \57103 , \57099 , \56643 );
nor \U$56727 ( \57104 , \57102 , \57103 );
xnor \U$56728 ( \57105 , \56768 , \56740 );
not \U$56729 ( \57106 , \57105 );
not \U$56730 ( \57107 , \56714 );
and \U$56731 ( \57108 , \57106 , \57107 );
and \U$56732 ( \57109 , \57105 , \56714 );
nor \U$56733 ( \57110 , \57108 , \57109 );
xor \U$56734 ( \57111 , \57104 , \57110 );
not \U$56735 ( \57112 , \56778 );
not \U$56736 ( \57113 , \56788 );
or \U$56737 ( \57114 , \57112 , \57113 );
or \U$56738 ( \57115 , \56788 , \56778 );
nand \U$56739 ( \57116 , \57114 , \57115 );
not \U$56740 ( \57117 , \57116 );
not \U$56741 ( \57118 , \56773 );
and \U$56742 ( \57119 , \57117 , \57118 );
and \U$56743 ( \57120 , \57116 , \56773 );
nor \U$56744 ( \57121 , \57119 , \57120 );
and \U$56745 ( \57122 , \57111 , \57121 );
and \U$56746 ( \57123 , \57104 , \57110 );
or \U$56747 ( \57124 , \57122 , \57123 );
and \U$56748 ( \57125 , \57094 , \57124 );
and \U$56749 ( \57126 , \57065 , \57093 );
nor \U$56750 ( \57127 , \57125 , \57126 );
not \U$56751 ( \57128 , \56806 );
not \U$56752 ( \57129 , \56803 );
or \U$56753 ( \57130 , \57128 , \57129 );
or \U$56754 ( \57131 , \56803 , \56806 );
nand \U$56755 ( \57132 , \57130 , \57131 );
not \U$56756 ( \57133 , \57132 );
xor \U$56757 ( \57134 , \56699 , \56770 );
xor \U$56758 ( \57135 , \57134 , \56790 );
not \U$56759 ( \57136 , \57135 );
or \U$56760 ( \57137 , \57133 , \57136 );
or \U$56761 ( \57138 , \57135 , \57132 );
not \U$56762 ( \57139 , \56818 );
xor \U$56763 ( \57140 , \56842 , \56821 );
not \U$56764 ( \57141 , \57140 );
or \U$56765 ( \57142 , \57139 , \57141 );
or \U$56766 ( \57143 , \57140 , \56818 );
nand \U$56767 ( \57144 , \57142 , \57143 );
nand \U$56768 ( \57145 , \57138 , \57144 );
nand \U$56769 ( \57146 , \57137 , \57145 );
xor \U$56770 ( \57147 , \57127 , \57146 );
xor \U$56771 ( \57148 , \56362 , \56364 );
xor \U$56772 ( \57149 , \57148 , \56371 );
xor \U$56773 ( \57150 , \56852 , \56857 );
xor \U$56774 ( \57151 , \57149 , \57150 );
and \U$56775 ( \57152 , \57147 , \57151 );
and \U$56776 ( \57153 , \57127 , \57146 );
or \U$56777 ( \57154 , \57152 , \57153 );
nand \U$56778 ( \57155 , \56897 , \57154 );
nand \U$56779 ( \57156 , \56894 , \57155 );
and \U$56780 ( \57157 , \56886 , \57156 );
xor \U$56781 ( \57158 , \57156 , \56886 );
not \U$56782 ( \57159 , \56888 );
not \U$56783 ( \57160 , \57154 );
and \U$56784 ( \57161 , \57159 , \57160 );
and \U$56785 ( \57162 , \56888 , \57154 );
nor \U$56786 ( \57163 , \57161 , \57162 );
xnor \U$56787 ( \57164 , \57163 , \56893 );
xor \U$56788 ( \57165 , \57127 , \57146 );
xor \U$56789 ( \57166 , \57165 , \57151 );
not \U$56790 ( \57167 , \57166 );
xor \U$56791 ( \57168 , \56793 , \56807 );
xor \U$56792 ( \57169 , \57168 , \56844 );
nand \U$56793 ( \57170 , \57167 , \57169 );
xor \U$56794 ( \57171 , \57065 , \57093 );
xor \U$56795 ( \57172 , \57171 , \57124 );
xnor \U$56796 ( \57173 , \57060 , \57055 );
not \U$56797 ( \57174 , \57173 );
not \U$56798 ( \57175 , \57052 );
and \U$56799 ( \57176 , \57174 , \57175 );
and \U$56800 ( \57177 , \57173 , \57052 );
nor \U$56801 ( \57178 , \57176 , \57177 );
not \U$56802 ( \57179 , \57178 );
xor \U$56803 ( \57180 , \56920 , \56947 );
xor \U$56804 ( \57181 , \57180 , \56975 );
not \U$56805 ( \57182 , \57181 );
and \U$56806 ( \57183 , \57179 , \57182 );
and \U$56807 ( \57184 , \57178 , \57181 );
xor \U$56808 ( \57185 , \57083 , \57085 );
xor \U$56809 ( \57186 , \57185 , \57088 );
nor \U$56810 ( \57187 , \57184 , \57186 );
nor \U$56811 ( \57188 , \57183 , \57187 );
not \U$56812 ( \57189 , \56927 );
xor \U$56813 ( \57190 , \56935 , \56945 );
not \U$56814 ( \57191 , \57190 );
or \U$56815 ( \57192 , \57189 , \57191 );
or \U$56816 ( \57193 , \57190 , \56927 );
nand \U$56817 ( \57194 , \57192 , \57193 );
not \U$56818 ( \57195 , \56955 );
xor \U$56819 ( \57196 , \56963 , \56973 );
not \U$56820 ( \57197 , \57196 );
or \U$56821 ( \57198 , \57195 , \57197 );
or \U$56822 ( \57199 , \57196 , \56955 );
nand \U$56823 ( \57200 , \57198 , \57199 );
xor \U$56824 ( \57201 , \57194 , \57200 );
xor \U$56825 ( \57202 , \56985 , \56992 );
xor \U$56826 ( \57203 , \57202 , \57000 );
and \U$56827 ( \57204 , \57201 , \57203 );
and \U$56828 ( \57205 , \57194 , \57200 );
or \U$56829 ( \57206 , \57204 , \57205 );
and \U$56830 ( \57207 , \11470 , RIae78260_106);
and \U$56831 ( \57208 , RIae78620_114, \11468 );
nor \U$56832 ( \57209 , \57207 , \57208 );
and \U$56833 ( \57210 , \57209 , \10936 );
not \U$56834 ( \57211 , \57209 );
and \U$56835 ( \57212 , \57211 , \11474 );
nor \U$56836 ( \57213 , \57210 , \57212 );
and \U$56837 ( \57214 , \12180 , RIae78440_110);
and \U$56838 ( \57215 , RIae784b8_111, \12178 );
nor \U$56839 ( \57216 , \57214 , \57215 );
and \U$56840 ( \57217 , \57216 , \12184 );
not \U$56841 ( \57218 , \57216 );
and \U$56842 ( \57219 , \57218 , \11827 );
nor \U$56843 ( \57220 , \57217 , \57219 );
xor \U$56844 ( \57221 , \57213 , \57220 );
and \U$56845 ( \57222 , \13059 , RIae77cc0_94);
and \U$56846 ( \57223 , RIae77bd0_92, \13057 );
nor \U$56847 ( \57224 , \57222 , \57223 );
and \U$56848 ( \57225 , \57224 , \13063 );
not \U$56849 ( \57226 , \57224 );
and \U$56850 ( \57227 , \57226 , \12718 );
nor \U$56851 ( \57228 , \57225 , \57227 );
and \U$56852 ( \57229 , \57221 , \57228 );
and \U$56853 ( \57230 , \57213 , \57220 );
or \U$56854 ( \57231 , \57229 , \57230 );
and \U$56855 ( \57232 , \14964 , RIae789e0_122);
and \U$56856 ( \57233 , RIae788f0_120, \14962 );
nor \U$56857 ( \57234 , \57232 , \57233 );
and \U$56858 ( \57235 , \57234 , \14463 );
not \U$56859 ( \57236 , \57234 );
and \U$56860 ( \57237 , \57236 , \14462 );
nor \U$56861 ( \57238 , \57235 , \57237 );
and \U$56862 ( \57239 , \15726 , RIae78800_118);
and \U$56863 ( \57240 , RIae78710_116, RIae7aab0_192);
nor \U$56864 ( \57241 , \57239 , \57240 );
and \U$56865 ( \57242 , \57241 , \14959 );
not \U$56866 ( \57243 , \57241 );
and \U$56867 ( \57244 , \57243 , RIae7aa38_191);
nor \U$56868 ( \57245 , \57242 , \57244 );
xor \U$56869 ( \57246 , \57238 , \57245 );
and \U$56870 ( \57247 , \14059 , RIae77db0_96);
and \U$56871 ( \57248 , RIae77ea0_98, \14057 );
nor \U$56872 ( \57249 , \57247 , \57248 );
and \U$56873 ( \57250 , \57249 , \13502 );
not \U$56874 ( \57251 , \57249 );
and \U$56875 ( \57252 , \57251 , \14063 );
nor \U$56876 ( \57253 , \57250 , \57252 );
and \U$56877 ( \57254 , \57246 , \57253 );
and \U$56878 ( \57255 , \57238 , \57245 );
or \U$56879 ( \57256 , \57254 , \57255 );
xor \U$56880 ( \57257 , \57231 , \57256 );
and \U$56881 ( \57258 , \8966 , RIae77270_72);
and \U$56882 ( \57259 , RIae77360_74, \8964 );
nor \U$56883 ( \57260 , \57258 , \57259 );
and \U$56884 ( \57261 , \57260 , \8799 );
not \U$56885 ( \57262 , \57260 );
and \U$56886 ( \57263 , \57262 , \8789 );
nor \U$56887 ( \57264 , \57261 , \57263 );
and \U$56888 ( \57265 , \9760 , RIae78350_108);
and \U$56889 ( \57266 , RIae78170_104, \9758 );
nor \U$56890 ( \57267 , \57265 , \57266 );
and \U$56891 ( \57268 , \57267 , \9273 );
not \U$56892 ( \57269 , \57267 );
and \U$56893 ( \57270 , \57269 , \9764 );
nor \U$56894 ( \57271 , \57268 , \57270 );
xor \U$56895 ( \57272 , \57264 , \57271 );
and \U$56896 ( \57273 , \10548 , RIae77f90_100);
and \U$56897 ( \57274 , RIae78080_102, \10546 );
nor \U$56898 ( \57275 , \57273 , \57274 );
and \U$56899 ( \57276 , \57275 , \10421 );
not \U$56900 ( \57277 , \57275 );
and \U$56901 ( \57278 , \57277 , \10118 );
nor \U$56902 ( \57279 , \57276 , \57278 );
and \U$56903 ( \57280 , \57272 , \57279 );
and \U$56904 ( \57281 , \57264 , \57271 );
or \U$56905 ( \57282 , \57280 , \57281 );
and \U$56906 ( \57283 , \57257 , \57282 );
and \U$56907 ( \57284 , \57231 , \57256 );
or \U$56908 ( \57285 , \57283 , \57284 );
xor \U$56909 ( \57286 , \57206 , \57285 );
xor \U$56910 ( \57287 , \56904 , \56909 );
xor \U$56911 ( \57288 , \57287 , \56917 );
and \U$56912 ( \57289 , \7633 , RIae76dc0_62);
and \U$56913 ( \57290 , RIae76cd0_60, \7631 );
nor \U$56914 ( \57291 , \57289 , \57290 );
and \U$56915 ( \57292 , \57291 , \7206 );
not \U$56916 ( \57293 , \57291 );
and \U$56917 ( \57294 , \57293 , \7205 );
nor \U$56918 ( \57295 , \57292 , \57294 );
and \U$56919 ( \57296 , \8371 , RIae77108_69);
and \U$56920 ( \57297 , RIae77090_68, \8369 );
nor \U$56921 ( \57298 , \57296 , \57297 );
and \U$56922 ( \57299 , \57298 , \8020 );
not \U$56923 ( \57300 , \57298 );
and \U$56924 ( \57301 , \57300 , \8019 );
nor \U$56925 ( \57302 , \57299 , \57301 );
xor \U$56926 ( \57303 , \57295 , \57302 );
and \U$56927 ( \57304 , \6941 , RIae76fa0_66);
and \U$56928 ( \57305 , RIae76eb0_64, \6939 );
nor \U$56929 ( \57306 , \57304 , \57305 );
and \U$56930 ( \57307 , \57306 , \6314 );
not \U$56931 ( \57308 , \57306 );
and \U$56932 ( \57309 , \57308 , \6945 );
nor \U$56933 ( \57310 , \57307 , \57309 );
and \U$56934 ( \57311 , \57303 , \57310 );
and \U$56935 ( \57312 , \57295 , \57302 );
nor \U$56936 ( \57313 , \57311 , \57312 );
or \U$56937 ( \57314 , \57288 , \57313 );
not \U$56938 ( \57315 , \57313 );
not \U$56939 ( \57316 , \57288 );
or \U$56940 ( \57317 , \57315 , \57316 );
and \U$56941 ( \57318 , \5399 , RIae776a8_81);
and \U$56942 ( \57319 , RIae77450_76, \5397 );
nor \U$56943 ( \57320 , \57318 , \57319 );
and \U$56944 ( \57321 , \57320 , \5016 );
not \U$56945 ( \57322 , \57320 );
and \U$56946 ( \57323 , \57322 , \5403 );
nor \U$56947 ( \57324 , \57321 , \57323 );
and \U$56948 ( \57325 , \5896 , RIae77ae0_90);
and \U$56949 ( \57326 , RIae779f0_88, \5894 );
nor \U$56950 ( \57327 , \57325 , \57326 );
and \U$56951 ( \57328 , \57327 , \5590 );
not \U$56952 ( \57329 , \57327 );
and \U$56953 ( \57330 , \57329 , \5589 );
nor \U$56954 ( \57331 , \57328 , \57330 );
xor \U$56955 ( \57332 , \57324 , \57331 );
and \U$56956 ( \57333 , \6172 , RIae77810_84);
and \U$56957 ( \57334 , RIae77900_86, \6170 );
nor \U$56958 ( \57335 , \57333 , \57334 );
and \U$56959 ( \57336 , \57335 , \6176 );
not \U$56960 ( \57337 , \57335 );
and \U$56961 ( \57338 , \57337 , \6175 );
nor \U$56962 ( \57339 , \57336 , \57338 );
and \U$56963 ( \57340 , \57332 , \57339 );
and \U$56964 ( \57341 , \57324 , \57331 );
or \U$56965 ( \57342 , \57340 , \57341 );
nand \U$56966 ( \57343 , \57317 , \57342 );
nand \U$56967 ( \57344 , \57314 , \57343 );
and \U$56968 ( \57345 , \57286 , \57344 );
and \U$56969 ( \57346 , \57206 , \57285 );
nor \U$56970 ( \57347 , \57345 , \57346 );
xor \U$56971 ( \57348 , \57188 , \57347 );
xor \U$56972 ( \57349 , \57104 , \57110 );
xor \U$56973 ( \57350 , \57349 , \57121 );
and \U$56974 ( \57351 , \57348 , \57350 );
and \U$56975 ( \57352 , \57188 , \57347 );
or \U$56976 ( \57353 , \57351 , \57352 );
xor \U$56977 ( \57354 , \57172 , \57353 );
xnor \U$56978 ( \57355 , \57135 , \57144 );
not \U$56979 ( \57356 , \57355 );
not \U$56980 ( \57357 , \57132 );
and \U$56981 ( \57358 , \57356 , \57357 );
and \U$56982 ( \57359 , \57355 , \57132 );
nor \U$56983 ( \57360 , \57358 , \57359 );
and \U$56984 ( \57361 , \57354 , \57360 );
and \U$56985 ( \57362 , \57172 , \57353 );
nor \U$56986 ( \57363 , \57361 , \57362 );
and \U$56987 ( \57364 , \57170 , \57363 );
not \U$56988 ( \57365 , \57169 );
and \U$56989 ( \57366 , \57365 , \57166 );
nor \U$56990 ( \57367 , \57364 , \57366 );
or \U$56991 ( \57368 , \57164 , \57367 );
xnor \U$56992 ( \57369 , \57367 , \57164 );
not \U$56993 ( \57370 , \57166 );
not \U$56994 ( \57371 , \57363 );
not \U$56995 ( \57372 , \57169 );
and \U$56996 ( \57373 , \57371 , \57372 );
and \U$56997 ( \57374 , \57363 , \57169 );
nor \U$56998 ( \57375 , \57373 , \57374 );
not \U$56999 ( \57376 , \57375 );
or \U$57000 ( \57377 , \57370 , \57376 );
or \U$57001 ( \57378 , \57375 , \57166 );
nand \U$57002 ( \57379 , \57377 , \57378 );
xor \U$57003 ( \57380 , \57172 , \57353 );
xor \U$57004 ( \57381 , \57380 , \57360 );
xor \U$57005 ( \57382 , \57188 , \57347 );
xor \U$57006 ( \57383 , \57382 , \57350 );
not \U$57007 ( \57384 , \57383 );
xor \U$57008 ( \57385 , \56978 , \57050 );
xor \U$57009 ( \57386 , \57385 , \57062 );
nand \U$57010 ( \57387 , \57384 , \57386 );
or \U$57011 ( \57388 , \57381 , \57387 );
not \U$57012 ( \57389 , \57387 );
not \U$57013 ( \57390 , \57381 );
or \U$57014 ( \57391 , \57389 , \57390 );
xor \U$57015 ( \57392 , \57029 , \57036 );
xor \U$57016 ( \57393 , \57392 , \57044 );
xor \U$57017 ( \57394 , \57010 , \4251 );
xor \U$57018 ( \57395 , \57394 , \57018 );
and \U$57019 ( \57396 , \57393 , \57395 );
xor \U$57020 ( \57397 , \57194 , \57200 );
xor \U$57021 ( \57398 , \57397 , \57203 );
xor \U$57022 ( \57399 , \57010 , \4251 );
xor \U$57023 ( \57400 , \57399 , \57018 );
and \U$57024 ( \57401 , \57398 , \57400 );
and \U$57025 ( \57402 , \57393 , \57398 );
or \U$57026 ( \57403 , \57396 , \57401 , \57402 );
not \U$57027 ( \57404 , \57403 );
not \U$57028 ( \57405 , \57342 );
not \U$57029 ( \57406 , \57313 );
or \U$57030 ( \57407 , \57405 , \57406 );
or \U$57031 ( \57408 , \57313 , \57342 );
nand \U$57032 ( \57409 , \57407 , \57408 );
not \U$57033 ( \57410 , \57409 );
not \U$57034 ( \57411 , \57288 );
and \U$57035 ( \57412 , \57410 , \57411 );
and \U$57036 ( \57413 , \57409 , \57288 );
nor \U$57037 ( \57414 , \57412 , \57413 );
not \U$57038 ( \57415 , \57414 );
xor \U$57039 ( \57416 , \57231 , \57256 );
xor \U$57040 ( \57417 , \57416 , \57282 );
nand \U$57041 ( \57418 , \57415 , \57417 );
or \U$57042 ( \57419 , \57404 , \57418 );
and \U$57043 ( \57420 , \57404 , \57418 );
and \U$57044 ( \57421 , \11470 , RIae78080_102);
and \U$57045 ( \57422 , RIae78260_106, \11468 );
nor \U$57046 ( \57423 , \57421 , \57422 );
and \U$57047 ( \57424 , \57423 , \10936 );
not \U$57048 ( \57425 , \57423 );
and \U$57049 ( \57426 , \57425 , \11474 );
nor \U$57050 ( \57427 , \57424 , \57426 );
and \U$57051 ( \57428 , \9760 , RIae77360_74);
and \U$57052 ( \57429 , RIae78350_108, \9758 );
nor \U$57053 ( \57430 , \57428 , \57429 );
and \U$57054 ( \57431 , \57430 , \9273 );
not \U$57055 ( \57432 , \57430 );
and \U$57056 ( \57433 , \57432 , \9272 );
nor \U$57057 ( \57434 , \57431 , \57433 );
xor \U$57058 ( \57435 , \57427 , \57434 );
and \U$57059 ( \57436 , \10548 , RIae78170_104);
and \U$57060 ( \57437 , RIae77f90_100, \10546 );
nor \U$57061 ( \57438 , \57436 , \57437 );
and \U$57062 ( \57439 , \57438 , \10421 );
not \U$57063 ( \57440 , \57438 );
and \U$57064 ( \57441 , \57440 , \10118 );
nor \U$57065 ( \57442 , \57439 , \57441 );
and \U$57066 ( \57443 , \57435 , \57442 );
and \U$57067 ( \57444 , \57427 , \57434 );
or \U$57068 ( \57445 , \57443 , \57444 );
and \U$57069 ( \57446 , \15726 , RIae788f0_120);
and \U$57070 ( \57447 , RIae78800_118, RIae7aab0_192);
nor \U$57071 ( \57448 , \57446 , \57447 );
and \U$57072 ( \57449 , \57448 , \14959 );
not \U$57073 ( \57450 , \57448 );
and \U$57074 ( \57451 , \57450 , RIae7aa38_191);
nor \U$57075 ( \57452 , \57449 , \57451 );
xor \U$57076 ( \57453 , \57452 , \4482 );
and \U$57077 ( \57454 , \14964 , RIae77ea0_98);
and \U$57078 ( \57455 , RIae789e0_122, \14962 );
nor \U$57079 ( \57456 , \57454 , \57455 );
and \U$57080 ( \57457 , \57456 , \14463 );
not \U$57081 ( \57458 , \57456 );
and \U$57082 ( \57459 , \57458 , \14462 );
nor \U$57083 ( \57460 , \57457 , \57459 );
and \U$57084 ( \57461 , \57453 , \57460 );
and \U$57085 ( \57462 , \57452 , \4482 );
or \U$57086 ( \57463 , \57461 , \57462 );
xor \U$57087 ( \57464 , \57445 , \57463 );
and \U$57088 ( \57465 , \12180 , RIae78620_114);
and \U$57089 ( \57466 , RIae78440_110, \12178 );
nor \U$57090 ( \57467 , \57465 , \57466 );
and \U$57091 ( \57468 , \57467 , \12184 );
not \U$57092 ( \57469 , \57467 );
and \U$57093 ( \57470 , \57469 , \11827 );
nor \U$57094 ( \57471 , \57468 , \57470 );
and \U$57095 ( \57472 , \13059 , RIae784b8_111);
and \U$57096 ( \57473 , RIae77cc0_94, \13057 );
nor \U$57097 ( \57474 , \57472 , \57473 );
and \U$57098 ( \57475 , \57474 , \13063 );
not \U$57099 ( \57476 , \57474 );
and \U$57100 ( \57477 , \57476 , \12718 );
nor \U$57101 ( \57478 , \57475 , \57477 );
xor \U$57102 ( \57479 , \57471 , \57478 );
and \U$57103 ( \57480 , \14059 , RIae77bd0_92);
and \U$57104 ( \57481 , RIae77db0_96, \14057 );
nor \U$57105 ( \57482 , \57480 , \57481 );
and \U$57106 ( \57483 , \57482 , \13502 );
not \U$57107 ( \57484 , \57482 );
and \U$57108 ( \57485 , \57484 , \14063 );
nor \U$57109 ( \57486 , \57483 , \57485 );
and \U$57110 ( \57487 , \57479 , \57486 );
and \U$57111 ( \57488 , \57471 , \57478 );
or \U$57112 ( \57489 , \57487 , \57488 );
and \U$57113 ( \57490 , \57464 , \57489 );
and \U$57114 ( \57491 , \57445 , \57463 );
or \U$57115 ( \57492 , \57490 , \57491 );
and \U$57116 ( \57493 , \5896 , RIae77450_76);
and \U$57117 ( \57494 , RIae77ae0_90, \5894 );
nor \U$57118 ( \57495 , \57493 , \57494 );
and \U$57119 ( \57496 , \57495 , \5590 );
not \U$57120 ( \57497 , \57495 );
and \U$57121 ( \57498 , \57497 , \5589 );
nor \U$57122 ( \57499 , \57496 , \57498 );
and \U$57123 ( \57500 , \6172 , RIae779f0_88);
and \U$57124 ( \57501 , RIae77810_84, \6170 );
nor \U$57125 ( \57502 , \57500 , \57501 );
and \U$57126 ( \57503 , \57502 , \6176 );
not \U$57127 ( \57504 , \57502 );
and \U$57128 ( \57505 , \57504 , \6175 );
nor \U$57129 ( \57506 , \57503 , \57505 );
xor \U$57130 ( \57507 , \57499 , \57506 );
and \U$57131 ( \57508 , \6941 , RIae77900_86);
and \U$57132 ( \57509 , RIae76fa0_66, \6939 );
nor \U$57133 ( \57510 , \57508 , \57509 );
and \U$57134 ( \57511 , \57510 , \6314 );
not \U$57135 ( \57512 , \57510 );
and \U$57136 ( \57513 , \57512 , \6945 );
nor \U$57137 ( \57514 , \57511 , \57513 );
and \U$57138 ( \57515 , \57507 , \57514 );
and \U$57139 ( \57516 , \57499 , \57506 );
or \U$57140 ( \57517 , \57515 , \57516 );
and \U$57141 ( \57518 , \4688 , RIae77630_80);
and \U$57142 ( \57519 , RIae77540_78, \4686 );
nor \U$57143 ( \57520 , \57518 , \57519 );
and \U$57144 ( \57521 , \57520 , \4481 );
not \U$57145 ( \57522 , \57520 );
and \U$57146 ( \57523 , \57522 , \4482 );
nor \U$57147 ( \57524 , \57521 , \57523 );
xor \U$57148 ( \57525 , \57517 , \57524 );
and \U$57149 ( \57526 , \8966 , RIae77090_68);
and \U$57150 ( \57527 , RIae77270_72, \8964 );
nor \U$57151 ( \57528 , \57526 , \57527 );
and \U$57152 ( \57529 , \57528 , \8799 );
not \U$57153 ( \57530 , \57528 );
and \U$57154 ( \57531 , \57530 , \8789 );
nor \U$57155 ( \57532 , \57529 , \57531 );
and \U$57156 ( \57533 , \7633 , RIae76eb0_64);
and \U$57157 ( \57534 , RIae76dc0_62, \7631 );
nor \U$57158 ( \57535 , \57533 , \57534 );
and \U$57159 ( \57536 , \57535 , \7206 );
not \U$57160 ( \57537 , \57535 );
and \U$57161 ( \57538 , \57537 , \7205 );
nor \U$57162 ( \57539 , \57536 , \57538 );
xor \U$57163 ( \57540 , \57532 , \57539 );
and \U$57164 ( \57541 , \8371 , RIae76cd0_60);
and \U$57165 ( \57542 , RIae77108_69, \8369 );
nor \U$57166 ( \57543 , \57541 , \57542 );
and \U$57167 ( \57544 , \57543 , \8020 );
not \U$57168 ( \57545 , \57543 );
and \U$57169 ( \57546 , \57545 , \8019 );
nor \U$57170 ( \57547 , \57544 , \57546 );
and \U$57171 ( \57548 , \57540 , \57547 );
and \U$57172 ( \57549 , \57532 , \57539 );
or \U$57173 ( \57550 , \57548 , \57549 );
and \U$57174 ( \57551 , \57525 , \57550 );
and \U$57175 ( \57552 , \57517 , \57524 );
or \U$57176 ( \57553 , \57551 , \57552 );
xor \U$57177 ( \57554 , \57492 , \57553 );
xor \U$57178 ( \57555 , \57324 , \57331 );
xor \U$57179 ( \57556 , \57555 , \57339 );
xor \U$57180 ( \57557 , \57264 , \57271 );
xor \U$57181 ( \57558 , \57557 , \57279 );
and \U$57182 ( \57559 , \57556 , \57558 );
xor \U$57183 ( \57560 , \57295 , \57302 );
xor \U$57184 ( \57561 , \57560 , \57310 );
xor \U$57185 ( \57562 , \57264 , \57271 );
xor \U$57186 ( \57563 , \57562 , \57279 );
and \U$57187 ( \57564 , \57561 , \57563 );
and \U$57188 ( \57565 , \57556 , \57561 );
or \U$57189 ( \57566 , \57559 , \57564 , \57565 );
and \U$57190 ( \57567 , \57554 , \57566 );
and \U$57191 ( \57568 , \57492 , \57553 );
nor \U$57192 ( \57569 , \57567 , \57568 );
nor \U$57193 ( \57570 , \57420 , \57569 );
not \U$57194 ( \57571 , \57570 );
nand \U$57195 ( \57572 , \57419 , \57571 );
not \U$57196 ( \57573 , \57067 );
xor \U$57197 ( \57574 , \57078 , \57091 );
not \U$57198 ( \57575 , \57574 );
or \U$57199 ( \57576 , \57573 , \57575 );
or \U$57200 ( \57577 , \57574 , \57067 );
nand \U$57201 ( \57578 , \57576 , \57577 );
xor \U$57202 ( \57579 , \57572 , \57578 );
xor \U$57203 ( \57580 , \57206 , \57285 );
xor \U$57204 ( \57581 , \57580 , \57344 );
xor \U$57205 ( \57582 , \57003 , \57021 );
xor \U$57206 ( \57583 , \57582 , \57047 );
xor \U$57207 ( \57584 , \57581 , \57583 );
not \U$57208 ( \57585 , \57178 );
xor \U$57209 ( \57586 , \57181 , \57186 );
not \U$57210 ( \57587 , \57586 );
or \U$57211 ( \57588 , \57585 , \57587 );
or \U$57212 ( \57589 , \57586 , \57178 );
nand \U$57213 ( \57590 , \57588 , \57589 );
and \U$57214 ( \57591 , \57584 , \57590 );
and \U$57215 ( \57592 , \57581 , \57583 );
or \U$57216 ( \57593 , \57591 , \57592 );
and \U$57217 ( \57594 , \57579 , \57593 );
and \U$57218 ( \57595 , \57572 , \57578 );
or \U$57219 ( \57596 , \57594 , \57595 );
nand \U$57220 ( \57597 , \57391 , \57596 );
nand \U$57221 ( \57598 , \57388 , \57597 );
and \U$57222 ( \57599 , \57379 , \57598 );
xor \U$57223 ( \57600 , \57598 , \57379 );
not \U$57224 ( \57601 , \57386 );
not \U$57225 ( \57602 , \57383 );
or \U$57226 ( \57603 , \57601 , \57602 );
or \U$57227 ( \57604 , \57383 , \57386 );
nand \U$57228 ( \57605 , \57603 , \57604 );
xor \U$57229 ( \57606 , \57010 , \4251 );
xor \U$57230 ( \57607 , \57606 , \57018 );
xor \U$57231 ( \57608 , \57393 , \57398 );
xor \U$57232 ( \57609 , \57607 , \57608 );
not \U$57233 ( \57610 , \57414 );
not \U$57234 ( \57611 , \57417 );
or \U$57235 ( \57612 , \57610 , \57611 );
or \U$57236 ( \57613 , \57417 , \57414 );
nand \U$57237 ( \57614 , \57612 , \57613 );
xor \U$57238 ( \57615 , \57609 , \57614 );
xor \U$57239 ( \57616 , \57492 , \57553 );
xor \U$57240 ( \57617 , \57616 , \57566 );
and \U$57241 ( \57618 , \57615 , \57617 );
and \U$57242 ( \57619 , \57609 , \57614 );
or \U$57243 ( \57620 , \57618 , \57619 );
not \U$57244 ( \57621 , \57620 );
xor \U$57245 ( \57622 , \57581 , \57583 );
xor \U$57246 ( \57623 , \57622 , \57590 );
not \U$57247 ( \57624 , \57623 );
or \U$57248 ( \57625 , \57621 , \57624 );
or \U$57249 ( \57626 , \57623 , \57620 );
and \U$57250 ( \57627 , \9760 , RIae77270_72);
and \U$57251 ( \57628 , RIae77360_74, \9758 );
nor \U$57252 ( \57629 , \57627 , \57628 );
and \U$57253 ( \57630 , \57629 , \9273 );
not \U$57254 ( \57631 , \57629 );
and \U$57255 ( \57632 , \57631 , \9764 );
nor \U$57256 ( \57633 , \57630 , \57632 );
and \U$57257 ( \57634 , \10548 , RIae78350_108);
and \U$57258 ( \57635 , RIae78170_104, \10546 );
nor \U$57259 ( \57636 , \57634 , \57635 );
and \U$57260 ( \57637 , \57636 , \10421 );
not \U$57261 ( \57638 , \57636 );
and \U$57262 ( \57639 , \57638 , \10118 );
nor \U$57263 ( \57640 , \57637 , \57639 );
xor \U$57264 ( \57641 , \57633 , \57640 );
and \U$57265 ( \57642 , \8966 , RIae77108_69);
and \U$57266 ( \57643 , RIae77090_68, \8964 );
nor \U$57267 ( \57644 , \57642 , \57643 );
and \U$57268 ( \57645 , \57644 , \8799 );
not \U$57269 ( \57646 , \57644 );
and \U$57270 ( \57647 , \57646 , \8789 );
nor \U$57271 ( \57648 , \57645 , \57647 );
and \U$57272 ( \57649 , \57641 , \57648 );
and \U$57273 ( \57650 , \57633 , \57640 );
nor \U$57274 ( \57651 , \57649 , \57650 );
and \U$57275 ( \57652 , \11470 , RIae77f90_100);
and \U$57276 ( \57653 , RIae78080_102, \11468 );
nor \U$57277 ( \57654 , \57652 , \57653 );
and \U$57278 ( \57655 , \57654 , \11474 );
not \U$57279 ( \57656 , \57654 );
and \U$57280 ( \57657 , \57656 , \10936 );
nor \U$57281 ( \57658 , \57655 , \57657 );
and \U$57282 ( \57659 , \12180 , RIae78260_106);
and \U$57283 ( \57660 , RIae78620_114, \12178 );
nor \U$57284 ( \57661 , \57659 , \57660 );
and \U$57285 ( \57662 , \57661 , \11827 );
not \U$57286 ( \57663 , \57661 );
and \U$57287 ( \57664 , \57663 , \12184 );
nor \U$57288 ( \57665 , \57662 , \57664 );
xor \U$57289 ( \57666 , \57658 , \57665 );
and \U$57290 ( \57667 , \13059 , RIae78440_110);
and \U$57291 ( \57668 , RIae784b8_111, \13057 );
nor \U$57292 ( \57669 , \57667 , \57668 );
and \U$57293 ( \57670 , \57669 , \12718 );
not \U$57294 ( \57671 , \57669 );
and \U$57295 ( \57672 , \57671 , \13063 );
nor \U$57296 ( \57673 , \57670 , \57672 );
and \U$57297 ( \57674 , \57666 , \57673 );
and \U$57298 ( \57675 , \57658 , \57665 );
or \U$57299 ( \57676 , \57674 , \57675 );
xor \U$57300 ( \57677 , \57651 , \57676 );
and \U$57301 ( \57678 , \14059 , RIae77cc0_94);
and \U$57302 ( \57679 , RIae77bd0_92, \14057 );
nor \U$57303 ( \57680 , \57678 , \57679 );
and \U$57304 ( \57681 , \57680 , \14063 );
not \U$57305 ( \57682 , \57680 );
and \U$57306 ( \57683 , \57682 , \13502 );
nor \U$57307 ( \57684 , \57681 , \57683 );
and \U$57308 ( \57685 , \15726 , RIae789e0_122);
and \U$57309 ( \57686 , RIae788f0_120, RIae7aab0_192);
nor \U$57310 ( \57687 , \57685 , \57686 );
and \U$57311 ( \57688 , \57687 , RIae7aa38_191);
not \U$57312 ( \57689 , \57687 );
and \U$57313 ( \57690 , \57689 , \14959 );
nor \U$57314 ( \57691 , \57688 , \57690 );
xor \U$57315 ( \57692 , \57684 , \57691 );
and \U$57316 ( \57693 , \14964 , RIae77db0_96);
and \U$57317 ( \57694 , RIae77ea0_98, \14962 );
nor \U$57318 ( \57695 , \57693 , \57694 );
and \U$57319 ( \57696 , \57695 , \14462 );
not \U$57320 ( \57697 , \57695 );
and \U$57321 ( \57698 , \57697 , \14463 );
nor \U$57322 ( \57699 , \57696 , \57698 );
and \U$57323 ( \57700 , \57692 , \57699 );
and \U$57324 ( \57701 , \57684 , \57691 );
or \U$57325 ( \57702 , \57700 , \57701 );
and \U$57326 ( \57703 , \57677 , \57702 );
and \U$57327 ( \57704 , \57651 , \57676 );
nor \U$57328 ( \57705 , \57703 , \57704 );
and \U$57329 ( \57706 , \6941 , RIae77810_84);
and \U$57330 ( \57707 , RIae77900_86, \6939 );
nor \U$57331 ( \57708 , \57706 , \57707 );
and \U$57332 ( \57709 , \57708 , \6945 );
not \U$57333 ( \57710 , \57708 );
and \U$57334 ( \57711 , \57710 , \6314 );
nor \U$57335 ( \57712 , \57709 , \57711 );
and \U$57336 ( \57713 , \8371 , RIae76dc0_62);
and \U$57337 ( \57714 , RIae76cd0_60, \8369 );
nor \U$57338 ( \57715 , \57713 , \57714 );
and \U$57339 ( \57716 , \57715 , \8019 );
not \U$57340 ( \57717 , \57715 );
and \U$57341 ( \57718 , \57717 , \8020 );
nor \U$57342 ( \57719 , \57716 , \57718 );
or \U$57343 ( \57720 , \57712 , \57719 );
not \U$57344 ( \57721 , \57719 );
not \U$57345 ( \57722 , \57712 );
or \U$57346 ( \57723 , \57721 , \57722 );
and \U$57347 ( \57724 , \7633 , RIae76fa0_66);
and \U$57348 ( \57725 , RIae76eb0_64, \7631 );
nor \U$57349 ( \57726 , \57724 , \57725 );
and \U$57350 ( \57727 , \57726 , \7206 );
not \U$57351 ( \57728 , \57726 );
and \U$57352 ( \57729 , \57728 , \7205 );
nor \U$57353 ( \57730 , \57727 , \57729 );
nand \U$57354 ( \57731 , \57723 , \57730 );
nand \U$57355 ( \57732 , \57720 , \57731 );
and \U$57356 ( \57733 , \5399 , RIae77540_78);
and \U$57357 ( \57734 , RIae776a8_81, \5397 );
nor \U$57358 ( \57735 , \57733 , \57734 );
and \U$57359 ( \57736 , \57735 , \5016 );
not \U$57360 ( \57737 , \57735 );
and \U$57361 ( \57738 , \57737 , \5403 );
nor \U$57362 ( \57739 , \57736 , \57738 );
xor \U$57363 ( \57740 , \57732 , \57739 );
and \U$57364 ( \57741 , \5399 , RIae77630_80);
and \U$57365 ( \57742 , RIae77540_78, \5397 );
nor \U$57366 ( \57743 , \57741 , \57742 );
and \U$57367 ( \57744 , \57743 , \5403 );
not \U$57368 ( \57745 , \57743 );
and \U$57369 ( \57746 , \57745 , \5016 );
nor \U$57370 ( \57747 , \57744 , \57746 );
and \U$57371 ( \57748 , \5896 , RIae776a8_81);
and \U$57372 ( \57749 , RIae77450_76, \5894 );
nor \U$57373 ( \57750 , \57748 , \57749 );
and \U$57374 ( \57751 , \57750 , \5589 );
not \U$57375 ( \57752 , \57750 );
and \U$57376 ( \57753 , \57752 , \5590 );
nor \U$57377 ( \57754 , \57751 , \57753 );
or \U$57378 ( \57755 , \57747 , \57754 );
not \U$57379 ( \57756 , \57754 );
not \U$57380 ( \57757 , \57747 );
or \U$57381 ( \57758 , \57756 , \57757 );
and \U$57382 ( \57759 , \6172 , RIae77ae0_90);
and \U$57383 ( \57760 , RIae779f0_88, \6170 );
nor \U$57384 ( \57761 , \57759 , \57760 );
and \U$57385 ( \57762 , \57761 , \6176 );
not \U$57386 ( \57763 , \57761 );
and \U$57387 ( \57764 , \57763 , \6175 );
nor \U$57388 ( \57765 , \57762 , \57764 );
nand \U$57389 ( \57766 , \57758 , \57765 );
nand \U$57390 ( \57767 , \57755 , \57766 );
and \U$57391 ( \57768 , \57740 , \57767 );
and \U$57392 ( \57769 , \57732 , \57739 );
or \U$57393 ( \57770 , \57768 , \57769 );
xor \U$57394 ( \57771 , \57705 , \57770 );
nand \U$57395 ( \57772 , RIae77630_80, \4686 );
and \U$57396 ( \57773 , \57772 , \4481 );
not \U$57397 ( \57774 , \57772 );
and \U$57398 ( \57775 , \57774 , \4482 );
nor \U$57399 ( \57776 , \57773 , \57775 );
xor \U$57400 ( \57777 , \57499 , \57506 );
xor \U$57401 ( \57778 , \57777 , \57514 );
and \U$57402 ( \57779 , \57776 , \57778 );
xor \U$57403 ( \57780 , \57532 , \57539 );
xor \U$57404 ( \57781 , \57780 , \57547 );
xor \U$57405 ( \57782 , \57499 , \57506 );
xor \U$57406 ( \57783 , \57782 , \57514 );
and \U$57407 ( \57784 , \57781 , \57783 );
and \U$57408 ( \57785 , \57776 , \57781 );
or \U$57409 ( \57786 , \57779 , \57784 , \57785 );
and \U$57410 ( \57787 , \57771 , \57786 );
and \U$57411 ( \57788 , \57705 , \57770 );
or \U$57412 ( \57789 , \57787 , \57788 );
xor \U$57413 ( \57790 , \57238 , \57245 );
xor \U$57414 ( \57791 , \57790 , \57253 );
xor \U$57415 ( \57792 , \57213 , \57220 );
xor \U$57416 ( \57793 , \57792 , \57228 );
and \U$57417 ( \57794 , \57791 , \57793 );
xor \U$57418 ( \57795 , \57427 , \57434 );
xor \U$57419 ( \57796 , \57795 , \57442 );
xor \U$57420 ( \57797 , \57471 , \57478 );
xor \U$57421 ( \57798 , \57797 , \57486 );
xor \U$57422 ( \57799 , \57796 , \57798 );
xor \U$57423 ( \57800 , \57452 , \4482 );
xor \U$57424 ( \57801 , \57800 , \57460 );
and \U$57425 ( \57802 , \57799 , \57801 );
and \U$57426 ( \57803 , \57796 , \57798 );
or \U$57427 ( \57804 , \57802 , \57803 );
xor \U$57428 ( \57805 , \57213 , \57220 );
xor \U$57429 ( \57806 , \57805 , \57228 );
and \U$57430 ( \57807 , \57804 , \57806 );
and \U$57431 ( \57808 , \57791 , \57804 );
or \U$57432 ( \57809 , \57794 , \57807 , \57808 );
xor \U$57433 ( \57810 , \57789 , \57809 );
xor \U$57434 ( \57811 , \57517 , \57524 );
xor \U$57435 ( \57812 , \57811 , \57550 );
xor \U$57436 ( \57813 , \57445 , \57463 );
xor \U$57437 ( \57814 , \57813 , \57489 );
and \U$57438 ( \57815 , \57812 , \57814 );
xor \U$57439 ( \57816 , \57264 , \57271 );
xor \U$57440 ( \57817 , \57816 , \57279 );
xor \U$57441 ( \57818 , \57556 , \57561 );
xor \U$57442 ( \57819 , \57817 , \57818 );
xor \U$57443 ( \57820 , \57445 , \57463 );
xor \U$57444 ( \57821 , \57820 , \57489 );
and \U$57445 ( \57822 , \57819 , \57821 );
and \U$57446 ( \57823 , \57812 , \57819 );
or \U$57447 ( \57824 , \57815 , \57822 , \57823 );
and \U$57448 ( \57825 , \57810 , \57824 );
and \U$57449 ( \57826 , \57789 , \57809 );
or \U$57450 ( \57827 , \57825 , \57826 );
nand \U$57451 ( \57828 , \57626 , \57827 );
nand \U$57452 ( \57829 , \57625 , \57828 );
xor \U$57453 ( \57830 , \57605 , \57829 );
xor \U$57454 ( \57831 , \57572 , \57578 );
xor \U$57455 ( \57832 , \57831 , \57593 );
xor \U$57456 ( \57833 , \57830 , \57832 );
xnor \U$57457 ( \57834 , \57827 , \57620 );
not \U$57458 ( \57835 , \57834 );
not \U$57459 ( \57836 , \57623 );
and \U$57460 ( \57837 , \57835 , \57836 );
and \U$57461 ( \57838 , \57834 , \57623 );
nor \U$57462 ( \57839 , \57837 , \57838 );
not \U$57463 ( \57840 , \57403 );
not \U$57464 ( \57841 , \57569 );
or \U$57465 ( \57842 , \57840 , \57841 );
or \U$57466 ( \57843 , \57569 , \57403 );
nand \U$57467 ( \57844 , \57842 , \57843 );
not \U$57468 ( \57845 , \57844 );
not \U$57469 ( \57846 , \57418 );
and \U$57470 ( \57847 , \57845 , \57846 );
and \U$57471 ( \57848 , \57844 , \57418 );
nor \U$57472 ( \57849 , \57847 , \57848 );
or \U$57473 ( \57850 , \57839 , \57849 );
not \U$57474 ( \57851 , \57849 );
not \U$57475 ( \57852 , \57839 );
or \U$57476 ( \57853 , \57851 , \57852 );
xor \U$57477 ( \57854 , \57732 , \57739 );
xor \U$57478 ( \57855 , \57854 , \57767 );
xor \U$57479 ( \57856 , \57796 , \57798 );
xor \U$57480 ( \57857 , \57856 , \57801 );
and \U$57481 ( \57858 , \57855 , \57857 );
xor \U$57482 ( \57859 , \57499 , \57506 );
xor \U$57483 ( \57860 , \57859 , \57514 );
xor \U$57484 ( \57861 , \57776 , \57781 );
xor \U$57485 ( \57862 , \57860 , \57861 );
xor \U$57486 ( \57863 , \57796 , \57798 );
xor \U$57487 ( \57864 , \57863 , \57801 );
and \U$57488 ( \57865 , \57862 , \57864 );
and \U$57489 ( \57866 , \57855 , \57862 );
or \U$57490 ( \57867 , \57858 , \57865 , \57866 );
not \U$57491 ( \57868 , \57754 );
not \U$57492 ( \57869 , \57765 );
or \U$57493 ( \57870 , \57868 , \57869 );
or \U$57494 ( \57871 , \57754 , \57765 );
nand \U$57495 ( \57872 , \57870 , \57871 );
not \U$57496 ( \57873 , \57872 );
not \U$57497 ( \57874 , \57747 );
and \U$57498 ( \57875 , \57873 , \57874 );
and \U$57499 ( \57876 , \57872 , \57747 );
nor \U$57500 ( \57877 , \57875 , \57876 );
and \U$57501 ( \57878 , \8371 , RIae76eb0_64);
and \U$57502 ( \57879 , RIae76dc0_62, \8369 );
nor \U$57503 ( \57880 , \57878 , \57879 );
and \U$57504 ( \57881 , \57880 , \8020 );
not \U$57505 ( \57882 , \57880 );
and \U$57506 ( \57883 , \57882 , \8019 );
nor \U$57507 ( \57884 , \57881 , \57883 );
and \U$57508 ( \57885 , \8966 , RIae76cd0_60);
and \U$57509 ( \57886 , RIae77108_69, \8964 );
nor \U$57510 ( \57887 , \57885 , \57886 );
and \U$57511 ( \57888 , \57887 , \8799 );
not \U$57512 ( \57889 , \57887 );
and \U$57513 ( \57890 , \57889 , \8789 );
nor \U$57514 ( \57891 , \57888 , \57890 );
xor \U$57515 ( \57892 , \57884 , \57891 );
and \U$57516 ( \57893 , \7633 , RIae77900_86);
and \U$57517 ( \57894 , RIae76fa0_66, \7631 );
nor \U$57518 ( \57895 , \57893 , \57894 );
and \U$57519 ( \57896 , \57895 , \7206 );
not \U$57520 ( \57897 , \57895 );
and \U$57521 ( \57898 , \57897 , \7205 );
nor \U$57522 ( \57899 , \57896 , \57898 );
and \U$57523 ( \57900 , \57892 , \57899 );
and \U$57524 ( \57901 , \57884 , \57891 );
nor \U$57525 ( \57902 , \57900 , \57901 );
or \U$57526 ( \57903 , \57877 , \57902 );
not \U$57527 ( \57904 , \57902 );
not \U$57528 ( \57905 , \57877 );
or \U$57529 ( \57906 , \57904 , \57905 );
and \U$57530 ( \57907 , \6172 , RIae77450_76);
and \U$57531 ( \57908 , RIae77ae0_90, \6170 );
nor \U$57532 ( \57909 , \57907 , \57908 );
and \U$57533 ( \57910 , \57909 , \6176 );
not \U$57534 ( \57911 , \57909 );
and \U$57535 ( \57912 , \57911 , \6175 );
nor \U$57536 ( \57913 , \57910 , \57912 );
and \U$57537 ( \57914 , \5896 , RIae77540_78);
and \U$57538 ( \57915 , RIae776a8_81, \5894 );
nor \U$57539 ( \57916 , \57914 , \57915 );
and \U$57540 ( \57917 , \57916 , \5590 );
not \U$57541 ( \57918 , \57916 );
and \U$57542 ( \57919 , \57918 , \5589 );
nor \U$57543 ( \57920 , \57917 , \57919 );
xor \U$57544 ( \57921 , \57913 , \57920 );
and \U$57545 ( \57922 , \6941 , RIae779f0_88);
and \U$57546 ( \57923 , RIae77810_84, \6939 );
nor \U$57547 ( \57924 , \57922 , \57923 );
and \U$57548 ( \57925 , \57924 , \6314 );
not \U$57549 ( \57926 , \57924 );
and \U$57550 ( \57927 , \57926 , \6945 );
nor \U$57551 ( \57928 , \57925 , \57927 );
and \U$57552 ( \57929 , \57921 , \57928 );
and \U$57553 ( \57930 , \57913 , \57920 );
or \U$57554 ( \57931 , \57929 , \57930 );
nand \U$57555 ( \57932 , \57906 , \57931 );
nand \U$57556 ( \57933 , \57903 , \57932 );
and \U$57557 ( \57934 , \11470 , RIae78170_104);
and \U$57558 ( \57935 , RIae77f90_100, \11468 );
nor \U$57559 ( \57936 , \57934 , \57935 );
and \U$57560 ( \57937 , \57936 , \10936 );
not \U$57561 ( \57938 , \57936 );
and \U$57562 ( \57939 , \57938 , \11474 );
nor \U$57563 ( \57940 , \57937 , \57939 );
and \U$57564 ( \57941 , \9760 , RIae77090_68);
and \U$57565 ( \57942 , RIae77270_72, \9758 );
nor \U$57566 ( \57943 , \57941 , \57942 );
and \U$57567 ( \57944 , \57943 , \9273 );
not \U$57568 ( \57945 , \57943 );
and \U$57569 ( \57946 , \57945 , \9272 );
nor \U$57570 ( \57947 , \57944 , \57946 );
xor \U$57571 ( \57948 , \57940 , \57947 );
and \U$57572 ( \57949 , \10548 , RIae77360_74);
and \U$57573 ( \57950 , RIae78350_108, \10546 );
nor \U$57574 ( \57951 , \57949 , \57950 );
and \U$57575 ( \57952 , \57951 , \10421 );
not \U$57576 ( \57953 , \57951 );
and \U$57577 ( \57954 , \57953 , \10118 );
nor \U$57578 ( \57955 , \57952 , \57954 );
and \U$57579 ( \57956 , \57948 , \57955 );
and \U$57580 ( \57957 , \57940 , \57947 );
or \U$57581 ( \57958 , \57956 , \57957 );
and \U$57582 ( \57959 , \15726 , RIae77ea0_98);
and \U$57583 ( \57960 , RIae789e0_122, RIae7aab0_192);
nor \U$57584 ( \57961 , \57959 , \57960 );
and \U$57585 ( \57962 , \57961 , \14959 );
not \U$57586 ( \57963 , \57961 );
and \U$57587 ( \57964 , \57963 , RIae7aa38_191);
nor \U$57588 ( \57965 , \57962 , \57964 );
xor \U$57589 ( \57966 , \57965 , \5403 );
and \U$57590 ( \57967 , \14964 , RIae77bd0_92);
and \U$57591 ( \57968 , RIae77db0_96, \14962 );
nor \U$57592 ( \57969 , \57967 , \57968 );
and \U$57593 ( \57970 , \57969 , \14463 );
not \U$57594 ( \57971 , \57969 );
and \U$57595 ( \57972 , \57971 , \14462 );
nor \U$57596 ( \57973 , \57970 , \57972 );
and \U$57597 ( \57974 , \57966 , \57973 );
and \U$57598 ( \57975 , \57965 , \5403 );
or \U$57599 ( \57976 , \57974 , \57975 );
xor \U$57600 ( \57977 , \57958 , \57976 );
and \U$57601 ( \57978 , \14059 , RIae784b8_111);
and \U$57602 ( \57979 , RIae77cc0_94, \14057 );
nor \U$57603 ( \57980 , \57978 , \57979 );
and \U$57604 ( \57981 , \57980 , \13502 );
not \U$57605 ( \57982 , \57980 );
and \U$57606 ( \57983 , \57982 , \14063 );
nor \U$57607 ( \57984 , \57981 , \57983 );
and \U$57608 ( \57985 , \12180 , RIae78080_102);
and \U$57609 ( \57986 , RIae78260_106, \12178 );
nor \U$57610 ( \57987 , \57985 , \57986 );
and \U$57611 ( \57988 , \57987 , \12184 );
not \U$57612 ( \57989 , \57987 );
and \U$57613 ( \57990 , \57989 , \11827 );
nor \U$57614 ( \57991 , \57988 , \57990 );
xor \U$57615 ( \57992 , \57984 , \57991 );
and \U$57616 ( \57993 , \13059 , RIae78620_114);
and \U$57617 ( \57994 , RIae78440_110, \13057 );
nor \U$57618 ( \57995 , \57993 , \57994 );
and \U$57619 ( \57996 , \57995 , \13063 );
not \U$57620 ( \57997 , \57995 );
and \U$57621 ( \57998 , \57997 , \12718 );
nor \U$57622 ( \57999 , \57996 , \57998 );
and \U$57623 ( \58000 , \57992 , \57999 );
and \U$57624 ( \58001 , \57984 , \57991 );
or \U$57625 ( \58002 , \58000 , \58001 );
and \U$57626 ( \58003 , \57977 , \58002 );
and \U$57627 ( \58004 , \57958 , \57976 );
or \U$57628 ( \58005 , \58003 , \58004 );
xor \U$57629 ( \58006 , \57933 , \58005 );
not \U$57630 ( \58007 , \57719 );
not \U$57631 ( \58008 , \57730 );
or \U$57632 ( \58009 , \58007 , \58008 );
or \U$57633 ( \58010 , \57719 , \57730 );
nand \U$57634 ( \58011 , \58009 , \58010 );
not \U$57635 ( \58012 , \58011 );
not \U$57636 ( \58013 , \57712 );
and \U$57637 ( \58014 , \58012 , \58013 );
and \U$57638 ( \58015 , \58011 , \57712 );
nor \U$57639 ( \58016 , \58014 , \58015 );
xor \U$57640 ( \58017 , \57658 , \57665 );
xor \U$57641 ( \58018 , \58017 , \57673 );
or \U$57642 ( \58019 , \58016 , \58018 );
not \U$57643 ( \58020 , \58018 );
not \U$57644 ( \58021 , \58016 );
or \U$57645 ( \58022 , \58020 , \58021 );
xor \U$57646 ( \58023 , \57633 , \57640 );
xor \U$57647 ( \58024 , \58023 , \57648 );
nand \U$57648 ( \58025 , \58022 , \58024 );
nand \U$57649 ( \58026 , \58019 , \58025 );
and \U$57650 ( \58027 , \58006 , \58026 );
and \U$57651 ( \58028 , \57933 , \58005 );
or \U$57652 ( \58029 , \58027 , \58028 );
xor \U$57653 ( \58030 , \57867 , \58029 );
xor \U$57654 ( \58031 , \57445 , \57463 );
xor \U$57655 ( \58032 , \58031 , \57489 );
xor \U$57656 ( \58033 , \57812 , \57819 );
xor \U$57657 ( \58034 , \58032 , \58033 );
and \U$57658 ( \58035 , \58030 , \58034 );
and \U$57659 ( \58036 , \57867 , \58029 );
or \U$57660 ( \58037 , \58035 , \58036 );
xor \U$57661 ( \58038 , \57705 , \57770 );
xor \U$57662 ( \58039 , \58038 , \57786 );
xor \U$57663 ( \58040 , \57213 , \57220 );
xor \U$57664 ( \58041 , \58040 , \57228 );
xor \U$57665 ( \58042 , \57791 , \57804 );
xor \U$57666 ( \58043 , \58041 , \58042 );
and \U$57667 ( \58044 , \58039 , \58043 );
xor \U$57668 ( \58045 , \58037 , \58044 );
xor \U$57669 ( \58046 , \57609 , \57614 );
xor \U$57670 ( \58047 , \58046 , \57617 );
and \U$57671 ( \58048 , \58045 , \58047 );
and \U$57672 ( \58049 , \58037 , \58044 );
or \U$57673 ( \58050 , \58048 , \58049 );
nand \U$57674 ( \58051 , \57853 , \58050 );
nand \U$57675 ( \58052 , \57850 , \58051 );
and \U$57676 ( \58053 , \57833 , \58052 );
xor \U$57677 ( \58054 , \58052 , \57833 );
and \U$57678 ( \58055 , \9760 , RIae76cd0_60);
and \U$57679 ( \58056 , RIae77108_69, \9758 );
nor \U$57680 ( \58057 , \58055 , \58056 );
and \U$57681 ( \58058 , \58057 , \9273 );
not \U$57682 ( \58059 , \58057 );
and \U$57683 ( \58060 , \58059 , \9764 );
nor \U$57684 ( \58061 , \58058 , \58060 );
and \U$57685 ( \58062 , \10548 , RIae77090_68);
and \U$57686 ( \58063 , RIae77270_72, \10546 );
nor \U$57687 ( \58064 , \58062 , \58063 );
and \U$57688 ( \58065 , \58064 , \10421 );
not \U$57689 ( \58066 , \58064 );
and \U$57690 ( \58067 , \58066 , \10118 );
nor \U$57691 ( \58068 , \58065 , \58067 );
xor \U$57692 ( \58069 , \58061 , \58068 );
and \U$57693 ( \58070 , \11470 , RIae77360_74);
and \U$57694 ( \58071 , RIae78350_108, \11468 );
nor \U$57695 ( \58072 , \58070 , \58071 );
and \U$57696 ( \58073 , \58072 , \10936 );
not \U$57697 ( \58074 , \58072 );
and \U$57698 ( \58075 , \58074 , \11474 );
nor \U$57699 ( \58076 , \58073 , \58075 );
and \U$57700 ( \58077 , \58069 , \58076 );
and \U$57701 ( \58078 , \58061 , \58068 );
or \U$57702 ( \58079 , \58077 , \58078 );
and \U$57703 ( \58080 , \15726 , RIae77bd0_92);
and \U$57704 ( \58081 , RIae77db0_96, RIae7aab0_192);
nor \U$57705 ( \58082 , \58080 , \58081 );
and \U$57706 ( \58083 , \58082 , \14959 );
not \U$57707 ( \58084 , \58082 );
and \U$57708 ( \58085 , \58084 , RIae7aa38_191);
nor \U$57709 ( \58086 , \58083 , \58085 );
xor \U$57710 ( \58087 , \58086 , \5589 );
and \U$57711 ( \58088 , \14964 , RIae784b8_111);
and \U$57712 ( \58089 , RIae77cc0_94, \14962 );
nor \U$57713 ( \58090 , \58088 , \58089 );
and \U$57714 ( \58091 , \58090 , \14463 );
not \U$57715 ( \58092 , \58090 );
and \U$57716 ( \58093 , \58092 , \14462 );
nor \U$57717 ( \58094 , \58091 , \58093 );
and \U$57718 ( \58095 , \58087 , \58094 );
and \U$57719 ( \58096 , \58086 , \5589 );
or \U$57720 ( \58097 , \58095 , \58096 );
xor \U$57721 ( \58098 , \58079 , \58097 );
and \U$57722 ( \58099 , \14059 , RIae78620_114);
and \U$57723 ( \58100 , RIae78440_110, \14057 );
nor \U$57724 ( \58101 , \58099 , \58100 );
and \U$57725 ( \58102 , \58101 , \13502 );
not \U$57726 ( \58103 , \58101 );
and \U$57727 ( \58104 , \58103 , \14063 );
nor \U$57728 ( \58105 , \58102 , \58104 );
and \U$57729 ( \58106 , \12180 , RIae78170_104);
and \U$57730 ( \58107 , RIae77f90_100, \12178 );
nor \U$57731 ( \58108 , \58106 , \58107 );
and \U$57732 ( \58109 , \58108 , \12184 );
not \U$57733 ( \58110 , \58108 );
and \U$57734 ( \58111 , \58110 , \11827 );
nor \U$57735 ( \58112 , \58109 , \58111 );
xor \U$57736 ( \58113 , \58105 , \58112 );
and \U$57737 ( \58114 , \13059 , RIae78080_102);
and \U$57738 ( \58115 , RIae78260_106, \13057 );
nor \U$57739 ( \58116 , \58114 , \58115 );
and \U$57740 ( \58117 , \58116 , \13063 );
not \U$57741 ( \58118 , \58116 );
and \U$57742 ( \58119 , \58118 , \12718 );
nor \U$57743 ( \58120 , \58117 , \58119 );
and \U$57744 ( \58121 , \58113 , \58120 );
and \U$57745 ( \58122 , \58105 , \58112 );
or \U$57746 ( \58123 , \58121 , \58122 );
and \U$57747 ( \58124 , \58098 , \58123 );
and \U$57748 ( \58125 , \58079 , \58097 );
or \U$57749 ( \58126 , \58124 , \58125 );
and \U$57750 ( \58127 , \6941 , RIae77450_76);
and \U$57751 ( \58128 , RIae77ae0_90, \6939 );
nor \U$57752 ( \58129 , \58127 , \58128 );
and \U$57753 ( \58130 , \58129 , \6314 );
not \U$57754 ( \58131 , \58129 );
and \U$57755 ( \58132 , \58131 , \6945 );
nor \U$57756 ( \58133 , \58130 , \58132 );
nand \U$57757 ( \58134 , RIae77630_80, \5894 );
and \U$57758 ( \58135 , \58134 , \5590 );
not \U$57759 ( \58136 , \58134 );
and \U$57760 ( \58137 , \58136 , \5589 );
nor \U$57761 ( \58138 , \58135 , \58137 );
xor \U$57762 ( \58139 , \58133 , \58138 );
and \U$57763 ( \58140 , \6172 , RIae77540_78);
and \U$57764 ( \58141 , RIae776a8_81, \6170 );
nor \U$57765 ( \58142 , \58140 , \58141 );
and \U$57766 ( \58143 , \58142 , \6176 );
not \U$57767 ( \58144 , \58142 );
and \U$57768 ( \58145 , \58144 , \6175 );
nor \U$57769 ( \58146 , \58143 , \58145 );
and \U$57770 ( \58147 , \58139 , \58146 );
and \U$57771 ( \58148 , \58133 , \58138 );
or \U$57772 ( \58149 , \58147 , \58148 );
and \U$57773 ( \58150 , \6172 , RIae776a8_81);
and \U$57774 ( \58151 , RIae77450_76, \6170 );
nor \U$57775 ( \58152 , \58150 , \58151 );
and \U$57776 ( \58153 , \58152 , \6176 );
not \U$57777 ( \58154 , \58152 );
and \U$57778 ( \58155 , \58154 , \6175 );
nor \U$57779 ( \58156 , \58153 , \58155 );
xor \U$57780 ( \58157 , \58149 , \58156 );
and \U$57781 ( \58158 , \7633 , RIae779f0_88);
and \U$57782 ( \58159 , RIae77810_84, \7631 );
nor \U$57783 ( \58160 , \58158 , \58159 );
and \U$57784 ( \58161 , \58160 , \7206 );
not \U$57785 ( \58162 , \58160 );
and \U$57786 ( \58163 , \58162 , \7205 );
nor \U$57787 ( \58164 , \58161 , \58163 );
and \U$57788 ( \58165 , \8371 , RIae77900_86);
and \U$57789 ( \58166 , RIae76fa0_66, \8369 );
nor \U$57790 ( \58167 , \58165 , \58166 );
and \U$57791 ( \58168 , \58167 , \8020 );
not \U$57792 ( \58169 , \58167 );
and \U$57793 ( \58170 , \58169 , \8019 );
nor \U$57794 ( \58171 , \58168 , \58170 );
xor \U$57795 ( \58172 , \58164 , \58171 );
and \U$57796 ( \58173 , \8966 , RIae76eb0_64);
and \U$57797 ( \58174 , RIae76dc0_62, \8964 );
nor \U$57798 ( \58175 , \58173 , \58174 );
and \U$57799 ( \58176 , \58175 , \8799 );
not \U$57800 ( \58177 , \58175 );
and \U$57801 ( \58178 , \58177 , \8789 );
nor \U$57802 ( \58179 , \58176 , \58178 );
and \U$57803 ( \58180 , \58172 , \58179 );
and \U$57804 ( \58181 , \58164 , \58171 );
or \U$57805 ( \58182 , \58180 , \58181 );
and \U$57806 ( \58183 , \58157 , \58182 );
and \U$57807 ( \58184 , \58149 , \58156 );
or \U$57808 ( \58185 , \58183 , \58184 );
xor \U$57809 ( \58186 , \58126 , \58185 );
and \U$57810 ( \58187 , \5896 , RIae77630_80);
and \U$57811 ( \58188 , RIae77540_78, \5894 );
nor \U$57812 ( \58189 , \58187 , \58188 );
and \U$57813 ( \58190 , \58189 , \5590 );
not \U$57814 ( \58191 , \58189 );
and \U$57815 ( \58192 , \58191 , \5589 );
nor \U$57816 ( \58193 , \58190 , \58192 );
and \U$57817 ( \58194 , \6941 , RIae77ae0_90);
and \U$57818 ( \58195 , RIae779f0_88, \6939 );
nor \U$57819 ( \58196 , \58194 , \58195 );
and \U$57820 ( \58197 , \58196 , \6314 );
not \U$57821 ( \58198 , \58196 );
and \U$57822 ( \58199 , \58198 , \6945 );
nor \U$57823 ( \58200 , \58197 , \58199 );
and \U$57824 ( \58201 , \7633 , RIae77810_84);
and \U$57825 ( \58202 , RIae77900_86, \7631 );
nor \U$57826 ( \58203 , \58201 , \58202 );
and \U$57827 ( \58204 , \58203 , \7206 );
not \U$57828 ( \58205 , \58203 );
and \U$57829 ( \58206 , \58205 , \7205 );
nor \U$57830 ( \58207 , \58204 , \58206 );
xor \U$57831 ( \58208 , \58200 , \58207 );
and \U$57832 ( \58209 , \8371 , RIae76fa0_66);
and \U$57833 ( \58210 , RIae76eb0_64, \8369 );
nor \U$57834 ( \58211 , \58209 , \58210 );
and \U$57835 ( \58212 , \58211 , \8020 );
not \U$57836 ( \58213 , \58211 );
and \U$57837 ( \58214 , \58213 , \8019 );
nor \U$57838 ( \58215 , \58212 , \58214 );
xor \U$57839 ( \58216 , \58208 , \58215 );
and \U$57840 ( \58217 , \58193 , \58216 );
and \U$57841 ( \58218 , \8966 , RIae76dc0_62);
and \U$57842 ( \58219 , RIae76cd0_60, \8964 );
nor \U$57843 ( \58220 , \58218 , \58219 );
and \U$57844 ( \58221 , \58220 , \8799 );
not \U$57845 ( \58222 , \58220 );
and \U$57846 ( \58223 , \58222 , \8789 );
nor \U$57847 ( \58224 , \58221 , \58223 );
and \U$57848 ( \58225 , \9760 , RIae77108_69);
and \U$57849 ( \58226 , RIae77090_68, \9758 );
nor \U$57850 ( \58227 , \58225 , \58226 );
and \U$57851 ( \58228 , \58227 , \9273 );
not \U$57852 ( \58229 , \58227 );
and \U$57853 ( \58230 , \58229 , \9764 );
nor \U$57854 ( \58231 , \58228 , \58230 );
xor \U$57855 ( \58232 , \58224 , \58231 );
and \U$57856 ( \58233 , \10548 , RIae77270_72);
and \U$57857 ( \58234 , RIae77360_74, \10546 );
nor \U$57858 ( \58235 , \58233 , \58234 );
and \U$57859 ( \58236 , \58235 , \10421 );
not \U$57860 ( \58237 , \58235 );
and \U$57861 ( \58238 , \58237 , \10118 );
nor \U$57862 ( \58239 , \58236 , \58238 );
xor \U$57863 ( \58240 , \58232 , \58239 );
xor \U$57864 ( \58241 , \58200 , \58207 );
xor \U$57865 ( \58242 , \58241 , \58215 );
and \U$57866 ( \58243 , \58240 , \58242 );
and \U$57867 ( \58244 , \58193 , \58240 );
or \U$57868 ( \58245 , \58217 , \58243 , \58244 );
xor \U$57869 ( \58246 , \58186 , \58245 );
and \U$57870 ( \58247 , \11470 , RIae78350_108);
and \U$57871 ( \58248 , RIae78170_104, \11468 );
nor \U$57872 ( \58249 , \58247 , \58248 );
and \U$57873 ( \58250 , \58249 , \10936 );
not \U$57874 ( \58251 , \58249 );
and \U$57875 ( \58252 , \58251 , \11474 );
nor \U$57876 ( \58253 , \58250 , \58252 );
and \U$57877 ( \58254 , \12180 , RIae77f90_100);
and \U$57878 ( \58255 , RIae78080_102, \12178 );
nor \U$57879 ( \58256 , \58254 , \58255 );
and \U$57880 ( \58257 , \58256 , \12184 );
not \U$57881 ( \58258 , \58256 );
and \U$57882 ( \58259 , \58258 , \11827 );
nor \U$57883 ( \58260 , \58257 , \58259 );
xor \U$57884 ( \58261 , \58253 , \58260 );
and \U$57885 ( \58262 , \13059 , RIae78260_106);
and \U$57886 ( \58263 , RIae78620_114, \13057 );
nor \U$57887 ( \58264 , \58262 , \58263 );
and \U$57888 ( \58265 , \58264 , \13063 );
not \U$57889 ( \58266 , \58264 );
and \U$57890 ( \58267 , \58266 , \12718 );
nor \U$57891 ( \58268 , \58265 , \58267 );
xor \U$57892 ( \58269 , \58261 , \58268 );
and \U$57893 ( \58270 , \14964 , RIae77cc0_94);
and \U$57894 ( \58271 , RIae77bd0_92, \14962 );
nor \U$57895 ( \58272 , \58270 , \58271 );
and \U$57896 ( \58273 , \58272 , \14463 );
not \U$57897 ( \58274 , \58272 );
and \U$57898 ( \58275 , \58274 , \14462 );
nor \U$57899 ( \58276 , \58273 , \58275 );
and \U$57900 ( \58277 , \15726 , RIae77db0_96);
and \U$57901 ( \58278 , RIae77ea0_98, RIae7aab0_192);
nor \U$57902 ( \58279 , \58277 , \58278 );
and \U$57903 ( \58280 , \58279 , \14959 );
not \U$57904 ( \58281 , \58279 );
and \U$57905 ( \58282 , \58281 , RIae7aa38_191);
nor \U$57906 ( \58283 , \58280 , \58282 );
xor \U$57907 ( \58284 , \58276 , \58283 );
and \U$57908 ( \58285 , \14059 , RIae78440_110);
and \U$57909 ( \58286 , RIae784b8_111, \14057 );
nor \U$57910 ( \58287 , \58285 , \58286 );
and \U$57911 ( \58288 , \58287 , \13502 );
not \U$57912 ( \58289 , \58287 );
and \U$57913 ( \58290 , \58289 , \14063 );
nor \U$57914 ( \58291 , \58288 , \58290 );
xor \U$57915 ( \58292 , \58284 , \58291 );
xor \U$57916 ( \58293 , \58269 , \58292 );
xor \U$57917 ( \58294 , \58200 , \58207 );
xor \U$57918 ( \58295 , \58294 , \58215 );
xor \U$57919 ( \58296 , \58193 , \58240 );
xor \U$57920 ( \58297 , \58295 , \58296 );
and \U$57921 ( \58298 , \58293 , \58297 );
and \U$57922 ( \58299 , \58269 , \58292 );
or \U$57923 ( \58300 , \58298 , \58299 );
xor \U$57924 ( \58301 , \58224 , \58231 );
and \U$57925 ( \58302 , \58301 , \58239 );
and \U$57926 ( \58303 , \58224 , \58231 );
or \U$57927 ( \58304 , \58302 , \58303 );
xor \U$57928 ( \58305 , \58276 , \58283 );
and \U$57929 ( \58306 , \58305 , \58291 );
and \U$57930 ( \58307 , \58276 , \58283 );
or \U$57931 ( \58308 , \58306 , \58307 );
xor \U$57932 ( \58309 , \58304 , \58308 );
xor \U$57933 ( \58310 , \58253 , \58260 );
and \U$57934 ( \58311 , \58310 , \58268 );
and \U$57935 ( \58312 , \58253 , \58260 );
or \U$57936 ( \58313 , \58311 , \58312 );
xor \U$57937 ( \58314 , \58309 , \58313 );
xor \U$57938 ( \58315 , \58300 , \58314 );
xor \U$57939 ( \58316 , \58133 , \58138 );
xor \U$57940 ( \58317 , \58316 , \58146 );
and \U$57941 ( \58318 , \6941 , RIae776a8_81);
and \U$57942 ( \58319 , RIae77450_76, \6939 );
nor \U$57943 ( \58320 , \58318 , \58319 );
and \U$57944 ( \58321 , \58320 , \6945 );
not \U$57945 ( \58322 , \58320 );
and \U$57946 ( \58323 , \58322 , \6314 );
nor \U$57947 ( \58324 , \58321 , \58323 );
and \U$57948 ( \58325 , \8371 , RIae77810_84);
and \U$57949 ( \58326 , RIae77900_86, \8369 );
nor \U$57950 ( \58327 , \58325 , \58326 );
and \U$57951 ( \58328 , \58327 , \8019 );
not \U$57952 ( \58329 , \58327 );
and \U$57953 ( \58330 , \58329 , \8020 );
nor \U$57954 ( \58331 , \58328 , \58330 );
or \U$57955 ( \58332 , \58324 , \58331 );
not \U$57956 ( \58333 , \58331 );
not \U$57957 ( \58334 , \58324 );
or \U$57958 ( \58335 , \58333 , \58334 );
and \U$57959 ( \58336 , \7633 , RIae77ae0_90);
and \U$57960 ( \58337 , RIae779f0_88, \7631 );
nor \U$57961 ( \58338 , \58336 , \58337 );
and \U$57962 ( \58339 , \58338 , \7206 );
not \U$57963 ( \58340 , \58338 );
and \U$57964 ( \58341 , \58340 , \7205 );
nor \U$57965 ( \58342 , \58339 , \58341 );
nand \U$57966 ( \58343 , \58335 , \58342 );
nand \U$57967 ( \58344 , \58332 , \58343 );
xor \U$57968 ( \58345 , \58317 , \58344 );
xor \U$57969 ( \58346 , \58164 , \58171 );
xor \U$57970 ( \58347 , \58346 , \58179 );
and \U$57971 ( \58348 , \58345 , \58347 );
and \U$57972 ( \58349 , \58317 , \58344 );
or \U$57973 ( \58350 , \58348 , \58349 );
and \U$57974 ( \58351 , \11470 , RIae77270_72);
and \U$57975 ( \58352 , RIae77360_74, \11468 );
nor \U$57976 ( \58353 , \58351 , \58352 );
and \U$57977 ( \58354 , \58353 , \11474 );
not \U$57978 ( \58355 , \58353 );
and \U$57979 ( \58356 , \58355 , \10936 );
nor \U$57980 ( \58357 , \58354 , \58356 );
and \U$57981 ( \58358 , \13059 , RIae77f90_100);
and \U$57982 ( \58359 , RIae78080_102, \13057 );
nor \U$57983 ( \58360 , \58358 , \58359 );
and \U$57984 ( \58361 , \58360 , \12718 );
not \U$57985 ( \58362 , \58360 );
and \U$57986 ( \58363 , \58362 , \13063 );
nor \U$57987 ( \58364 , \58361 , \58363 );
or \U$57988 ( \58365 , \58357 , \58364 );
not \U$57989 ( \58366 , \58364 );
not \U$57990 ( \58367 , \58357 );
or \U$57991 ( \58368 , \58366 , \58367 );
and \U$57992 ( \58369 , \12180 , RIae78350_108);
and \U$57993 ( \58370 , RIae78170_104, \12178 );
nor \U$57994 ( \58371 , \58369 , \58370 );
and \U$57995 ( \58372 , \58371 , \12184 );
not \U$57996 ( \58373 , \58371 );
and \U$57997 ( \58374 , \58373 , \11827 );
nor \U$57998 ( \58375 , \58372 , \58374 );
nand \U$57999 ( \58376 , \58368 , \58375 );
nand \U$58000 ( \58377 , \58365 , \58376 );
and \U$58001 ( \58378 , \15726 , RIae77cc0_94);
and \U$58002 ( \58379 , RIae77bd0_92, RIae7aab0_192);
nor \U$58003 ( \58380 , \58378 , \58379 );
and \U$58004 ( \58381 , \58380 , RIae7aa38_191);
not \U$58005 ( \58382 , \58380 );
and \U$58006 ( \58383 , \58382 , \14959 );
nor \U$58007 ( \58384 , \58381 , \58383 );
and \U$58008 ( \58385 , \14964 , RIae78440_110);
and \U$58009 ( \58386 , RIae784b8_111, \14962 );
nor \U$58010 ( \58387 , \58385 , \58386 );
and \U$58011 ( \58388 , \58387 , \14462 );
not \U$58012 ( \58389 , \58387 );
and \U$58013 ( \58390 , \58389 , \14463 );
nor \U$58014 ( \58391 , \58388 , \58390 );
xor \U$58015 ( \58392 , \58384 , \58391 );
and \U$58016 ( \58393 , \14059 , RIae78260_106);
and \U$58017 ( \58394 , RIae78620_114, \14057 );
nor \U$58018 ( \58395 , \58393 , \58394 );
and \U$58019 ( \58396 , \58395 , \14063 );
not \U$58020 ( \58397 , \58395 );
and \U$58021 ( \58398 , \58397 , \13502 );
nor \U$58022 ( \58399 , \58396 , \58398 );
and \U$58023 ( \58400 , \58392 , \58399 );
and \U$58024 ( \58401 , \58384 , \58391 );
nor \U$58025 ( \58402 , \58400 , \58401 );
xor \U$58026 ( \58403 , \58377 , \58402 );
and \U$58027 ( \58404 , \8966 , RIae76fa0_66);
and \U$58028 ( \58405 , RIae76eb0_64, \8964 );
nor \U$58029 ( \58406 , \58404 , \58405 );
and \U$58030 ( \58407 , \58406 , \8789 );
not \U$58031 ( \58408 , \58406 );
and \U$58032 ( \58409 , \58408 , \8799 );
nor \U$58033 ( \58410 , \58407 , \58409 );
and \U$58034 ( \58411 , \10548 , RIae77108_69);
and \U$58035 ( \58412 , RIae77090_68, \10546 );
nor \U$58036 ( \58413 , \58411 , \58412 );
and \U$58037 ( \58414 , \58413 , \10118 );
not \U$58038 ( \58415 , \58413 );
and \U$58039 ( \58416 , \58415 , \10421 );
nor \U$58040 ( \58417 , \58414 , \58416 );
or \U$58041 ( \58418 , \58410 , \58417 );
not \U$58042 ( \58419 , \58417 );
not \U$58043 ( \58420 , \58410 );
or \U$58044 ( \58421 , \58419 , \58420 );
and \U$58045 ( \58422 , \9760 , RIae76dc0_62);
and \U$58046 ( \58423 , RIae76cd0_60, \9758 );
nor \U$58047 ( \58424 , \58422 , \58423 );
and \U$58048 ( \58425 , \58424 , \9273 );
not \U$58049 ( \58426 , \58424 );
and \U$58050 ( \58427 , \58426 , \9272 );
nor \U$58051 ( \58428 , \58425 , \58427 );
nand \U$58052 ( \58429 , \58421 , \58428 );
nand \U$58053 ( \58430 , \58418 , \58429 );
and \U$58054 ( \58431 , \58403 , \58430 );
and \U$58055 ( \58432 , \58377 , \58402 );
or \U$58056 ( \58433 , \58431 , \58432 );
xor \U$58057 ( \58434 , \58350 , \58433 );
xor \U$58058 ( \58435 , \58105 , \58112 );
xor \U$58059 ( \58436 , \58435 , \58120 );
xor \U$58060 ( \58437 , \58061 , \58068 );
xor \U$58061 ( \58438 , \58437 , \58076 );
and \U$58062 ( \58439 , \58436 , \58438 );
xor \U$58063 ( \58440 , \58086 , \5589 );
xor \U$58064 ( \58441 , \58440 , \58094 );
xor \U$58065 ( \58442 , \58061 , \58068 );
xor \U$58066 ( \58443 , \58442 , \58076 );
and \U$58067 ( \58444 , \58441 , \58443 );
and \U$58068 ( \58445 , \58436 , \58441 );
or \U$58069 ( \58446 , \58439 , \58444 , \58445 );
and \U$58070 ( \58447 , \58434 , \58446 );
and \U$58071 ( \58448 , \58350 , \58433 );
or \U$58072 ( \58449 , \58447 , \58448 );
xor \U$58073 ( \58450 , \58315 , \58449 );
xor \U$58074 ( \58451 , \58246 , \58450 );
xor \U$58075 ( \58452 , \58079 , \58097 );
xor \U$58076 ( \58453 , \58452 , \58123 );
xor \U$58077 ( \58454 , \58269 , \58292 );
xor \U$58078 ( \58455 , \58454 , \58297 );
and \U$58079 ( \58456 , \58453 , \58455 );
xor \U$58080 ( \58457 , \58350 , \58433 );
xor \U$58081 ( \58458 , \58457 , \58446 );
xor \U$58082 ( \58459 , \58269 , \58292 );
xor \U$58083 ( \58460 , \58459 , \58297 );
and \U$58084 ( \58461 , \58458 , \58460 );
and \U$58085 ( \58462 , \58453 , \58458 );
or \U$58086 ( \58463 , \58456 , \58461 , \58462 );
xor \U$58087 ( \58464 , \58200 , \58207 );
and \U$58088 ( \58465 , \58464 , \58215 );
and \U$58089 ( \58466 , \58200 , \58207 );
or \U$58090 ( \58467 , \58465 , \58466 );
nand \U$58091 ( \58468 , RIae77630_80, \5397 );
and \U$58092 ( \58469 , \58468 , \5016 );
not \U$58093 ( \58470 , \58468 );
and \U$58094 ( \58471 , \58470 , \5403 );
nor \U$58095 ( \58472 , \58469 , \58471 );
xor \U$58096 ( \58473 , \58467 , \58472 );
xor \U$58097 ( \58474 , \57913 , \57920 );
xor \U$58098 ( \58475 , \58474 , \57928 );
xor \U$58099 ( \58476 , \58473 , \58475 );
xor \U$58100 ( \58477 , \57965 , \5403 );
xor \U$58101 ( \58478 , \58477 , \57973 );
xor \U$58102 ( \58479 , \57940 , \57947 );
xor \U$58103 ( \58480 , \58479 , \57955 );
xor \U$58104 ( \58481 , \57884 , \57891 );
xor \U$58105 ( \58482 , \58481 , \57899 );
xor \U$58106 ( \58483 , \57984 , \57991 );
xor \U$58107 ( \58484 , \58483 , \57999 );
xor \U$58108 ( \58485 , \58482 , \58484 );
xor \U$58109 ( \58486 , \58480 , \58485 );
xor \U$58110 ( \58487 , \58478 , \58486 );
xor \U$58111 ( \58488 , \58476 , \58487 );
xor \U$58112 ( \58489 , \58463 , \58488 );
and \U$58113 ( \58490 , \12180 , RIae77360_74);
and \U$58114 ( \58491 , RIae78350_108, \12178 );
nor \U$58115 ( \58492 , \58490 , \58491 );
and \U$58116 ( \58493 , \58492 , \12184 );
not \U$58117 ( \58494 , \58492 );
and \U$58118 ( \58495 , \58494 , \11827 );
nor \U$58119 ( \58496 , \58493 , \58495 );
and \U$58120 ( \58497 , \13059 , RIae78170_104);
and \U$58121 ( \58498 , RIae77f90_100, \13057 );
nor \U$58122 ( \58499 , \58497 , \58498 );
and \U$58123 ( \58500 , \58499 , \13063 );
not \U$58124 ( \58501 , \58499 );
and \U$58125 ( \58502 , \58501 , \12718 );
nor \U$58126 ( \58503 , \58500 , \58502 );
xor \U$58127 ( \58504 , \58496 , \58503 );
and \U$58128 ( \58505 , \14059 , RIae78080_102);
and \U$58129 ( \58506 , RIae78260_106, \14057 );
nor \U$58130 ( \58507 , \58505 , \58506 );
and \U$58131 ( \58508 , \58507 , \13502 );
not \U$58132 ( \58509 , \58507 );
and \U$58133 ( \58510 , \58509 , \14063 );
nor \U$58134 ( \58511 , \58508 , \58510 );
and \U$58135 ( \58512 , \58504 , \58511 );
and \U$58136 ( \58513 , \58496 , \58503 );
or \U$58137 ( \58514 , \58512 , \58513 );
and \U$58138 ( \58515 , \15726 , RIae784b8_111);
and \U$58139 ( \58516 , RIae77cc0_94, RIae7aab0_192);
nor \U$58140 ( \58517 , \58515 , \58516 );
and \U$58141 ( \58518 , \58517 , \14959 );
not \U$58142 ( \58519 , \58517 );
and \U$58143 ( \58520 , \58519 , RIae7aa38_191);
nor \U$58144 ( \58521 , \58518 , \58520 );
xor \U$58145 ( \58522 , \58521 , \6175 );
and \U$58146 ( \58523 , \14964 , RIae78620_114);
and \U$58147 ( \58524 , RIae78440_110, \14962 );
nor \U$58148 ( \58525 , \58523 , \58524 );
and \U$58149 ( \58526 , \58525 , \14463 );
not \U$58150 ( \58527 , \58525 );
and \U$58151 ( \58528 , \58527 , \14462 );
nor \U$58152 ( \58529 , \58526 , \58528 );
and \U$58153 ( \58530 , \58522 , \58529 );
and \U$58154 ( \58531 , \58521 , \6175 );
or \U$58155 ( \58532 , \58530 , \58531 );
xor \U$58156 ( \58533 , \58514 , \58532 );
and \U$58157 ( \58534 , \11470 , RIae77090_68);
and \U$58158 ( \58535 , RIae77270_72, \11468 );
nor \U$58159 ( \58536 , \58534 , \58535 );
and \U$58160 ( \58537 , \58536 , \10936 );
not \U$58161 ( \58538 , \58536 );
and \U$58162 ( \58539 , \58538 , \11474 );
nor \U$58163 ( \58540 , \58537 , \58539 );
and \U$58164 ( \58541 , \9760 , RIae76eb0_64);
and \U$58165 ( \58542 , RIae76dc0_62, \9758 );
nor \U$58166 ( \58543 , \58541 , \58542 );
and \U$58167 ( \58544 , \58543 , \9273 );
not \U$58168 ( \58545 , \58543 );
and \U$58169 ( \58546 , \58545 , \9272 );
nor \U$58170 ( \58547 , \58544 , \58546 );
xor \U$58171 ( \58548 , \58540 , \58547 );
and \U$58172 ( \58549 , \10548 , RIae76cd0_60);
and \U$58173 ( \58550 , RIae77108_69, \10546 );
nor \U$58174 ( \58551 , \58549 , \58550 );
and \U$58175 ( \58552 , \58551 , \10421 );
not \U$58176 ( \58553 , \58551 );
and \U$58177 ( \58554 , \58553 , \10118 );
nor \U$58178 ( \58555 , \58552 , \58554 );
and \U$58179 ( \58556 , \58548 , \58555 );
and \U$58180 ( \58557 , \58540 , \58547 );
or \U$58181 ( \58558 , \58556 , \58557 );
and \U$58182 ( \58559 , \58533 , \58558 );
and \U$58183 ( \58560 , \58514 , \58532 );
or \U$58184 ( \58561 , \58559 , \58560 );
and \U$58185 ( \58562 , \6172 , RIae77630_80);
and \U$58186 ( \58563 , RIae77540_78, \6170 );
nor \U$58187 ( \58564 , \58562 , \58563 );
and \U$58188 ( \58565 , \58564 , \6176 );
not \U$58189 ( \58566 , \58564 );
and \U$58190 ( \58567 , \58566 , \6175 );
nor \U$58191 ( \58568 , \58565 , \58567 );
not \U$58192 ( \58569 , \58568 );
nand \U$58193 ( \58570 , RIae77630_80, \6170 );
and \U$58194 ( \58571 , \58570 , \6176 );
not \U$58195 ( \58572 , \58570 );
and \U$58196 ( \58573 , \58572 , \6175 );
nor \U$58197 ( \58574 , \58571 , \58573 );
and \U$58198 ( \58575 , \6941 , RIae77540_78);
and \U$58199 ( \58576 , RIae776a8_81, \6939 );
nor \U$58200 ( \58577 , \58575 , \58576 );
and \U$58201 ( \58578 , \58577 , \6314 );
not \U$58202 ( \58579 , \58577 );
and \U$58203 ( \58580 , \58579 , \6945 );
nor \U$58204 ( \58581 , \58578 , \58580 );
and \U$58205 ( \58582 , \58574 , \58581 );
not \U$58206 ( \58583 , \58582 );
or \U$58207 ( \58584 , \58569 , \58583 );
or \U$58208 ( \58585 , \58582 , \58568 );
and \U$58209 ( \58586 , \8371 , RIae779f0_88);
and \U$58210 ( \58587 , RIae77810_84, \8369 );
nor \U$58211 ( \58588 , \58586 , \58587 );
and \U$58212 ( \58589 , \58588 , \8020 );
not \U$58213 ( \58590 , \58588 );
and \U$58214 ( \58591 , \58590 , \8019 );
nor \U$58215 ( \58592 , \58589 , \58591 );
and \U$58216 ( \58593 , \7633 , RIae77450_76);
and \U$58217 ( \58594 , RIae77ae0_90, \7631 );
nor \U$58218 ( \58595 , \58593 , \58594 );
and \U$58219 ( \58596 , \58595 , \7206 );
not \U$58220 ( \58597 , \58595 );
and \U$58221 ( \58598 , \58597 , \7205 );
nor \U$58222 ( \58599 , \58596 , \58598 );
xor \U$58223 ( \58600 , \58592 , \58599 );
and \U$58224 ( \58601 , \8966 , RIae77900_86);
and \U$58225 ( \58602 , RIae76fa0_66, \8964 );
nor \U$58226 ( \58603 , \58601 , \58602 );
and \U$58227 ( \58604 , \58603 , \8799 );
not \U$58228 ( \58605 , \58603 );
and \U$58229 ( \58606 , \58605 , \8789 );
nor \U$58230 ( \58607 , \58604 , \58606 );
and \U$58231 ( \58608 , \58600 , \58607 );
and \U$58232 ( \58609 , \58592 , \58599 );
or \U$58233 ( \58610 , \58608 , \58609 );
nand \U$58234 ( \58611 , \58585 , \58610 );
nand \U$58235 ( \58612 , \58584 , \58611 );
xor \U$58236 ( \58613 , \58561 , \58612 );
not \U$58237 ( \58614 , \58331 );
not \U$58238 ( \58615 , \58342 );
or \U$58239 ( \58616 , \58614 , \58615 );
or \U$58240 ( \58617 , \58331 , \58342 );
nand \U$58241 ( \58618 , \58616 , \58617 );
not \U$58242 ( \58619 , \58618 );
not \U$58243 ( \58620 , \58324 );
and \U$58244 ( \58621 , \58619 , \58620 );
and \U$58245 ( \58622 , \58618 , \58324 );
nor \U$58246 ( \58623 , \58621 , \58622 );
not \U$58247 ( \58624 , \58364 );
not \U$58248 ( \58625 , \58375 );
or \U$58249 ( \58626 , \58624 , \58625 );
or \U$58250 ( \58627 , \58364 , \58375 );
nand \U$58251 ( \58628 , \58626 , \58627 );
not \U$58252 ( \58629 , \58628 );
not \U$58253 ( \58630 , \58357 );
and \U$58254 ( \58631 , \58629 , \58630 );
and \U$58255 ( \58632 , \58628 , \58357 );
nor \U$58256 ( \58633 , \58631 , \58632 );
xor \U$58257 ( \58634 , \58623 , \58633 );
not \U$58258 ( \58635 , \58417 );
not \U$58259 ( \58636 , \58428 );
or \U$58260 ( \58637 , \58635 , \58636 );
or \U$58261 ( \58638 , \58417 , \58428 );
nand \U$58262 ( \58639 , \58637 , \58638 );
not \U$58263 ( \58640 , \58639 );
not \U$58264 ( \58641 , \58410 );
and \U$58265 ( \58642 , \58640 , \58641 );
and \U$58266 ( \58643 , \58639 , \58410 );
nor \U$58267 ( \58644 , \58642 , \58643 );
and \U$58268 ( \58645 , \58634 , \58644 );
and \U$58269 ( \58646 , \58623 , \58633 );
nor \U$58270 ( \58647 , \58645 , \58646 );
and \U$58271 ( \58648 , \58613 , \58647 );
and \U$58272 ( \58649 , \58561 , \58612 );
or \U$58273 ( \58650 , \58648 , \58649 );
xor \U$58274 ( \58651 , \58149 , \58156 );
xor \U$58275 ( \58652 , \58651 , \58182 );
xor \U$58276 ( \58653 , \58650 , \58652 );
xor \U$58277 ( \58654 , \58377 , \58402 );
xor \U$58278 ( \58655 , \58654 , \58430 );
xor \U$58279 ( \58656 , \58317 , \58344 );
xor \U$58280 ( \58657 , \58656 , \58347 );
and \U$58281 ( \58658 , \58655 , \58657 );
xor \U$58282 ( \58659 , \58061 , \58068 );
xor \U$58283 ( \58660 , \58659 , \58076 );
xor \U$58284 ( \58661 , \58436 , \58441 );
xor \U$58285 ( \58662 , \58660 , \58661 );
xor \U$58286 ( \58663 , \58317 , \58344 );
xor \U$58287 ( \58664 , \58663 , \58347 );
and \U$58288 ( \58665 , \58662 , \58664 );
and \U$58289 ( \58666 , \58655 , \58662 );
or \U$58290 ( \58667 , \58658 , \58665 , \58666 );
and \U$58291 ( \58668 , \58653 , \58667 );
and \U$58292 ( \58669 , \58650 , \58652 );
or \U$58293 ( \58670 , \58668 , \58669 );
xor \U$58294 ( \58671 , \58489 , \58670 );
xor \U$58295 ( \58672 , \58451 , \58671 );
xor \U$58296 ( \58673 , \58384 , \58391 );
xor \U$58297 ( \58674 , \58673 , \58399 );
xnor \U$58298 ( \58675 , \58610 , \58582 );
not \U$58299 ( \58676 , \58675 );
not \U$58300 ( \58677 , \58568 );
and \U$58301 ( \58678 , \58676 , \58677 );
and \U$58302 ( \58679 , \58675 , \58568 );
nor \U$58303 ( \58680 , \58678 , \58679 );
xor \U$58304 ( \58681 , \58674 , \58680 );
xor \U$58305 ( \58682 , \58623 , \58633 );
xor \U$58306 ( \58683 , \58682 , \58644 );
and \U$58307 ( \58684 , \58681 , \58683 );
and \U$58308 ( \58685 , \58674 , \58680 );
nor \U$58309 ( \58686 , \58684 , \58685 );
not \U$58310 ( \58687 , \58686 );
xor \U$58311 ( \58688 , \58317 , \58344 );
xor \U$58312 ( \58689 , \58688 , \58347 );
xor \U$58313 ( \58690 , \58655 , \58662 );
xor \U$58314 ( \58691 , \58689 , \58690 );
not \U$58315 ( \58692 , \58691 );
or \U$58316 ( \58693 , \58687 , \58692 );
or \U$58317 ( \58694 , \58691 , \58686 );
and \U$58318 ( \58695 , \6941 , RIae77630_80);
and \U$58319 ( \58696 , RIae77540_78, \6939 );
nor \U$58320 ( \58697 , \58695 , \58696 );
and \U$58321 ( \58698 , \58697 , \6945 );
not \U$58322 ( \58699 , \58697 );
and \U$58323 ( \58700 , \58699 , \6314 );
nor \U$58324 ( \58701 , \58698 , \58700 );
and \U$58325 ( \58702 , \8371 , RIae77ae0_90);
and \U$58326 ( \58703 , RIae779f0_88, \8369 );
nor \U$58327 ( \58704 , \58702 , \58703 );
and \U$58328 ( \58705 , \58704 , \8019 );
not \U$58329 ( \58706 , \58704 );
and \U$58330 ( \58707 , \58706 , \8020 );
nor \U$58331 ( \58708 , \58705 , \58707 );
or \U$58332 ( \58709 , \58701 , \58708 );
not \U$58333 ( \58710 , \58708 );
not \U$58334 ( \58711 , \58701 );
or \U$58335 ( \58712 , \58710 , \58711 );
and \U$58336 ( \58713 , \7633 , RIae776a8_81);
and \U$58337 ( \58714 , RIae77450_76, \7631 );
nor \U$58338 ( \58715 , \58713 , \58714 );
and \U$58339 ( \58716 , \58715 , \7206 );
not \U$58340 ( \58717 , \58715 );
and \U$58341 ( \58718 , \58717 , \7205 );
nor \U$58342 ( \58719 , \58716 , \58718 );
nand \U$58343 ( \58720 , \58712 , \58719 );
nand \U$58344 ( \58721 , \58709 , \58720 );
xor \U$58345 ( \58722 , \58574 , \58581 );
xor \U$58346 ( \58723 , \58721 , \58722 );
xor \U$58347 ( \58724 , \58592 , \58599 );
xor \U$58348 ( \58725 , \58724 , \58607 );
and \U$58349 ( \58726 , \58723 , \58725 );
and \U$58350 ( \58727 , \58721 , \58722 );
or \U$58351 ( \58728 , \58726 , \58727 );
and \U$58352 ( \58729 , \8966 , RIae77810_84);
and \U$58353 ( \58730 , RIae77900_86, \8964 );
nor \U$58354 ( \58731 , \58729 , \58730 );
and \U$58355 ( \58732 , \58731 , \8789 );
not \U$58356 ( \58733 , \58731 );
and \U$58357 ( \58734 , \58733 , \8799 );
nor \U$58358 ( \58735 , \58732 , \58734 );
and \U$58359 ( \58736 , \9760 , RIae76fa0_66);
and \U$58360 ( \58737 , RIae76eb0_64, \9758 );
nor \U$58361 ( \58738 , \58736 , \58737 );
and \U$58362 ( \58739 , \58738 , \9272 );
not \U$58363 ( \58740 , \58738 );
and \U$58364 ( \58741 , \58740 , \9273 );
nor \U$58365 ( \58742 , \58739 , \58741 );
or \U$58366 ( \58743 , \58735 , \58742 );
not \U$58367 ( \58744 , \58742 );
not \U$58368 ( \58745 , \58735 );
or \U$58369 ( \58746 , \58744 , \58745 );
and \U$58370 ( \58747 , \10548 , RIae76dc0_62);
and \U$58371 ( \58748 , RIae76cd0_60, \10546 );
nor \U$58372 ( \58749 , \58747 , \58748 );
and \U$58373 ( \58750 , \58749 , \10421 );
not \U$58374 ( \58751 , \58749 );
and \U$58375 ( \58752 , \58751 , \10118 );
nor \U$58376 ( \58753 , \58750 , \58752 );
nand \U$58377 ( \58754 , \58746 , \58753 );
nand \U$58378 ( \58755 , \58743 , \58754 );
and \U$58379 ( \58756 , \15726 , RIae78440_110);
and \U$58380 ( \58757 , RIae784b8_111, RIae7aab0_192);
nor \U$58381 ( \58758 , \58756 , \58757 );
and \U$58382 ( \58759 , \58758 , RIae7aa38_191);
not \U$58383 ( \58760 , \58758 );
and \U$58384 ( \58761 , \58760 , \14959 );
nor \U$58385 ( \58762 , \58759 , \58761 );
and \U$58386 ( \58763 , \14964 , RIae78260_106);
and \U$58387 ( \58764 , RIae78620_114, \14962 );
nor \U$58388 ( \58765 , \58763 , \58764 );
and \U$58389 ( \58766 , \58765 , \14462 );
not \U$58390 ( \58767 , \58765 );
and \U$58391 ( \58768 , \58767 , \14463 );
nor \U$58392 ( \58769 , \58766 , \58768 );
xor \U$58393 ( \58770 , \58762 , \58769 );
and \U$58394 ( \58771 , \14059 , RIae77f90_100);
and \U$58395 ( \58772 , RIae78080_102, \14057 );
nor \U$58396 ( \58773 , \58771 , \58772 );
and \U$58397 ( \58774 , \58773 , \14063 );
not \U$58398 ( \58775 , \58773 );
and \U$58399 ( \58776 , \58775 , \13502 );
nor \U$58400 ( \58777 , \58774 , \58776 );
and \U$58401 ( \58778 , \58770 , \58777 );
and \U$58402 ( \58779 , \58762 , \58769 );
nor \U$58403 ( \58780 , \58778 , \58779 );
xor \U$58404 ( \58781 , \58755 , \58780 );
and \U$58405 ( \58782 , \11470 , RIae77108_69);
and \U$58406 ( \58783 , RIae77090_68, \11468 );
nor \U$58407 ( \58784 , \58782 , \58783 );
and \U$58408 ( \58785 , \58784 , \10936 );
not \U$58409 ( \58786 , \58784 );
and \U$58410 ( \58787 , \58786 , \11474 );
nor \U$58411 ( \58788 , \58785 , \58787 );
and \U$58412 ( \58789 , \12180 , RIae77270_72);
and \U$58413 ( \58790 , RIae77360_74, \12178 );
nor \U$58414 ( \58791 , \58789 , \58790 );
and \U$58415 ( \58792 , \58791 , \12184 );
not \U$58416 ( \58793 , \58791 );
and \U$58417 ( \58794 , \58793 , \11827 );
nor \U$58418 ( \58795 , \58792 , \58794 );
xor \U$58419 ( \58796 , \58788 , \58795 );
and \U$58420 ( \58797 , \13059 , RIae78350_108);
and \U$58421 ( \58798 , RIae78170_104, \13057 );
nor \U$58422 ( \58799 , \58797 , \58798 );
and \U$58423 ( \58800 , \58799 , \13063 );
not \U$58424 ( \58801 , \58799 );
and \U$58425 ( \58802 , \58801 , \12718 );
nor \U$58426 ( \58803 , \58800 , \58802 );
and \U$58427 ( \58804 , \58796 , \58803 );
and \U$58428 ( \58805 , \58788 , \58795 );
or \U$58429 ( \58806 , \58804 , \58805 );
and \U$58430 ( \58807 , \58781 , \58806 );
and \U$58431 ( \58808 , \58755 , \58780 );
or \U$58432 ( \58809 , \58807 , \58808 );
xor \U$58433 ( \58810 , \58728 , \58809 );
xor \U$58434 ( \58811 , \58540 , \58547 );
xor \U$58435 ( \58812 , \58811 , \58555 );
xor \U$58436 ( \58813 , \58496 , \58503 );
xor \U$58437 ( \58814 , \58813 , \58511 );
and \U$58438 ( \58815 , \58812 , \58814 );
xor \U$58439 ( \58816 , \58521 , \6175 );
xor \U$58440 ( \58817 , \58816 , \58529 );
xor \U$58441 ( \58818 , \58496 , \58503 );
xor \U$58442 ( \58819 , \58818 , \58511 );
and \U$58443 ( \58820 , \58817 , \58819 );
and \U$58444 ( \58821 , \58812 , \58817 );
or \U$58445 ( \58822 , \58815 , \58820 , \58821 );
and \U$58446 ( \58823 , \58810 , \58822 );
and \U$58447 ( \58824 , \58728 , \58809 );
or \U$58448 ( \58825 , \58823 , \58824 );
nand \U$58449 ( \58826 , \58694 , \58825 );
nand \U$58450 ( \58827 , \58693 , \58826 );
xor \U$58451 ( \58828 , \58650 , \58652 );
xor \U$58452 ( \58829 , \58828 , \58667 );
and \U$58453 ( \58830 , \58827 , \58829 );
xor \U$58454 ( \58831 , \58269 , \58292 );
xor \U$58455 ( \58832 , \58831 , \58297 );
xor \U$58456 ( \58833 , \58453 , \58458 );
xor \U$58457 ( \58834 , \58832 , \58833 );
xor \U$58458 ( \58835 , \58650 , \58652 );
xor \U$58459 ( \58836 , \58835 , \58667 );
and \U$58460 ( \58837 , \58834 , \58836 );
and \U$58461 ( \58838 , \58827 , \58834 );
or \U$58462 ( \58839 , \58830 , \58837 , \58838 );
and \U$58463 ( \58840 , \58672 , \58839 );
and \U$58464 ( \58841 , \58451 , \58671 );
nor \U$58465 ( \58842 , \58840 , \58841 );
and \U$58466 ( \58843 , \58246 , \58450 );
xor \U$58467 ( \58844 , \58463 , \58488 );
and \U$58468 ( \58845 , \58844 , \58670 );
and \U$58469 ( \58846 , \58463 , \58488 );
or \U$58470 ( \58847 , \58845 , \58846 );
xnor \U$58471 ( \58848 , \58843 , \58847 );
not \U$58472 ( \58849 , \58848 );
xor \U$58473 ( \58850 , \57940 , \57947 );
xor \U$58474 ( \58851 , \58850 , \57955 );
and \U$58475 ( \58852 , \58482 , \58851 );
xor \U$58476 ( \58853 , \57940 , \57947 );
xor \U$58477 ( \58854 , \58853 , \57955 );
and \U$58478 ( \58855 , \58484 , \58854 );
and \U$58479 ( \58856 , \58482 , \58484 );
or \U$58480 ( \58857 , \58852 , \58855 , \58856 );
xor \U$58481 ( \58858 , \58304 , \58308 );
and \U$58482 ( \58859 , \58858 , \58313 );
and \U$58483 ( \58860 , \58304 , \58308 );
or \U$58484 ( \58861 , \58859 , \58860 );
xor \U$58485 ( \58862 , \58857 , \58861 );
xor \U$58486 ( \58863 , \58467 , \58472 );
and \U$58487 ( \58864 , \58863 , \58475 );
and \U$58488 ( \58865 , \58467 , \58472 );
or \U$58489 ( \58866 , \58864 , \58865 );
xor \U$58490 ( \58867 , \58862 , \58866 );
not \U$58491 ( \58868 , \58867 );
xor \U$58492 ( \58869 , \57684 , \57691 );
xor \U$58493 ( \58870 , \58869 , \57699 );
not \U$58494 ( \58871 , \57931 );
not \U$58495 ( \58872 , \57902 );
or \U$58496 ( \58873 , \58871 , \58872 );
or \U$58497 ( \58874 , \57902 , \57931 );
nand \U$58498 ( \58875 , \58873 , \58874 );
not \U$58499 ( \58876 , \58875 );
not \U$58500 ( \58877 , \57877 );
and \U$58501 ( \58878 , \58876 , \58877 );
and \U$58502 ( \58879 , \58875 , \57877 );
nor \U$58503 ( \58880 , \58878 , \58879 );
xor \U$58504 ( \58881 , \58870 , \58880 );
not \U$58505 ( \58882 , \58018 );
not \U$58506 ( \58883 , \58024 );
or \U$58507 ( \58884 , \58882 , \58883 );
or \U$58508 ( \58885 , \58018 , \58024 );
nand \U$58509 ( \58886 , \58884 , \58885 );
not \U$58510 ( \58887 , \58886 );
not \U$58511 ( \58888 , \58016 );
and \U$58512 ( \58889 , \58887 , \58888 );
and \U$58513 ( \58890 , \58886 , \58016 );
nor \U$58514 ( \58891 , \58889 , \58890 );
xor \U$58515 ( \58892 , \58881 , \58891 );
not \U$58516 ( \58893 , \58892 );
or \U$58517 ( \58894 , \58868 , \58893 );
or \U$58518 ( \58895 , \58892 , \58867 );
nand \U$58519 ( \58896 , \58894 , \58895 );
xor \U$58520 ( \58897 , \58300 , \58314 );
and \U$58521 ( \58898 , \58897 , \58449 );
and \U$58522 ( \58899 , \58300 , \58314 );
or \U$58523 ( \58900 , \58898 , \58899 );
xor \U$58524 ( \58901 , \58896 , \58900 );
xor \U$58525 ( \58902 , \58126 , \58185 );
and \U$58526 ( \58903 , \58902 , \58245 );
and \U$58527 ( \58904 , \58126 , \58185 );
or \U$58528 ( \58905 , \58903 , \58904 );
xor \U$58529 ( \58906 , \57958 , \57976 );
xor \U$58530 ( \58907 , \58906 , \58002 );
xor \U$58531 ( \58908 , \58905 , \58907 );
xor \U$58532 ( \58909 , \58467 , \58472 );
xor \U$58533 ( \58910 , \58909 , \58475 );
and \U$58534 ( \58911 , \58478 , \58910 );
xor \U$58535 ( \58912 , \58467 , \58472 );
xor \U$58536 ( \58913 , \58912 , \58475 );
and \U$58537 ( \58914 , \58486 , \58913 );
and \U$58538 ( \58915 , \58478 , \58486 );
or \U$58539 ( \58916 , \58911 , \58914 , \58915 );
xor \U$58540 ( \58917 , \58908 , \58916 );
xor \U$58541 ( \58918 , \58901 , \58917 );
not \U$58542 ( \58919 , \58918 );
and \U$58543 ( \58920 , \58849 , \58919 );
and \U$58544 ( \58921 , \58848 , \58918 );
nor \U$58545 ( \58922 , \58920 , \58921 );
or \U$58546 ( \58923 , \58842 , \58922 );
xnor \U$58547 ( \58924 , \58922 , \58842 );
xor \U$58548 ( \58925 , \58650 , \58652 );
xor \U$58549 ( \58926 , \58925 , \58667 );
xor \U$58550 ( \58927 , \58827 , \58834 );
xor \U$58551 ( \58928 , \58926 , \58927 );
not \U$58552 ( \58929 , \58928 );
xor \U$58553 ( \58930 , \58561 , \58612 );
xor \U$58554 ( \58931 , \58930 , \58647 );
not \U$58555 ( \58932 , \58931 );
xor \U$58556 ( \58933 , \58674 , \58680 );
xor \U$58557 ( \58934 , \58933 , \58683 );
not \U$58558 ( \58935 , \58934 );
xor \U$58559 ( \58936 , \58728 , \58809 );
xor \U$58560 ( \58937 , \58936 , \58822 );
nand \U$58561 ( \58938 , \58935 , \58937 );
nand \U$58562 ( \58939 , \58932 , \58938 );
and \U$58563 ( \58940 , \15726 , RIae78620_114);
and \U$58564 ( \58941 , RIae78440_110, RIae7aab0_192);
nor \U$58565 ( \58942 , \58940 , \58941 );
and \U$58566 ( \58943 , \58942 , \14959 );
not \U$58567 ( \58944 , \58942 );
and \U$58568 ( \58945 , \58944 , RIae7aa38_191);
nor \U$58569 ( \58946 , \58943 , \58945 );
xor \U$58570 ( \58947 , \58946 , \6945 );
and \U$58571 ( \58948 , \14964 , RIae78080_102);
and \U$58572 ( \58949 , RIae78260_106, \14962 );
nor \U$58573 ( \58950 , \58948 , \58949 );
and \U$58574 ( \58951 , \58950 , \14463 );
not \U$58575 ( \58952 , \58950 );
and \U$58576 ( \58953 , \58952 , \14462 );
nor \U$58577 ( \58954 , \58951 , \58953 );
and \U$58578 ( \58955 , \58947 , \58954 );
and \U$58579 ( \58956 , \58946 , \6945 );
or \U$58580 ( \58957 , \58955 , \58956 );
and \U$58581 ( \58958 , \13059 , RIae77360_74);
and \U$58582 ( \58959 , RIae78350_108, \13057 );
nor \U$58583 ( \58960 , \58958 , \58959 );
and \U$58584 ( \58961 , \58960 , \13063 );
not \U$58585 ( \58962 , \58960 );
and \U$58586 ( \58963 , \58962 , \12718 );
nor \U$58587 ( \58964 , \58961 , \58963 );
and \U$58588 ( \58965 , \12180 , RIae77090_68);
and \U$58589 ( \58966 , RIae77270_72, \12178 );
nor \U$58590 ( \58967 , \58965 , \58966 );
and \U$58591 ( \58968 , \58967 , \12184 );
not \U$58592 ( \58969 , \58967 );
and \U$58593 ( \58970 , \58969 , \11827 );
nor \U$58594 ( \58971 , \58968 , \58970 );
xor \U$58595 ( \58972 , \58964 , \58971 );
and \U$58596 ( \58973 , \14059 , RIae78170_104);
and \U$58597 ( \58974 , RIae77f90_100, \14057 );
nor \U$58598 ( \58975 , \58973 , \58974 );
and \U$58599 ( \58976 , \58975 , \13502 );
not \U$58600 ( \58977 , \58975 );
and \U$58601 ( \58978 , \58977 , \14063 );
nor \U$58602 ( \58979 , \58976 , \58978 );
and \U$58603 ( \58980 , \58972 , \58979 );
and \U$58604 ( \58981 , \58964 , \58971 );
or \U$58605 ( \58982 , \58980 , \58981 );
xor \U$58606 ( \58983 , \58957 , \58982 );
and \U$58607 ( \58984 , \11470 , RIae76cd0_60);
and \U$58608 ( \58985 , RIae77108_69, \11468 );
nor \U$58609 ( \58986 , \58984 , \58985 );
and \U$58610 ( \58987 , \58986 , \10936 );
not \U$58611 ( \58988 , \58986 );
and \U$58612 ( \58989 , \58988 , \11474 );
nor \U$58613 ( \58990 , \58987 , \58989 );
and \U$58614 ( \58991 , \9760 , RIae77900_86);
and \U$58615 ( \58992 , RIae76fa0_66, \9758 );
nor \U$58616 ( \58993 , \58991 , \58992 );
and \U$58617 ( \58994 , \58993 , \9273 );
not \U$58618 ( \58995 , \58993 );
and \U$58619 ( \58996 , \58995 , \9272 );
nor \U$58620 ( \58997 , \58994 , \58996 );
xor \U$58621 ( \58998 , \58990 , \58997 );
and \U$58622 ( \58999 , \10548 , RIae76eb0_64);
and \U$58623 ( \59000 , RIae76dc0_62, \10546 );
nor \U$58624 ( \59001 , \58999 , \59000 );
and \U$58625 ( \59002 , \59001 , \10421 );
not \U$58626 ( \59003 , \59001 );
and \U$58627 ( \59004 , \59003 , \10118 );
nor \U$58628 ( \59005 , \59002 , \59004 );
and \U$58629 ( \59006 , \58998 , \59005 );
and \U$58630 ( \59007 , \58990 , \58997 );
or \U$58631 ( \59008 , \59006 , \59007 );
and \U$58632 ( \59009 , \58983 , \59008 );
and \U$58633 ( \59010 , \58957 , \58982 );
nor \U$58634 ( \59011 , \59009 , \59010 );
not \U$58635 ( \59012 , \59011 );
xor \U$58636 ( \59013 , \58762 , \58769 );
xor \U$58637 ( \59014 , \59013 , \58777 );
not \U$58638 ( \59015 , \59014 );
xor \U$58639 ( \59016 , \58788 , \58795 );
xor \U$58640 ( \59017 , \59016 , \58803 );
nand \U$58641 ( \59018 , \59015 , \59017 );
not \U$58642 ( \59019 , \59018 );
and \U$58643 ( \59020 , \59012 , \59019 );
and \U$58644 ( \59021 , \59011 , \59018 );
not \U$58645 ( \59022 , \58708 );
not \U$58646 ( \59023 , \58719 );
or \U$58647 ( \59024 , \59022 , \59023 );
or \U$58648 ( \59025 , \58708 , \58719 );
nand \U$58649 ( \59026 , \59024 , \59025 );
not \U$58650 ( \59027 , \59026 );
not \U$58651 ( \59028 , \58701 );
and \U$58652 ( \59029 , \59027 , \59028 );
and \U$58653 ( \59030 , \59026 , \58701 );
nor \U$58654 ( \59031 , \59029 , \59030 );
not \U$58655 ( \59032 , \59031 );
not \U$58656 ( \59033 , \58742 );
not \U$58657 ( \59034 , \58753 );
or \U$58658 ( \59035 , \59033 , \59034 );
or \U$58659 ( \59036 , \58742 , \58753 );
nand \U$58660 ( \59037 , \59035 , \59036 );
not \U$58661 ( \59038 , \59037 );
not \U$58662 ( \59039 , \58735 );
and \U$58663 ( \59040 , \59038 , \59039 );
and \U$58664 ( \59041 , \59037 , \58735 );
nor \U$58665 ( \59042 , \59040 , \59041 );
not \U$58666 ( \59043 , \59042 );
and \U$58667 ( \59044 , \59032 , \59043 );
and \U$58668 ( \59045 , \59042 , \59031 );
and \U$58669 ( \59046 , \7633 , RIae77540_78);
and \U$58670 ( \59047 , RIae776a8_81, \7631 );
nor \U$58671 ( \59048 , \59046 , \59047 );
and \U$58672 ( \59049 , \59048 , \7205 );
not \U$58673 ( \59050 , \59048 );
and \U$58674 ( \59051 , \59050 , \7206 );
nor \U$58675 ( \59052 , \59049 , \59051 );
not \U$58676 ( \59053 , \59052 );
and \U$58677 ( \59054 , \8371 , RIae77450_76);
and \U$58678 ( \59055 , RIae77ae0_90, \8369 );
nor \U$58679 ( \59056 , \59054 , \59055 );
and \U$58680 ( \59057 , \59056 , \8019 );
not \U$58681 ( \59058 , \59056 );
and \U$58682 ( \59059 , \59058 , \8020 );
nor \U$58683 ( \59060 , \59057 , \59059 );
not \U$58684 ( \59061 , \59060 );
and \U$58685 ( \59062 , \59053 , \59061 );
and \U$58686 ( \59063 , \59060 , \59052 );
and \U$58687 ( \59064 , \8966 , RIae779f0_88);
and \U$58688 ( \59065 , RIae77810_84, \8964 );
nor \U$58689 ( \59066 , \59064 , \59065 );
and \U$58690 ( \59067 , \59066 , \8789 );
not \U$58691 ( \59068 , \59066 );
and \U$58692 ( \59069 , \59068 , \8799 );
nor \U$58693 ( \59070 , \59067 , \59069 );
nor \U$58694 ( \59071 , \59063 , \59070 );
nor \U$58695 ( \59072 , \59062 , \59071 );
nor \U$58696 ( \59073 , \59045 , \59072 );
nor \U$58697 ( \59074 , \59044 , \59073 );
nor \U$58698 ( \59075 , \59021 , \59074 );
nor \U$58699 ( \59076 , \59020 , \59075 );
xor \U$58700 ( \59077 , \58514 , \58532 );
xor \U$58701 ( \59078 , \59077 , \58558 );
not \U$58702 ( \59079 , \59078 );
or \U$58703 ( \59080 , \59076 , \59079 );
not \U$58704 ( \59081 , \59079 );
not \U$58705 ( \59082 , \59076 );
or \U$58706 ( \59083 , \59081 , \59082 );
xor \U$58707 ( \59084 , \58755 , \58780 );
xor \U$58708 ( \59085 , \59084 , \58806 );
xor \U$58709 ( \59086 , \58721 , \58722 );
xor \U$58710 ( \59087 , \59086 , \58725 );
and \U$58711 ( \59088 , \59085 , \59087 );
xor \U$58712 ( \59089 , \58496 , \58503 );
xor \U$58713 ( \59090 , \59089 , \58511 );
xor \U$58714 ( \59091 , \58812 , \58817 );
xor \U$58715 ( \59092 , \59090 , \59091 );
xor \U$58716 ( \59093 , \58721 , \58722 );
xor \U$58717 ( \59094 , \59093 , \58725 );
and \U$58718 ( \59095 , \59092 , \59094 );
and \U$58719 ( \59096 , \59085 , \59092 );
or \U$58720 ( \59097 , \59088 , \59095 , \59096 );
nand \U$58721 ( \59098 , \59083 , \59097 );
nand \U$58722 ( \59099 , \59080 , \59098 );
and \U$58723 ( \59100 , \58939 , \59099 );
not \U$58724 ( \59101 , \58938 );
and \U$58725 ( \59102 , \58931 , \59101 );
nor \U$58726 ( \59103 , \59100 , \59102 );
not \U$58727 ( \59104 , \59103 );
and \U$58728 ( \59105 , \58929 , \59104 );
and \U$58729 ( \59106 , \58928 , \59103 );
nor \U$58730 ( \59107 , \59105 , \59106 );
xnor \U$58731 ( \59108 , \58686 , \58825 );
not \U$58732 ( \59109 , \59108 );
not \U$58733 ( \59110 , \58691 );
and \U$58734 ( \59111 , \59109 , \59110 );
and \U$58735 ( \59112 , \59108 , \58691 );
nor \U$58736 ( \59113 , \59111 , \59112 );
not \U$58737 ( \59114 , \59113 );
not \U$58738 ( \59115 , \58931 );
not \U$58739 ( \59116 , \59099 );
not \U$58740 ( \59117 , \58938 );
and \U$58741 ( \59118 , \59116 , \59117 );
and \U$58742 ( \59119 , \59099 , \58938 );
nor \U$58743 ( \59120 , \59118 , \59119 );
not \U$58744 ( \59121 , \59120 );
or \U$58745 ( \59122 , \59115 , \59121 );
or \U$58746 ( \59123 , \59120 , \58931 );
nand \U$58747 ( \59124 , \59122 , \59123 );
nand \U$58748 ( \59125 , \59114 , \59124 );
or \U$58749 ( \59126 , \59107 , \59125 );
xnor \U$58750 ( \59127 , \59125 , \59107 );
xor \U$58751 ( \59128 , \58957 , \58982 );
xor \U$58752 ( \59129 , \59128 , \59008 );
not \U$58753 ( \59130 , \59017 );
not \U$58754 ( \59131 , \59014 );
or \U$58755 ( \59132 , \59130 , \59131 );
or \U$58756 ( \59133 , \59014 , \59017 );
nand \U$58757 ( \59134 , \59132 , \59133 );
xor \U$58758 ( \59135 , \59129 , \59134 );
not \U$58759 ( \59136 , \59031 );
xor \U$58760 ( \59137 , \59072 , \59042 );
not \U$58761 ( \59138 , \59137 );
or \U$58762 ( \59139 , \59136 , \59138 );
or \U$58763 ( \59140 , \59137 , \59031 );
nand \U$58764 ( \59141 , \59139 , \59140 );
and \U$58765 ( \59142 , \59135 , \59141 );
and \U$58766 ( \59143 , \59129 , \59134 );
or \U$58767 ( \59144 , \59142 , \59143 );
and \U$58768 ( \59145 , \8966 , RIae77ae0_90);
and \U$58769 ( \59146 , RIae779f0_88, \8964 );
nor \U$58770 ( \59147 , \59145 , \59146 );
and \U$58771 ( \59148 , \59147 , \8799 );
not \U$58772 ( \59149 , \59147 );
and \U$58773 ( \59150 , \59149 , \8789 );
nor \U$58774 ( \59151 , \59148 , \59150 );
and \U$58775 ( \59152 , \9760 , RIae77810_84);
and \U$58776 ( \59153 , RIae77900_86, \9758 );
nor \U$58777 ( \59154 , \59152 , \59153 );
and \U$58778 ( \59155 , \59154 , \9273 );
not \U$58779 ( \59156 , \59154 );
and \U$58780 ( \59157 , \59156 , \9764 );
nor \U$58781 ( \59158 , \59155 , \59157 );
xor \U$58782 ( \59159 , \59151 , \59158 );
and \U$58783 ( \59160 , \10548 , RIae76fa0_66);
and \U$58784 ( \59161 , RIae76eb0_64, \10546 );
nor \U$58785 ( \59162 , \59160 , \59161 );
and \U$58786 ( \59163 , \59162 , \10421 );
not \U$58787 ( \59164 , \59162 );
and \U$58788 ( \59165 , \59164 , \10118 );
nor \U$58789 ( \59166 , \59163 , \59165 );
and \U$58790 ( \59167 , \59159 , \59166 );
and \U$58791 ( \59168 , \59151 , \59158 );
or \U$58792 ( \59169 , \59167 , \59168 );
and \U$58793 ( \59170 , \14964 , RIae77f90_100);
and \U$58794 ( \59171 , RIae78080_102, \14962 );
nor \U$58795 ( \59172 , \59170 , \59171 );
and \U$58796 ( \59173 , \59172 , \14463 );
not \U$58797 ( \59174 , \59172 );
and \U$58798 ( \59175 , \59174 , \14462 );
nor \U$58799 ( \59176 , \59173 , \59175 );
and \U$58800 ( \59177 , \15726 , RIae78260_106);
and \U$58801 ( \59178 , RIae78620_114, RIae7aab0_192);
nor \U$58802 ( \59179 , \59177 , \59178 );
and \U$58803 ( \59180 , \59179 , \14959 );
not \U$58804 ( \59181 , \59179 );
and \U$58805 ( \59182 , \59181 , RIae7aa38_191);
nor \U$58806 ( \59183 , \59180 , \59182 );
xor \U$58807 ( \59184 , \59176 , \59183 );
and \U$58808 ( \59185 , \14059 , RIae78350_108);
and \U$58809 ( \59186 , RIae78170_104, \14057 );
nor \U$58810 ( \59187 , \59185 , \59186 );
and \U$58811 ( \59188 , \59187 , \13502 );
not \U$58812 ( \59189 , \59187 );
and \U$58813 ( \59190 , \59189 , \14063 );
nor \U$58814 ( \59191 , \59188 , \59190 );
and \U$58815 ( \59192 , \59184 , \59191 );
and \U$58816 ( \59193 , \59176 , \59183 );
or \U$58817 ( \59194 , \59192 , \59193 );
xor \U$58818 ( \59195 , \59169 , \59194 );
and \U$58819 ( \59196 , \11470 , RIae76dc0_62);
and \U$58820 ( \59197 , RIae76cd0_60, \11468 );
nor \U$58821 ( \59198 , \59196 , \59197 );
and \U$58822 ( \59199 , \59198 , \10936 );
not \U$58823 ( \59200 , \59198 );
and \U$58824 ( \59201 , \59200 , \11474 );
nor \U$58825 ( \59202 , \59199 , \59201 );
and \U$58826 ( \59203 , \12180 , RIae77108_69);
and \U$58827 ( \59204 , RIae77090_68, \12178 );
nor \U$58828 ( \59205 , \59203 , \59204 );
and \U$58829 ( \59206 , \59205 , \12184 );
not \U$58830 ( \59207 , \59205 );
and \U$58831 ( \59208 , \59207 , \11827 );
nor \U$58832 ( \59209 , \59206 , \59208 );
xor \U$58833 ( \59210 , \59202 , \59209 );
and \U$58834 ( \59211 , \13059 , RIae77270_72);
and \U$58835 ( \59212 , RIae77360_74, \13057 );
nor \U$58836 ( \59213 , \59211 , \59212 );
and \U$58837 ( \59214 , \59213 , \13063 );
not \U$58838 ( \59215 , \59213 );
and \U$58839 ( \59216 , \59215 , \12718 );
nor \U$58840 ( \59217 , \59214 , \59216 );
and \U$58841 ( \59218 , \59210 , \59217 );
and \U$58842 ( \59219 , \59202 , \59209 );
or \U$58843 ( \59220 , \59218 , \59219 );
and \U$58844 ( \59221 , \59195 , \59220 );
and \U$58845 ( \59222 , \59169 , \59194 );
or \U$58846 ( \59223 , \59221 , \59222 );
xor \U$58847 ( \59224 , \58964 , \58971 );
xor \U$58848 ( \59225 , \59224 , \58979 );
xor \U$58849 ( \59226 , \58946 , \6945 );
xor \U$58850 ( \59227 , \59226 , \58954 );
and \U$58851 ( \59228 , \59225 , \59227 );
xor \U$58852 ( \59229 , \59223 , \59228 );
nand \U$58853 ( \59230 , RIae77630_80, \6939 );
and \U$58854 ( \59231 , \59230 , \6314 );
not \U$58855 ( \59232 , \59230 );
and \U$58856 ( \59233 , \59232 , \6945 );
nor \U$58857 ( \59234 , \59231 , \59233 );
xor \U$58858 ( \59235 , \58990 , \58997 );
xor \U$58859 ( \59236 , \59235 , \59005 );
and \U$58860 ( \59237 , \59234 , \59236 );
not \U$58861 ( \59238 , \59052 );
xor \U$58862 ( \59239 , \59060 , \59070 );
not \U$58863 ( \59240 , \59239 );
or \U$58864 ( \59241 , \59238 , \59240 );
or \U$58865 ( \59242 , \59239 , \59052 );
nand \U$58866 ( \59243 , \59241 , \59242 );
xor \U$58867 ( \59244 , \58990 , \58997 );
xor \U$58868 ( \59245 , \59244 , \59005 );
and \U$58869 ( \59246 , \59243 , \59245 );
and \U$58870 ( \59247 , \59234 , \59243 );
or \U$58871 ( \59248 , \59237 , \59246 , \59247 );
and \U$58872 ( \59249 , \59229 , \59248 );
and \U$58873 ( \59250 , \59223 , \59228 );
or \U$58874 ( \59251 , \59249 , \59250 );
xor \U$58875 ( \59252 , \59144 , \59251 );
xor \U$58876 ( \59253 , \58721 , \58722 );
xor \U$58877 ( \59254 , \59253 , \58725 );
xor \U$58878 ( \59255 , \59085 , \59092 );
xor \U$58879 ( \59256 , \59254 , \59255 );
and \U$58880 ( \59257 , \59252 , \59256 );
and \U$58881 ( \59258 , \59144 , \59251 );
or \U$58882 ( \59259 , \59257 , \59258 );
not \U$58883 ( \59260 , \59259 );
not \U$58884 ( \59261 , \59097 );
not \U$58885 ( \59262 , \59076 );
and \U$58886 ( \59263 , \59261 , \59262 );
and \U$58887 ( \59264 , \59097 , \59076 );
nor \U$58888 ( \59265 , \59263 , \59264 );
not \U$58889 ( \59266 , \59265 );
not \U$58890 ( \59267 , \59078 );
and \U$58891 ( \59268 , \59266 , \59267 );
and \U$58892 ( \59269 , \59265 , \59078 );
nor \U$58893 ( \59270 , \59268 , \59269 );
not \U$58894 ( \59271 , \59270 );
or \U$58895 ( \59272 , \59260 , \59271 );
or \U$58896 ( \59273 , \59270 , \59259 );
nand \U$58897 ( \59274 , \59272 , \59273 );
not \U$58898 ( \59275 , \59274 );
not \U$58899 ( \59276 , \58937 );
not \U$58900 ( \59277 , \58934 );
and \U$58901 ( \59278 , \59276 , \59277 );
and \U$58902 ( \59279 , \58937 , \58934 );
nor \U$58903 ( \59280 , \59278 , \59279 );
not \U$58904 ( \59281 , \59280 );
and \U$58905 ( \59282 , \59275 , \59281 );
and \U$58906 ( \59283 , \59274 , \59280 );
nor \U$58907 ( \59284 , \59282 , \59283 );
xor \U$58908 ( \59285 , \59144 , \59251 );
xor \U$58909 ( \59286 , \59285 , \59256 );
not \U$58910 ( \59287 , \59018 );
xor \U$58911 ( \59288 , \59011 , \59074 );
not \U$58912 ( \59289 , \59288 );
or \U$58913 ( \59290 , \59287 , \59289 );
or \U$58914 ( \59291 , \59288 , \59018 );
nand \U$58915 ( \59292 , \59290 , \59291 );
xor \U$58916 ( \59293 , \59286 , \59292 );
xor \U$58917 ( \59294 , \59225 , \59227 );
xor \U$58918 ( \59295 , \59169 , \59194 );
xor \U$58919 ( \59296 , \59295 , \59220 );
and \U$58920 ( \59297 , \59294 , \59296 );
xor \U$58921 ( \59298 , \58990 , \58997 );
xor \U$58922 ( \59299 , \59298 , \59005 );
xor \U$58923 ( \59300 , \59234 , \59243 );
xor \U$58924 ( \59301 , \59299 , \59300 );
xor \U$58925 ( \59302 , \59169 , \59194 );
xor \U$58926 ( \59303 , \59302 , \59220 );
and \U$58927 ( \59304 , \59301 , \59303 );
and \U$58928 ( \59305 , \59294 , \59301 );
or \U$58929 ( \59306 , \59297 , \59304 , \59305 );
and \U$58930 ( \59307 , \14059 , RIae77360_74);
and \U$58931 ( \59308 , RIae78350_108, \14057 );
nor \U$58932 ( \59309 , \59307 , \59308 );
and \U$58933 ( \59310 , \59309 , \13502 );
not \U$58934 ( \59311 , \59309 );
and \U$58935 ( \59312 , \59311 , \14063 );
nor \U$58936 ( \59313 , \59310 , \59312 );
and \U$58937 ( \59314 , \12180 , RIae76cd0_60);
and \U$58938 ( \59315 , RIae77108_69, \12178 );
nor \U$58939 ( \59316 , \59314 , \59315 );
and \U$58940 ( \59317 , \59316 , \12184 );
not \U$58941 ( \59318 , \59316 );
and \U$58942 ( \59319 , \59318 , \11827 );
nor \U$58943 ( \59320 , \59317 , \59319 );
xor \U$58944 ( \59321 , \59313 , \59320 );
and \U$58945 ( \59322 , \13059 , RIae77090_68);
and \U$58946 ( \59323 , RIae77270_72, \13057 );
nor \U$58947 ( \59324 , \59322 , \59323 );
and \U$58948 ( \59325 , \59324 , \13063 );
not \U$58949 ( \59326 , \59324 );
and \U$58950 ( \59327 , \59326 , \12718 );
nor \U$58951 ( \59328 , \59325 , \59327 );
and \U$58952 ( \59329 , \59321 , \59328 );
and \U$58953 ( \59330 , \59313 , \59320 );
or \U$58954 ( \59331 , \59329 , \59330 );
and \U$58955 ( \59332 , \15726 , RIae78080_102);
and \U$58956 ( \59333 , RIae78260_106, RIae7aab0_192);
nor \U$58957 ( \59334 , \59332 , \59333 );
and \U$58958 ( \59335 , \59334 , \14959 );
not \U$58959 ( \59336 , \59334 );
and \U$58960 ( \59337 , \59336 , RIae7aa38_191);
nor \U$58961 ( \59338 , \59335 , \59337 );
xor \U$58962 ( \59339 , \59338 , \7205 );
and \U$58963 ( \59340 , \14964 , RIae78170_104);
and \U$58964 ( \59341 , RIae77f90_100, \14962 );
nor \U$58965 ( \59342 , \59340 , \59341 );
and \U$58966 ( \59343 , \59342 , \14463 );
not \U$58967 ( \59344 , \59342 );
and \U$58968 ( \59345 , \59344 , \14462 );
nor \U$58969 ( \59346 , \59343 , \59345 );
and \U$58970 ( \59347 , \59339 , \59346 );
and \U$58971 ( \59348 , \59338 , \7205 );
or \U$58972 ( \59349 , \59347 , \59348 );
xor \U$58973 ( \59350 , \59331 , \59349 );
and \U$58974 ( \59351 , \11470 , RIae76eb0_64);
and \U$58975 ( \59352 , RIae76dc0_62, \11468 );
nor \U$58976 ( \59353 , \59351 , \59352 );
and \U$58977 ( \59354 , \59353 , \10936 );
not \U$58978 ( \59355 , \59353 );
and \U$58979 ( \59356 , \59355 , \11474 );
nor \U$58980 ( \59357 , \59354 , \59356 );
and \U$58981 ( \59358 , \9760 , RIae779f0_88);
and \U$58982 ( \59359 , RIae77810_84, \9758 );
nor \U$58983 ( \59360 , \59358 , \59359 );
and \U$58984 ( \59361 , \59360 , \9273 );
not \U$58985 ( \59362 , \59360 );
and \U$58986 ( \59363 , \59362 , \9272 );
nor \U$58987 ( \59364 , \59361 , \59363 );
xor \U$58988 ( \59365 , \59357 , \59364 );
and \U$58989 ( \59366 , \10548 , RIae77900_86);
and \U$58990 ( \59367 , RIae76fa0_66, \10546 );
nor \U$58991 ( \59368 , \59366 , \59367 );
and \U$58992 ( \59369 , \59368 , \10421 );
not \U$58993 ( \59370 , \59368 );
and \U$58994 ( \59371 , \59370 , \10118 );
nor \U$58995 ( \59372 , \59369 , \59371 );
and \U$58996 ( \59373 , \59365 , \59372 );
and \U$58997 ( \59374 , \59357 , \59364 );
or \U$58998 ( \59375 , \59373 , \59374 );
and \U$58999 ( \59376 , \59350 , \59375 );
and \U$59000 ( \59377 , \59331 , \59349 );
or \U$59001 ( \59378 , \59376 , \59377 );
and \U$59002 ( \59379 , \8371 , RIae776a8_81);
and \U$59003 ( \59380 , RIae77450_76, \8369 );
nor \U$59004 ( \59381 , \59379 , \59380 );
and \U$59005 ( \59382 , \59381 , \8020 );
not \U$59006 ( \59383 , \59381 );
and \U$59007 ( \59384 , \59383 , \8019 );
nor \U$59008 ( \59385 , \59382 , \59384 );
and \U$59009 ( \59386 , \7633 , RIae77630_80);
and \U$59010 ( \59387 , RIae77540_78, \7631 );
nor \U$59011 ( \59388 , \59386 , \59387 );
and \U$59012 ( \59389 , \59388 , \7206 );
not \U$59013 ( \59390 , \59388 );
and \U$59014 ( \59391 , \59390 , \7205 );
nor \U$59015 ( \59392 , \59389 , \59391 );
xor \U$59016 ( \59393 , \59385 , \59392 );
and \U$59017 ( \59394 , \8966 , RIae77450_76);
and \U$59018 ( \59395 , RIae77ae0_90, \8964 );
nor \U$59019 ( \59396 , \59394 , \59395 );
and \U$59020 ( \59397 , \59396 , \8799 );
not \U$59021 ( \59398 , \59396 );
and \U$59022 ( \59399 , \59398 , \8789 );
nor \U$59023 ( \59400 , \59397 , \59399 );
nand \U$59024 ( \59401 , RIae77630_80, \7631 );
and \U$59025 ( \59402 , \59401 , \7206 );
not \U$59026 ( \59403 , \59401 );
and \U$59027 ( \59404 , \59403 , \7205 );
nor \U$59028 ( \59405 , \59402 , \59404 );
xor \U$59029 ( \59406 , \59400 , \59405 );
and \U$59030 ( \59407 , \8371 , RIae77540_78);
and \U$59031 ( \59408 , RIae776a8_81, \8369 );
nor \U$59032 ( \59409 , \59407 , \59408 );
and \U$59033 ( \59410 , \59409 , \8020 );
not \U$59034 ( \59411 , \59409 );
and \U$59035 ( \59412 , \59411 , \8019 );
nor \U$59036 ( \59413 , \59410 , \59412 );
and \U$59037 ( \59414 , \59406 , \59413 );
and \U$59038 ( \59415 , \59400 , \59405 );
or \U$59039 ( \59416 , \59414 , \59415 );
and \U$59040 ( \59417 , \59393 , \59416 );
and \U$59041 ( \59418 , \59385 , \59392 );
or \U$59042 ( \59419 , \59417 , \59418 );
xor \U$59043 ( \59420 , \59378 , \59419 );
xor \U$59044 ( \59421 , \59176 , \59183 );
xor \U$59045 ( \59422 , \59421 , \59191 );
xor \U$59046 ( \59423 , \59151 , \59158 );
xor \U$59047 ( \59424 , \59423 , \59166 );
and \U$59048 ( \59425 , \59422 , \59424 );
xor \U$59049 ( \59426 , \59202 , \59209 );
xor \U$59050 ( \59427 , \59426 , \59217 );
xor \U$59051 ( \59428 , \59151 , \59158 );
xor \U$59052 ( \59429 , \59428 , \59166 );
and \U$59053 ( \59430 , \59427 , \59429 );
and \U$59054 ( \59431 , \59422 , \59427 );
or \U$59055 ( \59432 , \59425 , \59430 , \59431 );
and \U$59056 ( \59433 , \59420 , \59432 );
and \U$59057 ( \59434 , \59378 , \59419 );
or \U$59058 ( \59435 , \59433 , \59434 );
xor \U$59059 ( \59436 , \59306 , \59435 );
xor \U$59060 ( \59437 , \59129 , \59134 );
xor \U$59061 ( \59438 , \59437 , \59141 );
and \U$59062 ( \59439 , \59436 , \59438 );
and \U$59063 ( \59440 , \59306 , \59435 );
or \U$59064 ( \59441 , \59439 , \59440 );
and \U$59065 ( \59442 , \59293 , \59441 );
and \U$59066 ( \59443 , \59286 , \59292 );
nor \U$59067 ( \59444 , \59442 , \59443 );
or \U$59068 ( \59445 , \59284 , \59444 );
xnor \U$59069 ( \59446 , \59444 , \59284 );
xor \U$59070 ( \59447 , \59286 , \59292 );
xor \U$59071 ( \59448 , \59447 , \59441 );
xor \U$59072 ( \59449 , \59223 , \59228 );
xor \U$59073 ( \59450 , \59449 , \59248 );
not \U$59074 ( \59451 , \59450 );
xor \U$59075 ( \59452 , \59306 , \59435 );
xor \U$59076 ( \59453 , \59452 , \59438 );
not \U$59077 ( \59454 , \59453 );
or \U$59078 ( \59455 , \59451 , \59454 );
or \U$59079 ( \59456 , \59453 , \59450 );
xor \U$59080 ( \59457 , \59400 , \59405 );
xor \U$59081 ( \59458 , \59457 , \59413 );
xor \U$59082 ( \59459 , \59313 , \59320 );
xor \U$59083 ( \59460 , \59459 , \59328 );
and \U$59084 ( \59461 , \59458 , \59460 );
xor \U$59085 ( \59462 , \59357 , \59364 );
xor \U$59086 ( \59463 , \59462 , \59372 );
xor \U$59087 ( \59464 , \59313 , \59320 );
xor \U$59088 ( \59465 , \59464 , \59328 );
and \U$59089 ( \59466 , \59463 , \59465 );
and \U$59090 ( \59467 , \59458 , \59463 );
or \U$59091 ( \59468 , \59461 , \59466 , \59467 );
and \U$59092 ( \59469 , \12180 , RIae76dc0_62);
and \U$59093 ( \59470 , RIae76cd0_60, \12178 );
nor \U$59094 ( \59471 , \59469 , \59470 );
and \U$59095 ( \59472 , \59471 , \11827 );
not \U$59096 ( \59473 , \59471 );
and \U$59097 ( \59474 , \59473 , \12184 );
nor \U$59098 ( \59475 , \59472 , \59474 );
and \U$59099 ( \59476 , \13059 , RIae77108_69);
and \U$59100 ( \59477 , RIae77090_68, \13057 );
nor \U$59101 ( \59478 , \59476 , \59477 );
and \U$59102 ( \59479 , \59478 , \12718 );
not \U$59103 ( \59480 , \59478 );
and \U$59104 ( \59481 , \59480 , \13063 );
nor \U$59105 ( \59482 , \59479 , \59481 );
xor \U$59106 ( \59483 , \59475 , \59482 );
and \U$59107 ( \59484 , \11470 , RIae76fa0_66);
and \U$59108 ( \59485 , RIae76eb0_64, \11468 );
nor \U$59109 ( \59486 , \59484 , \59485 );
and \U$59110 ( \59487 , \59486 , \11474 );
not \U$59111 ( \59488 , \59486 );
and \U$59112 ( \59489 , \59488 , \10936 );
nor \U$59113 ( \59490 , \59487 , \59489 );
and \U$59114 ( \59491 , \59483 , \59490 );
and \U$59115 ( \59492 , \59475 , \59482 );
nor \U$59116 ( \59493 , \59491 , \59492 );
and \U$59117 ( \59494 , \14059 , RIae77270_72);
and \U$59118 ( \59495 , RIae77360_74, \14057 );
nor \U$59119 ( \59496 , \59494 , \59495 );
and \U$59120 ( \59497 , \59496 , \13502 );
not \U$59121 ( \59498 , \59496 );
and \U$59122 ( \59499 , \59498 , \14063 );
nor \U$59123 ( \59500 , \59497 , \59499 );
and \U$59124 ( \59501 , \15726 , RIae77f90_100);
and \U$59125 ( \59502 , RIae78080_102, RIae7aab0_192);
nor \U$59126 ( \59503 , \59501 , \59502 );
and \U$59127 ( \59504 , \59503 , \14959 );
not \U$59128 ( \59505 , \59503 );
and \U$59129 ( \59506 , \59505 , RIae7aa38_191);
nor \U$59130 ( \59507 , \59504 , \59506 );
xor \U$59131 ( \59508 , \59500 , \59507 );
and \U$59132 ( \59509 , \14964 , RIae78350_108);
and \U$59133 ( \59510 , RIae78170_104, \14962 );
nor \U$59134 ( \59511 , \59509 , \59510 );
and \U$59135 ( \59512 , \59511 , \14463 );
not \U$59136 ( \59513 , \59511 );
and \U$59137 ( \59514 , \59513 , \14462 );
nor \U$59138 ( \59515 , \59512 , \59514 );
and \U$59139 ( \59516 , \59508 , \59515 );
and \U$59140 ( \59517 , \59500 , \59507 );
or \U$59141 ( \59518 , \59516 , \59517 );
xor \U$59142 ( \59519 , \59493 , \59518 );
and \U$59143 ( \59520 , \9760 , RIae77ae0_90);
and \U$59144 ( \59521 , RIae779f0_88, \9758 );
nor \U$59145 ( \59522 , \59520 , \59521 );
and \U$59146 ( \59523 , \59522 , \9272 );
not \U$59147 ( \59524 , \59522 );
and \U$59148 ( \59525 , \59524 , \9273 );
nor \U$59149 ( \59526 , \59523 , \59525 );
and \U$59150 ( \59527 , \10548 , RIae77810_84);
and \U$59151 ( \59528 , RIae77900_86, \10546 );
nor \U$59152 ( \59529 , \59527 , \59528 );
and \U$59153 ( \59530 , \59529 , \10118 );
not \U$59154 ( \59531 , \59529 );
and \U$59155 ( \59532 , \59531 , \10421 );
nor \U$59156 ( \59533 , \59530 , \59532 );
xor \U$59157 ( \59534 , \59526 , \59533 );
and \U$59158 ( \59535 , \8966 , RIae776a8_81);
and \U$59159 ( \59536 , RIae77450_76, \8964 );
nor \U$59160 ( \59537 , \59535 , \59536 );
and \U$59161 ( \59538 , \59537 , \8789 );
not \U$59162 ( \59539 , \59537 );
and \U$59163 ( \59540 , \59539 , \8799 );
nor \U$59164 ( \59541 , \59538 , \59540 );
and \U$59165 ( \59542 , \59534 , \59541 );
and \U$59166 ( \59543 , \59526 , \59533 );
nor \U$59167 ( \59544 , \59542 , \59543 );
and \U$59168 ( \59545 , \59519 , \59544 );
and \U$59169 ( \59546 , \59493 , \59518 );
or \U$59170 ( \59547 , \59545 , \59546 );
xor \U$59171 ( \59548 , \59468 , \59547 );
xor \U$59172 ( \59549 , \59151 , \59158 );
xor \U$59173 ( \59550 , \59549 , \59166 );
xor \U$59174 ( \59551 , \59422 , \59427 );
xor \U$59175 ( \59552 , \59550 , \59551 );
and \U$59176 ( \59553 , \59548 , \59552 );
and \U$59177 ( \59554 , \59468 , \59547 );
or \U$59178 ( \59555 , \59553 , \59554 );
xor \U$59179 ( \59556 , \59378 , \59419 );
xor \U$59180 ( \59557 , \59556 , \59432 );
and \U$59181 ( \59558 , \59555 , \59557 );
xor \U$59182 ( \59559 , \59169 , \59194 );
xor \U$59183 ( \59560 , \59559 , \59220 );
xor \U$59184 ( \59561 , \59294 , \59301 );
xor \U$59185 ( \59562 , \59560 , \59561 );
xor \U$59186 ( \59563 , \59378 , \59419 );
xor \U$59187 ( \59564 , \59563 , \59432 );
and \U$59188 ( \59565 , \59562 , \59564 );
and \U$59189 ( \59566 , \59555 , \59562 );
or \U$59190 ( \59567 , \59558 , \59565 , \59566 );
nand \U$59191 ( \59568 , \59456 , \59567 );
nand \U$59192 ( \59569 , \59455 , \59568 );
and \U$59193 ( \59570 , \59448 , \59569 );
xor \U$59194 ( \59571 , \59569 , \59448 );
xnor \U$59195 ( \59572 , \59450 , \59567 );
not \U$59196 ( \59573 , \59572 );
not \U$59197 ( \59574 , \59453 );
and \U$59198 ( \59575 , \59573 , \59574 );
and \U$59199 ( \59576 , \59572 , \59453 );
nor \U$59200 ( \59577 , \59575 , \59576 );
xor \U$59201 ( \59578 , \59378 , \59419 );
xor \U$59202 ( \59579 , \59578 , \59432 );
xor \U$59203 ( \59580 , \59555 , \59562 );
xor \U$59204 ( \59581 , \59579 , \59580 );
xor \U$59205 ( \59582 , \59493 , \59518 );
xor \U$59206 ( \59583 , \59582 , \59544 );
xor \U$59207 ( \59584 , \59313 , \59320 );
xor \U$59208 ( \59585 , \59584 , \59328 );
xor \U$59209 ( \59586 , \59458 , \59463 );
xor \U$59210 ( \59587 , \59585 , \59586 );
and \U$59211 ( \59588 , \59583 , \59587 );
xor \U$59212 ( \59589 , \59385 , \59392 );
xor \U$59213 ( \59590 , \59589 , \59416 );
xor \U$59214 ( \59591 , \59588 , \59590 );
and \U$59215 ( \59592 , \9760 , RIae77450_76);
and \U$59216 ( \59593 , RIae77ae0_90, \9758 );
nor \U$59217 ( \59594 , \59592 , \59593 );
and \U$59218 ( \59595 , \59594 , \9273 );
not \U$59219 ( \59596 , \59594 );
and \U$59220 ( \59597 , \59596 , \9272 );
nor \U$59221 ( \59598 , \59595 , \59597 );
and \U$59222 ( \59599 , \10548 , RIae779f0_88);
and \U$59223 ( \59600 , RIae77810_84, \10546 );
nor \U$59224 ( \59601 , \59599 , \59600 );
and \U$59225 ( \59602 , \59601 , \10421 );
not \U$59226 ( \59603 , \59601 );
and \U$59227 ( \59604 , \59603 , \10118 );
nor \U$59228 ( \59605 , \59602 , \59604 );
xor \U$59229 ( \59606 , \59598 , \59605 );
and \U$59230 ( \59607 , \11470 , RIae77900_86);
and \U$59231 ( \59608 , RIae76fa0_66, \11468 );
nor \U$59232 ( \59609 , \59607 , \59608 );
and \U$59233 ( \59610 , \59609 , \10936 );
not \U$59234 ( \59611 , \59609 );
and \U$59235 ( \59612 , \59611 , \11474 );
nor \U$59236 ( \59613 , \59610 , \59612 );
and \U$59237 ( \59614 , \59606 , \59613 );
and \U$59238 ( \59615 , \59598 , \59605 );
or \U$59239 ( \59616 , \59614 , \59615 );
and \U$59240 ( \59617 , \15726 , RIae78170_104);
and \U$59241 ( \59618 , RIae77f90_100, RIae7aab0_192);
nor \U$59242 ( \59619 , \59617 , \59618 );
and \U$59243 ( \59620 , \59619 , \14959 );
not \U$59244 ( \59621 , \59619 );
and \U$59245 ( \59622 , \59621 , RIae7aa38_191);
nor \U$59246 ( \59623 , \59620 , \59622 );
xor \U$59247 ( \59624 , \59623 , \8019 );
and \U$59248 ( \59625 , \14964 , RIae77360_74);
and \U$59249 ( \59626 , RIae78350_108, \14962 );
nor \U$59250 ( \59627 , \59625 , \59626 );
and \U$59251 ( \59628 , \59627 , \14463 );
not \U$59252 ( \59629 , \59627 );
and \U$59253 ( \59630 , \59629 , \14462 );
nor \U$59254 ( \59631 , \59628 , \59630 );
and \U$59255 ( \59632 , \59624 , \59631 );
and \U$59256 ( \59633 , \59623 , \8019 );
or \U$59257 ( \59634 , \59632 , \59633 );
xor \U$59258 ( \59635 , \59616 , \59634 );
and \U$59259 ( \59636 , \14059 , RIae77090_68);
and \U$59260 ( \59637 , RIae77270_72, \14057 );
nor \U$59261 ( \59638 , \59636 , \59637 );
and \U$59262 ( \59639 , \59638 , \13502 );
not \U$59263 ( \59640 , \59638 );
and \U$59264 ( \59641 , \59640 , \14063 );
nor \U$59265 ( \59642 , \59639 , \59641 );
and \U$59266 ( \59643 , \12180 , RIae76eb0_64);
and \U$59267 ( \59644 , RIae76dc0_62, \12178 );
nor \U$59268 ( \59645 , \59643 , \59644 );
and \U$59269 ( \59646 , \59645 , \12184 );
not \U$59270 ( \59647 , \59645 );
and \U$59271 ( \59648 , \59647 , \11827 );
nor \U$59272 ( \59649 , \59646 , \59648 );
xor \U$59273 ( \59650 , \59642 , \59649 );
and \U$59274 ( \59651 , \13059 , RIae76cd0_60);
and \U$59275 ( \59652 , RIae77108_69, \13057 );
nor \U$59276 ( \59653 , \59651 , \59652 );
and \U$59277 ( \59654 , \59653 , \13063 );
not \U$59278 ( \59655 , \59653 );
and \U$59279 ( \59656 , \59655 , \12718 );
nor \U$59280 ( \59657 , \59654 , \59656 );
and \U$59281 ( \59658 , \59650 , \59657 );
and \U$59282 ( \59659 , \59642 , \59649 );
or \U$59283 ( \59660 , \59658 , \59659 );
and \U$59284 ( \59661 , \59635 , \59660 );
and \U$59285 ( \59662 , \59616 , \59634 );
or \U$59286 ( \59663 , \59661 , \59662 );
xor \U$59287 ( \59664 , \59338 , \7205 );
xor \U$59288 ( \59665 , \59664 , \59346 );
xor \U$59289 ( \59666 , \59663 , \59665 );
and \U$59290 ( \59667 , \8371 , RIae77630_80);
and \U$59291 ( \59668 , RIae77540_78, \8369 );
nor \U$59292 ( \59669 , \59667 , \59668 );
and \U$59293 ( \59670 , \59669 , \8019 );
not \U$59294 ( \59671 , \59669 );
and \U$59295 ( \59672 , \59671 , \8020 );
nor \U$59296 ( \59673 , \59670 , \59672 );
xor \U$59297 ( \59674 , \59526 , \59533 );
xor \U$59298 ( \59675 , \59674 , \59541 );
xor \U$59299 ( \59676 , \59673 , \59675 );
xor \U$59300 ( \59677 , \59475 , \59482 );
xor \U$59301 ( \59678 , \59677 , \59490 );
and \U$59302 ( \59679 , \59676 , \59678 );
and \U$59303 ( \59680 , \59673 , \59675 );
nor \U$59304 ( \59681 , \59679 , \59680 );
and \U$59305 ( \59682 , \59666 , \59681 );
and \U$59306 ( \59683 , \59663 , \59665 );
or \U$59307 ( \59684 , \59682 , \59683 );
and \U$59308 ( \59685 , \59591 , \59684 );
and \U$59309 ( \59686 , \59588 , \59590 );
or \U$59310 ( \59687 , \59685 , \59686 );
xor \U$59311 ( \59688 , \59581 , \59687 );
xor \U$59312 ( \59689 , \59331 , \59349 );
xor \U$59313 ( \59690 , \59689 , \59375 );
xor \U$59314 ( \59691 , \59468 , \59547 );
xor \U$59315 ( \59692 , \59691 , \59552 );
and \U$59316 ( \59693 , \59690 , \59692 );
and \U$59317 ( \59694 , \59688 , \59693 );
and \U$59318 ( \59695 , \59581 , \59687 );
nor \U$59319 ( \59696 , \59694 , \59695 );
or \U$59320 ( \59697 , \59577 , \59696 );
xnor \U$59321 ( \59698 , \59696 , \59577 );
and \U$59322 ( \59699 , \9760 , RIae77630_80);
and \U$59323 ( \59700 , RIae77540_78, \9758 );
nor \U$59324 ( \59701 , \59699 , \59700 );
and \U$59325 ( \59702 , \59701 , \9272 );
not \U$59326 ( \59703 , \59701 );
and \U$59327 ( \59704 , \59703 , \9273 );
nor \U$59328 ( \59705 , \59702 , \59704 );
not \U$59329 ( \59706 , \59705 );
and \U$59330 ( \59707 , \10548 , RIae776a8_81);
and \U$59331 ( \59708 , RIae77450_76, \10546 );
nor \U$59332 ( \59709 , \59707 , \59708 );
and \U$59333 ( \59710 , \59709 , \10421 );
not \U$59334 ( \59711 , \59709 );
and \U$59335 ( \59712 , \59711 , \10118 );
nor \U$59336 ( \59713 , \59710 , \59712 );
nand \U$59337 ( \59714 , \59706 , \59713 );
not \U$59338 ( \59715 , \59714 );
and \U$59339 ( \59716 , \14964 , RIae77108_69);
and \U$59340 ( \59717 , RIae77090_68, \14962 );
nor \U$59341 ( \59718 , \59716 , \59717 );
and \U$59342 ( \59719 , \59718 , \14463 );
not \U$59343 ( \59720 , \59718 );
and \U$59344 ( \59721 , \59720 , \14462 );
nor \U$59345 ( \59722 , \59719 , \59721 );
and \U$59346 ( \59723 , \15726 , RIae77270_72);
and \U$59347 ( \59724 , RIae77360_74, RIae7aab0_192);
nor \U$59348 ( \59725 , \59723 , \59724 );
and \U$59349 ( \59726 , \59725 , \14959 );
not \U$59350 ( \59727 , \59725 );
and \U$59351 ( \59728 , \59727 , RIae7aa38_191);
nor \U$59352 ( \59729 , \59726 , \59728 );
xor \U$59353 ( \59730 , \59722 , \59729 );
and \U$59354 ( \59731 , \14059 , RIae76dc0_62);
and \U$59355 ( \59732 , RIae76cd0_60, \14057 );
nor \U$59356 ( \59733 , \59731 , \59732 );
and \U$59357 ( \59734 , \59733 , \13502 );
not \U$59358 ( \59735 , \59733 );
and \U$59359 ( \59736 , \59735 , \14063 );
nor \U$59360 ( \59737 , \59734 , \59736 );
and \U$59361 ( \59738 , \59730 , \59737 );
and \U$59362 ( \59739 , \59722 , \59729 );
nor \U$59363 ( \59740 , \59738 , \59739 );
and \U$59364 ( \59741 , \11470 , RIae77ae0_90);
and \U$59365 ( \59742 , RIae779f0_88, \11468 );
nor \U$59366 ( \59743 , \59741 , \59742 );
and \U$59367 ( \59744 , \59743 , \11474 );
not \U$59368 ( \59745 , \59743 );
and \U$59369 ( \59746 , \59745 , \10936 );
nor \U$59370 ( \59747 , \59744 , \59746 );
not \U$59371 ( \59748 , \59747 );
and \U$59372 ( \59749 , \12180 , RIae77810_84);
and \U$59373 ( \59750 , RIae77900_86, \12178 );
nor \U$59374 ( \59751 , \59749 , \59750 );
and \U$59375 ( \59752 , \59751 , \11827 );
not \U$59376 ( \59753 , \59751 );
and \U$59377 ( \59754 , \59753 , \12184 );
nor \U$59378 ( \59755 , \59752 , \59754 );
not \U$59379 ( \59756 , \59755 );
and \U$59380 ( \59757 , \59748 , \59756 );
and \U$59381 ( \59758 , \59755 , \59747 );
and \U$59382 ( \59759 , \13059 , RIae76fa0_66);
and \U$59383 ( \59760 , RIae76eb0_64, \13057 );
nor \U$59384 ( \59761 , \59759 , \59760 );
and \U$59385 ( \59762 , \59761 , \12718 );
not \U$59386 ( \59763 , \59761 );
and \U$59387 ( \59764 , \59763 , \13063 );
nor \U$59388 ( \59765 , \59762 , \59764 );
nor \U$59389 ( \59766 , \59758 , \59765 );
nor \U$59390 ( \59767 , \59757 , \59766 );
xor \U$59391 ( \59768 , \59740 , \59767 );
not \U$59392 ( \59769 , \59768 );
or \U$59393 ( \59770 , \59715 , \59769 );
or \U$59394 ( \59771 , \59768 , \59714 );
nand \U$59395 ( \59772 , \59770 , \59771 );
and \U$59396 ( \59773 , \9760 , RIae77540_78);
and \U$59397 ( \59774 , RIae776a8_81, \9758 );
nor \U$59398 ( \59775 , \59773 , \59774 );
and \U$59399 ( \59776 , \59775 , \9273 );
not \U$59400 ( \59777 , \59775 );
and \U$59401 ( \59778 , \59777 , \9272 );
nor \U$59402 ( \59779 , \59776 , \59778 );
and \U$59403 ( \59780 , \10548 , RIae77450_76);
and \U$59404 ( \59781 , RIae77ae0_90, \10546 );
nor \U$59405 ( \59782 , \59780 , \59781 );
and \U$59406 ( \59783 , \59782 , \10421 );
not \U$59407 ( \59784 , \59782 );
and \U$59408 ( \59785 , \59784 , \10118 );
nor \U$59409 ( \59786 , \59783 , \59785 );
xor \U$59410 ( \59787 , \59779 , \59786 );
and \U$59411 ( \59788 , \11470 , RIae779f0_88);
and \U$59412 ( \59789 , RIae77810_84, \11468 );
nor \U$59413 ( \59790 , \59788 , \59789 );
and \U$59414 ( \59791 , \59790 , \10936 );
not \U$59415 ( \59792 , \59790 );
and \U$59416 ( \59793 , \59792 , \11474 );
nor \U$59417 ( \59794 , \59791 , \59793 );
xor \U$59418 ( \59795 , \59787 , \59794 );
nand \U$59419 ( \59796 , RIae77630_80, \8964 );
and \U$59420 ( \59797 , \59796 , \8799 );
not \U$59421 ( \59798 , \59796 );
and \U$59422 ( \59799 , \59798 , \8789 );
nor \U$59423 ( \59800 , \59797 , \59799 );
xor \U$59424 ( \59801 , \59795 , \59800 );
and \U$59425 ( \59802 , \13059 , RIae76eb0_64);
and \U$59426 ( \59803 , RIae76dc0_62, \13057 );
nor \U$59427 ( \59804 , \59802 , \59803 );
and \U$59428 ( \59805 , \59804 , \13063 );
not \U$59429 ( \59806 , \59804 );
and \U$59430 ( \59807 , \59806 , \12718 );
nor \U$59431 ( \59808 , \59805 , \59807 );
and \U$59432 ( \59809 , \12180 , RIae77900_86);
and \U$59433 ( \59810 , RIae76fa0_66, \12178 );
nor \U$59434 ( \59811 , \59809 , \59810 );
and \U$59435 ( \59812 , \59811 , \12184 );
not \U$59436 ( \59813 , \59811 );
and \U$59437 ( \59814 , \59813 , \11827 );
nor \U$59438 ( \59815 , \59812 , \59814 );
xor \U$59439 ( \59816 , \59808 , \59815 );
and \U$59440 ( \59817 , \14059 , RIae76cd0_60);
and \U$59441 ( \59818 , RIae77108_69, \14057 );
nor \U$59442 ( \59819 , \59817 , \59818 );
and \U$59443 ( \59820 , \59819 , \13502 );
not \U$59444 ( \59821 , \59819 );
and \U$59445 ( \59822 , \59821 , \14063 );
nor \U$59446 ( \59823 , \59820 , \59822 );
xor \U$59447 ( \59824 , \59816 , \59823 );
xor \U$59448 ( \59825 , \59801 , \59824 );
and \U$59449 ( \59826 , \59772 , \59825 );
xor \U$59450 ( \59827 , \59808 , \59815 );
and \U$59451 ( \59828 , \59827 , \59823 );
and \U$59452 ( \59829 , \59808 , \59815 );
or \U$59453 ( \59830 , \59828 , \59829 );
and \U$59454 ( \59831 , \15726 , RIae77360_74);
and \U$59455 ( \59832 , RIae78350_108, RIae7aab0_192);
nor \U$59456 ( \59833 , \59831 , \59832 );
and \U$59457 ( \59834 , \59833 , \14959 );
not \U$59458 ( \59835 , \59833 );
and \U$59459 ( \59836 , \59835 , RIae7aa38_191);
nor \U$59460 ( \59837 , \59834 , \59836 );
xor \U$59461 ( \59838 , \59837 , \8789 );
and \U$59462 ( \59839 , \14964 , RIae77090_68);
and \U$59463 ( \59840 , RIae77270_72, \14962 );
nor \U$59464 ( \59841 , \59839 , \59840 );
and \U$59465 ( \59842 , \59841 , \14463 );
not \U$59466 ( \59843 , \59841 );
and \U$59467 ( \59844 , \59843 , \14462 );
nor \U$59468 ( \59845 , \59842 , \59844 );
and \U$59469 ( \59846 , \59838 , \59845 );
and \U$59470 ( \59847 , \59837 , \8789 );
or \U$59471 ( \59848 , \59846 , \59847 );
xor \U$59472 ( \59849 , \59830 , \59848 );
xor \U$59473 ( \59850 , \59779 , \59786 );
and \U$59474 ( \59851 , \59850 , \59794 );
and \U$59475 ( \59852 , \59779 , \59786 );
or \U$59476 ( \59853 , \59851 , \59852 );
xor \U$59477 ( \59854 , \59849 , \59853 );
xor \U$59478 ( \59855 , \59826 , \59854 );
and \U$59479 ( \59856 , \12180 , RIae779f0_88);
and \U$59480 ( \59857 , RIae77810_84, \12178 );
nor \U$59481 ( \59858 , \59856 , \59857 );
and \U$59482 ( \59859 , \59858 , \11827 );
not \U$59483 ( \59860 , \59858 );
and \U$59484 ( \59861 , \59860 , \12184 );
nor \U$59485 ( \59862 , \59859 , \59861 );
and \U$59486 ( \59863 , \13059 , RIae77900_86);
and \U$59487 ( \59864 , RIae76fa0_66, \13057 );
nor \U$59488 ( \59865 , \59863 , \59864 );
and \U$59489 ( \59866 , \59865 , \12718 );
not \U$59490 ( \59867 , \59865 );
and \U$59491 ( \59868 , \59867 , \13063 );
nor \U$59492 ( \59869 , \59866 , \59868 );
xor \U$59493 ( \59870 , \59862 , \59869 );
and \U$59494 ( \59871 , \14059 , RIae76eb0_64);
and \U$59495 ( \59872 , RIae76dc0_62, \14057 );
nor \U$59496 ( \59873 , \59871 , \59872 );
and \U$59497 ( \59874 , \59873 , \14063 );
not \U$59498 ( \59875 , \59873 );
and \U$59499 ( \59876 , \59875 , \13502 );
nor \U$59500 ( \59877 , \59874 , \59876 );
and \U$59501 ( \59878 , \59870 , \59877 );
and \U$59502 ( \59879 , \59862 , \59869 );
or \U$59503 ( \59880 , \59878 , \59879 );
and \U$59504 ( \59881 , \15726 , RIae77090_68);
and \U$59505 ( \59882 , RIae77270_72, RIae7aab0_192);
nor \U$59506 ( \59883 , \59881 , \59882 );
and \U$59507 ( \59884 , \59883 , \14959 );
not \U$59508 ( \59885 , \59883 );
and \U$59509 ( \59886 , \59885 , RIae7aa38_191);
nor \U$59510 ( \59887 , \59884 , \59886 );
and \U$59511 ( \59888 , \59887 , \9764 );
not \U$59512 ( \59889 , \59887 );
not \U$59513 ( \59890 , \9272 );
and \U$59514 ( \59891 , \59889 , \59890 );
and \U$59515 ( \59892 , \14964 , RIae76cd0_60);
and \U$59516 ( \59893 , RIae77108_69, \14962 );
nor \U$59517 ( \59894 , \59892 , \59893 );
and \U$59518 ( \59895 , \59894 , \14462 );
not \U$59519 ( \59896 , \59894 );
and \U$59520 ( \59897 , \59896 , \14463 );
nor \U$59521 ( \59898 , \59895 , \59897 );
nor \U$59522 ( \59899 , \59891 , \59898 );
nor \U$59523 ( \59900 , \59888 , \59899 );
or \U$59524 ( \59901 , \59880 , \59900 );
not \U$59525 ( \59902 , \59900 );
not \U$59526 ( \59903 , \59880 );
or \U$59527 ( \59904 , \59902 , \59903 );
and \U$59528 ( \59905 , \10548 , RIae77540_78);
and \U$59529 ( \59906 , RIae776a8_81, \10546 );
nor \U$59530 ( \59907 , \59905 , \59906 );
and \U$59531 ( \59908 , \59907 , \10421 );
not \U$59532 ( \59909 , \59907 );
and \U$59533 ( \59910 , \59909 , \10118 );
nor \U$59534 ( \59911 , \59908 , \59910 );
nand \U$59535 ( \59912 , RIae77630_80, \9758 );
and \U$59536 ( \59913 , \59912 , \9273 );
not \U$59537 ( \59914 , \59912 );
and \U$59538 ( \59915 , \59914 , \9764 );
nor \U$59539 ( \59916 , \59913 , \59915 );
xor \U$59540 ( \59917 , \59911 , \59916 );
and \U$59541 ( \59918 , \11470 , RIae77450_76);
and \U$59542 ( \59919 , RIae77ae0_90, \11468 );
nor \U$59543 ( \59920 , \59918 , \59919 );
and \U$59544 ( \59921 , \59920 , \10936 );
not \U$59545 ( \59922 , \59920 );
and \U$59546 ( \59923 , \59922 , \11474 );
nor \U$59547 ( \59924 , \59921 , \59923 );
and \U$59548 ( \59925 , \59917 , \59924 );
and \U$59549 ( \59926 , \59911 , \59916 );
or \U$59550 ( \59927 , \59925 , \59926 );
nand \U$59551 ( \59928 , \59904 , \59927 );
nand \U$59552 ( \59929 , \59901 , \59928 );
xor \U$59553 ( \59930 , \59837 , \8789 );
xor \U$59554 ( \59931 , \59930 , \59845 );
xor \U$59555 ( \59932 , \59929 , \59931 );
not \U$59556 ( \59933 , \59705 );
not \U$59557 ( \59934 , \59713 );
or \U$59558 ( \59935 , \59933 , \59934 );
or \U$59559 ( \59936 , \59705 , \59713 );
nand \U$59560 ( \59937 , \59935 , \59936 );
not \U$59561 ( \59938 , \59937 );
not \U$59562 ( \59939 , \59747 );
xor \U$59563 ( \59940 , \59755 , \59765 );
not \U$59564 ( \59941 , \59940 );
or \U$59565 ( \59942 , \59939 , \59941 );
or \U$59566 ( \59943 , \59940 , \59747 );
nand \U$59567 ( \59944 , \59942 , \59943 );
not \U$59568 ( \59945 , \59944 );
or \U$59569 ( \59946 , \59938 , \59945 );
or \U$59570 ( \59947 , \59944 , \59937 );
xor \U$59571 ( \59948 , \59722 , \59729 );
xor \U$59572 ( \59949 , \59948 , \59737 );
nand \U$59573 ( \59950 , \59947 , \59949 );
nand \U$59574 ( \59951 , \59946 , \59950 );
and \U$59575 ( \59952 , \59932 , \59951 );
and \U$59576 ( \59953 , \59929 , \59931 );
or \U$59577 ( \59954 , \59952 , \59953 );
xor \U$59578 ( \59955 , \59855 , \59954 );
not \U$59579 ( \59956 , \59955 );
not \U$59580 ( \59957 , \59740 );
not \U$59581 ( \59958 , \59714 );
and \U$59582 ( \59959 , \59957 , \59958 );
and \U$59583 ( \59960 , \59740 , \59714 );
nor \U$59584 ( \59961 , \59960 , \59767 );
nor \U$59585 ( \59962 , \59959 , \59961 );
xor \U$59586 ( \59963 , \59795 , \59800 );
and \U$59587 ( \59964 , \59963 , \59824 );
and \U$59588 ( \59965 , \59795 , \59800 );
nor \U$59589 ( \59966 , \59964 , \59965 );
xor \U$59590 ( \59967 , \59962 , \59966 );
and \U$59591 ( \59968 , \11470 , RIae77810_84);
and \U$59592 ( \59969 , RIae77900_86, \11468 );
nor \U$59593 ( \59970 , \59968 , \59969 );
and \U$59594 ( \59971 , \59970 , \11474 );
not \U$59595 ( \59972 , \59970 );
and \U$59596 ( \59973 , \59972 , \10936 );
nor \U$59597 ( \59974 , \59971 , \59973 );
not \U$59598 ( \59975 , \59974 );
and \U$59599 ( \59976 , \12180 , RIae76fa0_66);
and \U$59600 ( \59977 , RIae76eb0_64, \12178 );
nor \U$59601 ( \59978 , \59976 , \59977 );
and \U$59602 ( \59979 , \59978 , \11827 );
not \U$59603 ( \59980 , \59978 );
and \U$59604 ( \59981 , \59980 , \12184 );
nor \U$59605 ( \59982 , \59979 , \59981 );
and \U$59606 ( \59983 , \13059 , RIae76dc0_62);
and \U$59607 ( \59984 , RIae76cd0_60, \13057 );
nor \U$59608 ( \59985 , \59983 , \59984 );
and \U$59609 ( \59986 , \59985 , \12718 );
not \U$59610 ( \59987 , \59985 );
and \U$59611 ( \59988 , \59987 , \13063 );
nor \U$59612 ( \59989 , \59986 , \59988 );
xor \U$59613 ( \59990 , \59982 , \59989 );
not \U$59614 ( \59991 , \59990 );
or \U$59615 ( \59992 , \59975 , \59991 );
or \U$59616 ( \59993 , \59990 , \59974 );
nand \U$59617 ( \59994 , \59992 , \59993 );
not \U$59618 ( \59995 , \59994 );
and \U$59619 ( \59996 , \14964 , RIae77270_72);
and \U$59620 ( \59997 , RIae77360_74, \14962 );
nor \U$59621 ( \59998 , \59996 , \59997 );
and \U$59622 ( \59999 , \59998 , \14462 );
not \U$59623 ( \60000 , \59998 );
and \U$59624 ( \60001 , \60000 , \14463 );
nor \U$59625 ( \60002 , \59999 , \60001 );
and \U$59626 ( \60003 , \15726 , RIae78350_108);
and \U$59627 ( \60004 , RIae78170_104, RIae7aab0_192);
nor \U$59628 ( \60005 , \60003 , \60004 );
and \U$59629 ( \60006 , \60005 , RIae7aa38_191);
not \U$59630 ( \60007 , \60005 );
and \U$59631 ( \60008 , \60007 , \14959 );
nor \U$59632 ( \60009 , \60006 , \60008 );
xor \U$59633 ( \60010 , \60002 , \60009 );
and \U$59634 ( \60011 , \14059 , RIae77108_69);
and \U$59635 ( \60012 , RIae77090_68, \14057 );
nor \U$59636 ( \60013 , \60011 , \60012 );
and \U$59637 ( \60014 , \60013 , \14063 );
not \U$59638 ( \60015 , \60013 );
and \U$59639 ( \60016 , \60015 , \13502 );
nor \U$59640 ( \60017 , \60014 , \60016 );
xor \U$59641 ( \60018 , \60010 , \60017 );
not \U$59642 ( \60019 , \60018 );
or \U$59643 ( \60020 , \59995 , \60019 );
or \U$59644 ( \60021 , \60018 , \59994 );
nand \U$59645 ( \60022 , \60020 , \60021 );
not \U$59646 ( \60023 , \60022 );
and \U$59647 ( \60024 , \8966 , RIae77630_80);
and \U$59648 ( \60025 , RIae77540_78, \8964 );
nor \U$59649 ( \60026 , \60024 , \60025 );
and \U$59650 ( \60027 , \60026 , \8789 );
not \U$59651 ( \60028 , \60026 );
and \U$59652 ( \60029 , \60028 , \8799 );
nor \U$59653 ( \60030 , \60027 , \60029 );
and \U$59654 ( \60031 , \9760 , RIae776a8_81);
and \U$59655 ( \60032 , RIae77450_76, \9758 );
nor \U$59656 ( \60033 , \60031 , \60032 );
and \U$59657 ( \60034 , \60033 , \9272 );
not \U$59658 ( \60035 , \60033 );
and \U$59659 ( \60036 , \60035 , \9273 );
nor \U$59660 ( \60037 , \60034 , \60036 );
xor \U$59661 ( \60038 , \60030 , \60037 );
and \U$59662 ( \60039 , \10548 , RIae77ae0_90);
and \U$59663 ( \60040 , RIae779f0_88, \10546 );
nor \U$59664 ( \60041 , \60039 , \60040 );
and \U$59665 ( \60042 , \60041 , \10118 );
not \U$59666 ( \60043 , \60041 );
and \U$59667 ( \60044 , \60043 , \10421 );
nor \U$59668 ( \60045 , \60042 , \60044 );
xor \U$59669 ( \60046 , \60038 , \60045 );
not \U$59670 ( \60047 , \60046 );
and \U$59671 ( \60048 , \60023 , \60047 );
and \U$59672 ( \60049 , \60022 , \60046 );
nor \U$59673 ( \60050 , \60048 , \60049 );
xor \U$59674 ( \60051 , \59967 , \60050 );
not \U$59675 ( \60052 , \60051 );
and \U$59676 ( \60053 , \59956 , \60052 );
and \U$59677 ( \60054 , \59955 , \60051 );
nor \U$59678 ( \60055 , \60053 , \60054 );
xor \U$59679 ( \60056 , \59929 , \59931 );
xor \U$59680 ( \60057 , \60056 , \59951 );
xor \U$59681 ( \60058 , \59772 , \59825 );
and \U$59682 ( \60059 , \60057 , \60058 );
not \U$59683 ( \60060 , \60057 );
not \U$59684 ( \60061 , \60058 );
and \U$59685 ( \60062 , \60060 , \60061 );
and \U$59686 ( \60063 , \11470 , RIae776a8_81);
and \U$59687 ( \60064 , RIae77450_76, \11468 );
nor \U$59688 ( \60065 , \60063 , \60064 );
and \U$59689 ( \60066 , \60065 , \10936 );
not \U$59690 ( \60067 , \60065 );
and \U$59691 ( \60068 , \60067 , \11474 );
nor \U$59692 ( \60069 , \60066 , \60068 );
and \U$59693 ( \60070 , \12180 , RIae77ae0_90);
and \U$59694 ( \60071 , RIae779f0_88, \12178 );
nor \U$59695 ( \60072 , \60070 , \60071 );
and \U$59696 ( \60073 , \60072 , \12184 );
not \U$59697 ( \60074 , \60072 );
and \U$59698 ( \60075 , \60074 , \11827 );
nor \U$59699 ( \60076 , \60073 , \60075 );
xor \U$59700 ( \60077 , \60069 , \60076 );
and \U$59701 ( \60078 , \13059 , RIae77810_84);
and \U$59702 ( \60079 , RIae77900_86, \13057 );
nor \U$59703 ( \60080 , \60078 , \60079 );
and \U$59704 ( \60081 , \60080 , \13063 );
not \U$59705 ( \60082 , \60080 );
and \U$59706 ( \60083 , \60082 , \12718 );
nor \U$59707 ( \60084 , \60081 , \60083 );
and \U$59708 ( \60085 , \60077 , \60084 );
and \U$59709 ( \60086 , \60069 , \60076 );
or \U$59710 ( \60087 , \60085 , \60086 );
and \U$59711 ( \60088 , \14964 , RIae76dc0_62);
and \U$59712 ( \60089 , RIae76cd0_60, \14962 );
nor \U$59713 ( \60090 , \60088 , \60089 );
and \U$59714 ( \60091 , \60090 , \14463 );
not \U$59715 ( \60092 , \60090 );
and \U$59716 ( \60093 , \60092 , \14462 );
nor \U$59717 ( \60094 , \60091 , \60093 );
and \U$59718 ( \60095 , \15726 , RIae77108_69);
and \U$59719 ( \60096 , RIae77090_68, RIae7aab0_192);
nor \U$59720 ( \60097 , \60095 , \60096 );
and \U$59721 ( \60098 , \60097 , \14959 );
not \U$59722 ( \60099 , \60097 );
and \U$59723 ( \60100 , \60099 , RIae7aa38_191);
nor \U$59724 ( \60101 , \60098 , \60100 );
xor \U$59725 ( \60102 , \60094 , \60101 );
and \U$59726 ( \60103 , \14059 , RIae76fa0_66);
and \U$59727 ( \60104 , RIae76eb0_64, \14057 );
nor \U$59728 ( \60105 , \60103 , \60104 );
and \U$59729 ( \60106 , \60105 , \13502 );
not \U$59730 ( \60107 , \60105 );
and \U$59731 ( \60108 , \60107 , \14063 );
nor \U$59732 ( \60109 , \60106 , \60108 );
and \U$59733 ( \60110 , \60102 , \60109 );
and \U$59734 ( \60111 , \60094 , \60101 );
or \U$59735 ( \60112 , \60110 , \60111 );
xor \U$59736 ( \60113 , \60087 , \60112 );
xor \U$59737 ( \60114 , \59911 , \59916 );
xor \U$59738 ( \60115 , \60114 , \59924 );
and \U$59739 ( \60116 , \60113 , \60115 );
and \U$59740 ( \60117 , \60087 , \60112 );
nor \U$59741 ( \60118 , \60116 , \60117 );
xor \U$59742 ( \60119 , \59862 , \59869 );
xor \U$59743 ( \60120 , \60119 , \59877 );
not \U$59744 ( \60121 , \60120 );
not \U$59745 ( \60122 , \9273 );
not \U$59746 ( \60123 , \59887 );
not \U$59747 ( \60124 , \59898 );
or \U$59748 ( \60125 , \60123 , \60124 );
or \U$59749 ( \60126 , \59898 , \59887 );
nand \U$59750 ( \60127 , \60125 , \60126 );
not \U$59751 ( \60128 , \60127 );
or \U$59752 ( \60129 , \60122 , \60128 );
or \U$59753 ( \60130 , \60127 , \9273 );
nand \U$59754 ( \60131 , \60129 , \60130 );
nand \U$59755 ( \60132 , \60121 , \60131 );
xor \U$59756 ( \60133 , \60118 , \60132 );
xnor \U$59757 ( \60134 , \59949 , \59944 );
not \U$59758 ( \60135 , \60134 );
not \U$59759 ( \60136 , \59937 );
and \U$59760 ( \60137 , \60135 , \60136 );
and \U$59761 ( \60138 , \60134 , \59937 );
nor \U$59762 ( \60139 , \60137 , \60138 );
and \U$59763 ( \60140 , \60133 , \60139 );
and \U$59764 ( \60141 , \60118 , \60132 );
or \U$59765 ( \60142 , \60140 , \60141 );
nor \U$59766 ( \60143 , \60062 , \60142 );
nor \U$59767 ( \60144 , \60059 , \60143 );
or \U$59768 ( \60145 , \60055 , \60144 );
xnor \U$59769 ( \60146 , \60144 , \60055 );
not \U$59770 ( \60147 , \60058 );
not \U$59771 ( \60148 , \60142 );
not \U$59772 ( \60149 , \60057 );
and \U$59773 ( \60150 , \60148 , \60149 );
and \U$59774 ( \60151 , \60142 , \60057 );
nor \U$59775 ( \60152 , \60150 , \60151 );
not \U$59776 ( \60153 , \60152 );
or \U$59777 ( \60154 , \60147 , \60153 );
or \U$59778 ( \60155 , \60152 , \60058 );
nand \U$59779 ( \60156 , \60154 , \60155 );
xor \U$59780 ( \60157 , \60118 , \60132 );
xor \U$59781 ( \60158 , \60157 , \60139 );
not \U$59782 ( \60159 , \59900 );
not \U$59783 ( \60160 , \59927 );
or \U$59784 ( \60161 , \60159 , \60160 );
or \U$59785 ( \60162 , \59927 , \59900 );
nand \U$59786 ( \60163 , \60161 , \60162 );
not \U$59787 ( \60164 , \60163 );
not \U$59788 ( \60165 , \59880 );
and \U$59789 ( \60166 , \60164 , \60165 );
and \U$59790 ( \60167 , \60163 , \59880 );
nor \U$59791 ( \60168 , \60166 , \60167 );
or \U$59792 ( \60169 , \60158 , \60168 );
not \U$59793 ( \60170 , \60168 );
not \U$59794 ( \60171 , \60158 );
or \U$59795 ( \60172 , \60170 , \60171 );
not \U$59796 ( \60173 , \60120 );
not \U$59797 ( \60174 , \60131 );
or \U$59798 ( \60175 , \60173 , \60174 );
or \U$59799 ( \60176 , \60131 , \60120 );
nand \U$59800 ( \60177 , \60175 , \60176 );
and \U$59801 ( \60178 , \15726 , RIae76cd0_60);
and \U$59802 ( \60179 , RIae77108_69, RIae7aab0_192);
nor \U$59803 ( \60180 , \60178 , \60179 );
and \U$59804 ( \60181 , \60180 , \14959 );
not \U$59805 ( \60182 , \60180 );
and \U$59806 ( \60183 , \60182 , RIae7aa38_191);
nor \U$59807 ( \60184 , \60181 , \60183 );
xor \U$59808 ( \60185 , \60184 , \10118 );
and \U$59809 ( \60186 , \14964 , RIae76eb0_64);
and \U$59810 ( \60187 , RIae76dc0_62, \14962 );
nor \U$59811 ( \60188 , \60186 , \60187 );
and \U$59812 ( \60189 , \60188 , \14463 );
not \U$59813 ( \60190 , \60188 );
and \U$59814 ( \60191 , \60190 , \14462 );
nor \U$59815 ( \60192 , \60189 , \60191 );
and \U$59816 ( \60193 , \60185 , \60192 );
and \U$59817 ( \60194 , \60184 , \10118 );
or \U$59818 ( \60195 , \60193 , \60194 );
and \U$59819 ( \60196 , \10548 , RIae77630_80);
and \U$59820 ( \60197 , RIae77540_78, \10546 );
nor \U$59821 ( \60198 , \60196 , \60197 );
and \U$59822 ( \60199 , \60198 , \10421 );
not \U$59823 ( \60200 , \60198 );
and \U$59824 ( \60201 , \60200 , \10118 );
nor \U$59825 ( \60202 , \60199 , \60201 );
xor \U$59826 ( \60203 , \60195 , \60202 );
and \U$59827 ( \60204 , \13059 , RIae779f0_88);
and \U$59828 ( \60205 , RIae77810_84, \13057 );
nor \U$59829 ( \60206 , \60204 , \60205 );
and \U$59830 ( \60207 , \60206 , \13063 );
not \U$59831 ( \60208 , \60206 );
and \U$59832 ( \60209 , \60208 , \12718 );
nor \U$59833 ( \60210 , \60207 , \60209 );
and \U$59834 ( \60211 , \12180 , RIae77450_76);
and \U$59835 ( \60212 , RIae77ae0_90, \12178 );
nor \U$59836 ( \60213 , \60211 , \60212 );
and \U$59837 ( \60214 , \60213 , \12184 );
not \U$59838 ( \60215 , \60213 );
and \U$59839 ( \60216 , \60215 , \11827 );
nor \U$59840 ( \60217 , \60214 , \60216 );
xor \U$59841 ( \60218 , \60210 , \60217 );
and \U$59842 ( \60219 , \14059 , RIae77900_86);
and \U$59843 ( \60220 , RIae76fa0_66, \14057 );
nor \U$59844 ( \60221 , \60219 , \60220 );
and \U$59845 ( \60222 , \60221 , \13502 );
not \U$59846 ( \60223 , \60221 );
and \U$59847 ( \60224 , \60223 , \14063 );
nor \U$59848 ( \60225 , \60222 , \60224 );
and \U$59849 ( \60226 , \60218 , \60225 );
and \U$59850 ( \60227 , \60210 , \60217 );
or \U$59851 ( \60228 , \60226 , \60227 );
and \U$59852 ( \60229 , \60203 , \60228 );
and \U$59853 ( \60230 , \60195 , \60202 );
or \U$59854 ( \60231 , \60229 , \60230 );
xor \U$59855 ( \60232 , \60177 , \60231 );
xor \U$59856 ( \60233 , \60087 , \60112 );
xor \U$59857 ( \60234 , \60233 , \60115 );
and \U$59858 ( \60235 , \60232 , \60234 );
and \U$59859 ( \60236 , \60177 , \60231 );
or \U$59860 ( \60237 , \60235 , \60236 );
nand \U$59861 ( \60238 , \60172 , \60237 );
nand \U$59862 ( \60239 , \60169 , \60238 );
and \U$59863 ( \60240 , \60156 , \60239 );
xor \U$59864 ( \60241 , \60239 , \60156 );
xor \U$59865 ( \60242 , \60094 , \60101 );
xor \U$59866 ( \60243 , \60242 , \60109 );
xor \U$59867 ( \60244 , \60195 , \60202 );
xor \U$59868 ( \60245 , \60244 , \60228 );
xor \U$59869 ( \60246 , \60243 , \60245 );
not \U$59870 ( \60247 , \60246 );
and \U$59871 ( \60248 , \15726 , RIae76dc0_62);
and \U$59872 ( \60249 , RIae76cd0_60, RIae7aab0_192);
nor \U$59873 ( \60250 , \60248 , \60249 );
and \U$59874 ( \60251 , \60250 , RIae7aa38_191);
not \U$59875 ( \60252 , \60250 );
and \U$59876 ( \60253 , \60252 , \14959 );
nor \U$59877 ( \60254 , \60251 , \60253 );
and \U$59878 ( \60255 , \14964 , RIae76fa0_66);
and \U$59879 ( \60256 , RIae76eb0_64, \14962 );
nor \U$59880 ( \60257 , \60255 , \60256 );
and \U$59881 ( \60258 , \60257 , \14462 );
not \U$59882 ( \60259 , \60257 );
and \U$59883 ( \60260 , \60259 , \14463 );
nor \U$59884 ( \60261 , \60258 , \60260 );
xor \U$59885 ( \60262 , \60254 , \60261 );
and \U$59886 ( \60263 , \14059 , RIae77810_84);
and \U$59887 ( \60264 , RIae77900_86, \14057 );
nor \U$59888 ( \60265 , \60263 , \60264 );
and \U$59889 ( \60266 , \60265 , \14063 );
not \U$59890 ( \60267 , \60265 );
and \U$59891 ( \60268 , \60267 , \13502 );
nor \U$59892 ( \60269 , \60266 , \60268 );
and \U$59893 ( \60270 , \60262 , \60269 );
and \U$59894 ( \60271 , \60254 , \60261 );
nor \U$59895 ( \60272 , \60270 , \60271 );
and \U$59896 ( \60273 , \11470 , RIae77540_78);
and \U$59897 ( \60274 , RIae776a8_81, \11468 );
nor \U$59898 ( \60275 , \60273 , \60274 );
and \U$59899 ( \60276 , \60275 , \10936 );
not \U$59900 ( \60277 , \60275 );
and \U$59901 ( \60278 , \60277 , \11474 );
nor \U$59902 ( \60279 , \60276 , \60278 );
xor \U$59903 ( \60280 , \60272 , \60279 );
and \U$59904 ( \60281 , \11470 , RIae77630_80);
and \U$59905 ( \60282 , RIae77540_78, \11468 );
nor \U$59906 ( \60283 , \60281 , \60282 );
and \U$59907 ( \60284 , \60283 , \11474 );
not \U$59908 ( \60285 , \60283 );
and \U$59909 ( \60286 , \60285 , \10936 );
nor \U$59910 ( \60287 , \60284 , \60286 );
and \U$59911 ( \60288 , \12180 , RIae776a8_81);
and \U$59912 ( \60289 , RIae77450_76, \12178 );
nor \U$59913 ( \60290 , \60288 , \60289 );
and \U$59914 ( \60291 , \60290 , \11827 );
not \U$59915 ( \60292 , \60290 );
and \U$59916 ( \60293 , \60292 , \12184 );
nor \U$59917 ( \60294 , \60291 , \60293 );
or \U$59918 ( \60295 , \60287 , \60294 );
not \U$59919 ( \60296 , \60294 );
not \U$59920 ( \60297 , \60287 );
or \U$59921 ( \60298 , \60296 , \60297 );
and \U$59922 ( \60299 , \13059 , RIae77ae0_90);
and \U$59923 ( \60300 , RIae779f0_88, \13057 );
nor \U$59924 ( \60301 , \60299 , \60300 );
and \U$59925 ( \60302 , \60301 , \13063 );
not \U$59926 ( \60303 , \60301 );
and \U$59927 ( \60304 , \60303 , \12718 );
nor \U$59928 ( \60305 , \60302 , \60304 );
nand \U$59929 ( \60306 , \60298 , \60305 );
nand \U$59930 ( \60307 , \60295 , \60306 );
and \U$59931 ( \60308 , \60280 , \60307 );
and \U$59932 ( \60309 , \60272 , \60279 );
or \U$59933 ( \60310 , \60308 , \60309 );
xor \U$59934 ( \60311 , \60069 , \60076 );
xor \U$59935 ( \60312 , \60311 , \60084 );
xor \U$59936 ( \60313 , \60310 , \60312 );
nand \U$59937 ( \60314 , RIae77630_80, \10546 );
and \U$59938 ( \60315 , \60314 , \10421 );
not \U$59939 ( \60316 , \60314 );
and \U$59940 ( \60317 , \60316 , \10118 );
nor \U$59941 ( \60318 , \60315 , \60317 );
xor \U$59942 ( \60319 , \60210 , \60217 );
xor \U$59943 ( \60320 , \60319 , \60225 );
and \U$59944 ( \60321 , \60318 , \60320 );
xor \U$59945 ( \60322 , \60184 , \10118 );
xor \U$59946 ( \60323 , \60322 , \60192 );
xor \U$59947 ( \60324 , \60210 , \60217 );
xor \U$59948 ( \60325 , \60324 , \60225 );
and \U$59949 ( \60326 , \60323 , \60325 );
and \U$59950 ( \60327 , \60318 , \60323 );
or \U$59951 ( \60328 , \60321 , \60326 , \60327 );
xor \U$59952 ( \60329 , \60313 , \60328 );
not \U$59953 ( \60330 , \60329 );
or \U$59954 ( \60331 , \60247 , \60330 );
or \U$59955 ( \60332 , \60329 , \60246 );
not \U$59956 ( \60333 , \60294 );
not \U$59957 ( \60334 , \60305 );
or \U$59958 ( \60335 , \60333 , \60334 );
or \U$59959 ( \60336 , \60294 , \60305 );
nand \U$59960 ( \60337 , \60335 , \60336 );
not \U$59961 ( \60338 , \60337 );
not \U$59962 ( \60339 , \60287 );
and \U$59963 ( \60340 , \60338 , \60339 );
and \U$59964 ( \60341 , \60337 , \60287 );
nor \U$59965 ( \60342 , \60340 , \60341 );
and \U$59966 ( \60343 , \15726 , RIae76eb0_64);
and \U$59967 ( \60344 , RIae76dc0_62, RIae7aab0_192);
nor \U$59968 ( \60345 , \60343 , \60344 );
and \U$59969 ( \60346 , \60345 , \14959 );
not \U$59970 ( \60347 , \60345 );
and \U$59971 ( \60348 , \60347 , RIae7aa38_191);
nor \U$59972 ( \60349 , \60346 , \60348 );
and \U$59973 ( \60350 , \60349 , \11474 );
not \U$59974 ( \60351 , \60349 );
not \U$59975 ( \60352 , \11474 );
and \U$59976 ( \60353 , \60351 , \60352 );
and \U$59977 ( \60354 , \14964 , RIae77900_86);
and \U$59978 ( \60355 , RIae76fa0_66, \14962 );
nor \U$59979 ( \60356 , \60354 , \60355 );
and \U$59980 ( \60357 , \60356 , \14462 );
not \U$59981 ( \60358 , \60356 );
and \U$59982 ( \60359 , \60358 , \14463 );
nor \U$59983 ( \60360 , \60357 , \60359 );
nor \U$59984 ( \60361 , \60353 , \60360 );
nor \U$59985 ( \60362 , \60350 , \60361 );
or \U$59986 ( \60363 , \60342 , \60362 );
not \U$59987 ( \60364 , \60362 );
not \U$59988 ( \60365 , \60342 );
or \U$59989 ( \60366 , \60364 , \60365 );
and \U$59990 ( \60367 , \12180 , RIae77540_78);
and \U$59991 ( \60368 , RIae776a8_81, \12178 );
nor \U$59992 ( \60369 , \60367 , \60368 );
and \U$59993 ( \60370 , \60369 , \11827 );
not \U$59994 ( \60371 , \60369 );
and \U$59995 ( \60372 , \60371 , \12184 );
nor \U$59996 ( \60373 , \60370 , \60372 );
and \U$59997 ( \60374 , \13059 , RIae77450_76);
and \U$59998 ( \60375 , RIae77ae0_90, \13057 );
nor \U$59999 ( \60376 , \60374 , \60375 );
and \U$60000 ( \60377 , \60376 , \12718 );
not \U$60001 ( \60378 , \60376 );
and \U$60002 ( \60379 , \60378 , \13063 );
nor \U$60003 ( \60380 , \60377 , \60379 );
or \U$60004 ( \60381 , \60373 , \60380 );
not \U$60005 ( \60382 , \60380 );
not \U$60006 ( \60383 , \60373 );
or \U$60007 ( \60384 , \60382 , \60383 );
and \U$60008 ( \60385 , \14059 , RIae779f0_88);
and \U$60009 ( \60386 , RIae77810_84, \14057 );
nor \U$60010 ( \60387 , \60385 , \60386 );
and \U$60011 ( \60388 , \60387 , \13502 );
not \U$60012 ( \60389 , \60387 );
and \U$60013 ( \60390 , \60389 , \14063 );
nor \U$60014 ( \60391 , \60388 , \60390 );
nand \U$60015 ( \60392 , \60384 , \60391 );
nand \U$60016 ( \60393 , \60381 , \60392 );
nand \U$60017 ( \60394 , \60366 , \60393 );
nand \U$60018 ( \60395 , \60363 , \60394 );
xor \U$60019 ( \60396 , \60272 , \60279 );
xor \U$60020 ( \60397 , \60396 , \60307 );
and \U$60021 ( \60398 , \60395 , \60397 );
xor \U$60022 ( \60399 , \60210 , \60217 );
xor \U$60023 ( \60400 , \60399 , \60225 );
xor \U$60024 ( \60401 , \60318 , \60323 );
xor \U$60025 ( \60402 , \60400 , \60401 );
xor \U$60026 ( \60403 , \60272 , \60279 );
xor \U$60027 ( \60404 , \60403 , \60307 );
and \U$60028 ( \60405 , \60402 , \60404 );
and \U$60029 ( \60406 , \60395 , \60402 );
or \U$60030 ( \60407 , \60398 , \60405 , \60406 );
nand \U$60031 ( \60408 , \60332 , \60407 );
nand \U$60032 ( \60409 , \60331 , \60408 );
xor \U$60033 ( \60410 , \60177 , \60231 );
xor \U$60034 ( \60411 , \60410 , \60234 );
and \U$60035 ( \60412 , \60243 , \60245 );
xor \U$60036 ( \60413 , \60411 , \60412 );
xor \U$60037 ( \60414 , \60310 , \60312 );
and \U$60038 ( \60415 , \60414 , \60328 );
and \U$60039 ( \60416 , \60310 , \60312 );
or \U$60040 ( \60417 , \60415 , \60416 );
xor \U$60041 ( \60418 , \60413 , \60417 );
and \U$60042 ( \60419 , \60409 , \60418 );
xor \U$60043 ( \60420 , \60418 , \60409 );
and \U$60044 ( \60421 , \14964 , RIae77810_84);
and \U$60045 ( \60422 , RIae77900_86, \14962 );
nor \U$60046 ( \60423 , \60421 , \60422 );
and \U$60047 ( \60424 , \60423 , \14463 );
not \U$60048 ( \60425 , \60423 );
and \U$60049 ( \60426 , \60425 , \14462 );
nor \U$60050 ( \60427 , \60424 , \60426 );
and \U$60051 ( \60428 , \15726 , RIae76fa0_66);
and \U$60052 ( \60429 , RIae76eb0_64, RIae7aab0_192);
nor \U$60053 ( \60430 , \60428 , \60429 );
and \U$60054 ( \60431 , \60430 , \14959 );
not \U$60055 ( \60432 , \60430 );
and \U$60056 ( \60433 , \60432 , RIae7aa38_191);
nor \U$60057 ( \60434 , \60431 , \60433 );
xor \U$60058 ( \60435 , \60427 , \60434 );
and \U$60059 ( \60436 , \14059 , RIae77ae0_90);
and \U$60060 ( \60437 , RIae779f0_88, \14057 );
nor \U$60061 ( \60438 , \60436 , \60437 );
and \U$60062 ( \60439 , \60438 , \13502 );
not \U$60063 ( \60440 , \60438 );
and \U$60064 ( \60441 , \60440 , \14063 );
nor \U$60065 ( \60442 , \60439 , \60441 );
and \U$60066 ( \60443 , \60435 , \60442 );
and \U$60067 ( \60444 , \60427 , \60434 );
nor \U$60068 ( \60445 , \60443 , \60444 );
nand \U$60069 ( \60446 , RIae77630_80, \11468 );
and \U$60070 ( \60447 , \60446 , \11474 );
not \U$60071 ( \60448 , \60446 );
and \U$60072 ( \60449 , \60448 , \10936 );
nor \U$60073 ( \60450 , \60447 , \60449 );
xor \U$60074 ( \60451 , \60445 , \60450 );
not \U$60075 ( \60452 , \60380 );
not \U$60076 ( \60453 , \60391 );
or \U$60077 ( \60454 , \60452 , \60453 );
or \U$60078 ( \60455 , \60380 , \60391 );
nand \U$60079 ( \60456 , \60454 , \60455 );
not \U$60080 ( \60457 , \60456 );
not \U$60081 ( \60458 , \60373 );
and \U$60082 ( \60459 , \60457 , \60458 );
and \U$60083 ( \60460 , \60456 , \60373 );
nor \U$60084 ( \60461 , \60459 , \60460 );
and \U$60085 ( \60462 , \60451 , \60461 );
and \U$60086 ( \60463 , \60445 , \60450 );
or \U$60087 ( \60464 , \60462 , \60463 );
xor \U$60088 ( \60465 , \60254 , \60261 );
xor \U$60089 ( \60466 , \60465 , \60269 );
xor \U$60090 ( \60467 , \60464 , \60466 );
not \U$60091 ( \60468 , \60362 );
not \U$60092 ( \60469 , \60393 );
or \U$60093 ( \60470 , \60468 , \60469 );
or \U$60094 ( \60471 , \60393 , \60362 );
nand \U$60095 ( \60472 , \60470 , \60471 );
not \U$60096 ( \60473 , \60472 );
not \U$60097 ( \60474 , \60342 );
and \U$60098 ( \60475 , \60473 , \60474 );
and \U$60099 ( \60476 , \60472 , \60342 );
nor \U$60100 ( \60477 , \60475 , \60476 );
xor \U$60101 ( \60478 , \60467 , \60477 );
not \U$60102 ( \60479 , \60478 );
and \U$60103 ( \60480 , \15726 , RIae77900_86);
and \U$60104 ( \60481 , RIae76fa0_66, RIae7aab0_192);
nor \U$60105 ( \60482 , \60480 , \60481 );
and \U$60106 ( \60483 , \60482 , \14959 );
not \U$60107 ( \60484 , \60482 );
and \U$60108 ( \60485 , \60484 , RIae7aa38_191);
nor \U$60109 ( \60486 , \60483 , \60485 );
and \U$60110 ( \60487 , \60486 , \11827 );
not \U$60111 ( \60488 , \60486 );
not \U$60112 ( \60489 , \11827 );
and \U$60113 ( \60490 , \60488 , \60489 );
and \U$60114 ( \60491 , \14964 , RIae779f0_88);
and \U$60115 ( \60492 , RIae77810_84, \14962 );
nor \U$60116 ( \60493 , \60491 , \60492 );
and \U$60117 ( \60494 , \60493 , \14462 );
not \U$60118 ( \60495 , \60493 );
and \U$60119 ( \60496 , \60495 , \14463 );
nor \U$60120 ( \60497 , \60494 , \60496 );
nor \U$60121 ( \60498 , \60490 , \60497 );
nor \U$60122 ( \60499 , \60487 , \60498 );
and \U$60123 ( \60500 , \13059 , RIae776a8_81);
and \U$60124 ( \60501 , RIae77450_76, \13057 );
nor \U$60125 ( \60502 , \60500 , \60501 );
and \U$60126 ( \60503 , \60502 , \12718 );
not \U$60127 ( \60504 , \60502 );
and \U$60128 ( \60505 , \60504 , \13063 );
nor \U$60129 ( \60506 , \60503 , \60505 );
or \U$60130 ( \60507 , \60499 , \60506 );
not \U$60131 ( \60508 , \60506 );
not \U$60132 ( \60509 , \60499 );
or \U$60133 ( \60510 , \60508 , \60509 );
and \U$60134 ( \60511 , \13059 , RIae77540_78);
and \U$60135 ( \60512 , RIae776a8_81, \13057 );
nor \U$60136 ( \60513 , \60511 , \60512 );
and \U$60137 ( \60514 , \60513 , \13063 );
not \U$60138 ( \60515 , \60513 );
and \U$60139 ( \60516 , \60515 , \12718 );
nor \U$60140 ( \60517 , \60514 , \60516 );
nand \U$60141 ( \60518 , RIae77630_80, \12178 );
and \U$60142 ( \60519 , \60518 , \12184 );
not \U$60143 ( \60520 , \60518 );
and \U$60144 ( \60521 , \60520 , \11827 );
nor \U$60145 ( \60522 , \60519 , \60521 );
xor \U$60146 ( \60523 , \60517 , \60522 );
and \U$60147 ( \60524 , \14059 , RIae77450_76);
and \U$60148 ( \60525 , RIae77ae0_90, \14057 );
nor \U$60149 ( \60526 , \60524 , \60525 );
and \U$60150 ( \60527 , \60526 , \13502 );
not \U$60151 ( \60528 , \60526 );
and \U$60152 ( \60529 , \60528 , \14063 );
nor \U$60153 ( \60530 , \60527 , \60529 );
and \U$60154 ( \60531 , \60523 , \60530 );
and \U$60155 ( \60532 , \60517 , \60522 );
or \U$60156 ( \60533 , \60531 , \60532 );
nand \U$60157 ( \60534 , \60510 , \60533 );
nand \U$60158 ( \60535 , \60507 , \60534 );
not \U$60159 ( \60536 , \10936 );
not \U$60160 ( \60537 , \60349 );
not \U$60161 ( \60538 , \60360 );
or \U$60162 ( \60539 , \60537 , \60538 );
or \U$60163 ( \60540 , \60360 , \60349 );
nand \U$60164 ( \60541 , \60539 , \60540 );
not \U$60165 ( \60542 , \60541 );
or \U$60166 ( \60543 , \60536 , \60542 );
or \U$60167 ( \60544 , \60541 , \10936 );
nand \U$60168 ( \60545 , \60543 , \60544 );
xor \U$60169 ( \60546 , \60535 , \60545 );
and \U$60170 ( \60547 , \12180 , RIae77630_80);
and \U$60171 ( \60548 , RIae77540_78, \12178 );
nor \U$60172 ( \60549 , \60547 , \60548 );
and \U$60173 ( \60550 , \60549 , \12184 );
not \U$60174 ( \60551 , \60549 );
and \U$60175 ( \60552 , \60551 , \11827 );
nor \U$60176 ( \60553 , \60550 , \60552 );
xor \U$60177 ( \60554 , \60427 , \60434 );
xor \U$60178 ( \60555 , \60554 , \60442 );
and \U$60179 ( \60556 , \60553 , \60555 );
and \U$60180 ( \60557 , \60546 , \60556 );
and \U$60181 ( \60558 , \60535 , \60545 );
or \U$60182 ( \60559 , \60557 , \60558 );
not \U$60183 ( \60560 , \60559 );
and \U$60184 ( \60561 , \60479 , \60560 );
and \U$60185 ( \60562 , \60478 , \60559 );
nor \U$60186 ( \60563 , \60561 , \60562 );
xor \U$60187 ( \60564 , \60445 , \60450 );
xor \U$60188 ( \60565 , \60564 , \60461 );
not \U$60189 ( \60566 , \60565 );
xor \U$60190 ( \60567 , \60535 , \60545 );
xor \U$60191 ( \60568 , \60567 , \60556 );
nand \U$60192 ( \60569 , \60566 , \60568 );
or \U$60193 ( \60570 , \60563 , \60569 );
xnor \U$60194 ( \60571 , \60569 , \60563 );
nand \U$60195 ( \60572 , RIae77630_80, \13057 );
and \U$60196 ( \60573 , \60572 , \13063 );
not \U$60197 ( \60574 , \60572 );
and \U$60198 ( \60575 , \60574 , \12718 );
nor \U$60199 ( \60576 , \60573 , \60575 );
not \U$60200 ( \60577 , \60576 );
and \U$60201 ( \60578 , \14059 , RIae77540_78);
and \U$60202 ( \60579 , RIae776a8_81, \14057 );
nor \U$60203 ( \60580 , \60578 , \60579 );
and \U$60204 ( \60581 , \60580 , \14063 );
not \U$60205 ( \60582 , \60580 );
and \U$60206 ( \60583 , \60582 , \13502 );
nor \U$60207 ( \60584 , \60581 , \60583 );
not \U$60208 ( \60585 , \60584 );
or \U$60209 ( \60586 , \60577 , \60585 );
or \U$60210 ( \60587 , \60584 , \60576 );
nand \U$60211 ( \60588 , \60586 , \60587 );
and \U$60212 ( \60589 , \14059 , RIae77630_80);
and \U$60213 ( \60590 , RIae77540_78, \14057 );
nor \U$60214 ( \60591 , \60589 , \60590 );
and \U$60215 ( \60592 , \60591 , \14063 );
not \U$60216 ( \60593 , \60591 );
and \U$60217 ( \60594 , \60593 , \13502 );
nor \U$60218 ( \60595 , \60592 , \60594 );
and \U$60219 ( \60596 , \15726 , RIae77ae0_90);
and \U$60220 ( \60597 , RIae779f0_88, RIae7aab0_192);
nor \U$60221 ( \60598 , \60596 , \60597 );
and \U$60222 ( \60599 , \60598 , RIae7aa38_191);
not \U$60223 ( \60600 , \60598 );
and \U$60224 ( \60601 , \60600 , \14959 );
nor \U$60225 ( \60602 , \60599 , \60601 );
or \U$60226 ( \60603 , \60595 , \60602 );
not \U$60227 ( \60604 , \60602 );
not \U$60228 ( \60605 , \60595 );
or \U$60229 ( \60606 , \60604 , \60605 );
and \U$60230 ( \60607 , \14964 , RIae776a8_81);
and \U$60231 ( \60608 , RIae77450_76, \14962 );
nor \U$60232 ( \60609 , \60607 , \60608 );
and \U$60233 ( \60610 , \60609 , \14463 );
not \U$60234 ( \60611 , \60609 );
and \U$60235 ( \60612 , \60611 , \14462 );
nor \U$60236 ( \60613 , \60610 , \60612 );
nand \U$60237 ( \60614 , \60606 , \60613 );
nand \U$60238 ( \60615 , \60603 , \60614 );
xor \U$60239 ( \60616 , \60588 , \60615 );
and \U$60240 ( \60617 , \15726 , RIae779f0_88);
and \U$60241 ( \60618 , RIae77810_84, RIae7aab0_192);
nor \U$60242 ( \60619 , \60617 , \60618 );
and \U$60243 ( \60620 , \60619 , \14959 );
not \U$60244 ( \60621 , \60619 );
and \U$60245 ( \60622 , \60621 , RIae7aa38_191);
nor \U$60246 ( \60623 , \60620 , \60622 );
xor \U$60247 ( \60624 , \60623 , \12718 );
and \U$60248 ( \60625 , \14964 , RIae77450_76);
and \U$60249 ( \60626 , RIae77ae0_90, \14962 );
nor \U$60250 ( \60627 , \60625 , \60626 );
and \U$60251 ( \60628 , \60627 , \14463 );
not \U$60252 ( \60629 , \60627 );
and \U$60253 ( \60630 , \60629 , \14462 );
nor \U$60254 ( \60631 , \60628 , \60630 );
xor \U$60255 ( \60632 , \60624 , \60631 );
and \U$60256 ( \60633 , \60616 , \60632 );
and \U$60257 ( \60634 , \60588 , \60615 );
nor \U$60258 ( \60635 , \60633 , \60634 );
and \U$60259 ( \60636 , \13059 , RIae77630_80);
and \U$60260 ( \60637 , RIae77540_78, \13057 );
nor \U$60261 ( \60638 , \60636 , \60637 );
and \U$60262 ( \60639 , \60638 , \12718 );
not \U$60263 ( \60640 , \60638 );
and \U$60264 ( \60641 , \60640 , \13063 );
nor \U$60265 ( \60642 , \60639 , \60641 );
not \U$60266 ( \60643 , \60642 );
not \U$60267 ( \60644 , \60584 );
nand \U$60268 ( \60645 , \60644 , \60576 );
not \U$60269 ( \60646 , \60645 );
xor \U$60270 ( \60647 , \60623 , \12718 );
and \U$60271 ( \60648 , \60647 , \60631 );
and \U$60272 ( \60649 , \60623 , \12718 );
or \U$60273 ( \60650 , \60648 , \60649 );
not \U$60274 ( \60651 , \60650 );
or \U$60275 ( \60652 , \60646 , \60651 );
or \U$60276 ( \60653 , \60650 , \60645 );
nand \U$60277 ( \60654 , \60652 , \60653 );
not \U$60278 ( \60655 , \60654 );
or \U$60279 ( \60656 , \60643 , \60655 );
or \U$60280 ( \60657 , \60654 , \60642 );
nand \U$60281 ( \60658 , \60656 , \60657 );
not \U$60282 ( \60659 , \60658 );
and \U$60283 ( \60660 , \15726 , RIae77810_84);
and \U$60284 ( \60661 , RIae77900_86, RIae7aab0_192);
nor \U$60285 ( \60662 , \60660 , \60661 );
and \U$60286 ( \60663 , \60662 , RIae7aa38_191);
not \U$60287 ( \60664 , \60662 );
and \U$60288 ( \60665 , \60664 , \14959 );
nor \U$60289 ( \60666 , \60663 , \60665 );
and \U$60290 ( \60667 , \14964 , RIae77ae0_90);
and \U$60291 ( \60668 , RIae779f0_88, \14962 );
nor \U$60292 ( \60669 , \60667 , \60668 );
and \U$60293 ( \60670 , \60669 , \14462 );
not \U$60294 ( \60671 , \60669 );
and \U$60295 ( \60672 , \60671 , \14463 );
nor \U$60296 ( \60673 , \60670 , \60672 );
xor \U$60297 ( \60674 , \60666 , \60673 );
and \U$60298 ( \60675 , \14059 , RIae776a8_81);
and \U$60299 ( \60676 , RIae77450_76, \14057 );
nor \U$60300 ( \60677 , \60675 , \60676 );
and \U$60301 ( \60678 , \60677 , \14063 );
not \U$60302 ( \60679 , \60677 );
and \U$60303 ( \60680 , \60679 , \13502 );
nor \U$60304 ( \60681 , \60678 , \60680 );
xor \U$60305 ( \60682 , \60674 , \60681 );
not \U$60306 ( \60683 , \60682 );
and \U$60307 ( \60684 , \60659 , \60683 );
and \U$60308 ( \60685 , \60658 , \60682 );
nor \U$60309 ( \60686 , \60684 , \60685 );
xor \U$60310 ( \60687 , \60635 , \60686 );
and \U$60311 ( \60688 , \14964 , RIae77630_80);
and \U$60312 ( \60689 , RIae77540_78, \14962 );
nor \U$60313 ( \60690 , \60688 , \60689 );
and \U$60314 ( \60691 , \60690 , \14463 );
not \U$60315 ( \60692 , \60690 );
and \U$60316 ( \60693 , \60692 , \14462 );
nor \U$60317 ( \60694 , \60691 , \60693 );
not \U$60318 ( \60695 , \60694 );
and \U$60319 ( \60696 , \15726 , RIae776a8_81);
and \U$60320 ( \60697 , RIae77450_76, RIae7aab0_192);
nor \U$60321 ( \60698 , \60696 , \60697 );
and \U$60322 ( \60699 , \60698 , RIae7aa38_191);
not \U$60323 ( \60700 , \60698 );
and \U$60324 ( \60701 , \60700 , \14959 );
nor \U$60325 ( \60702 , \60699 , \60701 );
nor \U$60326 ( \60703 , \60695 , \60702 );
nand \U$60327 ( \60704 , RIae77630_80, \14057 );
and \U$60328 ( \60705 , \60704 , \14063 );
not \U$60329 ( \60706 , \60704 );
and \U$60330 ( \60707 , \60706 , \13502 );
nor \U$60331 ( \60708 , \60705 , \60707 );
not \U$60332 ( \60709 , \60708 );
and \U$60333 ( \60710 , \15726 , RIae77450_76);
and \U$60334 ( \60711 , RIae77ae0_90, RIae7aab0_192);
nor \U$60335 ( \60712 , \60710 , \60711 );
and \U$60336 ( \60713 , \60712 , \14959 );
not \U$60337 ( \60714 , \60712 );
and \U$60338 ( \60715 , \60714 , RIae7aa38_191);
nor \U$60339 ( \60716 , \60713 , \60715 );
xor \U$60340 ( \60717 , \60716 , \14063 );
and \U$60341 ( \60718 , \14964 , RIae77540_78);
and \U$60342 ( \60719 , RIae776a8_81, \14962 );
nor \U$60343 ( \60720 , \60718 , \60719 );
and \U$60344 ( \60721 , \60720 , \14463 );
not \U$60345 ( \60722 , \60720 );
and \U$60346 ( \60723 , \60722 , \14462 );
nor \U$60347 ( \60724 , \60721 , \60723 );
xor \U$60348 ( \60725 , \60717 , \60724 );
not \U$60349 ( \60726 , \60725 );
or \U$60350 ( \60727 , \60709 , \60726 );
or \U$60351 ( \60728 , \60725 , \60708 );
nand \U$60352 ( \60729 , \60727 , \60728 );
xor \U$60353 ( \60730 , \60703 , \60729 );
and \U$60354 ( \60731 , \15726 , RIae77540_78);
and \U$60355 ( \60732 , RIae776a8_81, RIae7aab0_192);
nor \U$60356 ( \60733 , \60731 , \60732 );
and \U$60357 ( \60734 , \60733 , \14959 );
not \U$60358 ( \60735 , \60733 );
and \U$60359 ( \60736 , \60735 , RIae7aa38_191);
nor \U$60360 ( \60737 , \60734 , \60736 );
nand \U$60361 ( \60738 , \14462 , \60737 );
not \U$60362 ( \60739 , \60694 );
not \U$60363 ( \60740 , \60702 );
and \U$60364 ( \60741 , \60739 , \60740 );
and \U$60365 ( \60742 , \60694 , \60702 );
nor \U$60366 ( \60743 , \60741 , \60742 );
xnor \U$60367 ( \60744 , \60738 , \60743 );
nand \U$60368 ( \60745 , RIae77630_80, \14962 );
and \U$60369 ( \60746 , \60745 , \14463 );
not \U$60370 ( \60747 , \60745 );
and \U$60371 ( \60748 , \60747 , \14462 );
nor \U$60372 ( \60749 , \60746 , \60748 );
and \U$60373 ( \60750 , \60737 , \14462 );
not \U$60374 ( \60751 , \60737 );
and \U$60375 ( \60752 , \60751 , \14463 );
nor \U$60376 ( \60753 , \60750 , \60752 );
xor \U$60377 ( \60754 , \60749 , \60753 );
and \U$60378 ( \60755 , \15726 , RIae77630_80);
and \U$60379 ( \60756 , RIae77540_78, RIae7aab0_192);
nor \U$60380 ( \60757 , \60755 , \60756 );
and \U$60381 ( \60758 , \60757 , RIae7aa38_191);
not \U$60382 ( \60759 , \60757 );
and \U$60383 ( \60760 , \60759 , \14959 );
nor \U$60384 ( \60761 , \60758 , \60760 );
nand \U$60385 ( \60762 , RIae77630_80, RIae7aab0_192);
nand \U$60386 ( \60763 , RIae7aa38_191, \60762 );
nor \U$60387 ( \60764 , \60761 , \60763 );
and \U$60388 ( \60765 , \60754 , \60764 );
and \U$60389 ( \60766 , \60749 , \60753 );
nor \U$60390 ( \60767 , \60765 , \60766 );
or \U$60391 ( \60768 , \60744 , \60767 );
or \U$60392 ( \60769 , \60738 , \60743 );
nand \U$60393 ( \60770 , \60768 , \60769 );
and \U$60394 ( \60771 , \60730 , \60770 );
and \U$60395 ( \60772 , \60703 , \60729 );
nor \U$60396 ( \60773 , \60771 , \60772 );
not \U$60397 ( \60774 , \60708 );
nand \U$60398 ( \60775 , \60774 , \60725 );
not \U$60399 ( \60776 , \60602 );
not \U$60400 ( \60777 , \60613 );
or \U$60401 ( \60778 , \60776 , \60777 );
or \U$60402 ( \60779 , \60613 , \60602 );
nand \U$60403 ( \60780 , \60778 , \60779 );
not \U$60404 ( \60781 , \60780 );
not \U$60405 ( \60782 , \60595 );
and \U$60406 ( \60783 , \60781 , \60782 );
and \U$60407 ( \60784 , \60780 , \60595 );
nor \U$60408 ( \60785 , \60783 , \60784 );
not \U$60409 ( \60786 , \60785 );
xor \U$60410 ( \60787 , \60716 , \14063 );
and \U$60411 ( \60788 , \60787 , \60724 );
and \U$60412 ( \60789 , \60716 , \14063 );
or \U$60413 ( \60790 , \60788 , \60789 );
not \U$60414 ( \60791 , \60790 );
and \U$60415 ( \60792 , \60786 , \60791 );
and \U$60416 ( \60793 , \60785 , \60790 );
nor \U$60417 ( \60794 , \60792 , \60793 );
xnor \U$60418 ( \60795 , \60775 , \60794 );
or \U$60419 ( \60796 , \60773 , \60795 );
or \U$60420 ( \60797 , \60775 , \60794 );
nand \U$60421 ( \60798 , \60796 , \60797 );
not \U$60422 ( \60799 , \60790 );
nor \U$60423 ( \60800 , \60799 , \60785 );
xor \U$60424 ( \60801 , \60588 , \60615 );
xor \U$60425 ( \60802 , \60801 , \60632 );
xor \U$60426 ( \60803 , \60800 , \60802 );
and \U$60427 ( \60804 , \60798 , \60803 );
and \U$60428 ( \60805 , \60800 , \60802 );
nor \U$60429 ( \60806 , \60804 , \60805 );
and \U$60430 ( \60807 , \60687 , \60806 );
and \U$60431 ( \60808 , \60635 , \60686 );
nor \U$60432 ( \60809 , \60807 , \60808 );
not \U$60433 ( \60810 , \60658 );
nor \U$60434 ( \60811 , \60810 , \60682 );
not \U$60435 ( \60812 , \60645 );
not \U$60436 ( \60813 , \60642 );
and \U$60437 ( \60814 , \60812 , \60813 );
and \U$60438 ( \60815 , \60645 , \60642 );
not \U$60439 ( \60816 , \60650 );
nor \U$60440 ( \60817 , \60815 , \60816 );
nor \U$60441 ( \60818 , \60814 , \60817 );
not \U$60442 ( \60819 , \60818 );
not \U$60443 ( \60820 , \60486 );
not \U$60444 ( \60821 , \60497 );
or \U$60445 ( \60822 , \60820 , \60821 );
or \U$60446 ( \60823 , \60497 , \60486 );
nand \U$60447 ( \60824 , \60822 , \60823 );
and \U$60448 ( \60825 , \60824 , \11827 );
not \U$60449 ( \60826 , \60824 );
and \U$60450 ( \60827 , \60826 , \12184 );
nor \U$60451 ( \60828 , \60825 , \60827 );
xor \U$60452 ( \60829 , \60666 , \60673 );
and \U$60453 ( \60830 , \60829 , \60681 );
and \U$60454 ( \60831 , \60666 , \60673 );
nor \U$60455 ( \60832 , \60830 , \60831 );
xor \U$60456 ( \60833 , \60828 , \60832 );
xor \U$60457 ( \60834 , \60517 , \60522 );
xor \U$60458 ( \60835 , \60834 , \60530 );
xor \U$60459 ( \60836 , \60833 , \60835 );
not \U$60460 ( \60837 , \60836 );
or \U$60461 ( \60838 , \60819 , \60837 );
or \U$60462 ( \60839 , \60836 , \60818 );
nand \U$60463 ( \60840 , \60838 , \60839 );
xor \U$60464 ( \60841 , \60811 , \60840 );
and \U$60465 ( \60842 , \60809 , \60841 );
and \U$60466 ( \60843 , \60811 , \60840 );
nor \U$60467 ( \60844 , \60842 , \60843 );
not \U$60468 ( \60845 , \60818 );
nand \U$60469 ( \60846 , \60845 , \60836 );
not \U$60470 ( \60847 , \60499 );
not \U$60471 ( \60848 , \60533 );
or \U$60472 ( \60849 , \60847 , \60848 );
or \U$60473 ( \60850 , \60533 , \60499 );
nand \U$60474 ( \60851 , \60849 , \60850 );
not \U$60475 ( \60852 , \60851 );
not \U$60476 ( \60853 , \60506 );
and \U$60477 ( \60854 , \60852 , \60853 );
and \U$60478 ( \60855 , \60851 , \60506 );
nor \U$60479 ( \60856 , \60854 , \60855 );
not \U$60480 ( \60857 , \60856 );
xor \U$60481 ( \60858 , \60828 , \60832 );
and \U$60482 ( \60859 , \60858 , \60835 );
and \U$60483 ( \60860 , \60828 , \60832 );
or \U$60484 ( \60861 , \60859 , \60860 );
not \U$60485 ( \60862 , \60861 );
and \U$60486 ( \60863 , \60857 , \60862 );
and \U$60487 ( \60864 , \60856 , \60861 );
nor \U$60488 ( \60865 , \60863 , \60864 );
not \U$60489 ( \60866 , \60865 );
xor \U$60490 ( \60867 , \60553 , \60555 );
not \U$60491 ( \60868 , \60867 );
and \U$60492 ( \60869 , \60866 , \60868 );
and \U$60493 ( \60870 , \60865 , \60867 );
nor \U$60494 ( \60871 , \60869 , \60870 );
xnor \U$60495 ( \60872 , \60846 , \60871 );
or \U$60496 ( \60873 , \60844 , \60872 );
or \U$60497 ( \60874 , \60846 , \60871 );
nand \U$60498 ( \60875 , \60873 , \60874 );
not \U$60499 ( \60876 , \60867 );
or \U$60500 ( \60877 , \60856 , \60876 );
not \U$60501 ( \60878 , \60876 );
not \U$60502 ( \60879 , \60856 );
or \U$60503 ( \60880 , \60878 , \60879 );
nand \U$60504 ( \60881 , \60880 , \60861 );
nand \U$60505 ( \60882 , \60877 , \60881 );
not \U$60506 ( \60883 , \60565 );
not \U$60507 ( \60884 , \60568 );
or \U$60508 ( \60885 , \60883 , \60884 );
or \U$60509 ( \60886 , \60568 , \60565 );
nand \U$60510 ( \60887 , \60885 , \60886 );
xor \U$60511 ( \60888 , \60882 , \60887 );
and \U$60512 ( \60889 , \60875 , \60888 );
and \U$60513 ( \60890 , \60882 , \60887 );
nor \U$60514 ( \60891 , \60889 , \60890 );
or \U$60515 ( \60892 , \60571 , \60891 );
nand \U$60516 ( \60893 , \60570 , \60892 );
not \U$60517 ( \60894 , \60559 );
nor \U$60518 ( \60895 , \60894 , \60478 );
xor \U$60519 ( \60896 , \60464 , \60466 );
and \U$60520 ( \60897 , \60896 , \60477 );
and \U$60521 ( \60898 , \60464 , \60466 );
or \U$60522 ( \60899 , \60897 , \60898 );
not \U$60523 ( \60900 , \60899 );
xor \U$60524 ( \60901 , \60272 , \60279 );
xor \U$60525 ( \60902 , \60901 , \60307 );
xor \U$60526 ( \60903 , \60395 , \60402 );
xor \U$60527 ( \60904 , \60902 , \60903 );
not \U$60528 ( \60905 , \60904 );
or \U$60529 ( \60906 , \60900 , \60905 );
or \U$60530 ( \60907 , \60904 , \60899 );
nand \U$60531 ( \60908 , \60906 , \60907 );
xor \U$60532 ( \60909 , \60895 , \60908 );
and \U$60533 ( \60910 , \60893 , \60909 );
and \U$60534 ( \60911 , \60895 , \60908 );
nor \U$60535 ( \60912 , \60910 , \60911 );
not \U$60536 ( \60913 , \60899 );
nand \U$60537 ( \60914 , \60913 , \60904 );
xnor \U$60538 ( \60915 , \60407 , \60329 );
not \U$60539 ( \60916 , \60915 );
not \U$60540 ( \60917 , \60246 );
and \U$60541 ( \60918 , \60916 , \60917 );
and \U$60542 ( \60919 , \60915 , \60246 );
nor \U$60543 ( \60920 , \60918 , \60919 );
xnor \U$60544 ( \60921 , \60914 , \60920 );
or \U$60545 ( \60922 , \60912 , \60921 );
or \U$60546 ( \60923 , \60914 , \60920 );
nand \U$60547 ( \60924 , \60922 , \60923 );
and \U$60548 ( \60925 , \60420 , \60924 );
nor \U$60549 ( \60926 , \60419 , \60925 );
not \U$60550 ( \60927 , \60168 );
not \U$60551 ( \60928 , \60237 );
or \U$60552 ( \60929 , \60927 , \60928 );
or \U$60553 ( \60930 , \60237 , \60168 );
nand \U$60554 ( \60931 , \60929 , \60930 );
not \U$60555 ( \60932 , \60931 );
not \U$60556 ( \60933 , \60158 );
and \U$60557 ( \60934 , \60932 , \60933 );
and \U$60558 ( \60935 , \60931 , \60158 );
nor \U$60559 ( \60936 , \60934 , \60935 );
xor \U$60560 ( \60937 , \60411 , \60412 );
and \U$60561 ( \60938 , \60937 , \60417 );
and \U$60562 ( \60939 , \60411 , \60412 );
nor \U$60563 ( \60940 , \60938 , \60939 );
xnor \U$60564 ( \60941 , \60936 , \60940 );
or \U$60565 ( \60942 , \60926 , \60941 );
or \U$60566 ( \60943 , \60940 , \60936 );
nand \U$60567 ( \60944 , \60942 , \60943 );
and \U$60568 ( \60945 , \60241 , \60944 );
nor \U$60569 ( \60946 , \60240 , \60945 );
or \U$60570 ( \60947 , \60146 , \60946 );
nand \U$60571 ( \60948 , \60145 , \60947 );
not \U$60572 ( \60949 , \59955 );
nor \U$60573 ( \60950 , \60949 , \60051 );
xor \U$60574 ( \60951 , \59826 , \59854 );
and \U$60575 ( \60952 , \60951 , \59954 );
and \U$60576 ( \60953 , \59826 , \59854 );
or \U$60577 ( \60954 , \60952 , \60953 );
not \U$60578 ( \60955 , \60954 );
xor \U$60579 ( \60956 , \59830 , \59848 );
and \U$60580 ( \60957 , \60956 , \59853 );
and \U$60581 ( \60958 , \59830 , \59848 );
or \U$60582 ( \60959 , \60957 , \60958 );
xor \U$60583 ( \60960 , \59642 , \59649 );
xor \U$60584 ( \60961 , \60960 , \59657 );
xor \U$60585 ( \60962 , \60959 , \60961 );
or \U$60586 ( \60963 , \60018 , \60046 );
not \U$60587 ( \60964 , \60046 );
not \U$60588 ( \60965 , \60018 );
or \U$60589 ( \60966 , \60964 , \60965 );
nand \U$60590 ( \60967 , \60966 , \59994 );
nand \U$60591 ( \60968 , \60963 , \60967 );
xor \U$60592 ( \60969 , \60962 , \60968 );
xor \U$60593 ( \60970 , \59962 , \59966 );
and \U$60594 ( \60971 , \60970 , \60050 );
and \U$60595 ( \60972 , \59962 , \59966 );
nor \U$60596 ( \60973 , \60971 , \60972 );
xnor \U$60597 ( \60974 , \60969 , \60973 );
not \U$60598 ( \60975 , \60974 );
and \U$60599 ( \60976 , \8966 , RIae77540_78);
and \U$60600 ( \60977 , RIae776a8_81, \8964 );
nor \U$60601 ( \60978 , \60976 , \60977 );
and \U$60602 ( \60979 , \60978 , \8799 );
not \U$60603 ( \60980 , \60978 );
and \U$60604 ( \60981 , \60980 , \8789 );
nor \U$60605 ( \60982 , \60979 , \60981 );
nand \U$60606 ( \60983 , RIae77630_80, \8369 );
and \U$60607 ( \60984 , \60983 , \8020 );
not \U$60608 ( \60985 , \60983 );
and \U$60609 ( \60986 , \60985 , \8019 );
nor \U$60610 ( \60987 , \60984 , \60986 );
xor \U$60611 ( \60988 , \60982 , \60987 );
xor \U$60612 ( \60989 , \59598 , \59605 );
xor \U$60613 ( \60990 , \60989 , \59613 );
xor \U$60614 ( \60991 , \60988 , \60990 );
not \U$60615 ( \60992 , \60991 );
xor \U$60616 ( \60993 , \60002 , \60009 );
and \U$60617 ( \60994 , \60993 , \60017 );
and \U$60618 ( \60995 , \60002 , \60009 );
or \U$60619 ( \60996 , \60994 , \60995 );
not \U$60620 ( \60997 , \59974 );
not \U$60621 ( \60998 , \59989 );
and \U$60622 ( \60999 , \60997 , \60998 );
and \U$60623 ( \61000 , \59989 , \59974 );
nor \U$60624 ( \61001 , \61000 , \59982 );
nor \U$60625 ( \61002 , \60999 , \61001 );
xor \U$60626 ( \61003 , \60996 , \61002 );
xor \U$60627 ( \61004 , \60030 , \60037 );
and \U$60628 ( \61005 , \61004 , \60045 );
and \U$60629 ( \61006 , \60030 , \60037 );
or \U$60630 ( \61007 , \61005 , \61006 );
xor \U$60631 ( \61008 , \61003 , \61007 );
not \U$60632 ( \61009 , \61008 );
xor \U$60633 ( \61010 , \59623 , \8019 );
xor \U$60634 ( \61011 , \61010 , \59631 );
not \U$60635 ( \61012 , \61011 );
and \U$60636 ( \61013 , \61009 , \61012 );
and \U$60637 ( \61014 , \61008 , \61011 );
nor \U$60638 ( \61015 , \61013 , \61014 );
not \U$60639 ( \61016 , \61015 );
or \U$60640 ( \61017 , \60992 , \61016 );
or \U$60641 ( \61018 , \61015 , \60991 );
nand \U$60642 ( \61019 , \61017 , \61018 );
not \U$60643 ( \61020 , \61019 );
and \U$60644 ( \61021 , \60975 , \61020 );
and \U$60645 ( \61022 , \60974 , \61019 );
nor \U$60646 ( \61023 , \61021 , \61022 );
not \U$60647 ( \61024 , \61023 );
or \U$60648 ( \61025 , \60955 , \61024 );
or \U$60649 ( \61026 , \61023 , \60954 );
nand \U$60650 ( \61027 , \61025 , \61026 );
xor \U$60651 ( \61028 , \60950 , \61027 );
and \U$60652 ( \61029 , \60948 , \61028 );
and \U$60653 ( \61030 , \60950 , \61027 );
nor \U$60654 ( \61031 , \61029 , \61030 );
not \U$60655 ( \61032 , \61023 );
nand \U$60656 ( \61033 , \61032 , \60954 );
not \U$60657 ( \61034 , \60969 );
not \U$60658 ( \61035 , \61019 );
or \U$60659 ( \61036 , \61034 , \61035 );
or \U$60660 ( \61037 , \61019 , \60969 );
nand \U$60661 ( \61038 , \61037 , \60973 );
nand \U$60662 ( \61039 , \61036 , \61038 );
not \U$60663 ( \61040 , \61039 );
xor \U$60664 ( \61041 , \60959 , \60961 );
and \U$60665 ( \61042 , \61041 , \60968 );
and \U$60666 ( \61043 , \60959 , \60961 );
or \U$60667 ( \61044 , \61042 , \61043 );
not \U$60668 ( \61045 , \61044 );
and \U$60669 ( \61046 , \60991 , \61011 );
not \U$60670 ( \61047 , \60991 );
not \U$60671 ( \61048 , \61011 );
and \U$60672 ( \61049 , \61047 , \61048 );
nor \U$60673 ( \61050 , \61049 , \61008 );
nor \U$60674 ( \61051 , \61046 , \61050 );
not \U$60675 ( \61052 , \61051 );
or \U$60676 ( \61053 , \61045 , \61052 );
or \U$60677 ( \61054 , \61051 , \61044 );
nand \U$60678 ( \61055 , \61053 , \61054 );
not \U$60679 ( \61056 , \61055 );
xor \U$60680 ( \61057 , \59673 , \59675 );
xor \U$60681 ( \61058 , \61057 , \59678 );
not \U$60682 ( \61059 , \61058 );
and \U$60683 ( \61060 , \61056 , \61059 );
and \U$60684 ( \61061 , \61055 , \61058 );
nor \U$60685 ( \61062 , \61060 , \61061 );
not \U$60686 ( \61063 , \61062 );
and \U$60687 ( \61064 , \61040 , \61063 );
and \U$60688 ( \61065 , \61039 , \61062 );
nor \U$60689 ( \61066 , \61064 , \61065 );
not \U$60690 ( \61067 , \61066 );
xor \U$60691 ( \61068 , \59616 , \59634 );
xor \U$60692 ( \61069 , \61068 , \59660 );
xor \U$60693 ( \61070 , \60982 , \60987 );
and \U$60694 ( \61071 , \61070 , \60990 );
and \U$60695 ( \61072 , \60982 , \60987 );
or \U$60696 ( \61073 , \61071 , \61072 );
xor \U$60697 ( \61074 , \59500 , \59507 );
xor \U$60698 ( \61075 , \61074 , \59515 );
xor \U$60699 ( \61076 , \61073 , \61075 );
xor \U$60700 ( \61077 , \60996 , \61002 );
and \U$60701 ( \61078 , \61077 , \61007 );
and \U$60702 ( \61079 , \60996 , \61002 );
nor \U$60703 ( \61080 , \61078 , \61079 );
xor \U$60704 ( \61081 , \61076 , \61080 );
xor \U$60705 ( \61082 , \61069 , \61081 );
not \U$60706 ( \61083 , \61082 );
and \U$60707 ( \61084 , \61067 , \61083 );
and \U$60708 ( \61085 , \61066 , \61082 );
nor \U$60709 ( \61086 , \61084 , \61085 );
xnor \U$60710 ( \61087 , \61033 , \61086 );
or \U$60711 ( \61088 , \61031 , \61087 );
or \U$60712 ( \61089 , \61033 , \61086 );
nand \U$60713 ( \61090 , \61088 , \61089 );
not \U$60714 ( \61091 , \61082 );
or \U$60715 ( \61092 , \61062 , \61091 );
not \U$60716 ( \61093 , \61091 );
not \U$60717 ( \61094 , \61062 );
or \U$60718 ( \61095 , \61093 , \61094 );
nand \U$60719 ( \61096 , \61095 , \61039 );
nand \U$60720 ( \61097 , \61092 , \61096 );
xor \U$60721 ( \61098 , \59583 , \59587 );
xor \U$60722 ( \61099 , \61073 , \61075 );
and \U$60723 ( \61100 , \61099 , \61080 );
and \U$60724 ( \61101 , \61073 , \61075 );
or \U$60725 ( \61102 , \61100 , \61101 );
xor \U$60726 ( \61103 , \61098 , \61102 );
xor \U$60727 ( \61104 , \59663 , \59665 );
xor \U$60728 ( \61105 , \61104 , \59681 );
xor \U$60729 ( \61106 , \61103 , \61105 );
and \U$60730 ( \61107 , \61069 , \61081 );
xor \U$60731 ( \61108 , \61106 , \61107 );
or \U$60732 ( \61109 , \61051 , \61058 );
not \U$60733 ( \61110 , \61058 );
not \U$60734 ( \61111 , \61051 );
or \U$60735 ( \61112 , \61110 , \61111 );
nand \U$60736 ( \61113 , \61112 , \61044 );
nand \U$60737 ( \61114 , \61109 , \61113 );
xor \U$60738 ( \61115 , \61108 , \61114 );
xor \U$60739 ( \61116 , \61097 , \61115 );
and \U$60740 ( \61117 , \61090 , \61116 );
and \U$60741 ( \61118 , \61097 , \61115 );
nor \U$60742 ( \61119 , \61117 , \61118 );
xor \U$60743 ( \61120 , \61106 , \61107 );
and \U$60744 ( \61121 , \61120 , \61114 );
and \U$60745 ( \61122 , \61106 , \61107 );
nor \U$60746 ( \61123 , \61121 , \61122 );
xor \U$60747 ( \61124 , \59588 , \59590 );
xor \U$60748 ( \61125 , \61124 , \59684 );
xor \U$60749 ( \61126 , \61098 , \61102 );
and \U$60750 ( \61127 , \61126 , \61105 );
and \U$60751 ( \61128 , \61098 , \61102 );
or \U$60752 ( \61129 , \61127 , \61128 );
xnor \U$60753 ( \61130 , \61125 , \61129 );
not \U$60754 ( \61131 , \61130 );
xor \U$60755 ( \61132 , \59690 , \59692 );
not \U$60756 ( \61133 , \61132 );
and \U$60757 ( \61134 , \61131 , \61133 );
and \U$60758 ( \61135 , \61130 , \61132 );
nor \U$60759 ( \61136 , \61134 , \61135 );
xnor \U$60760 ( \61137 , \61123 , \61136 );
or \U$60761 ( \61138 , \61119 , \61137 );
or \U$60762 ( \61139 , \61123 , \61136 );
nand \U$60763 ( \61140 , \61138 , \61139 );
xor \U$60764 ( \61141 , \59581 , \59687 );
xor \U$60765 ( \61142 , \61141 , \59693 );
not \U$60766 ( \61143 , \61132 );
not \U$60767 ( \61144 , \61129 );
or \U$60768 ( \61145 , \61143 , \61144 );
or \U$60769 ( \61146 , \61129 , \61132 );
nand \U$60770 ( \61147 , \61146 , \61125 );
nand \U$60771 ( \61148 , \61145 , \61147 );
xor \U$60772 ( \61149 , \61142 , \61148 );
and \U$60773 ( \61150 , \61140 , \61149 );
and \U$60774 ( \61151 , \61142 , \61148 );
nor \U$60775 ( \61152 , \61150 , \61151 );
or \U$60776 ( \61153 , \59698 , \61152 );
nand \U$60777 ( \61154 , \59697 , \61153 );
and \U$60778 ( \61155 , \59571 , \61154 );
nor \U$60779 ( \61156 , \59570 , \61155 );
or \U$60780 ( \61157 , \59446 , \61156 );
nand \U$60781 ( \61158 , \59445 , \61157 );
or \U$60782 ( \61159 , \59270 , \59280 );
not \U$60783 ( \61160 , \59280 );
not \U$60784 ( \61161 , \59270 );
or \U$60785 ( \61162 , \61160 , \61161 );
nand \U$60786 ( \61163 , \61162 , \59259 );
nand \U$60787 ( \61164 , \61159 , \61163 );
not \U$60788 ( \61165 , \59113 );
not \U$60789 ( \61166 , \59124 );
or \U$60790 ( \61167 , \61165 , \61166 );
or \U$60791 ( \61168 , \59124 , \59113 );
nand \U$60792 ( \61169 , \61167 , \61168 );
xor \U$60793 ( \61170 , \61164 , \61169 );
and \U$60794 ( \61171 , \61158 , \61170 );
and \U$60795 ( \61172 , \61164 , \61169 );
nor \U$60796 ( \61173 , \61171 , \61172 );
or \U$60797 ( \61174 , \59127 , \61173 );
nand \U$60798 ( \61175 , \59126 , \61174 );
not \U$60799 ( \61176 , \58928 );
nor \U$60800 ( \61177 , \61176 , \59103 );
xor \U$60801 ( \61178 , \58451 , \58671 );
xor \U$60802 ( \61179 , \61178 , \58839 );
xor \U$60803 ( \61180 , \61177 , \61179 );
and \U$60804 ( \61181 , \61175 , \61180 );
and \U$60805 ( \61182 , \61177 , \61179 );
nor \U$60806 ( \61183 , \61181 , \61182 );
or \U$60807 ( \61184 , \58924 , \61183 );
nand \U$60808 ( \61185 , \58923 , \61184 );
not \U$60809 ( \61186 , \58843 );
not \U$60810 ( \61187 , \58918 );
or \U$60811 ( \61188 , \61186 , \61187 );
or \U$60812 ( \61189 , \58918 , \58843 );
nand \U$60813 ( \61190 , \61189 , \58847 );
nand \U$60814 ( \61191 , \61188 , \61190 );
xor \U$60815 ( \61192 , \57933 , \58005 );
xor \U$60816 ( \61193 , \61192 , \58026 );
not \U$60817 ( \61194 , \61193 );
xor \U$60818 ( \61195 , \58857 , \58861 );
and \U$60819 ( \61196 , \61195 , \58866 );
and \U$60820 ( \61197 , \58857 , \58861 );
nor \U$60821 ( \61198 , \61196 , \61197 );
not \U$60822 ( \61199 , \61198 );
xor \U$60823 ( \61200 , \58870 , \58880 );
and \U$60824 ( \61201 , \61200 , \58891 );
and \U$60825 ( \61202 , \58870 , \58880 );
nor \U$60826 ( \61203 , \61201 , \61202 );
not \U$60827 ( \61204 , \61203 );
or \U$60828 ( \61205 , \61199 , \61204 );
or \U$60829 ( \61206 , \61203 , \61198 );
nand \U$60830 ( \61207 , \61205 , \61206 );
not \U$60831 ( \61208 , \61207 );
xor \U$60832 ( \61209 , \57651 , \57676 );
xor \U$60833 ( \61210 , \61209 , \57702 );
not \U$60834 ( \61211 , \61210 );
and \U$60835 ( \61212 , \61208 , \61211 );
and \U$60836 ( \61213 , \61207 , \61210 );
nor \U$60837 ( \61214 , \61212 , \61213 );
not \U$60838 ( \61215 , \61214 );
or \U$60839 ( \61216 , \61194 , \61215 );
or \U$60840 ( \61217 , \61214 , \61193 );
nand \U$60841 ( \61218 , \61216 , \61217 );
xor \U$60842 ( \61219 , \58896 , \58900 );
and \U$60843 ( \61220 , \61219 , \58917 );
and \U$60844 ( \61221 , \58896 , \58900 );
or \U$60845 ( \61222 , \61220 , \61221 );
xor \U$60846 ( \61223 , \61218 , \61222 );
xor \U$60847 ( \61224 , \57796 , \57798 );
xor \U$60848 ( \61225 , \61224 , \57801 );
xor \U$60849 ( \61226 , \57855 , \57862 );
xor \U$60850 ( \61227 , \61225 , \61226 );
not \U$60851 ( \61228 , \61227 );
xor \U$60852 ( \61229 , \58905 , \58907 );
and \U$60853 ( \61230 , \61229 , \58916 );
and \U$60854 ( \61231 , \58905 , \58907 );
or \U$60855 ( \61232 , \61230 , \61231 );
not \U$60856 ( \61233 , \61232 );
not \U$60857 ( \61234 , \58892 );
nand \U$60858 ( \61235 , \61234 , \58867 );
not \U$60859 ( \61236 , \61235 );
and \U$60860 ( \61237 , \61233 , \61236 );
and \U$60861 ( \61238 , \61232 , \61235 );
nor \U$60862 ( \61239 , \61237 , \61238 );
not \U$60863 ( \61240 , \61239 );
or \U$60864 ( \61241 , \61228 , \61240 );
or \U$60865 ( \61242 , \61239 , \61227 );
nand \U$60866 ( \61243 , \61241 , \61242 );
xor \U$60867 ( \61244 , \61223 , \61243 );
xor \U$60868 ( \61245 , \61191 , \61244 );
and \U$60869 ( \61246 , \61185 , \61245 );
and \U$60870 ( \61247 , \61191 , \61244 );
nor \U$60871 ( \61248 , \61246 , \61247 );
or \U$60872 ( \61249 , \61198 , \61210 );
not \U$60873 ( \61250 , \61210 );
not \U$60874 ( \61251 , \61198 );
or \U$60875 ( \61252 , \61250 , \61251 );
nand \U$60876 ( \61253 , \61252 , \61203 );
nand \U$60877 ( \61254 , \61249 , \61253 );
xor \U$60878 ( \61255 , \58039 , \58043 );
xor \U$60879 ( \61256 , \61254 , \61255 );
xor \U$60880 ( \61257 , \57867 , \58029 );
xor \U$60881 ( \61258 , \61257 , \58034 );
xor \U$60882 ( \61259 , \61256 , \61258 );
not \U$60883 ( \61260 , \61259 );
not \U$60884 ( \61261 , \61214 );
nand \U$60885 ( \61262 , \61261 , \61193 );
not \U$60886 ( \61263 , \61235 );
and \U$60887 ( \61264 , \61263 , \61227 );
not \U$60888 ( \61265 , \61227 );
nand \U$60889 ( \61266 , \61265 , \61235 );
and \U$60890 ( \61267 , \61232 , \61266 );
nor \U$60891 ( \61268 , \61264 , \61267 );
xnor \U$60892 ( \61269 , \61262 , \61268 );
not \U$60893 ( \61270 , \61269 );
and \U$60894 ( \61271 , \61260 , \61270 );
and \U$60895 ( \61272 , \61269 , \61259 );
nor \U$60896 ( \61273 , \61271 , \61272 );
xor \U$60897 ( \61274 , \61218 , \61222 );
and \U$60898 ( \61275 , \61274 , \61243 );
and \U$60899 ( \61276 , \61218 , \61222 );
nor \U$60900 ( \61277 , \61275 , \61276 );
xnor \U$60901 ( \61278 , \61273 , \61277 );
or \U$60902 ( \61279 , \61248 , \61278 );
or \U$60903 ( \61280 , \61277 , \61273 );
nand \U$60904 ( \61281 , \61279 , \61280 );
or \U$60905 ( \61282 , \61268 , \61262 );
not \U$60906 ( \61283 , \61262 );
not \U$60907 ( \61284 , \61268 );
or \U$60908 ( \61285 , \61283 , \61284 );
nand \U$60909 ( \61286 , \61285 , \61259 );
nand \U$60910 ( \61287 , \61282 , \61286 );
xor \U$60911 ( \61288 , \58037 , \58044 );
xor \U$60912 ( \61289 , \61288 , \58047 );
xor \U$60913 ( \61290 , \57789 , \57809 );
xor \U$60914 ( \61291 , \61290 , \57824 );
xor \U$60915 ( \61292 , \61289 , \61291 );
xor \U$60916 ( \61293 , \61254 , \61255 );
and \U$60917 ( \61294 , \61293 , \61258 );
and \U$60918 ( \61295 , \61254 , \61255 );
or \U$60919 ( \61296 , \61294 , \61295 );
xor \U$60920 ( \61297 , \61292 , \61296 );
xor \U$60921 ( \61298 , \61287 , \61297 );
and \U$60922 ( \61299 , \61281 , \61298 );
and \U$60923 ( \61300 , \61287 , \61297 );
nor \U$60924 ( \61301 , \61299 , \61300 );
xor \U$60925 ( \61302 , \61289 , \61291 );
and \U$60926 ( \61303 , \61302 , \61296 );
and \U$60927 ( \61304 , \61289 , \61291 );
nor \U$60928 ( \61305 , \61303 , \61304 );
not \U$60929 ( \61306 , \57849 );
not \U$60930 ( \61307 , \58050 );
or \U$60931 ( \61308 , \61306 , \61307 );
or \U$60932 ( \61309 , \58050 , \57849 );
nand \U$60933 ( \61310 , \61308 , \61309 );
not \U$60934 ( \61311 , \61310 );
not \U$60935 ( \61312 , \57839 );
and \U$60936 ( \61313 , \61311 , \61312 );
and \U$60937 ( \61314 , \61310 , \57839 );
nor \U$60938 ( \61315 , \61313 , \61314 );
xnor \U$60939 ( \61316 , \61305 , \61315 );
or \U$60940 ( \61317 , \61301 , \61316 );
or \U$60941 ( \61318 , \61305 , \61315 );
nand \U$60942 ( \61319 , \61317 , \61318 );
and \U$60943 ( \61320 , \58054 , \61319 );
nor \U$60944 ( \61321 , \58053 , \61320 );
not \U$60945 ( \61322 , \57387 );
not \U$60946 ( \61323 , \57596 );
or \U$60947 ( \61324 , \61322 , \61323 );
or \U$60948 ( \61325 , \57596 , \57387 );
nand \U$60949 ( \61326 , \61324 , \61325 );
not \U$60950 ( \61327 , \61326 );
not \U$60951 ( \61328 , \57381 );
and \U$60952 ( \61329 , \61327 , \61328 );
and \U$60953 ( \61330 , \61326 , \57381 );
nor \U$60954 ( \61331 , \61329 , \61330 );
xor \U$60955 ( \61332 , \57605 , \57829 );
and \U$60956 ( \61333 , \61332 , \57832 );
and \U$60957 ( \61334 , \57605 , \57829 );
nor \U$60958 ( \61335 , \61333 , \61334 );
xnor \U$60959 ( \61336 , \61331 , \61335 );
or \U$60960 ( \61337 , \61321 , \61336 );
or \U$60961 ( \61338 , \61331 , \61335 );
nand \U$60962 ( \61339 , \61337 , \61338 );
and \U$60963 ( \61340 , \57600 , \61339 );
nor \U$60964 ( \61341 , \57599 , \61340 );
or \U$60965 ( \61342 , \57369 , \61341 );
nand \U$60966 ( \61343 , \57368 , \61342 );
and \U$60967 ( \61344 , \57158 , \61343 );
nor \U$60968 ( \61345 , \57157 , \61344 );
or \U$60969 ( \61346 , \56881 , \61345 );
nand \U$60970 ( \61347 , \56880 , \61346 );
not \U$60971 ( \61348 , \56604 );
nor \U$60972 ( \61349 , \61348 , \56869 );
xor \U$60973 ( \61350 , \56598 , \56600 );
and \U$60974 ( \61351 , \61350 , \56603 );
and \U$60975 ( \61352 , \56598 , \56600 );
or \U$60976 ( \61353 , \61351 , \61352 );
not \U$60977 ( \61354 , \61353 );
xnor \U$60978 ( \61355 , \56025 , \56312 );
not \U$60979 ( \61356 , \61355 );
not \U$60980 ( \61357 , \56030 );
and \U$60981 ( \61358 , \61356 , \61357 );
and \U$60982 ( \61359 , \61355 , \56030 );
nor \U$60983 ( \61360 , \61358 , \61359 );
not \U$60984 ( \61361 , \61360 );
or \U$60985 ( \61362 , \61354 , \61361 );
or \U$60986 ( \61363 , \61360 , \61353 );
nand \U$60987 ( \61364 , \61362 , \61363 );
xor \U$60988 ( \61365 , \61349 , \61364 );
and \U$60989 ( \61366 , \61347 , \61365 );
and \U$60990 ( \61367 , \61349 , \61364 );
nor \U$60991 ( \61368 , \61366 , \61367 );
not \U$60992 ( \61369 , \61360 );
nand \U$60993 ( \61370 , \61369 , \61353 );
xnor \U$60994 ( \61371 , \56314 , \56020 );
not \U$60995 ( \61372 , \61371 );
not \U$60996 ( \61373 , \55748 );
and \U$60997 ( \61374 , \61372 , \61373 );
and \U$60998 ( \61375 , \61371 , \55748 );
nor \U$60999 ( \61376 , \61374 , \61375 );
xnor \U$61000 ( \61377 , \61370 , \61376 );
or \U$61001 ( \61378 , \61368 , \61377 );
or \U$61002 ( \61379 , \61370 , \61376 );
nand \U$61003 ( \61380 , \61378 , \61379 );
and \U$61004 ( \61381 , \56340 , \61380 );
nor \U$61005 ( \61382 , \56339 , \61381 );
not \U$61006 ( \61383 , \56334 );
nand \U$61007 ( \61384 , \61383 , \56320 );
xor \U$61008 ( \61385 , \54826 , \54832 );
xor \U$61009 ( \61386 , \61385 , \54847 );
not \U$61010 ( \61387 , \56330 );
not \U$61011 ( \61388 , \56327 );
or \U$61012 ( \61389 , \61387 , \61388 );
or \U$61013 ( \61390 , \56327 , \56330 );
nand \U$61014 ( \61391 , \61390 , \56325 );
nand \U$61015 ( \61392 , \61389 , \61391 );
xnor \U$61016 ( \61393 , \61386 , \61392 );
not \U$61017 ( \61394 , \61393 );
xor \U$61018 ( \61395 , \55116 , \55123 );
xor \U$61019 ( \61396 , \61395 , \55128 );
not \U$61020 ( \61397 , \61396 );
and \U$61021 ( \61398 , \61394 , \61397 );
and \U$61022 ( \61399 , \61393 , \61396 );
nor \U$61023 ( \61400 , \61398 , \61399 );
xnor \U$61024 ( \61401 , \61384 , \61400 );
or \U$61025 ( \61402 , \61382 , \61401 );
or \U$61026 ( \61403 , \61384 , \61400 );
nand \U$61027 ( \61404 , \61402 , \61403 );
not \U$61028 ( \61405 , \61386 );
not \U$61029 ( \61406 , \61396 );
or \U$61030 ( \61407 , \61405 , \61406 );
or \U$61031 ( \61408 , \61396 , \61386 );
nand \U$61032 ( \61409 , \61408 , \61392 );
nand \U$61033 ( \61410 , \61407 , \61409 );
xor \U$61034 ( \61411 , \54362 , \54851 );
xor \U$61035 ( \61412 , \61411 , \55131 );
xor \U$61036 ( \61413 , \61410 , \61412 );
and \U$61037 ( \61414 , \61404 , \61413 );
and \U$61038 ( \61415 , \61410 , \61412 );
nor \U$61039 ( \61416 , \61414 , \61415 );
or \U$61040 ( \61417 , \55510 , \61416 );
nand \U$61041 ( \61418 , \55509 , \61417 );
or \U$61042 ( \61419 , \55504 , \55136 );
not \U$61043 ( \61420 , \55136 );
not \U$61044 ( \61421 , \55504 );
or \U$61045 ( \61422 , \61420 , \61421 );
nand \U$61046 ( \61423 , \61422 , \55141 );
nand \U$61047 ( \61424 , \61419 , \61423 );
not \U$61048 ( \61425 , \55286 );
not \U$61049 ( \61426 , \55276 );
and \U$61050 ( \61427 , \61425 , \61426 );
and \U$61051 ( \61428 , \55286 , \55276 );
nor \U$61052 ( \61429 , \61428 , \55295 );
nor \U$61053 ( \61430 , \61427 , \61429 );
xor \U$61054 ( \61431 , \55158 , \55162 );
and \U$61055 ( \61432 , \61431 , \55171 );
and \U$61056 ( \61433 , \55158 , \55162 );
nor \U$61057 ( \61434 , \61432 , \61433 );
xor \U$61058 ( \61435 , \61430 , \61434 );
not \U$61059 ( \61436 , \55387 );
not \U$61060 ( \61437 , \55419 );
and \U$61061 ( \61438 , \61436 , \61437 );
and \U$61062 ( \61439 , \55387 , \55419 );
nor \U$61063 ( \61440 , \61439 , \55492 );
nor \U$61064 ( \61441 , \61438 , \61440 );
xor \U$61065 ( \61442 , \61435 , \61441 );
not \U$61066 ( \61443 , \61442 );
xor \U$61067 ( \61444 , \55215 , \55229 );
xor \U$61068 ( \61445 , \61444 , \55244 );
and \U$61069 ( \61446 , \55300 , \61445 );
xor \U$61070 ( \61447 , \55215 , \55229 );
xor \U$61071 ( \61448 , \61447 , \55244 );
and \U$61072 ( \61449 , \55497 , \61448 );
and \U$61073 ( \61450 , \55300 , \55497 );
or \U$61074 ( \61451 , \61446 , \61449 , \61450 );
xor \U$61075 ( \61452 , \55188 , \55192 );
and \U$61076 ( \61453 , \61452 , \55197 );
and \U$61077 ( \61454 , \55188 , \55192 );
or \U$61078 ( \61455 , \61453 , \61454 );
xor \U$61079 ( \61456 , \61451 , \61455 );
or \U$61080 ( \61457 , \55488 , \55426 );
not \U$61081 ( \61458 , \55426 );
not \U$61082 ( \61459 , \55488 );
or \U$61083 ( \61460 , \61458 , \61459 );
nand \U$61084 ( \61461 , \61460 , \55450 );
nand \U$61085 ( \61462 , \61457 , \61461 );
and \U$61086 ( \61463 , \15726 , RIae751a0_2);
and \U$61087 ( \61464 , RIae75380_6, RIae7aab0_192);
nor \U$61088 ( \61465 , \61463 , \61464 );
and \U$61089 ( \61466 , \61465 , \14959 );
not \U$61090 ( \61467 , \61465 );
and \U$61091 ( \61468 , \61467 , RIae7aa38_191);
nor \U$61092 ( \61469 , \61466 , \61468 );
xor \U$61093 ( \61470 , \61469 , \1488 );
and \U$61094 ( \61471 , \14964 , RIae75740_14);
and \U$61095 ( \61472 , RIae75290_4, \14962 );
nor \U$61096 ( \61473 , \61471 , \61472 );
and \U$61097 ( \61474 , \61473 , \14463 );
not \U$61098 ( \61475 , \61473 );
and \U$61099 ( \61476 , \61475 , \14462 );
nor \U$61100 ( \61477 , \61474 , \61476 );
xor \U$61101 ( \61478 , \61470 , \61477 );
xor \U$61102 ( \61479 , \61462 , \61478 );
or \U$61103 ( \61480 , \55331 , \55383 );
not \U$61104 ( \61481 , \55383 );
not \U$61105 ( \61482 , \55331 );
or \U$61106 ( \61483 , \61481 , \61482 );
nand \U$61107 ( \61484 , \61483 , \55355 );
nand \U$61108 ( \61485 , \61480 , \61484 );
xor \U$61109 ( \61486 , \61479 , \61485 );
xor \U$61110 ( \61487 , \55219 , \55223 );
and \U$61111 ( \61488 , \61487 , \55228 );
and \U$61112 ( \61489 , \55219 , \55223 );
or \U$61113 ( \61490 , \61488 , \61489 );
xor \U$61114 ( \61491 , \55202 , \55209 );
and \U$61115 ( \61492 , \61491 , \55214 );
and \U$61116 ( \61493 , \55202 , \55209 );
or \U$61117 ( \61494 , \61492 , \61493 );
xor \U$61118 ( \61495 , \61490 , \61494 );
xor \U$61119 ( \61496 , \55234 , \55238 );
and \U$61120 ( \61497 , \61496 , \55243 );
and \U$61121 ( \61498 , \55234 , \55238 );
or \U$61122 ( \61499 , \61497 , \61498 );
xor \U$61123 ( \61500 , \61495 , \61499 );
and \U$61124 ( \61501 , \13059 , RIae75dd0_28);
and \U$61125 ( \61502 , RIae75650_12, \13057 );
nor \U$61126 ( \61503 , \61501 , \61502 );
and \U$61127 ( \61504 , \61503 , \13063 );
not \U$61128 ( \61505 , \61503 );
and \U$61129 ( \61506 , \61505 , \12718 );
nor \U$61130 ( \61507 , \61504 , \61506 );
and \U$61131 ( \61508 , \12180 , RIae75ec0_30);
and \U$61132 ( \61509 , RIae75ce0_26, \12178 );
nor \U$61133 ( \61510 , \61508 , \61509 );
and \U$61134 ( \61511 , \61510 , \12184 );
not \U$61135 ( \61512 , \61510 );
and \U$61136 ( \61513 , \61512 , \11827 );
nor \U$61137 ( \61514 , \61511 , \61513 );
xor \U$61138 ( \61515 , \61507 , \61514 );
and \U$61139 ( \61516 , \14059 , RIae75560_10);
and \U$61140 ( \61517 , RIae75830_16, \14057 );
nor \U$61141 ( \61518 , \61516 , \61517 );
and \U$61142 ( \61519 , \61518 , \13502 );
not \U$61143 ( \61520 , \61518 );
and \U$61144 ( \61521 , \61520 , \14063 );
nor \U$61145 ( \61522 , \61519 , \61521 );
xor \U$61146 ( \61523 , \61515 , \61522 );
and \U$61147 ( \61524 , \8966 , RIae788f0_120);
and \U$61148 ( \61525 , RIae78800_118, \8964 );
nor \U$61149 ( \61526 , \61524 , \61525 );
and \U$61150 ( \61527 , \61526 , \8799 );
not \U$61151 ( \61528 , \61526 );
and \U$61152 ( \61529 , \61528 , \8789 );
nor \U$61153 ( \61530 , \61527 , \61529 );
and \U$61154 ( \61531 , \7633 , RIae77bd0_92);
and \U$61155 ( \61532 , RIae77db0_96, \7631 );
nor \U$61156 ( \61533 , \61531 , \61532 );
and \U$61157 ( \61534 , \61533 , \7206 );
not \U$61158 ( \61535 , \61533 );
and \U$61159 ( \61536 , \61535 , \7205 );
nor \U$61160 ( \61537 , \61534 , \61536 );
xor \U$61161 ( \61538 , \61530 , \61537 );
and \U$61162 ( \61539 , \8371 , RIae77ea0_98);
and \U$61163 ( \61540 , RIae789e0_122, \8369 );
nor \U$61164 ( \61541 , \61539 , \61540 );
and \U$61165 ( \61542 , \61541 , \8020 );
not \U$61166 ( \61543 , \61541 );
and \U$61167 ( \61544 , \61543 , \8019 );
nor \U$61168 ( \61545 , \61542 , \61544 );
xor \U$61169 ( \61546 , \61538 , \61545 );
and \U$61170 ( \61547 , \9760 , RIae78710_116);
and \U$61171 ( \61548 , RIae75bf0_24, \9758 );
nor \U$61172 ( \61549 , \61547 , \61548 );
and \U$61173 ( \61550 , \61549 , \9273 );
not \U$61174 ( \61551 , \61549 );
and \U$61175 ( \61552 , \61551 , \9764 );
nor \U$61176 ( \61553 , \61550 , \61552 );
and \U$61177 ( \61554 , \10548 , RIae75b00_22);
and \U$61178 ( \61555 , RIae75a10_20, \10546 );
nor \U$61179 ( \61556 , \61554 , \61555 );
and \U$61180 ( \61557 , \61556 , \10421 );
not \U$61181 ( \61558 , \61556 );
and \U$61182 ( \61559 , \61558 , \10118 );
nor \U$61183 ( \61560 , \61557 , \61559 );
xor \U$61184 ( \61561 , \61553 , \61560 );
and \U$61185 ( \61562 , \11470 , RIae75920_18);
and \U$61186 ( \61563 , RIae75fb0_32, \11468 );
nor \U$61187 ( \61564 , \61562 , \61563 );
and \U$61188 ( \61565 , \61564 , \10936 );
not \U$61189 ( \61566 , \61564 );
and \U$61190 ( \61567 , \61566 , \11474 );
nor \U$61191 ( \61568 , \61565 , \61567 );
xor \U$61192 ( \61569 , \61561 , \61568 );
xor \U$61193 ( \61570 , \61546 , \61569 );
xor \U$61194 ( \61571 , \61523 , \61570 );
or \U$61195 ( \61572 , \55484 , \55463 );
not \U$61196 ( \61573 , \55463 );
not \U$61197 ( \61574 , \55484 );
or \U$61198 ( \61575 , \61573 , \61574 );
nand \U$61199 ( \61576 , \61575 , \55472 );
nand \U$61200 ( \61577 , \61572 , \61576 );
nand \U$61201 ( \61578 , RIae77630_80, \1591 );
and \U$61202 ( \61579 , \61578 , \1498 );
not \U$61203 ( \61580 , \61578 );
and \U$61204 ( \61581 , \61580 , \1488 );
nor \U$61205 ( \61582 , \61579 , \61581 );
xor \U$61206 ( \61583 , \61577 , \61582 );
and \U$61207 ( \61584 , \1939 , RIae77540_78);
and \U$61208 ( \61585 , RIae776a8_81, \1937 );
nor \U$61209 ( \61586 , \61584 , \61585 );
and \U$61210 ( \61587 , \61586 , \1734 );
not \U$61211 ( \61588 , \61586 );
and \U$61212 ( \61589 , \61588 , \1735 );
nor \U$61213 ( \61590 , \61587 , \61589 );
not \U$61214 ( \61591 , \61590 );
and \U$61215 ( \61592 , \2224 , RIae77450_76);
and \U$61216 ( \61593 , RIae77ae0_90, \2222 );
nor \U$61217 ( \61594 , \61592 , \61593 );
and \U$61218 ( \61595 , \61594 , \2060 );
not \U$61219 ( \61596 , \61594 );
and \U$61220 ( \61597 , \61596 , \2061 );
nor \U$61221 ( \61598 , \61595 , \61597 );
and \U$61222 ( \61599 , \2607 , RIae779f0_88);
and \U$61223 ( \61600 , RIae77810_84, \2605 );
nor \U$61224 ( \61601 , \61599 , \61600 );
and \U$61225 ( \61602 , \61601 , \2397 );
not \U$61226 ( \61603 , \61601 );
and \U$61227 ( \61604 , \61603 , \2611 );
nor \U$61228 ( \61605 , \61602 , \61604 );
xor \U$61229 ( \61606 , \61598 , \61605 );
not \U$61230 ( \61607 , \61606 );
or \U$61231 ( \61608 , \61591 , \61607 );
or \U$61232 ( \61609 , \61606 , \61590 );
nand \U$61233 ( \61610 , \61608 , \61609 );
xor \U$61234 ( \61611 , \61583 , \61610 );
xor \U$61235 ( \61612 , \61571 , \61611 );
and \U$61236 ( \61613 , \2783 , RIae77900_86);
and \U$61237 ( \61614 , RIae76fa0_66, \2781 );
nor \U$61238 ( \61615 , \61613 , \61614 );
not \U$61239 ( \61616 , \61615 );
not \U$61240 ( \61617 , \3089 );
and \U$61241 ( \61618 , \61616 , \61617 );
and \U$61242 ( \61619 , \61615 , \3089 );
nor \U$61243 ( \61620 , \61618 , \61619 );
not \U$61244 ( \61621 , \61620 );
and \U$61245 ( \61622 , \3214 , RIae76eb0_64);
and \U$61246 ( \61623 , RIae76dc0_62, \3212 );
nor \U$61247 ( \61624 , \61622 , \61623 );
not \U$61248 ( \61625 , \61624 );
not \U$61249 ( \61626 , \2774 );
and \U$61250 ( \61627 , \61625 , \61626 );
and \U$61251 ( \61628 , \61624 , \3218 );
nor \U$61252 ( \61629 , \61627 , \61628 );
and \U$61253 ( \61630 , \3730 , RIae76cd0_60);
and \U$61254 ( \61631 , RIae77108_69, \3728 );
nor \U$61255 ( \61632 , \61630 , \61631 );
and \U$61256 ( \61633 , \61632 , \3422 );
not \U$61257 ( \61634 , \61632 );
and \U$61258 ( \61635 , \61634 , \3732 );
nor \U$61259 ( \61636 , \61633 , \61635 );
xor \U$61260 ( \61637 , \61629 , \61636 );
not \U$61261 ( \61638 , \61637 );
or \U$61262 ( \61639 , \61621 , \61638 );
or \U$61263 ( \61640 , \61637 , \61620 );
nand \U$61264 ( \61641 , \61639 , \61640 );
and \U$61265 ( \61642 , \5896 , RIae78080_102);
and \U$61266 ( \61643 , RIae78260_106, \5894 );
nor \U$61267 ( \61644 , \61642 , \61643 );
and \U$61268 ( \61645 , \61644 , \5590 );
not \U$61269 ( \61646 , \61644 );
and \U$61270 ( \61647 , \61646 , \5589 );
nor \U$61271 ( \61648 , \61645 , \61647 );
and \U$61272 ( \61649 , \6172 , RIae78620_114);
and \U$61273 ( \61650 , RIae78440_110, \6170 );
nor \U$61274 ( \61651 , \61649 , \61650 );
and \U$61275 ( \61652 , \61651 , \6176 );
not \U$61276 ( \61653 , \61651 );
and \U$61277 ( \61654 , \61653 , \6175 );
nor \U$61278 ( \61655 , \61652 , \61654 );
xor \U$61279 ( \61656 , \61648 , \61655 );
and \U$61280 ( \61657 , \6941 , RIae784b8_111);
and \U$61281 ( \61658 , RIae77cc0_94, \6939 );
nor \U$61282 ( \61659 , \61657 , \61658 );
and \U$61283 ( \61660 , \61659 , \6314 );
not \U$61284 ( \61661 , \61659 );
and \U$61285 ( \61662 , \61661 , \6945 );
nor \U$61286 ( \61663 , \61660 , \61662 );
xor \U$61287 ( \61664 , \61656 , \61663 );
xor \U$61288 ( \61665 , \61641 , \61664 );
and \U$61289 ( \61666 , \5399 , RIae78170_104);
and \U$61290 ( \61667 , RIae77f90_100, \5397 );
nor \U$61291 ( \61668 , \61666 , \61667 );
and \U$61292 ( \61669 , \61668 , \5016 );
not \U$61293 ( \61670 , \61668 );
and \U$61294 ( \61671 , \61670 , \5403 );
nor \U$61295 ( \61672 , \61669 , \61671 );
and \U$61296 ( \61673 , \4247 , RIae77090_68);
and \U$61297 ( \61674 , RIae77270_72, \4245 );
nor \U$61298 ( \61675 , \61673 , \61674 );
and \U$61299 ( \61676 , \61675 , \3989 );
not \U$61300 ( \61677 , \61675 );
and \U$61301 ( \61678 , \61677 , \4251 );
nor \U$61302 ( \61679 , \61676 , \61678 );
xor \U$61303 ( \61680 , \61672 , \61679 );
and \U$61304 ( \61681 , \4688 , RIae77360_74);
and \U$61305 ( \61682 , RIae78350_108, \4686 );
nor \U$61306 ( \61683 , \61681 , \61682 );
and \U$61307 ( \61684 , \61683 , \4481 );
not \U$61308 ( \61685 , \61683 );
and \U$61309 ( \61686 , \61685 , \4482 );
nor \U$61310 ( \61687 , \61684 , \61686 );
xor \U$61311 ( \61688 , \61680 , \61687 );
xor \U$61312 ( \61689 , \61665 , \61688 );
xor \U$61313 ( \61690 , \61612 , \61689 );
xor \U$61314 ( \61691 , \61500 , \61690 );
xor \U$61315 ( \61692 , \61486 , \61691 );
xor \U$61316 ( \61693 , \61456 , \61692 );
not \U$61317 ( \61694 , \61693 );
or \U$61318 ( \61695 , \61443 , \61694 );
or \U$61319 ( \61696 , \61693 , \61442 );
nand \U$61320 ( \61697 , \61695 , \61696 );
not \U$61321 ( \61698 , \55500 );
not \U$61322 ( \61699 , \55182 );
or \U$61323 ( \61700 , \61698 , \61699 );
or \U$61324 ( \61701 , \55182 , \55500 );
nand \U$61325 ( \61702 , \61701 , \55150 );
nand \U$61326 ( \61703 , \61700 , \61702 );
xor \U$61327 ( \61704 , \61697 , \61703 );
and \U$61328 ( \61705 , \55198 , \55499 );
or \U$61329 ( \61706 , \55327 , \55307 );
not \U$61330 ( \61707 , \55307 );
not \U$61331 ( \61708 , \55327 );
or \U$61332 ( \61709 , \61707 , \61708 );
nand \U$61333 ( \61710 , \61709 , \55315 );
nand \U$61334 ( \61711 , \61706 , \61710 );
xor \U$61335 ( \61712 , \55434 , \55441 );
and \U$61336 ( \61713 , \61712 , \55449 );
and \U$61337 ( \61714 , \55434 , \55441 );
or \U$61338 ( \61715 , \61713 , \61714 );
xor \U$61339 ( \61716 , \61711 , \61715 );
xor \U$61340 ( \61717 , \55339 , \55346 );
and \U$61341 ( \61718 , \61717 , \55354 );
and \U$61342 ( \61719 , \55339 , \55346 );
or \U$61343 ( \61720 , \61718 , \61719 );
xor \U$61344 ( \61721 , \61716 , \61720 );
xor \U$61345 ( \61722 , \55367 , \55374 );
and \U$61346 ( \61723 , \61722 , \55382 );
and \U$61347 ( \61724 , \55367 , \55374 );
nor \U$61348 ( \61725 , \61723 , \61724 );
or \U$61349 ( \61726 , \55415 , \55395 );
not \U$61350 ( \61727 , \55395 );
not \U$61351 ( \61728 , \55415 );
or \U$61352 ( \61729 , \61727 , \61728 );
nand \U$61353 ( \61730 , \61729 , \55403 );
nand \U$61354 ( \61731 , \61726 , \61730 );
xor \U$61355 ( \61732 , \61725 , \61731 );
or \U$61356 ( \61733 , \55272 , \55252 );
not \U$61357 ( \61734 , \55252 );
not \U$61358 ( \61735 , \55272 );
or \U$61359 ( \61736 , \61734 , \61735 );
nand \U$61360 ( \61737 , \61736 , \55260 );
nand \U$61361 ( \61738 , \61733 , \61737 );
xor \U$61362 ( \61739 , \61732 , \61738 );
xor \U$61363 ( \61740 , \55215 , \55229 );
and \U$61364 ( \61741 , \61740 , \55244 );
and \U$61365 ( \61742 , \55215 , \55229 );
or \U$61366 ( \61743 , \61741 , \61742 );
xor \U$61367 ( \61744 , \61739 , \61743 );
xor \U$61368 ( \61745 , \61721 , \61744 );
xor \U$61369 ( \61746 , \61705 , \61745 );
xor \U$61370 ( \61747 , \55154 , \55172 );
and \U$61371 ( \61748 , \61747 , \55181 );
and \U$61372 ( \61749 , \55154 , \55172 );
or \U$61373 ( \61750 , \61748 , \61749 );
xor \U$61374 ( \61751 , \61746 , \61750 );
xor \U$61375 ( \61752 , \61704 , \61751 );
xor \U$61376 ( \61753 , \61424 , \61752 );
and \U$61377 ( \61754 , \61418 , \61753 );
and \U$61378 ( \61755 , \61424 , \61752 );
nor \U$61379 ( \61756 , \61754 , \61755 );
not \U$61380 ( \61757 , \61442 );
nand \U$61381 ( \61758 , \61757 , \61693 );
not \U$61382 ( \61759 , \61758 );
xor \U$61383 ( \61760 , \61705 , \61745 );
and \U$61384 ( \61761 , \61760 , \61750 );
and \U$61385 ( \61762 , \61705 , \61745 );
or \U$61386 ( \61763 , \61761 , \61762 );
not \U$61387 ( \61764 , \61763 );
and \U$61388 ( \61765 , \61759 , \61764 );
and \U$61389 ( \61766 , \61758 , \61763 );
nor \U$61390 ( \61767 , \61765 , \61766 );
not \U$61391 ( \61768 , \61767 );
xor \U$61392 ( \61769 , \61451 , \61455 );
and \U$61393 ( \61770 , \61769 , \61692 );
and \U$61394 ( \61771 , \61451 , \61455 );
or \U$61395 ( \61772 , \61770 , \61771 );
xor \U$61396 ( \61773 , \61430 , \61434 );
and \U$61397 ( \61774 , \61773 , \61441 );
and \U$61398 ( \61775 , \61430 , \61434 );
nor \U$61399 ( \61776 , \61774 , \61775 );
xor \U$61400 ( \61777 , \61711 , \61715 );
xor \U$61401 ( \61778 , \61777 , \61720 );
and \U$61402 ( \61779 , \61739 , \61778 );
xor \U$61403 ( \61780 , \61711 , \61715 );
xor \U$61404 ( \61781 , \61780 , \61720 );
and \U$61405 ( \61782 , \61743 , \61781 );
and \U$61406 ( \61783 , \61739 , \61743 );
or \U$61407 ( \61784 , \61779 , \61782 , \61783 );
xor \U$61408 ( \61785 , \61776 , \61784 );
xor \U$61409 ( \61786 , \61462 , \61478 );
xor \U$61410 ( \61787 , \61786 , \61485 );
and \U$61411 ( \61788 , \61500 , \61787 );
xor \U$61412 ( \61789 , \61462 , \61478 );
xor \U$61413 ( \61790 , \61789 , \61485 );
and \U$61414 ( \61791 , \61690 , \61790 );
and \U$61415 ( \61792 , \61500 , \61690 );
or \U$61416 ( \61793 , \61788 , \61791 , \61792 );
xor \U$61417 ( \61794 , \61785 , \61793 );
xor \U$61418 ( \61795 , \61772 , \61794 );
xor \U$61419 ( \61796 , \61648 , \61655 );
and \U$61420 ( \61797 , \61796 , \61663 );
and \U$61421 ( \61798 , \61648 , \61655 );
or \U$61422 ( \61799 , \61797 , \61798 );
xor \U$61423 ( \61800 , \61672 , \61679 );
and \U$61424 ( \61801 , \61800 , \61687 );
and \U$61425 ( \61802 , \61672 , \61679 );
or \U$61426 ( \61803 , \61801 , \61802 );
xor \U$61427 ( \61804 , \61799 , \61803 );
xor \U$61428 ( \61805 , \61530 , \61537 );
and \U$61429 ( \61806 , \61805 , \61545 );
and \U$61430 ( \61807 , \61530 , \61537 );
or \U$61431 ( \61808 , \61806 , \61807 );
xor \U$61432 ( \61809 , \61804 , \61808 );
xor \U$61433 ( \61810 , \61553 , \61560 );
and \U$61434 ( \61811 , \61810 , \61568 );
and \U$61435 ( \61812 , \61553 , \61560 );
or \U$61436 ( \61813 , \61811 , \61812 );
xor \U$61437 ( \61814 , \61469 , \1488 );
and \U$61438 ( \61815 , \61814 , \61477 );
and \U$61439 ( \61816 , \61469 , \1488 );
or \U$61440 ( \61817 , \61815 , \61816 );
xor \U$61441 ( \61818 , \61813 , \61817 );
xor \U$61442 ( \61819 , \61507 , \61514 );
and \U$61443 ( \61820 , \61819 , \61522 );
and \U$61444 ( \61821 , \61507 , \61514 );
or \U$61445 ( \61822 , \61820 , \61821 );
xor \U$61446 ( \61823 , \61818 , \61822 );
xor \U$61447 ( \61824 , \61809 , \61823 );
not \U$61448 ( \61825 , \61620 );
not \U$61449 ( \61826 , \61629 );
and \U$61450 ( \61827 , \61825 , \61826 );
and \U$61451 ( \61828 , \61629 , \61620 );
nor \U$61452 ( \61829 , \61828 , \61636 );
nor \U$61453 ( \61830 , \61827 , \61829 );
not \U$61454 ( \61831 , \61590 );
not \U$61455 ( \61832 , \61605 );
and \U$61456 ( \61833 , \61831 , \61832 );
and \U$61457 ( \61834 , \61605 , \61590 );
nor \U$61458 ( \61835 , \61834 , \61598 );
nor \U$61459 ( \61836 , \61833 , \61835 );
xor \U$61460 ( \61837 , \61830 , \61836 );
and \U$61461 ( \61838 , \1939 , RIae776a8_81);
and \U$61462 ( \61839 , RIae77450_76, \1937 );
nor \U$61463 ( \61840 , \61838 , \61839 );
and \U$61464 ( \61841 , \61840 , \1734 );
not \U$61465 ( \61842 , \61840 );
and \U$61466 ( \61843 , \61842 , \1735 );
nor \U$61467 ( \61844 , \61841 , \61843 );
and \U$61468 ( \61845 , \1593 , RIae77630_80);
and \U$61469 ( \61846 , RIae77540_78, \1591 );
nor \U$61470 ( \61847 , \61845 , \61846 );
and \U$61471 ( \61848 , \61847 , \1488 );
not \U$61472 ( \61849 , \61847 );
and \U$61473 ( \61850 , \61849 , \1498 );
nor \U$61474 ( \61851 , \61848 , \61850 );
xor \U$61475 ( \61852 , \61844 , \61851 );
and \U$61476 ( \61853 , \2224 , RIae77ae0_90);
and \U$61477 ( \61854 , RIae779f0_88, \2222 );
nor \U$61478 ( \61855 , \61853 , \61854 );
and \U$61479 ( \61856 , \61855 , \2060 );
not \U$61480 ( \61857 , \61855 );
and \U$61481 ( \61858 , \61857 , \2061 );
nor \U$61482 ( \61859 , \61856 , \61858 );
xor \U$61483 ( \61860 , \61852 , \61859 );
xor \U$61484 ( \61861 , \61837 , \61860 );
not \U$61485 ( \61862 , \61861 );
and \U$61486 ( \61863 , \2783 , RIae76fa0_66);
and \U$61487 ( \61864 , RIae76eb0_64, \2781 );
nor \U$61488 ( \61865 , \61863 , \61864 );
not \U$61489 ( \61866 , \61865 );
not \U$61490 ( \61867 , \3089 );
and \U$61491 ( \61868 , \61866 , \61867 );
and \U$61492 ( \61869 , \61865 , \2789 );
nor \U$61493 ( \61870 , \61868 , \61869 );
and \U$61494 ( \61871 , \3214 , RIae76dc0_62);
and \U$61495 ( \61872 , RIae76cd0_60, \3212 );
nor \U$61496 ( \61873 , \61871 , \61872 );
not \U$61497 ( \61874 , \61873 );
not \U$61498 ( \61875 , \2774 );
and \U$61499 ( \61876 , \61874 , \61875 );
and \U$61500 ( \61877 , \61873 , \3218 );
nor \U$61501 ( \61878 , \61876 , \61877 );
xor \U$61502 ( \61879 , \61870 , \61878 );
and \U$61503 ( \61880 , \2607 , RIae77810_84);
and \U$61504 ( \61881 , RIae77900_86, \2605 );
nor \U$61505 ( \61882 , \61880 , \61881 );
and \U$61506 ( \61883 , \61882 , \2397 );
not \U$61507 ( \61884 , \61882 );
and \U$61508 ( \61885 , \61884 , \2611 );
nor \U$61509 ( \61886 , \61883 , \61885 );
xor \U$61510 ( \61887 , \61879 , \61886 );
not \U$61511 ( \61888 , \61887 );
and \U$61512 ( \61889 , \5399 , RIae77f90_100);
and \U$61513 ( \61890 , RIae78080_102, \5397 );
nor \U$61514 ( \61891 , \61889 , \61890 );
and \U$61515 ( \61892 , \61891 , \5403 );
not \U$61516 ( \61893 , \61891 );
and \U$61517 ( \61894 , \61893 , \5016 );
nor \U$61518 ( \61895 , \61892 , \61894 );
not \U$61519 ( \61896 , \61895 );
and \U$61520 ( \61897 , \5896 , RIae78260_106);
and \U$61521 ( \61898 , RIae78620_114, \5894 );
nor \U$61522 ( \61899 , \61897 , \61898 );
and \U$61523 ( \61900 , \61899 , \5589 );
not \U$61524 ( \61901 , \61899 );
and \U$61525 ( \61902 , \61901 , \5590 );
nor \U$61526 ( \61903 , \61900 , \61902 );
and \U$61527 ( \61904 , \6172 , RIae78440_110);
and \U$61528 ( \61905 , RIae784b8_111, \6170 );
nor \U$61529 ( \61906 , \61904 , \61905 );
and \U$61530 ( \61907 , \61906 , \6175 );
not \U$61531 ( \61908 , \61906 );
and \U$61532 ( \61909 , \61908 , \6176 );
nor \U$61533 ( \61910 , \61907 , \61909 );
xor \U$61534 ( \61911 , \61903 , \61910 );
not \U$61535 ( \61912 , \61911 );
or \U$61536 ( \61913 , \61896 , \61912 );
or \U$61537 ( \61914 , \61911 , \61895 );
nand \U$61538 ( \61915 , \61913 , \61914 );
not \U$61539 ( \61916 , \61915 );
or \U$61540 ( \61917 , \61888 , \61916 );
or \U$61541 ( \61918 , \61887 , \61915 );
nand \U$61542 ( \61919 , \61917 , \61918 );
not \U$61543 ( \61920 , \61919 );
and \U$61544 ( \61921 , \4688 , RIae78350_108);
and \U$61545 ( \61922 , RIae78170_104, \4686 );
nor \U$61546 ( \61923 , \61921 , \61922 );
and \U$61547 ( \61924 , \61923 , \4482 );
not \U$61548 ( \61925 , \61923 );
and \U$61549 ( \61926 , \61925 , \4481 );
nor \U$61550 ( \61927 , \61924 , \61926 );
and \U$61551 ( \61928 , \3730 , RIae77108_69);
and \U$61552 ( \61929 , RIae77090_68, \3728 );
nor \U$61553 ( \61930 , \61928 , \61929 );
and \U$61554 ( \61931 , \61930 , \3422 );
not \U$61555 ( \61932 , \61930 );
and \U$61556 ( \61933 , \61932 , \3732 );
nor \U$61557 ( \61934 , \61931 , \61933 );
xor \U$61558 ( \61935 , \61927 , \61934 );
and \U$61559 ( \61936 , \4247 , RIae77270_72);
and \U$61560 ( \61937 , RIae77360_74, \4245 );
nor \U$61561 ( \61938 , \61936 , \61937 );
and \U$61562 ( \61939 , \61938 , \4251 );
not \U$61563 ( \61940 , \61938 );
and \U$61564 ( \61941 , \61940 , \3989 );
nor \U$61565 ( \61942 , \61939 , \61941 );
xor \U$61566 ( \61943 , \61935 , \61942 );
not \U$61567 ( \61944 , \61943 );
and \U$61568 ( \61945 , \61920 , \61944 );
and \U$61569 ( \61946 , \61919 , \61943 );
nor \U$61570 ( \61947 , \61945 , \61946 );
and \U$61571 ( \61948 , \8371 , RIae789e0_122);
and \U$61572 ( \61949 , RIae788f0_120, \8369 );
nor \U$61573 ( \61950 , \61948 , \61949 );
and \U$61574 ( \61951 , \61950 , \8019 );
not \U$61575 ( \61952 , \61950 );
and \U$61576 ( \61953 , \61952 , \8020 );
nor \U$61577 ( \61954 , \61951 , \61953 );
and \U$61578 ( \61955 , \6941 , RIae77cc0_94);
and \U$61579 ( \61956 , RIae77bd0_92, \6939 );
nor \U$61580 ( \61957 , \61955 , \61956 );
and \U$61581 ( \61958 , \61957 , \6945 );
not \U$61582 ( \61959 , \61957 );
and \U$61583 ( \61960 , \61959 , \6314 );
nor \U$61584 ( \61961 , \61958 , \61960 );
xor \U$61585 ( \61962 , \61954 , \61961 );
and \U$61586 ( \61963 , \7633 , RIae77db0_96);
and \U$61587 ( \61964 , RIae77ea0_98, \7631 );
nor \U$61588 ( \61965 , \61963 , \61964 );
and \U$61589 ( \61966 , \61965 , \7205 );
not \U$61590 ( \61967 , \61965 );
and \U$61591 ( \61968 , \61967 , \7206 );
nor \U$61592 ( \61969 , \61966 , \61968 );
xor \U$61593 ( \61970 , \61962 , \61969 );
not \U$61594 ( \61971 , \61970 );
and \U$61595 ( \61972 , \11470 , RIae75fb0_32);
and \U$61596 ( \61973 , RIae75ec0_30, \11468 );
nor \U$61597 ( \61974 , \61972 , \61973 );
and \U$61598 ( \61975 , \61974 , \11474 );
not \U$61599 ( \61976 , \61974 );
and \U$61600 ( \61977 , \61976 , \10936 );
nor \U$61601 ( \61978 , \61975 , \61977 );
not \U$61602 ( \61979 , \61978 );
and \U$61603 ( \61980 , \12180 , RIae75ce0_26);
and \U$61604 ( \61981 , RIae75dd0_28, \12178 );
nor \U$61605 ( \61982 , \61980 , \61981 );
and \U$61606 ( \61983 , \61982 , \11827 );
not \U$61607 ( \61984 , \61982 );
and \U$61608 ( \61985 , \61984 , \12184 );
nor \U$61609 ( \61986 , \61983 , \61985 );
and \U$61610 ( \61987 , \13059 , RIae75650_12);
and \U$61611 ( \61988 , RIae75560_10, \13057 );
nor \U$61612 ( \61989 , \61987 , \61988 );
and \U$61613 ( \61990 , \61989 , \12718 );
not \U$61614 ( \61991 , \61989 );
and \U$61615 ( \61992 , \61991 , \13063 );
nor \U$61616 ( \61993 , \61990 , \61992 );
xor \U$61617 ( \61994 , \61986 , \61993 );
not \U$61618 ( \61995 , \61994 );
or \U$61619 ( \61996 , \61979 , \61995 );
or \U$61620 ( \61997 , \61994 , \61978 );
nand \U$61621 ( \61998 , \61996 , \61997 );
not \U$61622 ( \61999 , \61998 );
or \U$61623 ( \62000 , \61971 , \61999 );
or \U$61624 ( \62001 , \61970 , \61998 );
nand \U$61625 ( \62002 , \62000 , \62001 );
not \U$61626 ( \62003 , \62002 );
and \U$61627 ( \62004 , \10548 , RIae75a10_20);
and \U$61628 ( \62005 , RIae75920_18, \10546 );
nor \U$61629 ( \62006 , \62004 , \62005 );
and \U$61630 ( \62007 , \62006 , \10118 );
not \U$61631 ( \62008 , \62006 );
and \U$61632 ( \62009 , \62008 , \10421 );
nor \U$61633 ( \62010 , \62007 , \62009 );
and \U$61634 ( \62011 , \8966 , RIae78800_118);
and \U$61635 ( \62012 , RIae78710_116, \8964 );
nor \U$61636 ( \62013 , \62011 , \62012 );
and \U$61637 ( \62014 , \62013 , \8789 );
not \U$61638 ( \62015 , \62013 );
and \U$61639 ( \62016 , \62015 , \8799 );
nor \U$61640 ( \62017 , \62014 , \62016 );
xor \U$61641 ( \62018 , \62010 , \62017 );
and \U$61642 ( \62019 , \9760 , RIae75bf0_24);
and \U$61643 ( \62020 , RIae75b00_22, \9758 );
nor \U$61644 ( \62021 , \62019 , \62020 );
and \U$61645 ( \62022 , \62021 , \9272 );
not \U$61646 ( \62023 , \62021 );
and \U$61647 ( \62024 , \62023 , \9273 );
nor \U$61648 ( \62025 , \62022 , \62024 );
xor \U$61649 ( \62026 , \62018 , \62025 );
not \U$61650 ( \62027 , \62026 );
and \U$61651 ( \62028 , \62003 , \62027 );
and \U$61652 ( \62029 , \62002 , \62026 );
nor \U$61653 ( \62030 , \62028 , \62029 );
xor \U$61654 ( \62031 , \61947 , \62030 );
not \U$61655 ( \62032 , \62031 );
or \U$61656 ( \62033 , \61862 , \62032 );
or \U$61657 ( \62034 , \62031 , \61861 );
nand \U$61658 ( \62035 , \62033 , \62034 );
xor \U$61659 ( \62036 , \61824 , \62035 );
xor \U$61660 ( \62037 , \61711 , \61715 );
and \U$61661 ( \62038 , \62037 , \61720 );
and \U$61662 ( \62039 , \61711 , \61715 );
or \U$61663 ( \62040 , \62038 , \62039 );
xor \U$61664 ( \62041 , \61725 , \61731 );
and \U$61665 ( \62042 , \62041 , \61738 );
and \U$61666 ( \62043 , \61725 , \61731 );
or \U$61667 ( \62044 , \62042 , \62043 );
xor \U$61668 ( \62045 , \62040 , \62044 );
xor \U$61669 ( \62046 , \61577 , \61582 );
and \U$61670 ( \62047 , \62046 , \61610 );
and \U$61671 ( \62048 , \61577 , \61582 );
or \U$61672 ( \62049 , \62047 , \62048 );
xor \U$61673 ( \62050 , \62045 , \62049 );
and \U$61674 ( \62051 , \14964 , RIae75290_4);
and \U$61675 ( \62052 , RIae751a0_2, \14962 );
nor \U$61676 ( \62053 , \62051 , \62052 );
and \U$61677 ( \62054 , \62053 , \14462 );
not \U$61678 ( \62055 , \62053 );
and \U$61679 ( \62056 , \62055 , \14463 );
nor \U$61680 ( \62057 , \62054 , \62056 );
and \U$61681 ( \62058 , \15726 , RIae75380_6);
and \U$61682 ( \62059 , RIae75470_8, RIae7aab0_192);
nor \U$61683 ( \62060 , \62058 , \62059 );
and \U$61684 ( \62061 , \62060 , RIae7aa38_191);
not \U$61685 ( \62062 , \62060 );
and \U$61686 ( \62063 , \62062 , \14959 );
nor \U$61687 ( \62064 , \62061 , \62063 );
xor \U$61688 ( \62065 , \62057 , \62064 );
and \U$61689 ( \62066 , \14059 , RIae75830_16);
and \U$61690 ( \62067 , RIae75740_14, \14057 );
nor \U$61691 ( \62068 , \62066 , \62067 );
and \U$61692 ( \62069 , \62068 , \14063 );
not \U$61693 ( \62070 , \62068 );
and \U$61694 ( \62071 , \62070 , \13502 );
nor \U$61695 ( \62072 , \62069 , \62071 );
xor \U$61696 ( \62073 , \62065 , \62072 );
not \U$61697 ( \62074 , \62073 );
xor \U$61698 ( \62075 , \61641 , \61664 );
and \U$61699 ( \62076 , \62075 , \61688 );
and \U$61700 ( \62077 , \61641 , \61664 );
nor \U$61701 ( \62078 , \62076 , \62077 );
xor \U$61702 ( \62079 , \61507 , \61514 );
xor \U$61703 ( \62080 , \62079 , \61522 );
and \U$61704 ( \62081 , \61546 , \62080 );
xor \U$61705 ( \62082 , \61507 , \61514 );
xor \U$61706 ( \62083 , \62082 , \61522 );
and \U$61707 ( \62084 , \61569 , \62083 );
and \U$61708 ( \62085 , \61546 , \61569 );
or \U$61709 ( \62086 , \62081 , \62084 , \62085 );
not \U$61710 ( \62087 , \62086 );
xor \U$61711 ( \62088 , \62078 , \62087 );
not \U$61712 ( \62089 , \62088 );
or \U$61713 ( \62090 , \62074 , \62089 );
or \U$61714 ( \62091 , \62088 , \62073 );
nand \U$61715 ( \62092 , \62090 , \62091 );
xor \U$61716 ( \62093 , \62050 , \62092 );
xor \U$61717 ( \62094 , \61462 , \61478 );
and \U$61718 ( \62095 , \62094 , \61485 );
and \U$61719 ( \62096 , \61462 , \61478 );
or \U$61720 ( \62097 , \62095 , \62096 );
xor \U$61721 ( \62098 , \61490 , \61494 );
and \U$61722 ( \62099 , \62098 , \61499 );
and \U$61723 ( \62100 , \61490 , \61494 );
or \U$61724 ( \62101 , \62099 , \62100 );
xor \U$61725 ( \62102 , \62097 , \62101 );
xor \U$61726 ( \62103 , \61571 , \61611 );
and \U$61727 ( \62104 , \62103 , \61689 );
and \U$61728 ( \62105 , \61571 , \61611 );
or \U$61729 ( \62106 , \62104 , \62105 );
xor \U$61730 ( \62107 , \62102 , \62106 );
xor \U$61731 ( \62108 , \62093 , \62107 );
xor \U$61732 ( \62109 , \62036 , \62108 );
xor \U$61733 ( \62110 , \61795 , \62109 );
not \U$61734 ( \62111 , \62110 );
and \U$61735 ( \62112 , \61768 , \62111 );
and \U$61736 ( \62113 , \61767 , \62110 );
nor \U$61737 ( \62114 , \62112 , \62113 );
xor \U$61738 ( \62115 , \61697 , \61703 );
and \U$61739 ( \62116 , \62115 , \61751 );
and \U$61740 ( \62117 , \61697 , \61703 );
nor \U$61741 ( \62118 , \62116 , \62117 );
xnor \U$61742 ( \62119 , \62114 , \62118 );
or \U$61743 ( \62120 , \61756 , \62119 );
or \U$61744 ( \62121 , \62114 , \62118 );
nand \U$61745 ( \62122 , \62120 , \62121 );
xor \U$61746 ( \62123 , \61776 , \61784 );
and \U$61747 ( \62124 , \62123 , \61793 );
and \U$61748 ( \62125 , \61776 , \61784 );
or \U$61749 ( \62126 , \62124 , \62125 );
xor \U$61750 ( \62127 , \61809 , \61823 );
xor \U$61751 ( \62128 , \62127 , \62035 );
and \U$61752 ( \62129 , \62093 , \62128 );
xor \U$61753 ( \62130 , \61809 , \61823 );
xor \U$61754 ( \62131 , \62130 , \62035 );
and \U$61755 ( \62132 , \62107 , \62131 );
and \U$61756 ( \62133 , \62093 , \62107 );
or \U$61757 ( \62134 , \62129 , \62132 , \62133 );
xor \U$61758 ( \62135 , \62126 , \62134 );
or \U$61759 ( \62136 , \61887 , \61943 );
not \U$61760 ( \62137 , \61943 );
not \U$61761 ( \62138 , \61887 );
or \U$61762 ( \62139 , \62137 , \62138 );
nand \U$61763 ( \62140 , \62139 , \61915 );
nand \U$61764 ( \62141 , \62136 , \62140 );
or \U$61765 ( \62142 , \61970 , \62026 );
not \U$61766 ( \62143 , \62026 );
not \U$61767 ( \62144 , \61970 );
or \U$61768 ( \62145 , \62143 , \62144 );
nand \U$61769 ( \62146 , \62145 , \61998 );
nand \U$61770 ( \62147 , \62142 , \62146 );
xor \U$61771 ( \62148 , \62141 , \62147 );
and \U$61772 ( \62149 , \11470 , RIae75ec0_30);
and \U$61773 ( \62150 , RIae75ce0_26, \11468 );
nor \U$61774 ( \62151 , \62149 , \62150 );
and \U$61775 ( \62152 , \62151 , \10936 );
not \U$61776 ( \62153 , \62151 );
and \U$61777 ( \62154 , \62153 , \11474 );
nor \U$61778 ( \62155 , \62152 , \62154 );
and \U$61779 ( \62156 , \9760 , RIae75b00_22);
and \U$61780 ( \62157 , RIae75a10_20, \9758 );
nor \U$61781 ( \62158 , \62156 , \62157 );
and \U$61782 ( \62159 , \62158 , \9273 );
not \U$61783 ( \62160 , \62158 );
and \U$61784 ( \62161 , \62160 , \9764 );
nor \U$61785 ( \62162 , \62159 , \62161 );
xor \U$61786 ( \62163 , \62155 , \62162 );
and \U$61787 ( \62164 , \10548 , RIae75920_18);
and \U$61788 ( \62165 , RIae75fb0_32, \10546 );
nor \U$61789 ( \62166 , \62164 , \62165 );
and \U$61790 ( \62167 , \62166 , \10421 );
not \U$61791 ( \62168 , \62166 );
and \U$61792 ( \62169 , \62168 , \10118 );
nor \U$61793 ( \62170 , \62167 , \62169 );
xor \U$61794 ( \62171 , \62163 , \62170 );
and \U$61795 ( \62172 , \15726 , RIae75470_8);
and \U$61796 ( \62173 , RIae76460_42, RIae7aab0_192);
nor \U$61797 ( \62174 , \62172 , \62173 );
and \U$61798 ( \62175 , \62174 , \14959 );
not \U$61799 ( \62176 , \62174 );
and \U$61800 ( \62177 , \62176 , RIae7aa38_191);
nor \U$61801 ( \62178 , \62175 , \62177 );
xor \U$61802 ( \62179 , \62178 , \1261 );
and \U$61803 ( \62180 , \14964 , RIae751a0_2);
and \U$61804 ( \62181 , RIae75380_6, \14962 );
nor \U$61805 ( \62182 , \62180 , \62181 );
and \U$61806 ( \62183 , \62182 , \14463 );
not \U$61807 ( \62184 , \62182 );
and \U$61808 ( \62185 , \62184 , \14462 );
nor \U$61809 ( \62186 , \62183 , \62185 );
xor \U$61810 ( \62187 , \62179 , \62186 );
and \U$61811 ( \62188 , \14059 , RIae75740_14);
and \U$61812 ( \62189 , RIae75290_4, \14057 );
nor \U$61813 ( \62190 , \62188 , \62189 );
and \U$61814 ( \62191 , \62190 , \13502 );
not \U$61815 ( \62192 , \62190 );
and \U$61816 ( \62193 , \62192 , \14063 );
nor \U$61817 ( \62194 , \62191 , \62193 );
and \U$61818 ( \62195 , \12180 , RIae75dd0_28);
and \U$61819 ( \62196 , RIae75650_12, \12178 );
nor \U$61820 ( \62197 , \62195 , \62196 );
and \U$61821 ( \62198 , \62197 , \12184 );
not \U$61822 ( \62199 , \62197 );
and \U$61823 ( \62200 , \62199 , \11827 );
nor \U$61824 ( \62201 , \62198 , \62200 );
xor \U$61825 ( \62202 , \62194 , \62201 );
and \U$61826 ( \62203 , \13059 , RIae75560_10);
and \U$61827 ( \62204 , RIae75830_16, \13057 );
nor \U$61828 ( \62205 , \62203 , \62204 );
and \U$61829 ( \62206 , \62205 , \13063 );
not \U$61830 ( \62207 , \62205 );
and \U$61831 ( \62208 , \62207 , \12718 );
nor \U$61832 ( \62209 , \62206 , \62208 );
xor \U$61833 ( \62210 , \62202 , \62209 );
xor \U$61834 ( \62211 , \62187 , \62210 );
xor \U$61835 ( \62212 , \62171 , \62211 );
xor \U$61836 ( \62213 , \62148 , \62212 );
not \U$61837 ( \62214 , \62213 );
xor \U$61838 ( \62215 , \61813 , \61817 );
and \U$61839 ( \62216 , \62215 , \61822 );
and \U$61840 ( \62217 , \61813 , \61817 );
nor \U$61841 ( \62218 , \62216 , \62217 );
xor \U$61842 ( \62219 , \61799 , \61803 );
and \U$61843 ( \62220 , \62219 , \61808 );
and \U$61844 ( \62221 , \61799 , \61803 );
nor \U$61845 ( \62222 , \62220 , \62221 );
xor \U$61846 ( \62223 , \62218 , \62222 );
xor \U$61847 ( \62224 , \61830 , \61836 );
and \U$61848 ( \62225 , \62224 , \61860 );
and \U$61849 ( \62226 , \61830 , \61836 );
or \U$61850 ( \62227 , \62225 , \62226 );
xor \U$61851 ( \62228 , \62223 , \62227 );
not \U$61852 ( \62229 , \62228 );
and \U$61853 ( \62230 , \62214 , \62229 );
and \U$61854 ( \62231 , \62213 , \62228 );
nor \U$61855 ( \62232 , \62230 , \62231 );
not \U$61856 ( \62233 , \62232 );
xor \U$61857 ( \62234 , \61927 , \61934 );
and \U$61858 ( \62235 , \62234 , \61942 );
and \U$61859 ( \62236 , \61927 , \61934 );
or \U$61860 ( \62237 , \62235 , \62236 );
not \U$61861 ( \62238 , \61895 );
not \U$61862 ( \62239 , \61903 );
and \U$61863 ( \62240 , \62238 , \62239 );
and \U$61864 ( \62241 , \61903 , \61895 );
nor \U$61865 ( \62242 , \62241 , \61910 );
nor \U$61866 ( \62243 , \62240 , \62242 );
xor \U$61867 ( \62244 , \62237 , \62243 );
xor \U$61868 ( \62245 , \61954 , \61961 );
and \U$61869 ( \62246 , \62245 , \61969 );
and \U$61870 ( \62247 , \61954 , \61961 );
or \U$61871 ( \62248 , \62246 , \62247 );
xor \U$61872 ( \62249 , \62244 , \62248 );
xor \U$61873 ( \62250 , \62057 , \62064 );
and \U$61874 ( \62251 , \62250 , \62072 );
and \U$61875 ( \62252 , \62057 , \62064 );
or \U$61876 ( \62253 , \62251 , \62252 );
not \U$61877 ( \62254 , \61978 );
not \U$61878 ( \62255 , \61986 );
and \U$61879 ( \62256 , \62254 , \62255 );
and \U$61880 ( \62257 , \61986 , \61978 );
nor \U$61881 ( \62258 , \62257 , \61993 );
nor \U$61882 ( \62259 , \62256 , \62258 );
xor \U$61883 ( \62260 , \62253 , \62259 );
xor \U$61884 ( \62261 , \62010 , \62017 );
and \U$61885 ( \62262 , \62261 , \62025 );
and \U$61886 ( \62263 , \62010 , \62017 );
or \U$61887 ( \62264 , \62262 , \62263 );
xor \U$61888 ( \62265 , \62260 , \62264 );
xor \U$61889 ( \62266 , \62249 , \62265 );
xor \U$61890 ( \62267 , \61870 , \61878 );
and \U$61891 ( \62268 , \62267 , \61886 );
and \U$61892 ( \62269 , \61870 , \61878 );
nor \U$61893 ( \62270 , \62268 , \62269 );
not \U$61894 ( \62271 , \62270 );
xor \U$61895 ( \62272 , \61844 , \61851 );
and \U$61896 ( \62273 , \62272 , \61859 );
and \U$61897 ( \62274 , \61844 , \61851 );
or \U$61898 ( \62275 , \62273 , \62274 );
not \U$61899 ( \62276 , \62275 );
or \U$61900 ( \62277 , \62271 , \62276 );
or \U$61901 ( \62278 , \62275 , \62270 );
nand \U$61902 ( \62279 , \62277 , \62278 );
not \U$61903 ( \62280 , \62279 );
and \U$61904 ( \62281 , \1593 , RIae77540_78);
and \U$61905 ( \62282 , RIae776a8_81, \1591 );
nor \U$61906 ( \62283 , \62281 , \62282 );
and \U$61907 ( \62284 , \62283 , \1488 );
not \U$61908 ( \62285 , \62283 );
and \U$61909 ( \62286 , \62285 , \1498 );
nor \U$61910 ( \62287 , \62284 , \62286 );
not \U$61911 ( \62288 , \62287 );
and \U$61912 ( \62289 , \62280 , \62288 );
and \U$61913 ( \62290 , \62279 , \62287 );
nor \U$61914 ( \62291 , \62289 , \62290 );
not \U$61915 ( \62292 , \62291 );
and \U$61916 ( \62293 , \3730 , RIae77090_68);
and \U$61917 ( \62294 , RIae77270_72, \3728 );
nor \U$61918 ( \62295 , \62293 , \62294 );
and \U$61919 ( \62296 , \62295 , \3732 );
not \U$61920 ( \62297 , \62295 );
and \U$61921 ( \62298 , \62297 , \3422 );
nor \U$61922 ( \62299 , \62296 , \62298 );
not \U$61923 ( \62300 , \2789 );
and \U$61924 ( \62301 , \2783 , RIae76eb0_64);
and \U$61925 ( \62302 , RIae76dc0_62, \2781 );
nor \U$61926 ( \62303 , \62301 , \62302 );
not \U$61927 ( \62304 , \62303 );
or \U$61928 ( \62305 , \62300 , \62304 );
or \U$61929 ( \62306 , \62303 , \3089 );
nand \U$61930 ( \62307 , \62305 , \62306 );
xor \U$61931 ( \62308 , \62299 , \62307 );
not \U$61932 ( \62309 , \2774 );
and \U$61933 ( \62310 , \3214 , RIae76cd0_60);
and \U$61934 ( \62311 , RIae77108_69, \3212 );
nor \U$61935 ( \62312 , \62310 , \62311 );
not \U$61936 ( \62313 , \62312 );
or \U$61937 ( \62314 , \62309 , \62313 );
or \U$61938 ( \62315 , \62312 , \3218 );
nand \U$61939 ( \62316 , \62314 , \62315 );
xor \U$61940 ( \62317 , \62308 , \62316 );
nand \U$61941 ( \62318 , RIae77630_80, \1374 );
and \U$61942 ( \62319 , \62318 , \1380 );
not \U$61943 ( \62320 , \62318 );
and \U$61944 ( \62321 , \62320 , \1261 );
nor \U$61945 ( \62322 , \62319 , \62321 );
and \U$61946 ( \62323 , \2607 , RIae77900_86);
and \U$61947 ( \62324 , RIae76fa0_66, \2605 );
nor \U$61948 ( \62325 , \62323 , \62324 );
and \U$61949 ( \62326 , \62325 , \2611 );
not \U$61950 ( \62327 , \62325 );
and \U$61951 ( \62328 , \62327 , \2397 );
nor \U$61952 ( \62329 , \62326 , \62328 );
and \U$61953 ( \62330 , \1939 , RIae77450_76);
and \U$61954 ( \62331 , RIae77ae0_90, \1937 );
nor \U$61955 ( \62332 , \62330 , \62331 );
and \U$61956 ( \62333 , \62332 , \1735 );
not \U$61957 ( \62334 , \62332 );
and \U$61958 ( \62335 , \62334 , \1734 );
nor \U$61959 ( \62336 , \62333 , \62335 );
xor \U$61960 ( \62337 , \62329 , \62336 );
and \U$61961 ( \62338 , \2224 , RIae779f0_88);
and \U$61962 ( \62339 , RIae77810_84, \2222 );
nor \U$61963 ( \62340 , \62338 , \62339 );
and \U$61964 ( \62341 , \62340 , \2061 );
not \U$61965 ( \62342 , \62340 );
and \U$61966 ( \62343 , \62342 , \2060 );
nor \U$61967 ( \62344 , \62341 , \62343 );
xor \U$61968 ( \62345 , \62337 , \62344 );
xor \U$61969 ( \62346 , \62322 , \62345 );
xor \U$61970 ( \62347 , \62317 , \62346 );
not \U$61971 ( \62348 , \62347 );
or \U$61972 ( \62349 , \62292 , \62348 );
or \U$61973 ( \62350 , \62347 , \62291 );
nand \U$61974 ( \62351 , \62349 , \62350 );
not \U$61975 ( \62352 , \62351 );
and \U$61976 ( \62353 , \8371 , RIae788f0_120);
and \U$61977 ( \62354 , RIae78800_118, \8369 );
nor \U$61978 ( \62355 , \62353 , \62354 );
and \U$61979 ( \62356 , \62355 , \8019 );
not \U$61980 ( \62357 , \62355 );
and \U$61981 ( \62358 , \62357 , \8020 );
nor \U$61982 ( \62359 , \62356 , \62358 );
not \U$61983 ( \62360 , \62359 );
and \U$61984 ( \62361 , \8966 , RIae78710_116);
and \U$61985 ( \62362 , RIae75bf0_24, \8964 );
nor \U$61986 ( \62363 , \62361 , \62362 );
and \U$61987 ( \62364 , \62363 , \8799 );
not \U$61988 ( \62365 , \62363 );
and \U$61989 ( \62366 , \62365 , \8789 );
nor \U$61990 ( \62367 , \62364 , \62366 );
not \U$61991 ( \62368 , \62367 );
or \U$61992 ( \62369 , \62360 , \62368 );
or \U$61993 ( \62370 , \62359 , \62367 );
nand \U$61994 ( \62371 , \62369 , \62370 );
not \U$61995 ( \62372 , \62371 );
and \U$61996 ( \62373 , \7633 , RIae77ea0_98);
and \U$61997 ( \62374 , RIae789e0_122, \7631 );
nor \U$61998 ( \62375 , \62373 , \62374 );
and \U$61999 ( \62376 , \62375 , \7205 );
not \U$62000 ( \62377 , \62375 );
and \U$62001 ( \62378 , \62377 , \7206 );
nor \U$62002 ( \62379 , \62376 , \62378 );
not \U$62003 ( \62380 , \62379 );
and \U$62004 ( \62381 , \62372 , \62380 );
and \U$62005 ( \62382 , \62371 , \62379 );
nor \U$62006 ( \62383 , \62381 , \62382 );
not \U$62007 ( \62384 , \62383 );
and \U$62008 ( \62385 , \6941 , RIae77bd0_92);
and \U$62009 ( \62386 , RIae77db0_96, \6939 );
nor \U$62010 ( \62387 , \62385 , \62386 );
and \U$62011 ( \62388 , \62387 , \6314 );
not \U$62012 ( \62389 , \62387 );
and \U$62013 ( \62390 , \62389 , \6945 );
nor \U$62014 ( \62391 , \62388 , \62390 );
and \U$62015 ( \62392 , \5896 , RIae78620_114);
and \U$62016 ( \62393 , RIae78440_110, \5894 );
nor \U$62017 ( \62394 , \62392 , \62393 );
and \U$62018 ( \62395 , \62394 , \5590 );
not \U$62019 ( \62396 , \62394 );
and \U$62020 ( \62397 , \62396 , \5589 );
nor \U$62021 ( \62398 , \62395 , \62397 );
xor \U$62022 ( \62399 , \62391 , \62398 );
and \U$62023 ( \62400 , \6172 , RIae784b8_111);
and \U$62024 ( \62401 , RIae77cc0_94, \6170 );
nor \U$62025 ( \62402 , \62400 , \62401 );
and \U$62026 ( \62403 , \62402 , \6176 );
not \U$62027 ( \62404 , \62402 );
and \U$62028 ( \62405 , \62404 , \6175 );
nor \U$62029 ( \62406 , \62403 , \62405 );
xor \U$62030 ( \62407 , \62399 , \62406 );
not \U$62031 ( \62408 , \62407 );
or \U$62032 ( \62409 , \62384 , \62408 );
or \U$62033 ( \62410 , \62383 , \62407 );
nand \U$62034 ( \62411 , \62409 , \62410 );
not \U$62035 ( \62412 , \62411 );
and \U$62036 ( \62413 , \4688 , RIae78170_104);
and \U$62037 ( \62414 , RIae77f90_100, \4686 );
nor \U$62038 ( \62415 , \62413 , \62414 );
and \U$62039 ( \62416 , \62415 , \4482 );
not \U$62040 ( \62417 , \62415 );
and \U$62041 ( \62418 , \62417 , \4481 );
nor \U$62042 ( \62419 , \62416 , \62418 );
not \U$62043 ( \62420 , \62419 );
and \U$62044 ( \62421 , \5399 , RIae78080_102);
and \U$62045 ( \62422 , RIae78260_106, \5397 );
nor \U$62046 ( \62423 , \62421 , \62422 );
and \U$62047 ( \62424 , \62423 , \5016 );
not \U$62048 ( \62425 , \62423 );
and \U$62049 ( \62426 , \62425 , \5403 );
nor \U$62050 ( \62427 , \62424 , \62426 );
not \U$62051 ( \62428 , \62427 );
or \U$62052 ( \62429 , \62420 , \62428 );
or \U$62053 ( \62430 , \62419 , \62427 );
nand \U$62054 ( \62431 , \62429 , \62430 );
not \U$62055 ( \62432 , \62431 );
and \U$62056 ( \62433 , \4247 , RIae77360_74);
and \U$62057 ( \62434 , RIae78350_108, \4245 );
nor \U$62058 ( \62435 , \62433 , \62434 );
and \U$62059 ( \62436 , \62435 , \4251 );
not \U$62060 ( \62437 , \62435 );
and \U$62061 ( \62438 , \62437 , \3989 );
nor \U$62062 ( \62439 , \62436 , \62438 );
not \U$62063 ( \62440 , \62439 );
and \U$62064 ( \62441 , \62432 , \62440 );
and \U$62065 ( \62442 , \62431 , \62439 );
nor \U$62066 ( \62443 , \62441 , \62442 );
not \U$62067 ( \62444 , \62443 );
and \U$62068 ( \62445 , \62412 , \62444 );
and \U$62069 ( \62446 , \62411 , \62443 );
nor \U$62070 ( \62447 , \62445 , \62446 );
not \U$62071 ( \62448 , \62447 );
and \U$62072 ( \62449 , \62352 , \62448 );
and \U$62073 ( \62450 , \62351 , \62447 );
nor \U$62074 ( \62451 , \62449 , \62450 );
xor \U$62075 ( \62452 , \62266 , \62451 );
xor \U$62076 ( \62453 , \62040 , \62044 );
and \U$62077 ( \62454 , \62453 , \62049 );
and \U$62078 ( \62455 , \62040 , \62044 );
nor \U$62079 ( \62456 , \62454 , \62455 );
not \U$62080 ( \62457 , \62078 );
not \U$62081 ( \62458 , \62073 );
and \U$62082 ( \62459 , \62457 , \62458 );
and \U$62083 ( \62460 , \62078 , \62073 );
nor \U$62084 ( \62461 , \62460 , \62087 );
nor \U$62085 ( \62462 , \62459 , \62461 );
xor \U$62086 ( \62463 , \62456 , \62462 );
not \U$62087 ( \62464 , \61947 );
not \U$62088 ( \62465 , \61861 );
and \U$62089 ( \62466 , \62464 , \62465 );
and \U$62090 ( \62467 , \61947 , \61861 );
nor \U$62091 ( \62468 , \62467 , \62030 );
nor \U$62092 ( \62469 , \62466 , \62468 );
xor \U$62093 ( \62470 , \62463 , \62469 );
xor \U$62094 ( \62471 , \62452 , \62470 );
not \U$62095 ( \62472 , \62471 );
or \U$62096 ( \62473 , \62233 , \62472 );
or \U$62097 ( \62474 , \62471 , \62232 );
nand \U$62098 ( \62475 , \62473 , \62474 );
xor \U$62099 ( \62476 , \62135 , \62475 );
and \U$62100 ( \62477 , \62050 , \62092 );
xor \U$62101 ( \62478 , \61809 , \61823 );
and \U$62102 ( \62479 , \62478 , \62035 );
and \U$62103 ( \62480 , \61809 , \61823 );
or \U$62104 ( \62481 , \62479 , \62480 );
xor \U$62105 ( \62482 , \62477 , \62481 );
xor \U$62106 ( \62483 , \62097 , \62101 );
and \U$62107 ( \62484 , \62483 , \62106 );
and \U$62108 ( \62485 , \62097 , \62101 );
or \U$62109 ( \62486 , \62484 , \62485 );
xor \U$62110 ( \62487 , \62482 , \62486 );
xor \U$62111 ( \62488 , \62476 , \62487 );
xor \U$62112 ( \62489 , \61772 , \61794 );
and \U$62113 ( \62490 , \62489 , \62109 );
and \U$62114 ( \62491 , \61772 , \61794 );
or \U$62115 ( \62492 , \62490 , \62491 );
xor \U$62116 ( \62493 , \62488 , \62492 );
not \U$62117 ( \62494 , \62110 );
or \U$62118 ( \62495 , \62494 , \61758 );
not \U$62119 ( \62496 , \61758 );
not \U$62120 ( \62497 , \62494 );
or \U$62121 ( \62498 , \62496 , \62497 );
nand \U$62122 ( \62499 , \62498 , \61763 );
nand \U$62123 ( \62500 , \62495 , \62499 );
xor \U$62124 ( \62501 , \62493 , \62500 );
and \U$62125 ( \62502 , \62122 , \62501 );
and \U$62126 ( \62503 , \62493 , \62500 );
nor \U$62127 ( \62504 , \62502 , \62503 );
xor \U$62128 ( \62505 , \62456 , \62462 );
and \U$62129 ( \62506 , \62505 , \62469 );
and \U$62130 ( \62507 , \62456 , \62462 );
nor \U$62131 ( \62508 , \62506 , \62507 );
not \U$62132 ( \62509 , \62508 );
xor \U$62133 ( \62510 , \62249 , \62265 );
and \U$62134 ( \62511 , \62510 , \62451 );
and \U$62135 ( \62512 , \62249 , \62265 );
or \U$62136 ( \62513 , \62511 , \62512 );
not \U$62137 ( \62514 , \62513 );
or \U$62138 ( \62515 , \62509 , \62514 );
or \U$62139 ( \62516 , \62513 , \62508 );
nand \U$62140 ( \62517 , \62515 , \62516 );
not \U$62141 ( \62518 , \62517 );
not \U$62142 ( \62519 , \62228 );
nand \U$62143 ( \62520 , \62519 , \62213 );
not \U$62144 ( \62521 , \62520 );
and \U$62145 ( \62522 , \62518 , \62521 );
and \U$62146 ( \62523 , \62517 , \62520 );
nor \U$62147 ( \62524 , \62522 , \62523 );
not \U$62148 ( \62525 , \62524 );
xor \U$62149 ( \62526 , \62126 , \62134 );
and \U$62150 ( \62527 , \62526 , \62475 );
and \U$62151 ( \62528 , \62126 , \62134 );
or \U$62152 ( \62529 , \62527 , \62528 );
not \U$62153 ( \62530 , \62529 );
or \U$62154 ( \62531 , \62525 , \62530 );
or \U$62155 ( \62532 , \62529 , \62524 );
nand \U$62156 ( \62533 , \62531 , \62532 );
not \U$62157 ( \62534 , \62533 );
xor \U$62158 ( \62535 , \62477 , \62481 );
and \U$62159 ( \62536 , \62535 , \62486 );
and \U$62160 ( \62537 , \62477 , \62481 );
nor \U$62161 ( \62538 , \62536 , \62537 );
not \U$62162 ( \62539 , \62470 );
not \U$62163 ( \62540 , \62232 );
and \U$62164 ( \62541 , \62539 , \62540 );
and \U$62165 ( \62542 , \62470 , \62232 );
nor \U$62166 ( \62543 , \62542 , \62452 );
nor \U$62167 ( \62544 , \62541 , \62543 );
xnor \U$62168 ( \62545 , \62538 , \62544 );
not \U$62169 ( \62546 , \62545 );
xor \U$62170 ( \62547 , \62141 , \62147 );
and \U$62171 ( \62548 , \62547 , \62212 );
and \U$62172 ( \62549 , \62141 , \62147 );
or \U$62173 ( \62550 , \62548 , \62549 );
xor \U$62174 ( \62551 , \62218 , \62222 );
and \U$62175 ( \62552 , \62551 , \62227 );
and \U$62176 ( \62553 , \62218 , \62222 );
nor \U$62177 ( \62554 , \62552 , \62553 );
xor \U$62178 ( \62555 , \62550 , \62554 );
or \U$62179 ( \62556 , \62447 , \62291 );
not \U$62180 ( \62557 , \62291 );
not \U$62181 ( \62558 , \62447 );
or \U$62182 ( \62559 , \62557 , \62558 );
nand \U$62183 ( \62560 , \62559 , \62347 );
nand \U$62184 ( \62561 , \62556 , \62560 );
xor \U$62185 ( \62562 , \62555 , \62561 );
xor \U$62186 ( \62563 , \62253 , \62259 );
and \U$62187 ( \62564 , \62563 , \62264 );
and \U$62188 ( \62565 , \62253 , \62259 );
nor \U$62189 ( \62566 , \62564 , \62565 );
or \U$62190 ( \62567 , \62275 , \62287 );
not \U$62191 ( \62568 , \62287 );
not \U$62192 ( \62569 , \62275 );
or \U$62193 ( \62570 , \62568 , \62569 );
nand \U$62194 ( \62571 , \62570 , \62270 );
nand \U$62195 ( \62572 , \62567 , \62571 );
xor \U$62196 ( \62573 , \62566 , \62572 );
xor \U$62197 ( \62574 , \62237 , \62243 );
and \U$62198 ( \62575 , \62574 , \62248 );
and \U$62199 ( \62576 , \62237 , \62243 );
nor \U$62200 ( \62577 , \62575 , \62576 );
xor \U$62201 ( \62578 , \62573 , \62577 );
xor \U$62202 ( \62579 , \62155 , \62162 );
xor \U$62203 ( \62580 , \62579 , \62170 );
and \U$62204 ( \62581 , \62187 , \62580 );
xor \U$62205 ( \62582 , \62155 , \62162 );
xor \U$62206 ( \62583 , \62582 , \62170 );
and \U$62207 ( \62584 , \62210 , \62583 );
and \U$62208 ( \62585 , \62187 , \62210 );
or \U$62209 ( \62586 , \62581 , \62584 , \62585 );
xor \U$62210 ( \62587 , \62299 , \62307 );
xor \U$62211 ( \62588 , \62587 , \62316 );
and \U$62212 ( \62589 , \62322 , \62588 );
xor \U$62213 ( \62590 , \62299 , \62307 );
xor \U$62214 ( \62591 , \62590 , \62316 );
and \U$62215 ( \62592 , \62345 , \62591 );
and \U$62216 ( \62593 , \62322 , \62345 );
or \U$62217 ( \62594 , \62589 , \62592 , \62593 );
xor \U$62218 ( \62595 , \62586 , \62594 );
or \U$62219 ( \62596 , \62443 , \62383 );
not \U$62220 ( \62597 , \62383 );
not \U$62221 ( \62598 , \62443 );
or \U$62222 ( \62599 , \62597 , \62598 );
nand \U$62223 ( \62600 , \62599 , \62407 );
nand \U$62224 ( \62601 , \62596 , \62600 );
xor \U$62225 ( \62602 , \62595 , \62601 );
xor \U$62226 ( \62603 , \62329 , \62336 );
and \U$62227 ( \62604 , \62603 , \62344 );
and \U$62228 ( \62605 , \62329 , \62336 );
or \U$62229 ( \62606 , \62604 , \62605 );
and \U$62230 ( \62607 , \1376 , RIae77630_80);
and \U$62231 ( \62608 , RIae77540_78, \1374 );
nor \U$62232 ( \62609 , \62607 , \62608 );
and \U$62233 ( \62610 , \62609 , \1380 );
not \U$62234 ( \62611 , \62609 );
and \U$62235 ( \62612 , \62611 , \1261 );
nor \U$62236 ( \62613 , \62610 , \62612 );
xor \U$62237 ( \62614 , \62606 , \62613 );
xor \U$62238 ( \62615 , \62299 , \62307 );
and \U$62239 ( \62616 , \62615 , \62316 );
and \U$62240 ( \62617 , \62299 , \62307 );
or \U$62241 ( \62618 , \62616 , \62617 );
xor \U$62242 ( \62619 , \62614 , \62618 );
xor \U$62243 ( \62620 , \62194 , \62201 );
and \U$62244 ( \62621 , \62620 , \62209 );
and \U$62245 ( \62622 , \62194 , \62201 );
or \U$62246 ( \62623 , \62621 , \62622 );
xor \U$62247 ( \62624 , \62178 , \1261 );
and \U$62248 ( \62625 , \62624 , \62186 );
and \U$62249 ( \62626 , \62178 , \1261 );
or \U$62250 ( \62627 , \62625 , \62626 );
xor \U$62251 ( \62628 , \62623 , \62627 );
xor \U$62252 ( \62629 , \62155 , \62162 );
and \U$62253 ( \62630 , \62629 , \62170 );
and \U$62254 ( \62631 , \62155 , \62162 );
or \U$62255 ( \62632 , \62630 , \62631 );
xor \U$62256 ( \62633 , \62628 , \62632 );
xor \U$62257 ( \62634 , \62391 , \62398 );
and \U$62258 ( \62635 , \62634 , \62406 );
and \U$62259 ( \62636 , \62391 , \62398 );
or \U$62260 ( \62637 , \62635 , \62636 );
or \U$62261 ( \62638 , \62439 , \62419 );
not \U$62262 ( \62639 , \62419 );
not \U$62263 ( \62640 , \62439 );
or \U$62264 ( \62641 , \62639 , \62640 );
nand \U$62265 ( \62642 , \62641 , \62427 );
nand \U$62266 ( \62643 , \62638 , \62642 );
xor \U$62267 ( \62644 , \62637 , \62643 );
or \U$62268 ( \62645 , \62379 , \62359 );
not \U$62269 ( \62646 , \62359 );
not \U$62270 ( \62647 , \62379 );
or \U$62271 ( \62648 , \62646 , \62647 );
nand \U$62272 ( \62649 , \62648 , \62367 );
nand \U$62273 ( \62650 , \62645 , \62649 );
xor \U$62274 ( \62651 , \62644 , \62650 );
xor \U$62275 ( \62652 , \62633 , \62651 );
xor \U$62276 ( \62653 , \62619 , \62652 );
xor \U$62277 ( \62654 , \53137 , \53144 );
xor \U$62278 ( \62655 , \62654 , \53152 );
xor \U$62279 ( \62656 , \53109 , \53116 );
xor \U$62280 ( \62657 , \62656 , \53124 );
xor \U$62281 ( \62658 , \62655 , \62657 );
xor \U$62282 ( \62659 , \53058 , \53065 );
xor \U$62283 ( \62660 , \62659 , \53073 );
xor \U$62284 ( \62661 , \62658 , \62660 );
xor \U$62285 ( \62662 , \53188 , \53195 );
xor \U$62286 ( \62663 , \62662 , \53203 );
xor \U$62287 ( \62664 , \53162 , \53169 );
xor \U$62288 ( \62665 , \62664 , \53177 );
xor \U$62289 ( \62666 , \62663 , \62665 );
xor \U$62290 ( \62667 , \53218 , \53225 );
xor \U$62291 ( \62668 , \62667 , \53234 );
xor \U$62292 ( \62669 , \53244 , \53251 );
xor \U$62293 ( \62670 , \62669 , \53259 );
xor \U$62294 ( \62671 , \53083 , \53090 );
xor \U$62295 ( \62672 , \62671 , \53098 );
xor \U$62296 ( \62673 , \62670 , \62672 );
xor \U$62297 ( \62674 , \62668 , \62673 );
xor \U$62298 ( \62675 , \62666 , \62674 );
xor \U$62299 ( \62676 , \62661 , \62675 );
xor \U$62300 ( \62677 , \62653 , \62676 );
xor \U$62301 ( \62678 , \62602 , \62677 );
xor \U$62302 ( \62679 , \62578 , \62678 );
xor \U$62303 ( \62680 , \62562 , \62679 );
not \U$62304 ( \62681 , \62680 );
and \U$62305 ( \62682 , \62546 , \62681 );
and \U$62306 ( \62683 , \62545 , \62680 );
nor \U$62307 ( \62684 , \62682 , \62683 );
not \U$62308 ( \62685 , \62684 );
and \U$62309 ( \62686 , \62534 , \62685 );
and \U$62310 ( \62687 , \62533 , \62684 );
nor \U$62311 ( \62688 , \62686 , \62687 );
xor \U$62312 ( \62689 , \62476 , \62487 );
and \U$62313 ( \62690 , \62689 , \62492 );
and \U$62314 ( \62691 , \62476 , \62487 );
nor \U$62315 ( \62692 , \62690 , \62691 );
xnor \U$62316 ( \62693 , \62688 , \62692 );
or \U$62317 ( \62694 , \62504 , \62693 );
or \U$62318 ( \62695 , \62692 , \62688 );
nand \U$62319 ( \62696 , \62694 , \62695 );
xor \U$62320 ( \62697 , \62550 , \62554 );
xor \U$62321 ( \62698 , \62697 , \62561 );
and \U$62322 ( \62699 , \62578 , \62698 );
xor \U$62323 ( \62700 , \62550 , \62554 );
xor \U$62324 ( \62701 , \62700 , \62561 );
and \U$62325 ( \62702 , \62678 , \62701 );
and \U$62326 ( \62703 , \62578 , \62678 );
or \U$62327 ( \62704 , \62699 , \62702 , \62703 );
or \U$62328 ( \62705 , \62513 , \62520 );
not \U$62329 ( \62706 , \62520 );
not \U$62330 ( \62707 , \62513 );
or \U$62331 ( \62708 , \62706 , \62707 );
nand \U$62332 ( \62709 , \62708 , \62508 );
nand \U$62333 ( \62710 , \62705 , \62709 );
xor \U$62334 ( \62711 , \62704 , \62710 );
xor \U$62335 ( \62712 , \62586 , \62594 );
and \U$62336 ( \62713 , \62712 , \62601 );
and \U$62337 ( \62714 , \62586 , \62594 );
or \U$62338 ( \62715 , \62713 , \62714 );
xor \U$62339 ( \62716 , \62566 , \62572 );
and \U$62340 ( \62717 , \62716 , \62577 );
and \U$62341 ( \62718 , \62566 , \62572 );
or \U$62342 ( \62719 , \62717 , \62718 );
xor \U$62343 ( \62720 , \62715 , \62719 );
xor \U$62344 ( \62721 , \62655 , \62657 );
xor \U$62345 ( \62722 , \62721 , \62660 );
and \U$62346 ( \62723 , \62666 , \62722 );
xor \U$62347 ( \62724 , \62655 , \62657 );
xor \U$62348 ( \62725 , \62724 , \62660 );
and \U$62349 ( \62726 , \62674 , \62725 );
and \U$62350 ( \62727 , \62666 , \62674 );
or \U$62351 ( \62728 , \62723 , \62726 , \62727 );
xor \U$62352 ( \62729 , \62720 , \62728 );
xor \U$62353 ( \62730 , \62606 , \62613 );
and \U$62354 ( \62731 , \62730 , \62618 );
and \U$62355 ( \62732 , \62606 , \62613 );
or \U$62356 ( \62733 , \62731 , \62732 );
xor \U$62357 ( \62734 , \62623 , \62627 );
and \U$62358 ( \62735 , \62734 , \62632 );
and \U$62359 ( \62736 , \62623 , \62627 );
or \U$62360 ( \62737 , \62735 , \62736 );
xor \U$62361 ( \62738 , \62733 , \62737 );
xor \U$62362 ( \62739 , \62637 , \62643 );
and \U$62363 ( \62740 , \62739 , \62650 );
and \U$62364 ( \62741 , \62637 , \62643 );
or \U$62365 ( \62742 , \62740 , \62741 );
xor \U$62366 ( \62743 , \62738 , \62742 );
xor \U$62367 ( \62744 , \62729 , \62743 );
xor \U$62368 ( \62745 , \53237 , \53262 );
xor \U$62369 ( \62746 , \62745 , \53265 );
xor \U$62370 ( \62747 , \53155 , \53180 );
xor \U$62371 ( \62748 , \62747 , \53206 );
xor \U$62372 ( \62749 , \53076 , \53101 );
xor \U$62373 ( \62750 , \62749 , \53127 );
xor \U$62374 ( \62751 , \62748 , \62750 );
xor \U$62375 ( \62752 , \62746 , \62751 );
xor \U$62376 ( \62753 , \62606 , \62613 );
xor \U$62377 ( \62754 , \62753 , \62618 );
and \U$62378 ( \62755 , \62633 , \62754 );
xor \U$62379 ( \62756 , \62606 , \62613 );
xor \U$62380 ( \62757 , \62756 , \62618 );
and \U$62381 ( \62758 , \62651 , \62757 );
and \U$62382 ( \62759 , \62633 , \62651 );
or \U$62383 ( \62760 , \62755 , \62758 , \62759 );
xor \U$62384 ( \62761 , \62752 , \62760 );
not \U$62385 ( \62762 , \53324 );
xor \U$62386 ( \62763 , \53332 , \53327 );
not \U$62387 ( \62764 , \62763 );
or \U$62388 ( \62765 , \62762 , \62764 );
or \U$62389 ( \62766 , \62763 , \53324 );
nand \U$62390 ( \62767 , \62765 , \62766 );
not \U$62391 ( \62768 , \53309 );
not \U$62392 ( \62769 , \53312 );
or \U$62393 ( \62770 , \62768 , \62769 );
or \U$62394 ( \62771 , \53312 , \53309 );
nand \U$62395 ( \62772 , \62770 , \62771 );
xor \U$62396 ( \62773 , \62767 , \62772 );
not \U$62397 ( \62774 , \53284 );
xor \U$62398 ( \62775 , \53297 , \53273 );
not \U$62399 ( \62776 , \62775 );
or \U$62400 ( \62777 , \62774 , \62776 );
or \U$62401 ( \62778 , \62775 , \53284 );
nand \U$62402 ( \62779 , \62777 , \62778 );
xor \U$62403 ( \62780 , \62773 , \62779 );
xor \U$62404 ( \62781 , \62761 , \62780 );
xor \U$62405 ( \62782 , \62744 , \62781 );
xor \U$62406 ( \62783 , \62711 , \62782 );
xor \U$62407 ( \62784 , \62550 , \62554 );
and \U$62408 ( \62785 , \62784 , \62561 );
and \U$62409 ( \62786 , \62550 , \62554 );
or \U$62410 ( \62787 , \62785 , \62786 );
xor \U$62411 ( \62788 , \53218 , \53225 );
xor \U$62412 ( \62789 , \62788 , \53234 );
and \U$62413 ( \62790 , \62670 , \62789 );
xor \U$62414 ( \62791 , \53218 , \53225 );
xor \U$62415 ( \62792 , \62791 , \53234 );
and \U$62416 ( \62793 , \62672 , \62792 );
and \U$62417 ( \62794 , \62670 , \62672 );
or \U$62418 ( \62795 , \62790 , \62793 , \62794 );
and \U$62419 ( \62796 , \62663 , \62665 );
xor \U$62420 ( \62797 , \62795 , \62796 );
xor \U$62421 ( \62798 , \62655 , \62657 );
and \U$62422 ( \62799 , \62798 , \62660 );
and \U$62423 ( \62800 , \62655 , \62657 );
or \U$62424 ( \62801 , \62799 , \62800 );
xor \U$62425 ( \62802 , \62797 , \62801 );
xor \U$62426 ( \62803 , \62787 , \62802 );
xor \U$62427 ( \62804 , \62586 , \62594 );
xor \U$62428 ( \62805 , \62804 , \62601 );
and \U$62429 ( \62806 , \62653 , \62805 );
xor \U$62430 ( \62807 , \62586 , \62594 );
xor \U$62431 ( \62808 , \62807 , \62601 );
and \U$62432 ( \62809 , \62676 , \62808 );
and \U$62433 ( \62810 , \62653 , \62676 );
or \U$62434 ( \62811 , \62806 , \62809 , \62810 );
xor \U$62435 ( \62812 , \62803 , \62811 );
xor \U$62436 ( \62813 , \62783 , \62812 );
or \U$62437 ( \62814 , \62544 , \62538 );
not \U$62438 ( \62815 , \62538 );
not \U$62439 ( \62816 , \62544 );
or \U$62440 ( \62817 , \62815 , \62816 );
nand \U$62441 ( \62818 , \62817 , \62680 );
nand \U$62442 ( \62819 , \62814 , \62818 );
xor \U$62443 ( \62820 , \62813 , \62819 );
or \U$62444 ( \62821 , \62684 , \62524 );
not \U$62445 ( \62822 , \62524 );
not \U$62446 ( \62823 , \62684 );
or \U$62447 ( \62824 , \62822 , \62823 );
nand \U$62448 ( \62825 , \62824 , \62529 );
nand \U$62449 ( \62826 , \62821 , \62825 );
xor \U$62450 ( \62827 , \62820 , \62826 );
and \U$62451 ( \62828 , \62696 , \62827 );
and \U$62452 ( \62829 , \62826 , \62820 );
nor \U$62453 ( \62830 , \62828 , \62829 );
xor \U$62454 ( \62831 , \62783 , \62812 );
and \U$62455 ( \62832 , \62831 , \62819 );
and \U$62456 ( \62833 , \62783 , \62812 );
nor \U$62457 ( \62834 , \62832 , \62833 );
xor \U$62458 ( \62835 , \62704 , \62710 );
and \U$62459 ( \62836 , \62835 , \62782 );
and \U$62460 ( \62837 , \62704 , \62710 );
or \U$62461 ( \62838 , \62836 , \62837 );
not \U$62462 ( \62839 , \62838 );
xor \U$62463 ( \62840 , \62715 , \62719 );
and \U$62464 ( \62841 , \62840 , \62728 );
and \U$62465 ( \62842 , \62715 , \62719 );
or \U$62466 ( \62843 , \62841 , \62842 );
not \U$62467 ( \62844 , \62843 );
xor \U$62468 ( \62845 , \62752 , \62760 );
and \U$62469 ( \62846 , \62845 , \62780 );
and \U$62470 ( \62847 , \62752 , \62760 );
nor \U$62471 ( \62848 , \62846 , \62847 );
not \U$62472 ( \62849 , \62848 );
or \U$62473 ( \62850 , \62844 , \62849 );
or \U$62474 ( \62851 , \62848 , \62843 );
nand \U$62475 ( \62852 , \62850 , \62851 );
not \U$62476 ( \62853 , \62852 );
xor \U$62477 ( \62854 , \53299 , \53313 );
xor \U$62478 ( \62855 , \62854 , \53334 );
not \U$62479 ( \62856 , \62855 );
and \U$62480 ( \62857 , \62853 , \62856 );
and \U$62481 ( \62858 , \62852 , \62855 );
nor \U$62482 ( \62859 , \62857 , \62858 );
not \U$62483 ( \62860 , \62859 );
and \U$62484 ( \62861 , \62839 , \62860 );
and \U$62485 ( \62862 , \62838 , \62859 );
nor \U$62486 ( \62863 , \62861 , \62862 );
not \U$62487 ( \62864 , \62863 );
xor \U$62488 ( \62865 , \62787 , \62802 );
and \U$62489 ( \62866 , \62865 , \62811 );
and \U$62490 ( \62867 , \62787 , \62802 );
or \U$62491 ( \62868 , \62866 , \62867 );
xor \U$62492 ( \62869 , \62729 , \62743 );
and \U$62493 ( \62870 , \62869 , \62781 );
and \U$62494 ( \62871 , \62729 , \62743 );
or \U$62495 ( \62872 , \62870 , \62871 );
xor \U$62496 ( \62873 , \62868 , \62872 );
xor \U$62497 ( \62874 , \62795 , \62796 );
and \U$62498 ( \62875 , \62874 , \62801 );
and \U$62499 ( \62876 , \62795 , \62796 );
or \U$62500 ( \62877 , \62875 , \62876 );
xor \U$62501 ( \62878 , \62733 , \62737 );
and \U$62502 ( \62879 , \62878 , \62742 );
and \U$62503 ( \62880 , \62733 , \62737 );
or \U$62504 ( \62881 , \62879 , \62880 );
xor \U$62505 ( \62882 , \62877 , \62881 );
xor \U$62506 ( \62883 , \62767 , \62772 );
and \U$62507 ( \62884 , \62883 , \62779 );
and \U$62508 ( \62885 , \62767 , \62772 );
or \U$62509 ( \62886 , \62884 , \62885 );
xor \U$62510 ( \62887 , \62882 , \62886 );
xor \U$62511 ( \62888 , \53130 , \53209 );
xor \U$62512 ( \62889 , \62888 , \53268 );
xor \U$62513 ( \62890 , \53033 , \53035 );
xor \U$62514 ( \62891 , \62890 , \53038 );
xor \U$62515 ( \62892 , \53237 , \53262 );
xor \U$62516 ( \62893 , \62892 , \53265 );
and \U$62517 ( \62894 , \62748 , \62893 );
xor \U$62518 ( \62895 , \53237 , \53262 );
xor \U$62519 ( \62896 , \62895 , \53265 );
and \U$62520 ( \62897 , \62750 , \62896 );
and \U$62521 ( \62898 , \62748 , \62750 );
or \U$62522 ( \62899 , \62894 , \62897 , \62898 );
not \U$62523 ( \62900 , \53348 );
xor \U$62524 ( \62901 , \53359 , \53372 );
not \U$62525 ( \62902 , \62901 );
or \U$62526 ( \62903 , \62900 , \62902 );
or \U$62527 ( \62904 , \62901 , \53348 );
nand \U$62528 ( \62905 , \62903 , \62904 );
xor \U$62529 ( \62906 , \62899 , \62905 );
xor \U$62530 ( \62907 , \62891 , \62906 );
xor \U$62531 ( \62908 , \62889 , \62907 );
xor \U$62532 ( \62909 , \62887 , \62908 );
xor \U$62533 ( \62910 , \62873 , \62909 );
not \U$62534 ( \62911 , \62910 );
and \U$62535 ( \62912 , \62864 , \62911 );
and \U$62536 ( \62913 , \62863 , \62910 );
nor \U$62537 ( \62914 , \62912 , \62913 );
xnor \U$62538 ( \62915 , \62834 , \62914 );
or \U$62539 ( \62916 , \62830 , \62915 );
or \U$62540 ( \62917 , \62834 , \62914 );
nand \U$62541 ( \62918 , \62916 , \62917 );
not \U$62542 ( \62919 , \62910 );
or \U$62543 ( \62920 , \62919 , \62859 );
not \U$62544 ( \62921 , \62859 );
not \U$62545 ( \62922 , \62919 );
or \U$62546 ( \62923 , \62921 , \62922 );
nand \U$62547 ( \62924 , \62923 , \62838 );
nand \U$62548 ( \62925 , \62920 , \62924 );
xor \U$62549 ( \62926 , \53271 , \53337 );
xor \U$62550 ( \62927 , \62926 , \53374 );
not \U$62551 ( \62928 , \62927 );
xor \U$62552 ( \62929 , \53033 , \53035 );
xor \U$62553 ( \62930 , \62929 , \53038 );
and \U$62554 ( \62931 , \62899 , \62930 );
xor \U$62555 ( \62932 , \53033 , \53035 );
xor \U$62556 ( \62933 , \62932 , \53038 );
and \U$62557 ( \62934 , \62905 , \62933 );
and \U$62558 ( \62935 , \62899 , \62905 );
or \U$62559 ( \62936 , \62931 , \62934 , \62935 );
xor \U$62560 ( \62937 , \62877 , \62881 );
and \U$62561 ( \62938 , \62937 , \62886 );
and \U$62562 ( \62939 , \62877 , \62881 );
or \U$62563 ( \62940 , \62938 , \62939 );
xor \U$62564 ( \62941 , \62936 , \62940 );
xor \U$62565 ( \62942 , \52628 , \52648 );
xor \U$62566 ( \62943 , \62942 , \52669 );
xor \U$62567 ( \62944 , \53380 , \53387 );
xor \U$62568 ( \62945 , \62943 , \62944 );
xor \U$62569 ( \62946 , \62941 , \62945 );
not \U$62570 ( \62947 , \62946 );
or \U$62571 ( \62948 , \62928 , \62947 );
or \U$62572 ( \62949 , \62946 , \62927 );
nand \U$62573 ( \62950 , \62948 , \62949 );
xor \U$62574 ( \62951 , \62868 , \62872 );
and \U$62575 ( \62952 , \62951 , \62909 );
and \U$62576 ( \62953 , \62868 , \62872 );
or \U$62577 ( \62954 , \62952 , \62953 );
xor \U$62578 ( \62955 , \62950 , \62954 );
not \U$62579 ( \62956 , \62843 );
or \U$62580 ( \62957 , \62956 , \62855 );
and \U$62581 ( \62958 , \62956 , \62855 );
nor \U$62582 ( \62959 , \62958 , \62848 );
not \U$62583 ( \62960 , \62959 );
nand \U$62584 ( \62961 , \62957 , \62960 );
xor \U$62585 ( \62962 , \53041 , \53043 );
xor \U$62586 ( \62963 , \62962 , \53048 );
xor \U$62587 ( \62964 , \62961 , \62963 );
xor \U$62588 ( \62965 , \62877 , \62881 );
xor \U$62589 ( \62966 , \62965 , \62886 );
and \U$62590 ( \62967 , \62889 , \62966 );
xor \U$62591 ( \62968 , \62877 , \62881 );
xor \U$62592 ( \62969 , \62968 , \62886 );
and \U$62593 ( \62970 , \62907 , \62969 );
and \U$62594 ( \62971 , \62889 , \62907 );
or \U$62595 ( \62972 , \62967 , \62970 , \62971 );
xor \U$62596 ( \62973 , \62964 , \62972 );
xor \U$62597 ( \62974 , \62955 , \62973 );
xor \U$62598 ( \62975 , \62925 , \62974 );
and \U$62599 ( \62976 , \62918 , \62975 );
and \U$62600 ( \62977 , \62925 , \62974 );
nor \U$62601 ( \62978 , \62976 , \62977 );
xor \U$62602 ( \62979 , \62961 , \62963 );
and \U$62603 ( \62980 , \62979 , \62972 );
and \U$62604 ( \62981 , \62961 , \62963 );
or \U$62605 ( \62982 , \62980 , \62981 );
not \U$62606 ( \62983 , \62982 );
not \U$62607 ( \62984 , \62927 );
nand \U$62608 ( \62985 , \62984 , \62946 );
not \U$62609 ( \62986 , \62985 );
and \U$62610 ( \62987 , \62983 , \62986 );
and \U$62611 ( \62988 , \62982 , \62985 );
nor \U$62612 ( \62989 , \62987 , \62988 );
not \U$62613 ( \62990 , \62989 );
xor \U$62614 ( \62991 , \53051 , \53377 );
xor \U$62615 ( \62992 , \62991 , \53392 );
xor \U$62616 ( \62993 , \62936 , \62940 );
and \U$62617 ( \62994 , \62993 , \62945 );
and \U$62618 ( \62995 , \62936 , \62940 );
or \U$62619 ( \62996 , \62994 , \62995 );
xor \U$62620 ( \62997 , \52672 , \52914 );
xor \U$62621 ( \62998 , \62997 , \52929 );
xor \U$62622 ( \62999 , \53396 , \53403 );
xor \U$62623 ( \63000 , \62998 , \62999 );
xor \U$62624 ( \63001 , \62996 , \63000 );
xor \U$62625 ( \63002 , \62992 , \63001 );
not \U$62626 ( \63003 , \63002 );
and \U$62627 ( \63004 , \62990 , \63003 );
and \U$62628 ( \63005 , \62989 , \63002 );
nor \U$62629 ( \63006 , \63004 , \63005 );
xor \U$62630 ( \63007 , \62950 , \62954 );
and \U$62631 ( \63008 , \63007 , \62973 );
and \U$62632 ( \63009 , \62950 , \62954 );
nor \U$62633 ( \63010 , \63008 , \63009 );
xnor \U$62634 ( \63011 , \63006 , \63010 );
or \U$62635 ( \63012 , \62978 , \63011 );
or \U$62636 ( \63013 , \63010 , \63006 );
nand \U$62637 ( \63014 , \63012 , \63013 );
not \U$62638 ( \63015 , \63002 );
or \U$62639 ( \63016 , \63015 , \62985 );
not \U$62640 ( \63017 , \62985 );
not \U$62641 ( \63018 , \63015 );
or \U$62642 ( \63019 , \63017 , \63018 );
nand \U$62643 ( \63020 , \63019 , \62982 );
nand \U$62644 ( \63021 , \63016 , \63020 );
xor \U$62645 ( \63022 , \53395 , \53408 );
xor \U$62646 ( \63023 , \63022 , \53413 );
xor \U$62647 ( \63024 , \52932 , \52937 );
xor \U$62648 ( \63025 , \63024 , \52964 );
xor \U$62649 ( \63026 , \63023 , \63025 );
xor \U$62650 ( \63027 , \53051 , \53377 );
xor \U$62651 ( \63028 , \63027 , \53392 );
and \U$62652 ( \63029 , \62996 , \63028 );
xor \U$62653 ( \63030 , \53051 , \53377 );
xor \U$62654 ( \63031 , \63030 , \53392 );
and \U$62655 ( \63032 , \63000 , \63031 );
and \U$62656 ( \63033 , \62996 , \63000 );
or \U$62657 ( \63034 , \63029 , \63032 , \63033 );
xor \U$62658 ( \63035 , \63026 , \63034 );
xor \U$62659 ( \63036 , \63021 , \63035 );
and \U$62660 ( \63037 , \63014 , \63036 );
and \U$62661 ( \63038 , \63021 , \63035 );
nor \U$62662 ( \63039 , \63037 , \63038 );
xor \U$62663 ( \63040 , \63023 , \63025 );
and \U$62664 ( \63041 , \63040 , \63034 );
and \U$62665 ( \63042 , \63023 , \63025 );
nor \U$62666 ( \63043 , \63041 , \63042 );
xnor \U$62667 ( \63044 , \53416 , \53028 );
not \U$62668 ( \63045 , \63044 );
not \U$62669 ( \63046 , \53025 );
and \U$62670 ( \63047 , \63045 , \63046 );
and \U$62671 ( \63048 , \63044 , \53025 );
nor \U$62672 ( \63049 , \63047 , \63048 );
xnor \U$62673 ( \63050 , \63043 , \63049 );
or \U$62674 ( \63051 , \63039 , \63050 );
or \U$62675 ( \63052 , \63043 , \63049 );
nand \U$62676 ( \63053 , \63051 , \63052 );
and \U$62677 ( \63054 , \53420 , \63053 );
nor \U$62678 ( \63055 , \53419 , \63054 );
or \U$62679 ( \63056 , \53015 , \63055 );
nand \U$62680 ( \63057 , \53014 , \63056 );
not \U$62681 ( \63058 , \52583 );
nor \U$62682 ( \63059 , \63058 , \52987 );
not \U$62683 ( \63060 , \52575 );
not \U$62684 ( \63061 , \52578 );
or \U$62685 ( \63062 , \63060 , \63061 );
or \U$62686 ( \63063 , \52578 , \52575 );
nand \U$62687 ( \63064 , \63062 , \63063 );
xor \U$62688 ( \63065 , \63059 , \63064 );
and \U$62689 ( \63066 , \63057 , \63065 );
and \U$62690 ( \63067 , \63059 , \63064 );
nor \U$62691 ( \63068 , \63066 , \63067 );
or \U$62692 ( \63069 , \52581 , \63068 );
nand \U$62693 ( \63070 , \52580 , \63069 );
not \U$62694 ( \63071 , \52201 );
nor \U$62695 ( \63072 , \63071 , \51829 );
xor \U$62696 ( \63073 , \50972 , \50984 );
xor \U$62697 ( \63074 , \63073 , \50989 );
xor \U$62698 ( \63075 , \50175 , \50523 );
xor \U$62699 ( \63076 , \63075 , \50566 );
or \U$62700 ( \63077 , \51388 , \51403 );
not \U$62701 ( \63078 , \51403 );
not \U$62702 ( \63079 , \51388 );
or \U$62703 ( \63080 , \63078 , \63079 );
nand \U$62704 ( \63081 , \63080 , \51375 );
nand \U$62705 ( \63082 , \63077 , \63081 );
xor \U$62706 ( \63083 , \63076 , \63082 );
xor \U$62707 ( \63084 , \50974 , \50976 );
xor \U$62708 ( \63085 , \63084 , \50981 );
and \U$62709 ( \63086 , \51821 , \63085 );
xor \U$62710 ( \63087 , \50974 , \50976 );
xor \U$62711 ( \63088 , \63087 , \50981 );
and \U$62712 ( \63089 , \51823 , \63088 );
and \U$62713 ( \63090 , \51821 , \51823 );
or \U$62714 ( \63091 , \63086 , \63089 , \63090 );
xor \U$62715 ( \63092 , \63083 , \63091 );
xor \U$62716 ( \63093 , \63074 , \63092 );
not \U$62717 ( \63094 , \51825 );
or \U$62718 ( \63095 , \63094 , \51407 );
not \U$62719 ( \63096 , \51407 );
not \U$62720 ( \63097 , \63094 );
or \U$62721 ( \63098 , \63096 , \63097 );
nand \U$62722 ( \63099 , \63098 , \51812 );
nand \U$62723 ( \63100 , \63095 , \63099 );
xor \U$62724 ( \63101 , \63093 , \63100 );
xor \U$62725 ( \63102 , \63072 , \63101 );
and \U$62726 ( \63103 , \63070 , \63102 );
and \U$62727 ( \63104 , \63072 , \63101 );
nor \U$62728 ( \63105 , \63103 , \63104 );
xor \U$62729 ( \63106 , \50610 , \50992 );
xor \U$62730 ( \63107 , \63106 , \50995 );
not \U$62731 ( \63108 , \63107 );
xor \U$62732 ( \63109 , \63076 , \63082 );
and \U$62733 ( \63110 , \63109 , \63091 );
and \U$62734 ( \63111 , \63076 , \63082 );
nor \U$62735 ( \63112 , \63110 , \63111 );
not \U$62736 ( \63113 , \63112 );
and \U$62737 ( \63114 , \63108 , \63113 );
and \U$62738 ( \63115 , \63107 , \63112 );
nor \U$62739 ( \63116 , \63114 , \63115 );
xor \U$62740 ( \63117 , \63074 , \63092 );
and \U$62741 ( \63118 , \63117 , \63100 );
and \U$62742 ( \63119 , \63074 , \63092 );
nor \U$62743 ( \63120 , \63118 , \63119 );
xnor \U$62744 ( \63121 , \63116 , \63120 );
or \U$62745 ( \63122 , \63105 , \63121 );
or \U$62746 ( \63123 , \63116 , \63120 );
nand \U$62747 ( \63124 , \63122 , \63123 );
not \U$62748 ( \63125 , \63107 );
nor \U$62749 ( \63126 , \63125 , \63112 );
not \U$62750 ( \63127 , \50998 );
not \U$62751 ( \63128 , \51003 );
or \U$62752 ( \63129 , \63127 , \63128 );
or \U$62753 ( \63130 , \51003 , \50998 );
nand \U$62754 ( \63131 , \63129 , \63130 );
xor \U$62755 ( \63132 , \63126 , \63131 );
and \U$62756 ( \63133 , \63124 , \63132 );
and \U$62757 ( \63134 , \63126 , \63131 );
nor \U$62758 ( \63135 , \63133 , \63134 );
or \U$62759 ( \63136 , \51006 , \63135 );
nand \U$62760 ( \63137 , \51005 , \63136 );
and \U$62761 ( \63138 , \50602 , \63137 );
nor \U$62762 ( \63139 , \50601 , \63138 );
not \U$62763 ( \63140 , \50593 );
nand \U$62764 ( \63141 , \63140 , \50596 );
xor \U$62765 ( \63142 , \49724 , \49729 );
xor \U$62766 ( \63143 , \63142 , \49736 );
and \U$62767 ( \63144 , \63141 , \63143 );
not \U$62768 ( \63145 , \63141 );
not \U$62769 ( \63146 , \63143 );
and \U$62770 ( \63147 , \63145 , \63146 );
nor \U$62771 ( \63148 , \63144 , \63147 );
or \U$62772 ( \63149 , \63139 , \63148 );
or \U$62773 ( \63150 , \63141 , \63146 );
nand \U$62774 ( \63151 , \63149 , \63150 );
and \U$62775 ( \63152 , \49741 , \63151 );
nor \U$62776 ( \63153 , \49740 , \63152 );
not \U$62777 ( \63154 , \48879 );
not \U$62778 ( \63155 , \48894 );
and \U$62779 ( \63156 , \63154 , \63155 );
and \U$62780 ( \63157 , \48879 , \48894 );
nor \U$62781 ( \63158 , \63157 , \49317 );
nor \U$62782 ( \63159 , \63156 , \63158 );
or \U$62783 ( \63160 , \48875 , \48856 );
not \U$62784 ( \63161 , \48875 );
not \U$62785 ( \63162 , \48856 );
or \U$62786 ( \63163 , \63161 , \63162 );
nand \U$62787 ( \63164 , \63163 , \48779 );
nand \U$62788 ( \63165 , \63160 , \63164 );
or \U$62789 ( \63166 , \48865 , \48863 );
not \U$62790 ( \63167 , \48863 );
not \U$62791 ( \63168 , \48865 );
or \U$62792 ( \63169 , \63167 , \63168 );
nand \U$62793 ( \63170 , \63169 , \48871 );
nand \U$62794 ( \63171 , \63166 , \63170 );
xor \U$62795 ( \63172 , \46581 , \46591 );
xor \U$62796 ( \63173 , \63172 , \46596 );
xor \U$62797 ( \63174 , \47492 , \47499 );
xor \U$62798 ( \63175 , \63173 , \63174 );
xor \U$62799 ( \63176 , \63171 , \63175 );
or \U$62800 ( \63177 , \48837 , \48852 );
not \U$62801 ( \63178 , \48852 );
not \U$62802 ( \63179 , \48837 );
or \U$62803 ( \63180 , \63178 , \63179 );
nand \U$62804 ( \63181 , \63180 , \48824 );
nand \U$62805 ( \63182 , \63177 , \63181 );
xor \U$62806 ( \63183 , \63176 , \63182 );
xnor \U$62807 ( \63184 , \63165 , \63183 );
not \U$62808 ( \63185 , \63184 );
xor \U$62809 ( \63186 , \47109 , \47469 );
xor \U$62810 ( \63187 , \63186 , \47484 );
xor \U$62811 ( \63188 , \47553 , \47555 );
xor \U$62812 ( \63189 , \63188 , \48012 );
xor \U$62813 ( \63190 , \63187 , \63189 );
not \U$62814 ( \63191 , \63190 );
and \U$62815 ( \63192 , \63185 , \63191 );
and \U$62816 ( \63193 , \63184 , \63190 );
nor \U$62817 ( \63194 , \63192 , \63193 );
xnor \U$62818 ( \63195 , \63159 , \63194 );
or \U$62819 ( \63196 , \63153 , \63195 );
or \U$62820 ( \63197 , \63159 , \63194 );
nand \U$62821 ( \63198 , \63196 , \63197 );
xnor \U$62822 ( \63199 , \48015 , \47536 );
not \U$62823 ( \63200 , \63199 );
not \U$62824 ( \63201 , \47533 );
and \U$62825 ( \63202 , \63200 , \63201 );
and \U$62826 ( \63203 , \63199 , \47533 );
nor \U$62827 ( \63204 , \63202 , \63203 );
not \U$62828 ( \63205 , \63204 );
and \U$62829 ( \63206 , \63187 , \63189 );
xor \U$62830 ( \63207 , \63171 , \63175 );
and \U$62831 ( \63208 , \63207 , \63182 );
and \U$62832 ( \63209 , \63171 , \63175 );
or \U$62833 ( \63210 , \63208 , \63209 );
xor \U$62834 ( \63211 , \63206 , \63210 );
not \U$62835 ( \63212 , \63211 );
or \U$62836 ( \63213 , \63205 , \63212 );
or \U$62837 ( \63214 , \63211 , \63204 );
nand \U$62838 ( \63215 , \63213 , \63214 );
not \U$62839 ( \63216 , \63190 );
not \U$62840 ( \63217 , \63183 );
or \U$62841 ( \63218 , \63216 , \63217 );
or \U$62842 ( \63219 , \63183 , \63190 );
nand \U$62843 ( \63220 , \63219 , \63165 );
nand \U$62844 ( \63221 , \63218 , \63220 );
xor \U$62845 ( \63222 , \63215 , \63221 );
and \U$62846 ( \63223 , \63198 , \63222 );
and \U$62847 ( \63224 , \63221 , \63215 );
nor \U$62848 ( \63225 , \63223 , \63224 );
and \U$62849 ( \63226 , \63210 , \63206 );
not \U$62850 ( \63227 , \63210 );
not \U$62851 ( \63228 , \63206 );
and \U$62852 ( \63229 , \63227 , \63228 );
nor \U$62853 ( \63230 , \63229 , \63204 );
nor \U$62854 ( \63231 , \63226 , \63230 );
xnor \U$62855 ( \63232 , \47529 , \48017 );
not \U$62856 ( \63233 , \63232 );
not \U$62857 ( \63234 , \47526 );
and \U$62858 ( \63235 , \63233 , \63234 );
and \U$62859 ( \63236 , \63232 , \47526 );
nor \U$62860 ( \63237 , \63235 , \63236 );
xnor \U$62861 ( \63238 , \63231 , \63237 );
or \U$62862 ( \63239 , \63225 , \63238 );
or \U$62863 ( \63240 , \63231 , \63237 );
nand \U$62864 ( \63241 , \63239 , \63240 );
and \U$62865 ( \63242 , \48021 , \63241 );
nor \U$62866 ( \63243 , \48020 , \63242 );
xnor \U$62867 ( \63244 , \47518 , \47521 );
or \U$62868 ( \63245 , \63243 , \63244 );
nand \U$62869 ( \63246 , \47523 , \63245 );
and \U$62870 ( \63247 , \47044 , \63246 );
nor \U$62871 ( \63248 , \47043 , \63247 );
xnor \U$62872 ( \63249 , \46548 , \46563 );
or \U$62873 ( \63250 , \63248 , \63249 );
nand \U$62874 ( \63251 , \46565 , \63250 );
not \U$62875 ( \63252 , \45663 );
not \U$62876 ( \63253 , \45666 );
or \U$62877 ( \63254 , \63252 , \63253 );
or \U$62878 ( \63255 , \45666 , \45663 );
nand \U$62879 ( \63256 , \63254 , \63255 );
xor \U$62880 ( \63257 , \46557 , \46559 );
and \U$62881 ( \63258 , \63257 , \46562 );
and \U$62882 ( \63259 , \46557 , \46559 );
or \U$62883 ( \63260 , \63258 , \63259 );
xor \U$62884 ( \63261 , \63256 , \63260 );
and \U$62885 ( \63262 , \63251 , \63261 );
and \U$62886 ( \63263 , \63256 , \63260 );
nor \U$62887 ( \63264 , \63262 , \63263 );
or \U$62888 ( \63265 , \45673 , \63264 );
nand \U$62889 ( \63266 , \45668 , \63265 );
and \U$62890 ( \63267 , \45251 , \63266 );
nor \U$62891 ( \63268 , \45250 , \63267 );
xnor \U$62892 ( \63269 , \44838 , \44420 );
or \U$62893 ( \63270 , \63268 , \63269 );
nand \U$62894 ( \63271 , \44840 , \63270 );
and \U$62895 ( \63272 , \44419 , \63271 );
nor \U$62896 ( \63273 , \44418 , \63272 );
not \U$62897 ( \63274 , \44015 );
nand \U$62898 ( \63275 , \63274 , \44004 );
not \U$62899 ( \63276 , \43613 );
not \U$62900 ( \63277 , \43610 );
and \U$62901 ( \63278 , \63276 , \63277 );
and \U$62902 ( \63279 , \43613 , \43610 );
nor \U$62903 ( \63280 , \63278 , \63279 );
xnor \U$62904 ( \63281 , \63275 , \63280 );
or \U$62905 ( \63282 , \63273 , \63281 );
or \U$62906 ( \63283 , \63275 , \63280 );
nand \U$62907 ( \63284 , \63282 , \63283 );
and \U$62908 ( \63285 , \43616 , \63284 );
nor \U$62909 ( \63286 , \43615 , \63285 );
or \U$62910 ( \63287 , \43205 , \63286 );
nand \U$62911 ( \63288 , \43204 , \63287 );
and \U$62912 ( \63289 , \42812 , \63288 );
nor \U$62913 ( \63290 , \42811 , \63289 );
xnor \U$62914 ( \63291 , \42421 , \42429 );
or \U$62915 ( \63292 , \63290 , \63291 );
nand \U$62916 ( \63293 , \42431 , \63292 );
not \U$62917 ( \63294 , \41649 );
not \U$62918 ( \63295 , \41288 );
or \U$62919 ( \63296 , \63294 , \63295 );
or \U$62920 ( \63297 , \41288 , \41649 );
nand \U$62921 ( \63298 , \63296 , \63297 );
and \U$62922 ( \63299 , \42426 , \42428 );
xor \U$62923 ( \63300 , \63298 , \63299 );
and \U$62924 ( \63301 , \63293 , \63300 );
and \U$62925 ( \63302 , \63299 , \63298 );
nor \U$62926 ( \63303 , \63301 , \63302 );
or \U$62927 ( \63304 , \41652 , \63303 );
nand \U$62928 ( \63305 , \41651 , \63304 );
not \U$62929 ( \63306 , \41274 );
nor \U$62930 ( \63307 , \63306 , \40914 );
not \U$62931 ( \63308 , \40898 );
not \U$62932 ( \63309 , \40909 );
or \U$62933 ( \63310 , \63308 , \63309 );
or \U$62934 ( \63311 , \40909 , \40898 );
nand \U$62935 ( \63312 , \63310 , \63311 );
xor \U$62936 ( \63313 , \63307 , \63312 );
and \U$62937 ( \63314 , \63305 , \63313 );
and \U$62938 ( \63315 , \63307 , \63312 );
nor \U$62939 ( \63316 , \63314 , \63315 );
or \U$62940 ( \63317 , \40912 , \63316 );
nand \U$62941 ( \63318 , \40911 , \63317 );
and \U$62942 ( \63319 , \40516 , \63318 );
nor \U$62943 ( \63320 , \40515 , \63319 );
or \U$62944 ( \63321 , \40130 , \63320 );
nand \U$62945 ( \63322 , \40125 , \63321 );
and \U$62946 ( \63323 , \39763 , \63322 );
nor \U$62947 ( \63324 , \39762 , \63323 );
or \U$62948 ( \63325 , \39406 , \63324 );
nand \U$62949 ( \63326 , \39401 , \63325 );
xor \U$62950 ( \63327 , \38174 , \38384 );
and \U$62951 ( \63328 , \63327 , \38481 );
and \U$62952 ( \63329 , \38174 , \38384 );
or \U$62953 ( \63330 , \63328 , \63329 );
xor \U$62954 ( \63331 , \38178 , \38182 );
and \U$62955 ( \63332 , \63331 , \38187 );
and \U$62956 ( \63333 , \38178 , \38182 );
or \U$62957 ( \63334 , \63332 , \63333 );
xor \U$62958 ( \63335 , \38205 , \38213 );
xor \U$62959 ( \63336 , \63335 , \38221 );
and \U$62960 ( \63337 , \38238 , \63336 );
xor \U$62961 ( \63338 , \38205 , \38213 );
xor \U$62962 ( \63339 , \63338 , \38221 );
and \U$62963 ( \63340 , \38262 , \63339 );
and \U$62964 ( \63341 , \38238 , \38262 );
or \U$62965 ( \63342 , \63337 , \63340 , \63341 );
not \U$62966 ( \63343 , \2774 );
and \U$62967 ( \63344 , \3214 , RIae76280_38);
and \U$62968 ( \63345 , RIae76af0_56, \3212 );
nor \U$62969 ( \63346 , \63344 , \63345 );
not \U$62970 ( \63347 , \63346 );
or \U$62971 ( \63348 , \63343 , \63347 );
or \U$62972 ( \63349 , \63346 , \3218 );
nand \U$62973 ( \63350 , \63348 , \63349 );
not \U$62974 ( \63351 , \3089 );
and \U$62975 ( \63352 , \2783 , RIae760a0_34);
and \U$62976 ( \63353 , RIae76370_40, \2781 );
nor \U$62977 ( \63354 , \63352 , \63353 );
not \U$62978 ( \63355 , \63354 );
or \U$62979 ( \63356 , \63351 , \63355 );
or \U$62980 ( \63357 , \63354 , \2789 );
nand \U$62981 ( \63358 , \63356 , \63357 );
xor \U$62982 ( \63359 , \63350 , \63358 );
and \U$62983 ( \63360 , \3730 , RIae76a00_54);
and \U$62984 ( \63361 , RIae76820_50, \3728 );
nor \U$62985 ( \63362 , \63360 , \63361 );
and \U$62986 ( \63363 , \63362 , \3732 );
not \U$62987 ( \63364 , \63362 );
and \U$62988 ( \63365 , \63364 , \3422 );
nor \U$62989 ( \63366 , \63363 , \63365 );
xor \U$62990 ( \63367 , \63359 , \63366 );
xor \U$62991 ( \63368 , \63342 , \63367 );
xor \U$62992 ( \63369 , \38312 , \38319 );
xor \U$62993 ( \63370 , \63369 , \38327 );
and \U$62994 ( \63371 , \38353 , \63370 );
xor \U$62995 ( \63372 , \38312 , \38319 );
xor \U$62996 ( \63373 , \63372 , \38327 );
and \U$62997 ( \63374 , \38377 , \63373 );
and \U$62998 ( \63375 , \38353 , \38377 );
or \U$62999 ( \63376 , \63371 , \63374 , \63375 );
xor \U$63000 ( \63377 , \63368 , \63376 );
xor \U$63001 ( \63378 , \63334 , \63377 );
xor \U$63002 ( \63379 , \38196 , \38197 );
xor \U$63003 ( \63380 , \63379 , \38264 );
and \U$63004 ( \63381 , \38279 , \63380 );
xor \U$63005 ( \63382 , \38196 , \38197 );
xor \U$63006 ( \63383 , \63382 , \38264 );
and \U$63007 ( \63384 , \38381 , \63383 );
and \U$63008 ( \63385 , \38279 , \38381 );
or \U$63009 ( \63386 , \63381 , \63384 , \63385 );
xor \U$63010 ( \63387 , \63378 , \63386 );
xor \U$63011 ( \63388 , \63330 , \63387 );
xor \U$63012 ( \63389 , \38457 , \38471 );
and \U$63013 ( \63390 , \63389 , \38480 );
and \U$63014 ( \63391 , \38457 , \38471 );
or \U$63015 ( \63392 , \63390 , \63391 );
and \U$63016 ( \63393 , \38188 , \38383 );
xor \U$63017 ( \63394 , \63392 , \63393 );
xor \U$63018 ( \63395 , \38246 , \38253 );
and \U$63019 ( \63396 , \63395 , \38261 );
and \U$63020 ( \63397 , \38246 , \38253 );
or \U$63021 ( \63398 , \63396 , \63397 );
xor \U$63022 ( \63399 , \38229 , \5590 );
and \U$63023 ( \63400 , \63399 , \38237 );
and \U$63024 ( \63401 , \38229 , \5590 );
or \U$63025 ( \63402 , \63400 , \63401 );
xor \U$63026 ( \63403 , \63398 , \63402 );
xor \U$63027 ( \63404 , \38205 , \38213 );
and \U$63028 ( \63405 , \63404 , \38221 );
and \U$63029 ( \63406 , \38205 , \38213 );
or \U$63030 ( \63407 , \63405 , \63406 );
xor \U$63031 ( \63408 , \63403 , \63407 );
xor \U$63032 ( \63409 , \38312 , \38319 );
and \U$63033 ( \63410 , \63409 , \38327 );
and \U$63034 ( \63411 , \38312 , \38319 );
or \U$63035 ( \63412 , \63410 , \63411 );
xor \U$63036 ( \63413 , \38335 , \38343 );
and \U$63037 ( \63414 , \63413 , \38352 );
and \U$63038 ( \63415 , \38335 , \38343 );
or \U$63039 ( \63416 , \63414 , \63415 );
xor \U$63040 ( \63417 , \63412 , \63416 );
xor \U$63041 ( \63418 , \38361 , \38368 );
and \U$63042 ( \63419 , \63418 , \38376 );
and \U$63043 ( \63420 , \38361 , \38368 );
or \U$63044 ( \63421 , \63419 , \63420 );
xor \U$63045 ( \63422 , \63417 , \63421 );
xor \U$63046 ( \63423 , \63408 , \63422 );
and \U$63047 ( \63424 , \436 , RIae78710_116);
and \U$63048 ( \63425 , RIae75bf0_24, \434 );
nor \U$63049 ( \63426 , \63424 , \63425 );
not \U$63050 ( \63427 , \63426 );
not \U$63051 ( \63428 , \402 );
and \U$63052 ( \63429 , \63427 , \63428 );
and \U$63053 ( \63430 , \63426 , \400 );
nor \U$63054 ( \63431 , \63429 , \63430 );
not \U$63055 ( \63432 , \63431 );
not \U$63056 ( \63433 , \471 );
and \U$63057 ( \63434 , \514 , RIae75b00_22);
and \U$63058 ( \63435 , RIae75a10_20, \512 );
nor \U$63059 ( \63436 , \63434 , \63435 );
not \U$63060 ( \63437 , \63436 );
or \U$63061 ( \63438 , \63433 , \63437 );
or \U$63062 ( \63439 , \63436 , \469 );
nand \U$63063 ( \63440 , \63438 , \63439 );
not \U$63064 ( \63441 , \63440 );
or \U$63065 ( \63442 , \63432 , \63441 );
or \U$63066 ( \63443 , \63431 , \63440 );
nand \U$63067 ( \63444 , \63442 , \63443 );
not \U$63068 ( \63445 , \63444 );
and \U$63069 ( \63446 , \384 , RIae788f0_120);
and \U$63070 ( \63447 , RIae78800_118, \382 );
nor \U$63071 ( \63448 , \63446 , \63447 );
not \U$63072 ( \63449 , \63448 );
not \U$63073 ( \63450 , \388 );
and \U$63074 ( \63451 , \63449 , \63450 );
and \U$63075 ( \63452 , \63448 , \388 );
nor \U$63076 ( \63453 , \63451 , \63452 );
not \U$63077 ( \63454 , \63453 );
and \U$63078 ( \63455 , \63445 , \63454 );
and \U$63079 ( \63456 , \63444 , \63453 );
nor \U$63080 ( \63457 , \63455 , \63456 );
nand \U$63081 ( \63458 , RIae789e0_122, RIae78b48_125);
or \U$63082 ( \63459 , \63457 , \63458 );
nand \U$63083 ( \63460 , \63458 , \63457 );
nand \U$63084 ( \63461 , \63459 , \63460 );
and \U$63085 ( \63462 , \4247 , RIae76910_52);
and \U$63086 ( \63463 , RIae76be0_58, \4245 );
nor \U$63087 ( \63464 , \63462 , \63463 );
and \U$63088 ( \63465 , \63464 , \3989 );
not \U$63089 ( \63466 , \63464 );
and \U$63090 ( \63467 , \63466 , \4251 );
nor \U$63091 ( \63468 , \63465 , \63467 );
nand \U$63092 ( \63469 , RIae78e18_131, \5399 );
and \U$63093 ( \63470 , \63469 , \5016 );
not \U$63094 ( \63471 , \63469 );
and \U$63095 ( \63472 , \63471 , \5403 );
nor \U$63096 ( \63473 , \63470 , \63472 );
xor \U$63097 ( \63474 , \63468 , \63473 );
and \U$63098 ( \63475 , \4688 , RIae78ad0_124);
and \U$63099 ( \63476 , RIae78d28_129, \4686 );
nor \U$63100 ( \63477 , \63475 , \63476 );
and \U$63101 ( \63478 , \63477 , \4481 );
not \U$63102 ( \63479 , \63477 );
and \U$63103 ( \63480 , \63479 , \4482 );
nor \U$63104 ( \63481 , \63478 , \63480 );
xor \U$63105 ( \63482 , \63474 , \63481 );
xor \U$63106 ( \63483 , \63461 , \63482 );
not \U$63107 ( \63484 , \789 );
and \U$63108 ( \63485 , \883 , RIae75dd0_28);
and \U$63109 ( \63486 , RIae75650_12, \881 );
nor \U$63110 ( \63487 , \63485 , \63486 );
not \U$63111 ( \63488 , \63487 );
or \U$63112 ( \63489 , \63484 , \63488 );
or \U$63113 ( \63490 , \63487 , \789 );
nand \U$63114 ( \63491 , \63489 , \63490 );
and \U$63115 ( \63492 , \558 , RIae75920_18);
and \U$63116 ( \63493 , RIae75fb0_32, \556 );
nor \U$63117 ( \63494 , \63492 , \63493 );
and \U$63118 ( \63495 , \63494 , \504 );
not \U$63119 ( \63496 , \63494 );
and \U$63120 ( \63497 , \63496 , \562 );
nor \U$63121 ( \63498 , \63495 , \63497 );
xor \U$63122 ( \63499 , \63491 , \63498 );
and \U$63123 ( \63500 , \672 , RIae75ec0_30);
and \U$63124 ( \63501 , RIae75ce0_26, \670 );
nor \U$63125 ( \63502 , \63500 , \63501 );
and \U$63126 ( \63503 , \63502 , \588 );
not \U$63127 ( \63504 , \63502 );
and \U$63128 ( \63505 , \63504 , \587 );
nor \U$63129 ( \63506 , \63503 , \63505 );
xor \U$63130 ( \63507 , \63499 , \63506 );
and \U$63131 ( \63508 , \1376 , RIae75740_14);
and \U$63132 ( \63509 , RIae75290_4, \1374 );
nor \U$63133 ( \63510 , \63508 , \63509 );
and \U$63134 ( \63511 , \63510 , \1380 );
not \U$63135 ( \63512 , \63510 );
and \U$63136 ( \63513 , \63512 , \1261 );
nor \U$63137 ( \63514 , \63511 , \63513 );
and \U$63138 ( \63515 , \1138 , RIae75560_10);
and \U$63139 ( \63516 , RIae75830_16, \1136 );
nor \U$63140 ( \63517 , \63515 , \63516 );
and \U$63141 ( \63518 , \63517 , \1012 );
not \U$63142 ( \63519 , \63517 );
and \U$63143 ( \63520 , \63519 , \1142 );
nor \U$63144 ( \63521 , \63518 , \63520 );
xor \U$63145 ( \63522 , \63514 , \63521 );
and \U$63146 ( \63523 , \1593 , RIae751a0_2);
and \U$63147 ( \63524 , RIae75380_6, \1591 );
nor \U$63148 ( \63525 , \63523 , \63524 );
and \U$63149 ( \63526 , \63525 , \1498 );
not \U$63150 ( \63527 , \63525 );
and \U$63151 ( \63528 , \63527 , \1488 );
nor \U$63152 ( \63529 , \63526 , \63528 );
xor \U$63153 ( \63530 , \63522 , \63529 );
and \U$63154 ( \63531 , \1939 , RIae75470_8);
and \U$63155 ( \63532 , RIae76460_42, \1937 );
nor \U$63156 ( \63533 , \63531 , \63532 );
and \U$63157 ( \63534 , \63533 , \1735 );
not \U$63158 ( \63535 , \63533 );
and \U$63159 ( \63536 , \63535 , \1734 );
nor \U$63160 ( \63537 , \63534 , \63536 );
and \U$63161 ( \63538 , \2224 , RIae76550_44);
and \U$63162 ( \63539 , RIae76730_48, \2222 );
nor \U$63163 ( \63540 , \63538 , \63539 );
and \U$63164 ( \63541 , \63540 , \2061 );
not \U$63165 ( \63542 , \63540 );
and \U$63166 ( \63543 , \63542 , \2060 );
nor \U$63167 ( \63544 , \63541 , \63543 );
xor \U$63168 ( \63545 , \63537 , \63544 );
and \U$63169 ( \63546 , \2607 , RIae76640_46);
and \U$63170 ( \63547 , RIae76190_36, \2605 );
nor \U$63171 ( \63548 , \63546 , \63547 );
and \U$63172 ( \63549 , \63548 , \2611 );
not \U$63173 ( \63550 , \63548 );
and \U$63174 ( \63551 , \63550 , \2397 );
nor \U$63175 ( \63552 , \63549 , \63551 );
xor \U$63176 ( \63553 , \63545 , \63552 );
xor \U$63177 ( \63554 , \63530 , \63553 );
xor \U$63178 ( \63555 , \63507 , \63554 );
xor \U$63179 ( \63556 , \63483 , \63555 );
xor \U$63180 ( \63557 , \63423 , \63556 );
xor \U$63181 ( \63558 , \38269 , \38273 );
and \U$63182 ( \63559 , \63558 , \38278 );
and \U$63183 ( \63560 , \38269 , \38273 );
or \U$63184 ( \63561 , \63559 , \63560 );
xor \U$63185 ( \63562 , \38301 , \38303 );
and \U$63186 ( \63563 , \63562 , \37997 );
and \U$63187 ( \63564 , \38301 , \38303 );
or \U$63188 ( \63565 , \63563 , \63564 );
xor \U$63189 ( \63566 , \63561 , \63565 );
xor \U$63190 ( \63567 , \38283 , \38287 );
and \U$63191 ( \63568 , \63567 , \38292 );
and \U$63192 ( \63569 , \38283 , \38287 );
or \U$63193 ( \63570 , \63568 , \63569 );
xor \U$63194 ( \63571 , \63566 , \63570 );
xor \U$63195 ( \63572 , \38283 , \38287 );
xor \U$63196 ( \63573 , \63572 , \38292 );
and \U$63197 ( \63574 , \38305 , \63573 );
xor \U$63198 ( \63575 , \38283 , \38287 );
xor \U$63199 ( \63576 , \63575 , \38292 );
and \U$63200 ( \63577 , \38379 , \63576 );
and \U$63201 ( \63578 , \38305 , \38379 );
or \U$63202 ( \63579 , \63574 , \63577 , \63578 );
xor \U$63203 ( \63580 , \38461 , \38465 );
and \U$63204 ( \63581 , \63580 , \38470 );
and \U$63205 ( \63582 , \38461 , \38465 );
or \U$63206 ( \63583 , \63581 , \63582 );
xor \U$63207 ( \63584 , \63579 , \63583 );
xor \U$63208 ( \63585 , \38196 , \38197 );
and \U$63209 ( \63586 , \63585 , \38264 );
and \U$63210 ( \63587 , \38196 , \38197 );
or \U$63211 ( \63588 , \63586 , \63587 );
xor \U$63212 ( \63589 , \63584 , \63588 );
xor \U$63213 ( \63590 , \63571 , \63589 );
xor \U$63214 ( \63591 , \63557 , \63590 );
xor \U$63215 ( \63592 , \63394 , \63591 );
xor \U$63216 ( \63593 , \63388 , \63592 );
xor \U$63217 ( \63594 , \38174 , \38384 );
xor \U$63218 ( \63595 , \63594 , \38481 );
and \U$63219 ( \63596 , \38759 , \63595 );
xor \U$63220 ( \63597 , \38174 , \38384 );
xor \U$63221 ( \63598 , \63597 , \38481 );
and \U$63222 ( \63599 , \39061 , \63598 );
and \U$63223 ( \63600 , \38759 , \39061 );
or \U$63224 ( \63601 , \63596 , \63599 , \63600 );
xor \U$63225 ( \63602 , \63593 , \63601 );
and \U$63226 ( \63603 , \63326 , \63602 );
and \U$63227 ( \63604 , \63593 , \63601 );
nor \U$63228 ( \63605 , \63603 , \63604 );
not \U$63229 ( \63606 , \63605 );
xor \U$63230 ( \63607 , \63330 , \63387 );
and \U$63231 ( \63608 , \63607 , \63592 );
and \U$63232 ( \63609 , \63330 , \63387 );
or \U$63233 ( \63610 , \63608 , \63609 );
xor \U$63234 ( \63611 , \63392 , \63393 );
and \U$63235 ( \63612 , \63611 , \63591 );
and \U$63236 ( \63613 , \63392 , \63393 );
or \U$63237 ( \63614 , \63612 , \63613 );
xor \U$63238 ( \63615 , \63579 , \63583 );
and \U$63239 ( \63616 , \63615 , \63588 );
and \U$63240 ( \63617 , \63579 , \63583 );
or \U$63241 ( \63618 , \63616 , \63617 );
xor \U$63242 ( \63619 , \63408 , \63422 );
and \U$63243 ( \63620 , \63619 , \63556 );
and \U$63244 ( \63621 , \63408 , \63422 );
or \U$63245 ( \63622 , \63620 , \63621 );
xor \U$63246 ( \63623 , \63618 , \63622 );
xor \U$63247 ( \63624 , \63491 , \63498 );
xor \U$63248 ( \63625 , \63624 , \63506 );
and \U$63249 ( \63626 , \63530 , \63625 );
xor \U$63250 ( \63627 , \63491 , \63498 );
xor \U$63251 ( \63628 , \63627 , \63506 );
and \U$63252 ( \63629 , \63553 , \63628 );
and \U$63253 ( \63630 , \63530 , \63553 );
or \U$63254 ( \63631 , \63626 , \63629 , \63630 );
xor \U$63255 ( \63632 , \37004 , \5016 );
xor \U$63256 ( \63633 , \63632 , \37012 );
xor \U$63257 ( \63634 , \63631 , \63633 );
xor \U$63258 ( \63635 , \37075 , \37082 );
xor \U$63259 ( \63636 , \63635 , \37090 );
xor \U$63260 ( \63637 , \36979 , \36986 );
xor \U$63261 ( \63638 , \63637 , \36994 );
xor \U$63262 ( \63639 , \37023 , \37031 );
xor \U$63263 ( \63640 , \63639 , \37040 );
xor \U$63264 ( \63641 , \63638 , \63640 );
xor \U$63265 ( \63642 , \63636 , \63641 );
xor \U$63266 ( \63643 , \63634 , \63642 );
xor \U$63267 ( \63644 , \63398 , \63402 );
and \U$63268 ( \63645 , \63644 , \63407 );
and \U$63269 ( \63646 , \63398 , \63402 );
or \U$63270 ( \63647 , \63645 , \63646 );
xor \U$63271 ( \63648 , \63647 , \63460 );
xor \U$63272 ( \63649 , \63412 , \63416 );
and \U$63273 ( \63650 , \63649 , \63421 );
and \U$63274 ( \63651 , \63412 , \63416 );
or \U$63275 ( \63652 , \63650 , \63651 );
xor \U$63276 ( \63653 , \63648 , \63652 );
xor \U$63277 ( \63654 , \63514 , \63521 );
and \U$63278 ( \63655 , \63654 , \63529 );
and \U$63279 ( \63656 , \63514 , \63521 );
or \U$63280 ( \63657 , \63655 , \63656 );
xor \U$63281 ( \63658 , \63491 , \63498 );
and \U$63282 ( \63659 , \63658 , \63506 );
and \U$63283 ( \63660 , \63491 , \63498 );
or \U$63284 ( \63661 , \63659 , \63660 );
xor \U$63285 ( \63662 , \63657 , \63661 );
or \U$63286 ( \63663 , \63453 , \63431 );
not \U$63287 ( \63664 , \63431 );
not \U$63288 ( \63665 , \63453 );
or \U$63289 ( \63666 , \63664 , \63665 );
nand \U$63290 ( \63667 , \63666 , \63440 );
nand \U$63291 ( \63668 , \63663 , \63667 );
xor \U$63292 ( \63669 , \63662 , \63668 );
xor \U$63293 ( \63670 , \63350 , \63358 );
and \U$63294 ( \63671 , \63670 , \63366 );
and \U$63295 ( \63672 , \63350 , \63358 );
or \U$63296 ( \63673 , \63671 , \63672 );
xor \U$63297 ( \63674 , \63468 , \63473 );
and \U$63298 ( \63675 , \63674 , \63481 );
and \U$63299 ( \63676 , \63468 , \63473 );
or \U$63300 ( \63677 , \63675 , \63676 );
xor \U$63301 ( \63678 , \63673 , \63677 );
xor \U$63302 ( \63679 , \63537 , \63544 );
and \U$63303 ( \63680 , \63679 , \63552 );
and \U$63304 ( \63681 , \63537 , \63544 );
or \U$63305 ( \63682 , \63680 , \63681 );
xor \U$63306 ( \63683 , \63678 , \63682 );
xor \U$63307 ( \63684 , \37128 , \37136 );
xor \U$63308 ( \63685 , \63684 , \37145 );
not \U$63309 ( \63686 , RIae788f0_120);
nor \U$63310 ( \63687 , \63686 , \491 );
xor \U$63311 ( \63688 , \37100 , \37107 );
xor \U$63312 ( \63689 , \63688 , \37116 );
xor \U$63313 ( \63690 , \63687 , \63689 );
xor \U$63314 ( \63691 , \63685 , \63690 );
xor \U$63315 ( \63692 , \63683 , \63691 );
xor \U$63316 ( \63693 , \63669 , \63692 );
xor \U$63317 ( \63694 , \63653 , \63693 );
xor \U$63318 ( \63695 , \63643 , \63694 );
xor \U$63319 ( \63696 , \63623 , \63695 );
xor \U$63320 ( \63697 , \63614 , \63696 );
xor \U$63321 ( \63698 , \63342 , \63367 );
and \U$63322 ( \63699 , \63698 , \63376 );
and \U$63323 ( \63700 , \63342 , \63367 );
or \U$63324 ( \63701 , \63699 , \63700 );
xor \U$63325 ( \63702 , \63561 , \63565 );
and \U$63326 ( \63703 , \63702 , \63570 );
and \U$63327 ( \63704 , \63561 , \63565 );
or \U$63328 ( \63705 , \63703 , \63704 );
xor \U$63329 ( \63706 , \63701 , \63705 );
xor \U$63330 ( \63707 , \63461 , \63482 );
and \U$63331 ( \63708 , \63707 , \63555 );
and \U$63332 ( \63709 , \63461 , \63482 );
or \U$63333 ( \63710 , \63708 , \63709 );
xor \U$63334 ( \63711 , \63706 , \63710 );
xor \U$63335 ( \63712 , \63408 , \63422 );
xor \U$63336 ( \63713 , \63712 , \63556 );
and \U$63337 ( \63714 , \63571 , \63713 );
xor \U$63338 ( \63715 , \63408 , \63422 );
xor \U$63339 ( \63716 , \63715 , \63556 );
and \U$63340 ( \63717 , \63589 , \63716 );
and \U$63341 ( \63718 , \63571 , \63589 );
or \U$63342 ( \63719 , \63714 , \63717 , \63718 );
xor \U$63343 ( \63720 , \63711 , \63719 );
xor \U$63344 ( \63721 , \63334 , \63377 );
and \U$63345 ( \63722 , \63721 , \63386 );
and \U$63346 ( \63723 , \63334 , \63377 );
or \U$63347 ( \63724 , \63722 , \63723 );
xor \U$63348 ( \63725 , \63720 , \63724 );
xor \U$63349 ( \63726 , \63697 , \63725 );
xor \U$63350 ( \63727 , \63610 , \63726 );
and \U$63351 ( \63728 , \63606 , \63727 );
and \U$63352 ( \63729 , \63610 , \63726 );
nor \U$63353 ( \63730 , \63728 , \63729 );
not \U$63354 ( \63731 , \63730 );
xor \U$63355 ( \63732 , \63711 , \63719 );
and \U$63356 ( \63733 , \63732 , \63724 );
and \U$63357 ( \63734 , \63711 , \63719 );
nor \U$63358 ( \63735 , \63733 , \63734 );
not \U$63359 ( \63736 , \63735 );
xor \U$63360 ( \63737 , \63618 , \63622 );
and \U$63361 ( \63738 , \63737 , \63695 );
and \U$63362 ( \63739 , \63618 , \63622 );
or \U$63363 ( \63740 , \63738 , \63739 );
xor \U$63364 ( \63741 , \63657 , \63661 );
xor \U$63365 ( \63742 , \63741 , \63668 );
and \U$63366 ( \63743 , \63683 , \63742 );
xor \U$63367 ( \63744 , \63657 , \63661 );
xor \U$63368 ( \63745 , \63744 , \63668 );
and \U$63369 ( \63746 , \63691 , \63745 );
and \U$63370 ( \63747 , \63683 , \63691 );
or \U$63371 ( \63748 , \63743 , \63746 , \63747 );
xor \U$63372 ( \63749 , \63647 , \63460 );
and \U$63373 ( \63750 , \63749 , \63652 );
and \U$63374 ( \63751 , \63647 , \63460 );
or \U$63375 ( \63752 , \63750 , \63751 );
xor \U$63376 ( \63753 , \63748 , \63752 );
xor \U$63377 ( \63754 , \63631 , \63633 );
and \U$63378 ( \63755 , \63754 , \63642 );
and \U$63379 ( \63756 , \63631 , \63633 );
or \U$63380 ( \63757 , \63755 , \63756 );
xor \U$63381 ( \63758 , \63753 , \63757 );
xor \U$63382 ( \63759 , \63740 , \63758 );
xor \U$63383 ( \63760 , \63631 , \63633 );
xor \U$63384 ( \63761 , \63760 , \63642 );
and \U$63385 ( \63762 , \63653 , \63761 );
xor \U$63386 ( \63763 , \63631 , \63633 );
xor \U$63387 ( \63764 , \63763 , \63642 );
and \U$63388 ( \63765 , \63693 , \63764 );
and \U$63389 ( \63766 , \63653 , \63693 );
or \U$63390 ( \63767 , \63762 , \63765 , \63766 );
xor \U$63391 ( \63768 , \63701 , \63705 );
and \U$63392 ( \63769 , \63768 , \63710 );
and \U$63393 ( \63770 , \63701 , \63705 );
or \U$63394 ( \63771 , \63769 , \63770 );
xor \U$63395 ( \63772 , \63767 , \63771 );
xor \U$63396 ( \63773 , \37075 , \37082 );
xor \U$63397 ( \63774 , \63773 , \37090 );
and \U$63398 ( \63775 , \63638 , \63774 );
xor \U$63399 ( \63776 , \37075 , \37082 );
xor \U$63400 ( \63777 , \63776 , \37090 );
and \U$63401 ( \63778 , \63640 , \63777 );
and \U$63402 ( \63779 , \63638 , \63640 );
or \U$63403 ( \63780 , \63775 , \63778 , \63779 );
xor \U$63404 ( \63781 , \36752 , \36757 );
xor \U$63405 ( \63782 , \63781 , \36765 );
xor \U$63406 ( \63783 , \63780 , \63782 );
xor \U$63407 ( \63784 , \36776 , \36784 );
xor \U$63408 ( \63785 , \63784 , \36793 );
xor \U$63409 ( \63786 , \37162 , \37167 );
xor \U$63410 ( \63787 , \63785 , \63786 );
xor \U$63411 ( \63788 , \63783 , \63787 );
xor \U$63412 ( \63789 , \63657 , \63661 );
and \U$63413 ( \63790 , \63789 , \63668 );
and \U$63414 ( \63791 , \63657 , \63661 );
or \U$63415 ( \63792 , \63790 , \63791 );
xor \U$63416 ( \63793 , \63673 , \63677 );
and \U$63417 ( \63794 , \63793 , \63682 );
and \U$63418 ( \63795 , \63673 , \63677 );
or \U$63419 ( \63796 , \63794 , \63795 );
xor \U$63420 ( \63797 , \63792 , \63796 );
xor \U$63421 ( \63798 , \37128 , \37136 );
xor \U$63422 ( \63799 , \63798 , \37145 );
and \U$63423 ( \63800 , \63687 , \63799 );
xor \U$63424 ( \63801 , \37128 , \37136 );
xor \U$63425 ( \63802 , \63801 , \37145 );
and \U$63426 ( \63803 , \63689 , \63802 );
and \U$63427 ( \63804 , \63687 , \63689 );
or \U$63428 ( \63805 , \63800 , \63803 , \63804 );
xor \U$63429 ( \63806 , \63797 , \63805 );
xor \U$63430 ( \63807 , \36997 , \37015 );
xor \U$63431 ( \63808 , \63807 , \37043 );
or \U$63432 ( \63809 , \37056 , \37066 );
nand \U$63433 ( \63810 , \63809 , \37067 );
xor \U$63434 ( \63811 , \37093 , \37119 );
xor \U$63435 ( \63812 , \63811 , \37148 );
xor \U$63436 ( \63813 , \63810 , \63812 );
xor \U$63437 ( \63814 , \63808 , \63813 );
xor \U$63438 ( \63815 , \63806 , \63814 );
xor \U$63439 ( \63816 , \63788 , \63815 );
xor \U$63440 ( \63817 , \63772 , \63816 );
xor \U$63441 ( \63818 , \63759 , \63817 );
not \U$63442 ( \63819 , \63818 );
or \U$63443 ( \63820 , \63736 , \63819 );
or \U$63444 ( \63821 , \63818 , \63735 );
nand \U$63445 ( \63822 , \63820 , \63821 );
xor \U$63446 ( \63823 , \63614 , \63696 );
and \U$63447 ( \63824 , \63823 , \63725 );
and \U$63448 ( \63825 , \63614 , \63696 );
or \U$63449 ( \63826 , \63824 , \63825 );
xor \U$63450 ( \63827 , \63822 , \63826 );
and \U$63451 ( \63828 , \63731 , \63827 );
and \U$63452 ( \63829 , \63822 , \63826 );
nor \U$63453 ( \63830 , \63828 , \63829 );
xor \U$63454 ( \63831 , \63740 , \63758 );
and \U$63455 ( \63832 , \63831 , \63817 );
and \U$63456 ( \63833 , \63740 , \63758 );
or \U$63457 ( \63834 , \63832 , \63833 );
xor \U$63458 ( \63835 , \63767 , \63771 );
and \U$63459 ( \63836 , \63835 , \63816 );
and \U$63460 ( \63837 , \63767 , \63771 );
or \U$63461 ( \63838 , \63836 , \63837 );
xor \U$63462 ( \63839 , \36997 , \37015 );
xor \U$63463 ( \63840 , \63839 , \37043 );
and \U$63464 ( \63841 , \63810 , \63840 );
xor \U$63465 ( \63842 , \36997 , \37015 );
xor \U$63466 ( \63843 , \63842 , \37043 );
and \U$63467 ( \63844 , \63812 , \63843 );
and \U$63468 ( \63845 , \63810 , \63812 );
or \U$63469 ( \63846 , \63841 , \63844 , \63845 );
xor \U$63470 ( \63847 , \63792 , \63796 );
and \U$63471 ( \63848 , \63847 , \63805 );
and \U$63472 ( \63849 , \63792 , \63796 );
or \U$63473 ( \63850 , \63848 , \63849 );
xor \U$63474 ( \63851 , \63846 , \63850 );
xor \U$63475 ( \63852 , \63780 , \63782 );
and \U$63476 ( \63853 , \63852 , \63787 );
and \U$63477 ( \63854 , \63780 , \63782 );
or \U$63478 ( \63855 , \63853 , \63854 );
xor \U$63479 ( \63856 , \63851 , \63855 );
xor \U$63480 ( \63857 , \63838 , \63856 );
xor \U$63481 ( \63858 , \63780 , \63782 );
xor \U$63482 ( \63859 , \63858 , \63787 );
and \U$63483 ( \63860 , \63806 , \63859 );
xor \U$63484 ( \63861 , \63780 , \63782 );
xor \U$63485 ( \63862 , \63861 , \63787 );
and \U$63486 ( \63863 , \63814 , \63862 );
and \U$63487 ( \63864 , \63806 , \63814 );
or \U$63488 ( \63865 , \63860 , \63863 , \63864 );
xor \U$63489 ( \63866 , \63748 , \63752 );
and \U$63490 ( \63867 , \63866 , \63757 );
and \U$63491 ( \63868 , \63748 , \63752 );
or \U$63492 ( \63869 , \63867 , \63868 );
xor \U$63493 ( \63870 , \63865 , \63869 );
xor \U$63494 ( \63871 , \37046 , \37067 );
xor \U$63495 ( \63872 , \63871 , \37151 );
xor \U$63496 ( \63873 , \37156 , \37158 );
xor \U$63497 ( \63874 , \36883 , \36885 );
xor \U$63498 ( \63875 , \63874 , \36888 );
xor \U$63499 ( \63876 , \37172 , \37179 );
xor \U$63500 ( \63877 , \63875 , \63876 );
xor \U$63501 ( \63878 , \63873 , \63877 );
xor \U$63502 ( \63879 , \63872 , \63878 );
xor \U$63503 ( \63880 , \63870 , \63879 );
xor \U$63504 ( \63881 , \63857 , \63880 );
xor \U$63505 ( \63882 , \63834 , \63881 );
not \U$63506 ( \63883 , \63882 );
not \U$63507 ( \63884 , \63735 );
nand \U$63508 ( \63885 , \63884 , \63818 );
not \U$63509 ( \63886 , \63885 );
and \U$63510 ( \63887 , \63883 , \63886 );
and \U$63511 ( \63888 , \63882 , \63885 );
nor \U$63512 ( \63889 , \63887 , \63888 );
or \U$63513 ( \63890 , \63830 , \63889 );
not \U$63514 ( \63891 , \63882 );
or \U$63515 ( \63892 , \63885 , \63891 );
nand \U$63516 ( \63893 , \63890 , \63892 );
and \U$63517 ( \63894 , \63834 , \63881 );
xor \U$63518 ( \63895 , \63838 , \63856 );
and \U$63519 ( \63896 , \63895 , \63880 );
and \U$63520 ( \63897 , \63838 , \63856 );
or \U$63521 ( \63898 , \63896 , \63897 );
xor \U$63522 ( \63899 , \63865 , \63869 );
and \U$63523 ( \63900 , \63899 , \63879 );
and \U$63524 ( \63901 , \63865 , \63869 );
or \U$63525 ( \63902 , \63900 , \63901 );
xor \U$63526 ( \63903 , \37154 , \37159 );
xor \U$63527 ( \63904 , \63903 , \37184 );
xor \U$63528 ( \63905 , \63902 , \63904 );
xor \U$63529 ( \63906 , \63846 , \63850 );
and \U$63530 ( \63907 , \63906 , \63855 );
and \U$63531 ( \63908 , \63846 , \63850 );
or \U$63532 ( \63909 , \63907 , \63908 );
xor \U$63533 ( \63910 , \37046 , \37067 );
xor \U$63534 ( \63911 , \63910 , \37151 );
and \U$63535 ( \63912 , \63873 , \63911 );
xor \U$63536 ( \63913 , \37046 , \37067 );
xor \U$63537 ( \63914 , \63913 , \37151 );
and \U$63538 ( \63915 , \63877 , \63914 );
and \U$63539 ( \63916 , \63873 , \63877 );
or \U$63540 ( \63917 , \63912 , \63915 , \63916 );
xor \U$63541 ( \63918 , \63909 , \63917 );
xor \U$63542 ( \63919 , \36799 , \36880 );
xor \U$63543 ( \63920 , \63919 , \36891 );
xor \U$63544 ( \63921 , \36959 , \36966 );
xor \U$63545 ( \63922 , \63920 , \63921 );
xor \U$63546 ( \63923 , \63918 , \63922 );
xor \U$63547 ( \63924 , \63905 , \63923 );
xor \U$63548 ( \63925 , \63898 , \63924 );
xor \U$63549 ( \63926 , \63894 , \63925 );
and \U$63550 ( \63927 , \63893 , \63926 );
and \U$63551 ( \63928 , \63894 , \63925 );
nor \U$63552 ( \63929 , \63927 , \63928 );
nand \U$63553 ( \63930 , \63898 , \63924 );
xor \U$63554 ( \63931 , \63909 , \63917 );
and \U$63555 ( \63932 , \63931 , \63922 );
and \U$63556 ( \63933 , \63909 , \63917 );
or \U$63557 ( \63934 , \63932 , \63933 );
not \U$63558 ( \63935 , \63934 );
xnor \U$63559 ( \63936 , \36894 , \36919 );
not \U$63560 ( \63937 , \63936 );
not \U$63561 ( \63938 , \36719 );
and \U$63562 ( \63939 , \63937 , \63938 );
and \U$63563 ( \63940 , \63936 , \36719 );
nor \U$63564 ( \63941 , \63939 , \63940 );
not \U$63565 ( \63942 , \63941 );
and \U$63566 ( \63943 , \63935 , \63942 );
and \U$63567 ( \63944 , \63934 , \63941 );
nor \U$63568 ( \63945 , \63943 , \63944 );
not \U$63569 ( \63946 , \63945 );
xor \U$63570 ( \63947 , \36958 , \36971 );
xor \U$63571 ( \63948 , \63947 , \37187 );
not \U$63572 ( \63949 , \63948 );
and \U$63573 ( \63950 , \63946 , \63949 );
and \U$63574 ( \63951 , \63945 , \63948 );
nor \U$63575 ( \63952 , \63950 , \63951 );
not \U$63576 ( \63953 , \63952 );
xor \U$63577 ( \63954 , \63902 , \63904 );
and \U$63578 ( \63955 , \63954 , \63923 );
and \U$63579 ( \63956 , \63902 , \63904 );
or \U$63580 ( \63957 , \63955 , \63956 );
not \U$63581 ( \63958 , \63957 );
and \U$63582 ( \63959 , \63953 , \63958 );
and \U$63583 ( \63960 , \63952 , \63957 );
nor \U$63584 ( \63961 , \63959 , \63960 );
xnor \U$63585 ( \63962 , \63930 , \63961 );
or \U$63586 ( \63963 , \63929 , \63962 );
or \U$63587 ( \63964 , \63930 , \63961 );
nand \U$63588 ( \63965 , \63963 , \63964 );
not \U$63589 ( \63966 , \63957 );
nor \U$63590 ( \63967 , \63966 , \63952 );
not \U$63591 ( \63968 , \63948 );
or \U$63592 ( \63969 , \63968 , \63941 );
not \U$63593 ( \63970 , \63941 );
not \U$63594 ( \63971 , \63968 );
or \U$63595 ( \63972 , \63970 , \63971 );
nand \U$63596 ( \63973 , \63972 , \63934 );
nand \U$63597 ( \63974 , \63969 , \63973 );
not \U$63598 ( \63975 , \63974 );
xor \U$63599 ( \63976 , \36945 , \36955 );
xor \U$63600 ( \63977 , \63976 , \37190 );
not \U$63601 ( \63978 , \63977 );
or \U$63602 ( \63979 , \63975 , \63978 );
or \U$63603 ( \63980 , \63977 , \63974 );
nand \U$63604 ( \63981 , \63979 , \63980 );
xor \U$63605 ( \63982 , \63967 , \63981 );
and \U$63606 ( \63983 , \63965 , \63982 );
and \U$63607 ( \63984 , \63967 , \63981 );
nor \U$63608 ( \63985 , \63983 , \63984 );
not \U$63609 ( \63986 , \63977 );
nand \U$63610 ( \63987 , \63986 , \63974 );
not \U$63611 ( \63988 , \36938 );
not \U$63612 ( \63989 , \37193 );
and \U$63613 ( \63990 , \63988 , \63989 );
and \U$63614 ( \63991 , \36938 , \37193 );
nor \U$63615 ( \63992 , \63990 , \63991 );
xnor \U$63616 ( \63993 , \63987 , \63992 );
or \U$63617 ( \63994 , \63985 , \63993 );
or \U$63618 ( \63995 , \63987 , \63992 );
nand \U$63619 ( \63996 , \63994 , \63995 );
and \U$63620 ( \63997 , \37196 , \63996 );
nor \U$63621 ( \63998 , \37195 , \63997 );
or \U$63622 ( \63999 , \36933 , \63998 );
nand \U$63623 ( \64000 , \36932 , \63999 );
not \U$63624 ( \64001 , \36680 );
nor \U$63625 ( \64002 , \64001 , \36426 );
xor \U$63626 ( \64003 , \36387 , \36389 );
and \U$63627 ( \64004 , \64003 , \36425 );
and \U$63628 ( \64005 , \36387 , \36389 );
or \U$63629 ( \64006 , \64004 , \64005 );
not \U$63630 ( \64007 , \64006 );
not \U$63631 ( \64008 , \35687 );
not \U$63632 ( \64009 , \35698 );
or \U$63633 ( \64010 , \64008 , \64009 );
or \U$63634 ( \64011 , \35698 , \35687 );
nand \U$63635 ( \64012 , \64010 , \64011 );
not \U$63636 ( \64013 , \35716 );
not \U$63637 ( \64014 , \35712 );
not \U$63638 ( \64015 , \35927 );
and \U$63639 ( \64016 , \64014 , \64015 );
and \U$63640 ( \64017 , \35712 , \35927 );
nor \U$63641 ( \64018 , \64016 , \64017 );
not \U$63642 ( \64019 , \64018 );
or \U$63643 ( \64020 , \64013 , \64019 );
or \U$63644 ( \64021 , \64018 , \35716 );
nand \U$63645 ( \64022 , \64020 , \64021 );
xor \U$63646 ( \64023 , \64012 , \64022 );
or \U$63647 ( \64024 , \36421 , \36414 );
not \U$63648 ( \64025 , \36414 );
not \U$63649 ( \64026 , \36421 );
or \U$63650 ( \64027 , \64025 , \64026 );
nand \U$63651 ( \64028 , \64027 , \36405 );
nand \U$63652 ( \64029 , \64024 , \64028 );
xor \U$63653 ( \64030 , \64023 , \64029 );
not \U$63654 ( \64031 , \64030 );
or \U$63655 ( \64032 , \64007 , \64031 );
or \U$63656 ( \64033 , \64030 , \64006 );
nand \U$63657 ( \64034 , \64032 , \64033 );
xor \U$63658 ( \64035 , \64002 , \64034 );
and \U$63659 ( \64036 , \64000 , \64035 );
and \U$63660 ( \64037 , \64002 , \64034 );
nor \U$63661 ( \64038 , \64036 , \64037 );
not \U$63662 ( \64039 , \64006 );
nand \U$63663 ( \64040 , \64039 , \64030 );
not \U$63664 ( \64041 , \35684 );
xor \U$63665 ( \64042 , \35699 , \35929 );
not \U$63666 ( \64043 , \64042 );
or \U$63667 ( \64044 , \64041 , \64043 );
or \U$63668 ( \64045 , \64042 , \35684 );
nand \U$63669 ( \64046 , \64044 , \64045 );
not \U$63670 ( \64047 , \64046 );
xor \U$63671 ( \64048 , \64012 , \64022 );
and \U$63672 ( \64049 , \64048 , \64029 );
and \U$63673 ( \64050 , \64012 , \64022 );
nor \U$63674 ( \64051 , \64049 , \64050 );
not \U$63675 ( \64052 , \64051 );
and \U$63676 ( \64053 , \64047 , \64052 );
and \U$63677 ( \64054 , \64046 , \64051 );
nor \U$63678 ( \64055 , \64053 , \64054 );
xnor \U$63679 ( \64056 , \64040 , \64055 );
or \U$63680 ( \64057 , \64038 , \64056 );
or \U$63681 ( \64058 , \64040 , \64055 );
nand \U$63682 ( \64059 , \64057 , \64058 );
not \U$63683 ( \64060 , \64046 );
nor \U$63684 ( \64061 , \64060 , \64051 );
not \U$63685 ( \64062 , \35931 );
not \U$63686 ( \64063 , \35942 );
or \U$63687 ( \64064 , \64062 , \64063 );
or \U$63688 ( \64065 , \35942 , \35931 );
nand \U$63689 ( \64066 , \64064 , \64065 );
xor \U$63690 ( \64067 , \64061 , \64066 );
and \U$63691 ( \64068 , \64059 , \64067 );
and \U$63692 ( \64069 , \64061 , \64066 );
nor \U$63693 ( \64070 , \64068 , \64069 );
or \U$63694 ( \64071 , \35945 , \64070 );
nand \U$63695 ( \64072 , \35944 , \64071 );
and \U$63696 ( \64073 , \35672 , \64072 );
nor \U$63697 ( \64074 , \35671 , \64073 );
or \U$63698 ( \64075 , \35244 , \64074 );
nand \U$63699 ( \64076 , \35243 , \64075 );
not \U$63700 ( \64077 , \35230 );
nor \U$63701 ( \64078 , \64077 , \35238 );
xor \U$63702 ( \64079 , \35208 , \35218 );
and \U$63703 ( \64080 , \64079 , \35229 );
and \U$63704 ( \64081 , \35208 , \35218 );
or \U$63705 ( \64082 , \64080 , \64081 );
not \U$63706 ( \64083 , \64082 );
xor \U$63707 ( \64084 , \34664 , \34666 );
xor \U$63708 ( \64085 , \64084 , \34669 );
not \U$63709 ( \64086 , \64085 );
or \U$63710 ( \64087 , \64083 , \64086 );
or \U$63711 ( \64088 , \64085 , \64082 );
nand \U$63712 ( \64089 , \64087 , \64088 );
xor \U$63713 ( \64090 , \64078 , \64089 );
and \U$63714 ( \64091 , \64076 , \64090 );
and \U$63715 ( \64092 , \64078 , \64089 );
nor \U$63716 ( \64093 , \64091 , \64092 );
not \U$63717 ( \64094 , \64085 );
nand \U$63718 ( \64095 , \64094 , \64082 );
not \U$63719 ( \64096 , \34503 );
not \U$63720 ( \64097 , \34672 );
and \U$63721 ( \64098 , \64096 , \64097 );
and \U$63722 ( \64099 , \34503 , \34672 );
nor \U$63723 ( \64100 , \64098 , \64099 );
xnor \U$63724 ( \64101 , \64095 , \64100 );
or \U$63725 ( \64102 , \64093 , \64101 );
or \U$63726 ( \64103 , \64095 , \64100 );
nand \U$63727 ( \64104 , \64102 , \64103 );
and \U$63728 ( \64105 , \34675 , \64104 );
nor \U$63729 ( \64106 , \34674 , \64105 );
or \U$63730 ( \64107 , \34492 , \64106 );
nand \U$63731 ( \64108 , \34491 , \64107 );
and \U$63732 ( \64109 , \34300 , \64108 );
nor \U$63733 ( \64110 , \34299 , \64109 );
or \U$63734 ( \64111 , \34125 , \64110 );
nand \U$63735 ( \64112 , \34124 , \64111 );
and \U$63736 ( \64113 , \33941 , \64112 );
nor \U$63737 ( \64114 , \33940 , \64113 );
xor \U$63738 ( \64115 , \33355 , \33378 );
and \U$63739 ( \64116 , \64115 , \33498 );
and \U$63740 ( \64117 , \33355 , \33378 );
or \U$63741 ( \64118 , \64116 , \64117 );
not \U$63742 ( \64119 , \64118 );
or \U$63743 ( \64120 , \33454 , \33479 );
not \U$63744 ( \64121 , \33479 );
not \U$63745 ( \64122 , \33454 );
or \U$63746 ( \64123 , \64121 , \64122 );
nand \U$63747 ( \64124 , \64123 , \33493 );
nand \U$63748 ( \64125 , \64120 , \64124 );
or \U$63749 ( \64126 , \33374 , \33365 );
not \U$63750 ( \64127 , \33365 );
not \U$63751 ( \64128 , \33374 );
or \U$63752 ( \64129 , \64127 , \64128 );
nand \U$63753 ( \64130 , \64129 , \33360 );
nand \U$63754 ( \64131 , \64126 , \64130 );
xor \U$63755 ( \64132 , \64125 , \64131 );
xor \U$63756 ( \64133 , \33081 , \1012 );
xor \U$63757 ( \64134 , \64133 , \33090 );
xor \U$63758 ( \64135 , \33095 , \33103 );
xor \U$63759 ( \64136 , \33113 , \33121 );
xor \U$63760 ( \64137 , \64136 , \33129 );
xor \U$63761 ( \64138 , \64135 , \64137 );
xor \U$63762 ( \64139 , \64134 , \64138 );
xor \U$63763 ( \64140 , \64132 , \64139 );
not \U$63764 ( \64141 , \64140 );
xor \U$63765 ( \64142 , \33387 , \33423 );
and \U$63766 ( \64143 , \64142 , \33497 );
and \U$63767 ( \64144 , \33387 , \33423 );
or \U$63768 ( \64145 , \64143 , \64144 );
not \U$63769 ( \64146 , \64145 );
or \U$63770 ( \64147 , \33450 , \33438 );
not \U$63771 ( \64148 , \33438 );
not \U$63772 ( \64149 , \33450 );
or \U$63773 ( \64150 , \64148 , \64149 );
nand \U$63774 ( \64151 , \64150 , \33429 );
nand \U$63775 ( \64152 , \64147 , \64151 );
xor \U$63776 ( \64153 , \64152 , \33492 );
xor \U$63777 ( \64154 , \33462 , \33469 );
and \U$63778 ( \64155 , \64154 , \33478 );
and \U$63779 ( \64156 , \33462 , \33469 );
nor \U$63780 ( \64157 , \64155 , \64156 );
xor \U$63781 ( \64158 , \64153 , \64157 );
not \U$63782 ( \64159 , \64158 );
and \U$63783 ( \64160 , \64146 , \64159 );
and \U$63784 ( \64161 , \64145 , \64158 );
nor \U$63785 ( \64162 , \64160 , \64161 );
not \U$63786 ( \64163 , \64162 );
or \U$63787 ( \64164 , \64141 , \64163 );
or \U$63788 ( \64165 , \64162 , \64140 );
nand \U$63789 ( \64166 , \64164 , \64165 );
not \U$63790 ( \64167 , \64166 );
and \U$63791 ( \64168 , \64119 , \64167 );
and \U$63792 ( \64169 , \64118 , \64166 );
nor \U$63793 ( \64170 , \64168 , \64169 );
not \U$63794 ( \64171 , \33499 );
not \U$63795 ( \64172 , \33612 );
and \U$63796 ( \64173 , \64171 , \64172 );
and \U$63797 ( \64174 , \33499 , \33612 );
not \U$63798 ( \64175 , \33756 );
nor \U$63799 ( \64176 , \64174 , \64175 );
nor \U$63800 ( \64177 , \64173 , \64176 );
xnor \U$63801 ( \64178 , \64170 , \64177 );
or \U$63802 ( \64179 , \64114 , \64178 );
or \U$63803 ( \64180 , \64170 , \64177 );
nand \U$63804 ( \64181 , \64179 , \64180 );
not \U$63805 ( \64182 , \64166 );
nor \U$63806 ( \64183 , \64182 , \64118 );
and \U$63807 ( \64184 , \64140 , \64158 );
not \U$63808 ( \64185 , \64140 );
not \U$63809 ( \64186 , \64158 );
and \U$63810 ( \64187 , \64185 , \64186 );
nor \U$63811 ( \64188 , \64187 , \64145 );
nor \U$63812 ( \64189 , \64184 , \64188 );
not \U$63813 ( \64190 , \64189 );
xor \U$63814 ( \64191 , \64125 , \64131 );
and \U$63815 ( \64192 , \64191 , \64139 );
and \U$63816 ( \64193 , \64125 , \64131 );
or \U$63817 ( \64194 , \64192 , \64193 );
xor \U$63818 ( \64195 , \33093 , \33104 );
xor \U$63819 ( \64196 , \64195 , \33132 );
xor \U$63820 ( \64197 , \64194 , \64196 );
xor \U$63821 ( \64198 , \33081 , \1012 );
xor \U$63822 ( \64199 , \64198 , \33090 );
and \U$63823 ( \64200 , \64135 , \64199 );
xor \U$63824 ( \64201 , \33081 , \1012 );
xor \U$63825 ( \64202 , \64201 , \33090 );
and \U$63826 ( \64203 , \64137 , \64202 );
and \U$63827 ( \64204 , \64135 , \64137 );
or \U$63828 ( \64205 , \64200 , \64203 , \64204 );
xor \U$63829 ( \64206 , \64152 , \33492 );
and \U$63830 ( \64207 , \64206 , \64157 );
and \U$63831 ( \64208 , \64152 , \33492 );
or \U$63832 ( \64209 , \64207 , \64208 );
xor \U$63833 ( \64210 , \64205 , \64209 );
xor \U$63834 ( \64211 , \32956 , \32964 );
xor \U$63835 ( \64212 , \64211 , \32973 );
xor \U$63836 ( \64213 , \33002 , \33069 );
xor \U$63837 ( \64214 , \64212 , \64213 );
xor \U$63838 ( \64215 , \64210 , \64214 );
xor \U$63839 ( \64216 , \64197 , \64215 );
not \U$63840 ( \64217 , \64216 );
or \U$63841 ( \64218 , \64190 , \64217 );
or \U$63842 ( \64219 , \64216 , \64189 );
nand \U$63843 ( \64220 , \64218 , \64219 );
xor \U$63844 ( \64221 , \64183 , \64220 );
and \U$63845 ( \64222 , \64181 , \64221 );
and \U$63846 ( \64223 , \64183 , \64220 );
nor \U$63847 ( \64224 , \64222 , \64223 );
not \U$63848 ( \64225 , \64189 );
nand \U$63849 ( \64226 , \64225 , \64216 );
xor \U$63850 ( \64227 , \32976 , \33000 );
not \U$63851 ( \64228 , \33002 );
xor \U$63852 ( \64229 , \64227 , \64228 );
xor \U$63853 ( \64230 , \64205 , \64209 );
and \U$63854 ( \64231 , \64230 , \64214 );
and \U$63855 ( \64232 , \64205 , \64209 );
or \U$63856 ( \64233 , \64231 , \64232 );
xnor \U$63857 ( \64234 , \64229 , \64233 );
not \U$63858 ( \64235 , \64234 );
not \U$63859 ( \64236 , \33143 );
xor \U$63860 ( \64237 , \33135 , \33074 );
not \U$63861 ( \64238 , \64237 );
or \U$63862 ( \64239 , \64236 , \64238 );
or \U$63863 ( \64240 , \64237 , \33143 );
nand \U$63864 ( \64241 , \64239 , \64240 );
not \U$63865 ( \64242 , \64241 );
and \U$63866 ( \64243 , \64235 , \64242 );
and \U$63867 ( \64244 , \64234 , \64241 );
nor \U$63868 ( \64245 , \64243 , \64244 );
not \U$63869 ( \64246 , \64245 );
xor \U$63870 ( \64247 , \64194 , \64196 );
and \U$63871 ( \64248 , \64247 , \64215 );
and \U$63872 ( \64249 , \64194 , \64196 );
or \U$63873 ( \64250 , \64248 , \64249 );
not \U$63874 ( \64251 , \64250 );
and \U$63875 ( \64252 , \64246 , \64251 );
and \U$63876 ( \64253 , \64245 , \64250 );
nor \U$63877 ( \64254 , \64252 , \64253 );
xnor \U$63878 ( \64255 , \64226 , \64254 );
or \U$63879 ( \64256 , \64224 , \64255 );
or \U$63880 ( \64257 , \64226 , \64254 );
nand \U$63881 ( \64258 , \64256 , \64257 );
not \U$63882 ( \64259 , \64250 );
nor \U$63883 ( \64260 , \64259 , \64245 );
not \U$63884 ( \64261 , \64229 );
not \U$63885 ( \64262 , \64241 );
or \U$63886 ( \64263 , \64261 , \64262 );
or \U$63887 ( \64264 , \64241 , \64229 );
nand \U$63888 ( \64265 , \64264 , \64233 );
nand \U$63889 ( \64266 , \64263 , \64265 );
not \U$63890 ( \64267 , \64266 );
xor \U$63891 ( \64268 , \33145 , \33150 );
xor \U$63892 ( \64269 , \64268 , \33153 );
not \U$63893 ( \64270 , \64269 );
or \U$63894 ( \64271 , \64267 , \64270 );
or \U$63895 ( \64272 , \64269 , \64266 );
nand \U$63896 ( \64273 , \64271 , \64272 );
xor \U$63897 ( \64274 , \64260 , \64273 );
and \U$63898 ( \64275 , \64258 , \64274 );
and \U$63899 ( \64276 , \64260 , \64273 );
nor \U$63900 ( \64277 , \64275 , \64276 );
not \U$63901 ( \64278 , \33156 );
not \U$63902 ( \64279 , \33063 );
and \U$63903 ( \64280 , \64278 , \64279 );
and \U$63904 ( \64281 , \33156 , \33063 );
nor \U$63905 ( \64282 , \64280 , \64281 );
not \U$63906 ( \64283 , \64269 );
nand \U$63907 ( \64284 , \64283 , \64266 );
xnor \U$63908 ( \64285 , \64282 , \64284 );
or \U$63909 ( \64286 , \64277 , \64285 );
or \U$63910 ( \64287 , \64284 , \64282 );
nand \U$63911 ( \64288 , \64286 , \64287 );
and \U$63912 ( \64289 , \33159 , \64288 );
nor \U$63913 ( \64290 , \33158 , \64289 );
or \U$63914 ( \64291 , \33043 , \64290 );
nand \U$63915 ( \64292 , \33042 , \64291 );
and \U$63916 ( \64293 , \32855 , \64292 );
nor \U$63917 ( \64294 , \32854 , \64293 );
or \U$63918 ( \64295 , \32761 , \64294 );
nand \U$63919 ( \64296 , \32760 , \64295 );
not \U$63920 ( \64297 , \32694 );
nor \U$63921 ( \64298 , \64297 , \32635 );
or \U$63922 ( \64299 , \32555 , \32553 );
nand \U$63923 ( \64300 , \64299 , \32556 );
or \U$63924 ( \64301 , \32631 , \32561 );
not \U$63925 ( \64302 , \32561 );
not \U$63926 ( \64303 , \32631 );
or \U$63927 ( \64304 , \64302 , \64303 );
nand \U$63928 ( \64305 , \64304 , \32611 );
nand \U$63929 ( \64306 , \64301 , \64305 );
xor \U$63930 ( \64307 , \64300 , \64306 );
or \U$63931 ( \64308 , \32583 , \32627 );
not \U$63932 ( \64309 , \32627 );
not \U$63933 ( \64310 , \32583 );
or \U$63934 ( \64311 , \64309 , \64310 );
nand \U$63935 ( \64312 , \64311 , \32621 );
nand \U$63936 ( \64313 , \64308 , \64312 );
xor \U$63937 ( \64314 , \64307 , \64313 );
xor \U$63938 ( \64315 , \64298 , \64314 );
and \U$63939 ( \64316 , \64296 , \64315 );
and \U$63940 ( \64317 , \64298 , \64314 );
nor \U$63941 ( \64318 , \64316 , \64317 );
not \U$63942 ( \64319 , \32529 );
not \U$63943 ( \64320 , \32556 );
or \U$63944 ( \64321 , \64319 , \64320 );
or \U$63945 ( \64322 , \32556 , \32529 );
nand \U$63946 ( \64323 , \64321 , \64322 );
not \U$63947 ( \64324 , \64323 );
not \U$63948 ( \64325 , \32510 );
and \U$63949 ( \64326 , \64324 , \64325 );
and \U$63950 ( \64327 , \64323 , \32510 );
nor \U$63951 ( \64328 , \64326 , \64327 );
xor \U$63952 ( \64329 , \64300 , \64306 );
and \U$63953 ( \64330 , \64329 , \64313 );
and \U$63954 ( \64331 , \64300 , \64306 );
nor \U$63955 ( \64332 , \64330 , \64331 );
xnor \U$63956 ( \64333 , \64328 , \64332 );
or \U$63957 ( \64334 , \64318 , \64333 );
or \U$63958 ( \64335 , \64328 , \64332 );
nand \U$63959 ( \64336 , \64334 , \64335 );
and \U$63960 ( \64337 , \32559 , \64336 );
and \U$63961 ( \64338 , \32558 , \32500 );
and \U$63962 ( \64339 , \32484 , \32499 );
nor \U$63963 ( \64340 , \64337 , \64338 , \64339 );
not \U$63964 ( \64341 , \64340 );
nand \U$63965 ( \64342 , RIae78b48_125, RIae78da0_130);
not \U$63966 ( \64343 , \64342 );
not \U$63967 ( \64344 , \397 );
or \U$63968 ( \64345 , \64343 , \64344 );
or \U$63969 ( \64346 , \397 , \64342 );
nand \U$63970 ( \64347 , \64345 , \64346 );
not \U$63971 ( \64348 , \64347 );
xor \U$63972 ( \64349 , \489 , \32458 );
xor \U$63973 ( \64350 , \32559 , \64336 );
and \U$63974 ( \64351 , \64349 , \64350 );
not \U$63975 ( \64352 , \64349 );
not \U$63976 ( \64353 , \64350 );
and \U$63977 ( \64354 , \64352 , \64353 );
xor \U$63978 ( \64355 , \32455 , \32440 );
xor \U$63979 ( \64356 , \64333 , \64318 );
and \U$63980 ( \64357 , \64355 , \64356 );
not \U$63981 ( \64358 , \64356 );
not \U$63982 ( \64359 , \64355 );
and \U$63983 ( \64360 , \64358 , \64359 );
xor \U$63984 ( \64361 , \32437 , \32418 );
xor \U$63985 ( \64362 , \64315 , \64296 );
and \U$63986 ( \64363 , \64361 , \64362 );
not \U$63987 ( \64364 , \64362 );
not \U$63988 ( \64365 , \64361 );
and \U$63989 ( \64366 , \64364 , \64365 );
xor \U$63990 ( \64367 , \32415 , \32372 );
xor \U$63991 ( \64368 , \32761 , \64294 );
and \U$63992 ( \64369 , \64367 , \64368 );
not \U$63993 ( \64370 , \64368 );
not \U$63994 ( \64371 , \64367 );
and \U$63995 ( \64372 , \64370 , \64371 );
xor \U$63996 ( \64373 , \768 , \32370 );
xor \U$63997 ( \64374 , \32855 , \64292 );
and \U$63998 ( \64375 , \64373 , \64374 );
not \U$63999 ( \64376 , \64374 );
not \U$64000 ( \64377 , \64373 );
and \U$64001 ( \64378 , \64376 , \64377 );
xor \U$64002 ( \64379 , \954 , \32368 );
xor \U$64003 ( \64380 , \33043 , \64290 );
and \U$64004 ( \64381 , \64379 , \64380 );
not \U$64005 ( \64382 , \64380 );
not \U$64006 ( \64383 , \64379 );
and \U$64007 ( \64384 , \64382 , \64383 );
and \U$64008 ( \64385 , \1081 , \32366 );
not \U$64009 ( \64386 , \1081 );
and \U$64010 ( \64387 , \64386 , \32365 );
nor \U$64011 ( \64388 , \64385 , \64387 );
xor \U$64012 ( \64389 , \33159 , \64288 );
and \U$64013 ( \64390 , \64388 , \64389 );
not \U$64014 ( \64391 , \64389 );
not \U$64015 ( \64392 , \64388 );
and \U$64016 ( \64393 , \64391 , \64392 );
xor \U$64017 ( \64394 , \32362 , \32358 );
xor \U$64018 ( \64395 , \64285 , \64277 );
and \U$64019 ( \64396 , \64394 , \64395 );
not \U$64020 ( \64397 , \64394 );
not \U$64021 ( \64398 , \64395 );
and \U$64022 ( \64399 , \64397 , \64398 );
xor \U$64023 ( \64400 , \1321 , \32356 );
xor \U$64024 ( \64401 , \64274 , \64258 );
and \U$64025 ( \64402 , \64400 , \64401 );
not \U$64026 ( \64403 , \64401 );
not \U$64027 ( \64404 , \64400 );
and \U$64028 ( \64405 , \64403 , \64404 );
xor \U$64029 ( \64406 , \1450 , \32354 );
xor \U$64030 ( \64407 , \64255 , \64224 );
and \U$64031 ( \64408 , \64406 , \64407 );
not \U$64032 ( \64409 , \64407 );
not \U$64033 ( \64410 , \64406 );
and \U$64034 ( \64411 , \64409 , \64410 );
xor \U$64035 ( \64412 , \64221 , \64181 );
xor \U$64036 ( \64413 , \32351 , \32343 );
and \U$64037 ( \64414 , \64412 , \64413 );
not \U$64038 ( \64415 , \64413 );
not \U$64039 ( \64416 , \64412 );
and \U$64040 ( \64417 , \64415 , \64416 );
xor \U$64041 ( \64418 , \64178 , \64114 );
xor \U$64042 ( \64419 , \1830 , \32341 );
and \U$64043 ( \64420 , \64418 , \64419 );
not \U$64044 ( \64421 , \64419 );
not \U$64045 ( \64422 , \64418 );
and \U$64046 ( \64423 , \64421 , \64422 );
xor \U$64047 ( \64424 , \33941 , \64112 );
xor \U$64048 ( \64425 , \2011 , \32339 );
and \U$64049 ( \64426 , \64424 , \64425 );
not \U$64050 ( \64427 , \64425 );
not \U$64051 ( \64428 , \64424 );
and \U$64052 ( \64429 , \64427 , \64428 );
xor \U$64053 ( \64430 , \34125 , \64110 );
xor \U$64054 ( \64431 , \2170 , \32337 );
and \U$64055 ( \64432 , \64430 , \64431 );
not \U$64056 ( \64433 , \64431 );
not \U$64057 ( \64434 , \64430 );
and \U$64058 ( \64435 , \64433 , \64434 );
xor \U$64059 ( \64436 , \34300 , \64108 );
xor \U$64060 ( \64437 , \32334 , \32326 );
and \U$64061 ( \64438 , \64436 , \64437 );
not \U$64062 ( \64439 , \64437 );
not \U$64063 ( \64440 , \64436 );
and \U$64064 ( \64441 , \64439 , \64440 );
xor \U$64065 ( \64442 , \32323 , \32307 );
xor \U$64066 ( \64443 , \34492 , \64106 );
and \U$64067 ( \64444 , \64442 , \64443 );
not \U$64068 ( \64445 , \64442 );
not \U$64069 ( \64446 , \64443 );
and \U$64070 ( \64447 , \64445 , \64446 );
xor \U$64071 ( \64448 , \2698 , \32305 );
xor \U$64072 ( \64449 , \34675 , \64104 );
and \U$64073 ( \64450 , \64448 , \64449 );
not \U$64074 ( \64451 , \64448 );
not \U$64075 ( \64452 , \64449 );
and \U$64076 ( \64453 , \64451 , \64452 );
xor \U$64077 ( \64454 , \32302 , \32294 );
xor \U$64078 ( \64455 , \64101 , \64093 );
and \U$64079 ( \64456 , \64454 , \64455 );
not \U$64080 ( \64457 , \64455 );
not \U$64081 ( \64458 , \64454 );
and \U$64082 ( \64459 , \64457 , \64458 );
xor \U$64083 ( \64460 , \32291 , \32277 );
xor \U$64084 ( \64461 , \64090 , \64076 );
and \U$64085 ( \64462 , \64460 , \64461 );
not \U$64086 ( \64463 , \64461 );
not \U$64087 ( \64464 , \64460 );
and \U$64088 ( \64465 , \64463 , \64464 );
xor \U$64089 ( \64466 , \32274 , \32247 );
xor \U$64090 ( \64467 , \35244 , \64074 );
and \U$64091 ( \64468 , \64466 , \64467 );
not \U$64092 ( \64469 , \64466 );
not \U$64093 ( \64470 , \64467 );
and \U$64094 ( \64471 , \64469 , \64470 );
xor \U$64095 ( \64472 , \32244 , \32197 );
xor \U$64096 ( \64473 , \35672 , \64072 );
and \U$64097 ( \64474 , \64472 , \64473 );
not \U$64098 ( \64475 , \64472 );
not \U$64099 ( \64476 , \64473 );
and \U$64100 ( \64477 , \64475 , \64476 );
xor \U$64101 ( \64478 , \32194 , \32113 );
xor \U$64102 ( \64479 , \35945 , \64070 );
and \U$64103 ( \64480 , \64478 , \64479 );
not \U$64104 ( \64481 , \64478 );
not \U$64105 ( \64482 , \64479 );
and \U$64106 ( \64483 , \64481 , \64482 );
xor \U$64107 ( \64484 , \4184 , \32111 );
xor \U$64108 ( \64485 , \64067 , \64059 );
and \U$64109 ( \64486 , \64484 , \64485 );
not \U$64110 ( \64487 , \64485 );
not \U$64111 ( \64488 , \64484 );
and \U$64112 ( \64489 , \64487 , \64488 );
xor \U$64113 ( \64490 , \4439 , \32109 );
xor \U$64114 ( \64491 , \64056 , \64038 );
and \U$64115 ( \64492 , \64490 , \64491 );
not \U$64116 ( \64493 , \64490 );
not \U$64117 ( \64494 , \64491 );
and \U$64118 ( \64495 , \64493 , \64494 );
xor \U$64119 ( \64496 , \32106 , \32098 );
xor \U$64120 ( \64497 , \64035 , \64000 );
and \U$64121 ( \64498 , \64496 , \64497 );
not \U$64122 ( \64499 , \64497 );
not \U$64123 ( \64500 , \64496 );
and \U$64124 ( \64501 , \64499 , \64500 );
not \U$64125 ( \64502 , \32095 );
not \U$64126 ( \64503 , \32081 );
or \U$64127 ( \64504 , \64502 , \64503 );
or \U$64128 ( \64505 , \32081 , \32095 );
nand \U$64129 ( \64506 , \64504 , \64505 );
xor \U$64130 ( \64507 , \36933 , \63998 );
and \U$64131 ( \64508 , \64506 , \64507 );
not \U$64132 ( \64509 , \64507 );
not \U$64133 ( \64510 , \64506 );
and \U$64134 ( \64511 , \64509 , \64510 );
xor \U$64135 ( \64512 , \5217 , \32079 );
xor \U$64136 ( \64513 , \37196 , \63996 );
and \U$64137 ( \64514 , \64512 , \64513 );
not \U$64138 ( \64515 , \64512 );
not \U$64139 ( \64516 , \64513 );
and \U$64140 ( \64517 , \64515 , \64516 );
xor \U$64141 ( \64518 , \5500 , \32077 );
xor \U$64142 ( \64519 , \63993 , \63985 );
and \U$64143 ( \64520 , \64518 , \64519 );
not \U$64144 ( \64521 , \64518 );
not \U$64145 ( \64522 , \64519 );
and \U$64146 ( \64523 , \64521 , \64522 );
xor \U$64147 ( \64524 , \5769 , \32075 );
xor \U$64148 ( \64525 , \63982 , \63965 );
and \U$64149 ( \64526 , \64524 , \64525 );
not \U$64150 ( \64527 , \64524 );
not \U$64151 ( \64528 , \64525 );
and \U$64152 ( \64529 , \64527 , \64528 );
xor \U$64153 ( \64530 , \6060 , \32073 );
xor \U$64154 ( \64531 , \63962 , \63929 );
and \U$64155 ( \64532 , \64530 , \64531 );
not \U$64156 ( \64533 , \64530 );
not \U$64157 ( \64534 , \64531 );
and \U$64158 ( \64535 , \64533 , \64534 );
xor \U$64159 ( \64536 , \32070 , \32063 );
xor \U$64160 ( \64537 , \63926 , \63893 );
and \U$64161 ( \64538 , \64536 , \64537 );
not \U$64162 ( \64539 , \64536 );
not \U$64163 ( \64540 , \64537 );
and \U$64164 ( \64541 , \64539 , \64540 );
xor \U$64165 ( \64542 , \63889 , \63830 );
xor \U$64166 ( \64543 , \32059 , \32045 );
and \U$64167 ( \64544 , \64542 , \64543 );
not \U$64168 ( \64545 , \64543 );
not \U$64169 ( \64546 , \64542 );
and \U$64170 ( \64547 , \64545 , \64546 );
and \U$64171 ( \64548 , \6926 , \32043 );
not \U$64172 ( \64549 , \6926 );
and \U$64173 ( \64550 , \64549 , \32042 );
nor \U$64174 ( \64551 , \64548 , \64550 );
not \U$64175 ( \64552 , \63827 );
not \U$64176 ( \64553 , \63730 );
or \U$64177 ( \64554 , \64552 , \64553 );
or \U$64178 ( \64555 , \63730 , \63827 );
nand \U$64179 ( \64556 , \64554 , \64555 );
and \U$64180 ( \64557 , \64551 , \64556 );
not \U$64181 ( \64558 , \64556 );
not \U$64182 ( \64559 , \64551 );
and \U$64183 ( \64560 , \64558 , \64559 );
and \U$64184 ( \64561 , \63727 , \63606 );
not \U$64185 ( \64562 , \63727 );
and \U$64186 ( \64563 , \64562 , \63605 );
nor \U$64187 ( \64564 , \64561 , \64563 );
not \U$64188 ( \64565 , \32039 );
not \U$64189 ( \64566 , \32031 );
or \U$64190 ( \64567 , \64565 , \64566 );
or \U$64191 ( \64568 , \32031 , \32039 );
nand \U$64192 ( \64569 , \64567 , \64568 );
and \U$64193 ( \64570 , \64564 , \64569 );
not \U$64194 ( \64571 , \64564 );
not \U$64195 ( \64572 , \64569 );
and \U$64196 ( \64573 , \64571 , \64572 );
and \U$64197 ( \64574 , \7865 , \32029 );
not \U$64198 ( \64575 , \7865 );
and \U$64199 ( \64576 , \64575 , \32028 );
nor \U$64200 ( \64577 , \64574 , \64576 );
xor \U$64201 ( \64578 , \63602 , \63326 );
and \U$64202 ( \64579 , \64577 , \64578 );
not \U$64203 ( \64580 , \64577 );
not \U$64204 ( \64581 , \64578 );
and \U$64205 ( \64582 , \64580 , \64581 );
xor \U$64206 ( \64583 , \8215 , \32026 );
xor \U$64207 ( \64584 , \39406 , \63324 );
and \U$64208 ( \64585 , \64583 , \64584 );
not \U$64209 ( \64586 , \64584 );
not \U$64210 ( \64587 , \64583 );
and \U$64211 ( \64588 , \64586 , \64587 );
xor \U$64212 ( \64589 , \8580 , \32024 );
xor \U$64213 ( \64590 , \39763 , \63322 );
and \U$64214 ( \64591 , \64589 , \64590 );
not \U$64215 ( \64592 , \64589 );
not \U$64216 ( \64593 , \64590 );
and \U$64217 ( \64594 , \64592 , \64593 );
xor \U$64218 ( \64595 , \32021 , \32013 );
xor \U$64219 ( \64596 , \40130 , \63320 );
and \U$64220 ( \64597 , \64595 , \64596 );
not \U$64221 ( \64598 , \64596 );
not \U$64222 ( \64599 , \64595 );
and \U$64223 ( \64600 , \64598 , \64599 );
xor \U$64224 ( \64601 , \32010 , \31991 );
xor \U$64225 ( \64602 , \40516 , \63318 );
and \U$64226 ( \64603 , \64601 , \64602 );
not \U$64227 ( \64604 , \64601 );
not \U$64228 ( \64605 , \64602 );
and \U$64229 ( \64606 , \64604 , \64605 );
not \U$64230 ( \64607 , \31988 );
not \U$64231 ( \64608 , \31966 );
or \U$64232 ( \64609 , \64607 , \64608 );
or \U$64233 ( \64610 , \31966 , \31988 );
nand \U$64234 ( \64611 , \64609 , \64610 );
xor \U$64235 ( \64612 , \40912 , \63316 );
and \U$64236 ( \64613 , \64611 , \64612 );
not \U$64237 ( \64614 , \64612 );
not \U$64238 ( \64615 , \64611 );
and \U$64239 ( \64616 , \64614 , \64615 );
xor \U$64240 ( \64617 , \10044 , \31964 );
xor \U$64241 ( \64618 , \63313 , \63305 );
and \U$64242 ( \64619 , \64617 , \64618 );
not \U$64243 ( \64620 , \64618 );
not \U$64244 ( \64621 , \64617 );
and \U$64245 ( \64622 , \64620 , \64621 );
xor \U$64246 ( \64623 , \31961 , \31953 );
xor \U$64247 ( \64624 , \41652 , \63303 );
and \U$64248 ( \64625 , \64623 , \64624 );
not \U$64249 ( \64626 , \64623 );
not \U$64250 ( \64627 , \64624 );
and \U$64251 ( \64628 , \64626 , \64627 );
not \U$64252 ( \64629 , \10818 );
not \U$64253 ( \64630 , \31950 );
or \U$64254 ( \64631 , \64629 , \64630 );
or \U$64255 ( \64632 , \31950 , \10818 );
nand \U$64256 ( \64633 , \64631 , \64632 );
xor \U$64257 ( \64634 , \63300 , \63293 );
and \U$64258 ( \64635 , \64633 , \64634 );
not \U$64259 ( \64636 , \64633 );
not \U$64260 ( \64637 , \64634 );
and \U$64261 ( \64638 , \64636 , \64637 );
xor \U$64262 ( \64639 , \11204 , \31948 );
xor \U$64263 ( \64640 , \63291 , \63290 );
and \U$64264 ( \64641 , \64639 , \64640 );
not \U$64265 ( \64642 , \64639 );
not \U$64266 ( \64643 , \64640 );
and \U$64267 ( \64644 , \64642 , \64643 );
xor \U$64268 ( \64645 , \31944 , \31936 );
xor \U$64269 ( \64646 , \42812 , \63288 );
and \U$64270 ( \64647 , \64645 , \64646 );
not \U$64271 ( \64648 , \64645 );
not \U$64272 ( \64649 , \64646 );
and \U$64273 ( \64650 , \64648 , \64649 );
xor \U$64274 ( \64651 , \12004 , \31934 );
xor \U$64275 ( \64652 , \43205 , \63286 );
and \U$64276 ( \64653 , \64651 , \64652 );
not \U$64277 ( \64654 , \64651 );
not \U$64278 ( \64655 , \64652 );
and \U$64279 ( \64656 , \64654 , \64655 );
xor \U$64280 ( \64657 , \31931 , \31923 );
xor \U$64281 ( \64658 , \43616 , \63284 );
and \U$64282 ( \64659 , \64657 , \64658 );
not \U$64283 ( \64660 , \64658 );
not \U$64284 ( \64661 , \64657 );
and \U$64285 ( \64662 , \64660 , \64661 );
xor \U$64286 ( \64663 , \12898 , \31921 );
xor \U$64287 ( \64664 , \63281 , \63273 );
and \U$64288 ( \64665 , \64663 , \64664 );
not \U$64289 ( \64666 , \64663 );
not \U$64290 ( \64667 , \64664 );
and \U$64291 ( \64668 , \64666 , \64667 );
xor \U$64292 ( \64669 , \31918 , \31910 );
xor \U$64293 ( \64670 , \44419 , \63271 );
and \U$64294 ( \64671 , \64669 , \64670 );
not \U$64295 ( \64672 , \64670 );
not \U$64296 ( \64673 , \64669 );
and \U$64297 ( \64674 , \64672 , \64673 );
and \U$64298 ( \64675 , \31907 , \31887 );
not \U$64299 ( \64676 , \31907 );
and \U$64300 ( \64677 , \64676 , \31886 );
nor \U$64301 ( \64678 , \64675 , \64677 );
xor \U$64302 ( \64679 , \63269 , \63268 );
and \U$64303 ( \64680 , \64678 , \64679 );
not \U$64304 ( \64681 , \64678 );
not \U$64305 ( \64682 , \64679 );
and \U$64306 ( \64683 , \64681 , \64682 );
xor \U$64307 ( \64684 , \31883 , \31854 );
xor \U$64308 ( \64685 , \45251 , \63266 );
and \U$64309 ( \64686 , \64684 , \64685 );
not \U$64310 ( \64687 , \64685 );
not \U$64311 ( \64688 , \64684 );
and \U$64312 ( \64689 , \64687 , \64688 );
xor \U$64313 ( \64690 , \14715 , \31852 );
xor \U$64314 ( \64691 , \45673 , \63264 );
and \U$64315 ( \64692 , \64690 , \64691 );
not \U$64316 ( \64693 , \64691 );
not \U$64317 ( \64694 , \64690 );
and \U$64318 ( \64695 , \64693 , \64694 );
xor \U$64319 ( \64696 , \15171 , \31850 );
xor \U$64320 ( \64697 , \63261 , \63251 );
and \U$64321 ( \64698 , \64696 , \64697 );
not \U$64322 ( \64699 , \64696 );
not \U$64323 ( \64700 , \64697 );
and \U$64324 ( \64701 , \64699 , \64700 );
xor \U$64325 ( \64702 , \31847 , \31834 );
xor \U$64326 ( \64703 , \63249 , \63248 );
and \U$64327 ( \64704 , \64702 , \64703 );
not \U$64328 ( \64705 , \64702 );
not \U$64329 ( \64706 , \64703 );
and \U$64330 ( \64707 , \64705 , \64706 );
xor \U$64331 ( \64708 , \31831 , \31807 );
xor \U$64332 ( \64709 , \47044 , \63246 );
and \U$64333 ( \64710 , \64708 , \64709 );
not \U$64334 ( \64711 , \64709 );
not \U$64335 ( \64712 , \64708 );
and \U$64336 ( \64713 , \64711 , \64712 );
xor \U$64337 ( \64714 , \31805 , \31804 );
xor \U$64338 ( \64715 , \63244 , \63243 );
and \U$64339 ( \64716 , \64714 , \64715 );
not \U$64340 ( \64717 , \64714 );
not \U$64341 ( \64718 , \64715 );
and \U$64342 ( \64719 , \64717 , \64718 );
xor \U$64343 ( \64720 , \17070 , \31802 );
xor \U$64344 ( \64721 , \48021 , \63241 );
and \U$64345 ( \64722 , \64720 , \64721 );
not \U$64346 ( \64723 , \64720 );
not \U$64347 ( \64724 , \64721 );
and \U$64348 ( \64725 , \64723 , \64724 );
xor \U$64349 ( \64726 , \31799 , \31786 );
xor \U$64350 ( \64727 , \63238 , \63225 );
and \U$64351 ( \64728 , \64726 , \64727 );
not \U$64352 ( \64729 , \64726 );
not \U$64353 ( \64730 , \64727 );
and \U$64354 ( \64731 , \64729 , \64730 );
xor \U$64355 ( \64732 , \31783 , \31757 );
xor \U$64356 ( \64733 , \63222 , \63198 );
and \U$64357 ( \64734 , \64732 , \64733 );
not \U$64358 ( \64735 , \64732 );
not \U$64359 ( \64736 , \64733 );
and \U$64360 ( \64737 , \64735 , \64736 );
xor \U$64361 ( \64738 , \31754 , \31703 );
xor \U$64362 ( \64739 , \63195 , \63153 );
and \U$64363 ( \64740 , \64738 , \64739 );
not \U$64364 ( \64741 , \64738 );
not \U$64365 ( \64742 , \64739 );
and \U$64366 ( \64743 , \64741 , \64742 );
xor \U$64367 ( \64744 , \18768 , \31701 );
xor \U$64368 ( \64745 , \49741 , \63151 );
and \U$64369 ( \64746 , \64744 , \64745 );
not \U$64370 ( \64747 , \64744 );
not \U$64371 ( \64748 , \64745 );
and \U$64372 ( \64749 , \64747 , \64748 );
xor \U$64373 ( \64750 , \19176 , \31699 );
xor \U$64374 ( \64751 , \63148 , \63139 );
and \U$64375 ( \64752 , \64750 , \64751 );
not \U$64376 ( \64753 , \64750 );
not \U$64377 ( \64754 , \64751 );
and \U$64378 ( \64755 , \64753 , \64754 );
xor \U$64379 ( \64756 , \31696 , \31684 );
xor \U$64380 ( \64757 , \50602 , \63137 );
and \U$64381 ( \64758 , \64756 , \64757 );
not \U$64382 ( \64759 , \64756 );
not \U$64383 ( \64760 , \64757 );
and \U$64384 ( \64761 , \64759 , \64760 );
xor \U$64385 ( \64762 , \31681 , \31660 );
xor \U$64386 ( \64763 , \51006 , \63135 );
and \U$64387 ( \64764 , \64762 , \64763 );
not \U$64388 ( \64765 , \64762 );
not \U$64389 ( \64766 , \64763 );
and \U$64390 ( \64767 , \64765 , \64766 );
xor \U$64391 ( \64768 , \20407 , \31658 );
xor \U$64392 ( \64769 , \63132 , \63124 );
and \U$64393 ( \64770 , \64768 , \64769 );
not \U$64394 ( \64771 , \64768 );
not \U$64395 ( \64772 , \64769 );
and \U$64396 ( \64773 , \64771 , \64772 );
xor \U$64397 ( \64774 , \31655 , \31645 );
xor \U$64398 ( \64775 , \63121 , \63105 );
and \U$64399 ( \64776 , \64774 , \64775 );
not \U$64400 ( \64777 , \64774 );
not \U$64401 ( \64778 , \64775 );
and \U$64402 ( \64779 , \64777 , \64778 );
xor \U$64403 ( \64780 , \31642 , \31626 );
xor \U$64404 ( \64781 , \63102 , \63070 );
and \U$64405 ( \64782 , \64780 , \64781 );
not \U$64406 ( \64783 , \64780 );
not \U$64407 ( \64784 , \64781 );
and \U$64408 ( \64785 , \64783 , \64784 );
xor \U$64409 ( \64786 , \31623 , \31583 );
xor \U$64410 ( \64787 , \52581 , \63068 );
and \U$64411 ( \64788 , \64786 , \64787 );
not \U$64412 ( \64789 , \64786 );
not \U$64413 ( \64790 , \64787 );
and \U$64414 ( \64791 , \64789 , \64790 );
xor \U$64415 ( \64792 , \21934 , \31581 );
xor \U$64416 ( \64793 , \63065 , \63057 );
and \U$64417 ( \64794 , \64792 , \64793 );
not \U$64418 ( \64795 , \64792 );
not \U$64419 ( \64796 , \64793 );
and \U$64420 ( \64797 , \64795 , \64796 );
xor \U$64421 ( \64798 , \21963 , \31579 );
xor \U$64422 ( \64799 , \53015 , \63055 );
and \U$64423 ( \64800 , \64798 , \64799 );
not \U$64424 ( \64801 , \64798 );
not \U$64425 ( \64802 , \64799 );
and \U$64426 ( \64803 , \64801 , \64802 );
xor \U$64427 ( \64804 , \31576 , \31564 );
xor \U$64428 ( \64805 , \53420 , \63053 );
and \U$64429 ( \64806 , \64804 , \64805 );
not \U$64430 ( \64807 , \64804 );
not \U$64431 ( \64808 , \64805 );
and \U$64432 ( \64809 , \64807 , \64808 );
xor \U$64433 ( \64810 , \22662 , \31562 );
xor \U$64434 ( \64811 , \63050 , \63039 );
and \U$64435 ( \64812 , \64810 , \64811 );
not \U$64436 ( \64813 , \64810 );
not \U$64437 ( \64814 , \64811 );
and \U$64438 ( \64815 , \64813 , \64814 );
xor \U$64439 ( \64816 , \23018 , \31560 );
xor \U$64440 ( \64817 , \63036 , \63014 );
and \U$64441 ( \64818 , \64816 , \64817 );
not \U$64442 ( \64819 , \64816 );
not \U$64443 ( \64820 , \64817 );
and \U$64444 ( \64821 , \64819 , \64820 );
xor \U$64445 ( \64822 , \23355 , \31558 );
xor \U$64446 ( \64823 , \63011 , \62978 );
and \U$64447 ( \64824 , \64822 , \64823 );
not \U$64448 ( \64825 , \64822 );
not \U$64449 ( \64826 , \64823 );
and \U$64450 ( \64827 , \64825 , \64826 );
xor \U$64451 ( \64828 , \31555 , \31546 );
xor \U$64452 ( \64829 , \62975 , \62918 );
and \U$64453 ( \64830 , \64828 , \64829 );
not \U$64454 ( \64831 , \64828 );
not \U$64455 ( \64832 , \64829 );
and \U$64456 ( \64833 , \64831 , \64832 );
xor \U$64457 ( \64834 , \24015 , \31544 );
xor \U$64458 ( \64835 , \62915 , \62830 );
and \U$64459 ( \64836 , \64834 , \64835 );
not \U$64460 ( \64837 , \64834 );
not \U$64461 ( \64838 , \64835 );
and \U$64462 ( \64839 , \64837 , \64838 );
xor \U$64463 ( \64840 , \31541 , \31532 );
xor \U$64464 ( \64841 , \62827 , \62696 );
and \U$64465 ( \64842 , \64840 , \64841 );
not \U$64466 ( \64843 , \64840 );
not \U$64467 ( \64844 , \64841 );
and \U$64468 ( \64845 , \64843 , \64844 );
xor \U$64469 ( \64846 , \24639 , \31530 );
xor \U$64470 ( \64847 , \62693 , \62504 );
and \U$64471 ( \64848 , \64846 , \64847 );
not \U$64472 ( \64849 , \64846 );
not \U$64473 ( \64850 , \64847 );
and \U$64474 ( \64851 , \64849 , \64850 );
xor \U$64475 ( \64852 , \31527 , \31518 );
xor \U$64476 ( \64853 , \62501 , \62122 );
and \U$64477 ( \64854 , \64852 , \64853 );
not \U$64478 ( \64855 , \64852 );
not \U$64479 ( \64856 , \64853 );
and \U$64480 ( \64857 , \64855 , \64856 );
xor \U$64481 ( \64858 , \31515 , \31497 );
xor \U$64482 ( \64859 , \62119 , \61756 );
and \U$64483 ( \64860 , \64858 , \64859 );
not \U$64484 ( \64861 , \64858 );
not \U$64485 ( \64862 , \64859 );
and \U$64486 ( \64863 , \64861 , \64862 );
xor \U$64487 ( \64864 , \25446 , \31495 );
xor \U$64488 ( \64865 , \61753 , \61418 );
and \U$64489 ( \64866 , \64864 , \64865 );
not \U$64490 ( \64867 , \64864 );
not \U$64491 ( \64868 , \64865 );
and \U$64492 ( \64869 , \64867 , \64868 );
xor \U$64493 ( \64870 , \25740 , \31493 );
xor \U$64494 ( \64871 , \55510 , \61416 );
and \U$64495 ( \64872 , \64870 , \64871 );
not \U$64496 ( \64873 , \64870 );
not \U$64497 ( \64874 , \64871 );
and \U$64498 ( \64875 , \64873 , \64874 );
xor \U$64499 ( \64876 , \31490 , \31481 );
xor \U$64500 ( \64877 , \61413 , \61404 );
and \U$64501 ( \64878 , \64876 , \64877 );
not \U$64502 ( \64879 , \64876 );
not \U$64503 ( \64880 , \64877 );
and \U$64504 ( \64881 , \64879 , \64880 );
xor \U$64505 ( \64882 , \31478 , \31459 );
xor \U$64506 ( \64883 , \61401 , \61382 );
and \U$64507 ( \64884 , \64882 , \64883 );
not \U$64508 ( \64885 , \64882 );
not \U$64509 ( \64886 , \64883 );
and \U$64510 ( \64887 , \64885 , \64886 );
xor \U$64511 ( \64888 , \26522 , \31457 );
xor \U$64512 ( \64889 , \56340 , \61380 );
and \U$64513 ( \64890 , \64888 , \64889 );
not \U$64514 ( \64891 , \64888 );
not \U$64515 ( \64892 , \64889 );
and \U$64516 ( \64893 , \64891 , \64892 );
xor \U$64517 ( \64894 , \26778 , \31455 );
xor \U$64518 ( \64895 , \61377 , \61368 );
and \U$64519 ( \64896 , \64894 , \64895 );
not \U$64520 ( \64897 , \64894 );
not \U$64521 ( \64898 , \64895 );
and \U$64522 ( \64899 , \64897 , \64898 );
xor \U$64523 ( \64900 , \31452 , \31444 );
xor \U$64524 ( \64901 , \61365 , \61347 );
and \U$64525 ( \64902 , \64900 , \64901 );
not \U$64526 ( \64903 , \64900 );
not \U$64527 ( \64904 , \64901 );
and \U$64528 ( \64905 , \64903 , \64904 );
xor \U$64529 ( \64906 , \27045 , \31442 );
xor \U$64530 ( \64907 , \56881 , \61345 );
and \U$64531 ( \64908 , \64906 , \64907 );
not \U$64532 ( \64909 , \64906 );
not \U$64533 ( \64910 , \64907 );
and \U$64534 ( \64911 , \64909 , \64910 );
xor \U$64535 ( \64912 , \31439 , \31427 );
xor \U$64536 ( \64913 , \57158 , \61343 );
and \U$64537 ( \64914 , \64912 , \64913 );
not \U$64538 ( \64915 , \64912 );
not \U$64539 ( \64916 , \64913 );
and \U$64540 ( \64917 , \64915 , \64916 );
xor \U$64541 ( \64918 , \27504 , \31425 );
xor \U$64542 ( \64919 , \57369 , \61341 );
and \U$64543 ( \64920 , \64918 , \64919 );
not \U$64544 ( \64921 , \64918 );
not \U$64545 ( \64922 , \64919 );
and \U$64546 ( \64923 , \64921 , \64922 );
xor \U$64547 ( \64924 , \31422 , \31412 );
xor \U$64548 ( \64925 , \57600 , \61339 );
and \U$64549 ( \64926 , \64924 , \64925 );
not \U$64550 ( \64927 , \64924 );
not \U$64551 ( \64928 , \64925 );
and \U$64552 ( \64929 , \64927 , \64928 );
xor \U$64553 ( \64930 , \31409 , \31384 );
xor \U$64554 ( \64931 , \61336 , \61321 );
and \U$64555 ( \64932 , \64930 , \64931 );
not \U$64556 ( \64933 , \64930 );
not \U$64557 ( \64934 , \64931 );
and \U$64558 ( \64935 , \64933 , \64934 );
xor \U$64559 ( \64936 , \28125 , \31382 );
xor \U$64560 ( \64937 , \58054 , \61319 );
and \U$64561 ( \64938 , \64936 , \64937 );
not \U$64562 ( \64939 , \64936 );
not \U$64563 ( \64940 , \64937 );
and \U$64564 ( \64941 , \64939 , \64940 );
xor \U$64565 ( \64942 , \28303 , \31380 );
xor \U$64566 ( \64943 , \61316 , \61301 );
and \U$64567 ( \64944 , \64942 , \64943 );
not \U$64568 ( \64945 , \64942 );
not \U$64569 ( \64946 , \64943 );
and \U$64570 ( \64947 , \64945 , \64946 );
xor \U$64571 ( \64948 , \28521 , \31378 );
xor \U$64572 ( \64949 , \61298 , \61281 );
and \U$64573 ( \64950 , \64948 , \64949 );
not \U$64574 ( \64951 , \64949 );
not \U$64575 ( \64952 , \64948 );
and \U$64576 ( \64953 , \64951 , \64952 );
xor \U$64577 ( \64954 , \28709 , \31376 );
xor \U$64578 ( \64955 , \61278 , \61248 );
and \U$64579 ( \64956 , \64954 , \64955 );
not \U$64580 ( \64957 , \64955 );
not \U$64581 ( \64958 , \64954 );
and \U$64582 ( \64959 , \64957 , \64958 );
xor \U$64583 ( \64960 , \31373 , \31364 );
xor \U$64584 ( \64961 , \61245 , \61185 );
and \U$64585 ( \64962 , \64960 , \64961 );
not \U$64586 ( \64963 , \64961 );
not \U$64587 ( \64964 , \64960 );
and \U$64588 ( \64965 , \64963 , \64964 );
xor \U$64589 ( \64966 , \29087 , \31362 );
xor \U$64590 ( \64967 , \58924 , \61183 );
and \U$64591 ( \64968 , \64966 , \64967 );
not \U$64592 ( \64969 , \64966 );
not \U$64593 ( \64970 , \64967 );
and \U$64594 ( \64971 , \64969 , \64970 );
xor \U$64595 ( \64972 , \31359 , \31354 );
xor \U$64596 ( \64973 , \61180 , \61175 );
and \U$64597 ( \64974 , \64972 , \64973 );
not \U$64598 ( \64975 , \64972 );
not \U$64599 ( \64976 , \64973 );
and \U$64600 ( \64977 , \64975 , \64976 );
xor \U$64601 ( \64978 , \29280 , \31352 );
xor \U$64602 ( \64979 , \59127 , \61173 );
and \U$64603 ( \64980 , \64978 , \64979 );
not \U$64604 ( \64981 , \64978 );
not \U$64605 ( \64982 , \64979 );
and \U$64606 ( \64983 , \64981 , \64982 );
xor \U$64607 ( \64984 , \29436 , \31350 );
xor \U$64608 ( \64985 , \61170 , \61158 );
and \U$64609 ( \64986 , \64984 , \64985 );
not \U$64610 ( \64987 , \64984 );
not \U$64611 ( \64988 , \64985 );
and \U$64612 ( \64989 , \64987 , \64988 );
xor \U$64613 ( \64990 , \29608 , \31348 );
xor \U$64614 ( \64991 , \59446 , \61156 );
and \U$64615 ( \64992 , \64990 , \64991 );
not \U$64616 ( \64993 , \64991 );
not \U$64617 ( \64994 , \64990 );
and \U$64618 ( \64995 , \64993 , \64994 );
xor \U$64619 ( \64996 , \29733 , \31346 );
xor \U$64620 ( \64997 , \59571 , \61154 );
and \U$64621 ( \64998 , \64996 , \64997 );
not \U$64622 ( \64999 , \64997 );
not \U$64623 ( \65000 , \64996 );
and \U$64624 ( \65001 , \64999 , \65000 );
xor \U$64625 ( \65002 , \29862 , \31344 );
xor \U$64626 ( \65003 , \59698 , \61152 );
and \U$64627 ( \65004 , \65002 , \65003 );
not \U$64628 ( \65005 , \65003 );
not \U$64629 ( \65006 , \65002 );
and \U$64630 ( \65007 , \65005 , \65006 );
xor \U$64631 ( \65008 , \31341 , \31332 );
xor \U$64632 ( \65009 , \61149 , \61140 );
and \U$64633 ( \65010 , \65008 , \65009 );
not \U$64634 ( \65011 , \65008 );
not \U$64635 ( \65012 , \65009 );
and \U$64636 ( \65013 , \65011 , \65012 );
xor \U$64637 ( \65014 , \31329 , \31311 );
xor \U$64638 ( \65015 , \61137 , \61119 );
and \U$64639 ( \65016 , \65014 , \65015 );
not \U$64640 ( \65017 , \65014 );
not \U$64641 ( \65018 , \65015 );
and \U$64642 ( \65019 , \65017 , \65018 );
xor \U$64643 ( \65020 , \31308 , \31285 );
xor \U$64644 ( \65021 , \61116 , \61090 );
and \U$64645 ( \65022 , \65020 , \65021 );
not \U$64646 ( \65023 , \65020 );
not \U$64647 ( \65024 , \65021 );
and \U$64648 ( \65025 , \65023 , \65024 );
xor \U$64649 ( \65026 , \61087 , \61031 );
xor \U$64650 ( \65027 , \30339 , \31283 );
and \U$64651 ( \65028 , \65026 , \65027 );
not \U$64652 ( \65029 , \65027 );
not \U$64653 ( \65030 , \65026 );
and \U$64654 ( \65031 , \65029 , \65030 );
xor \U$64655 ( \65032 , \61028 , \60948 );
xor \U$64656 ( \65033 , \30360 , \31281 );
and \U$64657 ( \65034 , \65032 , \65033 );
not \U$64658 ( \65035 , \65033 );
not \U$64659 ( \65036 , \65032 );
and \U$64660 ( \65037 , \65035 , \65036 );
xor \U$64661 ( \65038 , \60146 , \60946 );
xor \U$64662 ( \65039 , \30466 , \31279 );
and \U$64663 ( \65040 , \65038 , \65039 );
not \U$64664 ( \65041 , \65039 );
not \U$64665 ( \65042 , \65038 );
and \U$64666 ( \65043 , \65041 , \65042 );
xor \U$64667 ( \65044 , \60241 , \60944 );
xor \U$64668 ( \65045 , \31276 , \31259 );
and \U$64669 ( \65046 , \65044 , \65045 );
not \U$64670 ( \65047 , \65044 );
not \U$64671 ( \65048 , \65045 );
and \U$64672 ( \65049 , \65047 , \65048 );
xor \U$64673 ( \65050 , \31256 , \31225 );
xor \U$64674 ( \65051 , \60941 , \60926 );
and \U$64675 ( \65052 , \65050 , \65051 );
not \U$64676 ( \65053 , \65050 );
not \U$64677 ( \65054 , \65051 );
and \U$64678 ( \65055 , \65053 , \65054 );
xor \U$64679 ( \65056 , \30735 , \31223 );
xor \U$64680 ( \65057 , \60420 , \60924 );
and \U$64681 ( \65058 , \65056 , \65057 );
not \U$64682 ( \65059 , \65057 );
not \U$64683 ( \65060 , \65056 );
and \U$64684 ( \65061 , \65059 , \65060 );
xor \U$64685 ( \65062 , \31220 , \31207 );
xor \U$64686 ( \65063 , \60921 , \60912 );
and \U$64687 ( \65064 , \65062 , \65063 );
not \U$64688 ( \65065 , \65062 );
not \U$64689 ( \65066 , \65063 );
and \U$64690 ( \65067 , \65065 , \65066 );
xor \U$64691 ( \65068 , \60909 , \60893 );
xor \U$64692 ( \65069 , \31204 , \31190 );
and \U$64693 ( \65070 , \65068 , \65069 );
not \U$64694 ( \65071 , \65069 );
not \U$64695 ( \65072 , \65068 );
and \U$64696 ( \65073 , \65071 , \65072 );
xor \U$64697 ( \65074 , \30874 , \31188 );
xor \U$64698 ( \65075 , \60571 , \60891 );
and \U$64699 ( \65076 , \65074 , \65075 );
not \U$64700 ( \65077 , \65074 );
not \U$64701 ( \65078 , \65075 );
and \U$64702 ( \65079 , \65077 , \65078 );
xor \U$64703 ( \65080 , \60888 , \60875 );
xor \U$64704 ( \65081 , \31185 , \31173 );
and \U$64705 ( \65082 , \65080 , \65081 );
not \U$64706 ( \65083 , \65081 );
not \U$64707 ( \65084 , \65080 );
and \U$64708 ( \65085 , \65083 , \65084 );
xor \U$64709 ( \65086 , \60872 , \60844 );
xor \U$64710 ( \65087 , \31170 , \31150 );
and \U$64711 ( \65088 , \65086 , \65087 );
not \U$64712 ( \65089 , \65087 );
not \U$64713 ( \65090 , \65086 );
and \U$64714 ( \65091 , \65089 , \65090 );
xor \U$64715 ( \65092 , \60841 , \60809 );
xor \U$64716 ( \65093 , \31147 , \31120 );
and \U$64717 ( \65094 , \65092 , \65093 );
xor \U$64718 ( \65095 , \30938 , \30997 );
xor \U$64719 ( \65096 , \65095 , \31117 );
xor \U$64720 ( \65097 , \60635 , \60686 );
xor \U$64721 ( \65098 , \65097 , \60806 );
or \U$64722 ( \65099 , \65096 , \65098 );
xnor \U$64723 ( \65100 , \60803 , \60798 );
xnor \U$64724 ( \65101 , \31114 , \31101 );
or \U$64725 ( \65102 , \65100 , \65101 );
xor \U$64726 ( \65103 , \31098 , \31084 );
xor \U$64727 ( \65104 , \60795 , \60773 );
or \U$64728 ( \65105 , \65103 , \65104 );
nand \U$64729 ( \65106 , \65101 , \65100 );
xnor \U$64730 ( \65107 , \60770 , \60730 );
xnor \U$64731 ( \65108 , \31081 , \31041 );
and \U$64732 ( \65109 , \65107 , \65108 );
xor \U$64733 ( \65110 , \31078 , \31055 );
xor \U$64734 ( \65111 , \60767 , \60744 );
and \U$64735 ( \65112 , \65110 , \65111 );
not \U$64736 ( \65113 , \65110 );
not \U$64737 ( \65114 , \65111 );
and \U$64738 ( \65115 , \65113 , \65114 );
xor \U$64739 ( \65116 , \31075 , \31065 );
xor \U$64740 ( \65117 , \60764 , \60754 );
and \U$64741 ( \65118 , \65116 , \65117 );
not \U$64742 ( \65119 , \65116 );
not \U$64743 ( \65120 , \65117 );
and \U$64744 ( \65121 , \65119 , \65120 );
xor \U$64745 ( \65122 , \31067 , \31074 );
nor \U$64746 ( \65123 , \31066 , \60762 );
and \U$64747 ( \65124 , \65122 , \65123 );
and \U$64748 ( \65125 , \60761 , \60763 );
nor \U$64749 ( \65126 , \65122 , \65123 );
nor \U$64750 ( \65127 , \65125 , \65126 , \60764 );
nor \U$64751 ( \65128 , \65124 , \65127 );
nor \U$64752 ( \65129 , \65121 , \65128 );
nor \U$64753 ( \65130 , \65118 , \65129 );
nor \U$64754 ( \65131 , \65115 , \65130 );
nor \U$64755 ( \65132 , \65112 , \65131 );
or \U$64756 ( \65133 , \65109 , \65132 );
or \U$64757 ( \65134 , \65107 , \65108 );
nand \U$64758 ( \65135 , \65103 , \65104 );
nand \U$64759 ( \65136 , \65133 , \65134 , \65135 );
nand \U$64760 ( \65137 , \65105 , \65106 , \65136 );
nand \U$64761 ( \65138 , \65099 , \65102 , \65137 );
not \U$64762 ( \65139 , \65093 );
not \U$64763 ( \65140 , \65092 );
and \U$64764 ( \65141 , \65139 , \65140 );
and \U$64765 ( \65142 , \65098 , \65096 );
nor \U$64766 ( \65143 , \65141 , \65142 );
and \U$64767 ( \65144 , \65138 , \65143 );
nor \U$64768 ( \65145 , \65094 , \65144 );
nor \U$64769 ( \65146 , \65091 , \65145 );
nor \U$64770 ( \65147 , \65088 , \65146 );
nor \U$64771 ( \65148 , \65085 , \65147 );
nor \U$64772 ( \65149 , \65082 , \65148 );
nor \U$64773 ( \65150 , \65079 , \65149 );
nor \U$64774 ( \65151 , \65076 , \65150 );
nor \U$64775 ( \65152 , \65073 , \65151 );
nor \U$64776 ( \65153 , \65070 , \65152 );
nor \U$64777 ( \65154 , \65067 , \65153 );
nor \U$64778 ( \65155 , \65064 , \65154 );
nor \U$64779 ( \65156 , \65061 , \65155 );
nor \U$64780 ( \65157 , \65058 , \65156 );
nor \U$64781 ( \65158 , \65055 , \65157 );
nor \U$64782 ( \65159 , \65052 , \65158 );
nor \U$64783 ( \65160 , \65049 , \65159 );
nor \U$64784 ( \65161 , \65046 , \65160 );
nor \U$64785 ( \65162 , \65043 , \65161 );
nor \U$64786 ( \65163 , \65040 , \65162 );
nor \U$64787 ( \65164 , \65037 , \65163 );
nor \U$64788 ( \65165 , \65034 , \65164 );
nor \U$64789 ( \65166 , \65031 , \65165 );
nor \U$64790 ( \65167 , \65028 , \65166 );
nor \U$64791 ( \65168 , \65025 , \65167 );
nor \U$64792 ( \65169 , \65022 , \65168 );
nor \U$64793 ( \65170 , \65019 , \65169 );
nor \U$64794 ( \65171 , \65016 , \65170 );
nor \U$64795 ( \65172 , \65013 , \65171 );
nor \U$64796 ( \65173 , \65010 , \65172 );
nor \U$64797 ( \65174 , \65007 , \65173 );
nor \U$64798 ( \65175 , \65004 , \65174 );
nor \U$64799 ( \65176 , \65001 , \65175 );
nor \U$64800 ( \65177 , \64998 , \65176 );
nor \U$64801 ( \65178 , \64995 , \65177 );
nor \U$64802 ( \65179 , \64992 , \65178 );
nor \U$64803 ( \65180 , \64989 , \65179 );
nor \U$64804 ( \65181 , \64986 , \65180 );
nor \U$64805 ( \65182 , \64983 , \65181 );
nor \U$64806 ( \65183 , \64980 , \65182 );
nor \U$64807 ( \65184 , \64977 , \65183 );
nor \U$64808 ( \65185 , \64974 , \65184 );
nor \U$64809 ( \65186 , \64971 , \65185 );
nor \U$64810 ( \65187 , \64968 , \65186 );
nor \U$64811 ( \65188 , \64965 , \65187 );
nor \U$64812 ( \65189 , \64962 , \65188 );
nor \U$64813 ( \65190 , \64959 , \65189 );
nor \U$64814 ( \65191 , \64956 , \65190 );
nor \U$64815 ( \65192 , \64953 , \65191 );
nor \U$64816 ( \65193 , \64950 , \65192 );
nor \U$64817 ( \65194 , \64947 , \65193 );
nor \U$64818 ( \65195 , \64944 , \65194 );
nor \U$64819 ( \65196 , \64941 , \65195 );
nor \U$64820 ( \65197 , \64938 , \65196 );
nor \U$64821 ( \65198 , \64935 , \65197 );
nor \U$64822 ( \65199 , \64932 , \65198 );
nor \U$64823 ( \65200 , \64929 , \65199 );
nor \U$64824 ( \65201 , \64926 , \65200 );
nor \U$64825 ( \65202 , \64923 , \65201 );
nor \U$64826 ( \65203 , \64920 , \65202 );
nor \U$64827 ( \65204 , \64917 , \65203 );
nor \U$64828 ( \65205 , \64914 , \65204 );
nor \U$64829 ( \65206 , \64911 , \65205 );
nor \U$64830 ( \65207 , \64908 , \65206 );
nor \U$64831 ( \65208 , \64905 , \65207 );
nor \U$64832 ( \65209 , \64902 , \65208 );
nor \U$64833 ( \65210 , \64899 , \65209 );
nor \U$64834 ( \65211 , \64896 , \65210 );
nor \U$64835 ( \65212 , \64893 , \65211 );
nor \U$64836 ( \65213 , \64890 , \65212 );
nor \U$64837 ( \65214 , \64887 , \65213 );
nor \U$64838 ( \65215 , \64884 , \65214 );
nor \U$64839 ( \65216 , \64881 , \65215 );
nor \U$64840 ( \65217 , \64878 , \65216 );
nor \U$64841 ( \65218 , \64875 , \65217 );
nor \U$64842 ( \65219 , \64872 , \65218 );
nor \U$64843 ( \65220 , \64869 , \65219 );
nor \U$64844 ( \65221 , \64866 , \65220 );
nor \U$64845 ( \65222 , \64863 , \65221 );
nor \U$64846 ( \65223 , \64860 , \65222 );
nor \U$64847 ( \65224 , \64857 , \65223 );
nor \U$64848 ( \65225 , \64854 , \65224 );
nor \U$64849 ( \65226 , \64851 , \65225 );
nor \U$64850 ( \65227 , \64848 , \65226 );
nor \U$64851 ( \65228 , \64845 , \65227 );
nor \U$64852 ( \65229 , \64842 , \65228 );
nor \U$64853 ( \65230 , \64839 , \65229 );
nor \U$64854 ( \65231 , \64836 , \65230 );
nor \U$64855 ( \65232 , \64833 , \65231 );
nor \U$64856 ( \65233 , \64830 , \65232 );
nor \U$64857 ( \65234 , \64827 , \65233 );
nor \U$64858 ( \65235 , \64824 , \65234 );
nor \U$64859 ( \65236 , \64821 , \65235 );
nor \U$64860 ( \65237 , \64818 , \65236 );
nor \U$64861 ( \65238 , \64815 , \65237 );
nor \U$64862 ( \65239 , \64812 , \65238 );
nor \U$64863 ( \65240 , \64809 , \65239 );
nor \U$64864 ( \65241 , \64806 , \65240 );
nor \U$64865 ( \65242 , \64803 , \65241 );
nor \U$64866 ( \65243 , \64800 , \65242 );
nor \U$64867 ( \65244 , \64797 , \65243 );
nor \U$64868 ( \65245 , \64794 , \65244 );
nor \U$64869 ( \65246 , \64791 , \65245 );
nor \U$64870 ( \65247 , \64788 , \65246 );
nor \U$64871 ( \65248 , \64785 , \65247 );
nor \U$64872 ( \65249 , \64782 , \65248 );
nor \U$64873 ( \65250 , \64779 , \65249 );
nor \U$64874 ( \65251 , \64776 , \65250 );
nor \U$64875 ( \65252 , \64773 , \65251 );
nor \U$64876 ( \65253 , \64770 , \65252 );
nor \U$64877 ( \65254 , \64767 , \65253 );
nor \U$64878 ( \65255 , \64764 , \65254 );
nor \U$64879 ( \65256 , \64761 , \65255 );
nor \U$64880 ( \65257 , \64758 , \65256 );
nor \U$64881 ( \65258 , \64755 , \65257 );
nor \U$64882 ( \65259 , \64752 , \65258 );
nor \U$64883 ( \65260 , \64749 , \65259 );
nor \U$64884 ( \65261 , \64746 , \65260 );
nor \U$64885 ( \65262 , \64743 , \65261 );
nor \U$64886 ( \65263 , \64740 , \65262 );
nor \U$64887 ( \65264 , \64737 , \65263 );
nor \U$64888 ( \65265 , \64734 , \65264 );
nor \U$64889 ( \65266 , \64731 , \65265 );
nor \U$64890 ( \65267 , \64728 , \65266 );
nor \U$64891 ( \65268 , \64725 , \65267 );
nor \U$64892 ( \65269 , \64722 , \65268 );
nor \U$64893 ( \65270 , \64719 , \65269 );
nor \U$64894 ( \65271 , \64716 , \65270 );
nor \U$64895 ( \65272 , \64713 , \65271 );
nor \U$64896 ( \65273 , \64710 , \65272 );
nor \U$64897 ( \65274 , \64707 , \65273 );
nor \U$64898 ( \65275 , \64704 , \65274 );
nor \U$64899 ( \65276 , \64701 , \65275 );
nor \U$64900 ( \65277 , \64698 , \65276 );
nor \U$64901 ( \65278 , \64695 , \65277 );
nor \U$64902 ( \65279 , \64692 , \65278 );
nor \U$64903 ( \65280 , \64689 , \65279 );
nor \U$64904 ( \65281 , \64686 , \65280 );
nor \U$64905 ( \65282 , \64683 , \65281 );
nor \U$64906 ( \65283 , \64680 , \65282 );
nor \U$64907 ( \65284 , \64674 , \65283 );
nor \U$64908 ( \65285 , \64671 , \65284 );
nor \U$64909 ( \65286 , \64668 , \65285 );
nor \U$64910 ( \65287 , \64665 , \65286 );
nor \U$64911 ( \65288 , \64662 , \65287 );
nor \U$64912 ( \65289 , \64659 , \65288 );
nor \U$64913 ( \65290 , \64656 , \65289 );
nor \U$64914 ( \65291 , \64653 , \65290 );
nor \U$64915 ( \65292 , \64650 , \65291 );
nor \U$64916 ( \65293 , \64647 , \65292 );
nor \U$64917 ( \65294 , \64644 , \65293 );
nor \U$64918 ( \65295 , \64641 , \65294 );
nor \U$64919 ( \65296 , \64638 , \65295 );
nor \U$64920 ( \65297 , \64635 , \65296 );
nor \U$64921 ( \65298 , \64628 , \65297 );
nor \U$64922 ( \65299 , \64625 , \65298 );
nor \U$64923 ( \65300 , \64622 , \65299 );
nor \U$64924 ( \65301 , \64619 , \65300 );
nor \U$64925 ( \65302 , \64616 , \65301 );
nor \U$64926 ( \65303 , \64613 , \65302 );
nor \U$64927 ( \65304 , \64606 , \65303 );
nor \U$64928 ( \65305 , \64603 , \65304 );
nor \U$64929 ( \65306 , \64600 , \65305 );
nor \U$64930 ( \65307 , \64597 , \65306 );
nor \U$64931 ( \65308 , \64594 , \65307 );
nor \U$64932 ( \65309 , \64591 , \65308 );
nor \U$64933 ( \65310 , \64588 , \65309 );
nor \U$64934 ( \65311 , \64585 , \65310 );
nor \U$64935 ( \65312 , \64582 , \65311 );
nor \U$64936 ( \65313 , \64579 , \65312 );
nor \U$64937 ( \65314 , \64573 , \65313 );
nor \U$64938 ( \65315 , \64570 , \65314 );
nor \U$64939 ( \65316 , \64560 , \65315 );
nor \U$64940 ( \65317 , \64557 , \65316 );
nor \U$64941 ( \65318 , \64547 , \65317 );
nor \U$64942 ( \65319 , \64544 , \65318 );
nor \U$64943 ( \65320 , \64541 , \65319 );
nor \U$64944 ( \65321 , \64538 , \65320 );
nor \U$64945 ( \65322 , \64535 , \65321 );
nor \U$64946 ( \65323 , \64532 , \65322 );
nor \U$64947 ( \65324 , \64529 , \65323 );
nor \U$64948 ( \65325 , \64526 , \65324 );
nor \U$64949 ( \65326 , \64523 , \65325 );
nor \U$64950 ( \65327 , \64520 , \65326 );
nor \U$64951 ( \65328 , \64517 , \65327 );
nor \U$64952 ( \65329 , \64514 , \65328 );
nor \U$64953 ( \65330 , \64511 , \65329 );
nor \U$64954 ( \65331 , \64508 , \65330 );
nor \U$64955 ( \65332 , \64501 , \65331 );
nor \U$64956 ( \65333 , \64498 , \65332 );
nor \U$64957 ( \65334 , \64495 , \65333 );
nor \U$64958 ( \65335 , \64492 , \65334 );
nor \U$64959 ( \65336 , \64489 , \65335 );
nor \U$64960 ( \65337 , \64486 , \65336 );
nor \U$64961 ( \65338 , \64483 , \65337 );
nor \U$64962 ( \65339 , \64480 , \65338 );
nor \U$64963 ( \65340 , \64477 , \65339 );
nor \U$64964 ( \65341 , \64474 , \65340 );
nor \U$64965 ( \65342 , \64471 , \65341 );
nor \U$64966 ( \65343 , \64468 , \65342 );
nor \U$64967 ( \65344 , \64465 , \65343 );
nor \U$64968 ( \65345 , \64462 , \65344 );
nor \U$64969 ( \65346 , \64459 , \65345 );
nor \U$64970 ( \65347 , \64456 , \65346 );
nor \U$64971 ( \65348 , \64453 , \65347 );
nor \U$64972 ( \65349 , \64450 , \65348 );
nor \U$64973 ( \65350 , \64447 , \65349 );
nor \U$64974 ( \65351 , \64444 , \65350 );
nor \U$64975 ( \65352 , \64441 , \65351 );
nor \U$64976 ( \65353 , \64438 , \65352 );
nor \U$64977 ( \65354 , \64435 , \65353 );
nor \U$64978 ( \65355 , \64432 , \65354 );
nor \U$64979 ( \65356 , \64429 , \65355 );
nor \U$64980 ( \65357 , \64426 , \65356 );
nor \U$64981 ( \65358 , \64423 , \65357 );
nor \U$64982 ( \65359 , \64420 , \65358 );
nor \U$64983 ( \65360 , \64417 , \65359 );
nor \U$64984 ( \65361 , \64414 , \65360 );
nor \U$64985 ( \65362 , \64411 , \65361 );
nor \U$64986 ( \65363 , \64408 , \65362 );
nor \U$64987 ( \65364 , \64405 , \65363 );
nor \U$64988 ( \65365 , \64402 , \65364 );
nor \U$64989 ( \65366 , \64399 , \65365 );
nor \U$64990 ( \65367 , \64396 , \65366 );
nor \U$64991 ( \65368 , \64393 , \65367 );
nor \U$64992 ( \65369 , \64390 , \65368 );
nor \U$64993 ( \65370 , \64384 , \65369 );
nor \U$64994 ( \65371 , \64381 , \65370 );
nor \U$64995 ( \65372 , \64378 , \65371 );
nor \U$64996 ( \65373 , \64375 , \65372 );
nor \U$64997 ( \65374 , \64372 , \65373 );
nor \U$64998 ( \65375 , \64369 , \65374 );
nor \U$64999 ( \65376 , \64366 , \65375 );
nor \U$65000 ( \65377 , \64363 , \65376 );
nor \U$65001 ( \65378 , \64360 , \65377 );
nor \U$65002 ( \65379 , \64357 , \65378 );
nor \U$65003 ( \65380 , \64354 , \65379 );
nor \U$65004 ( \65381 , \64351 , \65380 );
not \U$65005 ( \65382 , \65381 );
or \U$65006 ( \65383 , \64348 , \65382 );
or \U$65007 ( \65384 , \65381 , \64347 );
nand \U$65008 ( \65385 , \65383 , \65384 );
not \U$65009 ( \65386 , \65385 );
or \U$65010 ( \65387 , \64341 , \65386 );
or \U$65011 ( \65388 , \65385 , \64340 );
nand \U$65012 ( \65389 , \65387 , \65388 );
not \U$65013 ( \65390 , \65389 );
or \U$65014 ( \65391 , \32482 , \65390 );
or \U$65015 ( \65392 , \65389 , \32481 );
nand \U$65016 ( \65393 , \65391 , \65392 );
xnor \U$65017 ( \65394 , RIae7c8b0_256, RIae7bfc8_237);
not \U$65018 ( \65395 , \65394 );
xor \U$65019 ( \65396 , RIae7c298_243, RIae7c838_255);
not \U$65020 ( \65397 , \65396 );
and \U$65021 ( \65398 , \65395 , \65397 );
and \U$65022 ( \65399 , \65394 , \65396 );
nor \U$65023 ( \65400 , \65398 , \65399 );
not \U$65024 ( \65401 , \65400 );
xor \U$65025 ( \65402 , RIae7b9b0_224, RIae7ab28_193);
not \U$65026 ( \65403 , \65402 );
xnor \U$65027 ( \65404 , RIae7b398_211, RIae7c658_251);
not \U$65028 ( \65405 , \65404 );
or \U$65029 ( \65406 , \65403 , \65405 );
or \U$65030 ( \65407 , \65404 , \65402 );
nand \U$65031 ( \65408 , \65406 , \65407 );
not \U$65032 ( \65409 , \65408 );
and \U$65033 ( \65410 , \65401 , \65409 );
and \U$65034 ( \65411 , \65400 , \65408 );
nor \U$65035 ( \65412 , \65410 , \65411 );
not \U$65036 ( \65413 , \65412 );
xor \U$65037 ( \65414 , RIae7b578_215, RIae7b6e0_218);
not \U$65038 ( \65415 , \65414 );
xnor \U$65039 ( \65416 , RIae7b2a8_209, RIae7bf50_236);
not \U$65040 ( \65417 , \65416 );
or \U$65041 ( \65418 , \65415 , \65417 );
or \U$65042 ( \65419 , \65416 , \65414 );
nand \U$65043 ( \65420 , \65418 , \65419 );
not \U$65044 ( \65421 , \65420 );
xnor \U$65045 ( \65422 , RIae7b848_221, RIae7b938_223);
not \U$65046 ( \65423 , \65422 );
xor \U$65047 ( \65424 , RIae7bb90_228, RIae7afd8_203);
not \U$65048 ( \65425 , \65424 );
and \U$65049 ( \65426 , \65423 , \65425 );
and \U$65050 ( \65427 , \65422 , \65424 );
nor \U$65051 ( \65428 , \65426 , \65427 );
not \U$65052 ( \65429 , \65428 );
or \U$65053 ( \65430 , \65421 , \65429 );
or \U$65054 ( \65431 , \65428 , \65420 );
nand \U$65055 ( \65432 , \65430 , \65431 );
not \U$65056 ( \65433 , \65432 );
and \U$65057 ( \65434 , \65413 , \65433 );
and \U$65058 ( \65435 , \65412 , \65432 );
nor \U$65059 ( \65436 , \65434 , \65435 );
not \U$65060 ( \65437 , \65436 );
xor \U$65061 ( \65438 , RIae7c7c0_254, RIae7bc80_230);
not \U$65062 ( \65439 , \65438 );
xnor \U$65063 ( \65440 , RIae7b8c0_222, RIae7b500_214);
not \U$65064 ( \65441 , \65440 );
or \U$65065 ( \65442 , \65439 , \65441 );
or \U$65066 ( \65443 , \65440 , \65438 );
nand \U$65067 ( \65444 , \65442 , \65443 );
not \U$65068 ( \65445 , \65444 );
xnor \U$65069 ( \65446 , RIae7b410_212, RIae7c400_246);
not \U$65070 ( \65447 , \65446 );
xor \U$65071 ( \65448 , RIae7be60_234, RIae7c130_240);
not \U$65072 ( \65449 , \65448 );
and \U$65073 ( \65450 , \65447 , \65449 );
and \U$65074 ( \65451 , \65446 , \65448 );
nor \U$65075 ( \65452 , \65450 , \65451 );
not \U$65076 ( \65453 , \65452 );
or \U$65077 ( \65454 , \65445 , \65453 );
or \U$65078 ( \65455 , \65452 , \65444 );
nand \U$65079 ( \65456 , \65454 , \65455 );
not \U$65080 ( \65457 , \65456 );
xnor \U$65081 ( \65458 , RIae7c310_244, RIae7c568_249);
not \U$65082 ( \65459 , \65458 );
xor \U$65083 ( \65460 , RIae7aba0_194, RIae7c6d0_252);
not \U$65084 ( \65461 , \65460 );
and \U$65085 ( \65462 , \65459 , \65461 );
and \U$65086 ( \65463 , \65458 , \65460 );
nor \U$65087 ( \65464 , \65462 , \65463 );
not \U$65088 ( \65465 , \65464 );
xor \U$65089 ( \65466 , RIae7ad80_198, RIae7b140_206);
not \U$65090 ( \65467 , \65466 );
xnor \U$65091 ( \65468 , RIae7b050_204, RIae7c0b8_239);
not \U$65092 ( \65469 , \65468 );
or \U$65093 ( \65470 , \65467 , \65469 );
or \U$65094 ( \65471 , \65468 , \65466 );
nand \U$65095 ( \65472 , \65470 , \65471 );
not \U$65096 ( \65473 , \65472 );
and \U$65097 ( \65474 , \65465 , \65473 );
and \U$65098 ( \65475 , \65464 , \65472 );
nor \U$65099 ( \65476 , \65474 , \65475 );
not \U$65100 ( \65477 , \65476 );
or \U$65101 ( \65478 , \65457 , \65477 );
or \U$65102 ( \65479 , \65476 , \65456 );
nand \U$65103 ( \65480 , \65478 , \65479 );
not \U$65104 ( \65481 , \65480 );
or \U$65105 ( \65482 , \65437 , \65481 );
or \U$65106 ( \65483 , \65436 , \65480 );
nand \U$65107 ( \65484 , \65482 , \65483 );
xnor \U$65108 ( \65485 , RIae7bc08_229, RIae7c748_253);
not \U$65109 ( \65486 , \65485 );
xor \U$65110 ( \65487 , RIae7c388_245, RIae7b488_213);
not \U$65111 ( \65488 , \65487 );
and \U$65112 ( \65489 , \65486 , \65488 );
and \U$65113 ( \65490 , \65485 , \65487 );
nor \U$65114 ( \65491 , \65489 , \65490 );
not \U$65115 ( \65492 , \65491 );
xor \U$65116 ( \65493 , RIae7b5f0_216, RIae7ac90_196);
not \U$65117 ( \65494 , \65493 );
xnor \U$65118 ( \65495 , RIae7c040_238, RIae7c5e0_250);
not \U$65119 ( \65496 , \65495 );
or \U$65120 ( \65497 , \65494 , \65496 );
or \U$65121 ( \65498 , \65495 , \65493 );
nand \U$65122 ( \65499 , \65497 , \65498 );
not \U$65123 ( \65500 , \65499 );
and \U$65124 ( \65501 , \65492 , \65500 );
and \U$65125 ( \65502 , \65491 , \65499 );
nor \U$65126 ( \65503 , \65501 , \65502 );
not \U$65127 ( \65504 , \65503 );
xor \U$65128 ( \65505 , RIae7c478_247, RIae7b320_210);
not \U$65129 ( \65506 , \65505 );
xnor \U$65130 ( \65507 , RIae7adf8_199, RIae7af60_202);
not \U$65131 ( \65508 , \65507 );
or \U$65132 ( \65509 , \65506 , \65508 );
or \U$65133 ( \65510 , \65507 , \65505 );
nand \U$65134 ( \65511 , \65509 , \65510 );
not \U$65135 ( \65512 , \65511 );
xnor \U$65136 ( \65513 , RIae7b758_219, RIae7bcf8_231);
not \U$65137 ( \65514 , \65513 );
xor \U$65138 ( \65515 , RIae7b668_217, RIae7ad08_197);
not \U$65139 ( \65516 , \65515 );
and \U$65140 ( \65517 , \65514 , \65516 );
and \U$65141 ( \65518 , \65513 , \65515 );
nor \U$65142 ( \65519 , \65517 , \65518 );
not \U$65143 ( \65520 , \65519 );
or \U$65144 ( \65521 , \65512 , \65520 );
or \U$65145 ( \65522 , \65519 , \65511 );
nand \U$65146 ( \65523 , \65521 , \65522 );
not \U$65147 ( \65524 , \65523 );
and \U$65148 ( \65525 , \65504 , \65524 );
and \U$65149 ( \65526 , \65503 , \65523 );
nor \U$65150 ( \65527 , \65525 , \65526 );
not \U$65151 ( \65528 , \65527 );
xor \U$65152 ( \65529 , RIae7ac18_195, RIae7bd70_232);
not \U$65153 ( \65530 , \65529 );
xnor \U$65154 ( \65531 , RIae7b7d0_220, RIae7aee8_201);
not \U$65155 ( \65532 , \65531 );
or \U$65156 ( \65533 , \65530 , \65532 );
or \U$65157 ( \65534 , \65531 , \65529 );
nand \U$65158 ( \65535 , \65533 , \65534 );
not \U$65159 ( \65536 , \65535 );
xnor \U$65160 ( \65537 , RIae7c1a8_241, RIae7b1b8_207);
not \U$65161 ( \65538 , \65537 );
xor \U$65162 ( \65539 , RIae7ae70_200, RIae7c4f0_248);
not \U$65163 ( \65540 , \65539 );
and \U$65164 ( \65541 , \65538 , \65540 );
and \U$65165 ( \65542 , \65537 , \65539 );
nor \U$65166 ( \65543 , \65541 , \65542 );
not \U$65167 ( \65544 , \65543 );
or \U$65168 ( \65545 , \65536 , \65544 );
or \U$65169 ( \65546 , \65543 , \65535 );
nand \U$65170 ( \65547 , \65545 , \65546 );
not \U$65171 ( \65548 , \65547 );
xnor \U$65172 ( \65549 , RIae7bde8_233, RIae7c220_242);
not \U$65173 ( \65550 , \65549 );
xor \U$65174 ( \65551 , RIae7bed8_235, RIae7b0c8_205);
not \U$65175 ( \65552 , \65551 );
and \U$65176 ( \65553 , \65550 , \65552 );
and \U$65177 ( \65554 , \65549 , \65551 );
nor \U$65178 ( \65555 , \65553 , \65554 );
not \U$65179 ( \65556 , \65555 );
xor \U$65180 ( \65557 , RIae7bb18_227, RIae7ba28_225);
not \U$65181 ( \65558 , \65557 );
xnor \U$65182 ( \65559 , RIae7baa0_226, RIae7b230_208);
not \U$65183 ( \65560 , \65559 );
or \U$65184 ( \65561 , \65558 , \65560 );
or \U$65185 ( \65562 , \65559 , \65557 );
nand \U$65186 ( \65563 , \65561 , \65562 );
not \U$65187 ( \65564 , \65563 );
and \U$65188 ( \65565 , \65556 , \65564 );
and \U$65189 ( \65566 , \65555 , \65563 );
nor \U$65190 ( \65567 , \65565 , \65566 );
not \U$65191 ( \65568 , \65567 );
or \U$65192 ( \65569 , \65548 , \65568 );
or \U$65193 ( \65570 , \65567 , \65547 );
nand \U$65194 ( \65571 , \65569 , \65570 );
not \U$65195 ( \65572 , \65571 );
and \U$65196 ( \65573 , \65528 , \65572 );
and \U$65197 ( \65574 , \65527 , \65571 );
nor \U$65198 ( \65575 , \65573 , \65574 );
not \U$65199 ( \65576 , \65575 );
and \U$65200 ( \65577 , \65484 , \65576 );
not \U$65201 ( \65578 , \65484 );
and \U$65202 ( \65579 , \65578 , \65575 );
or \U$65203 ( \65580 , \65577 , \65579 );
_DC g10344 ( \65581_nG10344 , \65393 , \65580 );
buf \U$65204 ( \65582 , \65581_nG10344 );
not \U$65205 ( \65583 , \65379 );
xor \U$65206 ( \65584 , \64350 , \64349 );
not \U$65207 ( \65585 , \65584 );
or \U$65208 ( \65586 , \65583 , \65585 );
or \U$65209 ( \65587 , \65584 , \65379 );
nand \U$65210 ( \65588 , \65586 , \65587 );
_DC g10315 ( \65589_nG10315 , \65588 , \65580 );
buf \U$65211 ( \65590 , \65589_nG10315 );
not \U$65212 ( \65591 , \65377 );
xor \U$65213 ( \65592 , \64355 , \64356 );
not \U$65214 ( \65593 , \65592 );
or \U$65215 ( \65594 , \65591 , \65593 );
or \U$65216 ( \65595 , \65592 , \65377 );
nand \U$65217 ( \65596 , \65594 , \65595 );
_DC g102d0 ( \65597_nG102d0 , \65596 , \65580 );
buf \U$65218 ( \65598 , \65597_nG102d0 );
not \U$65219 ( \65599 , \65375 );
xor \U$65220 ( \65600 , \64361 , \64362 );
not \U$65221 ( \65601 , \65600 );
or \U$65222 ( \65602 , \65599 , \65601 );
or \U$65223 ( \65603 , \65600 , \65375 );
nand \U$65224 ( \65604 , \65602 , \65603 );
_DC g1026f ( \65605_nG1026f , \65604 , \65580 );
buf \U$65225 ( \65606 , \65605_nG1026f );
not \U$65226 ( \65607 , \65373 );
xor \U$65227 ( \65608 , \64367 , \64368 );
not \U$65228 ( \65609 , \65608 );
or \U$65229 ( \65610 , \65607 , \65609 );
or \U$65230 ( \65611 , \65608 , \65373 );
nand \U$65231 ( \65612 , \65610 , \65611 );
_DC g10201 ( \65613_nG10201 , \65612 , \65580 );
buf \U$65232 ( \65614 , \65613_nG10201 );
not \U$65233 ( \65615 , \65371 );
xor \U$65234 ( \65616 , \64373 , \64374 );
not \U$65235 ( \65617 , \65616 );
or \U$65236 ( \65618 , \65615 , \65617 );
or \U$65237 ( \65619 , \65616 , \65371 );
nand \U$65238 ( \65620 , \65618 , \65619 );
_DC g10176 ( \65621_nG10176 , \65620 , \65580 );
buf \U$65239 ( \65622 , \65621_nG10176 );
not \U$65240 ( \65623 , \65369 );
xor \U$65241 ( \65624 , \64380 , \64379 );
not \U$65242 ( \65625 , \65624 );
or \U$65243 ( \65626 , \65623 , \65625 );
or \U$65244 ( \65627 , \65624 , \65369 );
nand \U$65245 ( \65628 , \65626 , \65627 );
_DC g100f9 ( \65629_nG100f9 , \65628 , \65580 );
buf \U$65246 ( \65630 , \65629_nG100f9 );
not \U$65247 ( \65631 , \65367 );
xor \U$65248 ( \65632 , \64388 , \64389 );
not \U$65249 ( \65633 , \65632 );
or \U$65250 ( \65634 , \65631 , \65633 );
or \U$65251 ( \65635 , \65632 , \65367 );
nand \U$65252 ( \65636 , \65634 , \65635 );
_DC g1005e ( \65637_nG1005e , \65636 , \65580 );
buf \U$65253 ( \65638 , \65637_nG1005e );
not \U$65254 ( \65639 , \65365 );
xor \U$65255 ( \65640 , \64395 , \64394 );
not \U$65256 ( \65641 , \65640 );
or \U$65257 ( \65642 , \65639 , \65641 );
or \U$65258 ( \65643 , \65640 , \65365 );
nand \U$65259 ( \65644 , \65642 , \65643 );
_DC gff9a ( \65645_nGff9a , \65644 , \65580 );
buf \U$65260 ( \65646 , \65645_nGff9a );
not \U$65261 ( \65647 , \65363 );
xor \U$65262 ( \65648 , \64400 , \64401 );
not \U$65263 ( \65649 , \65648 );
or \U$65264 ( \65650 , \65647 , \65649 );
or \U$65265 ( \65651 , \65648 , \65363 );
nand \U$65266 ( \65652 , \65650 , \65651 );
_DC gfed3 ( \65653_nGfed3 , \65652 , \65580 );
buf \U$65267 ( \65654 , \65653_nGfed3 );
not \U$65268 ( \65655 , \65361 );
xor \U$65269 ( \65656 , \64407 , \64406 );
not \U$65270 ( \65657 , \65656 );
or \U$65271 ( \65658 , \65655 , \65657 );
or \U$65272 ( \65659 , \65656 , \65361 );
nand \U$65273 ( \65660 , \65658 , \65659 );
_DC gfded ( \65661_nGfded , \65660 , \65580 );
buf \U$65274 ( \65662 , \65661_nGfded );
not \U$65275 ( \65663 , \65359 );
xor \U$65276 ( \65664 , \64413 , \64412 );
not \U$65277 ( \65665 , \65664 );
or \U$65278 ( \65666 , \65663 , \65665 );
or \U$65279 ( \65667 , \65664 , \65359 );
nand \U$65280 ( \65668 , \65666 , \65667 );
_DC gfd15 ( \65669_nGfd15 , \65668 , \65580 );
buf \U$65281 ( \65670 , \65669_nGfd15 );
not \U$65282 ( \65671 , \65357 );
xor \U$65283 ( \65672 , \64418 , \64419 );
not \U$65284 ( \65673 , \65672 );
or \U$65285 ( \65674 , \65671 , \65673 );
or \U$65286 ( \65675 , \65672 , \65357 );
nand \U$65287 ( \65676 , \65674 , \65675 );
_DC gfc38 ( \65677_nGfc38 , \65676 , \65580 );
buf \U$65288 ( \65678 , \65677_nGfc38 );
not \U$65289 ( \65679 , \65355 );
xor \U$65290 ( \65680 , \64424 , \64425 );
not \U$65291 ( \65681 , \65680 );
or \U$65292 ( \65682 , \65679 , \65681 );
or \U$65293 ( \65683 , \65680 , \65355 );
nand \U$65294 ( \65684 , \65682 , \65683 );
_DC gfb46 ( \65685_nGfb46 , \65684 , \65580 );
buf \U$65295 ( \65686 , \65685_nGfb46 );
not \U$65296 ( \65687 , \65353 );
xor \U$65297 ( \65688 , \64430 , \64431 );
not \U$65298 ( \65689 , \65688 );
or \U$65299 ( \65690 , \65687 , \65689 );
or \U$65300 ( \65691 , \65688 , \65353 );
nand \U$65301 ( \65692 , \65690 , \65691 );
_DC gfa24 ( \65693_nGfa24 , \65692 , \65580 );
buf \U$65302 ( \65694 , \65693_nGfa24 );
not \U$65303 ( \65695 , \65351 );
xor \U$65304 ( \65696 , \64437 , \64436 );
not \U$65305 ( \65697 , \65696 );
or \U$65306 ( \65698 , \65695 , \65697 );
or \U$65307 ( \65699 , \65696 , \65351 );
nand \U$65308 ( \65700 , \65698 , \65699 );
_DC gf914 ( \65701_nGf914 , \65700 , \65580 );
buf \U$65309 ( \65702 , \65701_nGf914 );
not \U$65310 ( \65703 , \65349 );
xor \U$65311 ( \65704 , \64443 , \64442 );
not \U$65312 ( \65705 , \65704 );
or \U$65313 ( \65706 , \65703 , \65705 );
or \U$65314 ( \65707 , \65704 , \65349 );
nand \U$65315 ( \65708 , \65706 , \65707 );
_DC gf7e6 ( \65709_nGf7e6 , \65708 , \65580 );
buf \U$65316 ( \65710 , \65709_nGf7e6 );
not \U$65317 ( \65711 , \65347 );
xor \U$65318 ( \65712 , \64449 , \64448 );
not \U$65319 ( \65713 , \65712 );
or \U$65320 ( \65714 , \65711 , \65713 );
or \U$65321 ( \65715 , \65712 , \65347 );
nand \U$65322 ( \65716 , \65714 , \65715 );
_DC gf6c6 ( \65717_nGf6c6 , \65716 , \65580 );
buf \U$65323 ( \65718 , \65717_nGf6c6 );
not \U$65324 ( \65719 , \65345 );
xor \U$65325 ( \65720 , \64454 , \64455 );
not \U$65326 ( \65721 , \65720 );
or \U$65327 ( \65722 , \65719 , \65721 );
or \U$65328 ( \65723 , \65720 , \65345 );
nand \U$65329 ( \65724 , \65722 , \65723 );
_DC gf581 ( \65725_nGf581 , \65724 , \65580 );
buf \U$65330 ( \65726 , \65725_nGf581 );
not \U$65331 ( \65727 , \65343 );
xor \U$65332 ( \65728 , \64460 , \64461 );
not \U$65333 ( \65729 , \65728 );
or \U$65334 ( \65730 , \65727 , \65729 );
or \U$65335 ( \65731 , \65728 , \65343 );
nand \U$65336 ( \65732 , \65730 , \65731 );
_DC gf429 ( \65733_nGf429 , \65732 , \65580 );
buf \U$65337 ( \65734 , \65733_nGf429 );
not \U$65338 ( \65735 , \65341 );
xor \U$65339 ( \65736 , \64467 , \64466 );
not \U$65340 ( \65737 , \65736 );
or \U$65341 ( \65738 , \65735 , \65737 );
or \U$65342 ( \65739 , \65736 , \65341 );
nand \U$65343 ( \65740 , \65738 , \65739 );
_DC gf2c7 ( \65741_nGf2c7 , \65740 , \65580 );
buf \U$65344 ( \65742 , \65741_nGf2c7 );
not \U$65345 ( \65743 , \65339 );
xor \U$65346 ( \65744 , \64473 , \64472 );
not \U$65347 ( \65745 , \65744 );
or \U$65348 ( \65746 , \65743 , \65745 );
or \U$65349 ( \65747 , \65744 , \65339 );
nand \U$65350 ( \65748 , \65746 , \65747 );
_DC gf156 ( \65749_nGf156 , \65748 , \65580 );
buf \U$65351 ( \65750 , \65749_nGf156 );
not \U$65352 ( \65751 , \65337 );
xor \U$65353 ( \65752 , \64479 , \64478 );
not \U$65354 ( \65753 , \65752 );
or \U$65355 ( \65754 , \65751 , \65753 );
or \U$65356 ( \65755 , \65752 , \65337 );
nand \U$65357 ( \65756 , \65754 , \65755 );
_DC gefd8 ( \65757_nGefd8 , \65756 , \65580 );
buf \U$65358 ( \65758 , \65757_nGefd8 );
not \U$65359 ( \65759 , \65335 );
xor \U$65360 ( \65760 , \64484 , \64485 );
not \U$65361 ( \65761 , \65760 );
or \U$65362 ( \65762 , \65759 , \65761 );
or \U$65363 ( \65763 , \65760 , \65335 );
nand \U$65364 ( \65764 , \65762 , \65763 );
_DC gee3c ( \65765_nGee3c , \65764 , \65580 );
buf \U$65365 ( \65766 , \65765_nGee3c );
not \U$65366 ( \65767 , \65333 );
xor \U$65367 ( \65768 , \64491 , \64490 );
not \U$65368 ( \65769 , \65768 );
or \U$65369 ( \65770 , \65767 , \65769 );
or \U$65370 ( \65771 , \65768 , \65333 );
nand \U$65371 ( \65772 , \65770 , \65771 );
_DC gec7d ( \65773_nGec7d , \65772 , \65580 );
buf \U$65372 ( \65774 , \65773_nGec7d );
not \U$65373 ( \65775 , \65331 );
xor \U$65374 ( \65776 , \64496 , \64497 );
not \U$65375 ( \65777 , \65776 );
or \U$65376 ( \65778 , \65775 , \65777 );
or \U$65377 ( \65779 , \65776 , \65331 );
nand \U$65378 ( \65780 , \65778 , \65779 );
_DC gea87 ( \65781_nGea87 , \65780 , \65580 );
buf \U$65379 ( \65782 , \65781_nGea87 );
not \U$65380 ( \65783 , \65329 );
xor \U$65381 ( \65784 , \64506 , \64507 );
not \U$65382 ( \65785 , \65784 );
or \U$65383 ( \65786 , \65783 , \65785 );
or \U$65384 ( \65787 , \65784 , \65329 );
nand \U$65385 ( \65788 , \65786 , \65787 );
_DC ge8b1 ( \65789_nGe8b1 , \65788 , \65580 );
buf \U$65386 ( \65790 , \65789_nGe8b1 );
not \U$65387 ( \65791 , \65327 );
xor \U$65388 ( \65792 , \64513 , \64512 );
not \U$65389 ( \65793 , \65792 );
or \U$65390 ( \65794 , \65791 , \65793 );
or \U$65391 ( \65795 , \65792 , \65327 );
nand \U$65392 ( \65796 , \65794 , \65795 );
_DC ge6d4 ( \65797_nGe6d4 , \65796 , \65580 );
buf \U$65393 ( \65798 , \65797_nGe6d4 );
not \U$65394 ( \65799 , \65325 );
xor \U$65395 ( \65800 , \64519 , \64518 );
not \U$65396 ( \65801 , \65800 );
or \U$65397 ( \65802 , \65799 , \65801 );
or \U$65398 ( \65803 , \65800 , \65325 );
nand \U$65399 ( \65804 , \65802 , \65803 );
_DC ge4e7 ( \65805_nGe4e7 , \65804 , \65580 );
buf \U$65400 ( \65806 , \65805_nGe4e7 );
not \U$65401 ( \65807 , \65323 );
xor \U$65402 ( \65808 , \64525 , \64524 );
not \U$65403 ( \65809 , \65808 );
or \U$65404 ( \65810 , \65807 , \65809 );
or \U$65405 ( \65811 , \65808 , \65323 );
nand \U$65406 ( \65812 , \65810 , \65811 );
_DC ge2e5 ( \65813_nGe2e5 , \65812 , \65580 );
buf \U$65407 ( \65814 , \65813_nGe2e5 );
not \U$65408 ( \65815 , \65321 );
xor \U$65409 ( \65816 , \64530 , \64531 );
not \U$65410 ( \65817 , \65816 );
or \U$65411 ( \65818 , \65815 , \65817 );
or \U$65412 ( \65819 , \65816 , \65321 );
nand \U$65413 ( \65820 , \65818 , \65819 );
_DC ge0da ( \65821_nGe0da , \65820 , \65580 );
buf \U$65414 ( \65822 , \65821_nGe0da );
not \U$65415 ( \65823 , \65319 );
xor \U$65416 ( \65824 , \64537 , \64536 );
not \U$65417 ( \65825 , \65824 );
or \U$65418 ( \65826 , \65823 , \65825 );
or \U$65419 ( \65827 , \65824 , \65319 );
nand \U$65420 ( \65828 , \65826 , \65827 );
_DC gdec8 ( \65829_nGdec8 , \65828 , \65580 );
buf \U$65421 ( \65830 , \65829_nGdec8 );
not \U$65422 ( \65831 , \65317 );
xor \U$65423 ( \65832 , \64542 , \64543 );
not \U$65424 ( \65833 , \65832 );
or \U$65425 ( \65834 , \65831 , \65833 );
or \U$65426 ( \65835 , \65832 , \65317 );
nand \U$65427 ( \65836 , \65834 , \65835 );
_DC gdcc3 ( \65837_nGdcc3 , \65836 , \65580 );
buf \U$65428 ( \65838 , \65837_nGdcc3 );
not \U$65429 ( \65839 , \65315 );
xor \U$65430 ( \65840 , \64556 , \64551 );
not \U$65431 ( \65841 , \65840 );
or \U$65432 ( \65842 , \65839 , \65841 );
or \U$65433 ( \65843 , \65840 , \65315 );
nand \U$65434 ( \65844 , \65842 , \65843 );
_DC gda9d ( \65845_nGda9d , \65844 , \65580 );
buf \U$65435 ( \65846 , \65845_nGda9d );
not \U$65436 ( \65847 , \65313 );
xor \U$65437 ( \65848 , \64569 , \64564 );
not \U$65438 ( \65849 , \65848 );
or \U$65439 ( \65850 , \65847 , \65849 );
or \U$65440 ( \65851 , \65848 , \65313 );
nand \U$65441 ( \65852 , \65850 , \65851 );
_DC gd85e ( \65853_nGd85e , \65852 , \65580 );
buf \U$65442 ( \65854 , \65853_nGd85e );
not \U$65443 ( \65855 , \65311 );
xor \U$65444 ( \65856 , \64578 , \64577 );
not \U$65445 ( \65857 , \65856 );
or \U$65446 ( \65858 , \65855 , \65857 );
or \U$65447 ( \65859 , \65856 , \65311 );
nand \U$65448 ( \65860 , \65858 , \65859 );
_DC gd657 ( \65861_nGd657 , \65860 , \65580 );
buf \U$65449 ( \65862 , \65861_nGd657 );
not \U$65450 ( \65863 , \65309 );
xor \U$65451 ( \65864 , \64583 , \64584 );
not \U$65452 ( \65865 , \65864 );
or \U$65453 ( \65866 , \65863 , \65865 );
or \U$65454 ( \65867 , \65864 , \65309 );
nand \U$65455 ( \65868 , \65866 , \65867 );
_DC gd41d ( \65869_nGd41d , \65868 , \65580 );
buf \U$65456 ( \65870 , \65869_nGd41d );
not \U$65457 ( \65871 , \65307 );
xor \U$65458 ( \65872 , \64590 , \64589 );
not \U$65459 ( \65873 , \65872 );
or \U$65460 ( \65874 , \65871 , \65873 );
or \U$65461 ( \65875 , \65872 , \65307 );
nand \U$65462 ( \65876 , \65874 , \65875 );
_DC gd1fd ( \65877_nGd1fd , \65876 , \65580 );
buf \U$65463 ( \65878 , \65877_nGd1fd );
not \U$65464 ( \65879 , \65305 );
xor \U$65465 ( \65880 , \64595 , \64596 );
not \U$65466 ( \65881 , \65880 );
or \U$65467 ( \65882 , \65879 , \65881 );
or \U$65468 ( \65883 , \65880 , \65305 );
nand \U$65469 ( \65884 , \65882 , \65883 );
_DC gcfa1 ( \65885_nGcfa1 , \65884 , \65580 );
buf \U$65470 ( \65886 , \65885_nGcfa1 );
not \U$65471 ( \65887 , \65303 );
xor \U$65472 ( \65888 , \64602 , \64601 );
not \U$65473 ( \65889 , \65888 );
or \U$65474 ( \65890 , \65887 , \65889 );
or \U$65475 ( \65891 , \65888 , \65303 );
nand \U$65476 ( \65892 , \65890 , \65891 );
_DC gcd2c ( \65893_nGcd2c , \65892 , \65580 );
buf \U$65477 ( \65894 , \65893_nGcd2c );
not \U$65478 ( \65895 , \65301 );
xor \U$65479 ( \65896 , \64611 , \64612 );
not \U$65480 ( \65897 , \65896 );
or \U$65481 ( \65898 , \65895 , \65897 );
or \U$65482 ( \65899 , \65896 , \65301 );
nand \U$65483 ( \65900 , \65898 , \65899 );
_DC gca99 ( \65901_nGca99 , \65900 , \65580 );
buf \U$65484 ( \65902 , \65901_nGca99 );
not \U$65485 ( \65903 , \65299 );
xor \U$65486 ( \65904 , \64617 , \64618 );
not \U$65487 ( \65905 , \65904 );
or \U$65488 ( \65906 , \65903 , \65905 );
or \U$65489 ( \65907 , \65904 , \65299 );
nand \U$65490 ( \65908 , \65906 , \65907 );
_DC gc812 ( \65909_nGc812 , \65908 , \65580 );
buf \U$65491 ( \65910 , \65909_nGc812 );
not \U$65492 ( \65911 , \65297 );
xor \U$65493 ( \65912 , \64624 , \64623 );
not \U$65494 ( \65913 , \65912 );
or \U$65495 ( \65914 , \65911 , \65913 );
or \U$65496 ( \65915 , \65912 , \65297 );
nand \U$65497 ( \65916 , \65914 , \65915 );
_DC gc589 ( \65917_nGc589 , \65916 , \65580 );
buf \U$65498 ( \65918 , \65917_nGc589 );
not \U$65499 ( \65919 , \65295 );
xor \U$65500 ( \65920 , \64634 , \64633 );
not \U$65501 ( \65921 , \65920 );
or \U$65502 ( \65922 , \65919 , \65921 );
or \U$65503 ( \65923 , \65920 , \65295 );
nand \U$65504 ( \65924 , \65922 , \65923 );
_DC gc2e5 ( \65925_nGc2e5 , \65924 , \65580 );
buf \U$65505 ( \65926 , \65925_nGc2e5 );
not \U$65506 ( \65927 , \65293 );
xor \U$65507 ( \65928 , \64640 , \64639 );
not \U$65508 ( \65929 , \65928 );
or \U$65509 ( \65930 , \65927 , \65929 );
or \U$65510 ( \65931 , \65928 , \65293 );
nand \U$65511 ( \65932 , \65930 , \65931 );
_DC gbff1 ( \65933_nGbff1 , \65932 , \65580 );
buf \U$65512 ( \65934 , \65933_nGbff1 );
not \U$65513 ( \65935 , \65291 );
xor \U$65514 ( \65936 , \64645 , \64646 );
not \U$65515 ( \65937 , \65936 );
or \U$65516 ( \65938 , \65935 , \65937 );
or \U$65517 ( \65939 , \65936 , \65291 );
nand \U$65518 ( \65940 , \65938 , \65939 );
_DC gbcf3 ( \65941_nGbcf3 , \65940 , \65580 );
buf \U$65519 ( \65942 , \65941_nGbcf3 );
not \U$65520 ( \65943 , \65289 );
xor \U$65521 ( \65944 , \64652 , \64651 );
not \U$65522 ( \65945 , \65944 );
or \U$65523 ( \65946 , \65943 , \65945 );
or \U$65524 ( \65947 , \65944 , \65289 );
nand \U$65525 ( \65948 , \65946 , \65947 );
_DC gba17 ( \65949_nGba17 , \65948 , \65580 );
buf \U$65526 ( \65950 , \65949_nGba17 );
not \U$65527 ( \65951 , \65287 );
xor \U$65528 ( \65952 , \64657 , \64658 );
not \U$65529 ( \65953 , \65952 );
or \U$65530 ( \65954 , \65951 , \65953 );
or \U$65531 ( \65955 , \65952 , \65287 );
nand \U$65532 ( \65956 , \65954 , \65955 );
_DC gb727 ( \65957_nGb727 , \65956 , \65580 );
buf \U$65533 ( \65958 , \65957_nGb727 );
not \U$65534 ( \65959 , \65285 );
xor \U$65535 ( \65960 , \64663 , \64664 );
not \U$65536 ( \65961 , \65960 );
or \U$65537 ( \65962 , \65959 , \65961 );
or \U$65538 ( \65963 , \65960 , \65285 );
nand \U$65539 ( \65964 , \65962 , \65963 );
_DC gb43a ( \65965_nGb43a , \65964 , \65580 );
buf \U$65540 ( \65966 , \65965_nGb43a );
not \U$65541 ( \65967 , \65283 );
xor \U$65542 ( \65968 , \64669 , \64670 );
not \U$65543 ( \65969 , \65968 );
or \U$65544 ( \65970 , \65967 , \65969 );
or \U$65545 ( \65971 , \65968 , \65283 );
nand \U$65546 ( \65972 , \65970 , \65971 );
_DC gb150 ( \65973_nGb150 , \65972 , \65580 );
buf \U$65547 ( \65974 , \65973_nGb150 );
not \U$65548 ( \65975 , \65281 );
xor \U$65549 ( \65976 , \64679 , \64678 );
not \U$65550 ( \65977 , \65976 );
or \U$65551 ( \65978 , \65975 , \65977 );
or \U$65552 ( \65979 , \65976 , \65281 );
nand \U$65553 ( \65980 , \65978 , \65979 );
_DC gae24 ( \65981_nGae24 , \65980 , \65580 );
buf \U$65554 ( \65982 , \65981_nGae24 );
not \U$65555 ( \65983 , \65279 );
xor \U$65556 ( \65984 , \64684 , \64685 );
not \U$65557 ( \65985 , \65984 );
or \U$65558 ( \65986 , \65983 , \65985 );
or \U$65559 ( \65987 , \65984 , \65279 );
nand \U$65560 ( \65988 , \65986 , \65987 );
_DC gaae2 ( \65989_nGaae2 , \65988 , \65580 );
buf \U$65561 ( \65990 , \65989_nGaae2 );
not \U$65562 ( \65991 , \65277 );
xor \U$65563 ( \65992 , \64691 , \64690 );
not \U$65564 ( \65993 , \65992 );
or \U$65565 ( \65994 , \65991 , \65993 );
or \U$65566 ( \65995 , \65992 , \65277 );
nand \U$65567 ( \65996 , \65994 , \65995 );
_DC ga7c6 ( \65997_nGa7c6 , \65996 , \65580 );
buf \U$65568 ( \65998 , \65997_nGa7c6 );
not \U$65569 ( \65999 , \65275 );
xor \U$65570 ( \66000 , \64697 , \64696 );
not \U$65571 ( \66001 , \66000 );
or \U$65572 ( \66002 , \65999 , \66001 );
or \U$65573 ( \66003 , \66000 , \65275 );
nand \U$65574 ( \66004 , \66002 , \66003 );
_DC ga4a9 ( \66005_nGa4a9 , \66004 , \65580 );
buf \U$65575 ( \66006 , \66005_nGa4a9 );
not \U$65576 ( \66007 , \65273 );
xor \U$65577 ( \66008 , \64703 , \64702 );
not \U$65578 ( \66009 , \66008 );
or \U$65579 ( \66010 , \66007 , \66009 );
or \U$65580 ( \66011 , \66008 , \65273 );
nand \U$65581 ( \66012 , \66010 , \66011 );
_DC ga14c ( \66013_nGa14c , \66012 , \65580 );
buf \U$65582 ( \66014 , \66013_nGa14c );
not \U$65583 ( \66015 , \65271 );
xor \U$65584 ( \66016 , \64708 , \64709 );
not \U$65585 ( \66017 , \66016 );
or \U$65586 ( \66018 , \66015 , \66017 );
or \U$65587 ( \66019 , \66016 , \65271 );
nand \U$65588 ( \66020 , \66018 , \66019 );
_DC g9ddd ( \66021_nG9ddd , \66020 , \65580 );
buf \U$65589 ( \66022 , \66021_nG9ddd );
not \U$65590 ( \66023 , \65269 );
xor \U$65591 ( \66024 , \64715 , \64714 );
not \U$65592 ( \66025 , \66024 );
or \U$65593 ( \66026 , \66023 , \66025 );
or \U$65594 ( \66027 , \66024 , \65269 );
nand \U$65595 ( \66028 , \66026 , \66027 );
_DC g9a6c ( \66029_nG9a6c , \66028 , \65580 );
buf \U$65596 ( \66030 , \66029_nG9a6c );
not \U$65597 ( \66031 , \65267 );
xor \U$65598 ( \66032 , \64721 , \64720 );
not \U$65599 ( \66033 , \66032 );
or \U$65600 ( \66034 , \66031 , \66033 );
or \U$65601 ( \66035 , \66032 , \65267 );
nand \U$65602 ( \66036 , \66034 , \66035 );
_DC g9704 ( \66037_nG9704 , \66036 , \65580 );
buf \U$65603 ( \66038 , \66037_nG9704 );
not \U$65604 ( \66039 , \65265 );
xor \U$65605 ( \66040 , \64727 , \64726 );
not \U$65606 ( \66041 , \66040 );
or \U$65607 ( \66042 , \66039 , \66041 );
or \U$65608 ( \66043 , \66040 , \65265 );
nand \U$65609 ( \66044 , \66042 , \66043 );
_DC g9381 ( \66045_nG9381 , \66044 , \65580 );
buf \U$65610 ( \66046 , \66045_nG9381 );
not \U$65611 ( \66047 , \65263 );
xor \U$65612 ( \66048 , \64733 , \64732 );
not \U$65613 ( \66049 , \66048 );
or \U$65614 ( \66050 , \66047 , \66049 );
or \U$65615 ( \66051 , \66048 , \65263 );
nand \U$65616 ( \66052 , \66050 , \66051 );
_DC g8ff4 ( \66053_nG8ff4 , \66052 , \65580 );
buf \U$65617 ( \66054 , \66053_nG8ff4 );
not \U$65618 ( \66055 , \65261 );
xor \U$65619 ( \66056 , \64739 , \64738 );
not \U$65620 ( \66057 , \66056 );
or \U$65621 ( \66058 , \66055 , \66057 );
or \U$65622 ( \66059 , \66056 , \65261 );
nand \U$65623 ( \66060 , \66058 , \66059 );
_DC g8c7b ( \66061_nG8c7b , \66060 , \65580 );
buf \U$65624 ( \66062 , \66061_nG8c7b );
not \U$65625 ( \66063 , \65259 );
xor \U$65626 ( \66064 , \64745 , \64744 );
not \U$65627 ( \66065 , \66064 );
or \U$65628 ( \66066 , \66063 , \66065 );
or \U$65629 ( \66067 , \66064 , \65259 );
nand \U$65630 ( \66068 , \66066 , \66067 );
_DC g88e4 ( \66069_nG88e4 , \66068 , \65580 );
buf \U$65631 ( \66070 , \66069_nG88e4 );
not \U$65632 ( \66071 , \65257 );
xor \U$65633 ( \66072 , \64751 , \64750 );
not \U$65634 ( \66073 , \66072 );
or \U$65635 ( \66074 , \66071 , \66073 );
or \U$65636 ( \66075 , \66072 , \65257 );
nand \U$65637 ( \66076 , \66074 , \66075 );
_DC g850c ( \66077_nG850c , \66076 , \65580 );
buf \U$65638 ( \66078 , \66077_nG850c );
not \U$65639 ( \66079 , \65255 );
xor \U$65640 ( \66080 , \64757 , \64756 );
not \U$65641 ( \66081 , \66080 );
or \U$65642 ( \66082 , \66079 , \66081 );
or \U$65643 ( \66083 , \66080 , \65255 );
nand \U$65644 ( \66084 , \66082 , \66083 );
_DC g80dd ( \66085_nG80dd , \66084 , \65580 );
buf \U$65645 ( \66086 , \66085_nG80dd );
not \U$65646 ( \66087 , \65253 );
xor \U$65647 ( \66088 , \64763 , \64762 );
not \U$65648 ( \66089 , \66088 );
or \U$65649 ( \66090 , \66087 , \66089 );
or \U$65650 ( \66091 , \66088 , \65253 );
nand \U$65651 ( \66092 , \66090 , \66091 );
_DC g7cf2 ( \66093_nG7cf2 , \66092 , \65580 );
buf \U$65652 ( \66094 , \66093_nG7cf2 );
not \U$65653 ( \66095 , \65251 );
xor \U$65654 ( \66096 , \64769 , \64768 );
not \U$65655 ( \66097 , \66096 );
or \U$65656 ( \66098 , \66095 , \66097 );
or \U$65657 ( \66099 , \66096 , \65251 );
nand \U$65658 ( \66100 , \66098 , \66099 );
_DC g7913 ( \66101_nG7913 , \66100 , \65580 );
buf \U$65659 ( \66102 , \66101_nG7913 );
not \U$65660 ( \66103 , \65249 );
xor \U$65661 ( \66104 , \64775 , \64774 );
not \U$65662 ( \66105 , \66104 );
or \U$65663 ( \66106 , \66103 , \66105 );
or \U$65664 ( \66107 , \66104 , \65249 );
nand \U$65665 ( \66108 , \66106 , \66107 );
_DC g7586 ( \66109_nG7586 , \66108 , \65580 );
buf \U$65666 ( \66110 , \66109_nG7586 );
not \U$65667 ( \66111 , \65247 );
xor \U$65668 ( \66112 , \64781 , \64780 );
not \U$65669 ( \66113 , \66112 );
or \U$65670 ( \66114 , \66111 , \66113 );
or \U$65671 ( \66115 , \66112 , \65247 );
nand \U$65672 ( \66116 , \66114 , \66115 );
_DC g7216 ( \66117_nG7216 , \66116 , \65580 );
buf \U$65673 ( \66118 , \66117_nG7216 );
not \U$65674 ( \66119 , \65245 );
xor \U$65675 ( \66120 , \64787 , \64786 );
not \U$65676 ( \66121 , \66120 );
or \U$65677 ( \66122 , \66119 , \66121 );
or \U$65678 ( \66123 , \66120 , \65245 );
nand \U$65679 ( \66124 , \66122 , \66123 );
_DC g6ea7 ( \66125_nG6ea7 , \66124 , \65580 );
buf \U$65680 ( \66126 , \66125_nG6ea7 );
not \U$65681 ( \66127 , \65243 );
xor \U$65682 ( \66128 , \64793 , \64792 );
not \U$65683 ( \66129 , \66128 );
or \U$65684 ( \66130 , \66127 , \66129 );
or \U$65685 ( \66131 , \66128 , \65243 );
nand \U$65686 ( \66132 , \66130 , \66131 );
_DC g6b15 ( \66133_nG6b15 , \66132 , \65580 );
buf \U$65687 ( \66134 , \66133_nG6b15 );
not \U$65688 ( \66135 , \65241 );
xor \U$65689 ( \66136 , \64799 , \64798 );
not \U$65690 ( \66137 , \66136 );
or \U$65691 ( \66138 , \66135 , \66137 );
or \U$65692 ( \66139 , \66136 , \65241 );
nand \U$65693 ( \66140 , \66138 , \66139 );
_DC g6785 ( \66141_nG6785 , \66140 , \65580 );
buf \U$65694 ( \66142 , \66141_nG6785 );
not \U$65695 ( \66143 , \65239 );
xor \U$65696 ( \66144 , \64805 , \64804 );
not \U$65697 ( \66145 , \66144 );
or \U$65698 ( \66146 , \66143 , \66145 );
or \U$65699 ( \66147 , \66144 , \65239 );
nand \U$65700 ( \66148 , \66146 , \66147 );
_DC g642a ( \66149_nG642a , \66148 , \65580 );
buf \U$65701 ( \66150 , \66149_nG642a );
not \U$65702 ( \66151 , \65237 );
xor \U$65703 ( \66152 , \64811 , \64810 );
not \U$65704 ( \66153 , \66152 );
or \U$65705 ( \66154 , \66151 , \66153 );
or \U$65706 ( \66155 , \66152 , \65237 );
nand \U$65707 ( \66156 , \66154 , \66155 );
_DC g60ac ( \66157_nG60ac , \66156 , \65580 );
buf \U$65708 ( \66158 , \66157_nG60ac );
not \U$65709 ( \66159 , \65235 );
xor \U$65710 ( \66160 , \64817 , \64816 );
not \U$65711 ( \66161 , \66160 );
or \U$65712 ( \66162 , \66159 , \66161 );
or \U$65713 ( \66163 , \66160 , \65235 );
nand \U$65714 ( \66164 , \66162 , \66163 );
_DC g5d39 ( \66165_nG5d39 , \66164 , \65580 );
buf \U$65715 ( \66166 , \66165_nG5d39 );
not \U$65716 ( \66167 , \65233 );
xor \U$65717 ( \66168 , \64823 , \64822 );
not \U$65718 ( \66169 , \66168 );
or \U$65719 ( \66170 , \66167 , \66169 );
or \U$65720 ( \66171 , \66168 , \65233 );
nand \U$65721 ( \66172 , \66170 , \66171 );
_DC g5a0d ( \66173_nG5a0d , \66172 , \65580 );
buf \U$65722 ( \66174 , \66173_nG5a0d );
not \U$65723 ( \66175 , \65231 );
xor \U$65724 ( \66176 , \64829 , \64828 );
not \U$65725 ( \66177 , \66176 );
or \U$65726 ( \66178 , \66175 , \66177 );
or \U$65727 ( \66179 , \66176 , \65231 );
nand \U$65728 ( \66180 , \66178 , \66179 );
_DC g5705 ( \66181_nG5705 , \66180 , \65580 );
buf \U$65729 ( \66182 , \66181_nG5705 );
not \U$65730 ( \66183 , \65229 );
xor \U$65731 ( \66184 , \64835 , \64834 );
not \U$65732 ( \66185 , \66184 );
or \U$65733 ( \66186 , \66183 , \66185 );
or \U$65734 ( \66187 , \66184 , \65229 );
nand \U$65735 ( \66188 , \66186 , \66187 );
_DC g5400 ( \66189_nG5400 , \66188 , \65580 );
buf \U$65736 ( \66190 , \66189_nG5400 );
not \U$65737 ( \66191 , \65227 );
xor \U$65738 ( \66192 , \64841 , \64840 );
not \U$65739 ( \66193 , \66192 );
or \U$65740 ( \66194 , \66191 , \66193 );
or \U$65741 ( \66195 , \66192 , \65227 );
nand \U$65742 ( \66196 , \66194 , \66195 );
_DC g50b7 ( \66197_nG50b7 , \66196 , \65580 );
buf \U$65743 ( \66198 , \66197_nG50b7 );
not \U$65744 ( \66199 , \65225 );
xor \U$65745 ( \66200 , \64847 , \64846 );
not \U$65746 ( \66201 , \66200 );
or \U$65747 ( \66202 , \66199 , \66201 );
or \U$65748 ( \66203 , \66200 , \65225 );
nand \U$65749 ( \66204 , \66202 , \66203 );
_DC g4d9f ( \66205_nG4d9f , \66204 , \65580 );
buf \U$65750 ( \66206 , \66205_nG4d9f );
not \U$65751 ( \66207 , \65223 );
xor \U$65752 ( \66208 , \64853 , \64852 );
not \U$65753 ( \66209 , \66208 );
or \U$65754 ( \66210 , \66207 , \66209 );
or \U$65755 ( \66211 , \66208 , \65223 );
nand \U$65756 ( \66212 , \66210 , \66211 );
_DC g4aba ( \66213_nG4aba , \66212 , \65580 );
buf \U$65757 ( \66214 , \66213_nG4aba );
not \U$65758 ( \66215 , \65221 );
xor \U$65759 ( \66216 , \64859 , \64858 );
not \U$65760 ( \66217 , \66216 );
or \U$65761 ( \66218 , \66215 , \66217 );
or \U$65762 ( \66219 , \66216 , \65221 );
nand \U$65763 ( \66220 , \66218 , \66219 );
_DC g47cd ( \66221_nG47cd , \66220 , \65580 );
buf \U$65764 ( \66222 , \66221_nG47cd );
not \U$65765 ( \66223 , \65219 );
xor \U$65766 ( \66224 , \64865 , \64864 );
not \U$65767 ( \66225 , \66224 );
or \U$65768 ( \66226 , \66223 , \66225 );
or \U$65769 ( \66227 , \66224 , \65219 );
nand \U$65770 ( \66228 , \66226 , \66227 );
_DC g44fd ( \66229_nG44fd , \66228 , \65580 );
buf \U$65771 ( \66230 , \66229_nG44fd );
not \U$65772 ( \66231 , \65217 );
xor \U$65773 ( \66232 , \64871 , \64870 );
not \U$65774 ( \66233 , \66232 );
or \U$65775 ( \66234 , \66231 , \66233 );
or \U$65776 ( \66235 , \66232 , \65217 );
nand \U$65777 ( \66236 , \66234 , \66235 );
_DC g4250 ( \66237_nG4250 , \66236 , \65580 );
buf \U$65778 ( \66238 , \66237_nG4250 );
not \U$65779 ( \66239 , \65215 );
xor \U$65780 ( \66240 , \64877 , \64876 );
not \U$65781 ( \66241 , \66240 );
or \U$65782 ( \66242 , \66239 , \66241 );
or \U$65783 ( \66243 , \66240 , \65215 );
nand \U$65784 ( \66244 , \66242 , \66243 );
_DC g3f85 ( \66245_nG3f85 , \66244 , \65580 );
buf \U$65785 ( \66246 , \66245_nG3f85 );
not \U$65786 ( \66247 , \65213 );
xor \U$65787 ( \66248 , \64883 , \64882 );
not \U$65788 ( \66249 , \66248 );
or \U$65789 ( \66250 , \66247 , \66249 );
or \U$65790 ( \66251 , \66248 , \65213 );
nand \U$65791 ( \66252 , \66250 , \66251 );
_DC g3cff ( \66253_nG3cff , \66252 , \65580 );
buf \U$65792 ( \66254 , \66253_nG3cff );
not \U$65793 ( \66255 , \65211 );
xor \U$65794 ( \66256 , \64889 , \64888 );
not \U$65795 ( \66257 , \66256 );
or \U$65796 ( \66258 , \66255 , \66257 );
or \U$65797 ( \66259 , \66256 , \65211 );
nand \U$65798 ( \66260 , \66258 , \66259 );
_DC g3a58 ( \66261_nG3a58 , \66260 , \65580 );
buf \U$65799 ( \66262 , \66261_nG3a58 );
not \U$65800 ( \66263 , \65209 );
xor \U$65801 ( \66264 , \64895 , \64894 );
not \U$65802 ( \66265 , \66264 );
or \U$65803 ( \66266 , \66263 , \66265 );
or \U$65804 ( \66267 , \66264 , \65209 );
nand \U$65805 ( \66268 , \66266 , \66267 );
_DC g37d2 ( \66269_nG37d2 , \66268 , \65580 );
buf \U$65806 ( \66270 , \66269_nG37d2 );
not \U$65807 ( \66271 , \65207 );
xor \U$65808 ( \66272 , \64900 , \64901 );
not \U$65809 ( \66273 , \66272 );
or \U$65810 ( \66274 , \66271 , \66273 );
or \U$65811 ( \66275 , \66272 , \65207 );
nand \U$65812 ( \66276 , \66274 , \66275 );
_DC g3580 ( \66277_nG3580 , \66276 , \65580 );
buf \U$65813 ( \66278 , \66277_nG3580 );
not \U$65814 ( \66279 , \65205 );
xor \U$65815 ( \66280 , \64907 , \64906 );
not \U$65816 ( \66281 , \66280 );
or \U$65817 ( \66282 , \66279 , \66281 );
or \U$65818 ( \66283 , \66280 , \65205 );
nand \U$65819 ( \66284 , \66282 , \66283 );
_DC g3327 ( \66285_nG3327 , \66284 , \65580 );
buf \U$65820 ( \66286 , \66285_nG3327 );
not \U$65821 ( \66287 , \65203 );
xor \U$65822 ( \66288 , \64913 , \64912 );
not \U$65823 ( \66289 , \66288 );
or \U$65824 ( \66290 , \66287 , \66289 );
or \U$65825 ( \66291 , \66288 , \65203 );
nand \U$65826 ( \66292 , \66290 , \66291 );
_DC g30eb ( \66293_nG30eb , \66292 , \65580 );
buf \U$65827 ( \66294 , \66293_nG30eb );
not \U$65828 ( \66295 , \65201 );
xor \U$65829 ( \66296 , \64919 , \64918 );
not \U$65830 ( \66297 , \66296 );
or \U$65831 ( \66298 , \66295 , \66297 );
or \U$65832 ( \66299 , \66296 , \65201 );
nand \U$65833 ( \66300 , \66298 , \66299 );
_DC g2eb3 ( \66301_nG2eb3 , \66300 , \65580 );
buf \U$65834 ( \66302 , \66301_nG2eb3 );
not \U$65835 ( \66303 , \65199 );
xor \U$65836 ( \66304 , \64924 , \64925 );
not \U$65837 ( \66305 , \66304 );
or \U$65838 ( \66306 , \66303 , \66305 );
or \U$65839 ( \66307 , \66304 , \65199 );
nand \U$65840 ( \66308 , \66306 , \66307 );
_DC g2c54 ( \66309_nG2c54 , \66308 , \65580 );
buf \U$65841 ( \66310 , \66309_nG2c54 );
not \U$65842 ( \66311 , \65197 );
xor \U$65843 ( \66312 , \64931 , \64930 );
not \U$65844 ( \66313 , \66312 );
or \U$65845 ( \66314 , \66311 , \66313 );
or \U$65846 ( \66315 , \66312 , \65197 );
nand \U$65847 ( \66316 , \66314 , \66315 );
_DC g2a16 ( \66317_nG2a16 , \66316 , \65580 );
buf \U$65848 ( \66318 , \66317_nG2a16 );
not \U$65849 ( \66319 , \65195 );
xor \U$65850 ( \66320 , \64937 , \64936 );
not \U$65851 ( \66321 , \66320 );
or \U$65852 ( \66322 , \66319 , \66321 );
or \U$65853 ( \66323 , \66320 , \65195 );
nand \U$65854 ( \66324 , \66322 , \66323 );
_DC g27e2 ( \66325_nG27e2 , \66324 , \65580 );
buf \U$65855 ( \66326 , \66325_nG27e2 );
not \U$65856 ( \66327 , \65193 );
xor \U$65857 ( \66328 , \64943 , \64942 );
not \U$65858 ( \66329 , \66328 );
or \U$65859 ( \66330 , \66327 , \66329 );
or \U$65860 ( \66331 , \66328 , \65193 );
nand \U$65861 ( \66332 , \66330 , \66331 );
_DC g25af ( \66333_nG25af , \66332 , \65580 );
buf \U$65862 ( \66334 , \66333_nG25af );
not \U$65863 ( \66335 , \65191 );
xor \U$65864 ( \66336 , \64948 , \64949 );
not \U$65865 ( \66337 , \66336 );
or \U$65866 ( \66338 , \66335 , \66337 );
or \U$65867 ( \66339 , \66336 , \65191 );
nand \U$65868 ( \66340 , \66338 , \66339 );
_DC g23ac ( \66341_nG23ac , \66340 , \65580 );
buf \U$65869 ( \66342 , \66341_nG23ac );
not \U$65870 ( \66343 , \65189 );
xor \U$65871 ( \66344 , \64954 , \64955 );
not \U$65872 ( \66345 , \66344 );
or \U$65873 ( \66346 , \66343 , \66345 );
or \U$65874 ( \66347 , \66344 , \65189 );
nand \U$65875 ( \66348 , \66346 , \66347 );
_DC g21c1 ( \66349_nG21c1 , \66348 , \65580 );
buf \U$65876 ( \66350 , \66349_nG21c1 );
not \U$65877 ( \66351 , \65187 );
xor \U$65878 ( \66352 , \64960 , \64961 );
not \U$65879 ( \66353 , \66352 );
or \U$65880 ( \66354 , \66351 , \66353 );
or \U$65881 ( \66355 , \66352 , \65187 );
nand \U$65882 ( \66356 , \66354 , \66355 );
_DC g1ff9 ( \66357_nG1ff9 , \66356 , \65580 );
buf \U$65883 ( \66358 , \66357_nG1ff9 );
not \U$65884 ( \66359 , \65185 );
xor \U$65885 ( \66360 , \64967 , \64966 );
not \U$65886 ( \66361 , \66360 );
or \U$65887 ( \66362 , \66359 , \66361 );
or \U$65888 ( \66363 , \66360 , \65185 );
nand \U$65889 ( \66364 , \66362 , \66363 );
_DC g1e19 ( \66365_nG1e19 , \66364 , \65580 );
buf \U$65890 ( \66366 , \66365_nG1e19 );
not \U$65891 ( \66367 , \65183 );
xor \U$65892 ( \66368 , \64973 , \64972 );
not \U$65893 ( \66369 , \66368 );
or \U$65894 ( \66370 , \66367 , \66369 );
or \U$65895 ( \66371 , \66368 , \65183 );
nand \U$65896 ( \66372 , \66370 , \66371 );
_DC g1c46 ( \66373_nG1c46 , \66372 , \65580 );
buf \U$65897 ( \66374 , \66373_nG1c46 );
not \U$65898 ( \66375 , \65181 );
xor \U$65899 ( \66376 , \64979 , \64978 );
not \U$65900 ( \66377 , \66376 );
or \U$65901 ( \66378 , \66375 , \66377 );
or \U$65902 ( \66379 , \66376 , \65181 );
nand \U$65903 ( \66380 , \66378 , \66379 );
_DC g1aa2 ( \66381_nG1aa2 , \66380 , \65580 );
buf \U$65904 ( \66382 , \66381_nG1aa2 );
not \U$65905 ( \66383 , \65179 );
xor \U$65906 ( \66384 , \64985 , \64984 );
not \U$65907 ( \66385 , \66384 );
or \U$65908 ( \66386 , \66383 , \66385 );
or \U$65909 ( \66387 , \66384 , \65179 );
nand \U$65910 ( \66388 , \66386 , \66387 );
_DC g190e ( \66389_nG190e , \66388 , \65580 );
buf \U$65911 ( \66390 , \66389_nG190e );
not \U$65912 ( \66391 , \65177 );
xor \U$65913 ( \66392 , \64990 , \64991 );
not \U$65914 ( \66393 , \66392 );
or \U$65915 ( \66394 , \66391 , \66393 );
or \U$65916 ( \66395 , \66392 , \65177 );
nand \U$65917 ( \66396 , \66394 , \66395 );
_DC g176a ( \66397_nG176a , \66396 , \65580 );
buf \U$65918 ( \66398 , \66397_nG176a );
not \U$65919 ( \66399 , \65175 );
xor \U$65920 ( \66400 , \64996 , \64997 );
not \U$65921 ( \66401 , \66400 );
or \U$65922 ( \66402 , \66399 , \66401 );
or \U$65923 ( \66403 , \66400 , \65175 );
nand \U$65924 ( \66404 , \66402 , \66403 );
_DC g10367 ( \66405_nG10367 , \66404 , \65580 );
buf \U$65925 ( \66406 , \66405_nG10367 );
not \U$65926 ( \66407 , \65173 );
xor \U$65927 ( \66408 , \65002 , \65003 );
not \U$65928 ( \66409 , \66408 );
or \U$65929 ( \66410 , \66407 , \66409 );
or \U$65930 ( \66411 , \66408 , \65173 );
nand \U$65931 ( \66412 , \66410 , \66411 );
_DC g10360 ( \66413_nG10360 , \66412 , \65580 );
buf \U$65932 ( \66414 , \66413_nG10360 );
not \U$65933 ( \66415 , \65171 );
xor \U$65934 ( \66416 , \65008 , \65009 );
not \U$65935 ( \66417 , \66416 );
or \U$65936 ( \66418 , \66415 , \66417 );
or \U$65937 ( \66419 , \66416 , \65171 );
nand \U$65938 ( \66420 , \66418 , \66419 );
_DC g10359 ( \66421_nG10359 , \66420 , \65580 );
buf \U$65939 ( \66422 , \66421_nG10359 );
not \U$65940 ( \66423 , \65169 );
xor \U$65941 ( \66424 , \65015 , \65014 );
not \U$65942 ( \66425 , \66424 );
or \U$65943 ( \66426 , \66423 , \66425 );
or \U$65944 ( \66427 , \66424 , \65169 );
nand \U$65945 ( \66428 , \66426 , \66427 );
_DC g10352 ( \66429_nG10352 , \66428 , \65580 );
buf \U$65946 ( \66430 , \66429_nG10352 );
not \U$65947 ( \66431 , \65167 );
xor \U$65948 ( \66432 , \65021 , \65020 );
not \U$65949 ( \66433 , \66432 );
or \U$65950 ( \66434 , \66431 , \66433 );
or \U$65951 ( \66435 , \66432 , \65167 );
nand \U$65952 ( \66436 , \66434 , \66435 );
_DC g1034b ( \66437_nG1034b , \66436 , \65580 );
buf \U$65953 ( \66438 , \66437_nG1034b );
not \U$65954 ( \66439 , \65165 );
xor \U$65955 ( \66440 , \65026 , \65027 );
not \U$65956 ( \66441 , \66440 );
or \U$65957 ( \66442 , \66439 , \66441 );
or \U$65958 ( \66443 , \66440 , \65165 );
nand \U$65959 ( \66444 , \66442 , \66443 );
_DC g10208 ( \66445_nG10208 , \66444 , \65580 );
buf \U$65960 ( \66446 , \66445_nG10208 );
not \U$65961 ( \66447 , \65163 );
xor \U$65962 ( \66448 , \65032 , \65033 );
not \U$65963 ( \66449 , \66448 );
or \U$65964 ( \66450 , \66447 , \66449 );
or \U$65965 ( \66451 , \66448 , \65163 );
nand \U$65966 ( \66452 , \66450 , \66451 );
_DC gec84 ( \66453_nGec84 , \66452 , \65580 );
buf \U$65967 ( \66454 , \66453_nGec84 );
not \U$65968 ( \66455 , \65161 );
xor \U$65969 ( \66456 , \65038 , \65039 );
not \U$65970 ( \66457 , \66456 );
or \U$65971 ( \66458 , \66455 , \66457 );
or \U$65972 ( \66459 , \66456 , \65161 );
nand \U$65973 ( \66460 , \66458 , \66459 );
_DC gd865 ( \66461_nGd865 , \66460 , \65580 );
buf \U$65974 ( \66462 , \66461_nGd865 );
not \U$65975 ( \66463 , \65159 );
xor \U$65976 ( \66464 , \65045 , \65044 );
not \U$65977 ( \66465 , \66464 );
or \U$65978 ( \66466 , \66463 , \66465 );
or \U$65979 ( \66467 , \66464 , \65159 );
nand \U$65980 ( \66468 , \66466 , \66467 );
_DC gc819 ( \66469_nGc819 , \66468 , \65580 );
buf \U$65981 ( \66470 , \66469_nGc819 );
not \U$65982 ( \66471 , \65157 );
xor \U$65983 ( \66472 , \65051 , \65050 );
not \U$65984 ( \66473 , \66472 );
or \U$65985 ( \66474 , \66471 , \66473 );
or \U$65986 ( \66475 , \66472 , \65157 );
nand \U$65987 ( \66476 , \66474 , \66475 );
_DC gb441 ( \66477_nGb441 , \66476 , \65580 );
buf \U$65988 ( \66478 , \66477_nGb441 );
not \U$65989 ( \66479 , \65155 );
xor \U$65990 ( \66480 , \65056 , \65057 );
not \U$65991 ( \66481 , \66480 );
or \U$65992 ( \66482 , \66479 , \66481 );
or \U$65993 ( \66483 , \66480 , \65155 );
nand \U$65994 ( \66484 , \66482 , \66483 );
_DC ga4b0 ( \66485_nGa4b0 , \66484 , \65580 );
buf \U$65995 ( \66486 , \66485_nGa4b0 );
not \U$65996 ( \66487 , \65153 );
xor \U$65997 ( \66488 , \65063 , \65062 );
not \U$65998 ( \66489 , \66488 );
or \U$65999 ( \66490 , \66487 , \66489 );
or \U$66000 ( \66491 , \66488 , \65153 );
nand \U$66001 ( \66492 , \66490 , \66491 );
_DC g970b ( \66493_nG970b , \66492 , \65580 );
buf \U$66002 ( \66494 , \66493_nG970b );
not \U$66003 ( \66495 , \65151 );
xor \U$66004 ( \66496 , \65068 , \65069 );
not \U$66005 ( \66497 , \66496 );
or \U$66006 ( \66498 , \66495 , \66497 );
or \U$66007 ( \66499 , \66496 , \65151 );
nand \U$66008 ( \66500 , \66498 , \66499 );
_DC g88eb ( \66501_nG88eb , \66500 , \65580 );
buf \U$66009 ( \66502 , \66501_nG88eb );
not \U$66010 ( \66503 , \65149 );
xor \U$66011 ( \66504 , \65075 , \65074 );
not \U$66012 ( \66505 , \66504 );
or \U$66013 ( \66506 , \66503 , \66505 );
or \U$66014 ( \66507 , \66504 , \65149 );
nand \U$66015 ( \66508 , \66506 , \66507 );
_DC g791a ( \66509_nG791a , \66508 , \65580 );
buf \U$66016 ( \66510 , \66509_nG791a );
not \U$66017 ( \66511 , \65147 );
xor \U$66018 ( \66512 , \65080 , \65081 );
not \U$66019 ( \66513 , \66512 );
or \U$66020 ( \66514 , \66511 , \66513 );
or \U$66021 ( \66515 , \66512 , \65147 );
nand \U$66022 ( \66516 , \66514 , \66515 );
_DC g6eae ( \66517_nG6eae , \66516 , \65580 );
buf \U$66023 ( \66518 , \66517_nG6eae );
not \U$66024 ( \66519 , \65145 );
xor \U$66025 ( \66520 , \65086 , \65087 );
not \U$66026 ( \66521 , \66520 );
or \U$66027 ( \66522 , \66519 , \66521 );
or \U$66028 ( \66523 , \66520 , \65145 );
nand \U$66029 ( \66524 , \66522 , \66523 );
_DC g6431 ( \66525_nG6431 , \66524 , \65580 );
buf \U$66030 ( \66526 , \66525_nG6431 );
endmodule

