//
// Conformal-LEC Version 20.10-d214 (03-Sep-2020)
//
module top(RIb54a900_11,RIb54a888_10,RIb54a810_9,RIb54a798_8,RIb54a720_7,RIb54a6a8_6,RIb54a630_5,RIb54a5b8_4,RIb54a540_3,
        RIb54a4c8_2,RIb54a450_1,RIb5517a0_247,RIb551980_251,RIb54ab58_16,RIb54abd0_17,RIb54aae0_15,RIb54aa68_14,RIb54a9f0_13,RIb551908_250,
        RIb551b60_255,RIb551ae8_254,RIb551f98_264,RIb551f20_263,RIb551cc8_258,RIb551c50_257,RIb551bd8_256,RIb551890_249,RIb551818_248,RIb551ea8_262,
        RIb551e30_261,RIb551db8_260,RIb551d40_259,RIb5519f8_252,RIb551a70_253,RIb54ad38_20,RIb54acc0_19,RIb54af18_24,RIb54aea0_23,RIb54b350_33,
        RIb54b2d8_32,RIb54af90_25,RIb54b008_26,RIb54b080_27,RIb54ac48_18,RIb54a978_12,RIb54b260_31,RIb54b1e8_30,RIb54b170_29,RIb54b0f8_28,
        RIb54adb0_21,RIb54ae28_22,RIb54b968_46,RIb54b8f0_45,RIb54b710_41,RIb54b698_40,RIb54bb48_50,RIb54bad0_49,RIb54b788_42,RIb54b620_39,
        RIb54b878_44,RIb54b800_43,RIb54b3c8_34,RIb54b4b8_36,RIb54b440_35,RIb54ba58_48,RIb54b9e0_47,RIb54b5a8_38,RIb54b530_37,RIb54bf08_58,
        RIb54be90_57,RIb54c160_63,RIb54bda0_55,RIb54bd28_54,RIb54bc38_52,RIb54be18_56,RIb54bcb0_53,RIb54c340_67,RIb54c0e8_62,RIb54bbc0_51,
        RIb54c250_65,RIb54c1d8_64,RIb54c070_61,RIb54bff8_60,RIb54c2c8_66,RIb54bf80_59,RIb54c8e0_79,RIb54c700_75,RIb54c778_76,RIb54c610_73,
        RIb54c520_71,RIb54c430_69,RIb54c598_72,RIb54c4a8_70,RIb54c868_78,RIb54c7f0_77,RIb54c3b8_68,RIb54cb38_84,RIb54cac0_83,RIb54ca48_82,
        RIb54c9d0_81,RIb54c958_80,RIb54c688_74,RIb54cca0_87,RIb54cc28_86,RIb54cef8_92,RIb54ce80_91,RIb54cd90_89,RIb54cfe8_94,RIb54d240_99,
        RIb54ce08_90,RIb54d330_101,RIb54d2b8_100,RIb54cbb0_85,RIb54d150_97,RIb54d1c8_98,RIb54d0d8_96,RIb54d060_95,RIb54cf70_93,RIb54cd18_88,
        RIb54d498_104,RIb54d420_103,RIb54d6f0_109,RIb54d678_108,RIb54db28_118,RIb54dab0_117,RIb54d768_110,RIb54d510_105,RIb54d858_112,RIb54d7e0_111,
        RIb54d3a8_102,RIb54da38_116,RIb54d9c0_115,RIb54d948_114,RIb54d8d0_113,RIb54d588_106,RIb54d600_107,RIb54dee8_126,RIb54de70_125,RIb54e050_129,
        RIb54dfd8_128,RIb54e140_131,RIb54e0c8_130,RIb54df60_127,RIb54dd08_122,RIb54e230_133,RIb54e1b8_132,RIb54dba0_119,RIb54dc90_121,RIb54dc18_120,
        RIb54e320_135,RIb54e2a8_134,RIb54dd80_123,RIb54ddf8_124,RIb54e500_139,RIb54e488_138,RIb54e6e0_143,RIb54e668_142,RIb54eb18_152,RIb54eaa0_151,
        RIb54e758_144,RIb54e7d0_145,RIb54e848_146,RIb54e410_137,RIb54e398_136,RIb54ea28_150,RIb54e9b0_149,RIb54e938_148,RIb54e8c0_147,RIb54e578_140,
        RIb54e5f0_141,RIb54eed8_160,RIb54ee60_159,RIb54f040_163,RIb54efc8_162,RIb54f220_167,RIb54f1a8_166,RIb54ef50_161,RIb54ede8_158,RIb54f130_165,
        RIb54f0b8_164,RIb54eb90_153,RIb54ec80_155,RIb54ec08_154,RIb54f310_169,RIb54f298_168,RIb54ed70_157,RIb54ecf8_156,RIb54f6d0_177,RIb54f658_176,
        RIb54f838_180,RIb54f7c0_179,RIb54f478_172,RIb54f400_171,RIb54fa18_184,RIb54f9a0_183,RIb54f928_182,RIb54f8b0_181,RIb54f388_170,RIb54f748_178,
        RIb54f5e0_175,RIb54fb08_186,RIb54fa90_185,RIb54f568_174,RIb54f4f0_173,RIb54ff40_195,RIb54fdd8_192,RIb54fc70_189,RIb54fbf8_188,RIb550300_203,
        RIb550288_202,RIb54fd60_191,RIb54fce8_190,RIb54fec8_194,RIb54fe50_193,RIb54fb80_187,RIb550120_199,RIb5500a8_198,RIb550030_197,RIb54ffb8_196,
        RIb550210_201,RIb550198_200,RIb550990_217,RIb550918_216,RIb550738_212,RIb5506c0_211,RIb550b70_221,RIb550af8_220,RIb5505d0_209,RIb550558_208,
        RIb5504e0_207,RIb550468_206,RIb5503f0_205,RIb550a80_219,RIb550a08_218,RIb5508a0_215,RIb550828_214,RIb5507b0_213,RIb550648_210,RIb550378_204,
        RIb550e40_227,RIb550eb8_228,RIb550f30_229,RIb550fa8_230,RIb550c60_223,RIb550cd8_224,RIb550d50_225,RIb550dc8_226,RIb5515c0_243,RIb551728_246,
        RIb551458_240,RIb5513e0_239,RIb5516b0_245,RIb551548_242,RIb5514d0_241,RIb550be8_222,RIb551200_235,RIb551368_238,RIb5512f0_237,RIb551188_234,
        RIb551110_233,RIb551638_244,RIb551020_231,RIb551278_236,RIb551098_232,RIb552448_274,RIb5526a0_279,RIb552628_278,RIb552010_265,RIb552268_270,
        RIb5525b0_277,RIb552538_276,RIb5521f0_269,RIb552178_268,RIb552718_280,RIb5524c0_275,RIb552358_272,RIb5522e0_271,RIb552100_267,RIb552088_266,
        RIb552790_281,RIb5523d0_273,RIb552c40_291,RIb552e98_296,RIb552e20_295,RIb552808_282,RIb552a60_287,RIb552da8_294,RIb552d30_293,RIb5529e8_286,
        RIb552970_285,RIb552f10_297,RIb552cb8_292,RIb552b50_289,RIb552ad8_288,RIb5528f8_284,RIb552880_283,RIb552f88_298,RIb552bc8_290,RIb553c30_325,
        RIb553e88_330,RIb553e10_329,RIb5537f8_316,RIb553a50_321,RIb553d98_328,RIb553d20_327,RIb5539d8_320,RIb553960_319,RIb553f00_331,RIb553ca8_326,
        RIb553b40_323,RIb553ac8_322,RIb5538e8_318,RIb553870_317,RIb553f78_332,RIb553bb8_324,RIb553618_312,RIb553780_315,RIb5534b0_309,RIb553438_308,
        RIb553708_314,RIb5535a0_311,RIb553528_310,RIb553000_299,RIb553258_304,RIb5533c0_307,RIb553348_306,RIb5531e0_303,RIb553168_302,RIb553690_313,
        RIb553078_300,RIb5532d0_305,RIb5530f0_301,RIb554068_334,RIb554680_347,RIb554608_346,RIb553ff0_333,RIb554248_338,RIb554590_345,RIb554518_344,
        RIb5541d0_337,RIb554158_336,RIb5542c0_339,RIb5540e0_335,RIb5543b0_341,RIb554338_340,RIb5544a0_343,RIb554428_342,RIb554770_349,RIb5546f8_348,
        RIb554ba8_358,RIb554d88_362,RIb554e00_363,RIb5549c8_354,RIb554950_353,RIb554d10_361,RIb554c98_360,RIb5547e8_350,RIb554ef0_365,RIb554e78_364,
        RIb554c20_359,RIb554ab8_356,RIb554a40_355,RIb5548d8_352,RIb554860_351,RIb554f68_366,RIb554b30_357,RIb555058_368,RIb555670_381,RIb5555f8_380,
        RIb554fe0_367,RIb555238_372,RIb555580_379,RIb555508_378,RIb5551c0_371,RIb555148_370,RIb5552b0_373,RIb5550d0_369,RIb5553a0_375,RIb555328_374,
        RIb555490_377,RIb555418_376,RIb555760_383,RIb5556e8_382,RIb5565e8_414,RIb556750_417,RIb556480_411,RIb556408_410,RIb5566d8_416,RIb556570_413,
        RIb5564f8_412,RIb555fd0_401,RIb556228_406,RIb556390_409,RIb556318_408,RIb5561b0_405,RIb556138_404,RIb556660_415,RIb556048_402,RIb5562a0_407,
        RIb5560c0_403,RIb555940_387,RIb555ee0_399,RIb555e68_398,RIb555aa8_390,RIb555a30_389,RIb5558c8_386,RIb555850_385,RIb5557d8_384,RIb555df0_397,
        RIb555b20_391,RIb5559b8_388,RIb555b98_392,RIb555c10_393,RIb555d00_395,RIb555c88_394,RIb555f58_400,RIb555d78_396,RIb557308_442,RIb557560_447,
        RIb5575d8_448,RIb5571a0_439,RIb557128_438,RIb5574e8_446,RIb557470_445,RIb556fc0_435,RIb557650_449,RIb557380_443,RIb5573f8_444,RIb557290_441,
        RIb557218_440,RIb5570b0_437,RIb557038_436,RIb557740_451,RIb5576c8_450,RIb556c00_427,RIb556ed0_433,RIb556e58_432,RIb5569a8_422,RIb556930_421,
        RIb5567c8_418,RIb556a20_423,RIb556d68_430,RIb556de0_431,RIb556cf0_429,RIb556c78_428,RIb556b10_425,RIb556a98_424,RIb5568b8_420,RIb556840_419,
        RIb556f48_434,RIb556b88_426,RIb557fb0_469,RIb5580a0_471,RIb5585c8_482,RIb558028_470,RIb558370_477,RIb5582f8_476,RIb558280_475,RIb558208_474,
        RIb558730_485,RIb558640_483,RIb558550_481,RIb558190_473,RIb558118_472,RIb558460_479,RIb5583e8_478,RIb5586b8_484,RIb5584d8_480,RIb557b00_459,
        RIb557830_453,RIb557ce0_463,RIb557bf0_461,RIb557b78_460,RIb557c68_462,RIb557a88_458,RIb557a10_457,RIb557f38_468,RIb557d58_464,RIb557dd0_465,
        RIb557998_456,RIb557920_455,RIb5577b8_452,RIb5578a8_454,RIb557ec0_467,RIb557e48_466,RIb559180_507,RIb5591f8_508,RIb558fa0_503,RIb559018_504,
        RIb559108_506,RIb559090_505,RIb559540_515,RIb5595b8_516,RIb559720_519,RIb5596a8_518,RIb559630_517,RIb559360_511,RIb5593d8_512,RIb5594c8_514,
        RIb559450_513,RIb5592e8_510,RIb559270_509,RIb558a00_491,RIb558988_490,RIb558910_489,RIb5587a8_486,RIb558cd0_497,RIb558c58_496,RIb558be0_495,
        RIb558898_488,RIb558820_487,RIb558d48_498,RIb558dc0_499,RIb558e38_500,RIb558a78_492,RIb558b68_494,RIb558af0_493,RIb558f28_502,RIb558eb0_501,
        RIb55a4b8_548,RIb55a440_547,RIb55a080_539,RIb55a008_538,RIb55a350_545,RIb55a3c8_546,RIb559f90_537,RIb55a2d8_544,RIb55a710_553,RIb55a698_552,
        RIb55a0f8_540,RIb55a170_541,RIb55a1e8_542,RIb55a530_549,RIb55a260_543,RIb55a620_551,RIb55a5a8_550,RIb559d38_532,RIb559db0_533,RIb559978_524,
        RIb5599f0_525,RIb559ae0_527,RIb559a68_526,RIb559cc0_531,RIb559c48_530,RIb559f18_536,RIb559b58_528,RIb559bd0_529,RIb559900_523,RIb559888_522,
        RIb559798_520,RIb559810_521,RIb559ea0_535,RIb559e28_534,RIb55ab48_562,RIb55aad0_561,RIb55a968_558,RIb55a8f0_557,RIb55aa58_560,RIb55a9e0_559,
        RIb55a878_556,RIb55a800_555,RIb55af08_570,RIb55ad28_566,RIb55ada0_567,RIb55a788_554,RIb55abc0_563,RIb55acb0_565,RIb55ac38_564,RIb55ae90_569,
        RIb55ae18_568,RIb55af80_571,RIb55aff8_572,RIb55b160_575,RIb55b1d8_576,RIb55b2c8_578,RIb55b250_577,RIb55b4a8_582,RIb55b430_581,RIb55b700_587,
        RIb55b340_579,RIb55b3b8_580,RIb55b520_583,RIb55b598_584,RIb55b0e8_574,RIb55b070_573,RIb55b688_586,RIb55b610_585,RIb55b778_588,RIb55bca0_599,
        RIb55bc28_598,RIb55bbb0_597,RIb55bb38_596,RIb55bac0_595,RIb55ba48_594,RIb55b9d0_593,RIb55b958_592,RIb55b8e0_591,RIb55b868_590,RIb55b7f0_589,
        RIb55c3a8_614,RIb55be80_603,RIb55bef8_604,RIb55be08_602,RIb55bd90_601,RIb55bd18_600,RIb55bf70_605,RIb55bfe8_606,RIb55c060_607,RIb55c0d8_608,
        RIb55c150_609,RIb55c1c8_610,RIb55c240_611,RIb55c2b8_612,RIb55c330_613,R_267_b942f48,R_268_b942ff0,R_269_b943098,R_26a_b943140,R_26b_b9431e8,
        R_26c_b943290,R_26d_b943338,R_26e_b9433e0,R_26f_b943488,R_270_b943530,R_271_b9435d8,R_272_b943680,R_273_b943728,R_274_b9437d0,R_275_b943878,
        R_276_b943920,R_277_b9439c8,R_278_b943a70,R_279_b943b18,R_27a_b943bc0,R_27b_b943c68,R_27c_b943d10,R_27d_b943db8,R_27e_b943e60,R_27f_b943f08,
        R_280_b943fb0,R_281_b944058,R_289_b944598,R_28a_b944640,R_28b_b9446e8,R_28c_b944790,R_28d_b944838,R_28e_b9448e0,R_28f_b944988,R_290_b944a30,
        R_291_b944ad8,R_292_b944b80,R_293_b944c28,R_294_b944cd0,R_295_b944d78,R_296_b944e20,R_297_b944ec8,R_298_b944f70,R_299_b945018,R_29a_b9450c0,
        R_29b_b945168,R_29c_b945210,R_29d_b9452b8,R_29e_b945360,R_29f_b945408,R_2a0_b9454b0,R_2a1_b945558,R_2a2_b945600,R_2a3_b9456a8);
input RIb54a900_11,RIb54a888_10,RIb54a810_9,RIb54a798_8,RIb54a720_7,RIb54a6a8_6,RIb54a630_5,RIb54a5b8_4,RIb54a540_3,
        RIb54a4c8_2,RIb54a450_1,RIb5517a0_247,RIb551980_251,RIb54ab58_16,RIb54abd0_17,RIb54aae0_15,RIb54aa68_14,RIb54a9f0_13,RIb551908_250,
        RIb551b60_255,RIb551ae8_254,RIb551f98_264,RIb551f20_263,RIb551cc8_258,RIb551c50_257,RIb551bd8_256,RIb551890_249,RIb551818_248,RIb551ea8_262,
        RIb551e30_261,RIb551db8_260,RIb551d40_259,RIb5519f8_252,RIb551a70_253,RIb54ad38_20,RIb54acc0_19,RIb54af18_24,RIb54aea0_23,RIb54b350_33,
        RIb54b2d8_32,RIb54af90_25,RIb54b008_26,RIb54b080_27,RIb54ac48_18,RIb54a978_12,RIb54b260_31,RIb54b1e8_30,RIb54b170_29,RIb54b0f8_28,
        RIb54adb0_21,RIb54ae28_22,RIb54b968_46,RIb54b8f0_45,RIb54b710_41,RIb54b698_40,RIb54bb48_50,RIb54bad0_49,RIb54b788_42,RIb54b620_39,
        RIb54b878_44,RIb54b800_43,RIb54b3c8_34,RIb54b4b8_36,RIb54b440_35,RIb54ba58_48,RIb54b9e0_47,RIb54b5a8_38,RIb54b530_37,RIb54bf08_58,
        RIb54be90_57,RIb54c160_63,RIb54bda0_55,RIb54bd28_54,RIb54bc38_52,RIb54be18_56,RIb54bcb0_53,RIb54c340_67,RIb54c0e8_62,RIb54bbc0_51,
        RIb54c250_65,RIb54c1d8_64,RIb54c070_61,RIb54bff8_60,RIb54c2c8_66,RIb54bf80_59,RIb54c8e0_79,RIb54c700_75,RIb54c778_76,RIb54c610_73,
        RIb54c520_71,RIb54c430_69,RIb54c598_72,RIb54c4a8_70,RIb54c868_78,RIb54c7f0_77,RIb54c3b8_68,RIb54cb38_84,RIb54cac0_83,RIb54ca48_82,
        RIb54c9d0_81,RIb54c958_80,RIb54c688_74,RIb54cca0_87,RIb54cc28_86,RIb54cef8_92,RIb54ce80_91,RIb54cd90_89,RIb54cfe8_94,RIb54d240_99,
        RIb54ce08_90,RIb54d330_101,RIb54d2b8_100,RIb54cbb0_85,RIb54d150_97,RIb54d1c8_98,RIb54d0d8_96,RIb54d060_95,RIb54cf70_93,RIb54cd18_88,
        RIb54d498_104,RIb54d420_103,RIb54d6f0_109,RIb54d678_108,RIb54db28_118,RIb54dab0_117,RIb54d768_110,RIb54d510_105,RIb54d858_112,RIb54d7e0_111,
        RIb54d3a8_102,RIb54da38_116,RIb54d9c0_115,RIb54d948_114,RIb54d8d0_113,RIb54d588_106,RIb54d600_107,RIb54dee8_126,RIb54de70_125,RIb54e050_129,
        RIb54dfd8_128,RIb54e140_131,RIb54e0c8_130,RIb54df60_127,RIb54dd08_122,RIb54e230_133,RIb54e1b8_132,RIb54dba0_119,RIb54dc90_121,RIb54dc18_120,
        RIb54e320_135,RIb54e2a8_134,RIb54dd80_123,RIb54ddf8_124,RIb54e500_139,RIb54e488_138,RIb54e6e0_143,RIb54e668_142,RIb54eb18_152,RIb54eaa0_151,
        RIb54e758_144,RIb54e7d0_145,RIb54e848_146,RIb54e410_137,RIb54e398_136,RIb54ea28_150,RIb54e9b0_149,RIb54e938_148,RIb54e8c0_147,RIb54e578_140,
        RIb54e5f0_141,RIb54eed8_160,RIb54ee60_159,RIb54f040_163,RIb54efc8_162,RIb54f220_167,RIb54f1a8_166,RIb54ef50_161,RIb54ede8_158,RIb54f130_165,
        RIb54f0b8_164,RIb54eb90_153,RIb54ec80_155,RIb54ec08_154,RIb54f310_169,RIb54f298_168,RIb54ed70_157,RIb54ecf8_156,RIb54f6d0_177,RIb54f658_176,
        RIb54f838_180,RIb54f7c0_179,RIb54f478_172,RIb54f400_171,RIb54fa18_184,RIb54f9a0_183,RIb54f928_182,RIb54f8b0_181,RIb54f388_170,RIb54f748_178,
        RIb54f5e0_175,RIb54fb08_186,RIb54fa90_185,RIb54f568_174,RIb54f4f0_173,RIb54ff40_195,RIb54fdd8_192,RIb54fc70_189,RIb54fbf8_188,RIb550300_203,
        RIb550288_202,RIb54fd60_191,RIb54fce8_190,RIb54fec8_194,RIb54fe50_193,RIb54fb80_187,RIb550120_199,RIb5500a8_198,RIb550030_197,RIb54ffb8_196,
        RIb550210_201,RIb550198_200,RIb550990_217,RIb550918_216,RIb550738_212,RIb5506c0_211,RIb550b70_221,RIb550af8_220,RIb5505d0_209,RIb550558_208,
        RIb5504e0_207,RIb550468_206,RIb5503f0_205,RIb550a80_219,RIb550a08_218,RIb5508a0_215,RIb550828_214,RIb5507b0_213,RIb550648_210,RIb550378_204,
        RIb550e40_227,RIb550eb8_228,RIb550f30_229,RIb550fa8_230,RIb550c60_223,RIb550cd8_224,RIb550d50_225,RIb550dc8_226,RIb5515c0_243,RIb551728_246,
        RIb551458_240,RIb5513e0_239,RIb5516b0_245,RIb551548_242,RIb5514d0_241,RIb550be8_222,RIb551200_235,RIb551368_238,RIb5512f0_237,RIb551188_234,
        RIb551110_233,RIb551638_244,RIb551020_231,RIb551278_236,RIb551098_232,RIb552448_274,RIb5526a0_279,RIb552628_278,RIb552010_265,RIb552268_270,
        RIb5525b0_277,RIb552538_276,RIb5521f0_269,RIb552178_268,RIb552718_280,RIb5524c0_275,RIb552358_272,RIb5522e0_271,RIb552100_267,RIb552088_266,
        RIb552790_281,RIb5523d0_273,RIb552c40_291,RIb552e98_296,RIb552e20_295,RIb552808_282,RIb552a60_287,RIb552da8_294,RIb552d30_293,RIb5529e8_286,
        RIb552970_285,RIb552f10_297,RIb552cb8_292,RIb552b50_289,RIb552ad8_288,RIb5528f8_284,RIb552880_283,RIb552f88_298,RIb552bc8_290,RIb553c30_325,
        RIb553e88_330,RIb553e10_329,RIb5537f8_316,RIb553a50_321,RIb553d98_328,RIb553d20_327,RIb5539d8_320,RIb553960_319,RIb553f00_331,RIb553ca8_326,
        RIb553b40_323,RIb553ac8_322,RIb5538e8_318,RIb553870_317,RIb553f78_332,RIb553bb8_324,RIb553618_312,RIb553780_315,RIb5534b0_309,RIb553438_308,
        RIb553708_314,RIb5535a0_311,RIb553528_310,RIb553000_299,RIb553258_304,RIb5533c0_307,RIb553348_306,RIb5531e0_303,RIb553168_302,RIb553690_313,
        RIb553078_300,RIb5532d0_305,RIb5530f0_301,RIb554068_334,RIb554680_347,RIb554608_346,RIb553ff0_333,RIb554248_338,RIb554590_345,RIb554518_344,
        RIb5541d0_337,RIb554158_336,RIb5542c0_339,RIb5540e0_335,RIb5543b0_341,RIb554338_340,RIb5544a0_343,RIb554428_342,RIb554770_349,RIb5546f8_348,
        RIb554ba8_358,RIb554d88_362,RIb554e00_363,RIb5549c8_354,RIb554950_353,RIb554d10_361,RIb554c98_360,RIb5547e8_350,RIb554ef0_365,RIb554e78_364,
        RIb554c20_359,RIb554ab8_356,RIb554a40_355,RIb5548d8_352,RIb554860_351,RIb554f68_366,RIb554b30_357,RIb555058_368,RIb555670_381,RIb5555f8_380,
        RIb554fe0_367,RIb555238_372,RIb555580_379,RIb555508_378,RIb5551c0_371,RIb555148_370,RIb5552b0_373,RIb5550d0_369,RIb5553a0_375,RIb555328_374,
        RIb555490_377,RIb555418_376,RIb555760_383,RIb5556e8_382,RIb5565e8_414,RIb556750_417,RIb556480_411,RIb556408_410,RIb5566d8_416,RIb556570_413,
        RIb5564f8_412,RIb555fd0_401,RIb556228_406,RIb556390_409,RIb556318_408,RIb5561b0_405,RIb556138_404,RIb556660_415,RIb556048_402,RIb5562a0_407,
        RIb5560c0_403,RIb555940_387,RIb555ee0_399,RIb555e68_398,RIb555aa8_390,RIb555a30_389,RIb5558c8_386,RIb555850_385,RIb5557d8_384,RIb555df0_397,
        RIb555b20_391,RIb5559b8_388,RIb555b98_392,RIb555c10_393,RIb555d00_395,RIb555c88_394,RIb555f58_400,RIb555d78_396,RIb557308_442,RIb557560_447,
        RIb5575d8_448,RIb5571a0_439,RIb557128_438,RIb5574e8_446,RIb557470_445,RIb556fc0_435,RIb557650_449,RIb557380_443,RIb5573f8_444,RIb557290_441,
        RIb557218_440,RIb5570b0_437,RIb557038_436,RIb557740_451,RIb5576c8_450,RIb556c00_427,RIb556ed0_433,RIb556e58_432,RIb5569a8_422,RIb556930_421,
        RIb5567c8_418,RIb556a20_423,RIb556d68_430,RIb556de0_431,RIb556cf0_429,RIb556c78_428,RIb556b10_425,RIb556a98_424,RIb5568b8_420,RIb556840_419,
        RIb556f48_434,RIb556b88_426,RIb557fb0_469,RIb5580a0_471,RIb5585c8_482,RIb558028_470,RIb558370_477,RIb5582f8_476,RIb558280_475,RIb558208_474,
        RIb558730_485,RIb558640_483,RIb558550_481,RIb558190_473,RIb558118_472,RIb558460_479,RIb5583e8_478,RIb5586b8_484,RIb5584d8_480,RIb557b00_459,
        RIb557830_453,RIb557ce0_463,RIb557bf0_461,RIb557b78_460,RIb557c68_462,RIb557a88_458,RIb557a10_457,RIb557f38_468,RIb557d58_464,RIb557dd0_465,
        RIb557998_456,RIb557920_455,RIb5577b8_452,RIb5578a8_454,RIb557ec0_467,RIb557e48_466,RIb559180_507,RIb5591f8_508,RIb558fa0_503,RIb559018_504,
        RIb559108_506,RIb559090_505,RIb559540_515,RIb5595b8_516,RIb559720_519,RIb5596a8_518,RIb559630_517,RIb559360_511,RIb5593d8_512,RIb5594c8_514,
        RIb559450_513,RIb5592e8_510,RIb559270_509,RIb558a00_491,RIb558988_490,RIb558910_489,RIb5587a8_486,RIb558cd0_497,RIb558c58_496,RIb558be0_495,
        RIb558898_488,RIb558820_487,RIb558d48_498,RIb558dc0_499,RIb558e38_500,RIb558a78_492,RIb558b68_494,RIb558af0_493,RIb558f28_502,RIb558eb0_501,
        RIb55a4b8_548,RIb55a440_547,RIb55a080_539,RIb55a008_538,RIb55a350_545,RIb55a3c8_546,RIb559f90_537,RIb55a2d8_544,RIb55a710_553,RIb55a698_552,
        RIb55a0f8_540,RIb55a170_541,RIb55a1e8_542,RIb55a530_549,RIb55a260_543,RIb55a620_551,RIb55a5a8_550,RIb559d38_532,RIb559db0_533,RIb559978_524,
        RIb5599f0_525,RIb559ae0_527,RIb559a68_526,RIb559cc0_531,RIb559c48_530,RIb559f18_536,RIb559b58_528,RIb559bd0_529,RIb559900_523,RIb559888_522,
        RIb559798_520,RIb559810_521,RIb559ea0_535,RIb559e28_534,RIb55ab48_562,RIb55aad0_561,RIb55a968_558,RIb55a8f0_557,RIb55aa58_560,RIb55a9e0_559,
        RIb55a878_556,RIb55a800_555,RIb55af08_570,RIb55ad28_566,RIb55ada0_567,RIb55a788_554,RIb55abc0_563,RIb55acb0_565,RIb55ac38_564,RIb55ae90_569,
        RIb55ae18_568,RIb55af80_571,RIb55aff8_572,RIb55b160_575,RIb55b1d8_576,RIb55b2c8_578,RIb55b250_577,RIb55b4a8_582,RIb55b430_581,RIb55b700_587,
        RIb55b340_579,RIb55b3b8_580,RIb55b520_583,RIb55b598_584,RIb55b0e8_574,RIb55b070_573,RIb55b688_586,RIb55b610_585,RIb55b778_588,RIb55bca0_599,
        RIb55bc28_598,RIb55bbb0_597,RIb55bb38_596,RIb55bac0_595,RIb55ba48_594,RIb55b9d0_593,RIb55b958_592,RIb55b8e0_591,RIb55b868_590,RIb55b7f0_589,
        RIb55c3a8_614,RIb55be80_603,RIb55bef8_604,RIb55be08_602,RIb55bd90_601,RIb55bd18_600,RIb55bf70_605,RIb55bfe8_606,RIb55c060_607,RIb55c0d8_608,
        RIb55c150_609,RIb55c1c8_610,RIb55c240_611,RIb55c2b8_612,RIb55c330_613;
output R_267_b942f48,R_268_b942ff0,R_269_b943098,R_26a_b943140,R_26b_b9431e8,R_26c_b943290,R_26d_b943338,R_26e_b9433e0,R_26f_b943488,
        R_270_b943530,R_271_b9435d8,R_272_b943680,R_273_b943728,R_274_b9437d0,R_275_b943878,R_276_b943920,R_277_b9439c8,R_278_b943a70,R_279_b943b18,
        R_27a_b943bc0,R_27b_b943c68,R_27c_b943d10,R_27d_b943db8,R_27e_b943e60,R_27f_b943f08,R_280_b943fb0,R_281_b944058,R_289_b944598,R_28a_b944640,
        R_28b_b9446e8,R_28c_b944790,R_28d_b944838,R_28e_b9448e0,R_28f_b944988,R_290_b944a30,R_291_b944ad8,R_292_b944b80,R_293_b944c28,R_294_b944cd0,
        R_295_b944d78,R_296_b944e20,R_297_b944ec8,R_298_b944f70,R_299_b945018,R_29a_b9450c0,R_29b_b945168,R_29c_b945210,R_29d_b9452b8,R_29e_b945360,
        R_29f_b945408,R_2a0_b9454b0,R_2a1_b945558,R_2a2_b945600,R_2a3_b9456a8;

wire \669_ZERO , \670_ONE , \671 , \672 , \673 , \674 , \675 , \676 , \677 ,
         \678 , \679 , \680 , \681 , \682 , \683 , \684 , \685 , \686 , \687 ,
         \688 , \689 , \690 , \691 , \692 , \693 , \694 , \695 , \696 , \697 ,
         \698 , \699 , \700 , \701 , \702 , \703 , \704 , \705 , \706 , \707 ,
         \708 , \709 , \710 , \711 , \712 , \713 , \714 , \715 , \716 , \717 ,
         \718 , \719 , \720 , \721 , \722 , \723 , \724 , \725 , \726 , \727 ,
         \728 , \729 , \730 , \731 , \732 , \733 , \734 , \735 , \736 , \737 ,
         \738 , \739 , \740 , \741 , \742 , \743 , \744 , \745 , \746 , \747 ,
         \748 , \749 , \750 , \751 , \752 , \753 , \754 , \755 , \756 , \757 ,
         \758 , \759 , \760 , \761 , \762 , \763 , \764 , \765 , \766 , \767 ,
         \768_nR12c0 , \769 , \770 , \771 , \772 , \773 , \774 , \775 , \776 , \777 ,
         \778 , \779 , \780 , \781 , \782 , \783 , \784 , \785 , \786 , \787 ,
         \788 , \789 , \790 , \791 , \792 , \793 , \794 , \795 , \796 , \797 ,
         \798 , \799 , \800 , \801 , \802 , \803 , \804_nR10db , \805 , \806 , \807 ,
         \808 , \809 , \810 , \811 , \812 , \813 , \814 , \815 , \816 , \817 ,
         \818 , \819 , \820 , \821 , \822 , \823 , \824 , \825 , \826 , \827 ,
         \828 , \829 , \830 , \831 , \832 , \833 , \834 , \835 , \836 , \837 ,
         \838 , \839 , \840_nR10d9 , \841 , \842 , \843 , \844 , \845 , \846 , \847 ,
         \848 , \849 , \850 , \851 , \852 , \853 , \854 , \855 , \856 , \857 ,
         \858 , \859 , \860 , \861 , \862 , \863 , \864 , \865 , \866 , \867 ,
         \868 , \869 , \870 , \871 , \872 , \873 , \874 , \875 , \876_nRf20 , \877 ,
         \878 , \879 , \880 , \881 , \882 , \883 , \884 , \885 , \886 , \887 ,
         \888 , \889 , \890 , \891 , \892 , \893 , \894 , \895 , \896 , \897 ,
         \898 , \899 , \900 , \901 , \902 , \903 , \904 , \905 , \906 , \907 ,
         \908 , \909 , \910 , \911 , \912_nRf1e , \913 , \914 , \915 , \916 , \917 ,
         \918 , \919 , \920 , \921 , \922 , \923 , \924 , \925 , \926 , \927 ,
         \928 , \929 , \930 , \931 , \932 , \933 , \934 , \935 , \936 , \937 ,
         \938 , \939 , \940 , \941 , \942 , \943 , \944 , \945 , \946 , \947 ,
         \948_nRda0 , \949 , \950 , \951 , \952 , \953 , \954 , \955 , \956 , \957 ,
         \958 , \959 , \960 , \961 , \962 , \963 , \964 , \965 , \966 , \967 ,
         \968 , \969 , \970 , \971 , \972 , \973 , \974 , \975 , \976 , \977 ,
         \978 , \979 , \980 , \981 , \982 , \983 , \984_nRd9e , \985 , \986 , \987 ,
         \988 , \989 , \990 , \991 , \992 , \993 , \994 , \995 , \996 , \997 ,
         \998 , \999 , \1000 , \1001 , \1002 , \1003 , \1004 , \1005 , \1006 , \1007 ,
         \1008 , \1009 , \1010 , \1011 , \1012 , \1013 , \1014 , \1015 , \1016 , \1017 ,
         \1018 , \1019 , \1020_nRc66 , \1021 , \1022 , \1023 , \1024 , \1025 , \1026 , \1027 ,
         \1028 , \1029 , \1030 , \1031 , \1032 , \1033 , \1034 , \1035 , \1036 , \1037 ,
         \1038 , \1039 , \1040 , \1041 , \1042 , \1043 , \1044 , \1045 , \1046 , \1047 ,
         \1048 , \1049 , \1050 , \1051 , \1052 , \1053 , \1054 , \1055 , \1056_nRc64 , \1057 ,
         \1058 , \1059 , \1060 , \1061 , \1062 , \1063 , \1064 , \1065 , \1066 , \1067 ,
         \1068 , \1069 , \1070 , \1071 , \1072 , \1073 , \1074 , \1075 , \1076 , \1077 ,
         \1078 , \1079 , \1080 , \1081 , \1082 , \1083 , \1084 , \1085 , \1086 , \1087 ,
         \1088 , \1089 , \1090 , \1091 , \1092_nRb7a , \1093 , \1094 , \1095 , \1096 , \1097 ,
         \1098 , \1099 , \1100 , \1101 , \1102 , \1103 , \1104 , \1105 , \1106 , \1107 ,
         \1108 , \1109 , \1110 , \1111 , \1112 , \1113 , \1114 , \1115 , \1116 , \1117 ,
         \1118 , \1119 , \1120 , \1121 , \1122 , \1123 , \1124 , \1125 , \1126 , \1127 ,
         \1128_nRb7c , \1129 , \1130 , \1131 , \1132 , \1133 , \1134 , \1135 , \1136 , \1137 ,
         \1138 , \1139 , \1140 , \1141 , \1142 , \1143 , \1144 , \1145 , \1146 , \1147 ,
         \1148 , \1149 , \1150 , \1151 , \1152 , \1153 , \1154 , \1155 , \1156 , \1157 ,
         \1158 , \1159_nR9e7 , \1160 , \1161 , \1162 , \1163 , \1164 , \1165 , \1166 , \1167 ,
         \1168 , \1169 , \1170 , \1171 , \1172 , \1173 , \1174 , \1175 , \1176 , \1177 ,
         \1178 , \1179 , \1180 , \1181 , \1182 , \1183 , \1184 , \1185 , \1186 , \1187 ,
         \1188 , \1189 , \1190_nR9e5 , \1191 , \1192 , \1193 , \1194 , \1195 , \1196 , \1197 ,
         \1198 , \1199 , \1200 , \1201 , \1202 , \1203 , \1204 , \1205 , \1206 , \1207 ,
         \1208 , \1209 , \1210 , \1211 , \1212 , \1213 , \1214 , \1215 , \1216 , \1217 ,
         \1218 , \1219 , \1220 , \1221 , \1222 , \1223 , \1224 , \1225 , \1226 , \1227 ,
         \1228 , \1229 , \1230 , \1231 , \1232 , \1233 , \1234 , \1235 , \1236 , \1237 ,
         \1238 , \1239 , \1240 , \1241 , \1242 , \1243 , \1244 , \1245 , \1246 , \1247 ,
         \1248 , \1249 , \1250 , \1251 , \1252 , \1253 , \1254 , \1255 , \1256 , \1257 ,
         \1258 , \1259 , \1260 , \1261 , \1262 , \1263 , \1264 , \1265 , \1266 , \1267 ,
         \1268 , \1269 , \1270 , \1271 , \1272 , \1273 , \1274 , \1275 , \1276 , \1277 ,
         \1278 , \1279 , \1280 , \1281 , \1282 , \1283 , \1284 , \1285 , \1286 , \1287 ,
         \1288 , \1289 , \1290 , \1291 , \1292 , \1293 , \1294 , \1295 , \1296 , \1297 ,
         \1298 , \1299 , \1300 , \1301 , \1302 , \1303 , \1304 , \1305 , \1306 , \1307 ,
         \1308 , \1309 , \1310 , \1311 , \1312 , \1313 , \1314 , \1315 , \1316 , \1317 ,
         \1318 , \1319 , \1320 , \1321_nR1933 , \1322 , \1323 , \1324 , \1325 , \1326 , \1327 ,
         \1328 , \1329 , \1330 , \1331 , \1332 , \1333 , \1334 , \1335 , \1336 , \1337 ,
         \1338 , \1339 , \1340 , \1341 , \1342 , \1343 , \1344 , \1345 , \1346 , \1347 ,
         \1348 , \1349 , \1350 , \1351 , \1352 , \1353 , \1354 , \1355 , \1356 , \1357 ,
         \1358 , \1359 , \1360 , \1361 , \1362 , \1363 , \1364_nR1a4f , \1365 , \1366 , \1367 ,
         \1368 , \1369 , \1370 , \1371 , \1372 , \1373 , \1374 , \1375 , \1376 , \1377 ,
         \1378 , \1379 , \1380 , \1381 , \1382 , \1383 , \1384 , \1385 , \1386 , \1387 ,
         \1388 , \1389 , \1390 , \1391 , \1392 , \1393 , \1394 , \1395 , \1396 , \1397 ,
         \1398 , \1399 , \1400 , \1401 , \1402 , \1403 , \1404 , \1405 , \1406 , \1407 ,
         \1408 , \1409 , \1410 , \1411 , \1412 , \1413 , \1414 , \1415 , \1416 , \1417 ,
         \1418 , \1419 , \1420 , \1421 , \1422 , \1423_nR183c , \1424 , \1425 , \1426 , \1427 ,
         \1428 , \1429 , \1430 , \1431 , \1432 , \1433 , \1434 , \1435 , \1436 , \1437 ,
         \1438 , \1439 , \1440 , \1441 , \1442 , \1443 , \1444 , \1445 , \1446 , \1447 ,
         \1448 , \1449 , \1450 , \1451 , \1452 , \1453 , \1454 , \1455 , \1456 , \1457 ,
         \1458 , \1459 , \1460 , \1461 , \1462 , \1463 , \1464 , \1465 , \1466 , \1467 ,
         \1468 , \1469 , \1470 , \1471 , \1472 , \1473 , \1474 , \1475 , \1476 , \1477 ,
         \1478 , \1479 , \1480 , \1481 , \1482 , \1483 , \1484 , \1485 , \1486 , \1487 ,
         \1488 , \1489 , \1490 , \1491 , \1492 , \1493 , \1494_nR16fe , \1495 , \1496 , \1497 ,
         \1498 , \1499 , \1500 , \1501 , \1502 , \1503 , \1504 , \1505 , \1506 , \1507 ,
         \1508 , \1509 , \1510 , \1511 , \1512 , \1513 , \1514 , \1515 , \1516 , \1517 ,
         \1518 , \1519 , \1520 , \1521 , \1522 , \1523 , \1524 , \1525 , \1526 , \1527 ,
         \1528 , \1529 , \1530 , \1531 , \1532 , \1533 , \1534 , \1535 , \1536 , \1537 ,
         \1538 , \1539 , \1540 , \1541 , \1542 , \1543 , \1544 , \1545 , \1546 , \1547 ,
         \1548 , \1549 , \1550 , \1551 , \1552 , \1553 , \1554 , \1555 , \1556 , \1557 ,
         \1558 , \1559 , \1560 , \1561 , \1562 , \1563 , \1564 , \1565 , \1566 , \1567 ,
         \1568 , \1569 , \1570 , \1571 , \1572 , \1573 , \1574 , \1575 , \1576 , \1577 ,
         \1578_nR1611 , \1579 , \1580 , \1581 , \1582 , \1583 , \1584 , \1585 , \1586 , \1587 ,
         \1588 , \1589 , \1590 , \1591 , \1592 , \1593 , \1594 , \1595 , \1596 , \1597 ,
         \1598 , \1599 , \1600 , \1601 , \1602 , \1603 , \1604 , \1605 , \1606 , \1607 ,
         \1608 , \1609 , \1610 , \1611 , \1612 , \1613 , \1614 , \1615 , \1616 , \1617 ,
         \1618 , \1619 , \1620 , \1621 , \1622 , \1623 , \1624 , \1625 , \1626_nR14f1 , \1627 ,
         \1628 , \1629 , \1630 , \1631 , \1632 , \1633 , \1634 , \1635 , \1636 , \1637 ,
         \1638 , \1639 , \1640 , \1641 , \1642 , \1643 , \1644 , \1645 , \1646 , \1647 ,
         \1648 , \1649 , \1650 , \1651 , \1652 , \1653 , \1654 , \1655 , \1656 , \1657 ,
         \1658 , \1659 , \1660 , \1661 , \1662 , \1663 , \1664 , \1665 , \1666 , \1667 ,
         \1668 , \1669 , \1670 , \1671 , \1672 , \1673 , \1674 , \1675 , \1676 , \1677 ,
         \1678 , \1679 , \1680 , \1681 , \1682 , \1683 , \1684 , \1685 , \1686 , \1687 ,
         \1688 , \1689 , \1690 , \1691 , \1692 , \1693 , \1694 , \1695 , \1696 , \1697 ,
         \1698 , \1699 , \1700 , \1701 , \1702 , \1703 , \1704 , \1705 , \1706 , \1707 ,
         \1708 , \1709 , \1710 , \1711 , \1712 , \1713 , \1714 , \1715 , \1716 , \1717 ,
         \1718 , \1719 , \1720 , \1721 , \1722 , \1723 , \1724 , \1725 , \1726 , \1727 ,
         \1728_nR12de , \1729 , \1730 , \1731 , \1732 , \1733 , \1734 , \1735 , \1736 , \1737 ,
         \1738 , \1739 , \1740 , \1741 , \1742 , \1743 , \1744 , \1745 , \1746 , \1747 ,
         \1748 , \1749 , \1750 , \1751 , \1752 , \1753 , \1754 , \1755 , \1756 , \1757 ,
         \1758 , \1759 , \1760 , \1761_nR13ee , \1762 , \1763 , \1764 , \1765 , \1766 , \1767 ,
         \1768 , \1769 , \1770 , \1771 , \1772 , \1773 , \1774 , \1775 , \1776 , \1777 ,
         \1778 , \1779 , \1780 , \1781 , \1782 , \1783 , \1784 , \1785 , \1786 , \1787 ,
         \1788 , \1789 , \1790 , \1791 , \1792 , \1793 , \1794 , \1795 , \1796 , \1797 ,
         \1798 , \1799 , \1800 , \1801 , \1802 , \1803 , \1804 , \1805 , \1806 , \1807 ,
         \1808 , \1809 , \1810 , \1811 , \1812 , \1813 , \1814 , \1815 , \1816 , \1817 ,
         \1818 , \1819 , \1820 , \1821 , \1822 , \1823 , \1824 , \1825 , \1826 , \1827 ,
         \1828 , \1829 , \1830 , \1831 , \1832 , \1833 , \1834 , \1835 , \1836 , \1837 ,
         \1838 , \1839 , \1840 , \1841 , \1842 , \1843 , \1844 , \1845 , \1846 , \1847 ,
         \1848 , \1849 , \1850 , \1851 , \1852 , \1853 , \1854 , \1855 , \1856 , \1857 ,
         \1858 , \1859 , \1860 , \1861 , \1862 , \1863 , \1864 , \1865 , \1866 , \1867 ,
         \1868 , \1869 , \1870 , \1871 , \1872 , \1873 , \1874 , \1875 , \1876 , \1877 ,
         \1878 , \1879 , \1880 , \1881 , \1882 , \1883 , \1884 , \1885 , \1886 , \1887 ,
         \1888 , \1889 , \1890 , \1891 , \1892 , \1893 , \1894 , \1895 , \1896 , \1897 ,
         \1898 , \1899 , \1900 , \1901 , \1902 , \1903 , \1904 , \1905 , \1906 , \1907_nR1200 ,
         \1908 , \1909 , \1910 , \1911 , \1912 , \1913 , \1914 , \1915 , \1916 , \1917 ,
         \1918 , \1919 , \1920 , \1921 , \1922 , \1923 , \1924 , \1925 , \1926 , \1927 ,
         \1928 , \1929 , \1930 , \1931 , \1932 , \1933 , \1934 , \1935 , \1936 , \1937 ,
         \1938 , \1939 , \1940 , \1941 , \1942 , \1943 , \1944 , \1945 , \1946 , \1947 ,
         \1948 , \1949 , \1950 , \1951 , \1952 , \1953 , \1954 , \1955 , \1956 , \1957 ,
         \1958 , \1959 , \1960 , \1961 , \1962 , \1963 , \1964 , \1965 , \1966 , \1967 ,
         \1968 , \1969 , \1970 , \1971 , \1972 , \1973 , \1974 , \1975 , \1976 , \1977 ,
         \1978 , \1979 , \1980 , \1981 , \1982 , \1983 , \1984 , \1985 , \1986 , \1987 ,
         \1988 , \1989 , \1990 , \1991 , \1992 , \1993 , \1994 , \1995 , \1996 , \1997 ,
         \1998 , \1999 , \2000 , \2001 , \2002 , \2003 , \2004 , \2005 , \2006 , \2007 ,
         \2008 , \2009 , \2010 , \2011 , \2012 , \2013 , \2014 , \2015 , \2016 , \2017 ,
         \2018 , \2019 , \2020 , \2021 , \2022 , \2023 , \2024 , \2025 , \2026 , \2027 ,
         \2028 , \2029 , \2030 , \2031 , \2032 , \2033 , \2034 , \2035 , \2036 , \2037 ,
         \2038 , \2039 , \2040 , \2041 , \2042 , \2043 , \2044 , \2045 , \2046 , \2047 ,
         \2048 , \2049 , \2050 , \2051 , \2052 , \2053 , \2054 , \2055 , \2056 , \2057 ,
         \2058 , \2059 , \2060 , \2061 , \2062 , \2063 , \2064 , \2065 , \2066 , \2067 ,
         \2068 , \2069 , \2070 , \2071 , \2072 , \2073 , \2074 , \2075 , \2076 , \2077 ,
         \2078 , \2079 , \2080 , \2081 , \2082 , \2083 , \2084 , \2085 , \2086 , \2087 ,
         \2088 , \2089 , \2090 , \2091 , \2092 , \2093 , \2094 , \2095 , \2096 , \2097 ,
         \2098 , \2099 , \2100 , \2101 , \2102 , \2103 , \2104 , \2105 , \2106 , \2107 ,
         \2108 , \2109 , \2110 , \2111 , \2112 , \2113 , \2114 , \2115 , \2116 , \2117 ,
         \2118 , \2119 , \2120 , \2121 , \2122 , \2123 , \2124 , \2125 , \2126 , \2127 ,
         \2128 , \2129 , \2130 , \2131 , \2132_nR10f9 , \2133 , \2134 , \2135 , \2136 , \2137 ,
         \2138 , \2139 , \2140 , \2141 , \2142 , \2143 , \2144 , \2145 , \2146 , \2147 ,
         \2148 , \2149 , \2150 , \2151 , \2152 , \2153 , \2154 , \2155 , \2156 , \2157 ,
         \2158 , \2159 , \2160 , \2161 , \2162 , \2163 , \2164 , \2165 , \2166 , \2167 ,
         \2168 , \2169 , \2170 , \2171 , \2172 , \2173 , \2174 , \2175 , \2176 , \2177 ,
         \2178 , \2179 , \2180 , \2181 , \2182 , \2183 , \2184 , \2185 , \2186 , \2187 ,
         \2188 , \2189 , \2190 , \2191 , \2192 , \2193 , \2194 , \2195 , \2196 , \2197 ,
         \2198 , \2199 , \2200 , \2201 , \2202 , \2203 , \2204 , \2205 , \2206 , \2207 ,
         \2208 , \2209 , \2210 , \2211 , \2212 , \2213 , \2214 , \2215 , \2216 , \2217 ,
         \2218 , \2219 , \2220 , \2221 , \2222 , \2223 , \2224 , \2225 , \2226 , \2227 ,
         \2228 , \2229 , \2230 , \2231 , \2232 , \2233 , \2234 , \2235 , \2236 , \2237 ,
         \2238 , \2239 , \2240 , \2241 , \2242 , \2243 , \2244 , \2245 , \2246 , \2247 ,
         \2248 , \2249 , \2250 , \2251 , \2252 , \2253 , \2254 , \2255 , \2256 , \2257 ,
         \2258 , \2259 , \2260 , \2261 , \2262 , \2263 , \2264 , \2265 , \2266 , \2267 ,
         \2268 , \2269 , \2270 , \2271 , \2272 , \2273 , \2274 , \2275 , \2276 , \2277 ,
         \2278 , \2279 , \2280 , \2281 , \2282 , \2283_nR101a , \2284 , \2285 , \2286 , \2287 ,
         \2288 , \2289 , \2290 , \2291 , \2292 , \2293 , \2294 , \2295 , \2296 , \2297 ,
         \2298 , \2299 , \2300 , \2301 , \2302 , \2303 , \2304 , \2305 , \2306 , \2307 ,
         \2308 , \2309 , \2310 , \2311 , \2312 , \2313 , \2314 , \2315 , \2316 , \2317 ,
         \2318 , \2319 , \2320 , \2321 , \2322 , \2323 , \2324 , \2325 , \2326 , \2327 ,
         \2328 , \2329 , \2330 , \2331 , \2332 , \2333 , \2334 , \2335 , \2336 , \2337 ,
         \2338 , \2339 , \2340 , \2341 , \2342 , \2343 , \2344 , \2345 , \2346 , \2347 ,
         \2348 , \2349 , \2350 , \2351 , \2352 , \2353 , \2354 , \2355 , \2356 , \2357 ,
         \2358 , \2359 , \2360 , \2361 , \2362 , \2363 , \2364 , \2365 , \2366 , \2367 ,
         \2368 , \2369 , \2370 , \2371 , \2372 , \2373 , \2374 , \2375 , \2376 , \2377 ,
         \2378 , \2379 , \2380 , \2381 , \2382 , \2383 , \2384 , \2385 , \2386 , \2387 ,
         \2388 , \2389 , \2390 , \2391 , \2392 , \2393 , \2394 , \2395 , \2396 , \2397 ,
         \2398 , \2399 , \2400 , \2401 , \2402 , \2403 , \2404 , \2405 , \2406 , \2407_nRf3e ,
         \2408 , \2409 , \2410 , \2411 , \2412 , \2413 , \2414 , \2415 , \2416 , \2417 ,
         \2418 , \2419 , \2420 , \2421 , \2422 , \2423 , \2424 , \2425 , \2426 , \2427 ,
         \2428 , \2429 , \2430 , \2431 , \2432 , \2433 , \2434 , \2435 , \2436 , \2437 ,
         \2438 , \2439 , \2440 , \2441 , \2442 , \2443 , \2444 , \2445 , \2446 , \2447 ,
         \2448 , \2449 , \2450 , \2451 , \2452 , \2453 , \2454 , \2455 , \2456 , \2457 ,
         \2458 , \2459 , \2460 , \2461 , \2462 , \2463 , \2464 , \2465 , \2466 , \2467 ,
         \2468 , \2469 , \2470 , \2471 , \2472 , \2473 , \2474 , \2475 , \2476 , \2477 ,
         \2478 , \2479 , \2480_nRe8d , \2481 , \2482 , \2483 , \2484 , \2485 , \2486 , \2487 ,
         \2488 , \2489 , \2490 , \2491 , \2492 , \2493 , \2494 , \2495 , \2496 , \2497 ,
         \2498 , \2499 , \2500 , \2501 , \2502 , \2503 , \2504 , \2505 , \2506 , \2507 ,
         \2508 , \2509 , \2510 , \2511 , \2512 , \2513 , \2514 , \2515 , \2516 , \2517 ,
         \2518 , \2519 , \2520 , \2521 , \2522 , \2523 , \2524 , \2525 , \2526 , \2527 ,
         \2528 , \2529 , \2530 , \2531 , \2532 , \2533 , \2534 , \2535 , \2536 , \2537 ,
         \2538 , \2539 , \2540 , \2541 , \2542 , \2543 , \2544 , \2545 , \2546 , \2547 ,
         \2548 , \2549 , \2550 , \2551 , \2552 , \2553 , \2554 , \2555 , \2556 , \2557 ,
         \2558 , \2559 , \2560 , \2561 , \2562 , \2563 , \2564 , \2565 , \2566 , \2567 ,
         \2568 , \2569 , \2570_nRdbd , \2571 , \2572 , \2573 , \2574 , \2575 , \2576 , \2577 ,
         \2578 , \2579 , \2580 , \2581 , \2582 , \2583 , \2584 , \2585 , \2586 , \2587 ,
         \2588 , \2589 , \2590 , \2591 , \2592 , \2593 , \2594 , \2595 , \2596 , \2597 ,
         \2598 , \2599 , \2600 , \2601 , \2602 , \2603 , \2604 , \2605 , \2606 , \2607 ,
         \2608 , \2609 , \2610 , \2611 , \2612 , \2613 , \2614 , \2615 , \2616 , \2617 ,
         \2618 , \2619 , \2620 , \2621 , \2622 , \2623 , \2624 , \2625 , \2626 , \2627 ,
         \2628 , \2629 , \2630 , \2631 , \2632 , \2633 , \2634 , \2635 , \2636 , \2637 ,
         \2638 , \2639 , \2640 , \2641 , \2642 , \2643 , \2644 , \2645 , \2646 , \2647 ,
         \2648 , \2649 , \2650 , \2651 , \2652 , \2653 , \2654 , \2655 , \2656 , \2657 ,
         \2658 , \2659 , \2660 , \2661 , \2662 , \2663 , \2664 , \2665 , \2666 , \2667 ,
         \2668 , \2669 , \2670 , \2671 , \2672 , \2673 , \2674 , \2675 , \2676 , \2677 ,
         \2678 , \2679 , \2680 , \2681 , \2682 , \2683 , \2684 , \2685 , \2686 , \2687 ,
         \2688 , \2689 , \2690 , \2691 , \2692 , \2693 , \2694 , \2695 , \2696 , \2697 ,
         \2698 , \2699 , \2700 , \2701 , \2702 , \2703 , \2704 , \2705 , \2706 , \2707 ,
         \2708 , \2709 , \2710 , \2711 , \2712 , \2713 , \2714 , \2715 , \2716 , \2717 ,
         \2718 , \2719 , \2720 , \2721 , \2722 , \2723 , \2724 , \2725 , \2726 , \2727 ,
         \2728 , \2729 , \2730 , \2731 , \2732 , \2733 , \2734 , \2735 , \2736 , \2737 ,
         \2738 , \2739 , \2740 , \2741 , \2742 , \2743 , \2744 , \2745 , \2746 , \2747 ,
         \2748 , \2749 , \2750 , \2751 , \2752 , \2753 , \2754 , \2755 , \2756 , \2757 ,
         \2758 , \2759 , \2760 , \2761 , \2762 , \2763 , \2764_nRd2b , \2765 , \2766 , \2767 ,
         \2768 , \2769 , \2770 , \2771 , \2772 , \2773 , \2774 , \2775 , \2776 , \2777 ,
         \2778 , \2779 , \2780 , \2781 , \2782 , \2783 , \2784 , \2785 , \2786 , \2787 ,
         \2788 , \2789 , \2790 , \2791 , \2792 , \2793 , \2794 , \2795 , \2796 , \2797 ,
         \2798 , \2799 , \2800 , \2801 , \2802 , \2803 , \2804 , \2805 , \2806 , \2807 ,
         \2808 , \2809 , \2810 , \2811 , \2812 , \2813 , \2814 , \2815 , \2816 , \2817_nRc84 ,
         \2818 , \2819 , \2820 , \2821 , \2822 , \2823 , \2824 , \2825 , \2826 , \2827 ,
         \2828 , \2829 , \2830 , \2831 , \2832 , \2833 , \2834 , \2835 , \2836 , \2837 ,
         \2838 , \2839 , \2840 , \2841 , \2842 , \2843 , \2844 , \2845 , \2846 , \2847 ,
         \2848 , \2849 , \2850 , \2851 , \2852 , \2853 , \2854 , \2855 , \2856 , \2857 ,
         \2858 , \2859 , \2860 , \2861 , \2862 , \2863 , \2864 , \2865 , \2866 , \2867 ,
         \2868 , \2869 , \2870 , \2871 , \2872 , \2873 , \2874 , \2875 , \2876 , \2877 ,
         \2878 , \2879 , \2880 , \2881 , \2882 , \2883 , \2884 , \2885 , \2886 , \2887 ,
         \2888 , \2889 , \2890 , \2891 , \2892 , \2893 , \2894 , \2895 , \2896 , \2897 ,
         \2898 , \2899 , \2900 , \2901 , \2902 , \2903 , \2904 , \2905 , \2906 , \2907 ,
         \2908 , \2909 , \2910 , \2911 , \2912 , \2913 , \2914 , \2915 , \2916 , \2917 ,
         \2918 , \2919 , \2920 , \2921 , \2922 , \2923 , \2924 , \2925 , \2926 , \2927 ,
         \2928 , \2929 , \2930 , \2931 , \2932 , \2933 , \2934 , \2935 , \2936 , \2937 ,
         \2938 , \2939 , \2940 , \2941 , \2942 , \2943 , \2944 , \2945 , \2946 , \2947 ,
         \2948 , \2949 , \2950 , \2951 , \2952 , \2953 , \2954 , \2955 , \2956 , \2957 ,
         \2958 , \2959 , \2960 , \2961 , \2962 , \2963 , \2964 , \2965 , \2966 , \2967 ,
         \2968 , \2969 , \2970 , \2971 , \2972 , \2973 , \2974 , \2975 , \2976 , \2977 ,
         \2978 , \2979 , \2980 , \2981 , \2982 , \2983 , \2984 , \2985 , \2986 , \2987 ,
         \2988 , \2989 , \2990 , \2991 , \2992 , \2993 , \2994 , \2995 , \2996 , \2997 ,
         \2998 , \2999 , \3000 , \3001 , \3002 , \3003 , \3004 , \3005 , \3006 , \3007 ,
         \3008 , \3009 , \3010_nRc05 , \3011 , \3012 , \3013 , \3014 , \3015 , \3016 , \3017 ,
         \3018 , \3019 , \3020 , \3021 , \3022 , \3023 , \3024 , \3025 , \3026 , \3027 ,
         \3028 , \3029 , \3030 , \3031 , \3032 , \3033 , \3034 , \3035 , \3036 , \3037 ,
         \3038 , \3039 , \3040 , \3041 , \3042 , \3043 , \3044 , \3045 , \3046 , \3047 ,
         \3048 , \3049 , \3050 , \3051 , \3052 , \3053 , \3054 , \3055 , \3056 , \3057 ,
         \3058 , \3059 , \3060 , \3061 , \3062 , \3063 , \3064 , \3065 , \3066 , \3067 ,
         \3068 , \3069 , \3070 , \3071 , \3072 , \3073 , \3074 , \3075 , \3076 , \3077 ,
         \3078 , \3079 , \3080 , \3081 , \3082 , \3083 , \3084 , \3085 , \3086 , \3087 ,
         \3088 , \3089 , \3090 , \3091 , \3092 , \3093 , \3094 , \3095 , \3096 , \3097 ,
         \3098 , \3099 , \3100 , \3101 , \3102 , \3103 , \3104 , \3105 , \3106 , \3107 ,
         \3108 , \3109 , \3110 , \3111 , \3112 , \3113 , \3114 , \3115 , \3116 , \3117 ,
         \3118 , \3119 , \3120 , \3121 , \3122 , \3123 , \3124 , \3125 , \3126 , \3127_nRb78 ,
         \3128 , \3129 , \3130 , \3131 , \3132 , \3133 , \3134 , \3135 , \3136 , \3137 ,
         \3138 , \3139 , \3140 , \3141 , \3142 , \3143 , \3144 , \3145 , \3146 , \3147 ,
         \3148 , \3149 , \3150 , \3151 , \3152 , \3153 , \3154 , \3155 , \3156 , \3157 ,
         \3158 , \3159 , \3160 , \3161 , \3162 , \3163 , \3164 , \3165 , \3166 , \3167 ,
         \3168 , \3169 , \3170 , \3171 , \3172 , \3173 , \3174 , \3175 , \3176 , \3177 ,
         \3178 , \3179 , \3180 , \3181 , \3182 , \3183 , \3184 , \3185 , \3186 , \3187 ,
         \3188 , \3189 , \3190 , \3191 , \3192 , \3193 , \3194 , \3195 , \3196 , \3197 ,
         \3198 , \3199 , \3200 , \3201 , \3202 , \3203 , \3204 , \3205 , \3206 , \3207 ,
         \3208 , \3209 , \3210 , \3211 , \3212 , \3213 , \3214 , \3215 , \3216 , \3217 ,
         \3218 , \3219 , \3220 , \3221 , \3222 , \3223 , \3224 , \3225 , \3226 , \3227 ,
         \3228 , \3229 , \3230 , \3231 , \3232 , \3233 , \3234 , \3235 , \3236 , \3237 ,
         \3238 , \3239 , \3240 , \3241 , \3242 , \3243 , \3244 , \3245 , \3246 , \3247 ,
         \3248 , \3249 , \3250 , \3251 , \3252 , \3253 , \3254 , \3255 , \3256 , \3257 ,
         \3258 , \3259 , \3260 , \3261 , \3262 , \3263 , \3264 , \3265 , \3266 , \3267 ,
         \3268 , \3269 , \3270 , \3271 , \3272 , \3273 , \3274 , \3275 , \3276 , \3277 ,
         \3278 , \3279 , \3280 , \3281 , \3282 , \3283 , \3284 , \3285 , \3286 , \3287 ,
         \3288 , \3289 , \3290 , \3291 , \3292 , \3293 , \3294 , \3295 , \3296 , \3297 ,
         \3298 , \3299 , \3300 , \3301 , \3302 , \3303 , \3304 , \3305 , \3306_nRb1a , \3307 ,
         \3308 , \3309 , \3310 , \3311 , \3312 , \3313 , \3314 , \3315 , \3316 , \3317 ,
         \3318 , \3319 , \3320 , \3321 , \3322 , \3323 , \3324 , \3325 , \3326 , \3327 ,
         \3328 , \3329 , \3330 , \3331 , \3332 , \3333 , \3334 , \3335 , \3336 , \3337 ,
         \3338 , \3339 , \3340 , \3341 , \3342 , \3343 , \3344 , \3345 , \3346 , \3347 ,
         \3348 , \3349 , \3350 , \3351 , \3352 , \3353 , \3354 , \3355 , \3356 , \3357 ,
         \3358 , \3359 , \3360 , \3361 , \3362 , \3363 , \3364 , \3365 , \3366 , \3367 ,
         \3368 , \3369 , \3370 , \3371 , \3372 , \3373 , \3374 , \3375 , \3376 , \3377 ,
         \3378 , \3379 , \3380 , \3381 , \3382 , \3383 , \3384 , \3385 , \3386 , \3387 ,
         \3388 , \3389 , \3390 , \3391 , \3392 , \3393 , \3394 , \3395 , \3396 , \3397 ,
         \3398 , \3399 , \3400 , \3401 , \3402 , \3403 , \3404 , \3405 , \3406 , \3407 ,
         \3408 , \3409 , \3410 , \3411_nR9e2 , \3412 , \3413 , \3414 , \3415 , \3416 , \3417 ,
         \3418 , \3419 , \3420 , \3421 , \3422 , \3423 , \3424 , \3425 , \3426 , \3427 ,
         \3428 , \3429 , \3430 , \3431 , \3432 , \3433 , \3434 , \3435 , \3436 , \3437 ,
         \3438 , \3439 , \3440 , \3441 , \3442 , \3443 , \3444 , \3445 , \3446 , \3447 ,
         \3448 , \3449 , \3450 , \3451 , \3452 , \3453 , \3454 , \3455 , \3456 , \3457 ,
         \3458 , \3459 , \3460 , \3461 , \3462 , \3463 , \3464 , \3465 , \3466 , \3467 ,
         \3468 , \3469 , \3470 , \3471 , \3472 , \3473 , \3474 , \3475 , \3476 , \3477 ,
         \3478 , \3479 , \3480 , \3481 , \3482 , \3483 , \3484 , \3485 , \3486 , \3487 ,
         \3488 , \3489 , \3490 , \3491 , \3492 , \3493 , \3494 , \3495 , \3496 , \3497 ,
         \3498 , \3499 , \3500 , \3501 , \3502 , \3503 , \3504 , \3505 , \3506 , \3507 ,
         \3508 , \3509 , \3510 , \3511 , \3512 , \3513 , \3514 , \3515 , \3516 , \3517 ,
         \3518 , \3519 , \3520 , \3521 , \3522 , \3523 , \3524 , \3525 , \3526 , \3527 ,
         \3528 , \3529 , \3530 , \3531 , \3532 , \3533 , \3534 , \3535 , \3536 , \3537 ,
         \3538 , \3539 , \3540 , \3541 , \3542 , \3543 , \3544 , \3545 , \3546 , \3547 ,
         \3548 , \3549 , \3550 , \3551 , \3552 , \3553 , \3554 , \3555 , \3556 , \3557 ,
         \3558 , \3559 , \3560 , \3561 , \3562 , \3563 , \3564 , \3565 , \3566 , \3567 ,
         \3568 , \3569 , \3570 , \3571 , \3572 , \3573 , \3574 , \3575 , \3576 , \3577 ,
         \3578 , \3579 , \3580 , \3581 , \3582 , \3583 , \3584 , \3585 , \3586 , \3587 ,
         \3588 , \3589 , \3590 , \3591 , \3592 , \3593 , \3594 , \3595 , \3596 , \3597 ,
         \3598 , \3599 , \3600 , \3601 , \3602 , \3603 , \3604 , \3605 , \3606 , \3607 ,
         \3608 , \3609 , \3610 , \3611 , \3612 , \3613 , \3614 , \3615 , \3616 , \3617 ,
         \3618 , \3619 , \3620 , \3621 , \3622 , \3623 , \3624 , \3625 , \3626 , \3627 ,
         \3628 , \3629 , \3630 , \3631 , \3632 , \3633 , \3634 , \3635 , \3636 , \3637 ,
         \3638 , \3639 , \3640 , \3641 , \3642 , \3643 , \3644 , \3645 , \3646 , \3647 ,
         \3648 , \3649 , \3650 , \3651 , \3652 , \3653 , \3654 , \3655 , \3656 , \3657 ,
         \3658 , \3659 , \3660 , \3661 , \3662 , \3663 , \3664 , \3665 , \3666 , \3667 ,
         \3668 , \3669 , \3670 , \3671 , \3672 , \3673 , \3674 , \3675 , \3676 , \3677 ,
         \3678 , \3679 , \3680 , \3681 , \3682 , \3683 , \3684 , \3685 , \3686 , \3687 ,
         \3688 , \3689 , \3690 , \3691 , \3692 , \3693 , \3694 , \3695 , \3696 , \3697 ,
         \3698 , \3699 , \3700 , \3701 , \3702 , \3703 , \3704 , \3705 , \3706 , \3707 ,
         \3708 , \3709 , \3710 , \3711 , \3712 , \3713 , \3714 , \3715 , \3716 , \3717 ,
         \3718 , \3719 , \3720 , \3721 , \3722 , \3723 , \3724 , \3725 , \3726 , \3727 ,
         \3728 , \3729 , \3730 , \3731 , \3732 , \3733 , \3734 , \3735 , \3736 , \3737 ,
         \3738 , \3739 , \3740 , \3741 , \3742 , \3743 , \3744 , \3745 , \3746 , \3747 ,
         \3748 , \3749 , \3750 , \3751 , \3752 , \3753 , \3754 , \3755 , \3756 , \3757 ,
         \3758 , \3759 , \3760 , \3761 , \3762 , \3763 , \3764 , \3765 , \3766 , \3767 ,
         \3768 , \3769 , \3770 , \3771 , \3772 , \3773 , \3774 , \3775 , \3776 , \3777 ,
         \3778 , \3779 , \3780 , \3781 , \3782 , \3783 , \3784 , \3785 , \3786 , \3787 ,
         \3788 , \3789 , \3790 , \3791 , \3792 , \3793 , \3794 , \3795 , \3796 , \3797 ,
         \3798 , \3799 , \3800 , \3801 , \3802 , \3803 , \3804 , \3805 , \3806 , \3807 ,
         \3808 , \3809 , \3810 , \3811 , \3812 , \3813 , \3814 , \3815 , \3816 , \3817 ,
         \3818 , \3819 , \3820 , \3821 , \3822 , \3823 , \3824 , \3825 , \3826 , \3827 ,
         \3828 , \3829 , \3830 , \3831 , \3832 , \3833 , \3834 , \3835 , \3836 , \3837 ,
         \3838 , \3839 , \3840 , \3841 , \3842 , \3843 , \3844 , \3845 , \3846 , \3847 ,
         \3848 , \3849 , \3850 , \3851 , \3852 , \3853 , \3854 , \3855 , \3856 , \3857 ,
         \3858 , \3859 , \3860 , \3861 , \3862 , \3863 , \3864 , \3865 , \3866 , \3867 ,
         \3868 , \3869 , \3870 , \3871 , \3872 , \3873 , \3874 , \3875 , \3876 , \3877 ,
         \3878 , \3879 , \3880 , \3881 , \3882 , \3883 , \3884 , \3885 , \3886 , \3887 ,
         \3888 , \3889 , \3890 , \3891 , \3892 , \3893 , \3894 , \3895 , \3896 , \3897 ,
         \3898 , \3899 , \3900 , \3901 , \3902 , \3903 , \3904 , \3905 , \3906 , \3907 ,
         \3908 , \3909 , \3910 , \3911 , \3912 , \3913 , \3914 , \3915 , \3916 , \3917 ,
         \3918 , \3919 , \3920 , \3921 , \3922 , \3923 , \3924 , \3925 , \3926 , \3927 ,
         \3928 , \3929 , \3930 , \3931 , \3932 , \3933 , \3934 , \3935 , \3936 , \3937 ,
         \3938 , \3939 , \3940 , \3941 , \3942 , \3943 , \3944 , \3945 , \3946 , \3947 ,
         \3948 , \3949 , \3950 , \3951 , \3952 , \3953 , \3954 , \3955 , \3956 , \3957 ,
         \3958 , \3959 , \3960 , \3961 , \3962 , \3963 , \3964 , \3965 , \3966 , \3967 ,
         \3968 , \3969 , \3970 , \3971 , \3972 , \3973 , \3974 , \3975 , \3976 , \3977 ,
         \3978 , \3979 , \3980 , \3981 , \3982 , \3983 , \3984 , \3985 , \3986 , \3987 ,
         \3988 , \3989 , \3990 , \3991 , \3992 , \3993 , \3994 , \3995 , \3996 , \3997 ,
         \3998 , \3999 , \4000 , \4001 , \4002 , \4003 , \4004 , \4005 , \4006 , \4007 ,
         \4008 , \4009 , \4010 , \4011 , \4012 , \4013 , \4014 , \4015 , \4016 , \4017 ,
         \4018 , \4019 , \4020 , \4021 , \4022 , \4023 , \4024 , \4025 , \4026 , \4027 ,
         \4028 , \4029 , \4030 , \4031 , \4032 , \4033 , \4034 , \4035 , \4036 , \4037 ,
         \4038 , \4039 , \4040 , \4041 , \4042 , \4043 , \4044 , \4045 , \4046 , \4047 ,
         \4048 , \4049 , \4050 , \4051 , \4052 , \4053 , \4054 , \4055 , \4056 , \4057 ,
         \4058 , \4059 , \4060 , \4061 , \4062 , \4063 , \4064 , \4065 , \4066 , \4067 ,
         \4068 , \4069 , \4070 , \4071 , \4072 , \4073 , \4074 , \4075 , \4076 , \4077 ,
         \4078 , \4079 , \4080 , \4081 , \4082 , \4083 , \4084 , \4085 , \4086 , \4087 ,
         \4088 , \4089 , \4090 , \4091 , \4092 , \4093 , \4094 , \4095 , \4096 , \4097 ,
         \4098 , \4099 , \4100 , \4101 , \4102 , \4103 , \4104 , \4105 , \4106 , \4107 ,
         \4108 , \4109 , \4110 , \4111 , \4112 , \4113 , \4114 , \4115 , \4116 , \4117 ,
         \4118 , \4119 , \4120 , \4121 , \4122 , \4123 , \4124 , \4125 , \4126 , \4127 ,
         \4128 , \4129 , \4130 , \4131 , \4132 , \4133 , \4134 , \4135 , \4136 , \4137 ,
         \4138 , \4139 , \4140 , \4141 , \4142 , \4143 , \4144 , \4145 , \4146 , \4147 ,
         \4148 , \4149 , \4150 , \4151 , \4152 , \4153 , \4154 , \4155 , \4156 , \4157 ,
         \4158 , \4159 , \4160 , \4161 , \4162 , \4163 , \4164 , \4165 , \4166 , \4167 ,
         \4168 , \4169 , \4170 , \4171 , \4172 , \4173 , \4174 , \4175 , \4176 , \4177 ,
         \4178 , \4179 , \4180 , \4181 , \4182 , \4183 , \4184 , \4185 , \4186 , \4187 ,
         \4188 , \4189 , \4190 , \4191 , \4192 , \4193 , \4194 , \4195 , \4196 , \4197 ,
         \4198 , \4199 , \4200 , \4201 , \4202 , \4203 , \4204 , \4205 , \4206 , \4207 ,
         \4208 , \4209 , \4210 , \4211 , \4212 , \4213 , \4214 , \4215 , \4216 , \4217 ,
         \4218 , \4219 , \4220 , \4221 , \4222 , \4223 , \4224 , \4225 , \4226 , \4227 ,
         \4228 , \4229 , \4230 , \4231 , \4232 , \4233 , \4234 , \4235 , \4236 , \4237 ,
         \4238 , \4239 , \4240 , \4241 , \4242 , \4243 , \4244 , \4245 , \4246 , \4247 ,
         \4248 , \4249 , \4250 , \4251 , \4252 , \4253 , \4254 , \4255 , \4256 , \4257 ,
         \4258 , \4259 , \4260 , \4261 , \4262 , \4263 , \4264 , \4265 , \4266 , \4267 ,
         \4268 , \4269 , \4270 , \4271 , \4272 , \4273 , \4274 , \4275 , \4276 , \4277 ,
         \4278 , \4279 , \4280 , \4281 , \4282 , \4283 , \4284 , \4285 , \4286 , \4287 ,
         \4288 , \4289 , \4290 , \4291 , \4292 , \4293 , \4294 , \4295 , \4296_nR12e0 , \4297 ,
         \4298 , \4299 , \4300 , \4301 , \4302 , \4303 , \4304 , \4305 , \4306 , \4307 ,
         \4308 , \4309 , \4310 , \4311 , \4312 , \4313 , \4314 , \4315 , \4316 , \4317 ,
         \4318 , \4319 , \4320 , \4321 , \4322 , \4323 , \4324 , \4325 , \4326_nR10fd , \4327 ,
         \4328 , \4329 , \4330 , \4331 , \4332 , \4333 , \4334 , \4335 , \4336 , \4337 ,
         \4338 , \4339 , \4340 , \4341 , \4342 , \4343 , \4344 , \4345 , \4346 , \4347 ,
         \4348 , \4349 , \4350 , \4351 , \4352 , \4353 , \4354 , \4355 , \4356_nR10fb , \4357 ,
         \4358 , \4359 , \4360 , \4361 , \4362 , \4363 , \4364 , \4365 , \4366 , \4367 ,
         \4368 , \4369 , \4370 , \4371 , \4372 , \4373 , \4374 , \4375 , \4376 , \4377 ,
         \4378 , \4379 , \4380 , \4381 , \4382 , \4383 , \4384 , \4385 , \4386_nRf42 , \4387 ,
         \4388 , \4389 , \4390 , \4391 , \4392 , \4393 , \4394 , \4395 , \4396 , \4397 ,
         \4398 , \4399 , \4400 , \4401 , \4402 , \4403 , \4404 , \4405 , \4406 , \4407 ,
         \4408 , \4409 , \4410 , \4411 , \4412 , \4413 , \4414 , \4415 , \4416_nRf40 , \4417 ,
         \4418 , \4419 , \4420 , \4421 , \4422 , \4423 , \4424 , \4425 , \4426 , \4427 ,
         \4428 , \4429 , \4430 , \4431 , \4432 , \4433 , \4434 , \4435 , \4436 , \4437 ,
         \4438 , \4439 , \4440 , \4441 , \4442 , \4443 , \4444 , \4445 , \4446_nRdc1 , \4447 ,
         \4448 , \4449 , \4450 , \4451 , \4452 , \4453 , \4454 , \4455 , \4456 , \4457 ,
         \4458 , \4459 , \4460 , \4461 , \4462 , \4463 , \4464 , \4465 , \4466 , \4467 ,
         \4468 , \4469 , \4470 , \4471 , \4472 , \4473 , \4474 , \4475 , \4476_nRdbf , \4477 ,
         \4478 , \4479 , \4480 , \4481 , \4482 , \4483 , \4484 , \4485 , \4486 , \4487 ,
         \4488 , \4489 , \4490 , \4491 , \4492 , \4493 , \4494 , \4495 , \4496 , \4497 ,
         \4498 , \4499 , \4500 , \4501 , \4502 , \4503 , \4504 , \4505 , \4506_nRc88 , \4507 ,
         \4508 , \4509 , \4510 , \4511 , \4512 , \4513 , \4514 , \4515 , \4516 , \4517 ,
         \4518 , \4519 , \4520 , \4521 , \4522 , \4523 , \4524 , \4525 , \4526 , \4527 ,
         \4528 , \4529 , \4530 , \4531 , \4532 , \4533 , \4534 , \4535 , \4536_nRc86 , \4537 ,
         \4538 , \4539 , \4540 , \4541 , \4542 , \4543 , \4544 , \4545 , \4546 , \4547 ,
         \4548 , \4549 , \4550 , \4551 , \4552 , \4553 , \4554 , \4555 , \4556 , \4557 ,
         \4558 , \4559 , \4560 , \4561 , \4562 , \4563 , \4564 , \4565 , \4566_nRb9a , \4567 ,
         \4568 , \4569 , \4570 , \4571 , \4572 , \4573 , \4574 , \4575 , \4576 , \4577 ,
         \4578 , \4579 , \4580 , \4581 , \4582 , \4583 , \4584 , \4585 , \4586 , \4587 ,
         \4588 , \4589 , \4590 , \4591 , \4592 , \4593 , \4594 , \4595 , \4596_nRb9c , \4597 ,
         \4598 , \4599 , \4600 , \4601 , \4602 , \4603 , \4604 , \4605 , \4606 , \4607 ,
         \4608 , \4609 , \4610 , \4611 , \4612 , \4613 , \4614 , \4615 , \4616 , \4617 ,
         \4618 , \4619 , \4620 , \4621 , \4622 , \4623 , \4624 , \4625 , \4626_nRa38 , \4627 ,
         \4628 , \4629 , \4630 , \4631 , \4632 , \4633 , \4634 , \4635 , \4636 , \4637 ,
         \4638 , \4639 , \4640 , \4641 , \4642 , \4643 , \4644 , \4645 , \4646 , \4647 ,
         \4648 , \4649 , \4650 , \4651 , \4652 , \4653 , \4654 , \4655 , \4656_nRa36 , \4657 ,
         \4658 , \4659 , \4660 , \4661 , \4662 , \4663 , \4664 , \4665 , \4666 , \4667 ,
         \4668 , \4669 , \4670 , \4671 , \4672 , \4673 , \4674 , \4675 , \4676 , \4677 ,
         \4678 , \4679 , \4680 , \4681 , \4682 , \4683 , \4684 , \4685 , \4686 , \4687 ,
         \4688 , \4689 , \4690 , \4691 , \4692 , \4693 , \4694 , \4695 , \4696 , \4697 ,
         \4698 , \4699 , \4700 , \4701 , \4702 , \4703 , \4704 , \4705 , \4706 , \4707 ,
         \4708 , \4709 , \4710 , \4711 , \4712 , \4713 , \4714 , \4715 , \4716 , \4717 ,
         \4718 , \4719 , \4720 , \4721 , \4722 , \4723 , \4724 , \4725 , \4726 , \4727 ,
         \4728 , \4729 , \4730 , \4731 , \4732 , \4733 , \4734 , \4735 , \4736 , \4737 ,
         \4738 , \4739 , \4740 , \4741 , \4742 , \4743 , \4744 , \4745 , \4746 , \4747 ,
         \4748 , \4749 , \4750 , \4751 , \4752 , \4753 , \4754 , \4755 , \4756 , \4757 ,
         \4758 , \4759 , \4760 , \4761 , \4762 , \4763 , \4764 , \4765 , \4766 , \4767 ,
         \4768 , \4769 , \4770 , \4771 , \4772_nR194f , \4773 , \4774 , \4775 , \4776 , \4777 ,
         \4778 , \4779 , \4780 , \4781 , \4782 , \4783 , \4784 , \4785 , \4786 , \4787 ,
         \4788 , \4789 , \4790 , \4791 , \4792 , \4793 , \4794 , \4795 , \4796 , \4797 ,
         \4798 , \4799 , \4800 , \4801 , \4802 , \4803 , \4804 , \4805 , \4806 , \4807 ,
         \4808 , \4809 , \4810 , \4811 , \4812 , \4813 , \4814_nR1a6c , \4815 , \4816 , \4817 ,
         \4818 , \4819 , \4820 , \4821 , \4822 , \4823 , \4824 , \4825 , \4826 , \4827 ,
         \4828 , \4829 , \4830 , \4831 , \4832 , \4833 , \4834 , \4835 , \4836 , \4837 ,
         \4838 , \4839 , \4840 , \4841 , \4842 , \4843 , \4844 , \4845 , \4846 , \4847 ,
         \4848 , \4849 , \4850 , \4851 , \4852 , \4853 , \4854 , \4855 , \4856 , \4857 ,
         \4858 , \4859 , \4860 , \4861 , \4862 , \4863 , \4864 , \4865 , \4866 , \4867 ,
         \4868 , \4869 , \4870_nR1859 , \4871 , \4872 , \4873 , \4874 , \4875 , \4876 , \4877 ,
         \4878 , \4879 , \4880 , \4881 , \4882 , \4883 , \4884 , \4885 , \4886 , \4887 ,
         \4888 , \4889 , \4890 , \4891 , \4892 , \4893 , \4894 , \4895 , \4896 , \4897 ,
         \4898 , \4899 , \4900 , \4901 , \4902 , \4903 , \4904 , \4905 , \4906 , \4907 ,
         \4908 , \4909 , \4910 , \4911 , \4912 , \4913 , \4914 , \4915 , \4916 , \4917 ,
         \4918 , \4919 , \4920 , \4921 , \4922 , \4923 , \4924 , \4925 , \4926 , \4927 ,
         \4928 , \4929 , \4930 , \4931 , \4932 , \4933 , \4934 , \4935 , \4936 , \4937 ,
         \4938 , \4939 , \4940 , \4941 , \4942 , \4943 , \4944 , \4945 , \4946 , \4947 ,
         \4948 , \4949 , \4950 , \4951 , \4952 , \4953 , \4954 , \4955 , \4956 , \4957 ,
         \4958 , \4959 , \4960 , \4961 , \4962 , \4963 , \4964 , \4965 , \4966 , \4967 ,
         \4968_nR171b , \4969 , \4970 , \4971 , \4972 , \4973 , \4974 , \4975 , \4976 , \4977 ,
         \4978 , \4979 , \4980 , \4981 , \4982 , \4983 , \4984 , \4985 , \4986 , \4987 ,
         \4988 , \4989 , \4990 , \4991 , \4992 , \4993 , \4994 , \4995 , \4996 , \4997 ,
         \4998 , \4999 , \5000 , \5001 , \5002 , \5003 , \5004 , \5005 , \5006 , \5007 ,
         \5008 , \5009 , \5010 , \5011 , \5012 , \5013 , \5014 , \5015 , \5016 , \5017 ,
         \5018 , \5019 , \5020 , \5021 , \5022 , \5023 , \5024 , \5025 , \5026 , \5027 ,
         \5028_nR162d , \5029 , \5030 , \5031 , \5032 , \5033 , \5034 , \5035 , \5036 , \5037 ,
         \5038 , \5039 , \5040 , \5041 , \5042 , \5043 , \5044 , \5045 , \5046 , \5047 ,
         \5048 , \5049 , \5050 , \5051 , \5052 , \5053 , \5054 , \5055 , \5056 , \5057 ,
         \5058 , \5059 , \5060 , \5061 , \5062 , \5063_nR150e , \5064 , \5065 , \5066 , \5067 ,
         \5068 , \5069 , \5070 , \5071 , \5072 , \5073 , \5074 , \5075 , \5076 , \5077 ,
         \5078 , \5079 , \5080 , \5081 , \5082 , \5083 , \5084 , \5085 , \5086 , \5087 ,
         \5088 , \5089 , \5090 , \5091 , \5092 , \5093 , \5094 , \5095 , \5096 , \5097 ,
         \5098 , \5099 , \5100 , \5101 , \5102 , \5103 , \5104 , \5105 , \5106 , \5107 ,
         \5108 , \5109 , \5110 , \5111 , \5112 , \5113 , \5114 , \5115 , \5116 , \5117 ,
         \5118 , \5119 , \5120 , \5121 , \5122 , \5123 , \5124 , \5125 , \5126 , \5127 ,
         \5128 , \5129 , \5130 , \5131 , \5132 , \5133 , \5134 , \5135 , \5136 , \5137 ,
         \5138 , \5139 , \5140 , \5141 , \5142 , \5143 , \5144 , \5145 , \5146 , \5147 ,
         \5148 , \5149 , \5150 , \5151 , \5152 , \5153 , \5154 , \5155 , \5156 , \5157 ,
         \5158 , \5159 , \5160 , \5161 , \5162 , \5163 , \5164 , \5165 , \5166 , \5167_nR140b ,
         \5168 , \5169 , \5170 , \5171 , \5172 , \5173 , \5174 , \5175 , \5176 , \5177 ,
         \5178 , \5179 , \5180 , \5181 , \5182 , \5183 , \5184 , \5185 , \5186 , \5187 ,
         \5188 , \5189 , \5190 , \5191 , \5192 , \5193 , \5194 , \5195 , \5196 , \5197 ,
         \5198 , \5199 , \5200 , \5201 , \5202 , \5203 , \5204 , \5205 , \5206 , \5207 ,
         \5208 , \5209 , \5210 , \5211 , \5212 , \5213 , \5214 , \5215 , \5216 , \5217 ,
         \5218 , \5219 , \5220 , \5221 , \5222 , \5223 , \5224 , \5225 , \5226 , \5227 ,
         \5228 , \5229 , \5230 , \5231 , \5232 , \5233 , \5234 , \5235 , \5236 , \5237 ,
         \5238 , \5239 , \5240 , \5241 , \5242 , \5243 , \5244 , \5245 , \5246 , \5247 ,
         \5248 , \5249 , \5250 , \5251 , \5252 , \5253 , \5254 , \5255 , \5256 , \5257 ,
         \5258 , \5259 , \5260 , \5261_nR12fd , \5262 , \5263 , \5264 , \5265 , \5266 , \5267 ,
         \5268 , \5269 , \5270 , \5271 , \5272 , \5273 , \5274 , \5275 , \5276 , \5277 ,
         \5278 , \5279 , \5280 , \5281 , \5282 , \5283 , \5284 , \5285 , \5286 , \5287 ,
         \5288 , \5289 , \5290 , \5291 , \5292 , \5293 , \5294 , \5295 , \5296 , \5297 ,
         \5298 , \5299 , \5300 , \5301 , \5302 , \5303 , \5304 , \5305 , \5306 , \5307 ,
         \5308 , \5309 , \5310 , \5311 , \5312 , \5313 , \5314 , \5315 , \5316 , \5317 ,
         \5318 , \5319 , \5320 , \5321 , \5322 , \5323 , \5324 , \5325 , \5326 , \5327 ,
         \5328 , \5329 , \5330 , \5331 , \5332 , \5333 , \5334 , \5335 , \5336 , \5337 ,
         \5338 , \5339 , \5340 , \5341 , \5342 , \5343 , \5344 , \5345 , \5346 , \5347 ,
         \5348 , \5349 , \5350 , \5351 , \5352 , \5353 , \5354 , \5355 , \5356_nR121c , \5357 ,
         \5358 , \5359 , \5360 , \5361 , \5362 , \5363 , \5364 , \5365 , \5366 , \5367 ,
         \5368 , \5369 , \5370 , \5371 , \5372 , \5373 , \5374 , \5375 , \5376 , \5377 ,
         \5378 , \5379 , \5380 , \5381 , \5382 , \5383 , \5384 , \5385 , \5386 , \5387 ,
         \5388 , \5389 , \5390 , \5391 , \5392 , \5393 , \5394 , \5395 , \5396 , \5397 ,
         \5398 , \5399 , \5400 , \5401 , \5402 , \5403 , \5404 , \5405 , \5406 , \5407 ,
         \5408 , \5409 , \5410 , \5411 , \5412 , \5413 , \5414 , \5415 , \5416 , \5417 ,
         \5418 , \5419 , \5420 , \5421 , \5422 , \5423 , \5424 , \5425 , \5426 , \5427 ,
         \5428 , \5429 , \5430 , \5431 , \5432 , \5433 , \5434 , \5435 , \5436 , \5437 ,
         \5438 , \5439 , \5440 , \5441 , \5442 , \5443 , \5444 , \5445 , \5446 , \5447 ,
         \5448 , \5449 , \5450 , \5451 , \5452 , \5453 , \5454 , \5455 , \5456 , \5457 ,
         \5458 , \5459 , \5460 , \5461 , \5462 , \5463 , \5464 , \5465 , \5466 , \5467 ,
         \5468 , \5469 , \5470 , \5471 , \5472 , \5473 , \5474 , \5475 , \5476 , \5477 ,
         \5478 , \5479 , \5480 , \5481 , \5482 , \5483 , \5484 , \5485 , \5486 , \5487 ,
         \5488 , \5489 , \5490 , \5491 , \5492 , \5493 , \5494 , \5495 , \5496 , \5497 ,
         \5498 , \5499 , \5500 , \5501 , \5502 , \5503 , \5504 , \5505 , \5506 , \5507 ,
         \5508 , \5509 , \5510 , \5511 , \5512 , \5513 , \5514 , \5515 , \5516 , \5517 ,
         \5518 , \5519 , \5520 , \5521 , \5522 , \5523 , \5524 , \5525 , \5526 , \5527 ,
         \5528 , \5529 , \5530 , \5531 , \5532 , \5533 , \5534 , \5535 , \5536 , \5537 ,
         \5538 , \5539 , \5540 , \5541 , \5542 , \5543 , \5544 , \5545 , \5546 , \5547 ,
         \5548 , \5549 , \5550 , \5551 , \5552 , \5553 , \5554 , \5555 , \5556 , \5557 ,
         \5558 , \5559 , \5560 , \5561 , \5562 , \5563 , \5564 , \5565 , \5566 , \5567 ,
         \5568 , \5569 , \5570 , \5571 , \5572 , \5573 , \5574 , \5575 , \5576 , \5577 ,
         \5578 , \5579 , \5580 , \5581 , \5582 , \5583 , \5584 , \5585 , \5586 , \5587 ,
         \5588 , \5589 , \5590 , \5591 , \5592 , \5593 , \5594 , \5595_nR111a , \5596 , \5597 ,
         \5598 , \5599 , \5600 , \5601 , \5602 , \5603 , \5604 , \5605 , \5606 , \5607 ,
         \5608 , \5609 , \5610 , \5611 , \5612 , \5613 , \5614 , \5615 , \5616 , \5617 ,
         \5618 , \5619 , \5620 , \5621 , \5622 , \5623 , \5624 , \5625 , \5626 , \5627 ,
         \5628 , \5629 , \5630 , \5631 , \5632 , \5633 , \5634 , \5635 , \5636 , \5637 ,
         \5638 , \5639 , \5640 , \5641 , \5642 , \5643 , \5644 , \5645 , \5646 , \5647 ,
         \5648 , \5649 , \5650 , \5651 , \5652 , \5653 , \5654 , \5655 , \5656 , \5657 ,
         \5658 , \5659 , \5660 , \5661 , \5662 , \5663 , \5664 , \5665 , \5666 , \5667 ,
         \5668 , \5669 , \5670 , \5671 , \5672 , \5673 , \5674 , \5675 , \5676 , \5677 ,
         \5678 , \5679 , \5680 , \5681 , \5682 , \5683 , \5684 , \5685 , \5686 , \5687 ,
         \5688 , \5689 , \5690 , \5691 , \5692 , \5693 , \5694 , \5695 , \5696 , \5697 ,
         \5698 , \5699 , \5700 , \5701 , \5702 , \5703 , \5704 , \5705 , \5706 , \5707 ,
         \5708 , \5709 , \5710 , \5711 , \5712 , \5713 , \5714 , \5715 , \5716 , \5717 ,
         \5718 , \5719 , \5720 , \5721 , \5722 , \5723 , \5724 , \5725 , \5726 , \5727 ,
         \5728 , \5729 , \5730 , \5731 , \5732 , \5733 , \5734 , \5735 , \5736 , \5737 ,
         \5738 , \5739 , \5740 , \5741 , \5742 , \5743 , \5744 , \5745 , \5746 , \5747_nR1037 ,
         \5748 , \5749 , \5750 , \5751 , \5752 , \5753 , \5754 , \5755 , \5756 , \5757 ,
         \5758 , \5759 , \5760 , \5761 , \5762 , \5763 , \5764 , \5765 , \5766 , \5767 ,
         \5768 , \5769 , \5770 , \5771 , \5772 , \5773 , \5774 , \5775 , \5776 , \5777 ,
         \5778 , \5779 , \5780 , \5781 , \5782 , \5783 , \5784 , \5785 , \5786 , \5787 ,
         \5788 , \5789 , \5790 , \5791 , \5792 , \5793 , \5794 , \5795 , \5796 , \5797 ,
         \5798 , \5799 , \5800 , \5801 , \5802 , \5803 , \5804 , \5805 , \5806 , \5807 ,
         \5808 , \5809 , \5810 , \5811 , \5812 , \5813 , \5814 , \5815 , \5816 , \5817 ,
         \5818 , \5819 , \5820 , \5821 , \5822 , \5823 , \5824_nRf5f , \5825 , \5826 , \5827 ,
         \5828 , \5829 , \5830 , \5831 , \5832 , \5833 , \5834 , \5835 , \5836 , \5837 ,
         \5838 , \5839 , \5840 , \5841 , \5842 , \5843 , \5844 , \5845 , \5846 , \5847 ,
         \5848 , \5849 , \5850 , \5851 , \5852 , \5853 , \5854 , \5855 , \5856 , \5857 ,
         \5858 , \5859 , \5860 , \5861 , \5862 , \5863 , \5864 , \5865 , \5866 , \5867 ,
         \5868 , \5869 , \5870 , \5871 , \5872 , \5873 , \5874 , \5875 , \5876 , \5877 ,
         \5878 , \5879 , \5880 , \5881 , \5882 , \5883 , \5884 , \5885 , \5886 , \5887 ,
         \5888 , \5889 , \5890 , \5891 , \5892 , \5893 , \5894 , \5895 , \5896 , \5897 ,
         \5898 , \5899 , \5900 , \5901 , \5902 , \5903 , \5904 , \5905 , \5906 , \5907 ,
         \5908 , \5909 , \5910 , \5911 , \5912 , \5913 , \5914 , \5915 , \5916 , \5917 ,
         \5918 , \5919 , \5920 , \5921 , \5922 , \5923 , \5924 , \5925 , \5926 , \5927 ,
         \5928 , \5929 , \5930 , \5931 , \5932 , \5933 , \5934 , \5935 , \5936 , \5937 ,
         \5938 , \5939 , \5940 , \5941 , \5942 , \5943 , \5944 , \5945 , \5946 , \5947 ,
         \5948 , \5949 , \5950 , \5951 , \5952 , \5953 , \5954 , \5955 , \5956 , \5957 ,
         \5958 , \5959 , \5960 , \5961 , \5962 , \5963 , \5964 , \5965 , \5966 , \5967 ,
         \5968 , \5969 , \5970 , \5971 , \5972 , \5973 , \5974 , \5975 , \5976 , \5977 ,
         \5978 , \5979 , \5980 , \5981 , \5982 , \5983 , \5984 , \5985 , \5986 , \5987 ,
         \5988 , \5989_nRddd , \5990 , \5991 , \5992 , \5993 , \5994 , \5995 , \5996 , \5997 ,
         \5998 , \5999 , \6000 , \6001 , \6002 , \6003 , \6004 , \6005 , \6006 , \6007 ,
         \6008 , \6009 , \6010 , \6011 , \6012 , \6013 , \6014 , \6015 , \6016 , \6017 ,
         \6018 , \6019 , \6020_nRea9 , \6021 , \6022 , \6023 , \6024 , \6025 , \6026 , \6027 ,
         \6028 , \6029 , \6030 , \6031 , \6032 , \6033 , \6034 , \6035 , \6036 , \6037 ,
         \6038 , \6039 , \6040 , \6041 , \6042 , \6043 , \6044 , \6045 , \6046 , \6047 ,
         \6048 , \6049 , \6050 , \6051 , \6052 , \6053 , \6054 , \6055 , \6056 , \6057 ,
         \6058 , \6059 , \6060 , \6061 , \6062 , \6063 , \6064 , \6065 , \6066 , \6067 ,
         \6068 , \6069 , \6070 , \6071 , \6072 , \6073 , \6074 , \6075 , \6076 , \6077 ,
         \6078 , \6079 , \6080 , \6081 , \6082 , \6083 , \6084 , \6085 , \6086 , \6087 ,
         \6088 , \6089 , \6090 , \6091 , \6092 , \6093 , \6094 , \6095 , \6096 , \6097 ,
         \6098 , \6099 , \6100 , \6101 , \6102 , \6103 , \6104 , \6105 , \6106 , \6107 ,
         \6108 , \6109 , \6110 , \6111 , \6112 , \6113 , \6114 , \6115 , \6116 , \6117 ,
         \6118 , \6119 , \6120 , \6121 , \6122 , \6123 , \6124 , \6125 , \6126 , \6127 ,
         \6128 , \6129 , \6130 , \6131 , \6132 , \6133 , \6134 , \6135 , \6136 , \6137 ,
         \6138 , \6139 , \6140 , \6141 , \6142 , \6143 , \6144 , \6145 , \6146 , \6147 ,
         \6148 , \6149 , \6150 , \6151 , \6152 , \6153 , \6154 , \6155 , \6156 , \6157 ,
         \6158 , \6159 , \6160 , \6161 , \6162 , \6163 , \6164 , \6165 , \6166 , \6167 ,
         \6168 , \6169 , \6170 , \6171 , \6172 , \6173 , \6174 , \6175 , \6176 , \6177 ,
         \6178 , \6179 , \6180 , \6181 , \6182 , \6183 , \6184 , \6185 , \6186 , \6187 ,
         \6188 , \6189 , \6190 , \6191 , \6192 , \6193 , \6194 , \6195 , \6196 , \6197 ,
         \6198 , \6199 , \6200 , \6201 , \6202 , \6203 , \6204 , \6205 , \6206 , \6207 ,
         \6208 , \6209 , \6210 , \6211 , \6212 , \6213 , \6214_nRca5 , \6215 , \6216 , \6217 ,
         \6218 , \6219 , \6220 , \6221 , \6222 , \6223 , \6224 , \6225 , \6226 , \6227 ,
         \6228 , \6229 , \6230 , \6231 , \6232 , \6233 , \6234 , \6235 , \6236 , \6237 ,
         \6238 , \6239 , \6240 , \6241 , \6242 , \6243 , \6244 , \6245_nRd47 , \6246 , \6247 ,
         \6248 , \6249 , \6250 , \6251 , \6252 , \6253 , \6254 , \6255 , \6256 , \6257 ,
         \6258 , \6259 , \6260 , \6261 , \6262 , \6263 , \6264 , \6265 , \6266 , \6267 ,
         \6268 , \6269 , \6270 , \6271 , \6272 , \6273 , \6274 , \6275 , \6276 , \6277 ,
         \6278 , \6279 , \6280 , \6281 , \6282 , \6283 , \6284 , \6285 , \6286 , \6287 ,
         \6288 , \6289 , \6290 , \6291 , \6292 , \6293 , \6294 , \6295 , \6296 , \6297 ,
         \6298 , \6299 , \6300 , \6301 , \6302 , \6303 , \6304 , \6305 , \6306 , \6307 ,
         \6308 , \6309 , \6310 , \6311 , \6312 , \6313 , \6314 , \6315 , \6316 , \6317 ,
         \6318 , \6319 , \6320 , \6321 , \6322 , \6323 , \6324 , \6325 , \6326 , \6327 ,
         \6328 , \6329 , \6330 , \6331 , \6332 , \6333 , \6334 , \6335 , \6336 , \6337 ,
         \6338 , \6339 , \6340 , \6341 , \6342 , \6343 , \6344 , \6345 , \6346 , \6347 ,
         \6348 , \6349 , \6350 , \6351 , \6352 , \6353 , \6354 , \6355 , \6356 , \6357 ,
         \6358 , \6359 , \6360 , \6361 , \6362 , \6363 , \6364 , \6365 , \6366 , \6367 ,
         \6368 , \6369 , \6370 , \6371 , \6372 , \6373 , \6374 , \6375 , \6376 , \6377 ,
         \6378 , \6379 , \6380 , \6381 , \6382 , \6383 , \6384 , \6385 , \6386 , \6387 ,
         \6388 , \6389 , \6390 , \6391 , \6392 , \6393 , \6394 , \6395 , \6396 , \6397 ,
         \6398 , \6399 , \6400 , \6401 , \6402 , \6403 , \6404 , \6405 , \6406 , \6407 ,
         \6408 , \6409 , \6410 , \6411 , \6412 , \6413 , \6414 , \6415 , \6416 , \6417 ,
         \6418 , \6419 , \6420 , \6421 , \6422 , \6423 , \6424 , \6425 , \6426 , \6427 ,
         \6428 , \6429 , \6430 , \6431 , \6432 , \6433 , \6434 , \6435 , \6436 , \6437 ,
         \6438 , \6439 , \6440 , \6441 , \6442 , \6443 , \6444 , \6445 , \6446 , \6447 ,
         \6448 , \6449 , \6450 , \6451 , \6452 , \6453 , \6454 , \6455 , \6456 , \6457 ,
         \6458 , \6459 , \6460 , \6461 , \6462 , \6463_nRc21 , \6464 , \6465 , \6466 , \6467 ,
         \6468 , \6469 , \6470 , \6471 , \6472 , \6473 , \6474 , \6475 , \6476 , \6477 ,
         \6478 , \6479 , \6480 , \6481 , \6482 , \6483 , \6484 , \6485 , \6486 , \6487 ,
         \6488 , \6489 , \6490 , \6491 , \6492 , \6493 , \6494 , \6495 , \6496 , \6497 ,
         \6498 , \6499 , \6500 , \6501 , \6502 , \6503 , \6504 , \6505 , \6506 , \6507 ,
         \6508 , \6509 , \6510 , \6511 , \6512 , \6513 , \6514 , \6515 , \6516 , \6517 ,
         \6518 , \6519 , \6520 , \6521 , \6522 , \6523 , \6524 , \6525 , \6526 , \6527 ,
         \6528 , \6529 , \6530 , \6531 , \6532 , \6533 , \6534 , \6535 , \6536 , \6537 ,
         \6538 , \6539 , \6540 , \6541 , \6542 , \6543 , \6544 , \6545 , \6546 , \6547 ,
         \6548 , \6549 , \6550 , \6551 , \6552 , \6553 , \6554 , \6555 , \6556 , \6557 ,
         \6558 , \6559 , \6560 , \6561 , \6562 , \6563 , \6564 , \6565 , \6566 , \6567 ,
         \6568 , \6569 , \6570 , \6571 , \6572 , \6573_nRb98 , \6574 , \6575 , \6576 , \6577 ,
         \6578 , \6579 , \6580 , \6581 , \6582 , \6583 , \6584 , \6585 , \6586 , \6587 ,
         \6588 , \6589 , \6590 , \6591 , \6592 , \6593 , \6594 , \6595 , \6596 , \6597 ,
         \6598 , \6599 , \6600 , \6601 , \6602 , \6603 , \6604 , \6605 , \6606 , \6607 ,
         \6608 , \6609 , \6610 , \6611 , \6612 , \6613 , \6614 , \6615 , \6616 , \6617 ,
         \6618 , \6619 , \6620 , \6621 , \6622 , \6623 , \6624 , \6625 , \6626 , \6627 ,
         \6628 , \6629 , \6630 , \6631 , \6632 , \6633 , \6634 , \6635 , \6636 , \6637 ,
         \6638 , \6639 , \6640 , \6641 , \6642 , \6643 , \6644 , \6645 , \6646 , \6647 ,
         \6648 , \6649 , \6650 , \6651 , \6652 , \6653 , \6654 , \6655 , \6656 , \6657 ,
         \6658 , \6659 , \6660 , \6661 , \6662 , \6663 , \6664 , \6665 , \6666 , \6667 ,
         \6668 , \6669 , \6670 , \6671 , \6672 , \6673 , \6674 , \6675 , \6676 , \6677 ,
         \6678 , \6679 , \6680 , \6681 , \6682 , \6683 , \6684 , \6685 , \6686 , \6687 ,
         \6688 , \6689 , \6690 , \6691 , \6692 , \6693 , \6694 , \6695 , \6696 , \6697 ,
         \6698 , \6699 , \6700 , \6701 , \6702 , \6703 , \6704 , \6705 , \6706 , \6707 ,
         \6708 , \6709 , \6710 , \6711 , \6712 , \6713 , \6714 , \6715 , \6716 , \6717 ,
         \6718 , \6719 , \6720 , \6721 , \6722 , \6723 , \6724 , \6725 , \6726 , \6727 ,
         \6728 , \6729 , \6730 , \6731 , \6732 , \6733 , \6734 , \6735 , \6736 , \6737 ,
         \6738 , \6739 , \6740 , \6741 , \6742 , \6743 , \6744 , \6745 , \6746 , \6747 ,
         \6748 , \6749_nRb36 , \6750 , \6751 , \6752 , \6753 , \6754 , \6755 , \6756 , \6757 ,
         \6758 , \6759 , \6760 , \6761 , \6762 , \6763 , \6764 , \6765 , \6766 , \6767 ,
         \6768 , \6769 , \6770 , \6771 , \6772 , \6773 , \6774 , \6775 , \6776 , \6777 ,
         \6778 , \6779 , \6780 , \6781 , \6782 , \6783 , \6784 , \6785 , \6786 , \6787 ,
         \6788 , \6789 , \6790 , \6791 , \6792 , \6793 , \6794 , \6795 , \6796 , \6797 ,
         \6798 , \6799 , \6800 , \6801 , \6802 , \6803 , \6804 , \6805 , \6806 , \6807 ,
         \6808 , \6809 , \6810 , \6811 , \6812 , \6813 , \6814 , \6815 , \6816 , \6817 ,
         \6818 , \6819 , \6820 , \6821 , \6822 , \6823 , \6824 , \6825 , \6826 , \6827 ,
         \6828 , \6829 , \6830 , \6831 , \6832 , \6833 , \6834 , \6835 , \6836 , \6837 ,
         \6838 , \6839 , \6840 , \6841 , \6842 , \6843 , \6844 , \6845 , \6846 , \6847_nRa33 ,
         \6848 , \6849 , \6850 , \6851 , \6852 , \6853 , \6854 , \6855 , \6856 , \6857 ,
         \6858 , \6859 , \6860 , \6861 , \6862 , \6863 , \6864 , \6865 , \6866 , \6867 ,
         \6868 , \6869 , \6870 , \6871 , \6872 , \6873 , \6874 , \6875 , \6876 , \6877 ,
         \6878 , \6879 , \6880 , \6881 , \6882 , \6883 , \6884 , \6885 , \6886 , \6887 ,
         \6888 , \6889 , \6890 , \6891 , \6892 , \6893 , \6894 , \6895 , \6896 , \6897 ,
         \6898 , \6899 , \6900 , \6901 , \6902 , \6903 , \6904 , \6905 , \6906 , \6907 ,
         \6908 , \6909 , \6910 , \6911 , \6912 , \6913 , \6914 , \6915 , \6916 , \6917 ,
         \6918 , \6919 , \6920 , \6921 , \6922 , \6923 , \6924 , \6925 , \6926 , \6927 ,
         \6928 , \6929 , \6930 , \6931 , \6932 , \6933 , \6934 , \6935 , \6936 , \6937 ,
         \6938 , \6939 , \6940 , \6941 , \6942 , \6943 , \6944 , \6945 , \6946 , \6947 ,
         \6948 , \6949 , \6950 , \6951 , \6952 , \6953 , \6954 , \6955 , \6956 , \6957 ,
         \6958 , \6959 , \6960 , \6961 , \6962 , \6963 , \6964 , \6965 , \6966 , \6967 ,
         \6968 , \6969 , \6970 , \6971 , \6972 , \6973 , \6974 , \6975 , \6976 , \6977 ,
         \6978 , \6979 , \6980 , \6981 , \6982 , \6983 , \6984 , \6985 , \6986 , \6987 ,
         \6988 , \6989 , \6990 , \6991 , \6992 , \6993 , \6994 , \6995 , \6996 , \6997 ,
         \6998 , \6999 , \7000 , \7001 , \7002 , \7003 , \7004 , \7005 , \7006 , \7007 ,
         \7008 , \7009 , \7010 , \7011 , \7012 , \7013 , \7014 , \7015 , \7016 , \7017 ,
         \7018 , \7019 , \7020 , \7021 , \7022 , \7023 , \7024 , \7025 , \7026 , \7027 ,
         \7028 , \7029 , \7030 , \7031 , \7032 , \7033 , \7034 , \7035 , \7036 , \7037 ,
         \7038 , \7039 , \7040 , \7041 , \7042 , \7043 , \7044 , \7045 , \7046 , \7047 ,
         \7048 , \7049 , \7050 , \7051 , \7052 , \7053 , \7054 , \7055 , \7056 , \7057 ,
         \7058 , \7059 , \7060 , \7061 , \7062 , \7063 , \7064 , \7065 , \7066 , \7067 ,
         \7068 , \7069 , \7070 , \7071 , \7072 , \7073 , \7074 , \7075 , \7076 , \7077 ,
         \7078 , \7079 , \7080 , \7081 , \7082 , \7083 , \7084 , \7085 , \7086 , \7087 ,
         \7088 , \7089 , \7090 , \7091 , \7092 , \7093 , \7094 , \7095 , \7096 , \7097 ,
         \7098 , \7099 , \7100 , \7101 , \7102 , \7103 , \7104 , \7105 , \7106 , \7107 ,
         \7108 , \7109 , \7110 , \7111 , \7112 , \7113 , \7114 , \7115 , \7116 , \7117 ,
         \7118 , \7119 , \7120 , \7121 , \7122 , \7123 , \7124 , \7125 , \7126 , \7127 ,
         \7128 , \7129 , \7130 , \7131 , \7132 , \7133 , \7134 , \7135 , \7136 , \7137 ,
         \7138 , \7139 , \7140 , \7141 , \7142 , \7143 , \7144 , \7145 , \7146 , \7147 ,
         \7148 , \7149 , \7150 , \7151 , \7152 , \7153 , \7154 , \7155 , \7156 , \7157 ,
         \7158 , \7159 , \7160 , \7161 , \7162 , \7163 , \7164 , \7165 , \7166 , \7167 ,
         \7168 , \7169 , \7170 , \7171 , \7172 , \7173 , \7174 , \7175 , \7176 , \7177 ,
         \7178 , \7179 , \7180 , \7181 , \7182 , \7183 , \7184 , \7185 , \7186 , \7187 ,
         \7188 , \7189 , \7190 , \7191 , \7192 , \7193 , \7194 , \7195 , \7196 , \7197 ,
         \7198 , \7199 , \7200 , \7201 , \7202 , \7203 , \7204 , \7205 , \7206 , \7207 ,
         \7208 , \7209 , \7210 , \7211 , \7212 , \7213 , \7214 , \7215 , \7216 , \7217 ,
         \7218 , \7219 , \7220 , \7221 , \7222 , \7223 , \7224 , \7225 , \7226 , \7227 ,
         \7228 , \7229 , \7230 , \7231 , \7232 , \7233 , \7234 , \7235 , \7236 , \7237 ,
         \7238 , \7239 , \7240 , \7241 , \7242 , \7243 , \7244 , \7245 , \7246 , \7247 ,
         \7248 , \7249 , \7250 , \7251 , \7252 , \7253 , \7254 , \7255 , \7256 , \7257 ,
         \7258 , \7259 , \7260 , \7261 , \7262 , \7263 , \7264 , \7265 , \7266 , \7267 ,
         \7268 , \7269 , \7270 , \7271 , \7272 , \7273 , \7274 , \7275 , \7276 , \7277 ,
         \7278 , \7279 , \7280 , \7281 , \7282 , \7283 , \7284 , \7285 , \7286 , \7287 ,
         \7288 , \7289 , \7290 , \7291 , \7292 , \7293 , \7294 , \7295 , \7296 , \7297 ,
         \7298 , \7299 , \7300 , \7301 , \7302 , \7303 , \7304 , \7305 , \7306 , \7307 ,
         \7308 , \7309 , \7310 , \7311 , \7312 , \7313 , \7314 , \7315 , \7316 , \7317 ,
         \7318 , \7319 , \7320 , \7321 , \7322 , \7323 , \7324 , \7325 , \7326 , \7327 ,
         \7328 , \7329 , \7330 , \7331 , \7332 , \7333 , \7334 , \7335 , \7336 , \7337 ,
         \7338 , \7339 , \7340 , \7341 , \7342 , \7343 , \7344 , \7345 , \7346 , \7347 ,
         \7348 , \7349 , \7350 , \7351 , \7352 , \7353 , \7354 , \7355 , \7356 , \7357 ,
         \7358 , \7359 , \7360 , \7361 , \7362 , \7363 , \7364 , \7365 , \7366 , \7367 ,
         \7368 , \7369 , \7370 , \7371 , \7372 , \7373 , \7374 , \7375 , \7376 , \7377 ,
         \7378 , \7379 , \7380 , \7381 , \7382 , \7383 , \7384 , \7385 , \7386 , \7387 ,
         \7388 , \7389 , \7390 , \7391 , \7392 , \7393 , \7394 , \7395 , \7396 , \7397 ,
         \7398 , \7399 , \7400 , \7401 , \7402 , \7403 , \7404 , \7405 , \7406 , \7407 ,
         \7408 , \7409 , \7410 , \7411 , \7412 , \7413 , \7414 , \7415 , \7416 , \7417 ,
         \7418 , \7419 , \7420 , \7421 , \7422 , \7423 , \7424 , \7425 , \7426 , \7427 ,
         \7428 , \7429 , \7430 , \7431 , \7432 , \7433 , \7434 , \7435 , \7436 , \7437 ,
         \7438 , \7439 , \7440 , \7441 , \7442 , \7443 , \7444 , \7445 , \7446 , \7447 ,
         \7448 , \7449 , \7450 , \7451 , \7452 , \7453 , \7454 , \7455 , \7456 , \7457 ,
         \7458 , \7459 , \7460 , \7461 , \7462 , \7463 , \7464 , \7465 , \7466 , \7467 ,
         \7468 , \7469 , \7470 , \7471 , \7472 , \7473 , \7474 , \7475 , \7476 , \7477 ,
         \7478 , \7479 , \7480 , \7481 , \7482 , \7483 , \7484 , \7485 , \7486 , \7487 ,
         \7488 , \7489 , \7490 , \7491 , \7492 , \7493 , \7494 , \7495 , \7496 , \7497 ,
         \7498 , \7499 , \7500 , \7501 , \7502 , \7503 , \7504 , \7505 , \7506 , \7507 ,
         \7508 , \7509 , \7510 , \7511 , \7512 , \7513 , \7514 , \7515 , \7516 , \7517 ,
         \7518 , \7519 , \7520 , \7521 , \7522 , \7523 , \7524 , \7525 , \7526 , \7527 ,
         \7528 , \7529 , \7530 , \7531 , \7532 , \7533 , \7534 , \7535 , \7536 , \7537 ,
         \7538 , \7539 , \7540 , \7541 , \7542 , \7543 , \7544 , \7545 , \7546 , \7547 ,
         \7548 , \7549 , \7550 , \7551 , \7552 , \7553 , \7554 , \7555 , \7556 , \7557 ,
         \7558 , \7559 , \7560 , \7561 , \7562 , \7563 , \7564 , \7565 , \7566 , \7567 ,
         \7568 , \7569 , \7570 , \7571 , \7572 , \7573 , \7574 , \7575 , \7576 , \7577 ,
         \7578 , \7579 , \7580 , \7581 , \7582 , \7583 , \7584 , \7585 , \7586 , \7587 ,
         \7588 , \7589 , \7590 , \7591 , \7592 , \7593 , \7594 , \7595 , \7596 , \7597 ,
         \7598 , \7599 , \7600 , \7601 , \7602 , \7603 , \7604 , \7605 , \7606 , \7607 ,
         \7608 , \7609 , \7610 , \7611 , \7612 , \7613 , \7614 , \7615 , \7616 , \7617 ,
         \7618 , \7619 , \7620 , \7621 , \7622 , \7623 , \7624 , \7625 , \7626 , \7627 ,
         \7628 , \7629 , \7630 , \7631 , \7632 , \7633 , \7634 , \7635 , \7636 , \7637 ,
         \7638 , \7639 , \7640 , \7641 , \7642 , \7643 , \7644 , \7645 , \7646 , \7647 ,
         \7648 , \7649 , \7650 , \7651 , \7652 , \7653 , \7654 , \7655 , \7656 , \7657 ,
         \7658 , \7659 , \7660 , \7661 , \7662 , \7663 , \7664 , \7665 , \7666 , \7667 ,
         \7668 , \7669 , \7670 , \7671 , \7672 , \7673 , \7674 , \7675 , \7676 , \7677 ,
         \7678 , \7679 , \7680 , \7681 , \7682 , \7683 , \7684 , \7685 , \7686 , \7687 ,
         \7688 , \7689 , \7690 , \7691 , \7692 , \7693 , \7694 , \7695 , \7696 , \7697 ,
         \7698 , \7699 , \7700 , \7701 , \7702 , \7703 , \7704 , \7705 , \7706 , \7707 ,
         \7708 , \7709 , \7710 , \7711 , \7712 , \7713 , \7714 , \7715 , \7716 , \7717 ,
         \7718 , \7719 , \7720 , \7721_nR53c , \7722 , \7723 , \7724_nR55b , \7725 , \7726 , \7727 ,
         \7728_nR613 , \7729 , \7730 , \7731 , \7732_nR615 , \7733 , \7734 , \7735 , \7736_nR632 , \7737 ,
         \7738 , \7739_nR634 , \7740 , \7741 , \7742 , \7743 , \7744_nR5f6 , \7745 , \7746 , \7747 ,
         \7748_nR5f4 , \7749 , \7750 , \7751 , \7752 , \7753_nR5d7 , \7754 , \7755 , \7756 , \7757 ,
         \7758 , \7759_nR5d5 , \7760 , \7761 , \7762 , \7763_nR5b8 , \7764 , \7765 , \7766_nR5b6 , \7767 ,
         \7768 , \7769 , \7770 , \7771 , \7772_nR599 , \7773 , \7774 , \7775 , \7776 , \7777 ,
         \7778_nR597 , \7779 , \7780 , \7781 , \7782_nR57a , \7783 , \7784 , \7785_nR578 , \7786 , \7787 ,
         \7788 , \7789 , \7790 , \7791 , \7792 , \7793 , \7794_nR559 , \7795 , \7796 , \7797 ,
         \7798 , \7799 , \7800 , \7801_nR53a , \7802 , \7803 , \7804 , \7805_nR51d , \7806 , \7807 ,
         \7808 , \7809 , \7810 , \7811_nR51b , \7812 , \7813 , \7814 , \7815_nR4fe , \7816 , \7817 ,
         \7818_nR4fc , \7819 , \7820 , \7821 , \7822 , \7823 , \7824_nR4df , \7825 , \7826 , \7827 ,
         \7828 , \7829 , \7830_nR4c2 , \7831 , \7832 , \7833 , \7834_nR4a4 , \7835 , \7836 , \7837_nR486 ,
         \7838 , \7839 , \7840 , \7841 , \7842 , \7843 , \7844 , \7845 , \7846 , \7847 ,
         \7848 , \7849 , \7850 , \7851 , \7852 , \7853 , \7854 , \7855 , \7856 , \7857 ,
         \7858 , \7859 , \7860 , \7861 , \7862 , \7863 , \7864 , \7865_nRaa0 , \7866 , \7867 ,
         \7868_nRaa3 , \7869 , \7870 , \7871 , \7872 , \7873 , \7874 , \7875 , \7876 , \7877 ,
         \7878_nR35b , \7879 , \7880 , \7881 , \7882 , \7883 , \7884 , \7885_nR379 , \7886 , \7887 ,
         \7888_nR397 , \7889 , \7890 , \7891 , \7892 , \7893 , \7894 , \7895 , \7896_nR3b5 , \7897 ,
         \7898 , \7899_nR3d3 , \7900 , \7901 , \7902 , \7903 , \7904 , \7905 , \7906 , \7907_nR3f1 ,
         \7908 , \7909 , \7910_nR40f , \7911 , \7912 , \7913 , \7914 , \7915 , \7916_nR42d , \7917 ,
         \7918 , \7919_nR44b , \7920 , \7921 , \7922 , \7923 , \7924 , \7925 , \7926 , \7927 ,
         \7928 , \7929 , \7930 , \7931 , \7932 , \7933 , \7934 , \7935 , \7936 , \7937 ,
         \7938 , \7939 , \7940 , \7941 , \7942 , \7943 , \7944 , \7945 , \7946 , \7947 ,
         \7948 , \7949 , \7950 , \7951 , \7952 , \7953 , \7954 , \7955 , \7956 , \7957 ,
         \7958 , \7959 , \7960 , \7961_nR33d , \7962 , \7963 , \7964 , \7965 , \7966 , \7967 ,
         \7968 , \7969 , \7970_nR31f , \7971 , \7972 , \7973 , \7974 , \7975 , \7976 , \7977 ,
         \7978 , \7979_nR23b8 , \7980 , \7981 , \7982 , \7983 , \7984 , \7985 , \7986 , \7987 ,
         \7988 , \7989_nR237b , \7990 , \7991 , \7992 , \7993 , \7994 , \7995 , \7996_nR2348 , \7997 ,
         \7998 , \7999 , \8000 , \8001 , \8002 , \8003_nR2309 , \8004 , \8005 , \8006 , \8007 ,
         \8008 , \8009 , \8010 , \8011 , \8012 , \8013 , \8014_nR22a9 , \8015 , \8016 , \8017 ,
         \8018 , \8019 , \8020_nR2238 , \8021 , \8022 , \8023 , \8024 , \8025 , \8026_nR21a2 , \8027 ,
         \8028 , \8029 , \8030 , \8031 , \8032 , \8033 , \8034 , \8035 , \8036 , \8037_nR20fe ,
         \8038 , \8039 , \8040 , \8041 , \8042 , \8043 , \8044 , \8045 , \8046 , \8047 ,
         \8048 , \8049 , \8050 , \8051 , \8052_nR2046 , \8053 , \8054 , \8055 , \8056 , \8057 ,
         \8058 , \8059 , \8060 , \8061_nR1f79 , \8062 , \8063 , \8064 , \8065 , \8066 , \8067 ,
         \8068 , \8069 , \8070 , \8071_nR1eb0 , \8072 , \8073 , \8074 , \8075 , \8076 , \8077 ,
         \8078 , \8079 , \8080 , \8081 , \8082 , \8083 , \8084 , \8085 , \8086 , \8087 ,
         \8088_nR1dda , \8089 , \8090 , \8091 , \8092 , \8093 , \8094 , \8095 , \8096 , \8097 ,
         \8098 , \8099 , \8100 , \8101 , \8102_nR1cfd , \8103 , \8104 , \8105 , \8106 , \8107 ,
         \8108 , \8109 , \8110 , \8111 , \8112 , \8113_nR1c44 , \8114 , \8115 , \8116 , \8117 ,
         \8118 , \8119_nR1b4c , \8120 , \8121 , \8122 , \8123 , \8124 , \8125_nR1a31 , \8126 , \8127 ,
         \8128 , \8129 , \8130 , \8131_nR1915 , \8132 , \8133 , \8134 , \8135 , \8136 , \8137 ,
         \8138 , \8139 , \8140 , \8141_nR181e , \8142 , \8143 , \8144 , \8145 , \8146 , \8147 ,
         \8148 , \8149 , \8150 , \8151 , \8152 , \8153_nR16e0 , \8154 , \8155 , \8156 , \8157 ,
         \8158 , \8159 , \8160 , \8161 , \8162 , \8163 , \8164 , \8165 , \8166 , \8167 ,
         \8168 , \8169_nR15f3 , \8170 , \8171 , \8172 , \8173 , \8174 , \8175_nR14d3 , \8176 , \8177 ,
         \8178 , \8179 , \8180 , \8181_nR13d0 , \8182 , \8183 , \8184 , \8185 , \8186 , \8187_nR12be ,
         \8188 , \8189 , \8190 , \8191 , \8192 , \8193_nR11e2 , \8194 , \8195 , \8196 , \8197 ,
         \8198 , \8199_nR10d7 , \8200 , \8201 , \8202 , \8203 , \8204 , \8205_nRffc , \8206 , \8207 ,
         \8208 , \8209 , \8210 , \8211_nRf1c , \8212 , \8213 , \8214 , \8215 , \8216 , \8217 ,
         \8218 , \8219 , \8220 , \8221 , \8222 , \8223 , \8224 , \8225 , \8226 , \8227 ,
         \8228 , \8229 , \8230 , \8231 , \8232 , \8233 , \8234 , \8235 , \8236 , \8237 ,
         \8238 , \8239 , \8240 , \8241 , \8242 , \8243 , \8244 , \8245 , \8246 , \8247 ,
         \8248 , \8249 , \8250 , \8251 , \8252 , \8253 , \8254 , \8255 , \8256 , \8257 ,
         \8258 , \8259 , \8260 , \8261 , \8262 , \8263 , \8264 , \8265 , \8266 , \8267 ,
         \8268 , \8269 , \8270 , \8271 , \8272 , \8273 , \8274 , \8275 , \8276 , \8277 ,
         \8278 , \8279 , \8280 , \8281 , \8282 , \8283 , \8284 , \8285 , \8286 , \8287 ,
         \8288 , \8289 , \8290 , \8291 , \8292 , \8293 , \8294 , \8295 , \8296 , \8297 ,
         \8298 , \8299 , \8300 , \8301 , \8302 , \8303 , \8304 , \8305 , \8306 , \8307 ,
         \8308 , \8309_nR2ce1 , \8310 , \8311 , \8312 , \8313 , \8314 , \8315 , \8316 , \8317 ,
         \8318 , \8319 , \8320 , \8321 , \8322 , \8323 , \8324 , \8325 , \8326 , \8327 ,
         \8328 , \8329 , \8330 , \8331 , \8332 , \8333 , \8334 , \8335 , \8336 , \8337 ,
         \8338 , \8339 , \8340 , \8341 , \8342 , \8343 , \8344 , \8345_nR2af6 , \8346 , \8347 ,
         \8348 , \8349 , \8350 , \8351 , \8352 , \8353 , \8354 , \8355 , \8356 , \8357 ,
         \8358 , \8359 , \8360 , \8361 , \8362 , \8363 , \8364 , \8365 , \8366 , \8367 ,
         \8368 , \8369 , \8370 , \8371 , \8372 , \8373 , \8374 , \8375 , \8376 , \8377 ,
         \8378 , \8379 , \8380 , \8381_nR2af4 , \8382 , \8383 , \8384 , \8385 , \8386 , \8387 ,
         \8388 , \8389 , \8390 , \8391 , \8392 , \8393 , \8394 , \8395 , \8396 , \8397 ,
         \8398 , \8399 , \8400 , \8401 , \8402 , \8403 , \8404 , \8405 , \8406 , \8407 ,
         \8408 , \8409 , \8410 , \8411 , \8412 , \8413 , \8414 , \8415 , \8416 , \8417_nR293b ,
         \8418 , \8419 , \8420 , \8421 , \8422 , \8423 , \8424 , \8425 , \8426 , \8427 ,
         \8428 , \8429 , \8430 , \8431 , \8432 , \8433 , \8434 , \8435 , \8436 , \8437 ,
         \8438 , \8439 , \8440 , \8441 , \8442 , \8443 , \8444 , \8445 , \8446 , \8447 ,
         \8448 , \8449 , \8450 , \8451 , \8452 , \8453_nR2939 , \8454 , \8455 , \8456 , \8457 ,
         \8458 , \8459 , \8460 , \8461 , \8462 , \8463 , \8464 , \8465 , \8466 , \8467 ,
         \8468 , \8469 , \8470 , \8471 , \8472 , \8473 , \8474 , \8475 , \8476 , \8477 ,
         \8478 , \8479 , \8480 , \8481 , \8482 , \8483 , \8484 , \8485 , \8486 , \8487 ,
         \8488 , \8489_nR27af , \8490 , \8491 , \8492 , \8493 , \8494 , \8495 , \8496 , \8497 ,
         \8498 , \8499 , \8500 , \8501 , \8502 , \8503 , \8504 , \8505 , \8506 , \8507 ,
         \8508 , \8509 , \8510 , \8511 , \8512 , \8513 , \8514 , \8515 , \8516 , \8517 ,
         \8518 , \8519 , \8520 , \8521 , \8522 , \8523 , \8524 , \8525_nR27ad , \8526 , \8527 ,
         \8528 , \8529 , \8530 , \8531 , \8532 , \8533 , \8534 , \8535 , \8536 , \8537 ,
         \8538 , \8539 , \8540 , \8541 , \8542 , \8543 , \8544 , \8545 , \8546 , \8547 ,
         \8548 , \8549 , \8550 , \8551 , \8552 , \8553 , \8554 , \8555 , \8556 , \8557 ,
         \8558 , \8559 , \8560 , \8561_nR2667 , \8562 , \8563 , \8564 , \8565 , \8566 , \8567 ,
         \8568 , \8569 , \8570 , \8571 , \8572 , \8573 , \8574 , \8575 , \8576 , \8577 ,
         \8578 , \8579 , \8580 , \8581 , \8582 , \8583 , \8584 , \8585 , \8586 , \8587 ,
         \8588 , \8589 , \8590 , \8591 , \8592 , \8593 , \8594 , \8595 , \8596 , \8597_nR2665 ,
         \8598 , \8599 , \8600 , \8601 , \8602 , \8603 , \8604 , \8605 , \8606 , \8607 ,
         \8608 , \8609 , \8610 , \8611 , \8612 , \8613 , \8614 , \8615 , \8616 , \8617 ,
         \8618 , \8619 , \8620 , \8621 , \8622 , \8623 , \8624 , \8625 , \8626 , \8627 ,
         \8628 , \8629 , \8630 , \8631 , \8632 , \8633_nR2589 , \8634 , \8635 , \8636 , \8637 ,
         \8638 , \8639 , \8640 , \8641 , \8642 , \8643 , \8644 , \8645 , \8646 , \8647 ,
         \8648 , \8649 , \8650 , \8651 , \8652 , \8653 , \8654 , \8655 , \8656 , \8657 ,
         \8658 , \8659 , \8660 , \8661 , \8662 , \8663 , \8664 , \8665_nR258b , \8666 , \8667 ,
         \8668 , \8669 , \8670 , \8671 , \8672 , \8673 , \8674 , \8675 , \8676 , \8677 ,
         \8678 , \8679 , \8680 , \8681 , \8682 , \8683 , \8684 , \8685 , \8686 , \8687 ,
         \8688 , \8689 , \8690 , \8691 , \8692 , \8693 , \8694 , \8695 , \8696_nR23dd , \8697 ,
         \8698 , \8699 , \8700 , \8701 , \8702 , \8703 , \8704 , \8705 , \8706 , \8707 ,
         \8708 , \8709 , \8710 , \8711 , \8712 , \8713 , \8714 , \8715 , \8716 , \8717 ,
         \8718 , \8719 , \8720 , \8721 , \8722 , \8723 , \8724 , \8725 , \8726 , \8727 ,
         \8728_nR23df , \8729 , \8730 , \8731 , \8732 , \8733 , \8734 , \8735 , \8736 , \8737 ,
         \8738 , \8739 , \8740 , \8741 , \8742 , \8743 , \8744 , \8745 , \8746 , \8747 ,
         \8748 , \8749 , \8750 , \8751 , \8752 , \8753 , \8754 , \8755 , \8756 , \8757 ,
         \8758 , \8759 , \8760 , \8761 , \8762 , \8763 , \8764 , \8765 , \8766 , \8767 ,
         \8768 , \8769 , \8770 , \8771 , \8772 , \8773 , \8774 , \8775 , \8776 , \8777 ,
         \8778 , \8779 , \8780 , \8781 , \8782 , \8783 , \8784 , \8785 , \8786 , \8787 ,
         \8788 , \8789 , \8790 , \8791 , \8792 , \8793 , \8794 , \8795 , \8796 , \8797 ,
         \8798 , \8799 , \8800 , \8801 , \8802 , \8803 , \8804 , \8805 , \8806 , \8807 ,
         \8808 , \8809 , \8810 , \8811 , \8812 , \8813 , \8814 , \8815 , \8816 , \8817 ,
         \8818 , \8819 , \8820 , \8821 , \8822 , \8823 , \8824 , \8825 , \8826 , \8827 ,
         \8828 , \8829 , \8830 , \8831 , \8832 , \8833 , \8834 , \8835 , \8836 , \8837 ,
         \8838 , \8839 , \8840 , \8841 , \8842 , \8843 , \8844 , \8845 , \8846 , \8847 ,
         \8848 , \8849 , \8850 , \8851 , \8852 , \8853 , \8854 , \8855 , \8856 , \8857 ,
         \8858 , \8859 , \8860 , \8861 , \8862 , \8863 , \8864_nR335c , \8865 , \8866 , \8867 ,
         \8868 , \8869 , \8870 , \8871 , \8872 , \8873 , \8874 , \8875 , \8876 , \8877 ,
         \8878 , \8879 , \8880 , \8881 , \8882 , \8883 , \8884 , \8885 , \8886 , \8887 ,
         \8888 , \8889 , \8890 , \8891 , \8892 , \8893 , \8894 , \8895 , \8896 , \8897 ,
         \8898 , \8899 , \8900 , \8901 , \8902 , \8903 , \8904 , \8905 , \8906 , \8907_nR3482 ,
         \8908 , \8909 , \8910 , \8911 , \8912 , \8913 , \8914 , \8915 , \8916 , \8917 ,
         \8918 , \8919 , \8920 , \8921 , \8922 , \8923 , \8924 , \8925 , \8926 , \8927 ,
         \8928 , \8929 , \8930 , \8931 , \8932 , \8933 , \8934 , \8935 , \8936 , \8937 ,
         \8938 , \8939 , \8940 , \8941 , \8942 , \8943 , \8944 , \8945 , \8946 , \8947 ,
         \8948 , \8949 , \8950 , \8951 , \8952 , \8953 , \8954 , \8955 , \8956 , \8957 ,
         \8958 , \8959 , \8960 , \8961 , \8962 , \8963 , \8964 , \8965 , \8966_nR3254 , \8967 ,
         \8968 , \8969 , \8970 , \8971 , \8972 , \8973 , \8974 , \8975 , \8976 , \8977 ,
         \8978 , \8979 , \8980 , \8981 , \8982 , \8983 , \8984 , \8985 , \8986 , \8987 ,
         \8988 , \8989 , \8990 , \8991 , \8992 , \8993 , \8994 , \8995 , \8996 , \8997 ,
         \8998 , \8999 , \9000 , \9001 , \9002 , \9003 , \9004 , \9005 , \9006 , \9007 ,
         \9008 , \9009 , \9010 , \9011 , \9012 , \9013 , \9014 , \9015 , \9016 , \9017 ,
         \9018 , \9019 , \9020 , \9021 , \9022 , \9023 , \9024 , \9025 , \9026 , \9027 ,
         \9028 , \9029 , \9030 , \9031 , \9032 , \9033 , \9034 , \9035 , \9036 , \9037 ,
         \9038 , \9039 , \9040 , \9041 , \9042 , \9043 , \9044 , \9045 , \9046 , \9047 ,
         \9048 , \9049 , \9050 , \9051 , \9052 , \9053 , \9054 , \9055 , \9056 , \9057 ,
         \9058 , \9059 , \9060 , \9061 , \9062 , \9063_nR3133 , \9064 , \9065 , \9066 , \9067 ,
         \9068 , \9069 , \9070 , \9071 , \9072 , \9073 , \9074 , \9075 , \9076 , \9077 ,
         \9078 , \9079 , \9080 , \9081 , \9082 , \9083 , \9084 , \9085 , \9086 , \9087 ,
         \9088 , \9089 , \9090 , \9091 , \9092 , \9093 , \9094 , \9095 , \9096 , \9097 ,
         \9098 , \9099 , \9100 , \9101 , \9102 , \9103 , \9104 , \9105 , \9106 , \9107 ,
         \9108 , \9109 , \9110 , \9111 , \9112 , \9113 , \9114 , \9115 , \9116 , \9117 ,
         \9118 , \9119 , \9120 , \9121 , \9122_nR301c , \9123 , \9124 , \9125 , \9126 , \9127 ,
         \9128 , \9129 , \9130 , \9131 , \9132 , \9133 , \9134 , \9135 , \9136 , \9137 ,
         \9138 , \9139 , \9140 , \9141 , \9142 , \9143 , \9144 , \9145 , \9146 , \9147 ,
         \9148 , \9149 , \9150 , \9151 , \9152 , \9153 , \9154 , \9155 , \9156 , \9157 ,
         \9158 , \9159 , \9160 , \9161 , \9162 , \9163 , \9164 , \9165 , \9166 , \9167 ,
         \9168 , \9169 , \9170 , \9171 , \9172 , \9173 , \9174 , \9175 , \9176 , \9177_nR2f04 ,
         \9178 , \9179 , \9180 , \9181 , \9182 , \9183 , \9184 , \9185 , \9186 , \9187 ,
         \9188 , \9189 , \9190 , \9191 , \9192 , \9193 , \9194 , \9195 , \9196 , \9197 ,
         \9198 , \9199 , \9200 , \9201 , \9202 , \9203 , \9204 , \9205 , \9206 , \9207 ,
         \9208 , \9209 , \9210 , \9211 , \9212 , \9213 , \9214 , \9215 , \9216 , \9217 ,
         \9218 , \9219 , \9220 , \9221 , \9222 , \9223 , \9224 , \9225 , \9226 , \9227 ,
         \9228 , \9229 , \9230 , \9231 , \9232 , \9233 , \9234 , \9235 , \9236 , \9237 ,
         \9238 , \9239 , \9240 , \9241 , \9242 , \9243 , \9244 , \9245 , \9246 , \9247 ,
         \9248 , \9249 , \9250 , \9251 , \9252 , \9253 , \9254 , \9255 , \9256 , \9257 ,
         \9258 , \9259 , \9260 , \9261 , \9262 , \9263 , \9264 , \9265 , \9266 , \9267 ,
         \9268 , \9269 , \9270 , \9271_nR2e0d , \9272 , \9273 , \9274 , \9275 , \9276 , \9277 ,
         \9278 , \9279 , \9280 , \9281 , \9282 , \9283 , \9284 , \9285 , \9286 , \9287 ,
         \9288 , \9289 , \9290 , \9291 , \9292 , \9293 , \9294 , \9295 , \9296 , \9297 ,
         \9298 , \9299 , \9300 , \9301 , \9302 , \9303 , \9304 , \9305 , \9306 , \9307 ,
         \9308 , \9309 , \9310 , \9311 , \9312 , \9313 , \9314 , \9315 , \9316 , \9317 ,
         \9318 , \9319 , \9320 , \9321 , \9322 , \9323 , \9324 , \9325 , \9326 , \9327 ,
         \9328 , \9329 , \9330 , \9331 , \9332 , \9333 , \9334 , \9335 , \9336 , \9337 ,
         \9338 , \9339 , \9340 , \9341 , \9342 , \9343 , \9344 , \9345 , \9346 , \9347 ,
         \9348 , \9349 , \9350 , \9351 , \9352 , \9353 , \9354_nR2cff , \9355 , \9356 , \9357 ,
         \9358 , \9359 , \9360 , \9361 , \9362 , \9363 , \9364 , \9365 , \9366 , \9367 ,
         \9368 , \9369 , \9370 , \9371 , \9372 , \9373 , \9374 , \9375 , \9376 , \9377 ,
         \9378 , \9379 , \9380 , \9381 , \9382 , \9383 , \9384 , \9385 , \9386 , \9387 ,
         \9388 , \9389 , \9390 , \9391 , \9392 , \9393 , \9394 , \9395 , \9396 , \9397 ,
         \9398 , \9399 , \9400 , \9401 , \9402 , \9403 , \9404 , \9405 , \9406 , \9407 ,
         \9408 , \9409 , \9410 , \9411 , \9412 , \9413 , \9414 , \9415 , \9416 , \9417 ,
         \9418 , \9419 , \9420 , \9421 , \9422 , \9423 , \9424 , \9425 , \9426 , \9427 ,
         \9428 , \9429 , \9430 , \9431 , \9432 , \9433 , \9434 , \9435 , \9436 , \9437 ,
         \9438 , \9439 , \9440 , \9441 , \9442 , \9443 , \9444 , \9445 , \9446 , \9447 ,
         \9448 , \9449 , \9450 , \9451 , \9452 , \9453 , \9454 , \9455 , \9456 , \9457 ,
         \9458 , \9459 , \9460 , \9461 , \9462_nR2c1e , \9463 , \9464 , \9465 , \9466 , \9467 ,
         \9468 , \9469 , \9470 , \9471 , \9472 , \9473 , \9474 , \9475 , \9476 , \9477 ,
         \9478 , \9479 , \9480 , \9481 , \9482 , \9483 , \9484 , \9485 , \9486 , \9487 ,
         \9488 , \9489 , \9490 , \9491 , \9492 , \9493 , \9494 , \9495 , \9496 , \9497 ,
         \9498 , \9499 , \9500 , \9501 , \9502 , \9503 , \9504 , \9505 , \9506 , \9507 ,
         \9508 , \9509 , \9510 , \9511 , \9512 , \9513 , \9514 , \9515 , \9516 , \9517 ,
         \9518 , \9519 , \9520 , \9521 , \9522 , \9523 , \9524 , \9525 , \9526 , \9527 ,
         \9528 , \9529 , \9530 , \9531 , \9532 , \9533 , \9534 , \9535 , \9536 , \9537 ,
         \9538 , \9539 , \9540 , \9541 , \9542 , \9543 , \9544 , \9545 , \9546 , \9547 ,
         \9548 , \9549 , \9550 , \9551 , \9552 , \9553 , \9554 , \9555 , \9556 , \9557 ,
         \9558 , \9559 , \9560 , \9561 , \9562 , \9563 , \9564 , \9565 , \9566 , \9567 ,
         \9568 , \9569 , \9570 , \9571 , \9572 , \9573 , \9574 , \9575 , \9576 , \9577 ,
         \9578 , \9579 , \9580 , \9581 , \9582 , \9583 , \9584 , \9585 , \9586 , \9587 ,
         \9588 , \9589 , \9590 , \9591 , \9592 , \9593 , \9594 , \9595 , \9596 , \9597 ,
         \9598 , \9599 , \9600 , \9601 , \9602 , \9603 , \9604 , \9605 , \9606 , \9607 ,
         \9608 , \9609 , \9610 , \9611 , \9612 , \9613 , \9614 , \9615 , \9616 , \9617 ,
         \9618 , \9619 , \9620 , \9621 , \9622 , \9623 , \9624 , \9625 , \9626 , \9627 ,
         \9628 , \9629 , \9630 , \9631 , \9632 , \9633 , \9634 , \9635 , \9636 , \9637 ,
         \9638 , \9639 , \9640 , \9641 , \9642 , \9643 , \9644 , \9645 , \9646 , \9647 ,
         \9648 , \9649 , \9650 , \9651 , \9652 , \9653 , \9654 , \9655 , \9656 , \9657 ,
         \9658 , \9659 , \9660 , \9661 , \9662 , \9663 , \9664 , \9665 , \9666 , \9667 ,
         \9668 , \9669 , \9670 , \9671 , \9672 , \9673 , \9674 , \9675 , \9676 , \9677 ,
         \9678 , \9679 , \9680 , \9681 , \9682 , \9683 , \9684 , \9685 , \9686 , \9687_nR2b14 ,
         \9688 , \9689 , \9690 , \9691 , \9692 , \9693 , \9694 , \9695 , \9696 , \9697 ,
         \9698 , \9699 , \9700 , \9701 , \9702 , \9703 , \9704 , \9705 , \9706 , \9707 ,
         \9708 , \9709 , \9710 , \9711 , \9712 , \9713 , \9714 , \9715 , \9716 , \9717 ,
         \9718 , \9719 , \9720 , \9721 , \9722 , \9723 , \9724 , \9725 , \9726 , \9727 ,
         \9728 , \9729 , \9730 , \9731 , \9732 , \9733 , \9734 , \9735 , \9736 , \9737 ,
         \9738 , \9739 , \9740 , \9741 , \9742 , \9743 , \9744 , \9745 , \9746 , \9747 ,
         \9748 , \9749 , \9750 , \9751 , \9752 , \9753 , \9754 , \9755 , \9756 , \9757 ,
         \9758 , \9759 , \9760 , \9761 , \9762 , \9763 , \9764 , \9765 , \9766 , \9767 ,
         \9768 , \9769 , \9770 , \9771 , \9772 , \9773 , \9774 , \9775 , \9776 , \9777 ,
         \9778 , \9779 , \9780 , \9781 , \9782 , \9783 , \9784 , \9785 , \9786 , \9787 ,
         \9788 , \9789 , \9790 , \9791 , \9792 , \9793 , \9794 , \9795 , \9796 , \9797 ,
         \9798 , \9799 , \9800 , \9801 , \9802 , \9803 , \9804 , \9805 , \9806 , \9807 ,
         \9808 , \9809 , \9810 , \9811 , \9812 , \9813 , \9814 , \9815 , \9816 , \9817 ,
         \9818 , \9819 , \9820 , \9821 , \9822 , \9823 , \9824 , \9825 , \9826 , \9827 ,
         \9828 , \9829 , \9830 , \9831 , \9832 , \9833 , \9834 , \9835 , \9836 , \9837 ,
         \9838 , \9839 , \9840 , \9841 , \9842 , \9843_nR2a34 , \9844 , \9845 , \9846 , \9847 ,
         \9848 , \9849 , \9850 , \9851 , \9852 , \9853 , \9854 , \9855 , \9856 , \9857 ,
         \9858 , \9859 , \9860 , \9861 , \9862 , \9863 , \9864 , \9865 , \9866 , \9867 ,
         \9868 , \9869 , \9870 , \9871 , \9872 , \9873 , \9874 , \9875 , \9876 , \9877 ,
         \9878 , \9879 , \9880 , \9881 , \9882 , \9883 , \9884 , \9885 , \9886 , \9887 ,
         \9888 , \9889 , \9890 , \9891 , \9892 , \9893 , \9894 , \9895 , \9896 , \9897 ,
         \9898 , \9899_nR2959 , \9900 , \9901 , \9902 , \9903 , \9904 , \9905 , \9906 , \9907 ,
         \9908 , \9909 , \9910 , \9911 , \9912 , \9913 , \9914 , \9915 , \9916 , \9917 ,
         \9918 , \9919 , \9920 , \9921 , \9922 , \9923 , \9924 , \9925 , \9926 , \9927 ,
         \9928 , \9929 , \9930 , \9931 , \9932 , \9933 , \9934 , \9935 , \9936 , \9937 ,
         \9938 , \9939 , \9940 , \9941 , \9942 , \9943 , \9944 , \9945 , \9946 , \9947 ,
         \9948 , \9949 , \9950 , \9951 , \9952 , \9953 , \9954 , \9955 , \9956 , \9957 ,
         \9958 , \9959 , \9960 , \9961 , \9962 , \9963 , \9964 , \9965 , \9966 , \9967 ,
         \9968 , \9969 , \9970 , \9971 , \9972 , \9973 , \9974 , \9975 , \9976 , \9977 ,
         \9978 , \9979 , \9980 , \9981 , \9982 , \9983 , \9984 , \9985 , \9986 , \9987 ,
         \9988 , \9989 , \9990 , \9991 , \9992 , \9993 , \9994 , \9995 , \9996 , \9997 ,
         \9998 , \9999 , \10000 , \10001 , \10002 , \10003 , \10004 , \10005 , \10006 , \10007 ,
         \10008 , \10009 , \10010 , \10011 , \10012 , \10013 , \10014 , \10015 , \10016 , \10017 ,
         \10018 , \10019 , \10020 , \10021 , \10022 , \10023 , \10024 , \10025 , \10026 , \10027 ,
         \10028 , \10029 , \10030 , \10031 , \10032 , \10033 , \10034 , \10035 , \10036 , \10037 ,
         \10038 , \10039 , \10040 , \10041 , \10042 , \10043 , \10044 , \10045 , \10046 , \10047 ,
         \10048 , \10049 , \10050 , \10051 , \10052 , \10053 , \10054 , \10055 , \10056 , \10057 ,
         \10058 , \10059 , \10060 , \10061_nR27cd , \10062 , \10063 , \10064 , \10065 , \10066 , \10067 ,
         \10068 , \10069 , \10070 , \10071 , \10072 , \10073 , \10074 , \10075 , \10076 , \10077 ,
         \10078 , \10079 , \10080 , \10081 , \10082 , \10083 , \10084 , \10085 , \10086 , \10087 ,
         \10088 , \10089 , \10090 , \10091 , \10092 , \10093 , \10094_nR289e , \10095 , \10096 , \10097 ,
         \10098 , \10099 , \10100 , \10101 , \10102 , \10103 , \10104 , \10105 , \10106 , \10107 ,
         \10108 , \10109 , \10110 , \10111 , \10112 , \10113 , \10114 , \10115 , \10116 , \10117 ,
         \10118 , \10119 , \10120 , \10121 , \10122 , \10123 , \10124 , \10125 , \10126 , \10127 ,
         \10128 , \10129 , \10130 , \10131 , \10132 , \10133 , \10134 , \10135 , \10136 , \10137 ,
         \10138 , \10139 , \10140 , \10141 , \10142 , \10143 , \10144 , \10145 , \10146 , \10147 ,
         \10148 , \10149 , \10150 , \10151 , \10152 , \10153 , \10154 , \10155 , \10156 , \10157 ,
         \10158 , \10159 , \10160 , \10161 , \10162 , \10163 , \10164 , \10165 , \10166 , \10167 ,
         \10168 , \10169 , \10170 , \10171 , \10172 , \10173 , \10174 , \10175 , \10176 , \10177 ,
         \10178 , \10179 , \10180 , \10181 , \10182 , \10183 , \10184 , \10185 , \10186 , \10187 ,
         \10188 , \10189 , \10190 , \10191 , \10192 , \10193 , \10194 , \10195 , \10196 , \10197 ,
         \10198 , \10199 , \10200 , \10201 , \10202 , \10203 , \10204 , \10205 , \10206 , \10207 ,
         \10208 , \10209 , \10210 , \10211 , \10212 , \10213 , \10214 , \10215 , \10216 , \10217 ,
         \10218 , \10219 , \10220 , \10221 , \10222 , \10223 , \10224 , \10225 , \10226 , \10227 ,
         \10228 , \10229 , \10230 , \10231 , \10232 , \10233 , \10234 , \10235 , \10236 , \10237 ,
         \10238 , \10239 , \10240 , \10241 , \10242 , \10243 , \10244 , \10245 , \10246 , \10247 ,
         \10248 , \10249 , \10250 , \10251 , \10252 , \10253 , \10254 , \10255 , \10256 , \10257 ,
         \10258 , \10259 , \10260 , \10261 , \10262 , \10263 , \10264 , \10265 , \10266 , \10267 ,
         \10268 , \10269 , \10270 , \10271 , \10272 , \10273 , \10274 , \10275 , \10276 , \10277 ,
         \10278 , \10279 , \10280 , \10281 , \10282 , \10283 , \10284 , \10285 , \10286 , \10287 ,
         \10288 , \10289 , \10290 , \10291 , \10292 , \10293 , \10294 , \10295 , \10296 , \10297 ,
         \10298 , \10299 , \10300 , \10301 , \10302 , \10303 , \10304 , \10305 , \10306 , \10307 ,
         \10308 , \10309 , \10310 , \10311 , \10312 , \10313 , \10314_nR2685 , \10315 , \10316 , \10317 ,
         \10318 , \10319 , \10320 , \10321 , \10322 , \10323 , \10324 , \10325 , \10326 , \10327 ,
         \10328 , \10329 , \10330 , \10331 , \10332 , \10333 , \10334 , \10335 , \10336 , \10337 ,
         \10338 , \10339 , \10340 , \10341 , \10342 , \10343 , \10344 , \10345 , \10346 , \10347_nR272f ,
         \10348 , \10349 , \10350 , \10351 , \10352 , \10353 , \10354 , \10355 , \10356 , \10357 ,
         \10358 , \10359 , \10360 , \10361 , \10362 , \10363 , \10364 , \10365 , \10366 , \10367 ,
         \10368 , \10369 , \10370 , \10371 , \10372 , \10373 , \10374 , \10375 , \10376 , \10377 ,
         \10378 , \10379 , \10380 , \10381 , \10382 , \10383 , \10384 , \10385 , \10386 , \10387 ,
         \10388 , \10389 , \10390 , \10391 , \10392 , \10393 , \10394 , \10395 , \10396 , \10397 ,
         \10398 , \10399 , \10400 , \10401 , \10402 , \10403 , \10404 , \10405 , \10406 , \10407 ,
         \10408 , \10409 , \10410 , \10411 , \10412 , \10413 , \10414 , \10415 , \10416 , \10417 ,
         \10418 , \10419 , \10420 , \10421 , \10422 , \10423 , \10424 , \10425 , \10426 , \10427 ,
         \10428 , \10429 , \10430 , \10431 , \10432 , \10433 , \10434 , \10435 , \10436 , \10437 ,
         \10438 , \10439 , \10440 , \10441 , \10442 , \10443 , \10444 , \10445 , \10446 , \10447 ,
         \10448 , \10449 , \10450 , \10451 , \10452 , \10453 , \10454 , \10455 , \10456 , \10457 ,
         \10458 , \10459 , \10460 , \10461 , \10462 , \10463 , \10464 , \10465 , \10466 , \10467 ,
         \10468 , \10469 , \10470 , \10471 , \10472 , \10473 , \10474 , \10475 , \10476 , \10477 ,
         \10478 , \10479 , \10480 , \10481 , \10482 , \10483 , \10484 , \10485 , \10486 , \10487 ,
         \10488 , \10489 , \10490 , \10491 , \10492 , \10493 , \10494 , \10495 , \10496 , \10497 ,
         \10498 , \10499 , \10500 , \10501 , \10502 , \10503 , \10504 , \10505 , \10506 , \10507 ,
         \10508 , \10509 , \10510 , \10511 , \10512 , \10513 , \10514 , \10515 , \10516 , \10517 ,
         \10518 , \10519 , \10520 , \10521 , \10522 , \10523 , \10524 , \10525 , \10526 , \10527 ,
         \10528 , \10529 , \10530 , \10531 , \10532 , \10533 , \10534 , \10535 , \10536 , \10537 ,
         \10538 , \10539 , \10540 , \10541 , \10542 , \10543 , \10544 , \10545 , \10546 , \10547 ,
         \10548 , \10549 , \10550 , \10551 , \10552 , \10553 , \10554 , \10555 , \10556 , \10557 ,
         \10558 , \10559 , \10560 , \10561 , \10562 , \10563 , \10564 , \10565 , \10566 , \10567 ,
         \10568_nR260a , \10569 , \10570 , \10571 , \10572 , \10573 , \10574 , \10575 , \10576 , \10577 ,
         \10578 , \10579 , \10580 , \10581 , \10582 , \10583 , \10584 , \10585 , \10586 , \10587 ,
         \10588 , \10589 , \10590 , \10591 , \10592 , \10593 , \10594 , \10595 , \10596 , \10597 ,
         \10598 , \10599 , \10600 , \10601 , \10602 , \10603 , \10604 , \10605 , \10606 , \10607 ,
         \10608 , \10609 , \10610 , \10611 , \10612 , \10613 , \10614 , \10615 , \10616 , \10617 ,
         \10618 , \10619 , \10620 , \10621 , \10622 , \10623 , \10624 , \10625 , \10626 , \10627 ,
         \10628 , \10629 , \10630 , \10631 , \10632 , \10633 , \10634 , \10635 , \10636 , \10637 ,
         \10638 , \10639 , \10640 , \10641 , \10642 , \10643 , \10644 , \10645 , \10646 , \10647 ,
         \10648 , \10649 , \10650 , \10651 , \10652 , \10653 , \10654 , \10655 , \10656 , \10657 ,
         \10658 , \10659 , \10660 , \10661 , \10662 , \10663 , \10664 , \10665 , \10666 , \10667 ,
         \10668 , \10669 , \10670 , \10671 , \10672 , \10673 , \10674 , \10675 , \10676 , \10677 ,
         \10678 , \10679 , \10680 , \10681 , \10682 , \10683 , \10684 , \10685 , \10686_nR2587 , \10687 ,
         \10688 , \10689 , \10690 , \10691 , \10692 , \10693 , \10694 , \10695 , \10696 , \10697 ,
         \10698 , \10699 , \10700 , \10701 , \10702 , \10703 , \10704 , \10705 , \10706 , \10707 ,
         \10708 , \10709 , \10710 , \10711 , \10712 , \10713 , \10714 , \10715 , \10716 , \10717 ,
         \10718 , \10719 , \10720 , \10721 , \10722 , \10723 , \10724 , \10725 , \10726 , \10727 ,
         \10728 , \10729 , \10730 , \10731 , \10732 , \10733 , \10734 , \10735 , \10736 , \10737 ,
         \10738 , \10739 , \10740 , \10741 , \10742 , \10743 , \10744 , \10745 , \10746 , \10747 ,
         \10748 , \10749 , \10750 , \10751 , \10752 , \10753 , \10754 , \10755 , \10756 , \10757 ,
         \10758 , \10759 , \10760 , \10761 , \10762 , \10763 , \10764 , \10765 , \10766 , \10767 ,
         \10768 , \10769 , \10770 , \10771 , \10772 , \10773 , \10774 , \10775 , \10776 , \10777 ,
         \10778 , \10779 , \10780 , \10781 , \10782 , \10783 , \10784 , \10785 , \10786 , \10787 ,
         \10788 , \10789 , \10790 , \10791 , \10792 , \10793 , \10794 , \10795 , \10796 , \10797 ,
         \10798 , \10799 , \10800 , \10801 , \10802 , \10803 , \10804 , \10805 , \10806 , \10807 ,
         \10808 , \10809 , \10810 , \10811 , \10812 , \10813 , \10814 , \10815 , \10816 , \10817 ,
         \10818 , \10819 , \10820 , \10821 , \10822 , \10823 , \10824 , \10825 , \10826 , \10827 ,
         \10828 , \10829 , \10830 , \10831 , \10832 , \10833 , \10834 , \10835 , \10836 , \10837 ,
         \10838 , \10839 , \10840 , \10841 , \10842 , \10843 , \10844 , \10845 , \10846 , \10847 ,
         \10848 , \10849 , \10850 , \10851 , \10852 , \10853 , \10854 , \10855 , \10856 , \10857 ,
         \10858 , \10859 , \10860_nR251b , \10861 , \10862 , \10863 , \10864 , \10865 , \10866 , \10867 ,
         \10868 , \10869 , \10870 , \10871 , \10872 , \10873 , \10874 , \10875 , \10876 , \10877 ,
         \10878 , \10879 , \10880 , \10881 , \10882 , \10883 , \10884 , \10885 , \10886 , \10887 ,
         \10888 , \10889 , \10890 , \10891 , \10892 , \10893 , \10894 , \10895 , \10896 , \10897 ,
         \10898 , \10899 , \10900 , \10901 , \10902 , \10903 , \10904 , \10905 , \10906 , \10907 ,
         \10908 , \10909 , \10910 , \10911 , \10912 , \10913 , \10914 , \10915 , \10916 , \10917 ,
         \10918 , \10919 , \10920 , \10921 , \10922 , \10923 , \10924 , \10925 , \10926_nR23da , \10927 ,
         \10928 , \10929 , \10930 , \10931 , \10932 , \10933 , \10934 , \10935 , \10936 , \10937 ,
         \10938 , \10939 , \10940 , \10941 , \10942 , \10943 , \10944 , \10945 , \10946 , \10947 ,
         \10948 , \10949 , \10950 , \10951 , \10952 , \10953 , \10954 , \10955 , \10956 , \10957 ,
         \10958 , \10959 , \10960 , \10961 , \10962 , \10963 , \10964 , \10965 , \10966 , \10967 ,
         \10968 , \10969 , \10970 , \10971 , \10972 , \10973 , \10974 , \10975 , \10976 , \10977 ,
         \10978 , \10979 , \10980 , \10981 , \10982 , \10983 , \10984 , \10985 , \10986 , \10987 ,
         \10988 , \10989 , \10990 , \10991 , \10992 , \10993 , \10994 , \10995 , \10996 , \10997 ,
         \10998 , \10999 , \11000 , \11001 , \11002 , \11003 , \11004 , \11005 , \11006 , \11007 ,
         \11008 , \11009 , \11010 , \11011 , \11012 , \11013 , \11014 , \11015 , \11016 , \11017 ,
         \11018 , \11019 , \11020 , \11021 , \11022 , \11023 , \11024 , \11025 , \11026 , \11027 ,
         \11028 , \11029 , \11030 , \11031 , \11032 , \11033 , \11034 , \11035 , \11036 , \11037 ,
         \11038 , \11039 , \11040 , \11041 , \11042 , \11043 , \11044 , \11045 , \11046 , \11047 ,
         \11048 , \11049 , \11050 , \11051 , \11052 , \11053 , \11054 , \11055 , \11056 , \11057 ,
         \11058 , \11059 , \11060 , \11061 , \11062 , \11063 , \11064 , \11065 , \11066 , \11067 ,
         \11068 , \11069 , \11070 , \11071 , \11072 , \11073 , \11074 , \11075 , \11076 , \11077 ,
         \11078 , \11079 , \11080 , \11081 , \11082 , \11083 , \11084 , \11085 , \11086 , \11087 ,
         \11088 , \11089 , \11090 , \11091 , \11092 , \11093 , \11094 , \11095 , \11096 , \11097 ,
         \11098 , \11099 , \11100 , \11101 , \11102 , \11103 , \11104 , \11105 , \11106 , \11107 ,
         \11108 , \11109 , \11110 , \11111 , \11112 , \11113 , \11114 , \11115 , \11116 , \11117 ,
         \11118 , \11119 , \11120 , \11121 , \11122 , \11123 , \11124 , \11125 , \11126 , \11127 ,
         \11128 , \11129 , \11130 , \11131 , \11132 , \11133 , \11134 , \11135 , \11136 , \11137 ,
         \11138 , \11139 , \11140 , \11141 , \11142 , \11143 , \11144 , \11145 , \11146 , \11147 ,
         \11148 , \11149 , \11150 , \11151 , \11152 , \11153 , \11154 , \11155 , \11156 , \11157 ,
         \11158 , \11159 , \11160 , \11161 , \11162 , \11163 , \11164 , \11165 , \11166 , \11167 ,
         \11168 , \11169 , \11170 , \11171 , \11172 , \11173 , \11174 , \11175 , \11176 , \11177 ,
         \11178 , \11179 , \11180 , \11181 , \11182 , \11183 , \11184 , \11185 , \11186 , \11187 ,
         \11188 , \11189 , \11190 , \11191 , \11192 , \11193 , \11194 , \11195 , \11196 , \11197 ,
         \11198 , \11199 , \11200 , \11201 , \11202 , \11203 , \11204 , \11205 , \11206 , \11207 ,
         \11208 , \11209 , \11210 , \11211 , \11212 , \11213 , \11214 , \11215 , \11216 , \11217 ,
         \11218 , \11219 , \11220 , \11221 , \11222 , \11223 , \11224 , \11225 , \11226 , \11227 ,
         \11228 , \11229 , \11230 , \11231 , \11232 , \11233 , \11234 , \11235 , \11236 , \11237 ,
         \11238 , \11239 , \11240 , \11241 , \11242 , \11243 , \11244 , \11245 , \11246 , \11247 ,
         \11248 , \11249 , \11250 , \11251 , \11252 , \11253 , \11254 , \11255 , \11256 , \11257 ,
         \11258 , \11259 , \11260 , \11261 , \11262 , \11263 , \11264 , \11265 , \11266 , \11267 ,
         \11268 , \11269 , \11270 , \11271 , \11272 , \11273 , \11274 , \11275 , \11276 , \11277 ,
         \11278 , \11279 , \11280 , \11281 , \11282 , \11283 , \11284 , \11285 , \11286 , \11287 ,
         \11288 , \11289 , \11290 , \11291 , \11292 , \11293 , \11294 , \11295 , \11296 , \11297 ,
         \11298 , \11299 , \11300 , \11301 , \11302 , \11303 , \11304 , \11305 , \11306 , \11307 ,
         \11308 , \11309 , \11310 , \11311 , \11312 , \11313 , \11314 , \11315 , \11316 , \11317 ,
         \11318 , \11319 , \11320 , \11321 , \11322 , \11323 , \11324 , \11325 , \11326 , \11327 ,
         \11328 , \11329 , \11330 , \11331 , \11332 , \11333 , \11334 , \11335 , \11336 , \11337 ,
         \11338 , \11339 , \11340 , \11341 , \11342 , \11343 , \11344 , \11345 , \11346 , \11347 ,
         \11348 , \11349 , \11350 , \11351 , \11352 , \11353 , \11354 , \11355 , \11356 , \11357 ,
         \11358 , \11359 , \11360 , \11361 , \11362 , \11363 , \11364 , \11365 , \11366 , \11367 ,
         \11368 , \11369 , \11370 , \11371 , \11372 , \11373 , \11374 , \11375 , \11376 , \11377 ,
         \11378 , \11379 , \11380 , \11381 , \11382 , \11383 , \11384 , \11385 , \11386 , \11387 ,
         \11388 , \11389 , \11390 , \11391 , \11392 , \11393 , \11394 , \11395 , \11396 , \11397 ,
         \11398 , \11399 , \11400 , \11401 , \11402 , \11403 , \11404 , \11405 , \11406 , \11407 ,
         \11408 , \11409 , \11410 , \11411 , \11412 , \11413 , \11414 , \11415 , \11416 , \11417 ,
         \11418 , \11419 , \11420 , \11421 , \11422 , \11423 , \11424 , \11425 , \11426 , \11427 ,
         \11428 , \11429 , \11430 , \11431 , \11432 , \11433 , \11434 , \11435 , \11436 , \11437 ,
         \11438 , \11439 , \11440 , \11441 , \11442 , \11443 , \11444 , \11445 , \11446 , \11447 ,
         \11448 , \11449 , \11450 , \11451 , \11452 , \11453 , \11454 , \11455 , \11456 , \11457 ,
         \11458 , \11459 , \11460 , \11461 , \11462 , \11463 , \11464 , \11465 , \11466 , \11467 ,
         \11468 , \11469 , \11470 , \11471 , \11472 , \11473 , \11474 , \11475 , \11476 , \11477 ,
         \11478 , \11479 , \11480 , \11481 , \11482 , \11483 , \11484 , \11485 , \11486 , \11487 ,
         \11488 , \11489 , \11490 , \11491 , \11492 , \11493 , \11494 , \11495 , \11496 , \11497 ,
         \11498 , \11499 , \11500 , \11501 , \11502 , \11503 , \11504 , \11505 , \11506 , \11507 ,
         \11508 , \11509 , \11510 , \11511 , \11512 , \11513 , \11514 , \11515 , \11516 , \11517 ,
         \11518 , \11519 , \11520 , \11521 , \11522 , \11523 , \11524 , \11525 , \11526 , \11527 ,
         \11528 , \11529 , \11530 , \11531 , \11532 , \11533 , \11534 , \11535 , \11536 , \11537 ,
         \11538 , \11539 , \11540 , \11541 , \11542 , \11543 , \11544 , \11545 , \11546 , \11547 ,
         \11548 , \11549 , \11550 , \11551 , \11552 , \11553 , \11554 , \11555 , \11556 , \11557 ,
         \11558 , \11559 , \11560 , \11561 , \11562 , \11563 , \11564 , \11565 , \11566 , \11567 ,
         \11568 , \11569 , \11570 , \11571 , \11572 , \11573 , \11574 , \11575 , \11576 , \11577 ,
         \11578 , \11579 , \11580 , \11581 , \11582 , \11583 , \11584 , \11585 , \11586 , \11587 ,
         \11588 , \11589 , \11590 , \11591 , \11592 , \11593 , \11594 , \11595 , \11596 , \11597 ,
         \11598 , \11599 , \11600 , \11601 , \11602 , \11603 , \11604 , \11605 , \11606 , \11607 ,
         \11608 , \11609 , \11610 , \11611 , \11612 , \11613 , \11614 , \11615 , \11616 , \11617 ,
         \11618 , \11619 , \11620 , \11621 , \11622 , \11623 , \11624 , \11625 , \11626 , \11627 ,
         \11628 , \11629 , \11630 , \11631 , \11632 , \11633 , \11634 , \11635 , \11636 , \11637 ,
         \11638 , \11639 , \11640 , \11641 , \11642 , \11643 , \11644 , \11645 , \11646 , \11647 ,
         \11648 , \11649 , \11650 , \11651 , \11652 , \11653 , \11654 , \11655 , \11656 , \11657 ,
         \11658 , \11659 , \11660 , \11661 , \11662 , \11663 , \11664 , \11665 , \11666 , \11667 ,
         \11668 , \11669 , \11670 , \11671 , \11672 , \11673 , \11674 , \11675 , \11676 , \11677 ,
         \11678 , \11679 , \11680 , \11681 , \11682 , \11683 , \11684 , \11685 , \11686 , \11687 ,
         \11688 , \11689 , \11690 , \11691 , \11692 , \11693 , \11694 , \11695 , \11696 , \11697 ,
         \11698 , \11699 , \11700 , \11701 , \11702 , \11703 , \11704 , \11705 , \11706 , \11707 ,
         \11708 , \11709 , \11710 , \11711 , \11712 , \11713 , \11714 , \11715 , \11716 , \11717 ,
         \11718 , \11719 , \11720 , \11721 , \11722 , \11723 , \11724 , \11725 , \11726 , \11727 ,
         \11728 , \11729 , \11730 , \11731 , \11732 , \11733 , \11734 , \11735 , \11736 , \11737 ,
         \11738 , \11739 , \11740 , \11741 , \11742 , \11743 , \11744 , \11745 , \11746 , \11747 ,
         \11748 , \11749 , \11750 , \11751 , \11752 , \11753 , \11754 , \11755 , \11756 , \11757 ,
         \11758 , \11759 , \11760 , \11761 , \11762 , \11763 , \11764 , \11765 , \11766 , \11767 ,
         \11768 , \11769 , \11770 , \11771 , \11772 , \11773 , \11774 , \11775 , \11776 , \11777 ,
         \11778 , \11779 , \11780 , \11781 , \11782 , \11783 , \11784 , \11785 , \11786 , \11787 ,
         \11788 , \11789 , \11790 , \11791 , \11792 , \11793 , \11794 , \11795 , \11796 , \11797 ,
         \11798 , \11799 , \11800 , \11801 , \11802 , \11803 , \11804 , \11805 , \11806 , \11807 ,
         \11808 , \11809 , \11810 , \11811 , \11812 , \11813 , \11814 , \11815 , \11816 , \11817 ,
         \11818 , \11819 , \11820 , \11821 , \11822 , \11823 , \11824 , \11825 , \11826 , \11827 ,
         \11828 , \11829 , \11830 , \11831 , \11832 , \11833 , \11834 , \11835 , \11836 , \11837 ,
         \11838 , \11839 , \11840 , \11841 , \11842 , \11843 , \11844 , \11845 , \11846 , \11847 ,
         \11848 , \11849 , \11850 , \11851 , \11852 , \11853 , \11854 , \11855 , \11856 , \11857 ,
         \11858 , \11859 , \11860 , \11861 , \11862 , \11863 , \11864 , \11865 , \11866 , \11867 ,
         \11868 , \11869 , \11870 , \11871 , \11872 , \11873 , \11874 , \11875 , \11876 , \11877 ,
         \11878 , \11879 , \11880 , \11881 , \11882 , \11883 , \11884 , \11885 , \11886 , \11887 ,
         \11888 , \11889 , \11890_nR2d01 , \11891 , \11892 , \11893 , \11894 , \11895 , \11896 , \11897 ,
         \11898 , \11899 , \11900 , \11901 , \11902 , \11903 , \11904 , \11905 , \11906 , \11907 ,
         \11908 , \11909 , \11910 , \11911 , \11912 , \11913 , \11914 , \11915 , \11916 , \11917 ,
         \11918 , \11919 , \11920_nR2b18 , \11921 , \11922 , \11923 , \11924 , \11925 , \11926 , \11927 ,
         \11928 , \11929 , \11930 , \11931 , \11932 , \11933 , \11934 , \11935 , \11936 , \11937 ,
         \11938 , \11939 , \11940 , \11941 , \11942 , \11943 , \11944 , \11945 , \11946 , \11947 ,
         \11948 , \11949 , \11950_nR2b16 , \11951 , \11952 , \11953 , \11954 , \11955 , \11956 , \11957 ,
         \11958 , \11959 , \11960 , \11961 , \11962 , \11963 , \11964 , \11965 , \11966 , \11967 ,
         \11968 , \11969 , \11970 , \11971 , \11972 , \11973 , \11974 , \11975 , \11976 , \11977 ,
         \11978 , \11979 , \11980_nR295d , \11981 , \11982 , \11983 , \11984 , \11985 , \11986 , \11987 ,
         \11988 , \11989 , \11990 , \11991 , \11992 , \11993 , \11994 , \11995 , \11996 , \11997 ,
         \11998 , \11999 , \12000 , \12001 , \12002 , \12003 , \12004 , \12005 , \12006 , \12007 ,
         \12008 , \12009 , \12010_nR295b , \12011 , \12012 , \12013 , \12014 , \12015 , \12016 , \12017 ,
         \12018 , \12019 , \12020 , \12021 , \12022 , \12023 , \12024 , \12025 , \12026 , \12027 ,
         \12028 , \12029 , \12030 , \12031 , \12032 , \12033 , \12034 , \12035 , \12036 , \12037 ,
         \12038 , \12039 , \12040_nR27d1 , \12041 , \12042 , \12043 , \12044 , \12045 , \12046 , \12047 ,
         \12048 , \12049 , \12050 , \12051 , \12052 , \12053 , \12054 , \12055 , \12056 , \12057 ,
         \12058 , \12059 , \12060 , \12061 , \12062 , \12063 , \12064 , \12065 , \12066 , \12067 ,
         \12068 , \12069 , \12070_nR27cf , \12071 , \12072 , \12073 , \12074 , \12075 , \12076 , \12077 ,
         \12078 , \12079 , \12080 , \12081 , \12082 , \12083 , \12084 , \12085 , \12086 , \12087 ,
         \12088 , \12089 , \12090 , \12091 , \12092 , \12093 , \12094 , \12095 , \12096 , \12097 ,
         \12098 , \12099 , \12100_nR2689 , \12101 , \12102 , \12103 , \12104 , \12105 , \12106 , \12107 ,
         \12108 , \12109 , \12110 , \12111 , \12112 , \12113 , \12114 , \12115 , \12116 , \12117 ,
         \12118 , \12119 , \12120 , \12121 , \12122 , \12123 , \12124 , \12125 , \12126 , \12127 ,
         \12128 , \12129 , \12130_nR2687 , \12131 , \12132 , \12133 , \12134 , \12135 , \12136 , \12137 ,
         \12138 , \12139 , \12140 , \12141 , \12142 , \12143 , \12144 , \12145 , \12146 , \12147 ,
         \12148 , \12149 , \12150 , \12151 , \12152 , \12153 , \12154 , \12155 , \12156 , \12157 ,
         \12158 , \12159 , \12160_nR25a9 , \12161 , \12162 , \12163 , \12164 , \12165 , \12166 , \12167 ,
         \12168 , \12169 , \12170 , \12171 , \12172 , \12173 , \12174 , \12175 , \12176 , \12177 ,
         \12178 , \12179 , \12180 , \12181 , \12182 , \12183 , \12184 , \12185 , \12186 , \12187 ,
         \12188 , \12189 , \12190_nR25ab , \12191 , \12192 , \12193 , \12194 , \12195 , \12196 , \12197 ,
         \12198 , \12199 , \12200 , \12201 , \12202 , \12203 , \12204 , \12205 , \12206 , \12207 ,
         \12208 , \12209 , \12210 , \12211 , \12212 , \12213 , \12214 , \12215 , \12216 , \12217 ,
         \12218 , \12219 , \12220_nR2433 , \12221 , \12222 , \12223 , \12224 , \12225 , \12226 , \12227 ,
         \12228 , \12229 , \12230 , \12231 , \12232 , \12233 , \12234 , \12235 , \12236 , \12237 ,
         \12238 , \12239 , \12240 , \12241 , \12242 , \12243 , \12244 , \12245 , \12246 , \12247 ,
         \12248 , \12249 , \12250_nR2435 , \12251 , \12252 , \12253 , \12254 , \12255 , \12256 , \12257 ,
         \12258 , \12259 , \12260 , \12261 , \12262 , \12263 , \12264 , \12265 , \12266 , \12267 ,
         \12268 , \12269 , \12270 , \12271 , \12272 , \12273 , \12274 , \12275 , \12276 , \12277 ,
         \12278 , \12279 , \12280 , \12281 , \12282 , \12283 , \12284 , \12285 , \12286 , \12287 ,
         \12288 , \12289 , \12290 , \12291 , \12292 , \12293 , \12294 , \12295 , \12296 , \12297 ,
         \12298 , \12299 , \12300 , \12301 , \12302 , \12303 , \12304 , \12305 , \12306 , \12307 ,
         \12308 , \12309 , \12310 , \12311 , \12312 , \12313 , \12314 , \12315 , \12316 , \12317 ,
         \12318 , \12319 , \12320 , \12321 , \12322 , \12323 , \12324 , \12325 , \12326 , \12327 ,
         \12328 , \12329 , \12330 , \12331 , \12332 , \12333 , \12334 , \12335 , \12336 , \12337 ,
         \12338 , \12339 , \12340 , \12341 , \12342 , \12343 , \12344 , \12345 , \12346 , \12347 ,
         \12348 , \12349 , \12350 , \12351 , \12352 , \12353 , \12354 , \12355 , \12356 , \12357 ,
         \12358 , \12359 , \12360 , \12361 , \12362 , \12363 , \12364 , \12365 , \12366 , \12367 ,
         \12368 , \12369 , \12370_nR3379 , \12371 , \12372 , \12373 , \12374 , \12375 , \12376 , \12377 ,
         \12378 , \12379 , \12380 , \12381 , \12382 , \12383 , \12384 , \12385 , \12386 , \12387 ,
         \12388 , \12389 , \12390 , \12391 , \12392 , \12393 , \12394 , \12395 , \12396 , \12397 ,
         \12398 , \12399 , \12400 , \12401 , \12402 , \12403 , \12404 , \12405 , \12406 , \12407 ,
         \12408 , \12409 , \12410 , \12411 , \12412 , \12413 , \12414 , \12415 , \12416 , \12417 ,
         \12418_nR349f , \12419 , \12420 , \12421 , \12422 , \12423 , \12424 , \12425 , \12426 , \12427 ,
         \12428 , \12429 , \12430 , \12431 , \12432 , \12433 , \12434 , \12435 , \12436 , \12437 ,
         \12438 , \12439 , \12440 , \12441 , \12442 , \12443 , \12444 , \12445 , \12446 , \12447 ,
         \12448 , \12449 , \12450 , \12451 , \12452 , \12453 , \12454 , \12455 , \12456 , \12457 ,
         \12458 , \12459 , \12460 , \12461 , \12462 , \12463 , \12464 , \12465 , \12466 , \12467 ,
         \12468 , \12469 , \12470_nR3271 , \12471 , \12472 , \12473 , \12474 , \12475 , \12476 , \12477 ,
         \12478 , \12479 , \12480 , \12481 , \12482 , \12483 , \12484 , \12485 , \12486 , \12487 ,
         \12488 , \12489 , \12490 , \12491 , \12492 , \12493 , \12494 , \12495 , \12496 , \12497 ,
         \12498 , \12499 , \12500 , \12501 , \12502 , \12503 , \12504 , \12505 , \12506 , \12507 ,
         \12508 , \12509 , \12510 , \12511 , \12512 , \12513 , \12514 , \12515 , \12516 , \12517 ,
         \12518 , \12519 , \12520 , \12521 , \12522 , \12523 , \12524 , \12525 , \12526 , \12527 ,
         \12528 , \12529 , \12530 , \12531 , \12532 , \12533 , \12534 , \12535 , \12536 , \12537 ,
         \12538 , \12539 , \12540 , \12541 , \12542 , \12543 , \12544 , \12545 , \12546 , \12547 ,
         \12548 , \12549_nR3150 , \12550 , \12551 , \12552 , \12553 , \12554 , \12555 , \12556 , \12557 ,
         \12558 , \12559 , \12560 , \12561 , \12562 , \12563 , \12564 , \12565 , \12566 , \12567 ,
         \12568 , \12569 , \12570 , \12571 , \12572 , \12573 , \12574 , \12575 , \12576 , \12577 ,
         \12578 , \12579 , \12580 , \12581 , \12582 , \12583 , \12584 , \12585 , \12586 , \12587 ,
         \12588 , \12589 , \12590 , \12591 , \12592 , \12593 , \12594 , \12595 , \12596 , \12597 ,
         \12598 , \12599 , \12600 , \12601 , \12602 , \12603 , \12604 , \12605 , \12606 , \12607 ,
         \12608 , \12609 , \12610 , \12611 , \12612 , \12613 , \12614 , \12615 , \12616 , \12617 ,
         \12618 , \12619 , \12620 , \12621 , \12622 , \12623 , \12624 , \12625 , \12626 , \12627 ,
         \12628 , \12629 , \12630 , \12631_nR3038 , \12632 , \12633 , \12634 , \12635 , \12636 , \12637 ,
         \12638 , \12639 , \12640 , \12641 , \12642 , \12643 , \12644 , \12645 , \12646 , \12647 ,
         \12648 , \12649 , \12650 , \12651 , \12652 , \12653 , \12654 , \12655 , \12656 , \12657 ,
         \12658 , \12659 , \12660 , \12661 , \12662 , \12663 , \12664 , \12665 , \12666 , \12667 ,
         \12668 , \12669 , \12670 , \12671 , \12672 , \12673 , \12674 , \12675 , \12676 , \12677 ,
         \12678 , \12679 , \12680 , \12681 , \12682 , \12683 , \12684 , \12685 , \12686 , \12687 ,
         \12688 , \12689 , \12690_nR2f21 , \12691 , \12692 , \12693 , \12694 , \12695 , \12696 , \12697 ,
         \12698 , \12699 , \12700 , \12701 , \12702 , \12703 , \12704 , \12705 , \12706 , \12707 ,
         \12708 , \12709 , \12710 , \12711 , \12712 , \12713 , \12714 , \12715 , \12716 , \12717 ,
         \12718 , \12719 , \12720 , \12721 , \12722 , \12723 , \12724 , \12725 , \12726 , \12727 ,
         \12728 , \12729 , \12730 , \12731 , \12732 , \12733 , \12734 , \12735 , \12736 , \12737 ,
         \12738 , \12739 , \12740 , \12741 , \12742 , \12743 , \12744 , \12745 , \12746 , \12747 ,
         \12748 , \12749 , \12750 , \12751 , \12752 , \12753 , \12754 , \12755 , \12756 , \12757 ,
         \12758 , \12759 , \12760 , \12761 , \12762_nR2e29 , \12763 , \12764 , \12765 , \12766 , \12767 ,
         \12768 , \12769 , \12770 , \12771 , \12772 , \12773 , \12774 , \12775 , \12776 , \12777 ,
         \12778 , \12779 , \12780 , \12781 , \12782 , \12783 , \12784 , \12785 , \12786 , \12787 ,
         \12788 , \12789 , \12790 , \12791 , \12792 , \12793 , \12794 , \12795 , \12796 , \12797 ,
         \12798 , \12799 , \12800 , \12801 , \12802 , \12803 , \12804 , \12805 , \12806 , \12807 ,
         \12808 , \12809 , \12810 , \12811 , \12812 , \12813 , \12814 , \12815 , \12816 , \12817 ,
         \12818 , \12819 , \12820 , \12821 , \12822 , \12823 , \12824 , \12825 , \12826 , \12827 ,
         \12828 , \12829 , \12830 , \12831 , \12832 , \12833 , \12834 , \12835 , \12836 , \12837 ,
         \12838 , \12839 , \12840 , \12841 , \12842 , \12843_nR2d1d , \12844 , \12845 , \12846 , \12847 ,
         \12848 , \12849 , \12850 , \12851 , \12852 , \12853 , \12854 , \12855 , \12856 , \12857 ,
         \12858 , \12859 , \12860 , \12861 , \12862 , \12863 , \12864 , \12865 , \12866 , \12867 ,
         \12868 , \12869 , \12870 , \12871 , \12872 , \12873 , \12874 , \12875 , \12876 , \12877 ,
         \12878 , \12879 , \12880 , \12881 , \12882 , \12883 , \12884 , \12885 , \12886 , \12887 ,
         \12888 , \12889 , \12890 , \12891 , \12892 , \12893 , \12894 , \12895 , \12896 , \12897 ,
         \12898 , \12899 , \12900 , \12901 , \12902 , \12903 , \12904 , \12905 , \12906 , \12907 ,
         \12908 , \12909 , \12910 , \12911 , \12912 , \12913 , \12914 , \12915 , \12916 , \12917 ,
         \12918 , \12919 , \12920 , \12921 , \12922 , \12923 , \12924 , \12925 , \12926 , \12927 ,
         \12928 , \12929 , \12930 , \12931 , \12932 , \12933 , \12934 , \12935 , \12936 , \12937 ,
         \12938 , \12939 , \12940 , \12941 , \12942 , \12943 , \12944 , \12945 , \12946 , \12947 ,
         \12948 , \12949 , \12950 , \12951 , \12952_nR2c3a , \12953 , \12954 , \12955 , \12956 , \12957 ,
         \12958 , \12959 , \12960 , \12961 , \12962 , \12963 , \12964 , \12965 , \12966 , \12967 ,
         \12968 , \12969 , \12970 , \12971 , \12972 , \12973 , \12974 , \12975 , \12976 , \12977 ,
         \12978 , \12979 , \12980 , \12981 , \12982 , \12983 , \12984 , \12985 , \12986 , \12987 ,
         \12988 , \12989 , \12990 , \12991 , \12992 , \12993 , \12994 , \12995 , \12996 , \12997 ,
         \12998 , \12999 , \13000 , \13001 , \13002 , \13003 , \13004 , \13005 , \13006 , \13007 ,
         \13008 , \13009 , \13010 , \13011 , \13012 , \13013 , \13014 , \13015 , \13016 , \13017 ,
         \13018 , \13019 , \13020 , \13021 , \13022 , \13023 , \13024 , \13025 , \13026 , \13027 ,
         \13028 , \13029 , \13030 , \13031 , \13032 , \13033 , \13034 , \13035 , \13036 , \13037 ,
         \13038 , \13039 , \13040 , \13041 , \13042 , \13043 , \13044 , \13045 , \13046 , \13047 ,
         \13048 , \13049 , \13050 , \13051 , \13052 , \13053 , \13054 , \13055 , \13056 , \13057 ,
         \13058 , \13059 , \13060 , \13061 , \13062 , \13063 , \13064 , \13065 , \13066 , \13067 ,
         \13068 , \13069 , \13070 , \13071 , \13072 , \13073 , \13074 , \13075 , \13076 , \13077 ,
         \13078 , \13079 , \13080 , \13081 , \13082 , \13083 , \13084 , \13085 , \13086 , \13087 ,
         \13088 , \13089 , \13090 , \13091 , \13092 , \13093 , \13094 , \13095 , \13096 , \13097 ,
         \13098 , \13099 , \13100 , \13101 , \13102 , \13103 , \13104 , \13105 , \13106 , \13107 ,
         \13108 , \13109 , \13110 , \13111 , \13112 , \13113 , \13114 , \13115 , \13116 , \13117 ,
         \13118 , \13119 , \13120 , \13121 , \13122 , \13123 , \13124 , \13125 , \13126 , \13127 ,
         \13128 , \13129 , \13130 , \13131 , \13132 , \13133 , \13134 , \13135 , \13136 , \13137 ,
         \13138 , \13139 , \13140 , \13141 , \13142 , \13143 , \13144 , \13145 , \13146 , \13147 ,
         \13148 , \13149 , \13150 , \13151 , \13152 , \13153 , \13154 , \13155 , \13156 , \13157 ,
         \13158 , \13159 , \13160 , \13161 , \13162 , \13163 , \13164 , \13165 , \13166 , \13167 ,
         \13168 , \13169 , \13170 , \13171 , \13172 , \13173 , \13174 , \13175_nR2b34 , \13176 , \13177 ,
         \13178 , \13179 , \13180 , \13181 , \13182 , \13183 , \13184 , \13185 , \13186 , \13187 ,
         \13188 , \13189 , \13190 , \13191 , \13192 , \13193 , \13194 , \13195 , \13196 , \13197 ,
         \13198 , \13199 , \13200 , \13201 , \13202 , \13203 , \13204 , \13205 , \13206 , \13207 ,
         \13208 , \13209 , \13210 , \13211 , \13212 , \13213 , \13214 , \13215 , \13216 , \13217 ,
         \13218 , \13219 , \13220 , \13221 , \13222 , \13223 , \13224 , \13225 , \13226 , \13227 ,
         \13228 , \13229 , \13230 , \13231 , \13232 , \13233 , \13234 , \13235 , \13236 , \13237 ,
         \13238 , \13239 , \13240 , \13241 , \13242 , \13243 , \13244 , \13245 , \13246 , \13247 ,
         \13248 , \13249 , \13250 , \13251 , \13252 , \13253 , \13254 , \13255 , \13256 , \13257 ,
         \13258 , \13259 , \13260 , \13261 , \13262 , \13263 , \13264 , \13265 , \13266 , \13267 ,
         \13268 , \13269 , \13270 , \13271 , \13272 , \13273 , \13274 , \13275 , \13276 , \13277 ,
         \13278 , \13279 , \13280 , \13281 , \13282 , \13283 , \13284 , \13285 , \13286 , \13287 ,
         \13288 , \13289 , \13290 , \13291 , \13292 , \13293 , \13294 , \13295 , \13296 , \13297 ,
         \13298 , \13299 , \13300 , \13301 , \13302 , \13303 , \13304 , \13305 , \13306 , \13307 ,
         \13308 , \13309 , \13310 , \13311 , \13312 , \13313 , \13314 , \13315 , \13316 , \13317 ,
         \13318 , \13319 , \13320 , \13321 , \13322_nR2a51 , \13323 , \13324 , \13325 , \13326 , \13327 ,
         \13328 , \13329 , \13330 , \13331 , \13332 , \13333 , \13334 , \13335 , \13336 , \13337 ,
         \13338 , \13339 , \13340 , \13341 , \13342 , \13343 , \13344 , \13345 , \13346 , \13347 ,
         \13348 , \13349 , \13350 , \13351 , \13352 , \13353 , \13354 , \13355 , \13356 , \13357 ,
         \13358 , \13359 , \13360 , \13361 , \13362 , \13363 , \13364 , \13365 , \13366 , \13367 ,
         \13368 , \13369 , \13370 , \13371 , \13372 , \13373 , \13374 , \13375 , \13376 , \13377 ,
         \13378 , \13379 , \13380 , \13381 , \13382 , \13383 , \13384 , \13385 , \13386 , \13387 ,
         \13388_nR2979 , \13389 , \13390 , \13391 , \13392 , \13393 , \13394 , \13395 , \13396 , \13397 ,
         \13398 , \13399 , \13400 , \13401 , \13402 , \13403 , \13404 , \13405 , \13406 , \13407 ,
         \13408 , \13409 , \13410 , \13411 , \13412 , \13413 , \13414 , \13415 , \13416 , \13417 ,
         \13418 , \13419 , \13420 , \13421 , \13422 , \13423 , \13424 , \13425 , \13426 , \13427 ,
         \13428 , \13429 , \13430 , \13431 , \13432 , \13433 , \13434 , \13435 , \13436 , \13437 ,
         \13438 , \13439 , \13440 , \13441 , \13442 , \13443 , \13444 , \13445 , \13446 , \13447 ,
         \13448 , \13449 , \13450 , \13451 , \13452 , \13453 , \13454 , \13455 , \13456 , \13457 ,
         \13458 , \13459 , \13460 , \13461 , \13462 , \13463 , \13464 , \13465 , \13466 , \13467 ,
         \13468 , \13469 , \13470 , \13471 , \13472 , \13473 , \13474 , \13475 , \13476 , \13477 ,
         \13478 , \13479 , \13480 , \13481 , \13482 , \13483 , \13484 , \13485 , \13486 , \13487 ,
         \13488 , \13489 , \13490 , \13491 , \13492 , \13493 , \13494 , \13495 , \13496 , \13497 ,
         \13498 , \13499 , \13500 , \13501 , \13502 , \13503 , \13504 , \13505 , \13506 , \13507 ,
         \13508 , \13509 , \13510 , \13511 , \13512 , \13513 , \13514 , \13515 , \13516 , \13517 ,
         \13518 , \13519 , \13520 , \13521 , \13522 , \13523 , \13524 , \13525 , \13526 , \13527 ,
         \13528 , \13529 , \13530 , \13531 , \13532 , \13533 , \13534 , \13535 , \13536 , \13537 ,
         \13538 , \13539 , \13540 , \13541 , \13542 , \13543 , \13544 , \13545 , \13546 , \13547 ,
         \13548 , \13549 , \13550 , \13551 , \13552 , \13553 , \13554 , \13555 , \13556 , \13557 ,
         \13558 , \13559 , \13560 , \13561 , \13562 , \13563 , \13564 , \13565 , \13566 , \13567 ,
         \13568 , \13569 , \13570 , \13571 , \13572 , \13573 , \13574 , \13575_nR27ee , \13576 , \13577 ,
         \13578 , \13579 , \13580 , \13581 , \13582 , \13583 , \13584 , \13585 , \13586 , \13587 ,
         \13588 , \13589 , \13590 , \13591 , \13592 , \13593 , \13594 , \13595 , \13596 , \13597 ,
         \13598 , \13599 , \13600 , \13601 , \13602 , \13603 , \13604 , \13605 , \13606 , \13607_nR28bb ,
         \13608 , \13609 , \13610 , \13611 , \13612 , \13613 , \13614 , \13615 , \13616 , \13617 ,
         \13618 , \13619 , \13620 , \13621 , \13622 , \13623 , \13624 , \13625 , \13626 , \13627 ,
         \13628 , \13629 , \13630 , \13631 , \13632 , \13633 , \13634 , \13635 , \13636 , \13637 ,
         \13638 , \13639 , \13640 , \13641 , \13642 , \13643 , \13644 , \13645 , \13646 , \13647 ,
         \13648 , \13649 , \13650 , \13651 , \13652 , \13653 , \13654 , \13655 , \13656 , \13657 ,
         \13658 , \13659 , \13660 , \13661 , \13662 , \13663 , \13664 , \13665 , \13666 , \13667 ,
         \13668 , \13669 , \13670 , \13671 , \13672 , \13673 , \13674 , \13675 , \13676 , \13677 ,
         \13678 , \13679 , \13680 , \13681 , \13682 , \13683 , \13684 , \13685 , \13686 , \13687 ,
         \13688 , \13689 , \13690 , \13691 , \13692 , \13693 , \13694 , \13695 , \13696 , \13697 ,
         \13698 , \13699 , \13700 , \13701 , \13702 , \13703 , \13704 , \13705 , \13706 , \13707 ,
         \13708 , \13709 , \13710 , \13711 , \13712 , \13713 , \13714 , \13715 , \13716 , \13717 ,
         \13718 , \13719 , \13720 , \13721 , \13722 , \13723 , \13724 , \13725 , \13726 , \13727 ,
         \13728 , \13729 , \13730 , \13731 , \13732 , \13733 , \13734 , \13735 , \13736 , \13737 ,
         \13738 , \13739 , \13740 , \13741 , \13742 , \13743 , \13744 , \13745 , \13746 , \13747 ,
         \13748 , \13749 , \13750 , \13751 , \13752 , \13753 , \13754 , \13755 , \13756 , \13757 ,
         \13758 , \13759 , \13760 , \13761 , \13762 , \13763 , \13764 , \13765 , \13766 , \13767 ,
         \13768 , \13769 , \13770 , \13771 , \13772 , \13773 , \13774 , \13775 , \13776 , \13777 ,
         \13778 , \13779 , \13780 , \13781 , \13782 , \13783 , \13784 , \13785 , \13786 , \13787 ,
         \13788 , \13789 , \13790 , \13791 , \13792 , \13793 , \13794 , \13795 , \13796 , \13797 ,
         \13798 , \13799 , \13800 , \13801 , \13802 , \13803 , \13804 , \13805 , \13806 , \13807 ,
         \13808 , \13809 , \13810 , \13811 , \13812 , \13813 , \13814 , \13815 , \13816 , \13817 ,
         \13818 , \13819 , \13820 , \13821 , \13822 , \13823 , \13824 , \13825 , \13826_nR26a6 , \13827 ,
         \13828 , \13829 , \13830 , \13831 , \13832 , \13833 , \13834 , \13835 , \13836 , \13837 ,
         \13838 , \13839 , \13840 , \13841 , \13842 , \13843 , \13844 , \13845 , \13846 , \13847 ,
         \13848 , \13849 , \13850 , \13851 , \13852 , \13853 , \13854 , \13855 , \13856 , \13857 ,
         \13858_nR274c , \13859 , \13860 , \13861 , \13862 , \13863 , \13864 , \13865 , \13866 , \13867 ,
         \13868 , \13869 , \13870 , \13871 , \13872 , \13873 , \13874 , \13875 , \13876 , \13877 ,
         \13878 , \13879 , \13880 , \13881 , \13882 , \13883 , \13884 , \13885 , \13886 , \13887 ,
         \13888 , \13889 , \13890 , \13891 , \13892 , \13893 , \13894 , \13895 , \13896 , \13897 ,
         \13898 , \13899 , \13900 , \13901 , \13902 , \13903 , \13904 , \13905 , \13906 , \13907 ,
         \13908 , \13909 , \13910 , \13911 , \13912 , \13913 , \13914 , \13915 , \13916 , \13917 ,
         \13918 , \13919 , \13920 , \13921 , \13922 , \13923 , \13924 , \13925 , \13926 , \13927 ,
         \13928 , \13929 , \13930 , \13931 , \13932 , \13933 , \13934 , \13935 , \13936 , \13937 ,
         \13938 , \13939 , \13940 , \13941 , \13942 , \13943 , \13944 , \13945 , \13946 , \13947 ,
         \13948 , \13949 , \13950 , \13951 , \13952 , \13953 , \13954 , \13955 , \13956 , \13957 ,
         \13958 , \13959 , \13960 , \13961 , \13962 , \13963 , \13964 , \13965 , \13966 , \13967 ,
         \13968 , \13969 , \13970 , \13971 , \13972 , \13973 , \13974 , \13975 , \13976 , \13977 ,
         \13978 , \13979 , \13980 , \13981 , \13982 , \13983 , \13984 , \13985 , \13986 , \13987 ,
         \13988 , \13989 , \13990 , \13991 , \13992 , \13993 , \13994 , \13995 , \13996 , \13997 ,
         \13998 , \13999 , \14000 , \14001 , \14002 , \14003 , \14004 , \14005 , \14006 , \14007 ,
         \14008 , \14009 , \14010 , \14011 , \14012 , \14013 , \14014 , \14015 , \14016 , \14017 ,
         \14018 , \14019 , \14020 , \14021 , \14022 , \14023 , \14024 , \14025 , \14026 , \14027 ,
         \14028 , \14029 , \14030 , \14031 , \14032 , \14033 , \14034 , \14035 , \14036 , \14037 ,
         \14038 , \14039 , \14040 , \14041 , \14042 , \14043 , \14044 , \14045 , \14046 , \14047 ,
         \14048 , \14049 , \14050 , \14051 , \14052 , \14053 , \14054 , \14055 , \14056 , \14057 ,
         \14058 , \14059 , \14060 , \14061 , \14062 , \14063 , \14064 , \14065 , \14066 , \14067 ,
         \14068 , \14069_nR2626 , \14070 , \14071 , \14072 , \14073 , \14074 , \14075 , \14076 , \14077 ,
         \14078 , \14079 , \14080 , \14081 , \14082 , \14083 , \14084 , \14085 , \14086 , \14087 ,
         \14088 , \14089 , \14090 , \14091 , \14092 , \14093 , \14094 , \14095 , \14096 , \14097 ,
         \14098 , \14099 , \14100 , \14101 , \14102 , \14103 , \14104 , \14105 , \14106 , \14107 ,
         \14108 , \14109 , \14110 , \14111 , \14112 , \14113 , \14114 , \14115 , \14116 , \14117 ,
         \14118 , \14119 , \14120 , \14121 , \14122 , \14123 , \14124 , \14125 , \14126 , \14127 ,
         \14128 , \14129 , \14130 , \14131 , \14132 , \14133 , \14134 , \14135 , \14136 , \14137 ,
         \14138 , \14139 , \14140 , \14141 , \14142 , \14143 , \14144 , \14145 , \14146 , \14147 ,
         \14148 , \14149 , \14150 , \14151 , \14152 , \14153 , \14154 , \14155 , \14156 , \14157 ,
         \14158 , \14159 , \14160 , \14161 , \14162 , \14163 , \14164 , \14165 , \14166 , \14167 ,
         \14168 , \14169 , \14170 , \14171 , \14172_nR25a7 , \14173 , \14174 , \14175 , \14176 , \14177 ,
         \14178 , \14179 , \14180 , \14181 , \14182 , \14183 , \14184 , \14185 , \14186 , \14187 ,
         \14188 , \14189 , \14190 , \14191 , \14192 , \14193 , \14194 , \14195 , \14196 , \14197 ,
         \14198 , \14199 , \14200 , \14201 , \14202 , \14203 , \14204 , \14205 , \14206 , \14207 ,
         \14208 , \14209 , \14210 , \14211 , \14212 , \14213 , \14214 , \14215 , \14216 , \14217 ,
         \14218 , \14219 , \14220 , \14221 , \14222 , \14223 , \14224 , \14225 , \14226 , \14227 ,
         \14228 , \14229 , \14230 , \14231 , \14232 , \14233 , \14234 , \14235 , \14236 , \14237 ,
         \14238 , \14239 , \14240 , \14241 , \14242 , \14243 , \14244 , \14245 , \14246 , \14247 ,
         \14248 , \14249 , \14250 , \14251 , \14252 , \14253 , \14254 , \14255 , \14256 , \14257 ,
         \14258 , \14259 , \14260 , \14261 , \14262 , \14263 , \14264 , \14265 , \14266 , \14267 ,
         \14268 , \14269 , \14270 , \14271 , \14272 , \14273 , \14274 , \14275 , \14276 , \14277 ,
         \14278 , \14279 , \14280 , \14281 , \14282 , \14283 , \14284 , \14285 , \14286 , \14287 ,
         \14288 , \14289 , \14290 , \14291 , \14292 , \14293 , \14294 , \14295 , \14296 , \14297 ,
         \14298 , \14299 , \14300 , \14301 , \14302 , \14303 , \14304 , \14305 , \14306 , \14307 ,
         \14308 , \14309 , \14310 , \14311 , \14312 , \14313 , \14314 , \14315 , \14316 , \14317 ,
         \14318 , \14319 , \14320 , \14321 , \14322 , \14323 , \14324 , \14325 , \14326 , \14327 ,
         \14328 , \14329 , \14330 , \14331 , \14332 , \14333 , \14334 , \14335 , \14336 , \14337 ,
         \14338 , \14339 , \14340 , \14341 , \14342 , \14343 , \14344 , \14345 , \14346 , \14347 ,
         \14348 , \14349 , \14350 , \14351 , \14352 , \14353 , \14354 , \14355 , \14356 , \14357 ,
         \14358_nR2538 , \14359 , \14360 , \14361 , \14362 , \14363 , \14364 , \14365 , \14366 , \14367 ,
         \14368 , \14369 , \14370 , \14371 , \14372 , \14373 , \14374 , \14375 , \14376 , \14377 ,
         \14378 , \14379 , \14380 , \14381 , \14382 , \14383 , \14384 , \14385 , \14386 , \14387 ,
         \14388 , \14389 , \14390 , \14391 , \14392 , \14393 , \14394 , \14395 , \14396 , \14397 ,
         \14398 , \14399 , \14400 , \14401 , \14402 , \14403 , \14404 , \14405 , \14406 , \14407 ,
         \14408 , \14409 , \14410 , \14411 , \14412 , \14413_nR2430 , \14414 , \14415 , \14416 , \14417 ,
         \14418 , \14419 , \14420 , \14421 , \14422 , \14423 , \14424 , \14425 , \14426 , \14427 ,
         \14428 , \14429 , \14430 , \14431 , \14432 , \14433 , \14434 , \14435 , \14436 , \14437 ,
         \14438 , \14439 , \14440 , \14441 , \14442 , \14443 , \14444 , \14445 , \14446 , \14447 ,
         \14448 , \14449 , \14450 , \14451 , \14452 , \14453 , \14454 , \14455 , \14456 , \14457 ,
         \14458 , \14459 , \14460 , \14461 , \14462 , \14463 , \14464 , \14465 , \14466 , \14467 ,
         \14468 , \14469 , \14470 , \14471 , \14472 , \14473 , \14474 , \14475 , \14476 , \14477 ,
         \14478 , \14479 , \14480 , \14481 , \14482 , \14483 , \14484 , \14485 , \14486 , \14487 ,
         \14488 , \14489 , \14490 , \14491 , \14492 , \14493 , \14494 , \14495 , \14496 , \14497 ,
         \14498 , \14499 , \14500 , \14501 , \14502 , \14503 , \14504 , \14505 , \14506 , \14507 ,
         \14508 , \14509 , \14510 , \14511 , \14512 , \14513 , \14514 , \14515 , \14516 , \14517 ,
         \14518 , \14519 , \14520 , \14521 , \14522 , \14523 , \14524 , \14525 , \14526 , \14527 ,
         \14528 , \14529 , \14530 , \14531 , \14532 , \14533 , \14534 , \14535 , \14536 , \14537 ,
         \14538 , \14539 , \14540 , \14541 , \14542 , \14543 , \14544 , \14545 , \14546 , \14547 ,
         \14548 , \14549 , \14550 , \14551 , \14552 , \14553 , \14554 , \14555 , \14556 , \14557 ,
         \14558 , \14559 , \14560 , \14561 , \14562 , \14563 , \14564 , \14565 , \14566 , \14567 ,
         \14568 , \14569 , \14570 , \14571 , \14572 , \14573 , \14574 , \14575 , \14576 , \14577 ,
         \14578 , \14579 , \14580 , \14581 , \14582 , \14583 , \14584 , \14585 , \14586 , \14587 ,
         \14588 , \14589 , \14590 , \14591 , \14592 , \14593 , \14594 , \14595 , \14596 , \14597 ,
         \14598 , \14599 , \14600 , \14601 , \14602 , \14603 , \14604 , \14605 , \14606 , \14607 ,
         \14608 , \14609 , \14610 , \14611 , \14612 , \14613 , \14614 , \14615 , \14616 , \14617 ,
         \14618 , \14619 , \14620 , \14621 , \14622 , \14623 , \14624 , \14625 , \14626 , \14627 ,
         \14628 , \14629 , \14630 , \14631 , \14632 , \14633 , \14634 , \14635 , \14636 , \14637 ,
         \14638 , \14639 , \14640 , \14641 , \14642 , \14643 , \14644 , \14645 , \14646 , \14647 ,
         \14648 , \14649 , \14650 , \14651 , \14652 , \14653 , \14654 , \14655 , \14656 , \14657 ,
         \14658 , \14659 , \14660 , \14661 , \14662 , \14663 , \14664 , \14665 , \14666 , \14667 ,
         \14668 , \14669 , \14670 , \14671 , \14672 , \14673 , \14674 , \14675 , \14676 , \14677 ,
         \14678 , \14679 , \14680 , \14681 , \14682 , \14683 , \14684 , \14685 , \14686 , \14687 ,
         \14688 , \14689 , \14690 , \14691 , \14692 , \14693 , \14694 , \14695 , \14696 , \14697 ,
         \14698 , \14699 , \14700 , \14701 , \14702 , \14703 , \14704 , \14705 , \14706 , \14707 ,
         \14708 , \14709 , \14710 , \14711 , \14712 , \14713 , \14714 , \14715 , \14716 , \14717 ,
         \14718 , \14719 , \14720 , \14721 , \14722 , \14723 , \14724 , \14725 , \14726 , \14727 ,
         \14728 , \14729 , \14730 , \14731 , \14732 , \14733 , \14734 , \14735 , \14736 , \14737 ,
         \14738 , \14739 , \14740 , \14741 , \14742 , \14743 , \14744 , \14745 , \14746 , \14747 ,
         \14748 , \14749 , \14750 , \14751 , \14752 , \14753 , \14754 , \14755 , \14756 , \14757 ,
         \14758 , \14759 , \14760 , \14761 , \14762 , \14763 , \14764 , \14765 , \14766 , \14767 ,
         \14768 , \14769 , \14770 , \14771 , \14772 , \14773 , \14774 , \14775 , \14776 , \14777 ,
         \14778 , \14779 , \14780 , \14781 , \14782 , \14783 , \14784 , \14785 , \14786 , \14787 ,
         \14788 , \14789 , \14790 , \14791 , \14792 , \14793 , \14794 , \14795 , \14796 , \14797 ,
         \14798 , \14799 , \14800 , \14801 , \14802 , \14803 , \14804 , \14805 , \14806 , \14807 ,
         \14808 , \14809 , \14810 , \14811 , \14812 , \14813 , \14814 , \14815 , \14816 , \14817 ,
         \14818 , \14819 , \14820 , \14821 , \14822 , \14823 , \14824 , \14825 , \14826 , \14827 ,
         \14828 , \14829 , \14830 , \14831 , \14832 , \14833 , \14834 , \14835 , \14836 , \14837 ,
         \14838 , \14839 , \14840 , \14841 , \14842 , \14843 , \14844 , \14845 , \14846 , \14847 ,
         \14848 , \14849 , \14850 , \14851 , \14852 , \14853 , \14854 , \14855 , \14856 , \14857 ,
         \14858 , \14859 , \14860 , \14861 , \14862 , \14863 , \14864 , \14865 , \14866 , \14867 ,
         \14868 , \14869 , \14870 , \14871 , \14872 , \14873 , \14874 , \14875 , \14876 , \14877 ,
         \14878 , \14879 , \14880 , \14881 , \14882 , \14883 , \14884 , \14885 , \14886 , \14887 ,
         \14888 , \14889 , \14890 , \14891 , \14892 , \14893 , \14894 , \14895 , \14896 , \14897 ,
         \14898 , \14899 , \14900 , \14901 , \14902 , \14903 , \14904 , \14905 , \14906 , \14907 ,
         \14908 , \14909 , \14910 , \14911 , \14912 , \14913 , \14914 , \14915 , \14916 , \14917 ,
         \14918 , \14919 , \14920 , \14921 , \14922 , \14923 , \14924 , \14925 , \14926 , \14927 ,
         \14928 , \14929 , \14930 , \14931 , \14932 , \14933 , \14934 , \14935 , \14936 , \14937 ,
         \14938 , \14939 , \14940 , \14941 , \14942 , \14943 , \14944 , \14945 , \14946 , \14947 ,
         \14948 , \14949 , \14950 , \14951 , \14952 , \14953 , \14954 , \14955 , \14956 , \14957 ,
         \14958 , \14959 , \14960 , \14961 , \14962 , \14963 , \14964 , \14965 , \14966 , \14967 ,
         \14968 , \14969 , \14970 , \14971 , \14972 , \14973 , \14974 , \14975 , \14976 , \14977 ,
         \14978 , \14979 , \14980 , \14981 , \14982 , \14983 , \14984 , \14985 , \14986 , \14987 ,
         \14988 , \14989 , \14990 , \14991 , \14992 , \14993 , \14994 , \14995 , \14996 , \14997 ,
         \14998 , \14999 , \15000 , \15001 , \15002 , \15003 , \15004 , \15005 , \15006 , \15007 ,
         \15008 , \15009 , \15010 , \15011 , \15012 , \15013 , \15014 , \15015 , \15016 , \15017 ,
         \15018 , \15019 , \15020 , \15021 , \15022 , \15023 , \15024 , \15025 , \15026 , \15027 ,
         \15028 , \15029 , \15030 , \15031 , \15032 , \15033 , \15034 , \15035 , \15036 , \15037 ,
         \15038 , \15039 , \15040 , \15041 , \15042 , \15043 , \15044 , \15045 , \15046 , \15047 ,
         \15048 , \15049 , \15050 , \15051 , \15052 , \15053 , \15054 , \15055 , \15056 , \15057 ,
         \15058 , \15059 , \15060 , \15061 , \15062 , \15063 , \15064 , \15065 , \15066 , \15067 ,
         \15068 , \15069 , \15070 , \15071 , \15072 , \15073 , \15074 , \15075 , \15076 , \15077 ,
         \15078 , \15079 , \15080 , \15081 , \15082 , \15083 , \15084 , \15085 , \15086 , \15087 ,
         \15088 , \15089 , \15090 , \15091 , \15092 , \15093 , \15094 , \15095 , \15096 , \15097 ,
         \15098 , \15099 , \15100 , \15101 , \15102 , \15103 , \15104 , \15105 , \15106 , \15107 ,
         \15108 , \15109 , \15110 , \15111 , \15112 , \15113 , \15114 , \15115 , \15116 , \15117 ,
         \15118 , \15119 , \15120 , \15121 , \15122 , \15123 , \15124 , \15125 , \15126 , \15127 ,
         \15128 , \15129 , \15130 , \15131 , \15132 , \15133 , \15134 , \15135 , \15136 , \15137 ,
         \15138 , \15139 , \15140 , \15141 , \15142 , \15143 , \15144 , \15145 , \15146 , \15147 ,
         \15148 , \15149 , \15150 , \15151 , \15152 , \15153 , \15154 , \15155 , \15156 , \15157 ,
         \15158 , \15159 , \15160 , \15161 , \15162 , \15163 , \15164 , \15165 , \15166 , \15167 ,
         \15168 , \15169 , \15170 , \15171 , \15172 , \15173 , \15174 , \15175 , \15176 , \15177 ,
         \15178 , \15179 , \15180 , \15181 , \15182 , \15183 , \15184 , \15185 , \15186 , \15187 ,
         \15188 , \15189 , \15190 , \15191 , \15192 , \15193 , \15194 , \15195 , \15196 , \15197 ,
         \15198 , \15199 , \15200 , \15201 , \15202 , \15203 , \15204 , \15205 , \15206 , \15207 ,
         \15208 , \15209 , \15210 , \15211 , \15212 , \15213 , \15214 , \15215 , \15216 , \15217 ,
         \15218 , \15219 , \15220 , \15221 , \15222 , \15223 , \15224 , \15225 , \15226 , \15227 ,
         \15228 , \15229 , \15230 , \15231 , \15232 , \15233 , \15234 , \15235 , \15236 , \15237 ,
         \15238 , \15239 , \15240 , \15241 , \15242 , \15243 , \15244 , \15245 , \15246 , \15247 ,
         \15248 , \15249 , \15250 , \15251 , \15252 , \15253 , \15254 , \15255 , \15256 , \15257 ,
         \15258 , \15259 , \15260 , \15261 , \15262 , \15263 , \15264 , \15265 , \15266 , \15267 ,
         \15268 , \15269 , \15270 , \15271 , \15272 , \15273 , \15274 , \15275 , \15276 , \15277 ,
         \15278 , \15279 , \15280 , \15281 , \15282 , \15283 , \15284 , \15285 , \15286 , \15287 ,
         \15288 , \15289 , \15290 , \15291 , \15292 , \15293 , \15294 , \15295 , \15296 , \15297 ,
         \15298 , \15299 , \15300 , \15301 , \15302 , \15303 , \15304 , \15305 , \15306 , \15307 ,
         \15308 , \15309 , \15310 , \15311 , \15312 , \15313 , \15314 , \15315 , \15316 , \15317 ,
         \15318 , \15319 , \15320 , \15321 , \15322 , \15323 , \15324 , \15325 , \15326 , \15327_nR9a1 ,
         \15328 , \15329 , \15330 , \15331 , \15332_nR9a3 , \15333 , \15334 , \15335 , \15336_nR9c0 , \15337 ,
         \15338 , \15339_nR9c2 , \15340 , \15341 , \15342 , \15343 , \15344_nR984 , \15345 , \15346 , \15347 ,
         \15348_nR982 , \15349 , \15350 , \15351 , \15352 , \15353_nR965 , \15354 , \15355 , \15356 , \15357 ,
         \15358 , \15359_nR963 , \15360 , \15361 , \15362 , \15363_nR946 , \15364 , \15365 , \15366_nR944 , \15367 ,
         \15368 , \15369 , \15370 , \15371 , \15372_nR927 , \15373 , \15374 , \15375 , \15376 , \15377 ,
         \15378_nR925 , \15379 , \15380 , \15381 , \15382_nR906 , \15383 , \15384 , \15385 , \15386 , \15387 ,
         \15388_nR908 , \15389 , \15390 , \15391 , \15392_nR8e9 , \15393 , \15394 , \15395 , \15396 , \15397 ,
         \15398_nR8e7 , \15399 , \15400 , \15401 , \15402_nR8ca , \15403 , \15404 , \15405_nR8c8 , \15406 , \15407 ,
         \15408 , \15409 , \15410 , \15411_nR8ab , \15412 , \15413 , \15414 , \15415 , \15416 , \15417_nR8a9 ,
         \15418 , \15419 , \15420 , \15421_nR88c , \15422 , \15423 , \15424_nR88a , \15425 , \15426 , \15427 ,
         \15428 , \15429 , \15430_nR86d , \15431 , \15432 , \15433 , \15434 , \15435 , \15436_nR86b , \15437 ,
         \15438 , \15439 , \15440_nR84e , \15441 , \15442 , \15443_nR84b , \15444 , \15445 , \15446 , \15447 ,
         \15448 , \15449 , \15450 , \15451 , \15452 , \15453 , \15454 , \15455 , \15456 , \15457 ,
         \15458 , \15459 , \15460 , \15461 , \15462 , \15463 , \15464 , \15465 , \15466 , \15467 ,
         \15468 , \15469_nR6ad , \15470 , \15471 , \15472_nR6cb , \15473 , \15474 , \15475 , \15476 , \15477 ,
         \15478 , \15479 , \15480 , \15481 , \15482 , \15483_nR707 , \15484 , \15485 , \15486 , \15487 ,
         \15488 , \15489 , \15490 , \15491_nR725 , \15492 , \15493 , \15494 , \15495 , \15496 , \15497 ,
         \15498 , \15499 , \15500 , \15501 , \15502_nR743 , \15503 , \15504 , \15505 , \15506 , \15507 ,
         \15508 , \15509 , \15510_nR761 , \15511 , \15512 , \15513 , \15514 , \15515 , \15516 , \15517 ,
         \15518_nR77f , \15519 , \15520 , \15521 , \15522 , \15523 , \15524 , \15525 , \15526_nR79d , \15527 ,
         \15528 , \15529_nR7f7 , \15530 , \15531 , \15532_nR815 , \15533 , \15534 , \15535 , \15536 , \15537 ,
         \15538 , \15539 , \15540 , \15541 , \15542 , \15543_nR7d9 , \15544 , \15545 , \15546 , \15547 ,
         \15548 , \15549 , \15550 , \15551 , \15552 , \15553 , \15554 , \15555_nR7bb , \15556 , \15557 ,
         \15558 , \15559 , \15560 , \15561 , \15562 , \15563 , \15564 , \15565 , \15566 , \15567 ,
         \15568 , \15569 , \15570 , \15571 , \15572 , \15573 , \15574 , \15575 , \15576 , \15577 ,
         \15578 , \15579 , \15580 , \15581_nR6e9 , \15582 , \15583 , \15584 , \15585 , \15586 , \15587 ,
         \15588 , \15589 , \15590_nR3dc1 , \15591 , \15592 , \15593 , \15594 , \15595 , \15596 , \15597 ,
         \15598 , \15599 , \15600_nR3d84 , \15601 , \15602 , \15603 , \15604 , \15605 , \15606 , \15607 ,
         \15608 , \15609 , \15610 , \15611_nR3d54 , \15612 , \15613 , \15614 , \15615 , \15616 , \15617_nR3d07 ,
         \15618 , \15619 , \15620 , \15621 , \15622 , \15623_nR3c96 , \15624 , \15625 , \15626 , \15627 ,
         \15628 , \15629_nR3c30 , \15630 , \15631 , \15632 , \15633 , \15634 , \15635_nR3b9b , \15636 , \15637 ,
         \15638 , \15639 , \15640 , \15641_nR3afb , \15642 , \15643 , \15644 , \15645 , \15646 , \15647 ,
         \15648_nR3a4f , \15649 , \15650 , \15651 , \15652 , \15653 , \15654 , \15655 , \15656 , \15657 ,
         \15658 , \15659_nR3999 , \15660 , \15661 , \15662 , \15663 , \15664 , \15665_nR38e8 , \15666 , \15667 ,
         \15668 , \15669 , \15670 , \15671_nR381f , \15672 , \15673 , \15674 , \15675 , \15676 , \15677 ,
         \15678 , \15679 , \15680 , \15681 , \15682_nR374a , \15683 , \15684 , \15685 , \15686 , \15687 ,
         \15688_nR3678 , \15689 , \15690 , \15691 , \15692 , \15693 , \15694_nR3576 , \15695 , \15696 , \15697 ,
         \15698 , \15699 , \15700_nR3464 , \15701 , \15702 , \15703 , \15704 , \15705 , \15706_nR333e , \15707 ,
         \15708 , \15709 , \15710 , \15711 , \15712_nR3236 , \15713 , \15714 , \15715 , \15716 , \15717 ,
         \15718 , \15719 , \15720_nR3115 , \15721 , \15722 , \15723 , \15724 , \15725 , \15726 , \15727 ,
         \15728 , \15729 , \15730 , \15731 , \15732 , \15733 , \15734 , \15735 , \15736_nR2ffe , \15737 ,
         \15738 , \15739 , \15740 , \15741 , \15742_nR2ee6 , \15743 , \15744 , \15745 , \15746 , \15747 ,
         \15748_nR2def , \15749 , \15750 , \15751 , \15752 , \15753 , \15754_nR2cdf , \15755 , \15756 , \15757 ,
         \15758 , \15759 , \15760_nR2c00 , \15761 , \15762 , \15763 , \15764 , \15765 , \15766_nR2af2 , \15767 ,
         \15768 , \15769 , \15770 , \15771 , \15772_nR2a16 , \15773 , \15774 , \15775 , \15776 , \15777 ,
         \15778_nR2937 , \15779 ;
buf \U$labajz1652 ( R_267_b942f48, \7980 );
buf \U$labajz1653 ( R_268_b942ff0, \7990 );
buf \U$labajz1654 ( R_269_b943098, \7997 );
buf \U$labajz1655 ( R_26a_b943140, \8004 );
buf \U$labajz1656 ( R_26b_b9431e8, \8015 );
buf \U$labajz1657 ( R_26c_b943290, \8021 );
buf \U$labajz1658 ( R_26d_b943338, \8027 );
buf \U$labajz1659 ( R_26e_b9433e0, \8038 );
buf \U$labajz1660 ( R_26f_b943488, \8053 );
buf \U$labajz1661 ( R_270_b943530, \8062 );
buf \U$labajz1662 ( R_271_b9435d8, \8072 );
buf \U$labajz1663 ( R_272_b943680, \8089 );
buf \U$labajz1664 ( R_273_b943728, \8103 );
buf \U$labajz1665 ( R_274_b9437d0, \8114 );
buf \U$labajz1666 ( R_275_b943878, \8120 );
buf \U$labajz1667 ( R_276_b943920, \8126 );
buf \U$labajz1668 ( R_277_b9439c8, \8132 );
buf \U$labajz1669 ( R_278_b943a70, \8142 );
buf \U$labajz1670 ( R_279_b943b18, \8154 );
buf \U$labajz1671 ( R_27a_b943bc0, \8170 );
buf \U$labajz1672 ( R_27b_b943c68, \8176 );
buf \U$labajz1673 ( R_27c_b943d10, \8182 );
buf \U$labajz1674 ( R_27d_b943db8, \8188 );
buf \U$labajz1675 ( R_27e_b943e60, \8194 );
buf \U$labajz1676 ( R_27f_b943f08, \8200 );
buf \U$labajz1677 ( R_280_b943fb0, \8206 );
buf \U$labajz1678 ( R_281_b944058, \8212 );
buf \U$labajz1679 ( R_289_b944598, \15591 );
buf \U$labajz1680 ( R_28a_b944640, \15601 );
buf \U$labajz1681 ( R_28b_b9446e8, \15612 );
buf \U$labajz1682 ( R_28c_b944790, \15618 );
buf \U$labajz1683 ( R_28d_b944838, \15624 );
buf \U$labajz1684 ( R_28e_b9448e0, \15630 );
buf \U$labajz1685 ( R_28f_b944988, \15636 );
buf \U$labajz1686 ( R_290_b944a30, \15642 );
buf \U$labajz1687 ( R_291_b944ad8, \15649 );
buf \U$labajz1688 ( R_292_b944b80, \15660 );
buf \U$labajz1689 ( R_293_b944c28, \15666 );
buf \U$labajz1690 ( R_294_b944cd0, \15672 );
buf \U$labajz1691 ( R_295_b944d78, \15683 );
buf \U$labajz1692 ( R_296_b944e20, \15689 );
buf \U$labajz1693 ( R_297_b944ec8, \15695 );
buf \U$labajz1694 ( R_298_b944f70, \15701 );
buf \U$labajz1695 ( R_299_b945018, \15707 );
buf \U$labajz1696 ( R_29a_b9450c0, \15713 );
buf \U$labajz1697 ( R_29b_b945168, \15721 );
buf \U$labajz1698 ( R_29c_b945210, \15737 );
buf \U$labajz1699 ( R_29d_b9452b8, \15743 );
buf \U$labajz1700 ( R_29e_b945360, \15749 );
buf \U$labajz1701 ( R_29f_b945408, \15755 );
buf \U$labajz1702 ( R_2a0_b9454b0, \15761 );
buf \U$labajz1703 ( R_2a1_b945558, \15767 );
buf \U$labajz1704 ( R_2a2_b945600, \15773 );
buf \U$labajz1705 ( R_2a3_b9456a8, \15779 );
nand \U$1 ( \671 , RIb54a900_11, RIb54a888_10);
not \U$2 ( \672 , \671 );
nand \U$3 ( \673 , \672 , RIb54a810_9);
not \U$4 ( \674 , \673 );
nand \U$5 ( \675 , \674 , RIb54a798_8);
not \U$6 ( \676 , \675 );
nand \U$7 ( \677 , \676 , RIb54a720_7);
not \U$8 ( \678 , \677 );
nand \U$9 ( \679 , \678 , RIb54a6a8_6);
not \U$10 ( \680 , \679 );
nand \U$11 ( \681 , \680 , RIb54a630_5);
not \U$12 ( \682 , \681 );
nand \U$13 ( \683 , \682 , RIb54a5b8_4);
not \U$14 ( \684 , \683 );
nand \U$15 ( \685 , \684 , RIb54a540_3);
not \U$16 ( \686 , \685 );
nand \U$17 ( \687 , \686 , RIb54a4c8_2);
not \U$18 ( \688 , \687 );
nand \U$19 ( \689 , \688 , RIb54a450_1);
not \U$20 ( \690 , \689 );
not \U$21 ( \691 , RIb5517a0_247);
and \U$22 ( \692 , \690 , \691 );
and \U$23 ( \693 , \689 , RIb5517a0_247);
nor \U$24 ( \694 , \692 , \693 );
not \U$25 ( \695 , RIb54abd0_17);
nand \U$26 ( \696 , RIb54ab58_16, \695 );
not \U$27 ( \697 , \696 );
nand \U$28 ( \698 , \697 , RIb54aae0_15);
not \U$29 ( \699 , RIb54aa68_14);
nand \U$30 ( \700 , \699 , RIb54a9f0_13);
nor \U$31 ( \701 , \698 , \700 );
and \U$32 ( \702 , RIb551980_251, \701 );
not \U$33 ( \703 , RIb54a9f0_13);
nand \U$34 ( \704 , RIb54aa68_14, \703 );
nor \U$35 ( \705 , \698 , \704 );
and \U$36 ( \706 , RIb551908_250, \705 );
not \U$37 ( \707 , \696 );
not \U$38 ( \708 , RIb54aae0_15);
nand \U$39 ( \709 , \707 , \708 );
nor \U$40 ( \710 , \709 , \700 );
and \U$41 ( \711 , RIb551b60_255, \710 );
nor \U$42 ( \712 , \709 , \704 );
and \U$43 ( \713 , RIb551ae8_254, \712 );
nor \U$44 ( \714 , RIb54a9f0_13, RIb54aa68_14);
not \U$45 ( \715 , \714 );
nor \U$46 ( \716 , \715 , RIb54aae0_15);
nor \U$47 ( \717 , RIb54ab58_16, RIb54abd0_17);
and \U$48 ( \718 , \716 , \717 );
and \U$49 ( \719 , \718 , RIb551f98_264);
nand \U$50 ( \720 , \708 , \717 );
nor \U$51 ( \721 , \720 , \700 );
and \U$52 ( \722 , RIb551f20_263, \721 );
nor \U$53 ( \723 , \719 , \722 );
not \U$54 ( \724 , \723 );
nor \U$55 ( \725 , \711 , \713 , \724 );
nand \U$56 ( \726 , RIb54aae0_15, \717 );
nor \U$57 ( \727 , \726 , \704 );
and \U$58 ( \728 , \727 , RIb551cc8_258);
nand \U$59 ( \729 , RIb54aa68_14, RIb54a9f0_13);
nor \U$60 ( \730 , \729 , \708 );
and \U$61 ( \731 , \730 , \717 );
and \U$62 ( \732 , RIb551c50_257, \731 );
nor \U$63 ( \733 , \728 , \732 );
not \U$64 ( \734 , \716 );
nor \U$65 ( \735 , \734 , \696 );
and \U$66 ( \736 , \735 , RIb551bd8_256);
not \U$67 ( \737 , \730 );
nor \U$68 ( \738 , \737 , \696 );
and \U$69 ( \739 , RIb551890_249, \738 );
nor \U$70 ( \740 , \736 , \739 );
not \U$71 ( \741 , RIb54ab58_16);
nand \U$72 ( \742 , \741 , \716 );
nor \U$73 ( \743 , \742 , \695 );
nand \U$74 ( \744 , RIb551818_248, \743 );
nand \U$75 ( \745 , \725 , \733 , \740 , \744 );
nor \U$76 ( \746 , \702 , \706 , \745 );
nor \U$77 ( \747 , \720 , \704 );
and \U$78 ( \748 , \747 , RIb551ea8_262);
nor \U$79 ( \749 , \720 , \729 );
and \U$80 ( \750 , RIb551e30_261, \749 );
nor \U$81 ( \751 , \748 , \750 );
not \U$82 ( \752 , \714 );
nor \U$83 ( \753 , \752 , \726 );
and \U$84 ( \754 , \753 , RIb551db8_260);
nor \U$85 ( \755 , \726 , \700 );
and \U$86 ( \756 , RIb551d40_259, \755 );
nor \U$87 ( \757 , \754 , \756 );
not \U$88 ( \758 , \714 );
nor \U$89 ( \759 , \758 , \698 );
and \U$90 ( \760 , \759 , RIb5519f8_252);
nor \U$91 ( \761 , \709 , \729 );
and \U$92 ( \762 , RIb551a70_253, \761 );
nor \U$93 ( \763 , \760 , \762 );
nand \U$94 ( \764 , \746 , \751 , \757 , \763 );
buf \U$95 ( \765 , \764 );
and \U$96 ( \766 , \742 , RIb54abd0_17);
buf \U$97 ( \767 , \766 );
_DC r12c0 ( \768_nR12c0 , \765 , \767 );
xor \U$98 ( \769 , \694 , \768_nR12c0 );
not \U$99 ( \770 , \687 );
not \U$100 ( \771 , RIb54a450_1);
and \U$101 ( \772 , \770 , \771 );
and \U$102 ( \773 , \687 , RIb54a450_1);
nor \U$103 ( \774 , \772 , \773 );
and \U$104 ( \775 , RIb54ad38_20, \701 );
and \U$105 ( \776 , RIb54acc0_19, \705 );
and \U$106 ( \777 , RIb54af18_24, \710 );
and \U$107 ( \778 , RIb54aea0_23, \712 );
and \U$108 ( \779 , \718 , RIb54b350_33);
and \U$109 ( \780 , RIb54b2d8_32, \721 );
nor \U$110 ( \781 , \779 , \780 );
not \U$111 ( \782 , \781 );
nor \U$112 ( \783 , \777 , \778 , \782 );
and \U$113 ( \784 , \735 , RIb54af90_25);
and \U$114 ( \785 , RIb54b008_26, \731 );
nor \U$115 ( \786 , \784 , \785 );
and \U$116 ( \787 , \727 , RIb54b080_27);
and \U$117 ( \788 , RIb54ac48_18, \738 );
nor \U$118 ( \789 , \787 , \788 );
nand \U$119 ( \790 , RIb54a978_12, \743 );
nand \U$120 ( \791 , \783 , \786 , \789 , \790 );
nor \U$121 ( \792 , \775 , \776 , \791 );
and \U$122 ( \793 , \747 , RIb54b260_31);
and \U$123 ( \794 , RIb54b1e8_30, \749 );
nor \U$124 ( \795 , \793 , \794 );
and \U$125 ( \796 , \753 , RIb54b170_29);
and \U$126 ( \797 , RIb54b0f8_28, \755 );
nor \U$127 ( \798 , \796 , \797 );
and \U$128 ( \799 , \759 , RIb54adb0_21);
and \U$129 ( \800 , RIb54ae28_22, \761 );
nor \U$130 ( \801 , \799 , \800 );
nand \U$131 ( \802 , \792 , \795 , \798 , \801 );
buf \U$132 ( \803 , \802 );
_DC r10db ( \804_nR10db , \803 , \767 );
xor \U$133 ( \805 , \774 , \804_nR10db );
not \U$134 ( \806 , \685 );
not \U$135 ( \807 , RIb54a4c8_2);
and \U$136 ( \808 , \806 , \807 );
and \U$137 ( \809 , \685 , RIb54a4c8_2);
nor \U$138 ( \810 , \808 , \809 );
and \U$139 ( \811 , RIb54b968_46, \753 );
and \U$140 ( \812 , RIb54b8f0_45, \755 );
and \U$141 ( \813 , RIb54b710_41, \710 );
and \U$142 ( \814 , RIb54b698_40, \712 );
and \U$143 ( \815 , \718 , RIb54bb48_50);
and \U$144 ( \816 , RIb54bad0_49, \721 );
nor \U$145 ( \817 , \815 , \816 );
not \U$146 ( \818 , \817 );
nor \U$147 ( \819 , \813 , \814 , \818 );
and \U$148 ( \820 , \735 , RIb54b788_42);
and \U$149 ( \821 , RIb54b620_39, \761 );
nor \U$150 ( \822 , \820 , \821 );
and \U$151 ( \823 , \727 , RIb54b878_44);
and \U$152 ( \824 , RIb54b800_43, \731 );
nor \U$153 ( \825 , \823 , \824 );
nand \U$154 ( \826 , RIb54b3c8_34, \743 );
nand \U$155 ( \827 , \819 , \822 , \825 , \826 );
nor \U$156 ( \828 , \811 , \812 , \827 );
and \U$157 ( \829 , \705 , RIb54b4b8_36);
and \U$158 ( \830 , RIb54b440_35, \738 );
nor \U$159 ( \831 , \829 , \830 );
and \U$160 ( \832 , \747 , RIb54ba58_48);
and \U$161 ( \833 , RIb54b9e0_47, \749 );
nor \U$162 ( \834 , \832 , \833 );
and \U$163 ( \835 , \759 , RIb54b5a8_38);
and \U$164 ( \836 , RIb54b530_37, \701 );
nor \U$165 ( \837 , \835 , \836 );
nand \U$166 ( \838 , \828 , \831 , \834 , \837 );
buf \U$167 ( \839 , \838 );
_DC r10d9 ( \840_nR10d9 , \839 , \767 );
xor \U$168 ( \841 , \810 , \840_nR10d9 );
not \U$169 ( \842 , \683 );
not \U$170 ( \843 , RIb54a540_3);
and \U$171 ( \844 , \842 , \843 );
and \U$172 ( \845 , \683 , RIb54a540_3);
nor \U$173 ( \846 , \844 , \845 );
and \U$174 ( \847 , RIb54bf08_58, \710 );
and \U$175 ( \848 , RIb54be90_57, \712 );
and \U$176 ( \849 , RIb54c160_63, \753 );
and \U$177 ( \850 , RIb54bda0_55, \759 );
and \U$178 ( \851 , \701 , RIb54bd28_54);
and \U$179 ( \852 , RIb54bc38_52, \738 );
nor \U$180 ( \853 , \851 , \852 );
not \U$181 ( \854 , \853 );
nor \U$182 ( \855 , \849 , \850 , \854 );
and \U$183 ( \856 , \761 , RIb54be18_56);
and \U$184 ( \857 , RIb54bcb0_53, \705 );
nor \U$185 ( \858 , \856 , \857 );
and \U$186 ( \859 , \718 , RIb54c340_67);
and \U$187 ( \860 , RIb54c0e8_62, \755 );
nor \U$188 ( \861 , \859 , \860 );
nand \U$189 ( \862 , RIb54bbc0_51, \743 );
nand \U$190 ( \863 , \855 , \858 , \861 , \862 );
nor \U$191 ( \864 , \847 , \848 , \863 );
and \U$192 ( \865 , \747 , RIb54c250_65);
and \U$193 ( \866 , RIb54c1d8_64, \749 );
nor \U$194 ( \867 , \865 , \866 );
and \U$195 ( \868 , \727 , RIb54c070_61);
and \U$196 ( \869 , RIb54bff8_60, \731 );
nor \U$197 ( \870 , \868 , \869 );
and \U$198 ( \871 , \721 , RIb54c2c8_66);
and \U$199 ( \872 , RIb54bf80_59, \735 );
nor \U$200 ( \873 , \871 , \872 );
nand \U$201 ( \874 , \864 , \867 , \870 , \873 );
buf \U$202 ( \875 , \874 );
_DC rf20 ( \876_nRf20 , \875 , \767 );
xor \U$203 ( \877 , \846 , \876_nRf20 );
not \U$204 ( \878 , \681 );
not \U$205 ( \879 , RIb54a5b8_4);
and \U$206 ( \880 , \878 , \879 );
and \U$207 ( \881 , \681 , RIb54a5b8_4);
nor \U$208 ( \882 , \880 , \881 );
and \U$209 ( \883 , RIb54c8e0_79, \755 );
and \U$210 ( \884 , RIb54c700_75, \710 );
and \U$211 ( \885 , RIb54c778_76, \735 );
and \U$212 ( \886 , RIb54c610_73, \761 );
and \U$213 ( \887 , \701 , RIb54c520_71);
and \U$214 ( \888 , RIb54c430_69, \738 );
nor \U$215 ( \889 , \887 , \888 );
not \U$216 ( \890 , \889 );
nor \U$217 ( \891 , \885 , \886 , \890 );
and \U$218 ( \892 , \759 , RIb54c598_72);
and \U$219 ( \893 , RIb54c4a8_70, \705 );
nor \U$220 ( \894 , \892 , \893 );
and \U$221 ( \895 , \727 , RIb54c868_78);
and \U$222 ( \896 , RIb54c7f0_77, \731 );
nor \U$223 ( \897 , \895 , \896 );
nand \U$224 ( \898 , RIb54c3b8_68, \743 );
nand \U$225 ( \899 , \891 , \894 , \897 , \898 );
nor \U$226 ( \900 , \883 , \884 , \899 );
and \U$227 ( \901 , \718 , RIb54cb38_84);
and \U$228 ( \902 , RIb54cac0_83, \721 );
nor \U$229 ( \903 , \901 , \902 );
and \U$230 ( \904 , \747 , RIb54ca48_82);
and \U$231 ( \905 , RIb54c9d0_81, \749 );
nor \U$232 ( \906 , \904 , \905 );
and \U$233 ( \907 , \753 , RIb54c958_80);
and \U$234 ( \908 , RIb54c688_74, \712 );
nor \U$235 ( \909 , \907 , \908 );
nand \U$236 ( \910 , \900 , \903 , \906 , \909 );
buf \U$237 ( \911 , \910 );
_DC rf1e ( \912_nRf1e , \911 , \767 );
xor \U$238 ( \913 , \882 , \912_nRf1e );
not \U$239 ( \914 , \679 );
not \U$240 ( \915 , RIb54a630_5);
and \U$241 ( \916 , \914 , \915 );
and \U$242 ( \917 , \679 , RIb54a630_5);
nor \U$243 ( \918 , \916 , \917 );
and \U$244 ( \919 , RIb54cca0_87, \705 );
and \U$245 ( \920 , RIb54cc28_86, \738 );
and \U$246 ( \921 , RIb54cef8_92, \710 );
and \U$247 ( \922 , RIb54ce80_91, \712 );
and \U$248 ( \923 , \759 , RIb54cd90_89);
and \U$249 ( \924 , RIb54cfe8_94, \731 );
nor \U$250 ( \925 , \923 , \924 );
not \U$251 ( \926 , \925 );
nor \U$252 ( \927 , \921 , \922 , \926 );
and \U$253 ( \928 , \747 , RIb54d240_99);
and \U$254 ( \929 , RIb54ce08_90, \761 );
nor \U$255 ( \930 , \928 , \929 );
and \U$256 ( \931 , \718 , RIb54d330_101);
and \U$257 ( \932 , RIb54d2b8_100, \721 );
nor \U$258 ( \933 , \931 , \932 );
nand \U$259 ( \934 , RIb54cbb0_85, \743 );
nand \U$260 ( \935 , \927 , \930 , \933 , \934 );
nor \U$261 ( \936 , \919 , \920 , \935 );
and \U$262 ( \937 , \753 , RIb54d150_97);
and \U$263 ( \938 , RIb54d1c8_98, \749 );
nor \U$264 ( \939 , \937 , \938 );
and \U$265 ( \940 , \755 , RIb54d0d8_96);
and \U$266 ( \941 , RIb54d060_95, \727 );
nor \U$267 ( \942 , \940 , \941 );
and \U$268 ( \943 , \735 , RIb54cf70_93);
and \U$269 ( \944 , RIb54cd18_88, \701 );
nor \U$270 ( \945 , \943 , \944 );
nand \U$271 ( \946 , \936 , \939 , \942 , \945 );
buf \U$272 ( \947 , \946 );
_DC rda0 ( \948_nRda0 , \947 , \767 );
xor \U$273 ( \949 , \918 , \948_nRda0 );
not \U$274 ( \950 , \677 );
not \U$275 ( \951 , RIb54a6a8_6);
and \U$276 ( \952 , \950 , \951 );
and \U$277 ( \953 , \677 , RIb54a6a8_6);
nor \U$278 ( \954 , \952 , \953 );
and \U$279 ( \955 , RIb54d498_104, \705 );
and \U$280 ( \956 , RIb54d420_103, \738 );
and \U$281 ( \957 , RIb54d6f0_109, \710 );
and \U$282 ( \958 , RIb54d678_108, \712 );
and \U$283 ( \959 , \718 , RIb54db28_118);
and \U$284 ( \960 , RIb54dab0_117, \721 );
nor \U$285 ( \961 , \959 , \960 );
not \U$286 ( \962 , \961 );
nor \U$287 ( \963 , \957 , \958 , \962 );
and \U$288 ( \964 , \735 , RIb54d768_110);
and \U$289 ( \965 , RIb54d510_105, \701 );
nor \U$290 ( \966 , \964 , \965 );
and \U$291 ( \967 , \727 , RIb54d858_112);
and \U$292 ( \968 , RIb54d7e0_111, \731 );
nor \U$293 ( \969 , \967 , \968 );
nand \U$294 ( \970 , RIb54d3a8_102, \743 );
nand \U$295 ( \971 , \963 , \966 , \969 , \970 );
nor \U$296 ( \972 , \955 , \956 , \971 );
and \U$297 ( \973 , \747 , RIb54da38_116);
and \U$298 ( \974 , RIb54d9c0_115, \749 );
nor \U$299 ( \975 , \973 , \974 );
and \U$300 ( \976 , \753 , RIb54d948_114);
and \U$301 ( \977 , RIb54d8d0_113, \755 );
nor \U$302 ( \978 , \976 , \977 );
and \U$303 ( \979 , \759 , RIb54d588_106);
and \U$304 ( \980 , RIb54d600_107, \761 );
nor \U$305 ( \981 , \979 , \980 );
nand \U$306 ( \982 , \972 , \975 , \978 , \981 );
buf \U$307 ( \983 , \982 );
_DC rd9e ( \984_nRd9e , \983 , \767 );
xor \U$308 ( \985 , \954 , \984_nRd9e );
not \U$309 ( \986 , \675 );
not \U$310 ( \987 , RIb54a720_7);
and \U$311 ( \988 , \986 , \987 );
and \U$312 ( \989 , \675 , RIb54a720_7);
nor \U$313 ( \990 , \988 , \989 );
and \U$314 ( \991 , RIb54dee8_126, \710 );
and \U$315 ( \992 , RIb54de70_125, \712 );
and \U$316 ( \993 , RIb54e050_129, \727 );
and \U$317 ( \994 , RIb54dfd8_128, \731 );
and \U$318 ( \995 , \753 , RIb54e140_131);
and \U$319 ( \996 , RIb54e0c8_130, \755 );
nor \U$320 ( \997 , \995 , \996 );
not \U$321 ( \998 , \997 );
nor \U$322 ( \999 , \993 , \994 , \998 );
and \U$323 ( \1000 , \735 , RIb54df60_127);
and \U$324 ( \1001 , RIb54dd08_122, \701 );
nor \U$325 ( \1002 , \1000 , \1001 );
and \U$326 ( \1003 , \747 , RIb54e230_133);
and \U$327 ( \1004 , RIb54e1b8_132, \749 );
nor \U$328 ( \1005 , \1003 , \1004 );
nand \U$329 ( \1006 , RIb54dba0_119, \743 );
nand \U$330 ( \1007 , \999 , \1002 , \1005 , \1006 );
nor \U$331 ( \1008 , \991 , \992 , \1007 );
and \U$332 ( \1009 , \705 , RIb54dc90_121);
and \U$333 ( \1010 , RIb54dc18_120, \738 );
nor \U$334 ( \1011 , \1009 , \1010 );
and \U$335 ( \1012 , \718 , RIb54e320_135);
and \U$336 ( \1013 , RIb54e2a8_134, \721 );
nor \U$337 ( \1014 , \1012 , \1013 );
and \U$338 ( \1015 , \759 , RIb54dd80_123);
and \U$339 ( \1016 , RIb54ddf8_124, \761 );
nor \U$340 ( \1017 , \1015 , \1016 );
nand \U$341 ( \1018 , \1008 , \1011 , \1014 , \1017 );
buf \U$342 ( \1019 , \1018 );
_DC rc66 ( \1020_nRc66 , \1019 , \767 );
xor \U$343 ( \1021 , \990 , \1020_nRc66 );
not \U$344 ( \1022 , \673 );
not \U$345 ( \1023 , RIb54a798_8);
and \U$346 ( \1024 , \1022 , \1023 );
and \U$347 ( \1025 , \673 , RIb54a798_8);
nor \U$348 ( \1026 , \1024 , \1025 );
and \U$349 ( \1027 , RIb54e500_139, \701 );
and \U$350 ( \1028 , RIb54e488_138, \705 );
and \U$351 ( \1029 , RIb54e6e0_143, \710 );
and \U$352 ( \1030 , RIb54e668_142, \712 );
and \U$353 ( \1031 , \718 , RIb54eb18_152);
and \U$354 ( \1032 , RIb54eaa0_151, \721 );
nor \U$355 ( \1033 , \1031 , \1032 );
not \U$356 ( \1034 , \1033 );
nor \U$357 ( \1035 , \1029 , \1030 , \1034 );
and \U$358 ( \1036 , \735 , RIb54e758_144);
and \U$359 ( \1037 , RIb54e7d0_145, \731 );
nor \U$360 ( \1038 , \1036 , \1037 );
and \U$361 ( \1039 , \727 , RIb54e848_146);
and \U$362 ( \1040 , RIb54e410_137, \738 );
nor \U$363 ( \1041 , \1039 , \1040 );
nand \U$364 ( \1042 , RIb54e398_136, \743 );
nand \U$365 ( \1043 , \1035 , \1038 , \1041 , \1042 );
nor \U$366 ( \1044 , \1027 , \1028 , \1043 );
and \U$367 ( \1045 , \747 , RIb54ea28_150);
and \U$368 ( \1046 , RIb54e9b0_149, \749 );
nor \U$369 ( \1047 , \1045 , \1046 );
and \U$370 ( \1048 , \753 , RIb54e938_148);
and \U$371 ( \1049 , RIb54e8c0_147, \755 );
nor \U$372 ( \1050 , \1048 , \1049 );
and \U$373 ( \1051 , \759 , RIb54e578_140);
and \U$374 ( \1052 , RIb54e5f0_141, \761 );
nor \U$375 ( \1053 , \1051 , \1052 );
nand \U$376 ( \1054 , \1044 , \1047 , \1050 , \1053 );
buf \U$377 ( \1055 , \1054 );
_DC rc64 ( \1056_nRc64 , \1055 , \767 );
xor \U$378 ( \1057 , \1026 , \1056_nRc64 );
not \U$379 ( \1058 , \671 );
not \U$380 ( \1059 , RIb54a810_9);
and \U$381 ( \1060 , \1058 , \1059 );
and \U$382 ( \1061 , \671 , RIb54a810_9);
nor \U$383 ( \1062 , \1060 , \1061 );
and \U$384 ( \1063 , RIb54eed8_160, \710 );
and \U$385 ( \1064 , RIb54ee60_159, \712 );
and \U$386 ( \1065 , RIb54f040_163, \727 );
and \U$387 ( \1066 , RIb54efc8_162, \731 );
and \U$388 ( \1067 , \747 , RIb54f220_167);
and \U$389 ( \1068 , RIb54f1a8_166, \749 );
nor \U$390 ( \1069 , \1067 , \1068 );
not \U$391 ( \1070 , \1069 );
nor \U$392 ( \1071 , \1065 , \1066 , \1070 );
and \U$393 ( \1072 , \735 , RIb54ef50_161);
and \U$394 ( \1073 , RIb54ede8_158, \761 );
nor \U$395 ( \1074 , \1072 , \1073 );
and \U$396 ( \1075 , \753 , RIb54f130_165);
and \U$397 ( \1076 , RIb54f0b8_164, \755 );
nor \U$398 ( \1077 , \1075 , \1076 );
nand \U$399 ( \1078 , RIb54eb90_153, \743 );
nand \U$400 ( \1079 , \1071 , \1074 , \1077 , \1078 );
nor \U$401 ( \1080 , \1063 , \1064 , \1079 );
and \U$402 ( \1081 , \705 , RIb54ec80_155);
and \U$403 ( \1082 , RIb54ec08_154, \738 );
nor \U$404 ( \1083 , \1081 , \1082 );
and \U$405 ( \1084 , \718 , RIb54f310_169);
and \U$406 ( \1085 , RIb54f298_168, \721 );
nor \U$407 ( \1086 , \1084 , \1085 );
and \U$408 ( \1087 , \759 , RIb54ed70_157);
and \U$409 ( \1088 , RIb54ecf8_156, \701 );
nor \U$410 ( \1089 , \1087 , \1088 );
nand \U$411 ( \1090 , \1080 , \1083 , \1086 , \1089 );
buf \U$412 ( \1091 , \1090 );
_DC rb7a ( \1092_nRb7a , \1091 , \767 );
xor \U$413 ( \1093 , \1062 , \1092_nRb7a );
not \U$414 ( \1094 , RIb54a900_11);
and \U$415 ( \1095 , RIb54a888_10, \1094 );
not \U$416 ( \1096 , RIb54a888_10);
and \U$417 ( \1097 , \1096 , RIb54a900_11);
nor \U$418 ( \1098 , \1095 , \1097 );
and \U$419 ( \1099 , RIb54f6d0_177, \710 );
and \U$420 ( \1100 , RIb54f658_176, \712 );
and \U$421 ( \1101 , RIb54f838_180, \727 );
and \U$422 ( \1102 , RIb54f7c0_179, \731 );
and \U$423 ( \1103 , \705 , RIb54f478_172);
and \U$424 ( \1104 , RIb54f400_171, \738 );
nor \U$425 ( \1105 , \1103 , \1104 );
not \U$426 ( \1106 , \1105 );
nor \U$427 ( \1107 , \1101 , \1102 , \1106 );
and \U$428 ( \1108 , \747 , RIb54fa18_184);
and \U$429 ( \1109 , RIb54f9a0_183, \749 );
nor \U$430 ( \1110 , \1108 , \1109 );
and \U$431 ( \1111 , \753 , RIb54f928_182);
and \U$432 ( \1112 , RIb54f8b0_181, \755 );
nor \U$433 ( \1113 , \1111 , \1112 );
nand \U$434 ( \1114 , RIb54f388_170, \743 );
nand \U$435 ( \1115 , \1107 , \1110 , \1113 , \1114 );
nor \U$436 ( \1116 , \1099 , \1100 , \1115 );
and \U$437 ( \1117 , \735 , RIb54f748_178);
and \U$438 ( \1118 , RIb54f5e0_175, \761 );
nor \U$439 ( \1119 , \1117 , \1118 );
and \U$440 ( \1120 , \718 , RIb54fb08_186);
and \U$441 ( \1121 , RIb54fa90_185, \721 );
nor \U$442 ( \1122 , \1120 , \1121 );
and \U$443 ( \1123 , \759 , RIb54f568_174);
and \U$444 ( \1124 , RIb54f4f0_173, \701 );
nor \U$445 ( \1125 , \1123 , \1124 );
nand \U$446 ( \1126 , \1116 , \1119 , \1122 , \1125 );
buf \U$447 ( \1127 , \1126 );
_DC rb7c ( \1128_nRb7c , \1127 , \767 );
xor \U$448 ( \1129 , \1098 , \1128_nRb7c );
and \U$449 ( \1130 , RIb54ff40_195, \735 );
and \U$450 ( \1131 , RIb54fdd8_192, \761 );
and \U$451 ( \1132 , RIb54fc70_189, \705 );
and \U$452 ( \1133 , RIb54fbf8_188, \738 );
and \U$453 ( \1134 , \718 , RIb550300_203);
and \U$454 ( \1135 , RIb550288_202, \721 );
nor \U$455 ( \1136 , \1134 , \1135 );
not \U$456 ( \1137 , \1136 );
nor \U$457 ( \1138 , \1132 , \1133 , \1137 );
and \U$458 ( \1139 , \759 , RIb54fd60_191);
and \U$459 ( \1140 , RIb54fce8_190, \701 );
nor \U$460 ( \1141 , \1139 , \1140 );
and \U$461 ( \1142 , \710 , RIb54fec8_194);
and \U$462 ( \1143 , RIb54fe50_193, \712 );
nor \U$463 ( \1144 , \1142 , \1143 );
nand \U$464 ( \1145 , RIb54fb80_187, \743 );
nand \U$465 ( \1146 , \1138 , \1141 , \1144 , \1145 );
nor \U$466 ( \1147 , \1130 , \1131 , \1146 );
and \U$467 ( \1148 , \753 , RIb550120_199);
and \U$468 ( \1149 , RIb5500a8_198, \755 );
nor \U$469 ( \1150 , \1148 , \1149 );
and \U$470 ( \1151 , \727 , RIb550030_197);
and \U$471 ( \1152 , RIb54ffb8_196, \731 );
nor \U$472 ( \1153 , \1151 , \1152 );
and \U$473 ( \1154 , \747 , RIb550210_201);
and \U$474 ( \1155 , RIb550198_200, \749 );
nor \U$475 ( \1156 , \1154 , \1155 );
nand \U$476 ( \1157 , \1147 , \1150 , \1153 , \1156 );
buf \U$477 ( \1158 , \1157 );
_DC r9e7 ( \1159_nR9e7 , \1158 , \767 );
xor \U$478 ( \1160 , RIb54a900_11, \1159_nR9e7 );
and \U$479 ( \1161 , RIb550990_217, \753 );
and \U$480 ( \1162 , RIb550918_216, \755 );
and \U$481 ( \1163 , RIb550738_212, \710 );
and \U$482 ( \1164 , RIb5506c0_211, \712 );
and \U$483 ( \1165 , \718 , RIb550b70_221);
and \U$484 ( \1166 , RIb550af8_220, \721 );
nor \U$485 ( \1167 , \1165 , \1166 );
not \U$486 ( \1168 , \1167 );
nor \U$487 ( \1169 , \1163 , \1164 , \1168 );
and \U$488 ( \1170 , \759 , RIb5505d0_209);
and \U$489 ( \1171 , RIb550558_208, \701 );
nor \U$490 ( \1172 , \1170 , \1171 );
and \U$491 ( \1173 , \705 , RIb5504e0_207);
and \U$492 ( \1174 , RIb550468_206, \738 );
nor \U$493 ( \1175 , \1173 , \1174 );
nand \U$494 ( \1176 , RIb5503f0_205, \743 );
nand \U$495 ( \1177 , \1169 , \1172 , \1175 , \1176 );
nor \U$496 ( \1178 , \1161 , \1162 , \1177 );
and \U$497 ( \1179 , \747 , RIb550a80_219);
and \U$498 ( \1180 , RIb550a08_218, \749 );
nor \U$499 ( \1181 , \1179 , \1180 );
and \U$500 ( \1182 , \727 , RIb5508a0_215);
and \U$501 ( \1183 , RIb550828_214, \731 );
nor \U$502 ( \1184 , \1182 , \1183 );
and \U$503 ( \1185 , \735 , RIb5507b0_213);
and \U$504 ( \1186 , RIb550648_210, \761 );
nor \U$505 ( \1187 , \1185 , \1186 );
nand \U$506 ( \1188 , \1178 , \1181 , \1184 , \1187 );
buf \U$507 ( \1189 , \1188 );
_DC r9e5 ( \1190_nR9e5 , \1189 , \767 );
not \U$508 ( \1191 , RIb550378_204);
nand \U$509 ( \1192 , \1190_nR9e5 , \1191 );
not \U$510 ( \1193 , \1192 );
and \U$511 ( \1194 , \1160 , \1193 );
and \U$512 ( \1195 , RIb54a900_11, \1159_nR9e7 );
or \U$513 ( \1196 , \1194 , \1195 );
and \U$514 ( \1197 , \1129 , \1196 );
and \U$515 ( \1198 , \1098 , \1128_nRb7c );
or \U$516 ( \1199 , \1197 , \1198 );
and \U$517 ( \1200 , \1093 , \1199 );
and \U$518 ( \1201 , \1062 , \1092_nRb7a );
or \U$519 ( \1202 , \1200 , \1201 );
and \U$520 ( \1203 , \1057 , \1202 );
and \U$521 ( \1204 , \1026 , \1056_nRc64 );
or \U$522 ( \1205 , \1203 , \1204 );
and \U$523 ( \1206 , \1021 , \1205 );
and \U$524 ( \1207 , \990 , \1020_nRc66 );
or \U$525 ( \1208 , \1206 , \1207 );
and \U$526 ( \1209 , \985 , \1208 );
and \U$527 ( \1210 , \954 , \984_nRd9e );
or \U$528 ( \1211 , \1209 , \1210 );
and \U$529 ( \1212 , \949 , \1211 );
and \U$530 ( \1213 , \918 , \948_nRda0 );
or \U$531 ( \1214 , \1212 , \1213 );
and \U$532 ( \1215 , \913 , \1214 );
and \U$533 ( \1216 , \882 , \912_nRf1e );
or \U$534 ( \1217 , \1215 , \1216 );
and \U$535 ( \1218 , \877 , \1217 );
and \U$536 ( \1219 , \846 , \876_nRf20 );
or \U$537 ( \1220 , \1218 , \1219 );
and \U$538 ( \1221 , \841 , \1220 );
and \U$539 ( \1222 , \810 , \840_nR10d9 );
or \U$540 ( \1223 , \1221 , \1222 );
and \U$541 ( \1224 , \805 , \1223 );
and \U$542 ( \1225 , \774 , \804_nR10db );
or \U$543 ( \1226 , \1224 , \1225 );
and \U$544 ( \1227 , \769 , \1226 );
and \U$545 ( \1228 , \694 , \768_nR12c0 );
or \U$546 ( \1229 , \1227 , \1228 );
not \U$547 ( \1230 , \689 );
nand \U$548 ( \1231 , \1230 , RIb5517a0_247);
nor \U$549 ( \1232 , \1229 , \1231 );
not \U$550 ( \1233 , \1232 );
and \U$551 ( \1234 , \730 , RIb54ab58_16);
nor \U$552 ( \1235 , RIb550e40_227, RIb550eb8_228, RIb550f30_229, RIb550fa8_230);
nor \U$553 ( \1236 , RIb550c60_223, RIb550cd8_224, RIb550d50_225, RIb550dc8_226);
nand \U$554 ( \1237 , \1235 , \1236 , \695 );
nor \U$555 ( \1238 , \1234 , \1237 );
and \U$556 ( \1239 , \1238 , \730 );
not \U$557 ( \1240 , \1237 );
nand \U$558 ( \1241 , \730 , \1240 );
and \U$559 ( \1242 , RIb54ab58_16, \1241 );
nor \U$560 ( \1243 , \1239 , \1242 );
not \U$561 ( \1244 , \729 );
nand \U$562 ( \1245 , \1244 , \1240 );
and \U$563 ( \1246 , \1245 , RIb54aae0_15);
nor \U$564 ( \1247 , \1245 , RIb54aae0_15);
nor \U$565 ( \1248 , \1246 , \1247 );
and \U$566 ( \1249 , \1243 , \1248 );
not \U$567 ( \1250 , \1249 );
or \U$568 ( \1251 , \1241 , \741 );
nand \U$569 ( \1252 , \1251 , \695 );
nor \U$570 ( \1253 , \1250 , \1252 );
and \U$571 ( \1254 , \1237 , RIb54aa68_14);
nor \U$572 ( \1255 , \1237 , \700 );
nor \U$573 ( \1256 , \1254 , \1255 );
not \U$574 ( \1257 , \1256 );
not \U$575 ( \1258 , \704 );
or \U$576 ( \1259 , \1257 , \1258 );
not \U$577 ( \1260 , \1259 );
and \U$578 ( \1261 , \1240 , \703 );
and \U$579 ( \1262 , RIb54a9f0_13, \1237 );
nor \U$580 ( \1263 , \1261 , \1262 );
nor \U$581 ( \1264 , \1260 , \1263 );
and \U$582 ( \1265 , \1253 , \1264 );
and \U$583 ( \1266 , \1265 , RIb5515c0_243);
not \U$584 ( \1267 , \1263 );
nor \U$585 ( \1268 , \1267 , \1259 );
and \U$586 ( \1269 , \1253 , \1268 );
nand \U$587 ( \1270 , RIb551728_246, \1269 );
not \U$588 ( \1271 , \1243 );
nor \U$589 ( \1272 , \1271 , \1248 , \1252 );
and \U$590 ( \1273 , \1259 , \1263 );
and \U$591 ( \1274 , \1272 , \1273 );
and \U$592 ( \1275 , \1274 , RIb551458_240);
and \U$593 ( \1276 , \1272 , \1264 );
and \U$594 ( \1277 , RIb5513e0_239, \1276 );
nor \U$595 ( \1278 , \1275 , \1277 );
nor \U$596 ( \1279 , \1259 , \1263 );
and \U$597 ( \1280 , \1253 , \1279 );
nand \U$598 ( \1281 , RIb5516b0_245, \1280 );
nand \U$599 ( \1282 , \1270 , \1278 , \1281 );
and \U$600 ( \1283 , \1272 , \1268 );
and \U$601 ( \1284 , \1283 , RIb551548_242);
and \U$602 ( \1285 , \1272 , \1279 );
and \U$603 ( \1286 , RIb5514d0_241, \1285 );
nor \U$604 ( \1287 , \1284 , \1286 );
and \U$605 ( \1288 , \1268 , \1249 , \1252 );
and \U$606 ( \1289 , \1288 , RIb550be8_222);
not \U$607 ( \1290 , \1248 );
nor \U$608 ( \1291 , \1290 , \1243 , \1252 );
and \U$609 ( \1292 , \1291 , \1264 );
and \U$610 ( \1293 , RIb551200_235, \1292 );
nor \U$611 ( \1294 , \1289 , \1293 );
nand \U$612 ( \1295 , \1287 , \1294 );
nor \U$613 ( \1296 , \1266 , \1282 , \1295 );
and \U$614 ( \1297 , \1291 , \1268 );
and \U$615 ( \1298 , \1297 , RIb551368_238);
and \U$616 ( \1299 , \1291 , \1279 );
and \U$617 ( \1300 , RIb5512f0_237, \1299 );
nor \U$618 ( \1301 , \1298 , \1300 );
nor \U$619 ( \1302 , \1243 , \1248 , \1252 );
and \U$620 ( \1303 , \1302 , \1268 );
and \U$621 ( \1304 , \1303 , RIb551188_234);
and \U$622 ( \1305 , \1302 , \1279 );
and \U$623 ( \1306 , RIb551110_233, \1305 );
nor \U$624 ( \1307 , \1304 , \1306 );
and \U$625 ( \1308 , \1253 , \1273 );
and \U$626 ( \1309 , RIb551638_244, \1308 );
and \U$627 ( \1310 , \1302 , \1264 );
and \U$628 ( \1311 , RIb551020_231, \1310 );
and \U$629 ( \1312 , \1291 , \1273 );
and \U$630 ( \1313 , \1312 , RIb551278_236);
and \U$631 ( \1314 , \1302 , \1273 );
and \U$632 ( \1315 , RIb551098_232, \1314 );
nor \U$633 ( \1316 , \1313 , \1315 );
not \U$634 ( \1317 , \1316 );
nor \U$635 ( \1318 , \1309 , \1311 , \1317 );
nand \U$636 ( \1319 , \1296 , \1301 , \1307 , \1318 );
buf \U$637 ( \1320 , \766 );
_DC r1933 ( \1321_nR1933 , \1319 , \1320 );
not \U$638 ( \1322 , \1321_nR1933 );
nor \U$639 ( \1323 , \1233 , \1322 );
xor \U$640 ( \1324 , \694 , \768_nR12c0 );
xor \U$641 ( \1325 , \1324 , \1226 );
not \U$642 ( \1326 , \1325 );
xor \U$643 ( \1327 , \774 , \804_nR10db );
xor \U$644 ( \1328 , \1327 , \1223 );
not \U$645 ( \1329 , \1328 );
and \U$646 ( \1330 , \1326 , \1329 );
and \U$647 ( \1331 , \1229 , \1231 );
nor \U$648 ( \1332 , \1331 , \1232 );
nor \U$649 ( \1333 , \1330 , \1332 );
not \U$650 ( \1334 , \1333 );
and \U$651 ( \1335 , \1276 , RIb552448_274);
and \U$652 ( \1336 , \1308 , RIb5526a0_279);
and \U$653 ( \1337 , RIb552628_278, \1265 );
nor \U$654 ( \1338 , \1336 , \1337 );
and \U$655 ( \1339 , \1288 , RIb552010_265);
and \U$656 ( \1340 , RIb552268_270, \1292 );
nor \U$657 ( \1341 , \1339 , \1340 );
and \U$658 ( \1342 , \1283 , RIb5525b0_277);
and \U$659 ( \1343 , RIb552538_276, \1285 );
nor \U$660 ( \1344 , \1342 , \1343 );
and \U$661 ( \1345 , \1303 , RIb5521f0_269);
and \U$662 ( \1346 , RIb552178_268, \1305 );
nor \U$663 ( \1347 , \1345 , \1346 );
nand \U$664 ( \1348 , \1338 , \1341 , \1344 , \1347 );
and \U$665 ( \1349 , \1280 , RIb552718_280);
and \U$666 ( \1350 , RIb5524c0_275, \1274 );
nor \U$667 ( \1351 , \1349 , \1350 );
not \U$668 ( \1352 , \1351 );
nor \U$669 ( \1353 , \1335 , \1348 , \1352 );
and \U$670 ( \1354 , \1299 , RIb552358_272);
and \U$671 ( \1355 , RIb5522e0_271, \1312 );
nor \U$672 ( \1356 , \1354 , \1355 );
and \U$673 ( \1357 , \1314 , RIb552100_267);
and \U$674 ( \1358 , RIb552088_266, \1310 );
nor \U$675 ( \1359 , \1357 , \1358 );
and \U$676 ( \1360 , \1269 , RIb552790_281);
and \U$677 ( \1361 , RIb5523d0_273, \1297 );
nor \U$678 ( \1362 , \1360 , \1361 );
nand \U$679 ( \1363 , \1353 , \1356 , \1359 , \1362 );
_DC r1a4f ( \1364_nR1a4f , \1363 , \1320 );
or \U$680 ( \1365 , \1334 , \1364_nR1a4f );
not \U$681 ( \1366 , \1364_nR1a4f );
and \U$682 ( \1367 , \1332 , \1325 );
nor \U$683 ( \1368 , \1332 , \1325 );
xor \U$684 ( \1369 , \1325 , \1328 );
nor \U$685 ( \1370 , \1367 , \1368 , \1369 );
and \U$686 ( \1371 , \1370 , \1334 );
not \U$687 ( \1372 , \1371 );
or \U$688 ( \1373 , \1366 , \1372 );
or \U$689 ( \1374 , \1370 , \1334 );
nand \U$690 ( \1375 , \1365 , \1373 , \1374 );
xnor \U$691 ( \1376 , \1323 , \1375 );
not \U$692 ( \1377 , \1369 );
nor \U$693 ( \1378 , \1333 , \1377 );
not \U$694 ( \1379 , \1378 );
or \U$695 ( \1380 , \1379 , \1366 );
or \U$696 ( \1381 , \1322 , \1372 );
or \U$697 ( \1382 , \1377 , \1366 );
or \U$698 ( \1383 , \1334 , \1321_nR1933 );
nand \U$699 ( \1384 , \1383 , \1374 );
nand \U$700 ( \1385 , \1382 , \1384 );
nand \U$701 ( \1386 , \1380 , \1381 , \1385 );
xor \U$702 ( \1387 , \810 , \840_nR10d9 );
xor \U$703 ( \1388 , \1387 , \1220 );
xor \U$704 ( \1389 , \846 , \876_nRf20 );
xor \U$705 ( \1390 , \1389 , \1217 );
nor \U$706 ( \1391 , \1388 , \1390 );
or \U$707 ( \1392 , \1328 , \1391 );
and \U$708 ( \1393 , \1386 , \1392 );
and \U$709 ( \1394 , \1276 , RIb552c40_291);
and \U$710 ( \1395 , \1308 , RIb552e98_296);
and \U$711 ( \1396 , RIb552e20_295, \1265 );
nor \U$712 ( \1397 , \1395 , \1396 );
and \U$713 ( \1398 , \1288 , RIb552808_282);
and \U$714 ( \1399 , RIb552a60_287, \1292 );
nor \U$715 ( \1400 , \1398 , \1399 );
and \U$716 ( \1401 , \1283 , RIb552da8_294);
and \U$717 ( \1402 , RIb552d30_293, \1285 );
nor \U$718 ( \1403 , \1401 , \1402 );
and \U$719 ( \1404 , \1303 , RIb5529e8_286);
and \U$720 ( \1405 , RIb552970_285, \1305 );
nor \U$721 ( \1406 , \1404 , \1405 );
nand \U$722 ( \1407 , \1397 , \1400 , \1403 , \1406 );
and \U$723 ( \1408 , \1280 , RIb552f10_297);
and \U$724 ( \1409 , RIb552cb8_292, \1274 );
nor \U$725 ( \1410 , \1408 , \1409 );
not \U$726 ( \1411 , \1410 );
nor \U$727 ( \1412 , \1394 , \1407 , \1411 );
and \U$728 ( \1413 , \1299 , RIb552b50_289);
and \U$729 ( \1414 , RIb552ad8_288, \1312 );
nor \U$730 ( \1415 , \1413 , \1414 );
and \U$731 ( \1416 , \1314 , RIb5528f8_284);
and \U$732 ( \1417 , RIb552880_283, \1310 );
nor \U$733 ( \1418 , \1416 , \1417 );
and \U$734 ( \1419 , \1269 , RIb552f88_298);
and \U$735 ( \1420 , RIb552bc8_290, \1297 );
nor \U$736 ( \1421 , \1419 , \1420 );
nand \U$737 ( \1422 , \1412 , \1415 , \1418 , \1421 );
_DC r183c ( \1423_nR183c , \1422 , \1320 );
not \U$738 ( \1424 , \1423_nR183c );
nor \U$739 ( \1425 , \1233 , \1424 );
nor \U$740 ( \1426 , \1393 , \1425 );
xor \U$741 ( \1427 , \1376 , \1426 );
not \U$742 ( \1428 , \1427 );
or \U$743 ( \1429 , \1392 , \1364_nR1a4f );
and \U$744 ( \1430 , \1328 , \1388 );
nor \U$745 ( \1431 , \1328 , \1388 );
xor \U$746 ( \1432 , \1388 , \1390 );
nor \U$747 ( \1433 , \1430 , \1431 , \1432 );
and \U$748 ( \1434 , \1433 , \1392 );
not \U$749 ( \1435 , \1434 );
or \U$750 ( \1436 , \1366 , \1435 );
or \U$751 ( \1437 , \1433 , \1392 );
nand \U$752 ( \1438 , \1429 , \1436 , \1437 );
or \U$753 ( \1439 , \1379 , \1322 );
or \U$754 ( \1440 , \1424 , \1372 );
or \U$755 ( \1441 , \1377 , \1322 );
or \U$756 ( \1442 , \1334 , \1423_nR183c );
nand \U$757 ( \1443 , \1442 , \1374 );
nand \U$758 ( \1444 , \1441 , \1443 );
nand \U$759 ( \1445 , \1439 , \1440 , \1444 );
and \U$760 ( \1446 , \1438 , \1445 );
and \U$761 ( \1447 , \1386 , \1392 );
not \U$762 ( \1448 , \1386 );
not \U$763 ( \1449 , \1392 );
and \U$764 ( \1450 , \1448 , \1449 );
nor \U$765 ( \1451 , \1447 , \1450 );
xor \U$766 ( \1452 , \1425 , \1451 );
and \U$767 ( \1453 , \1446 , \1452 );
xor \U$768 ( \1454 , \1428 , \1453 );
nand \U$769 ( \1455 , \1364_nR1a4f , \1432 );
or \U$770 ( \1456 , \1392 , \1321_nR1933 );
nand \U$771 ( \1457 , \1456 , \1437 );
and \U$772 ( \1458 , \1455 , \1457 );
and \U$773 ( \1459 , \1434 , \1321_nR1933 );
not \U$774 ( \1460 , \1432 );
nor \U$775 ( \1461 , \1460 , \1449 );
and \U$776 ( \1462 , \1364_nR1a4f , \1461 );
nor \U$777 ( \1463 , \1458 , \1459 , \1462 );
and \U$778 ( \1464 , \1423_nR183c , \1378 );
and \U$779 ( \1465 , \1276 , RIb553c30_325);
and \U$780 ( \1466 , \1308 , RIb553e88_330);
and \U$781 ( \1467 , RIb553e10_329, \1265 );
nor \U$782 ( \1468 , \1466 , \1467 );
and \U$783 ( \1469 , \1288 , RIb5537f8_316);
and \U$784 ( \1470 , RIb553a50_321, \1292 );
nor \U$785 ( \1471 , \1469 , \1470 );
and \U$786 ( \1472 , \1283 , RIb553d98_328);
and \U$787 ( \1473 , RIb553d20_327, \1285 );
nor \U$788 ( \1474 , \1472 , \1473 );
and \U$789 ( \1475 , \1303 , RIb5539d8_320);
and \U$790 ( \1476 , RIb553960_319, \1305 );
nor \U$791 ( \1477 , \1475 , \1476 );
nand \U$792 ( \1478 , \1468 , \1471 , \1474 , \1477 );
and \U$793 ( \1479 , \1280 , RIb553f00_331);
and \U$794 ( \1480 , RIb553ca8_326, \1274 );
nor \U$795 ( \1481 , \1479 , \1480 );
not \U$796 ( \1482 , \1481 );
nor \U$797 ( \1483 , \1465 , \1478 , \1482 );
and \U$798 ( \1484 , \1299 , RIb553b40_323);
and \U$799 ( \1485 , RIb553ac8_322, \1312 );
nor \U$800 ( \1486 , \1484 , \1485 );
and \U$801 ( \1487 , \1314 , RIb5538e8_318);
and \U$802 ( \1488 , RIb553870_317, \1310 );
nor \U$803 ( \1489 , \1487 , \1488 );
and \U$804 ( \1490 , \1269 , RIb553f78_332);
and \U$805 ( \1491 , RIb553bb8_324, \1297 );
nor \U$806 ( \1492 , \1490 , \1491 );
nand \U$807 ( \1493 , \1483 , \1486 , \1489 , \1492 );
_DC r16fe ( \1494_nR16fe , \1493 , \1320 );
and \U$808 ( \1495 , \1371 , \1494_nR16fe );
nand \U$809 ( \1496 , \1423_nR183c , \1369 );
or \U$810 ( \1497 , \1334 , \1494_nR16fe );
nand \U$811 ( \1498 , \1497 , \1374 );
and \U$812 ( \1499 , \1496 , \1498 );
nor \U$813 ( \1500 , \1464 , \1495 , \1499 );
nand \U$814 ( \1501 , \1463 , \1500 );
xor \U$815 ( \1502 , \882 , \912_nRf1e );
xor \U$816 ( \1503 , \1502 , \1214 );
xor \U$817 ( \1504 , \918 , \948_nRda0 );
xor \U$818 ( \1505 , \1504 , \1211 );
nor \U$819 ( \1506 , \1503 , \1505 );
or \U$820 ( \1507 , \1390 , \1506 );
and \U$821 ( \1508 , \1501 , \1507 );
nor \U$822 ( \1509 , \1500 , \1463 );
nor \U$823 ( \1510 , \1508 , \1509 );
xor \U$824 ( \1511 , \1438 , \1445 );
not \U$825 ( \1512 , \1511 );
nand \U$826 ( \1513 , \1494_nR16fe , \1232 );
not \U$827 ( \1514 , \1513 );
and \U$828 ( \1515 , \1512 , \1514 );
and \U$829 ( \1516 , \1511 , \1513 );
nor \U$830 ( \1517 , \1515 , \1516 );
nand \U$831 ( \1518 , \1510 , \1517 );
xor \U$832 ( \1519 , \1446 , \1452 );
and \U$833 ( \1520 , \1518 , \1519 );
and \U$834 ( \1521 , \1454 , \1520 );
not \U$835 ( \1522 , \1521 );
and \U$836 ( \1523 , \1428 , \1453 );
or \U$837 ( \1524 , \1523 , \1333 );
and \U$838 ( \1525 , \1523 , \1333 );
and \U$839 ( \1526 , \1323 , \1375 );
nor \U$840 ( \1527 , \1525 , \1526 );
nand \U$841 ( \1528 , \1524 , \1527 );
not \U$842 ( \1529 , \1528 );
and \U$843 ( \1530 , \1232 , \1364_nR1a4f );
and \U$844 ( \1531 , \1376 , \1426 );
nor \U$845 ( \1532 , \1530 , \1531 );
not \U$846 ( \1533 , \1532 );
and \U$847 ( \1534 , \1529 , \1533 );
and \U$848 ( \1535 , \1528 , \1532 );
nor \U$849 ( \1536 , \1534 , \1535 );
not \U$850 ( \1537 , \1536 );
or \U$851 ( \1538 , \1522 , \1537 );
or \U$852 ( \1539 , \1536 , \1521 );
nand \U$853 ( \1540 , \1538 , \1539 );
not \U$854 ( \1541 , \1540 );
xor \U$855 ( \1542 , \1518 , \1519 );
not \U$856 ( \1543 , \1511 );
nor \U$857 ( \1544 , \1543 , \1513 );
xor \U$858 ( \1545 , \1542 , \1544 );
or \U$859 ( \1546 , \1517 , \1510 );
nand \U$860 ( \1547 , \1546 , \1518 );
not \U$861 ( \1548 , \1547 );
and \U$862 ( \1549 , \1265 , RIb553618_312);
nand \U$863 ( \1550 , RIb553780_315, \1269 );
and \U$864 ( \1551 , \1274 , RIb5534b0_309);
and \U$865 ( \1552 , RIb553438_308, \1276 );
nor \U$866 ( \1553 , \1551 , \1552 );
nand \U$867 ( \1554 , RIb553708_314, \1280 );
nand \U$868 ( \1555 , \1550 , \1553 , \1554 );
and \U$869 ( \1556 , \1283 , RIb5535a0_311);
and \U$870 ( \1557 , RIb553528_310, \1285 );
nor \U$871 ( \1558 , \1556 , \1557 );
and \U$872 ( \1559 , \1288 , RIb553000_299);
and \U$873 ( \1560 , RIb553258_304, \1292 );
nor \U$874 ( \1561 , \1559 , \1560 );
nand \U$875 ( \1562 , \1558 , \1561 );
nor \U$876 ( \1563 , \1549 , \1555 , \1562 );
and \U$877 ( \1564 , \1297 , RIb5533c0_307);
and \U$878 ( \1565 , RIb553348_306, \1299 );
nor \U$879 ( \1566 , \1564 , \1565 );
and \U$880 ( \1567 , \1303 , RIb5531e0_303);
and \U$881 ( \1568 , RIb553168_302, \1305 );
nor \U$882 ( \1569 , \1567 , \1568 );
and \U$883 ( \1570 , RIb553690_313, \1308 );
and \U$884 ( \1571 , RIb553078_300, \1310 );
and \U$885 ( \1572 , \1312 , RIb5532d0_305);
and \U$886 ( \1573 , RIb5530f0_301, \1314 );
nor \U$887 ( \1574 , \1572 , \1573 );
not \U$888 ( \1575 , \1574 );
nor \U$889 ( \1576 , \1570 , \1571 , \1575 );
nand \U$890 ( \1577 , \1563 , \1566 , \1569 , \1576 );
_DC r1611 ( \1578_nR1611 , \1577 , \1320 );
not \U$891 ( \1579 , \1578_nR1611 );
nor \U$892 ( \1580 , \1233 , \1579 );
not \U$893 ( \1581 , \1507 );
not \U$894 ( \1582 , \1509 );
nand \U$895 ( \1583 , \1582 , \1501 );
not \U$896 ( \1584 , \1583 );
or \U$897 ( \1585 , \1581 , \1584 );
or \U$898 ( \1586 , \1583 , \1507 );
nand \U$899 ( \1587 , \1585 , \1586 );
xnor \U$900 ( \1588 , \1580 , \1587 );
not \U$901 ( \1589 , \1588 );
and \U$902 ( \1590 , \1494_nR16fe , \1378 );
and \U$903 ( \1591 , \1371 , \1578_nR1611 );
nand \U$904 ( \1592 , \1494_nR16fe , \1369 );
or \U$905 ( \1593 , \1334 , \1578_nR1611 );
nand \U$906 ( \1594 , \1593 , \1374 );
and \U$907 ( \1595 , \1592 , \1594 );
nor \U$908 ( \1596 , \1590 , \1591 , \1595 );
and \U$909 ( \1597 , \1310 , RIb554068_334);
and \U$910 ( \1598 , \1308 , RIb554680_347);
and \U$911 ( \1599 , RIb554608_346, \1265 );
nor \U$912 ( \1600 , \1598 , \1599 );
and \U$913 ( \1601 , \1288 , RIb553ff0_333);
and \U$914 ( \1602 , RIb554248_338, \1292 );
nor \U$915 ( \1603 , \1601 , \1602 );
and \U$916 ( \1604 , \1283 , RIb554590_345);
and \U$917 ( \1605 , RIb554518_344, \1285 );
nor \U$918 ( \1606 , \1604 , \1605 );
and \U$919 ( \1607 , \1303 , RIb5541d0_337);
and \U$920 ( \1608 , RIb554158_336, \1305 );
nor \U$921 ( \1609 , \1607 , \1608 );
nand \U$922 ( \1610 , \1600 , \1603 , \1606 , \1609 );
and \U$923 ( \1611 , \1312 , RIb5542c0_339);
and \U$924 ( \1612 , RIb5540e0_335, \1314 );
nor \U$925 ( \1613 , \1611 , \1612 );
not \U$926 ( \1614 , \1613 );
nor \U$927 ( \1615 , \1597 , \1610 , \1614 );
and \U$928 ( \1616 , \1297 , RIb5543b0_341);
and \U$929 ( \1617 , RIb554338_340, \1299 );
nor \U$930 ( \1618 , \1616 , \1617 );
and \U$931 ( \1619 , \1274 , RIb5544a0_343);
and \U$932 ( \1620 , RIb554428_342, \1276 );
nor \U$933 ( \1621 , \1619 , \1620 );
and \U$934 ( \1622 , \1269 , RIb554770_349);
and \U$935 ( \1623 , RIb5546f8_348, \1280 );
nor \U$936 ( \1624 , \1622 , \1623 );
nand \U$937 ( \1625 , \1615 , \1618 , \1621 , \1624 );
_DC r14f1 ( \1626_nR14f1 , \1625 , \1320 );
nand \U$938 ( \1627 , \1626_nR14f1 , \1232 );
or \U$939 ( \1628 , \1596 , \1627 );
and \U$940 ( \1629 , \1390 , \1503 );
nor \U$941 ( \1630 , \1390 , \1503 );
xor \U$942 ( \1631 , \1503 , \1505 );
nor \U$943 ( \1632 , \1629 , \1630 , \1631 );
and \U$944 ( \1633 , \1632 , \1507 );
and \U$945 ( \1634 , \1364_nR1a4f , \1633 );
not \U$946 ( \1635 , \1507 );
and \U$947 ( \1636 , \1366 , \1635 );
or \U$948 ( \1637 , \1632 , \1507 );
not \U$949 ( \1638 , \1637 );
nor \U$950 ( \1639 , \1634 , \1636 , \1638 );
nand \U$951 ( \1640 , \1321_nR1933 , \1432 );
or \U$952 ( \1641 , \1392 , \1423_nR183c );
nand \U$953 ( \1642 , \1641 , \1437 );
and \U$954 ( \1643 , \1640 , \1642 );
and \U$955 ( \1644 , \1434 , \1423_nR183c );
and \U$956 ( \1645 , \1321_nR1933 , \1461 );
nor \U$957 ( \1646 , \1643 , \1644 , \1645 );
or \U$958 ( \1647 , \1639 , \1646 );
nand \U$959 ( \1648 , \1628 , \1647 );
nand \U$960 ( \1649 , \1589 , \1648 );
nor \U$961 ( \1650 , \1548 , \1649 );
and \U$962 ( \1651 , \1545 , \1650 );
and \U$963 ( \1652 , \1542 , \1544 );
or \U$964 ( \1653 , \1651 , \1652 );
xor \U$965 ( \1654 , \1454 , \1520 );
xor \U$966 ( \1655 , \1653 , \1654 );
xor \U$967 ( \1656 , \1542 , \1544 );
xor \U$968 ( \1657 , \1656 , \1650 );
and \U$969 ( \1658 , \1587 , \1580 );
not \U$970 ( \1659 , \1631 );
nor \U$971 ( \1660 , \1635 , \1659 );
not \U$972 ( \1661 , \1660 );
or \U$973 ( \1662 , \1661 , \1322 );
not \U$974 ( \1663 , \1633 );
or \U$975 ( \1664 , \1424 , \1663 );
or \U$976 ( \1665 , \1659 , \1322 );
or \U$977 ( \1666 , \1507 , \1423_nR183c );
nand \U$978 ( \1667 , \1666 , \1637 );
nand \U$979 ( \1668 , \1665 , \1667 );
nand \U$980 ( \1669 , \1662 , \1664 , \1668 );
not \U$981 ( \1670 , \1669 );
xor \U$982 ( \1671 , \954 , \984_nRd9e );
xor \U$983 ( \1672 , \1671 , \1208 );
xor \U$984 ( \1673 , \990 , \1020_nRc66 );
xor \U$985 ( \1674 , \1673 , \1205 );
nor \U$986 ( \1675 , \1672 , \1674 );
or \U$987 ( \1676 , \1505 , \1675 );
not \U$988 ( \1677 , \1676 );
not \U$989 ( \1678 , \1672 );
not \U$990 ( \1679 , \1505 );
or \U$991 ( \1680 , \1678 , \1679 );
or \U$992 ( \1681 , \1505 , \1672 );
nand \U$993 ( \1682 , \1680 , \1681 );
xor \U$994 ( \1683 , \1674 , \1672 );
nor \U$995 ( \1684 , \1682 , \1683 );
not \U$996 ( \1685 , \1684 );
nor \U$997 ( \1686 , \1677 , \1685 );
and \U$998 ( \1687 , \1686 , \1364_nR1a4f );
and \U$999 ( \1688 , \1684 , \1364_nR1a4f );
nor \U$1000 ( \1689 , \1688 , \1676 );
nor \U$1001 ( \1690 , \1687 , \1689 );
nor \U$1002 ( \1691 , \1670 , \1690 );
nand \U$1003 ( \1692 , \1494_nR16fe , \1432 );
or \U$1004 ( \1693 , \1392 , \1578_nR1611 );
nand \U$1005 ( \1694 , \1693 , \1437 );
and \U$1006 ( \1695 , \1692 , \1694 );
and \U$1007 ( \1696 , \1434 , \1578_nR1611 );
and \U$1008 ( \1697 , \1494_nR16fe , \1461 );
nor \U$1009 ( \1698 , \1695 , \1696 , \1697 );
and \U$1010 ( \1699 , \1297 , RIb554ba8_358);
and \U$1011 ( \1700 , \1283 , RIb554d88_362);
and \U$1012 ( \1701 , RIb554e00_363, \1265 );
nor \U$1013 ( \1702 , \1700 , \1701 );
and \U$1014 ( \1703 , \1303 , RIb5549c8_354);
and \U$1015 ( \1704 , RIb554950_353, \1305 );
nor \U$1016 ( \1705 , \1703 , \1704 );
and \U$1017 ( \1706 , \1285 , RIb554d10_361);
and \U$1018 ( \1707 , RIb554c98_360, \1274 );
nor \U$1019 ( \1708 , \1706 , \1707 );
and \U$1020 ( \1709 , \1288 , RIb5547e8_350);
and \U$1021 ( \1710 , RIb554ef0_365, \1280 );
nor \U$1022 ( \1711 , \1709 , \1710 );
nand \U$1023 ( \1712 , \1702 , \1705 , \1708 , \1711 );
and \U$1024 ( \1713 , \1308 , RIb554e78_364);
and \U$1025 ( \1714 , RIb554c20_359, \1276 );
nor \U$1026 ( \1715 , \1713 , \1714 );
not \U$1027 ( \1716 , \1715 );
nor \U$1028 ( \1717 , \1699 , \1712 , \1716 );
and \U$1029 ( \1718 , \1312 , RIb554ab8_356);
and \U$1030 ( \1719 , RIb554a40_355, \1292 );
nor \U$1031 ( \1720 , \1718 , \1719 );
and \U$1032 ( \1721 , \1314 , RIb5548d8_352);
and \U$1033 ( \1722 , RIb554860_351, \1310 );
nor \U$1034 ( \1723 , \1721 , \1722 );
and \U$1035 ( \1724 , \1269 , RIb554f68_366);
and \U$1036 ( \1725 , RIb554b30_357, \1299 );
nor \U$1037 ( \1726 , \1724 , \1725 );
nand \U$1038 ( \1727 , \1717 , \1720 , \1723 , \1726 );
_DC r12de ( \1728_nR12de , \1727 , \1320 );
nand \U$1039 ( \1729 , \1728_nR12de , \1232 );
and \U$1040 ( \1730 , \1698 , \1729 );
and \U$1041 ( \1731 , \1626_nR14f1 , \1378 );
and \U$1042 ( \1732 , \1310 , RIb555058_368);
and \U$1043 ( \1733 , \1308 , RIb555670_381);
and \U$1044 ( \1734 , RIb5555f8_380, \1265 );
nor \U$1045 ( \1735 , \1733 , \1734 );
and \U$1046 ( \1736 , \1288 , RIb554fe0_367);
and \U$1047 ( \1737 , RIb555238_372, \1292 );
nor \U$1048 ( \1738 , \1736 , \1737 );
and \U$1049 ( \1739 , \1283 , RIb555580_379);
and \U$1050 ( \1740 , RIb555508_378, \1285 );
nor \U$1051 ( \1741 , \1739 , \1740 );
and \U$1052 ( \1742 , \1303 , RIb5551c0_371);
and \U$1053 ( \1743 , RIb555148_370, \1305 );
nor \U$1054 ( \1744 , \1742 , \1743 );
nand \U$1055 ( \1745 , \1735 , \1738 , \1741 , \1744 );
and \U$1056 ( \1746 , \1312 , RIb5552b0_373);
and \U$1057 ( \1747 , RIb5550d0_369, \1314 );
nor \U$1058 ( \1748 , \1746 , \1747 );
not \U$1059 ( \1749 , \1748 );
nor \U$1060 ( \1750 , \1732 , \1745 , \1749 );
and \U$1061 ( \1751 , \1297 , RIb5553a0_375);
and \U$1062 ( \1752 , RIb555328_374, \1299 );
nor \U$1063 ( \1753 , \1751 , \1752 );
and \U$1064 ( \1754 , \1274 , RIb555490_377);
and \U$1065 ( \1755 , RIb555418_376, \1276 );
nor \U$1066 ( \1756 , \1754 , \1755 );
and \U$1067 ( \1757 , \1269 , RIb555760_383);
and \U$1068 ( \1758 , RIb5556e8_382, \1280 );
nor \U$1069 ( \1759 , \1757 , \1758 );
nand \U$1070 ( \1760 , \1750 , \1753 , \1756 , \1759 );
_DC r13ee ( \1761_nR13ee , \1760 , \1320 );
and \U$1071 ( \1762 , \1371 , \1761_nR13ee );
nand \U$1072 ( \1763 , \1626_nR14f1 , \1369 );
or \U$1073 ( \1764 , \1334 , \1761_nR13ee );
nand \U$1074 ( \1765 , \1764 , \1374 );
and \U$1075 ( \1766 , \1763 , \1765 );
nor \U$1076 ( \1767 , \1731 , \1762 , \1766 );
nor \U$1077 ( \1768 , \1730 , \1767 );
and \U$1078 ( \1769 , \1691 , \1768 );
not \U$1079 ( \1770 , \1676 );
nand \U$1080 ( \1771 , \1423_nR183c , \1432 );
or \U$1081 ( \1772 , \1392 , \1494_nR16fe );
nand \U$1082 ( \1773 , \1772 , \1437 );
and \U$1083 ( \1774 , \1771 , \1773 );
and \U$1084 ( \1775 , \1434 , \1494_nR16fe );
and \U$1085 ( \1776 , \1423_nR183c , \1461 );
nor \U$1086 ( \1777 , \1774 , \1775 , \1776 );
nand \U$1087 ( \1778 , \1364_nR1a4f , \1631 );
or \U$1088 ( \1779 , \1507 , \1321_nR1933 );
nand \U$1089 ( \1780 , \1779 , \1637 );
and \U$1090 ( \1781 , \1778 , \1780 );
and \U$1091 ( \1782 , \1633 , \1321_nR1933 );
and \U$1092 ( \1783 , \1364_nR1a4f , \1660 );
nor \U$1093 ( \1784 , \1781 , \1782 , \1783 );
nor \U$1094 ( \1785 , \1777 , \1784 );
not \U$1095 ( \1786 , \1785 );
nand \U$1096 ( \1787 , \1784 , \1777 );
nand \U$1097 ( \1788 , \1786 , \1787 );
not \U$1098 ( \1789 , \1788 );
or \U$1099 ( \1790 , \1770 , \1789 );
or \U$1100 ( \1791 , \1788 , \1676 );
nand \U$1101 ( \1792 , \1790 , \1791 );
not \U$1102 ( \1793 , \1792 );
and \U$1103 ( \1794 , \1578_nR1611 , \1378 );
and \U$1104 ( \1795 , \1371 , \1626_nR14f1 );
nand \U$1105 ( \1796 , \1578_nR1611 , \1369 );
or \U$1106 ( \1797 , \1334 , \1626_nR14f1 );
nand \U$1107 ( \1798 , \1797 , \1374 );
and \U$1108 ( \1799 , \1796 , \1798 );
nor \U$1109 ( \1800 , \1794 , \1795 , \1799 );
not \U$1110 ( \1801 , \1800 );
not \U$1111 ( \1802 , \1761_nR13ee );
nor \U$1112 ( \1803 , \1233 , \1802 );
not \U$1113 ( \1804 , \1803 );
and \U$1114 ( \1805 , \1801 , \1804 );
and \U$1115 ( \1806 , \1800 , \1803 );
nor \U$1116 ( \1807 , \1805 , \1806 );
nor \U$1117 ( \1808 , \1793 , \1807 );
and \U$1118 ( \1809 , \1769 , \1808 );
and \U$1119 ( \1810 , \1787 , \1676 );
not \U$1120 ( \1811 , \1803 );
nor \U$1121 ( \1812 , \1811 , \1800 );
nor \U$1122 ( \1813 , \1810 , \1812 , \1785 );
xor \U$1123 ( \1814 , \1627 , \1596 );
not \U$1124 ( \1815 , \1814 );
xnor \U$1125 ( \1816 , \1639 , \1646 );
not \U$1126 ( \1817 , \1816 );
and \U$1127 ( \1818 , \1815 , \1817 );
and \U$1128 ( \1819 , \1814 , \1816 );
nor \U$1129 ( \1820 , \1818 , \1819 );
nand \U$1130 ( \1821 , \1813 , \1820 );
xor \U$1131 ( \1822 , \1809 , \1821 );
not \U$1132 ( \1823 , \1648 );
not \U$1133 ( \1824 , \1588 );
or \U$1134 ( \1825 , \1823 , \1824 );
or \U$1135 ( \1826 , \1588 , \1648 );
nand \U$1136 ( \1827 , \1825 , \1826 );
and \U$1137 ( \1828 , \1822 , \1827 );
and \U$1138 ( \1829 , \1809 , \1821 );
or \U$1139 ( \1830 , \1828 , \1829 );
nor \U$1140 ( \1831 , \1658 , \1830 );
not \U$1141 ( \1832 , \1649 );
not \U$1142 ( \1833 , \1547 );
and \U$1143 ( \1834 , \1832 , \1833 );
and \U$1144 ( \1835 , \1649 , \1547 );
nor \U$1145 ( \1836 , \1834 , \1835 );
nor \U$1146 ( \1837 , \1831 , \1836 );
xor \U$1147 ( \1838 , \1657 , \1837 );
and \U$1148 ( \1839 , \1831 , \1836 );
nor \U$1149 ( \1840 , \1839 , \1837 );
and \U$1150 ( \1841 , \1321_nR1933 , \1686 );
or \U$1151 ( \1842 , \1676 , \1364_nR1a4f );
or \U$1152 ( \1843 , \1676 , \1683 );
nand \U$1153 ( \1844 , \1842 , \1843 );
nand \U$1154 ( \1845 , \1321_nR1933 , \1684 );
and \U$1155 ( \1846 , \1844 , \1845 );
and \U$1156 ( \1847 , \1676 , \1683 );
and \U$1157 ( \1848 , \1364_nR1a4f , \1847 );
nor \U$1158 ( \1849 , \1841 , \1846 , \1848 );
not \U$1159 ( \1850 , \1849 );
xor \U$1160 ( \1851 , \1026 , \1056_nRc64 );
xor \U$1161 ( \1852 , \1851 , \1202 );
xor \U$1162 ( \1853 , \1062 , \1092_nRb7a );
xor \U$1163 ( \1854 , \1853 , \1199 );
nor \U$1164 ( \1855 , \1852 , \1854 );
or \U$1165 ( \1856 , \1674 , \1855 );
not \U$1166 ( \1857 , \1856 );
not \U$1167 ( \1858 , \1857 );
and \U$1168 ( \1859 , \1850 , \1858 );
and \U$1169 ( \1860 , \1849 , \1857 );
nand \U$1170 ( \1861 , \1423_nR183c , \1631 );
or \U$1171 ( \1862 , \1507 , \1494_nR16fe );
nand \U$1172 ( \1863 , \1862 , \1637 );
and \U$1173 ( \1864 , \1861 , \1863 );
and \U$1174 ( \1865 , \1633 , \1494_nR16fe );
and \U$1175 ( \1866 , \1423_nR183c , \1660 );
nor \U$1176 ( \1867 , \1864 , \1865 , \1866 );
nor \U$1177 ( \1868 , \1860 , \1867 );
nor \U$1178 ( \1869 , \1859 , \1868 );
not \U$1179 ( \1870 , \1869 );
nand \U$1180 ( \1871 , \1578_nR1611 , \1432 );
or \U$1181 ( \1872 , \1392 , \1626_nR14f1 );
nand \U$1182 ( \1873 , \1872 , \1437 );
and \U$1183 ( \1874 , \1871 , \1873 );
and \U$1184 ( \1875 , \1434 , \1626_nR14f1 );
and \U$1185 ( \1876 , \1578_nR1611 , \1461 );
nor \U$1186 ( \1877 , \1874 , \1875 , \1876 );
and \U$1187 ( \1878 , \1265 , RIb5565e8_414);
nand \U$1188 ( \1879 , RIb556750_417, \1269 );
and \U$1189 ( \1880 , \1274 , RIb556480_411);
and \U$1190 ( \1881 , RIb556408_410, \1276 );
nor \U$1191 ( \1882 , \1880 , \1881 );
nand \U$1192 ( \1883 , RIb5566d8_416, \1280 );
nand \U$1193 ( \1884 , \1879 , \1882 , \1883 );
and \U$1194 ( \1885 , \1283 , RIb556570_413);
and \U$1195 ( \1886 , RIb5564f8_412, \1285 );
nor \U$1196 ( \1887 , \1885 , \1886 );
and \U$1197 ( \1888 , \1288 , RIb555fd0_401);
and \U$1198 ( \1889 , RIb556228_406, \1292 );
nor \U$1199 ( \1890 , \1888 , \1889 );
nand \U$1200 ( \1891 , \1887 , \1890 );
nor \U$1201 ( \1892 , \1878 , \1884 , \1891 );
and \U$1202 ( \1893 , \1297 , RIb556390_409);
and \U$1203 ( \1894 , RIb556318_408, \1299 );
nor \U$1204 ( \1895 , \1893 , \1894 );
and \U$1205 ( \1896 , \1303 , RIb5561b0_405);
and \U$1206 ( \1897 , RIb556138_404, \1305 );
nor \U$1207 ( \1898 , \1896 , \1897 );
and \U$1208 ( \1899 , RIb556660_415, \1308 );
and \U$1209 ( \1900 , RIb556048_402, \1310 );
and \U$1210 ( \1901 , \1312 , RIb5562a0_407);
and \U$1211 ( \1902 , RIb5560c0_403, \1314 );
nor \U$1212 ( \1903 , \1901 , \1902 );
not \U$1213 ( \1904 , \1903 );
nor \U$1214 ( \1905 , \1899 , \1900 , \1904 );
nand \U$1215 ( \1906 , \1892 , \1895 , \1898 , \1905 );
_DC r1200 ( \1907_nR1200 , \1906 , \1320 );
nand \U$1216 ( \1908 , \1907_nR1200 , \1232 );
and \U$1217 ( \1909 , \1877 , \1908 );
and \U$1218 ( \1910 , \1761_nR13ee , \1378 );
and \U$1219 ( \1911 , \1371 , \1728_nR12de );
nand \U$1220 ( \1912 , \1761_nR13ee , \1369 );
or \U$1221 ( \1913 , \1334 , \1728_nR12de );
nand \U$1222 ( \1914 , \1913 , \1374 );
and \U$1223 ( \1915 , \1912 , \1914 );
nor \U$1224 ( \1916 , \1910 , \1911 , \1915 );
nor \U$1225 ( \1917 , \1909 , \1916 );
nand \U$1226 ( \1918 , \1870 , \1917 );
not \U$1227 ( \1919 , \1918 );
not \U$1228 ( \1920 , \1729 );
not \U$1229 ( \1921 , \1767 );
not \U$1230 ( \1922 , \1698 );
and \U$1231 ( \1923 , \1921 , \1922 );
and \U$1232 ( \1924 , \1767 , \1698 );
nor \U$1233 ( \1925 , \1923 , \1924 );
not \U$1234 ( \1926 , \1925 );
or \U$1235 ( \1927 , \1920 , \1926 );
or \U$1236 ( \1928 , \1925 , \1729 );
nand \U$1237 ( \1929 , \1927 , \1928 );
not \U$1238 ( \1930 , \1929 );
not \U$1239 ( \1931 , \1669 );
not \U$1240 ( \1932 , \1690 );
and \U$1241 ( \1933 , \1931 , \1932 );
and \U$1242 ( \1934 , \1669 , \1690 );
nor \U$1243 ( \1935 , \1933 , \1934 );
nor \U$1244 ( \1936 , \1930 , \1935 );
nand \U$1245 ( \1937 , \1919 , \1936 );
not \U$1246 ( \1938 , \1807 );
not \U$1247 ( \1939 , \1792 );
and \U$1248 ( \1940 , \1938 , \1939 );
and \U$1249 ( \1941 , \1807 , \1792 );
nor \U$1250 ( \1942 , \1940 , \1941 );
not \U$1251 ( \1943 , \1942 );
xor \U$1252 ( \1944 , \1691 , \1768 );
nand \U$1253 ( \1945 , \1943 , \1944 );
and \U$1254 ( \1946 , \1937 , \1945 );
not \U$1255 ( \1947 , \1820 );
not \U$1256 ( \1948 , \1813 );
and \U$1257 ( \1949 , \1947 , \1948 );
not \U$1258 ( \1950 , \1821 );
nor \U$1259 ( \1951 , \1949 , \1950 );
nor \U$1260 ( \1952 , \1946 , \1951 );
not \U$1261 ( \1953 , \1814 );
nor \U$1262 ( \1954 , \1953 , \1816 );
xor \U$1263 ( \1955 , \1952 , \1954 );
xor \U$1264 ( \1956 , \1809 , \1821 );
xor \U$1265 ( \1957 , \1956 , \1827 );
and \U$1266 ( \1958 , \1955 , \1957 );
and \U$1267 ( \1959 , \1952 , \1954 );
or \U$1268 ( \1960 , \1958 , \1959 );
xor \U$1269 ( \1961 , \1840 , \1960 );
xor \U$1270 ( \1962 , \1952 , \1954 );
xor \U$1271 ( \1963 , \1962 , \1957 );
not \U$1272 ( \1964 , \1852 );
not \U$1273 ( \1965 , \1674 );
or \U$1274 ( \1966 , \1964 , \1965 );
or \U$1275 ( \1967 , \1674 , \1852 );
nand \U$1276 ( \1968 , \1966 , \1967 );
xor \U$1277 ( \1969 , \1854 , \1852 );
nor \U$1278 ( \1970 , \1968 , \1969 );
not \U$1279 ( \1971 , \1970 );
nor \U$1280 ( \1972 , \1971 , \1857 );
not \U$1281 ( \1973 , \1972 );
or \U$1282 ( \1974 , \1973 , \1366 );
or \U$1283 ( \1975 , \1971 , \1366 );
nand \U$1284 ( \1976 , \1975 , \1857 );
nand \U$1285 ( \1977 , \1974 , \1976 );
not \U$1286 ( \1978 , \1686 );
or \U$1287 ( \1979 , \1978 , \1424 );
not \U$1288 ( \1980 , \1847 );
or \U$1289 ( \1981 , \1322 , \1980 );
or \U$1290 ( \1982 , \1685 , \1424 );
or \U$1291 ( \1983 , \1676 , \1321_nR1933 );
nand \U$1292 ( \1984 , \1983 , \1843 );
nand \U$1293 ( \1985 , \1982 , \1984 );
nand \U$1294 ( \1986 , \1979 , \1981 , \1985 );
and \U$1295 ( \1987 , \1977 , \1986 );
nand \U$1296 ( \1988 , \1626_nR14f1 , \1432 );
or \U$1297 ( \1989 , \1392 , \1761_nR13ee );
nand \U$1298 ( \1990 , \1989 , \1437 );
and \U$1299 ( \1991 , \1988 , \1990 );
and \U$1300 ( \1992 , \1434 , \1761_nR13ee );
and \U$1301 ( \1993 , \1626_nR14f1 , \1461 );
nor \U$1302 ( \1994 , \1991 , \1992 , \1993 );
nand \U$1303 ( \1995 , \1494_nR16fe , \1631 );
or \U$1304 ( \1996 , \1507 , \1578_nR1611 );
nand \U$1305 ( \1997 , \1996 , \1637 );
and \U$1306 ( \1998 , \1995 , \1997 );
and \U$1307 ( \1999 , \1633 , \1578_nR1611 );
and \U$1308 ( \2000 , \1494_nR16fe , \1660 );
nor \U$1309 ( \2001 , \1998 , \1999 , \2000 );
xor \U$1310 ( \2002 , \1994 , \2001 );
and \U$1311 ( \2003 , \1728_nR12de , \1378 );
and \U$1312 ( \2004 , \1371 , \1907_nR1200 );
nand \U$1313 ( \2005 , \1728_nR12de , \1369 );
or \U$1314 ( \2006 , \1334 , \1907_nR1200 );
nand \U$1315 ( \2007 , \2006 , \1374 );
and \U$1316 ( \2008 , \2005 , \2007 );
nor \U$1317 ( \2009 , \2003 , \2004 , \2008 );
and \U$1318 ( \2010 , \2002 , \2009 );
and \U$1319 ( \2011 , \1994 , \2001 );
or \U$1320 ( \2012 , \2010 , \2011 );
not \U$1321 ( \2013 , \2012 );
and \U$1322 ( \2014 , \1987 , \2013 );
not \U$1323 ( \2015 , \1849 );
or \U$1324 ( \2016 , \1867 , \1856 );
nand \U$1325 ( \2017 , \1856 , \1867 );
nand \U$1326 ( \2018 , \2016 , \2017 );
not \U$1327 ( \2019 , \2018 );
or \U$1328 ( \2020 , \2015 , \2019 );
or \U$1329 ( \2021 , \2018 , \1849 );
nand \U$1330 ( \2022 , \2020 , \2021 );
not \U$1331 ( \2023 , \1908 );
not \U$1332 ( \2024 , \1916 );
not \U$1333 ( \2025 , \1877 );
and \U$1334 ( \2026 , \2024 , \2025 );
and \U$1335 ( \2027 , \1916 , \1877 );
nor \U$1336 ( \2028 , \2026 , \2027 );
not \U$1337 ( \2029 , \2028 );
or \U$1338 ( \2030 , \2023 , \2029 );
or \U$1339 ( \2031 , \2028 , \1908 );
nand \U$1340 ( \2032 , \2030 , \2031 );
and \U$1341 ( \2033 , \2022 , \2032 );
and \U$1342 ( \2034 , \2014 , \2033 );
not \U$1343 ( \2035 , \1917 );
not \U$1344 ( \2036 , \1869 );
and \U$1345 ( \2037 , \2035 , \2036 );
and \U$1346 ( \2038 , \1917 , \1869 );
nor \U$1347 ( \2039 , \2037 , \2038 );
not \U$1348 ( \2040 , \1929 );
not \U$1349 ( \2041 , \1935 );
and \U$1350 ( \2042 , \2040 , \2041 );
and \U$1351 ( \2043 , \1929 , \1935 );
nor \U$1352 ( \2044 , \2042 , \2043 );
nand \U$1353 ( \2045 , \2039 , \2044 );
xor \U$1354 ( \2046 , \2034 , \2045 );
not \U$1355 ( \2047 , \1944 );
not \U$1356 ( \2048 , \1942 );
or \U$1357 ( \2049 , \2047 , \2048 );
or \U$1358 ( \2050 , \1942 , \1944 );
nand \U$1359 ( \2051 , \2049 , \2050 );
and \U$1360 ( \2052 , \2046 , \2051 );
and \U$1361 ( \2053 , \2034 , \2045 );
or \U$1362 ( \2054 , \2052 , \2053 );
xor \U$1363 ( \2055 , \1769 , \1808 );
xor \U$1364 ( \2056 , \2054 , \2055 );
not \U$1365 ( \2057 , \1945 );
not \U$1366 ( \2058 , \1951 );
not \U$1367 ( \2059 , \1937 );
and \U$1368 ( \2060 , \2058 , \2059 );
and \U$1369 ( \2061 , \1951 , \1937 );
nor \U$1370 ( \2062 , \2060 , \2061 );
not \U$1371 ( \2063 , \2062 );
or \U$1372 ( \2064 , \2057 , \2063 );
or \U$1373 ( \2065 , \2062 , \1945 );
nand \U$1374 ( \2066 , \2064 , \2065 );
and \U$1375 ( \2067 , \2056 , \2066 );
and \U$1376 ( \2068 , \2054 , \2055 );
or \U$1377 ( \2069 , \2067 , \2068 );
xor \U$1378 ( \2070 , \1963 , \2069 );
not \U$1379 ( \2071 , \1918 );
not \U$1380 ( \2072 , \1936 );
or \U$1381 ( \2073 , \2071 , \2072 );
or \U$1382 ( \2074 , \1936 , \1918 );
nand \U$1383 ( \2075 , \2073 , \2074 );
xor \U$1384 ( \2076 , \2034 , \2045 );
xor \U$1385 ( \2077 , \2076 , \2051 );
and \U$1386 ( \2078 , \2075 , \2077 );
xor \U$1387 ( \2079 , \1987 , \2013 );
xor \U$1388 ( \2080 , \2022 , \2032 );
and \U$1389 ( \2081 , \2079 , \2080 );
xor \U$1390 ( \2082 , \1977 , \1986 );
not \U$1391 ( \2083 , \2082 );
xor \U$1392 ( \2084 , \1994 , \2001 );
xor \U$1393 ( \2085 , \2084 , \2009 );
nor \U$1394 ( \2086 , \2083 , \2085 );
nand \U$1395 ( \2087 , \1761_nR13ee , \1432 );
or \U$1396 ( \2088 , \1392 , \1728_nR12de );
nand \U$1397 ( \2089 , \2088 , \1437 );
and \U$1398 ( \2090 , \2087 , \2089 );
and \U$1399 ( \2091 , \1434 , \1728_nR12de );
and \U$1400 ( \2092 , \1761_nR13ee , \1461 );
nor \U$1401 ( \2093 , \2090 , \2091 , \2092 );
nand \U$1402 ( \2094 , \1578_nR1611 , \1631 );
or \U$1403 ( \2095 , \1507 , \1626_nR14f1 );
nand \U$1404 ( \2096 , \2095 , \1637 );
and \U$1405 ( \2097 , \2094 , \2096 );
and \U$1406 ( \2098 , \1633 , \1626_nR14f1 );
and \U$1407 ( \2099 , \1578_nR1611 , \1660 );
nor \U$1408 ( \2100 , \2097 , \2098 , \2099 );
xor \U$1409 ( \2101 , \2093 , \2100 );
and \U$1410 ( \2102 , \1907_nR1200 , \1378 );
and \U$1411 ( \2103 , \1305 , RIb555940_387);
and \U$1412 ( \2104 , \1280 , RIb555ee0_399);
and \U$1413 ( \2105 , RIb555e68_398, \1308 );
nor \U$1414 ( \2106 , \2104 , \2105 );
and \U$1415 ( \2107 , \1312 , RIb555aa8_390);
and \U$1416 ( \2108 , RIb555a30_389, \1292 );
nor \U$1417 ( \2109 , \2107 , \2108 );
and \U$1418 ( \2110 , \1314 , RIb5558c8_386);
and \U$1419 ( \2111 , RIb555850_385, \1310 );
nor \U$1420 ( \2112 , \2110 , \2111 );
and \U$1421 ( \2113 , \1288 , RIb5557d8_384);
and \U$1422 ( \2114 , RIb555df0_397, \1265 );
nor \U$1423 ( \2115 , \2113 , \2114 );
nand \U$1424 ( \2116 , \2106 , \2109 , \2112 , \2115 );
and \U$1425 ( \2117 , \1299 , RIb555b20_391);
and \U$1426 ( \2118 , RIb5559b8_388, \1303 );
nor \U$1427 ( \2119 , \2117 , \2118 );
not \U$1428 ( \2120 , \2119 );
nor \U$1429 ( \2121 , \2103 , \2116 , \2120 );
and \U$1430 ( \2122 , \1297 , RIb555b98_392);
and \U$1431 ( \2123 , RIb555c10_393, \1276 );
nor \U$1432 ( \2124 , \2122 , \2123 );
and \U$1433 ( \2125 , \1285 , RIb555d00_395);
and \U$1434 ( \2126 , RIb555c88_394, \1274 );
nor \U$1435 ( \2127 , \2125 , \2126 );
and \U$1436 ( \2128 , \1269 , RIb555f58_400);
and \U$1437 ( \2129 , RIb555d78_396, \1283 );
nor \U$1438 ( \2130 , \2128 , \2129 );
nand \U$1439 ( \2131 , \2121 , \2124 , \2127 , \2130 );
_DC r10f9 ( \2132_nR10f9 , \2131 , \1320 );
and \U$1440 ( \2133 , \1371 , \2132_nR10f9 );
nand \U$1441 ( \2134 , \1907_nR1200 , \1369 );
or \U$1442 ( \2135 , \1334 , \2132_nR10f9 );
nand \U$1443 ( \2136 , \2135 , \1374 );
and \U$1444 ( \2137 , \2134 , \2136 );
nor \U$1445 ( \2138 , \2102 , \2133 , \2137 );
and \U$1446 ( \2139 , \2101 , \2138 );
and \U$1447 ( \2140 , \2093 , \2100 );
or \U$1448 ( \2141 , \2139 , \2140 );
nand \U$1449 ( \2142 , \1321_nR1933 , \1970 );
or \U$1450 ( \2143 , \1856 , \1364_nR1a4f );
or \U$1451 ( \2144 , \1856 , \1969 );
nand \U$1452 ( \2145 , \2143 , \2144 );
and \U$1453 ( \2146 , \2142 , \2145 );
and \U$1454 ( \2147 , \1856 , \1969 );
and \U$1455 ( \2148 , \2147 , \1364_nR1a4f );
and \U$1456 ( \2149 , \1321_nR1933 , \1972 );
nor \U$1457 ( \2150 , \2146 , \2148 , \2149 );
and \U$1458 ( \2151 , \1494_nR16fe , \1686 );
or \U$1459 ( \2152 , \1676 , \1423_nR183c );
nand \U$1460 ( \2153 , \2152 , \1843 );
nand \U$1461 ( \2154 , \1494_nR16fe , \1684 );
and \U$1462 ( \2155 , \2153 , \2154 );
and \U$1463 ( \2156 , \1423_nR183c , \1847 );
nor \U$1464 ( \2157 , \2151 , \2155 , \2156 );
nand \U$1465 ( \2158 , \2150 , \2157 );
xor \U$1466 ( \2159 , \1098 , \1128_nRb7c );
xor \U$1467 ( \2160 , \2159 , \1196 );
not \U$1468 ( \2161 , \2160 );
xor \U$1469 ( \2162 , RIb54a900_11, \1159_nR9e7 );
xor \U$1470 ( \2163 , \2162 , \1193 );
not \U$1471 ( \2164 , \2163 );
and \U$1472 ( \2165 , \2161 , \2164 );
nor \U$1473 ( \2166 , \2165 , \1854 );
not \U$1474 ( \2167 , \2166 );
and \U$1475 ( \2168 , \2158 , \2167 );
nor \U$1476 ( \2169 , \2157 , \2150 );
nor \U$1477 ( \2170 , \2168 , \2169 );
nor \U$1478 ( \2171 , \2141 , \2170 );
and \U$1479 ( \2172 , \2086 , \2171 );
xor \U$1480 ( \2173 , \2081 , \2172 );
or \U$1481 ( \2174 , \2044 , \2039 );
nand \U$1482 ( \2175 , \2174 , \2045 );
and \U$1483 ( \2176 , \2173 , \2175 );
and \U$1484 ( \2177 , \2081 , \2172 );
or \U$1485 ( \2178 , \2176 , \2177 );
xor \U$1486 ( \2179 , \2034 , \2045 );
xor \U$1487 ( \2180 , \2179 , \2051 );
and \U$1488 ( \2181 , \2178 , \2180 );
and \U$1489 ( \2182 , \2075 , \2178 );
or \U$1490 ( \2183 , \2078 , \2181 , \2182 );
xor \U$1491 ( \2184 , \2054 , \2055 );
xor \U$1492 ( \2185 , \2184 , \2066 );
xor \U$1493 ( \2186 , \2183 , \2185 );
xor \U$1494 ( \2187 , \2034 , \2045 );
xor \U$1495 ( \2188 , \2187 , \2051 );
xor \U$1496 ( \2189 , \2075 , \2178 );
xor \U$1497 ( \2190 , \2188 , \2189 );
not \U$1498 ( \2191 , \2085 );
not \U$1499 ( \2192 , \2082 );
and \U$1500 ( \2193 , \2191 , \2192 );
and \U$1501 ( \2194 , \2085 , \2082 );
nor \U$1502 ( \2195 , \2193 , \2194 );
not \U$1503 ( \2196 , \2132_nR10f9 );
nor \U$1504 ( \2197 , \1233 , \2196 );
or \U$1505 ( \2198 , \2195 , \2197 );
xnor \U$1506 ( \2199 , \2170 , \2141 );
nand \U$1507 ( \2200 , \2198 , \2199 );
not \U$1508 ( \2201 , \2160 );
not \U$1509 ( \2202 , \1854 );
or \U$1510 ( \2203 , \2201 , \2202 );
or \U$1511 ( \2204 , \1854 , \2160 );
nand \U$1512 ( \2205 , \2203 , \2204 );
or \U$1513 ( \2206 , \2161 , \2163 );
or \U$1514 ( \2207 , \2164 , \2160 );
nand \U$1515 ( \2208 , \2206 , \2207 );
nor \U$1516 ( \2209 , \2205 , \2208 );
not \U$1517 ( \2210 , \2209 );
nor \U$1518 ( \2211 , \2210 , \2166 );
not \U$1519 ( \2212 , \2211 );
or \U$1520 ( \2213 , \2212 , \1366 );
or \U$1521 ( \2214 , \2210 , \1366 );
nand \U$1522 ( \2215 , \2214 , \2166 );
nand \U$1523 ( \2216 , \2213 , \2215 );
not \U$1524 ( \2217 , \2216 );
nand \U$1525 ( \2218 , \1423_nR183c , \1970 );
or \U$1526 ( \2219 , \1856 , \1321_nR1933 );
nand \U$1527 ( \2220 , \2219 , \2144 );
and \U$1528 ( \2221 , \2218 , \2220 );
and \U$1529 ( \2222 , \2147 , \1321_nR1933 );
and \U$1530 ( \2223 , \1423_nR183c , \1972 );
nor \U$1531 ( \2224 , \2221 , \2222 , \2223 );
nor \U$1532 ( \2225 , \2217 , \2224 );
not \U$1533 ( \2226 , \2225 );
nand \U$1534 ( \2227 , \1626_nR14f1 , \1631 );
or \U$1535 ( \2228 , \1507 , \1761_nR13ee );
nand \U$1536 ( \2229 , \2228 , \1637 );
and \U$1537 ( \2230 , \2227 , \2229 );
and \U$1538 ( \2231 , \1633 , \1761_nR13ee );
and \U$1539 ( \2232 , \1626_nR14f1 , \1660 );
nor \U$1540 ( \2233 , \2230 , \2231 , \2232 );
and \U$1541 ( \2234 , \1578_nR1611 , \1686 );
or \U$1542 ( \2235 , \1676 , \1494_nR16fe );
nand \U$1543 ( \2236 , \2235 , \1843 );
nand \U$1544 ( \2237 , \1578_nR1611 , \1684 );
and \U$1545 ( \2238 , \2236 , \2237 );
and \U$1546 ( \2239 , \1494_nR16fe , \1847 );
nor \U$1547 ( \2240 , \2234 , \2238 , \2239 );
xor \U$1548 ( \2241 , \2233 , \2240 );
nand \U$1549 ( \2242 , \1728_nR12de , \1432 );
or \U$1550 ( \2243 , \1392 , \1907_nR1200 );
nand \U$1551 ( \2244 , \2243 , \1437 );
and \U$1552 ( \2245 , \2242 , \2244 );
and \U$1553 ( \2246 , \1434 , \1907_nR1200 );
and \U$1554 ( \2247 , \1728_nR12de , \1461 );
nor \U$1555 ( \2248 , \2245 , \2246 , \2247 );
and \U$1556 ( \2249 , \2241 , \2248 );
and \U$1557 ( \2250 , \2233 , \2240 );
or \U$1558 ( \2251 , \2249 , \2250 );
nor \U$1559 ( \2252 , \2226 , \2251 );
not \U$1560 ( \2253 , \2252 );
and \U$1561 ( \2254 , \1299 , RIb557308_442);
and \U$1562 ( \2255 , \1283 , RIb557560_447);
and \U$1563 ( \2256 , RIb5575d8_448, \1265 );
nor \U$1564 ( \2257 , \2255 , \2256 );
and \U$1565 ( \2258 , \1303 , RIb5571a0_439);
and \U$1566 ( \2259 , RIb557128_438, \1305 );
nor \U$1567 ( \2260 , \2258 , \2259 );
and \U$1568 ( \2261 , \1285 , RIb5574e8_446);
and \U$1569 ( \2262 , RIb557470_445, \1274 );
nor \U$1570 ( \2263 , \2261 , \2262 );
and \U$1571 ( \2264 , \1288 , RIb556fc0_435);
and \U$1572 ( \2265 , RIb557650_449, \1308 );
nor \U$1573 ( \2266 , \2264 , \2265 );
nand \U$1574 ( \2267 , \2257 , \2260 , \2263 , \2266 );
and \U$1575 ( \2268 , \1297 , RIb557380_443);
and \U$1576 ( \2269 , RIb5573f8_444, \1276 );
nor \U$1577 ( \2270 , \2268 , \2269 );
not \U$1578 ( \2271 , \2270 );
nor \U$1579 ( \2272 , \2254 , \2267 , \2271 );
and \U$1580 ( \2273 , \1312 , RIb557290_441);
and \U$1581 ( \2274 , RIb557218_440, \1292 );
nor \U$1582 ( \2275 , \2273 , \2274 );
and \U$1583 ( \2276 , \1314 , RIb5570b0_437);
and \U$1584 ( \2277 , RIb557038_436, \1310 );
nor \U$1585 ( \2278 , \2276 , \2277 );
and \U$1586 ( \2279 , \1269 , RIb557740_451);
and \U$1587 ( \2280 , RIb5576c8_450, \1280 );
nor \U$1588 ( \2281 , \2279 , \2280 );
nand \U$1589 ( \2282 , \2272 , \2275 , \2278 , \2281 );
_DC r101a ( \2283_nR101a , \2282 , \1320 );
nand \U$1590 ( \2284 , \2283_nR101a , \1232 );
not \U$1591 ( \2285 , \2284 );
not \U$1592 ( \2286 , \2166 );
not \U$1593 ( \2287 , \2158 );
nor \U$1594 ( \2288 , \2287 , \2169 );
not \U$1595 ( \2289 , \2288 );
or \U$1596 ( \2290 , \2286 , \2289 );
or \U$1597 ( \2291 , \2288 , \2166 );
nand \U$1598 ( \2292 , \2290 , \2291 );
xor \U$1599 ( \2293 , \2093 , \2100 );
xor \U$1600 ( \2294 , \2293 , \2138 );
not \U$1601 ( \2295 , \2294 );
and \U$1602 ( \2296 , \2292 , \2295 );
nor \U$1603 ( \2297 , \2285 , \2296 );
nor \U$1604 ( \2298 , \2253 , \2297 );
xor \U$1605 ( \2299 , \2200 , \2298 );
xor \U$1606 ( \2300 , \2079 , \2080 );
and \U$1607 ( \2301 , \2299 , \2300 );
and \U$1608 ( \2302 , \2200 , \2298 );
or \U$1609 ( \2303 , \2301 , \2302 );
xor \U$1610 ( \2304 , \2014 , \2033 );
xor \U$1611 ( \2305 , \2303 , \2304 );
xor \U$1612 ( \2306 , \2081 , \2172 );
xor \U$1613 ( \2307 , \2306 , \2175 );
and \U$1614 ( \2308 , \2305 , \2307 );
and \U$1615 ( \2309 , \2303 , \2304 );
or \U$1616 ( \2310 , \2308 , \2309 );
xor \U$1617 ( \2311 , \2190 , \2310 );
xor \U$1618 ( \2312 , \2303 , \2304 );
xor \U$1619 ( \2313 , \2312 , \2307 );
xor \U$1620 ( \2314 , \2200 , \2298 );
xor \U$1621 ( \2315 , \2314 , \2300 );
not \U$1622 ( \2316 , \2315 );
not \U$1623 ( \2317 , \2199 );
xor \U$1624 ( \2318 , \2197 , \2195 );
not \U$1625 ( \2319 , \2318 );
or \U$1626 ( \2320 , \2317 , \2319 );
or \U$1627 ( \2321 , \2318 , \2199 );
nand \U$1628 ( \2322 , \2320 , \2321 );
nand \U$1629 ( \2323 , \1761_nR13ee , \1631 );
or \U$1630 ( \2324 , \1507 , \1728_nR12de );
nand \U$1631 ( \2325 , \2324 , \1637 );
and \U$1632 ( \2326 , \2323 , \2325 );
and \U$1633 ( \2327 , \1633 , \1728_nR12de );
and \U$1634 ( \2328 , \1761_nR13ee , \1660 );
nor \U$1635 ( \2329 , \2326 , \2327 , \2328 );
and \U$1636 ( \2330 , \1626_nR14f1 , \1686 );
or \U$1637 ( \2331 , \1676 , \1578_nR1611 );
nand \U$1638 ( \2332 , \2331 , \1843 );
nand \U$1639 ( \2333 , \1626_nR14f1 , \1684 );
and \U$1640 ( \2334 , \2332 , \2333 );
and \U$1641 ( \2335 , \1578_nR1611 , \1847 );
nor \U$1642 ( \2336 , \2330 , \2334 , \2335 );
xor \U$1643 ( \2337 , \2329 , \2336 );
nand \U$1644 ( \2338 , \1907_nR1200 , \1432 );
or \U$1645 ( \2339 , \1392 , \2132_nR10f9 );
nand \U$1646 ( \2340 , \2339 , \1437 );
and \U$1647 ( \2341 , \2338 , \2340 );
and \U$1648 ( \2342 , \1434 , \2132_nR10f9 );
and \U$1649 ( \2343 , \1907_nR1200 , \1461 );
nor \U$1650 ( \2344 , \2341 , \2342 , \2343 );
and \U$1651 ( \2345 , \2337 , \2344 );
and \U$1652 ( \2346 , \2329 , \2336 );
or \U$1653 ( \2347 , \2345 , \2346 );
nand \U$1654 ( \2348 , \1321_nR1933 , \2209 );
or \U$1655 ( \2349 , \2167 , \1364_nR1a4f );
or \U$1656 ( \2350 , \2167 , \2208 );
nand \U$1657 ( \2351 , \2349 , \2350 );
and \U$1658 ( \2352 , \2348 , \2351 );
and \U$1659 ( \2353 , \2167 , \2208 );
and \U$1660 ( \2354 , \2353 , \1364_nR1a4f );
and \U$1661 ( \2355 , \1321_nR1933 , \2211 );
nor \U$1662 ( \2356 , \2352 , \2354 , \2355 );
xor \U$1663 ( \2357 , \2356 , \2164 );
nand \U$1664 ( \2358 , \1494_nR16fe , \1970 );
or \U$1665 ( \2359 , \1856 , \1423_nR183c );
nand \U$1666 ( \2360 , \2359 , \2144 );
and \U$1667 ( \2361 , \2358 , \2360 );
and \U$1668 ( \2362 , \2147 , \1423_nR183c );
and \U$1669 ( \2363 , \1494_nR16fe , \1972 );
nor \U$1670 ( \2364 , \2361 , \2362 , \2363 );
and \U$1671 ( \2365 , \2357 , \2364 );
and \U$1672 ( \2366 , \2356 , \2164 );
or \U$1673 ( \2367 , \2365 , \2366 );
nor \U$1674 ( \2368 , \2347 , \2367 );
not \U$1675 ( \2369 , \2368 );
xor \U$1676 ( \2370 , \2233 , \2240 );
xor \U$1677 ( \2371 , \2370 , \2248 );
not \U$1678 ( \2372 , \2224 );
not \U$1679 ( \2373 , \2216 );
and \U$1680 ( \2374 , \2372 , \2373 );
and \U$1681 ( \2375 , \2224 , \2216 );
nor \U$1682 ( \2376 , \2374 , \2375 );
xor \U$1683 ( \2377 , \2371 , \2376 );
and \U$1684 ( \2378 , \1276 , RIb556c00_427);
and \U$1685 ( \2379 , \1280 , RIb556ed0_433);
and \U$1686 ( \2380 , RIb556e58_432, \1308 );
nor \U$1687 ( \2381 , \2379 , \2380 );
and \U$1688 ( \2382 , \1303 , RIb5569a8_422);
and \U$1689 ( \2383 , RIb556930_421, \1305 );
nor \U$1690 ( \2384 , \2382 , \2383 );
and \U$1691 ( \2385 , \1288 , RIb5567c8_418);
and \U$1692 ( \2386 , RIb556a20_423, \1292 );
nor \U$1693 ( \2387 , \2385 , \2386 );
and \U$1694 ( \2388 , \1283 , RIb556d68_430);
and \U$1695 ( \2389 , RIb556de0_431, \1265 );
nor \U$1696 ( \2390 , \2388 , \2389 );
nand \U$1697 ( \2391 , \2381 , \2384 , \2387 , \2390 );
and \U$1698 ( \2392 , \1285 , RIb556cf0_429);
and \U$1699 ( \2393 , RIb556c78_428, \1274 );
nor \U$1700 ( \2394 , \2392 , \2393 );
not \U$1701 ( \2395 , \2394 );
nor \U$1702 ( \2396 , \2378 , \2391 , \2395 );
and \U$1703 ( \2397 , \1299 , RIb556b10_425);
and \U$1704 ( \2398 , RIb556a98_424, \1312 );
nor \U$1705 ( \2399 , \2397 , \2398 );
and \U$1706 ( \2400 , \1314 , RIb5568b8_420);
and \U$1707 ( \2401 , RIb556840_419, \1310 );
nor \U$1708 ( \2402 , \2400 , \2401 );
and \U$1709 ( \2403 , \1269 , RIb556f48_434);
and \U$1710 ( \2404 , RIb556b88_426, \1297 );
nor \U$1711 ( \2405 , \2403 , \2404 );
nand \U$1712 ( \2406 , \2396 , \2399 , \2402 , \2405 );
_DC rf3e ( \2407_nRf3e , \2406 , \1320 );
nand \U$1713 ( \2408 , \2407_nRf3e , \1232 );
and \U$1714 ( \2409 , \2132_nR10f9 , \1378 );
and \U$1715 ( \2410 , \1371 , \2283_nR101a );
nand \U$1716 ( \2411 , \2132_nR10f9 , \1369 );
or \U$1717 ( \2412 , \1334 , \2283_nR101a );
nand \U$1718 ( \2413 , \2412 , \1374 );
and \U$1719 ( \2414 , \2411 , \2413 );
nor \U$1720 ( \2415 , \2409 , \2410 , \2414 );
xnor \U$1721 ( \2416 , \2408 , \2415 );
and \U$1722 ( \2417 , \2377 , \2416 );
and \U$1723 ( \2418 , \2371 , \2376 );
or \U$1724 ( \2419 , \2417 , \2418 );
nor \U$1725 ( \2420 , \2369 , \2419 );
nor \U$1726 ( \2421 , \2322 , \2420 );
xor \U$1727 ( \2422 , \2292 , \2295 );
not \U$1728 ( \2423 , \2422 );
not \U$1729 ( \2424 , \2284 );
and \U$1730 ( \2425 , \2423 , \2424 );
and \U$1731 ( \2426 , \2422 , \2284 );
nor \U$1732 ( \2427 , \2425 , \2426 );
not \U$1733 ( \2428 , \2427 );
or \U$1734 ( \2429 , \2251 , \2225 );
or \U$1735 ( \2430 , \2408 , \2415 );
nand \U$1736 ( \2431 , \2225 , \2251 );
nand \U$1737 ( \2432 , \2429 , \2430 , \2431 );
nand \U$1738 ( \2433 , \2428 , \2432 );
or \U$1739 ( \2434 , \2421 , \2433 );
nand \U$1740 ( \2435 , \2420 , \2322 );
nand \U$1741 ( \2436 , \2434 , \2435 );
nor \U$1742 ( \2437 , \2171 , \2197 );
not \U$1743 ( \2438 , \2437 );
not \U$1744 ( \2439 , \2086 );
or \U$1745 ( \2440 , \2438 , \2439 );
or \U$1746 ( \2441 , \2086 , \2437 );
nand \U$1747 ( \2442 , \2440 , \2441 );
or \U$1748 ( \2443 , \2436 , \2442 );
not \U$1749 ( \2444 , \2443 );
or \U$1750 ( \2445 , \2316 , \2444 );
nand \U$1751 ( \2446 , \2442 , \2436 );
nand \U$1752 ( \2447 , \2445 , \2446 );
and \U$1753 ( \2448 , \2313 , \2447 );
not \U$1754 ( \2449 , \2313 );
not \U$1755 ( \2450 , \2447 );
and \U$1756 ( \2451 , \2449 , \2450 );
and \U$1757 ( \2452 , RIb557fb0_469, \1288 );
and \U$1758 ( \2453 , RIb5580a0_471, \1314 );
and \U$1759 ( \2454 , RIb5585c8_482, \1265 );
and \U$1760 ( \2455 , RIb558028_470, \1310 );
and \U$1761 ( \2456 , \1297 , RIb558370_477);
and \U$1762 ( \2457 , RIb5582f8_476, \1299 );
nor \U$1763 ( \2458 , \2456 , \2457 );
not \U$1764 ( \2459 , \2458 );
nor \U$1765 ( \2460 , \2454 , \2455 , \2459 );
and \U$1766 ( \2461 , \1312 , RIb558280_475);
and \U$1767 ( \2462 , RIb558208_474, \1292 );
nor \U$1768 ( \2463 , \2461 , \2462 );
nand \U$1769 ( \2464 , RIb558730_485, \1269 );
and \U$1770 ( \2465 , \1308 , RIb558640_483);
and \U$1771 ( \2466 , RIb558550_481, \1283 );
nor \U$1772 ( \2467 , \2465 , \2466 );
nand \U$1773 ( \2468 , \2460 , \2463 , \2464 , \2467 );
nor \U$1774 ( \2469 , \2452 , \2453 , \2468 );
and \U$1775 ( \2470 , \1303 , RIb558190_473);
and \U$1776 ( \2471 , RIb558118_472, \1305 );
nor \U$1777 ( \2472 , \2470 , \2471 );
and \U$1778 ( \2473 , \1274 , RIb558460_479);
and \U$1779 ( \2474 , RIb5583e8_478, \1276 );
nor \U$1780 ( \2475 , \2473 , \2474 );
and \U$1781 ( \2476 , \1280 , RIb5586b8_484);
and \U$1782 ( \2477 , RIb5584d8_480, \1285 );
nor \U$1783 ( \2478 , \2476 , \2477 );
nand \U$1784 ( \2479 , \2469 , \2472 , \2475 , \2478 );
_DC re8d ( \2480_nRe8d , \2479 , \1320 );
nand \U$1785 ( \2481 , \2480_nRe8d , \1232 );
and \U$1786 ( \2482 , \2283_nR101a , \1378 );
and \U$1787 ( \2483 , \1371 , \2407_nRf3e );
nand \U$1788 ( \2484 , \2283_nR101a , \1369 );
or \U$1789 ( \2485 , \1334 , \2407_nRf3e );
nand \U$1790 ( \2486 , \2485 , \1374 );
and \U$1791 ( \2487 , \2484 , \2486 );
nor \U$1792 ( \2488 , \2482 , \2483 , \2487 );
xnor \U$1793 ( \2489 , \2481 , \2488 );
xor \U$1794 ( \2490 , \2371 , \2376 );
xor \U$1795 ( \2491 , \2490 , \2416 );
and \U$1796 ( \2492 , \2489 , \2491 );
and \U$1797 ( \2493 , \1761_nR13ee , \1686 );
or \U$1798 ( \2494 , \1676 , \1626_nR14f1 );
nand \U$1799 ( \2495 , \2494 , \1843 );
nand \U$1800 ( \2496 , \1761_nR13ee , \1684 );
and \U$1801 ( \2497 , \2495 , \2496 );
and \U$1802 ( \2498 , \1626_nR14f1 , \1847 );
nor \U$1803 ( \2499 , \2493 , \2497 , \2498 );
nand \U$1804 ( \2500 , \1578_nR1611 , \1970 );
or \U$1805 ( \2501 , \1856 , \1494_nR16fe );
nand \U$1806 ( \2502 , \2501 , \2144 );
and \U$1807 ( \2503 , \2500 , \2502 );
and \U$1808 ( \2504 , \2147 , \1494_nR16fe );
and \U$1809 ( \2505 , \1578_nR1611 , \1972 );
nor \U$1810 ( \2506 , \2503 , \2504 , \2505 );
xor \U$1811 ( \2507 , \2499 , \2506 );
nand \U$1812 ( \2508 , \1728_nR12de , \1631 );
or \U$1813 ( \2509 , \1507 , \1907_nR1200 );
nand \U$1814 ( \2510 , \2509 , \1637 );
and \U$1815 ( \2511 , \2508 , \2510 );
and \U$1816 ( \2512 , \1633 , \1907_nR1200 );
and \U$1817 ( \2513 , \1728_nR12de , \1660 );
nor \U$1818 ( \2514 , \2511 , \2512 , \2513 );
and \U$1819 ( \2515 , \2507 , \2514 );
and \U$1820 ( \2516 , \2499 , \2506 );
or \U$1821 ( \2517 , \2515 , \2516 );
nand \U$1822 ( \2518 , \1423_nR183c , \2209 );
or \U$1823 ( \2519 , \2167 , \1321_nR1933 );
nand \U$1824 ( \2520 , \2519 , \2350 );
and \U$1825 ( \2521 , \2518 , \2520 );
and \U$1826 ( \2522 , \2353 , \1321_nR1933 );
and \U$1827 ( \2523 , \1423_nR183c , \2211 );
nor \U$1828 ( \2524 , \2521 , \2522 , \2523 );
not \U$1829 ( \2525 , \2524 );
or \U$1830 ( \2526 , \2163 , \1364_nR1a4f );
or \U$1831 ( \2527 , \1191 , \1190_nR9e5 );
nand \U$1832 ( \2528 , \2527 , \1192 );
nor \U$1833 ( \2529 , \2163 , \2528 );
not \U$1834 ( \2530 , \2529 );
nand \U$1835 ( \2531 , \2164 , \2530 );
nand \U$1836 ( \2532 , \2526 , \2531 );
nand \U$1837 ( \2533 , \2525 , \2532 );
xor \U$1838 ( \2534 , \2517 , \2533 );
nand \U$1839 ( \2535 , \2132_nR10f9 , \1432 );
or \U$1840 ( \2536 , \1392 , \2283_nR101a );
nand \U$1841 ( \2537 , \2536 , \1437 );
and \U$1842 ( \2538 , \2535 , \2537 );
and \U$1843 ( \2539 , \1434 , \2283_nR101a );
and \U$1844 ( \2540 , \2132_nR10f9 , \1461 );
nor \U$1845 ( \2541 , \2538 , \2539 , \2540 );
and \U$1846 ( \2542 , RIb557b00_459, \1299 );
and \U$1847 ( \2543 , RIb557830_453, \1310 );
and \U$1848 ( \2544 , RIb557ce0_463, \1285 );
and \U$1849 ( \2545 , RIb557bf0_461, \1276 );
and \U$1850 ( \2546 , \1297 , RIb557b78_460);
and \U$1851 ( \2547 , RIb557c68_462, \1274 );
nor \U$1852 ( \2548 , \2546 , \2547 );
not \U$1853 ( \2549 , \2548 );
nor \U$1854 ( \2550 , \2544 , \2545 , \2549 );
and \U$1855 ( \2551 , \1312 , RIb557a88_458);
and \U$1856 ( \2552 , RIb557a10_457, \1292 );
nor \U$1857 ( \2553 , \2551 , \2552 );
nand \U$1858 ( \2554 , RIb557f38_468, \1269 );
and \U$1859 ( \2555 , \1283 , RIb557d58_464);
and \U$1860 ( \2556 , RIb557dd0_465, \1265 );
nor \U$1861 ( \2557 , \2555 , \2556 );
nand \U$1862 ( \2558 , \2550 , \2553 , \2554 , \2557 );
nor \U$1863 ( \2559 , \2542 , \2543 , \2558 );
and \U$1864 ( \2560 , \1303 , RIb557998_456);
and \U$1865 ( \2561 , RIb557920_455, \1305 );
nor \U$1866 ( \2562 , \2560 , \2561 );
and \U$1867 ( \2563 , \1288 , RIb5577b8_452);
and \U$1868 ( \2564 , RIb5578a8_454, \1314 );
nor \U$1869 ( \2565 , \2563 , \2564 );
and \U$1870 ( \2566 , \1280 , RIb557ec0_467);
and \U$1871 ( \2567 , RIb557e48_466, \1308 );
nor \U$1872 ( \2568 , \2566 , \2567 );
nand \U$1873 ( \2569 , \2559 , \2562 , \2565 , \2568 );
_DC rdbd ( \2570_nRdbd , \2569 , \1320 );
nand \U$1874 ( \2571 , \2570_nRdbd , \1232 );
and \U$1875 ( \2572 , \2541 , \2571 );
and \U$1876 ( \2573 , \2407_nRf3e , \1378 );
and \U$1877 ( \2574 , \1371 , \2480_nRe8d );
nand \U$1878 ( \2575 , \2407_nRf3e , \1369 );
or \U$1879 ( \2576 , \1334 , \2480_nRe8d );
nand \U$1880 ( \2577 , \2576 , \1374 );
and \U$1881 ( \2578 , \2575 , \2577 );
nor \U$1882 ( \2579 , \2573 , \2574 , \2578 );
nor \U$1883 ( \2580 , \2572 , \2579 );
not \U$1884 ( \2581 , \2580 );
and \U$1885 ( \2582 , \2534 , \2581 );
and \U$1886 ( \2583 , \2517 , \2533 );
or \U$1887 ( \2584 , \2582 , \2583 );
xor \U$1888 ( \2585 , \2371 , \2376 );
xor \U$1889 ( \2586 , \2585 , \2416 );
and \U$1890 ( \2587 , \2584 , \2586 );
and \U$1891 ( \2588 , \2489 , \2584 );
or \U$1892 ( \2589 , \2492 , \2587 , \2588 );
not \U$1893 ( \2590 , \2419 );
not \U$1894 ( \2591 , \2368 );
and \U$1895 ( \2592 , \2590 , \2591 );
and \U$1896 ( \2593 , \2419 , \2368 );
nor \U$1897 ( \2594 , \2592 , \2593 );
xor \U$1898 ( \2595 , \2589 , \2594 );
not \U$1899 ( \2596 , \2427 );
not \U$1900 ( \2597 , \2432 );
and \U$1901 ( \2598 , \2596 , \2597 );
and \U$1902 ( \2599 , \2427 , \2432 );
nor \U$1903 ( \2600 , \2598 , \2599 );
and \U$1904 ( \2601 , \2595 , \2600 );
and \U$1905 ( \2602 , \2589 , \2594 );
or \U$1906 ( \2603 , \2601 , \2602 );
not \U$1907 ( \2604 , \2297 );
not \U$1908 ( \2605 , \2252 );
and \U$1909 ( \2606 , \2604 , \2605 );
and \U$1910 ( \2607 , \2297 , \2252 );
nor \U$1911 ( \2608 , \2606 , \2607 );
nor \U$1912 ( \2609 , \2603 , \2608 );
and \U$1913 ( \2610 , \2603 , \2608 );
or \U$1914 ( \2611 , \2609 , \2610 );
not \U$1915 ( \2612 , \2611 );
not \U$1916 ( \2613 , \2435 );
nor \U$1917 ( \2614 , \2613 , \2421 );
not \U$1918 ( \2615 , \2614 );
not \U$1919 ( \2616 , \2433 );
and \U$1920 ( \2617 , \2615 , \2616 );
and \U$1921 ( \2618 , \2614 , \2433 );
nor \U$1922 ( \2619 , \2617 , \2618 );
not \U$1923 ( \2620 , \2619 );
and \U$1924 ( \2621 , \2612 , \2620 );
and \U$1925 ( \2622 , \2611 , \2619 );
nor \U$1926 ( \2623 , \2621 , \2622 );
not \U$1927 ( \2624 , \2489 );
xor \U$1928 ( \2625 , \2356 , \2164 );
xor \U$1929 ( \2626 , \2625 , \2364 );
xor \U$1930 ( \2627 , \2624 , \2626 );
xor \U$1931 ( \2628 , \2517 , \2533 );
xor \U$1932 ( \2629 , \2628 , \2581 );
and \U$1933 ( \2630 , \2627 , \2629 );
and \U$1934 ( \2631 , \2624 , \2626 );
or \U$1935 ( \2632 , \2630 , \2631 );
xor \U$1936 ( \2633 , \2329 , \2336 );
xor \U$1937 ( \2634 , \2633 , \2344 );
nand \U$1938 ( \2635 , \1494_nR16fe , \2209 );
or \U$1939 ( \2636 , \2167 , \1423_nR183c );
nand \U$1940 ( \2637 , \2636 , \2350 );
and \U$1941 ( \2638 , \2635 , \2637 );
and \U$1942 ( \2639 , \2353 , \1423_nR183c );
and \U$1943 ( \2640 , \1494_nR16fe , \2211 );
nor \U$1944 ( \2641 , \2638 , \2639 , \2640 );
not \U$1945 ( \2642 , \2531 );
and \U$1946 ( \2643 , \1366 , \2642 );
and \U$1947 ( \2644 , \2529 , \1322 );
nand \U$1948 ( \2645 , \2528 , \2163 );
not \U$1949 ( \2646 , \2645 );
and \U$1950 ( \2647 , \1364_nR1a4f , \2646 );
nor \U$1951 ( \2648 , \2643 , \2644 , \2647 );
xor \U$1952 ( \2649 , \2641 , \2648 );
nand \U$1953 ( \2650 , \1626_nR14f1 , \1970 );
or \U$1954 ( \2651 , \1856 , \1578_nR1611 );
nand \U$1955 ( \2652 , \2651 , \2144 );
and \U$1956 ( \2653 , \2650 , \2652 );
and \U$1957 ( \2654 , \2147 , \1578_nR1611 );
and \U$1958 ( \2655 , \1626_nR14f1 , \1972 );
nor \U$1959 ( \2656 , \2653 , \2654 , \2655 );
and \U$1960 ( \2657 , \2649 , \2656 );
and \U$1961 ( \2658 , \2641 , \2648 );
or \U$1962 ( \2659 , \2657 , \2658 );
not \U$1963 ( \2660 , \2659 );
nand \U$1964 ( \2661 , \1907_nR1200 , \1631 );
or \U$1965 ( \2662 , \1507 , \2132_nR10f9 );
nand \U$1966 ( \2663 , \2662 , \1637 );
and \U$1967 ( \2664 , \2661 , \2663 );
and \U$1968 ( \2665 , \1633 , \2132_nR10f9 );
and \U$1969 ( \2666 , \1907_nR1200 , \1660 );
nor \U$1970 ( \2667 , \2664 , \2665 , \2666 );
and \U$1971 ( \2668 , \1728_nR12de , \1686 );
or \U$1972 ( \2669 , \1676 , \1761_nR13ee );
nand \U$1973 ( \2670 , \2669 , \1843 );
nand \U$1974 ( \2671 , \1728_nR12de , \1684 );
and \U$1975 ( \2672 , \2670 , \2671 );
and \U$1976 ( \2673 , \1761_nR13ee , \1847 );
nor \U$1977 ( \2674 , \2668 , \2672 , \2673 );
xor \U$1978 ( \2675 , \2667 , \2674 );
nand \U$1979 ( \2676 , \2283_nR101a , \1432 );
or \U$1980 ( \2677 , \1392 , \2407_nRf3e );
nand \U$1981 ( \2678 , \2677 , \1437 );
and \U$1982 ( \2679 , \2676 , \2678 );
and \U$1983 ( \2680 , \1434 , \2407_nRf3e );
and \U$1984 ( \2681 , \2283_nR101a , \1461 );
nor \U$1985 ( \2682 , \2679 , \2680 , \2681 );
and \U$1986 ( \2683 , \2675 , \2682 );
and \U$1987 ( \2684 , \2667 , \2674 );
or \U$1988 ( \2685 , \2683 , \2684 );
not \U$1989 ( \2686 , \2685 );
nand \U$1990 ( \2687 , \2660 , \2686 );
xor \U$1991 ( \2688 , \2634 , \2687 );
xor \U$1992 ( \2689 , \2499 , \2506 );
xor \U$1993 ( \2690 , \2689 , \2514 );
not \U$1994 ( \2691 , \2690 );
not \U$1995 ( \2692 , \2571 );
not \U$1996 ( \2693 , \2579 );
not \U$1997 ( \2694 , \2541 );
and \U$1998 ( \2695 , \2693 , \2694 );
and \U$1999 ( \2696 , \2579 , \2541 );
nor \U$2000 ( \2697 , \2695 , \2696 );
not \U$2001 ( \2698 , \2697 );
or \U$2002 ( \2699 , \2692 , \2698 );
or \U$2003 ( \2700 , \2697 , \2571 );
nand \U$2004 ( \2701 , \2699 , \2700 );
nand \U$2005 ( \2702 , \2691 , \2701 );
and \U$2006 ( \2703 , \2688 , \2702 );
and \U$2007 ( \2704 , \2634 , \2687 );
or \U$2008 ( \2705 , \2703 , \2704 );
and \U$2009 ( \2706 , \2632 , \2705 );
xor \U$2010 ( \2707 , \2371 , \2376 );
xor \U$2011 ( \2708 , \2707 , \2416 );
xor \U$2012 ( \2709 , \2489 , \2584 );
xor \U$2013 ( \2710 , \2708 , \2709 );
not \U$2014 ( \2711 , \2710 );
not \U$2015 ( \2712 , \2367 );
or \U$2016 ( \2713 , \2347 , \2712 );
or \U$2017 ( \2714 , \2481 , \2488 );
not \U$2018 ( \2715 , \2347 );
or \U$2019 ( \2716 , \2367 , \2715 );
nand \U$2020 ( \2717 , \2713 , \2714 , \2716 );
nand \U$2021 ( \2718 , \2711 , \2717 );
xor \U$2022 ( \2719 , \2706 , \2718 );
xor \U$2023 ( \2720 , \2589 , \2594 );
xor \U$2024 ( \2721 , \2720 , \2600 );
and \U$2025 ( \2722 , \2719 , \2721 );
and \U$2026 ( \2723 , \2706 , \2718 );
nor \U$2027 ( \2724 , \2722 , \2723 );
xor \U$2028 ( \2725 , \2623 , \2724 );
not \U$2029 ( \2726 , \2710 );
not \U$2030 ( \2727 , \2717 );
and \U$2031 ( \2728 , \2726 , \2727 );
and \U$2032 ( \2729 , \2710 , \2717 );
nor \U$2033 ( \2730 , \2728 , \2729 );
xor \U$2034 ( \2731 , \2632 , \2705 );
xor \U$2035 ( \2732 , \2730 , \2731 );
xor \U$2036 ( \2733 , \2667 , \2674 );
xor \U$2037 ( \2734 , \2733 , \2682 );
not \U$2038 ( \2735 , \2734 );
and \U$2039 ( \2736 , RIb559180_507, \1303 );
and \U$2040 ( \2737 , RIb5591f8_508, \1292 );
and \U$2041 ( \2738 , RIb558fa0_503, \1288 );
and \U$2042 ( \2739 , RIb559018_504, \1310 );
and \U$2043 ( \2740 , \1305 , RIb559108_506);
and \U$2044 ( \2741 , RIb559090_505, \1314 );
nor \U$2045 ( \2742 , \2740 , \2741 );
not \U$2046 ( \2743 , \2742 );
nor \U$2047 ( \2744 , \2738 , \2739 , \2743 );
and \U$2048 ( \2745 , \1283 , RIb559540_515);
and \U$2049 ( \2746 , RIb5595b8_516, \1265 );
nor \U$2050 ( \2747 , \2745 , \2746 );
nand \U$2051 ( \2748 , RIb559720_519, \1269 );
and \U$2052 ( \2749 , \1280 , RIb5596a8_518);
and \U$2053 ( \2750 , RIb559630_517, \1308 );
nor \U$2054 ( \2751 , \2749 , \2750 );
nand \U$2055 ( \2752 , \2744 , \2747 , \2748 , \2751 );
nor \U$2056 ( \2753 , \2736 , \2737 , \2752 );
and \U$2057 ( \2754 , \1297 , RIb559360_511);
and \U$2058 ( \2755 , RIb5593d8_512, \1276 );
nor \U$2059 ( \2756 , \2754 , \2755 );
and \U$2060 ( \2757 , \1285 , RIb5594c8_514);
and \U$2061 ( \2758 , RIb559450_513, \1274 );
nor \U$2062 ( \2759 , \2757 , \2758 );
and \U$2063 ( \2760 , \1299 , RIb5592e8_510);
and \U$2064 ( \2761 , RIb559270_509, \1312 );
nor \U$2065 ( \2762 , \2760 , \2761 );
nand \U$2066 ( \2763 , \2753 , \2756 , \2759 , \2762 );
_DC rd2b ( \2764_nRd2b , \2763 , \1320 );
nand \U$2067 ( \2765 , \2764_nRd2b , \1232 );
and \U$2068 ( \2766 , \2480_nRe8d , \1378 );
and \U$2069 ( \2767 , \1371 , \2570_nRdbd );
nand \U$2070 ( \2768 , \2480_nRe8d , \1369 );
or \U$2071 ( \2769 , \1334 , \2570_nRdbd );
nand \U$2072 ( \2770 , \2769 , \1374 );
and \U$2073 ( \2771 , \2768 , \2770 );
nor \U$2074 ( \2772 , \2766 , \2767 , \2771 );
xor \U$2075 ( \2773 , \2765 , \2772 );
nand \U$2076 ( \2774 , \2735 , \2773 );
not \U$2077 ( \2775 , \2524 );
not \U$2078 ( \2776 , \2532 );
and \U$2079 ( \2777 , \2775 , \2776 );
and \U$2080 ( \2778 , \2524 , \2532 );
nor \U$2081 ( \2779 , \2777 , \2778 );
xor \U$2082 ( \2780 , \2774 , \2779 );
nand \U$2083 ( \2781 , \2407_nRf3e , \1432 );
or \U$2084 ( \2782 , \1392 , \2480_nRe8d );
nand \U$2085 ( \2783 , \2782 , \1437 );
and \U$2086 ( \2784 , \2781 , \2783 );
and \U$2087 ( \2785 , \1434 , \2480_nRe8d );
and \U$2088 ( \2786 , \2407_nRf3e , \1461 );
nor \U$2089 ( \2787 , \2784 , \2785 , \2786 );
and \U$2090 ( \2788 , \1292 , RIb558a00_491);
and \U$2091 ( \2789 , \1303 , RIb558988_490);
and \U$2092 ( \2790 , RIb558910_489, \1305 );
nor \U$2093 ( \2791 , \2789 , \2790 );
and \U$2094 ( \2792 , \1288 , RIb5587a8_486);
and \U$2095 ( \2793 , RIb558cd0_497, \1285 );
nor \U$2096 ( \2794 , \2792 , \2793 );
and \U$2097 ( \2795 , \1274 , RIb558c58_496);
and \U$2098 ( \2796 , RIb558be0_495, \1276 );
nor \U$2099 ( \2797 , \2795 , \2796 );
and \U$2100 ( \2798 , \1314 , RIb558898_488);
and \U$2101 ( \2799 , RIb558820_487, \1310 );
nor \U$2102 ( \2800 , \2798 , \2799 );
nand \U$2103 ( \2801 , \2791 , \2794 , \2797 , \2800 );
and \U$2104 ( \2802 , \1283 , RIb558d48_498);
and \U$2105 ( \2803 , RIb558dc0_499, \1265 );
nor \U$2106 ( \2804 , \2802 , \2803 );
not \U$2107 ( \2805 , \2804 );
nor \U$2108 ( \2806 , \2788 , \2801 , \2805 );
and \U$2109 ( \2807 , \1308 , RIb558e38_500);
and \U$2110 ( \2808 , RIb558a78_492, \1312 );
nor \U$2111 ( \2809 , \2807 , \2808 );
and \U$2112 ( \2810 , \1297 , RIb558b68_494);
and \U$2113 ( \2811 , RIb558af0_493, \1299 );
nor \U$2114 ( \2812 , \2810 , \2811 );
and \U$2115 ( \2813 , \1269 , RIb558f28_502);
and \U$2116 ( \2814 , RIb558eb0_501, \1280 );
nor \U$2117 ( \2815 , \2813 , \2814 );
nand \U$2118 ( \2816 , \2806 , \2809 , \2812 , \2815 );
_DC rc84 ( \2817_nRc84 , \2816 , \1320 );
nand \U$2119 ( \2818 , \2817_nRc84 , \1232 );
and \U$2120 ( \2819 , \2787 , \2818 );
and \U$2121 ( \2820 , \2570_nRdbd , \1378 );
and \U$2122 ( \2821 , \1371 , \2764_nRd2b );
nand \U$2123 ( \2822 , \2570_nRdbd , \1369 );
or \U$2124 ( \2823 , \1334 , \2764_nRd2b );
nand \U$2125 ( \2824 , \2823 , \1374 );
and \U$2126 ( \2825 , \2822 , \2824 );
nor \U$2127 ( \2826 , \2820 , \2821 , \2825 );
nor \U$2128 ( \2827 , \2819 , \2826 );
not \U$2129 ( \2828 , \2827 );
and \U$2130 ( \2829 , \1907_nR1200 , \1686 );
or \U$2131 ( \2830 , \1676 , \1728_nR12de );
nand \U$2132 ( \2831 , \2830 , \1843 );
nand \U$2133 ( \2832 , \1907_nR1200 , \1684 );
and \U$2134 ( \2833 , \2831 , \2832 );
and \U$2135 ( \2834 , \1728_nR12de , \1847 );
nor \U$2136 ( \2835 , \2829 , \2833 , \2834 );
nand \U$2137 ( \2836 , \1761_nR13ee , \1970 );
or \U$2138 ( \2837 , \1856 , \1626_nR14f1 );
nand \U$2139 ( \2838 , \2837 , \2144 );
and \U$2140 ( \2839 , \2836 , \2838 );
and \U$2141 ( \2840 , \2147 , \1626_nR14f1 );
and \U$2142 ( \2841 , \1761_nR13ee , \1972 );
nor \U$2143 ( \2842 , \2839 , \2840 , \2841 );
xor \U$2144 ( \2843 , \2835 , \2842 );
nand \U$2145 ( \2844 , \2132_nR10f9 , \1631 );
or \U$2146 ( \2845 , \1507 , \2283_nR101a );
nand \U$2147 ( \2846 , \2845 , \1637 );
and \U$2148 ( \2847 , \2844 , \2846 );
and \U$2149 ( \2848 , \1633 , \2283_nR101a );
and \U$2150 ( \2849 , \2132_nR10f9 , \1660 );
nor \U$2151 ( \2850 , \2847 , \2848 , \2849 );
and \U$2152 ( \2851 , \2843 , \2850 );
and \U$2153 ( \2852 , \2835 , \2842 );
or \U$2154 ( \2853 , \2851 , \2852 );
nand \U$2155 ( \2854 , \2828 , \2853 );
or \U$2156 ( \2855 , \2645 , \1322 );
or \U$2157 ( \2856 , \1321_nR1933 , \2531 );
or \U$2158 ( \2857 , \1423_nR183c , \2530 );
nand \U$2159 ( \2858 , \2855 , \2856 , \2857 );
not \U$2160 ( \2859 , \2858 );
nand \U$2161 ( \2860 , \1578_nR1611 , \2209 );
or \U$2162 ( \2861 , \2167 , \1494_nR16fe );
nand \U$2163 ( \2862 , \2861 , \2350 );
and \U$2164 ( \2863 , \2860 , \2862 );
and \U$2165 ( \2864 , \2353 , \1494_nR16fe );
and \U$2166 ( \2865 , \1578_nR1611 , \2211 );
nor \U$2167 ( \2866 , \2863 , \2864 , \2865 );
nor \U$2168 ( \2867 , \2859 , \2866 );
and \U$2169 ( \2868 , \2854 , \2867 );
not \U$2170 ( \2869 , \2827 );
nor \U$2171 ( \2870 , \2869 , \2853 );
nor \U$2172 ( \2871 , \2868 , \2870 );
and \U$2173 ( \2872 , \2780 , \2871 );
and \U$2174 ( \2873 , \2774 , \2779 );
or \U$2175 ( \2874 , \2872 , \2873 );
not \U$2176 ( \2875 , \2701 );
not \U$2177 ( \2876 , \2690 );
and \U$2178 ( \2877 , \2875 , \2876 );
and \U$2179 ( \2878 , \2701 , \2690 );
nor \U$2180 ( \2879 , \2877 , \2878 );
not \U$2181 ( \2880 , \2879 );
or \U$2182 ( \2881 , \2685 , \2660 );
or \U$2183 ( \2882 , \2765 , \2772 );
or \U$2184 ( \2883 , \2659 , \2686 );
nand \U$2185 ( \2884 , \2881 , \2882 , \2883 );
nand \U$2186 ( \2885 , \2880 , \2884 );
xor \U$2187 ( \2886 , \2874 , \2885 );
xor \U$2188 ( \2887 , \2624 , \2626 );
xor \U$2189 ( \2888 , \2887 , \2629 );
and \U$2190 ( \2889 , \2886 , \2888 );
and \U$2191 ( \2890 , \2874 , \2885 );
or \U$2192 ( \2891 , \2889 , \2890 );
and \U$2193 ( \2892 , \2732 , \2891 );
and \U$2194 ( \2893 , \2730 , \2731 );
or \U$2195 ( \2894 , \2892 , \2893 );
xor \U$2196 ( \2895 , \2706 , \2718 );
xor \U$2197 ( \2896 , \2895 , \2721 );
xor \U$2198 ( \2897 , \2894 , \2896 );
not \U$2199 ( \2898 , \2879 );
not \U$2200 ( \2899 , \2884 );
and \U$2201 ( \2900 , \2898 , \2899 );
and \U$2202 ( \2901 , \2879 , \2884 );
nor \U$2203 ( \2902 , \2900 , \2901 );
xor \U$2204 ( \2903 , \2641 , \2648 );
xor \U$2205 ( \2904 , \2903 , \2656 );
not \U$2206 ( \2905 , \2904 );
nand \U$2207 ( \2906 , \2283_nR101a , \1631 );
or \U$2208 ( \2907 , \1507 , \2407_nRf3e );
nand \U$2209 ( \2908 , \2907 , \1637 );
and \U$2210 ( \2909 , \2906 , \2908 );
and \U$2211 ( \2910 , \1633 , \2407_nRf3e );
and \U$2212 ( \2911 , \2283_nR101a , \1660 );
nor \U$2213 ( \2912 , \2909 , \2910 , \2911 );
and \U$2214 ( \2913 , \2132_nR10f9 , \1686 );
or \U$2215 ( \2914 , \1676 , \1907_nR1200 );
nand \U$2216 ( \2915 , \2914 , \1843 );
nand \U$2217 ( \2916 , \2132_nR10f9 , \1684 );
and \U$2218 ( \2917 , \2915 , \2916 );
and \U$2219 ( \2918 , \1907_nR1200 , \1847 );
nor \U$2220 ( \2919 , \2913 , \2917 , \2918 );
xor \U$2221 ( \2920 , \2912 , \2919 );
nand \U$2222 ( \2921 , \2480_nRe8d , \1432 );
or \U$2223 ( \2922 , \1392 , \2570_nRdbd );
nand \U$2224 ( \2923 , \2922 , \1437 );
and \U$2225 ( \2924 , \2921 , \2923 );
and \U$2226 ( \2925 , \1434 , \2570_nRdbd );
and \U$2227 ( \2926 , \2480_nRe8d , \1461 );
nor \U$2228 ( \2927 , \2924 , \2925 , \2926 );
and \U$2229 ( \2928 , \2920 , \2927 );
and \U$2230 ( \2929 , \2912 , \2919 );
or \U$2231 ( \2930 , \2928 , \2929 );
nand \U$2232 ( \2931 , \1626_nR14f1 , \2209 );
or \U$2233 ( \2932 , \2167 , \1578_nR1611 );
nand \U$2234 ( \2933 , \2932 , \2350 );
and \U$2235 ( \2934 , \2931 , \2933 );
and \U$2236 ( \2935 , \2353 , \1578_nR1611 );
and \U$2237 ( \2936 , \1626_nR14f1 , \2211 );
nor \U$2238 ( \2937 , \2934 , \2935 , \2936 );
and \U$2239 ( \2938 , \1424 , \2642 );
not \U$2240 ( \2939 , \1494_nR16fe );
and \U$2241 ( \2940 , \2529 , \2939 );
and \U$2242 ( \2941 , \1423_nR183c , \2646 );
nor \U$2243 ( \2942 , \2938 , \2940 , \2941 );
xor \U$2244 ( \2943 , \2937 , \2942 );
nand \U$2245 ( \2944 , \1728_nR12de , \1970 );
or \U$2246 ( \2945 , \1856 , \1761_nR13ee );
nand \U$2247 ( \2946 , \2945 , \2144 );
and \U$2248 ( \2947 , \2944 , \2946 );
and \U$2249 ( \2948 , \2147 , \1761_nR13ee );
and \U$2250 ( \2949 , \1728_nR12de , \1972 );
nor \U$2251 ( \2950 , \2947 , \2948 , \2949 );
and \U$2252 ( \2951 , \2943 , \2950 );
and \U$2253 ( \2952 , \2937 , \2942 );
or \U$2254 ( \2953 , \2951 , \2952 );
nor \U$2255 ( \2954 , \2930 , \2953 );
nand \U$2256 ( \2955 , \2905 , \2954 );
xor \U$2257 ( \2956 , \2902 , \2955 );
xor \U$2258 ( \2957 , \2774 , \2779 );
xor \U$2259 ( \2958 , \2957 , \2871 );
and \U$2260 ( \2959 , \2956 , \2958 );
and \U$2261 ( \2960 , \2902 , \2955 );
or \U$2262 ( \2961 , \2959 , \2960 );
xor \U$2263 ( \2962 , \2634 , \2687 );
xor \U$2264 ( \2963 , \2962 , \2702 );
xor \U$2265 ( \2964 , \2961 , \2963 );
xor \U$2266 ( \2965 , \2874 , \2885 );
xor \U$2267 ( \2966 , \2965 , \2888 );
and \U$2268 ( \2967 , \2964 , \2966 );
and \U$2269 ( \2968 , \2961 , \2963 );
or \U$2270 ( \2969 , \2967 , \2968 );
xor \U$2271 ( \2970 , \2730 , \2731 );
xor \U$2272 ( \2971 , \2970 , \2891 );
and \U$2273 ( \2972 , \2969 , \2971 );
not \U$2274 ( \2973 , \2930 );
and \U$2275 ( \2974 , \2973 , \2953 );
and \U$2276 ( \2975 , \2764_nRd2b , \1378 );
and \U$2277 ( \2976 , \1371 , \2817_nRc84 );
nand \U$2278 ( \2977 , \2764_nRd2b , \1369 );
or \U$2279 ( \2978 , \1334 , \2817_nRc84 );
nand \U$2280 ( \2979 , \2978 , \1374 );
and \U$2281 ( \2980 , \2977 , \2979 );
nor \U$2282 ( \2981 , \2975 , \2976 , \2980 );
and \U$2283 ( \2982 , RIb55a4b8_548, \1285 );
and \U$2284 ( \2983 , RIb55a440_547, \1274 );
and \U$2285 ( \2984 , RIb55a080_539, \1314 );
and \U$2286 ( \2985 , RIb55a008_538, \1310 );
and \U$2287 ( \2986 , \1297 , RIb55a350_545);
and \U$2288 ( \2987 , RIb55a3c8_546, \1276 );
nor \U$2289 ( \2988 , \2986 , \2987 );
not \U$2290 ( \2989 , \2988 );
nor \U$2291 ( \2990 , \2984 , \2985 , \2989 );
and \U$2292 ( \2991 , \1288 , RIb559f90_537);
and \U$2293 ( \2992 , RIb55a2d8_544, \1299 );
nor \U$2294 ( \2993 , \2991 , \2992 );
nand \U$2295 ( \2994 , RIb55a710_553, \1269 );
and \U$2296 ( \2995 , \1280 , RIb55a698_552);
and \U$2297 ( \2996 , RIb55a0f8_540, \1305 );
nor \U$2298 ( \2997 , \2995 , \2996 );
nand \U$2299 ( \2998 , \2990 , \2993 , \2994 , \2997 );
nor \U$2300 ( \2999 , \2982 , \2983 , \2998 );
and \U$2301 ( \3000 , \1303 , RIb55a170_541);
and \U$2302 ( \3001 , RIb55a1e8_542, \1292 );
nor \U$2303 ( \3002 , \3000 , \3001 );
and \U$2304 ( \3003 , \1283 , RIb55a530_549);
and \U$2305 ( \3004 , RIb55a260_543, \1312 );
nor \U$2306 ( \3005 , \3003 , \3004 );
and \U$2307 ( \3006 , \1308 , RIb55a620_551);
and \U$2308 ( \3007 , RIb55a5a8_550, \1265 );
nor \U$2309 ( \3008 , \3006 , \3007 );
nand \U$2310 ( \3009 , \2999 , \3002 , \3005 , \3008 );
_DC rc05 ( \3010_nRc05 , \3009 , \1320 );
nand \U$2311 ( \3011 , \3010_nRc05 , \1232 );
or \U$2312 ( \3012 , \2981 , \3011 );
or \U$2313 ( \3013 , \2953 , \2973 );
nand \U$2314 ( \3014 , \3012 , \3013 );
nor \U$2315 ( \3015 , \2974 , \3014 );
not \U$2316 ( \3016 , \2866 );
not \U$2317 ( \3017 , \2858 );
and \U$2318 ( \3018 , \3016 , \3017 );
and \U$2319 ( \3019 , \2866 , \2858 );
nor \U$2320 ( \3020 , \3018 , \3019 );
xor \U$2321 ( \3021 , \3015 , \3020 );
not \U$2322 ( \3022 , \2826 );
not \U$2323 ( \3023 , \2787 );
and \U$2324 ( \3024 , \3022 , \3023 );
and \U$2325 ( \3025 , \2826 , \2787 );
nor \U$2326 ( \3026 , \3024 , \3025 );
not \U$2327 ( \3027 , \3026 );
not \U$2328 ( \3028 , \2818 );
and \U$2329 ( \3029 , \3027 , \3028 );
and \U$2330 ( \3030 , \3026 , \2818 );
nor \U$2331 ( \3031 , \3029 , \3030 );
and \U$2332 ( \3032 , \3021 , \3031 );
and \U$2333 ( \3033 , \3015 , \3020 );
or \U$2334 ( \3034 , \3032 , \3033 );
not \U$2335 ( \3035 , \2773 );
not \U$2336 ( \3036 , \2734 );
and \U$2337 ( \3037 , \3035 , \3036 );
and \U$2338 ( \3038 , \2773 , \2734 );
nor \U$2339 ( \3039 , \3037 , \3038 );
xor \U$2340 ( \3040 , \3034 , \3039 );
xor \U$2341 ( \3041 , \2912 , \2919 );
xor \U$2342 ( \3042 , \3041 , \2927 );
xor \U$2343 ( \3043 , \2937 , \2942 );
xor \U$2344 ( \3044 , \3043 , \2950 );
xor \U$2345 ( \3045 , \3042 , \3044 );
xnor \U$2346 ( \3046 , \3011 , \2981 );
and \U$2347 ( \3047 , \3045 , \3046 );
and \U$2348 ( \3048 , \3042 , \3044 );
or \U$2349 ( \3049 , \3047 , \3048 );
xor \U$2350 ( \3050 , \2835 , \2842 );
xor \U$2351 ( \3051 , \3050 , \2850 );
xor \U$2352 ( \3052 , \3049 , \3051 );
and \U$2353 ( \3053 , \2283_nR101a , \1686 );
or \U$2354 ( \3054 , \1676 , \2132_nR10f9 );
nand \U$2355 ( \3055 , \3054 , \1843 );
nand \U$2356 ( \3056 , \2283_nR101a , \1684 );
and \U$2357 ( \3057 , \3055 , \3056 );
and \U$2358 ( \3058 , \2132_nR10f9 , \1847 );
nor \U$2359 ( \3059 , \3053 , \3057 , \3058 );
nand \U$2360 ( \3060 , \1907_nR1200 , \1970 );
or \U$2361 ( \3061 , \1856 , \1728_nR12de );
nand \U$2362 ( \3062 , \3061 , \2144 );
and \U$2363 ( \3063 , \3060 , \3062 );
and \U$2364 ( \3064 , \2147 , \1728_nR12de );
and \U$2365 ( \3065 , \1907_nR1200 , \1972 );
nor \U$2366 ( \3066 , \3063 , \3064 , \3065 );
xor \U$2367 ( \3067 , \3059 , \3066 );
nand \U$2368 ( \3068 , \2407_nRf3e , \1631 );
or \U$2369 ( \3069 , \1507 , \2480_nRe8d );
nand \U$2370 ( \3070 , \3069 , \1637 );
and \U$2371 ( \3071 , \3068 , \3070 );
and \U$2372 ( \3072 , \1633 , \2480_nRe8d );
and \U$2373 ( \3073 , \2407_nRf3e , \1660 );
nor \U$2374 ( \3074 , \3071 , \3072 , \3073 );
and \U$2375 ( \3075 , \3067 , \3074 );
and \U$2376 ( \3076 , \3059 , \3066 );
or \U$2377 ( \3077 , \3075 , \3076 );
nand \U$2378 ( \3078 , \1761_nR13ee , \2209 );
or \U$2379 ( \3079 , \2167 , \1626_nR14f1 );
nand \U$2380 ( \3080 , \3079 , \2350 );
and \U$2381 ( \3081 , \3078 , \3080 );
and \U$2382 ( \3082 , \2353 , \1626_nR14f1 );
and \U$2383 ( \3083 , \1761_nR13ee , \2211 );
nor \U$2384 ( \3084 , \3081 , \3082 , \3083 );
not \U$2385 ( \3085 , \3084 );
or \U$2386 ( \3086 , \2645 , \2939 );
or \U$2387 ( \3087 , \1494_nR16fe , \2531 );
or \U$2388 ( \3088 , \1578_nR1611 , \2530 );
nand \U$2389 ( \3089 , \3086 , \3087 , \3088 );
nand \U$2390 ( \3090 , \3085 , \3089 );
xor \U$2391 ( \3091 , \3077 , \3090 );
nand \U$2392 ( \3092 , \2570_nRdbd , \1432 );
or \U$2393 ( \3093 , \1392 , \2764_nRd2b );
nand \U$2394 ( \3094 , \3093 , \1437 );
and \U$2395 ( \3095 , \3092 , \3094 );
and \U$2396 ( \3096 , \1434 , \2764_nRd2b );
and \U$2397 ( \3097 , \2570_nRdbd , \1461 );
nor \U$2398 ( \3098 , \3095 , \3096 , \3097 );
and \U$2399 ( \3099 , RIb559d38_532, \1283 );
and \U$2400 ( \3100 , RIb559db0_533, \1265 );
and \U$2401 ( \3101 , RIb559978_524, \1303 );
and \U$2402 ( \3102 , RIb5599f0_525, \1292 );
and \U$2403 ( \3103 , \1299 , RIb559ae0_527);
and \U$2404 ( \3104 , RIb559a68_526, \1312 );
nor \U$2405 ( \3105 , \3103 , \3104 );
not \U$2406 ( \3106 , \3105 );
nor \U$2407 ( \3107 , \3101 , \3102 , \3106 );
and \U$2408 ( \3108 , \1285 , RIb559cc0_531);
and \U$2409 ( \3109 , RIb559c48_530, \1274 );
nor \U$2410 ( \3110 , \3108 , \3109 );
nand \U$2411 ( \3111 , RIb559f18_536, \1269 );
and \U$2412 ( \3112 , \1297 , RIb559b58_528);
and \U$2413 ( \3113 , RIb559bd0_529, \1276 );
nor \U$2414 ( \3114 , \3112 , \3113 );
nand \U$2415 ( \3115 , \3107 , \3110 , \3111 , \3114 );
nor \U$2416 ( \3116 , \3099 , \3100 , \3115 );
and \U$2417 ( \3117 , \1305 , RIb559900_523);
and \U$2418 ( \3118 , RIb559888_522, \1314 );
nor \U$2419 ( \3119 , \3117 , \3118 );
and \U$2420 ( \3120 , \1288 , RIb559798_520);
and \U$2421 ( \3121 , RIb559810_521, \1310 );
nor \U$2422 ( \3122 , \3120 , \3121 );
and \U$2423 ( \3123 , \1280 , RIb559ea0_535);
and \U$2424 ( \3124 , RIb559e28_534, \1308 );
nor \U$2425 ( \3125 , \3123 , \3124 );
nand \U$2426 ( \3126 , \3116 , \3119 , \3122 , \3125 );
_DC rb78 ( \3127_nRb78 , \3126 , \1320 );
nand \U$2427 ( \3128 , \3127_nRb78 , \1232 );
and \U$2428 ( \3129 , \3098 , \3128 );
and \U$2429 ( \3130 , \2817_nRc84 , \1378 );
and \U$2430 ( \3131 , \1371 , \3010_nRc05 );
nand \U$2431 ( \3132 , \2817_nRc84 , \1369 );
or \U$2432 ( \3133 , \1334 , \3010_nRc05 );
nand \U$2433 ( \3134 , \3133 , \1374 );
and \U$2434 ( \3135 , \3132 , \3134 );
nor \U$2435 ( \3136 , \3130 , \3131 , \3135 );
nor \U$2436 ( \3137 , \3129 , \3136 );
not \U$2437 ( \3138 , \3137 );
and \U$2438 ( \3139 , \3091 , \3138 );
and \U$2439 ( \3140 , \3077 , \3090 );
or \U$2440 ( \3141 , \3139 , \3140 );
and \U$2441 ( \3142 , \3052 , \3141 );
and \U$2442 ( \3143 , \3049 , \3051 );
or \U$2443 ( \3144 , \3142 , \3143 );
and \U$2444 ( \3145 , \3040 , \3144 );
and \U$2445 ( \3146 , \3034 , \3039 );
or \U$2446 ( \3147 , \3145 , \3146 );
not \U$2447 ( \3148 , \2954 );
not \U$2448 ( \3149 , \2904 );
and \U$2449 ( \3150 , \3148 , \3149 );
and \U$2450 ( \3151 , \2954 , \2904 );
nor \U$2451 ( \3152 , \3150 , \3151 );
not \U$2452 ( \3153 , \3152 );
not \U$2453 ( \3154 , \2867 );
not \U$2454 ( \3155 , \2870 );
nand \U$2455 ( \3156 , \3155 , \2854 );
not \U$2456 ( \3157 , \3156 );
or \U$2457 ( \3158 , \3154 , \3157 );
or \U$2458 ( \3159 , \3156 , \2867 );
nand \U$2459 ( \3160 , \3158 , \3159 );
nand \U$2460 ( \3161 , \3153 , \3160 );
xor \U$2461 ( \3162 , \3147 , \3161 );
xor \U$2462 ( \3163 , \2902 , \2955 );
xor \U$2463 ( \3164 , \3163 , \2958 );
and \U$2464 ( \3165 , \3162 , \3164 );
and \U$2465 ( \3166 , \3147 , \3161 );
or \U$2466 ( \3167 , \3165 , \3166 );
xor \U$2467 ( \3168 , \2961 , \2963 );
xor \U$2468 ( \3169 , \3168 , \2966 );
and \U$2469 ( \3170 , \3167 , \3169 );
not \U$2470 ( \3171 , \3152 );
not \U$2471 ( \3172 , \3160 );
or \U$2472 ( \3173 , \3171 , \3172 );
or \U$2473 ( \3174 , \3160 , \3152 );
nand \U$2474 ( \3175 , \3173 , \3174 );
not \U$2475 ( \3176 , \3175 );
nand \U$2476 ( \3177 , \1728_nR12de , \2209 );
or \U$2477 ( \3178 , \2167 , \1761_nR13ee );
nand \U$2478 ( \3179 , \3178 , \2350 );
and \U$2479 ( \3180 , \3177 , \3179 );
and \U$2480 ( \3181 , \2353 , \1761_nR13ee );
and \U$2481 ( \3182 , \1728_nR12de , \2211 );
nor \U$2482 ( \3183 , \3180 , \3181 , \3182 );
and \U$2483 ( \3184 , \1579 , \2642 );
not \U$2484 ( \3185 , \1626_nR14f1 );
and \U$2485 ( \3186 , \2529 , \3185 );
and \U$2486 ( \3187 , \1578_nR1611 , \2646 );
nor \U$2487 ( \3188 , \3184 , \3186 , \3187 );
xor \U$2488 ( \3189 , \3183 , \3188 );
nand \U$2489 ( \3190 , \2132_nR10f9 , \1970 );
or \U$2490 ( \3191 , \1856 , \1907_nR1200 );
nand \U$2491 ( \3192 , \3191 , \2144 );
and \U$2492 ( \3193 , \3190 , \3192 );
and \U$2493 ( \3194 , \2147 , \1907_nR1200 );
and \U$2494 ( \3195 , \2132_nR10f9 , \1972 );
nor \U$2495 ( \3196 , \3193 , \3194 , \3195 );
and \U$2496 ( \3197 , \3189 , \3196 );
and \U$2497 ( \3198 , \3183 , \3188 );
or \U$2498 ( \3199 , \3197 , \3198 );
not \U$2499 ( \3200 , \3199 );
nand \U$2500 ( \3201 , \2480_nRe8d , \1631 );
or \U$2501 ( \3202 , \1507 , \2570_nRdbd );
nand \U$2502 ( \3203 , \3202 , \1637 );
and \U$2503 ( \3204 , \3201 , \3203 );
and \U$2504 ( \3205 , \1633 , \2570_nRdbd );
and \U$2505 ( \3206 , \2480_nRe8d , \1660 );
nor \U$2506 ( \3207 , \3204 , \3205 , \3206 );
and \U$2507 ( \3208 , \2407_nRf3e , \1686 );
or \U$2508 ( \3209 , \1676 , \2283_nR101a );
nand \U$2509 ( \3210 , \3209 , \1843 );
nand \U$2510 ( \3211 , \2407_nRf3e , \1684 );
and \U$2511 ( \3212 , \3210 , \3211 );
and \U$2512 ( \3213 , \2283_nR101a , \1847 );
nor \U$2513 ( \3214 , \3208 , \3212 , \3213 );
xor \U$2514 ( \3215 , \3207 , \3214 );
nand \U$2515 ( \3216 , \2764_nRd2b , \1432 );
or \U$2516 ( \3217 , \1392 , \2817_nRc84 );
nand \U$2517 ( \3218 , \3217 , \1437 );
and \U$2518 ( \3219 , \3216 , \3218 );
and \U$2519 ( \3220 , \1434 , \2817_nRc84 );
and \U$2520 ( \3221 , \2764_nRd2b , \1461 );
nor \U$2521 ( \3222 , \3219 , \3220 , \3221 );
and \U$2522 ( \3223 , \3215 , \3222 );
and \U$2523 ( \3224 , \3207 , \3214 );
or \U$2524 ( \3225 , \3223 , \3224 );
not \U$2525 ( \3226 , \3225 );
nand \U$2526 ( \3227 , \3200 , \3226 );
xor \U$2527 ( \3228 , \3042 , \3044 );
xor \U$2528 ( \3229 , \3228 , \3046 );
and \U$2529 ( \3230 , \3227 , \3229 );
xor \U$2530 ( \3231 , \3059 , \3066 );
xor \U$2531 ( \3232 , \3231 , \3074 );
not \U$2532 ( \3233 , \3232 );
not \U$2533 ( \3234 , \3128 );
not \U$2534 ( \3235 , \3136 );
not \U$2535 ( \3236 , \3098 );
and \U$2536 ( \3237 , \3235 , \3236 );
and \U$2537 ( \3238 , \3136 , \3098 );
nor \U$2538 ( \3239 , \3237 , \3238 );
not \U$2539 ( \3240 , \3239 );
or \U$2540 ( \3241 , \3234 , \3240 );
or \U$2541 ( \3242 , \3239 , \3128 );
nand \U$2542 ( \3243 , \3241 , \3242 );
nand \U$2543 ( \3244 , \3233 , \3243 );
xor \U$2544 ( \3245 , \3042 , \3044 );
xor \U$2545 ( \3246 , \3245 , \3046 );
and \U$2546 ( \3247 , \3244 , \3246 );
and \U$2547 ( \3248 , \3227 , \3244 );
or \U$2548 ( \3249 , \3230 , \3247 , \3248 );
xor \U$2549 ( \3250 , \3015 , \3020 );
xor \U$2550 ( \3251 , \3250 , \3031 );
xor \U$2551 ( \3252 , \3249 , \3251 );
xor \U$2552 ( \3253 , \3049 , \3051 );
xor \U$2553 ( \3254 , \3253 , \3141 );
and \U$2554 ( \3255 , \3252 , \3254 );
and \U$2555 ( \3256 , \3249 , \3251 );
or \U$2556 ( \3257 , \3255 , \3256 );
nand \U$2557 ( \3258 , \3176 , \3257 );
not \U$2558 ( \3259 , \3257 );
nand \U$2559 ( \3260 , \3259 , \3175 );
nand \U$2560 ( \3261 , \3258 , \3260 );
not \U$2561 ( \3262 , \3261 );
xor \U$2562 ( \3263 , \3034 , \3039 );
xor \U$2563 ( \3264 , \3263 , \3144 );
not \U$2564 ( \3265 , \3264 );
and \U$2565 ( \3266 , \3262 , \3265 );
and \U$2566 ( \3267 , \3261 , \3264 );
nor \U$2567 ( \3268 , \3266 , \3267 );
xor \U$2568 ( \3269 , \3249 , \3251 );
xor \U$2569 ( \3270 , \3269 , \3254 );
not \U$2570 ( \3271 , \3243 );
not \U$2571 ( \3272 , \3232 );
and \U$2572 ( \3273 , \3271 , \3272 );
and \U$2573 ( \3274 , \3243 , \3232 );
nor \U$2574 ( \3275 , \3273 , \3274 );
not \U$2575 ( \3276 , \3275 );
or \U$2576 ( \3277 , \3225 , \3200 );
and \U$2577 ( \3278 , RIb55ab48_562, \1297 );
and \U$2578 ( \3279 , RIb55aad0_561, \1299 );
and \U$2579 ( \3280 , RIb55a968_558, \1303 );
and \U$2580 ( \3281 , RIb55a8f0_557, \1305 );
and \U$2581 ( \3282 , \1312 , RIb55aa58_560);
and \U$2582 ( \3283 , RIb55a9e0_559, \1292 );
nor \U$2583 ( \3284 , \3282 , \3283 );
not \U$2584 ( \3285 , \3284 );
nor \U$2585 ( \3286 , \3280 , \3281 , \3285 );
and \U$2586 ( \3287 , \1314 , RIb55a878_556);
and \U$2587 ( \3288 , RIb55a800_555, \1310 );
nor \U$2588 ( \3289 , \3287 , \3288 );
nand \U$2589 ( \3290 , RIb55af08_570, \1269 );
and \U$2590 ( \3291 , \1283 , RIb55ad28_566);
and \U$2591 ( \3292 , RIb55ada0_567, \1265 );
nor \U$2592 ( \3293 , \3291 , \3292 );
nand \U$2593 ( \3294 , \3286 , \3289 , \3290 , \3293 );
nor \U$2594 ( \3295 , \3278 , \3279 , \3294 );
and \U$2595 ( \3296 , \1288 , RIb55a788_554);
and \U$2596 ( \3297 , RIb55abc0_563, \1276 );
nor \U$2597 ( \3298 , \3296 , \3297 );
and \U$2598 ( \3299 , \1285 , RIb55acb0_565);
and \U$2599 ( \3300 , RIb55ac38_564, \1274 );
nor \U$2600 ( \3301 , \3299 , \3300 );
and \U$2601 ( \3302 , \1280 , RIb55ae90_569);
and \U$2602 ( \3303 , RIb55ae18_568, \1308 );
nor \U$2603 ( \3304 , \3302 , \3303 );
nand \U$2604 ( \3305 , \3295 , \3298 , \3301 , \3304 );
_DC rb1a ( \3306_nRb1a , \3305 , \1320 );
nand \U$2605 ( \3307 , \3306_nRb1a , \1232 );
and \U$2606 ( \3308 , \3010_nRc05 , \1378 );
and \U$2607 ( \3309 , \1371 , \3127_nRb78 );
nand \U$2608 ( \3310 , \3010_nRc05 , \1369 );
or \U$2609 ( \3311 , \1334 , \3127_nRb78 );
nand \U$2610 ( \3312 , \3311 , \1374 );
and \U$2611 ( \3313 , \3310 , \3312 );
nor \U$2612 ( \3314 , \3308 , \3309 , \3313 );
or \U$2613 ( \3315 , \3307 , \3314 );
or \U$2614 ( \3316 , \3199 , \3226 );
nand \U$2615 ( \3317 , \3277 , \3315 , \3316 );
nand \U$2616 ( \3318 , \3276 , \3317 );
xor \U$2617 ( \3319 , \3077 , \3090 );
xor \U$2618 ( \3320 , \3319 , \3138 );
xor \U$2619 ( \3321 , \3318 , \3320 );
xor \U$2620 ( \3322 , \3207 , \3214 );
xor \U$2621 ( \3323 , \3322 , \3222 );
xor \U$2622 ( \3324 , \3183 , \3188 );
xor \U$2623 ( \3325 , \3324 , \3196 );
xor \U$2624 ( \3326 , \3323 , \3325 );
xnor \U$2625 ( \3327 , \3307 , \3314 );
and \U$2626 ( \3328 , \3326 , \3327 );
and \U$2627 ( \3329 , \3323 , \3325 );
or \U$2628 ( \3330 , \3328 , \3329 );
not \U$2629 ( \3331 , \3084 );
not \U$2630 ( \3332 , \3089 );
and \U$2631 ( \3333 , \3331 , \3332 );
and \U$2632 ( \3334 , \3084 , \3089 );
nor \U$2633 ( \3335 , \3333 , \3334 );
xor \U$2634 ( \3336 , \3330 , \3335 );
and \U$2635 ( \3337 , \2480_nRe8d , \1686 );
or \U$2636 ( \3338 , \1676 , \2407_nRf3e );
nand \U$2637 ( \3339 , \3338 , \1843 );
nand \U$2638 ( \3340 , \2480_nRe8d , \1684 );
and \U$2639 ( \3341 , \3339 , \3340 );
and \U$2640 ( \3342 , \2407_nRf3e , \1847 );
nor \U$2641 ( \3343 , \3337 , \3341 , \3342 );
nand \U$2642 ( \3344 , \2283_nR101a , \1970 );
or \U$2643 ( \3345 , \1856 , \2132_nR10f9 );
nand \U$2644 ( \3346 , \3345 , \2144 );
and \U$2645 ( \3347 , \3344 , \3346 );
and \U$2646 ( \3348 , \2147 , \2132_nR10f9 );
and \U$2647 ( \3349 , \2283_nR101a , \1972 );
nor \U$2648 ( \3350 , \3347 , \3348 , \3349 );
xor \U$2649 ( \3351 , \3343 , \3350 );
nand \U$2650 ( \3352 , \2570_nRdbd , \1631 );
or \U$2651 ( \3353 , \1507 , \2764_nRd2b );
nand \U$2652 ( \3354 , \3353 , \1637 );
and \U$2653 ( \3355 , \3352 , \3354 );
and \U$2654 ( \3356 , \1633 , \2764_nRd2b );
and \U$2655 ( \3357 , \2570_nRdbd , \1660 );
nor \U$2656 ( \3358 , \3355 , \3356 , \3357 );
and \U$2657 ( \3359 , \3351 , \3358 );
and \U$2658 ( \3360 , \3343 , \3350 );
or \U$2659 ( \3361 , \3359 , \3360 );
nand \U$2660 ( \3362 , \1907_nR1200 , \2209 );
or \U$2661 ( \3363 , \2167 , \1728_nR12de );
nand \U$2662 ( \3364 , \3363 , \2350 );
and \U$2663 ( \3365 , \3362 , \3364 );
and \U$2664 ( \3366 , \2353 , \1728_nR12de );
and \U$2665 ( \3367 , \1907_nR1200 , \2211 );
nor \U$2666 ( \3368 , \3365 , \3366 , \3367 );
not \U$2667 ( \3369 , \3368 );
or \U$2668 ( \3370 , \2645 , \3185 );
or \U$2669 ( \3371 , \1626_nR14f1 , \2531 );
or \U$2670 ( \3372 , \1761_nR13ee , \2530 );
nand \U$2671 ( \3373 , \3370 , \3371 , \3372 );
nand \U$2672 ( \3374 , \3369 , \3373 );
xor \U$2673 ( \3375 , \3361 , \3374 );
nand \U$2674 ( \3376 , \2817_nRc84 , \1432 );
or \U$2675 ( \3377 , \1392 , \3010_nRc05 );
nand \U$2676 ( \3378 , \3377 , \1437 );
and \U$2677 ( \3379 , \3376 , \3378 );
and \U$2678 ( \3380 , \1434 , \3010_nRc05 );
and \U$2679 ( \3381 , \2817_nRc84 , \1461 );
nor \U$2680 ( \3382 , \3379 , \3380 , \3381 );
and \U$2681 ( \3383 , RIb55af80_571, \1288 );
and \U$2682 ( \3384 , RIb55aff8_572, \1310 );
and \U$2683 ( \3385 , RIb55b160_575, \1303 );
and \U$2684 ( \3386 , RIb55b1d8_576, \1292 );
and \U$2685 ( \3387 , \1299 , RIb55b2c8_578);
and \U$2686 ( \3388 , RIb55b250_577, \1312 );
nor \U$2687 ( \3389 , \3387 , \3388 );
not \U$2688 ( \3390 , \3389 );
nor \U$2689 ( \3391 , \3385 , \3386 , \3390 );
and \U$2690 ( \3392 , \1285 , RIb55b4a8_582);
and \U$2691 ( \3393 , RIb55b430_581, \1274 );
nor \U$2692 ( \3394 , \3392 , \3393 );
nand \U$2693 ( \3395 , RIb55b700_587, \1269 );
and \U$2694 ( \3396 , \1297 , RIb55b340_579);
and \U$2695 ( \3397 , RIb55b3b8_580, \1276 );
nor \U$2696 ( \3398 , \3396 , \3397 );
nand \U$2697 ( \3399 , \3391 , \3394 , \3395 , \3398 );
nor \U$2698 ( \3400 , \3383 , \3384 , \3399 );
and \U$2699 ( \3401 , \1283 , RIb55b520_583);
and \U$2700 ( \3402 , RIb55b598_584, \1265 );
nor \U$2701 ( \3403 , \3401 , \3402 );
and \U$2702 ( \3404 , \1305 , RIb55b0e8_574);
and \U$2703 ( \3405 , RIb55b070_573, \1314 );
nor \U$2704 ( \3406 , \3404 , \3405 );
and \U$2705 ( \3407 , \1280 , RIb55b688_586);
and \U$2706 ( \3408 , RIb55b610_585, \1308 );
nor \U$2707 ( \3409 , \3407 , \3408 );
nand \U$2708 ( \3410 , \3400 , \3403 , \3406 , \3409 );
_DC r9e2 ( \3411_nR9e2 , \3410 , \1320 );
nand \U$2709 ( \3412 , \3411_nR9e2 , \1232 );
and \U$2710 ( \3413 , \3382 , \3412 );
and \U$2711 ( \3414 , \3127_nRb78 , \1378 );
and \U$2712 ( \3415 , \1371 , \3306_nRb1a );
nand \U$2713 ( \3416 , \3127_nRb78 , \1369 );
or \U$2714 ( \3417 , \1334 , \3306_nRb1a );
nand \U$2715 ( \3418 , \3417 , \1374 );
and \U$2716 ( \3419 , \3416 , \3418 );
nor \U$2717 ( \3420 , \3414 , \3415 , \3419 );
nor \U$2718 ( \3421 , \3413 , \3420 );
not \U$2719 ( \3422 , \3421 );
and \U$2720 ( \3423 , \3375 , \3422 );
and \U$2721 ( \3424 , \3361 , \3374 );
or \U$2722 ( \3425 , \3423 , \3424 );
and \U$2723 ( \3426 , \3336 , \3425 );
and \U$2724 ( \3427 , \3330 , \3335 );
or \U$2725 ( \3428 , \3426 , \3427 );
and \U$2726 ( \3429 , \3321 , \3428 );
and \U$2727 ( \3430 , \3318 , \3320 );
or \U$2728 ( \3431 , \3429 , \3430 );
nor \U$2729 ( \3432 , \3270 , \3431 );
xor \U$2730 ( \3433 , \3268 , \3432 );
and \U$2731 ( \3434 , \3270 , \3431 );
nor \U$2732 ( \3435 , \3434 , \3432 );
xor \U$2733 ( \3436 , \3318 , \3320 );
xor \U$2734 ( \3437 , \3436 , \3428 );
xor \U$2735 ( \3438 , \3042 , \3044 );
xor \U$2736 ( \3439 , \3438 , \3046 );
xor \U$2737 ( \3440 , \3227 , \3244 );
xor \U$2738 ( \3441 , \3439 , \3440 );
nor \U$2739 ( \3442 , \3437 , \3441 );
xor \U$2740 ( \3443 , \3435 , \3442 );
and \U$2741 ( \3444 , \3437 , \3441 );
nor \U$2742 ( \3445 , \3444 , \3442 );
xor \U$2743 ( \3446 , \3330 , \3335 );
xor \U$2744 ( \3447 , \3446 , \3425 );
not \U$2745 ( \3448 , \3275 );
not \U$2746 ( \3449 , \3317 );
and \U$2747 ( \3450 , \3448 , \3449 );
and \U$2748 ( \3451 , \3275 , \3317 );
nor \U$2749 ( \3452 , \3450 , \3451 );
xor \U$2750 ( \3453 , \3447 , \3452 );
nand \U$2751 ( \3454 , \2764_nRd2b , \1631 );
or \U$2752 ( \3455 , \1507 , \2817_nRc84 );
nand \U$2753 ( \3456 , \3455 , \1637 );
and \U$2754 ( \3457 , \3454 , \3456 );
and \U$2755 ( \3458 , \1633 , \2817_nRc84 );
and \U$2756 ( \3459 , \2764_nRd2b , \1660 );
nor \U$2757 ( \3460 , \3457 , \3458 , \3459 );
and \U$2758 ( \3461 , \2570_nRdbd , \1686 );
or \U$2759 ( \3462 , \1676 , \2480_nRe8d );
nand \U$2760 ( \3463 , \3462 , \1843 );
nand \U$2761 ( \3464 , \2570_nRdbd , \1684 );
and \U$2762 ( \3465 , \3463 , \3464 );
and \U$2763 ( \3466 , \2480_nRe8d , \1847 );
nor \U$2764 ( \3467 , \3461 , \3465 , \3466 );
xor \U$2765 ( \3468 , \3460 , \3467 );
nand \U$2766 ( \3469 , \3010_nRc05 , \1432 );
or \U$2767 ( \3470 , \1392 , \3127_nRb78 );
nand \U$2768 ( \3471 , \3470 , \1437 );
and \U$2769 ( \3472 , \3469 , \3471 );
and \U$2770 ( \3473 , \1434 , \3127_nRb78 );
and \U$2771 ( \3474 , \3010_nRc05 , \1461 );
nor \U$2772 ( \3475 , \3472 , \3473 , \3474 );
and \U$2773 ( \3476 , \3468 , \3475 );
and \U$2774 ( \3477 , \3460 , \3467 );
or \U$2775 ( \3478 , \3476 , \3477 );
nand \U$2776 ( \3479 , \2132_nR10f9 , \2209 );
or \U$2777 ( \3480 , \2167 , \1907_nR1200 );
nand \U$2778 ( \3481 , \3480 , \2350 );
and \U$2779 ( \3482 , \3479 , \3481 );
and \U$2780 ( \3483 , \2353 , \1907_nR1200 );
and \U$2781 ( \3484 , \2132_nR10f9 , \2211 );
nor \U$2782 ( \3485 , \3482 , \3483 , \3484 );
and \U$2783 ( \3486 , \1802 , \2642 );
not \U$2784 ( \3487 , \1728_nR12de );
and \U$2785 ( \3488 , \2529 , \3487 );
and \U$2786 ( \3489 , \1761_nR13ee , \2646 );
nor \U$2787 ( \3490 , \3486 , \3488 , \3489 );
xor \U$2788 ( \3491 , \3485 , \3490 );
nand \U$2789 ( \3492 , \2407_nRf3e , \1970 );
or \U$2790 ( \3493 , \1856 , \2283_nR101a );
nand \U$2791 ( \3494 , \3493 , \2144 );
and \U$2792 ( \3495 , \3492 , \3494 );
and \U$2793 ( \3496 , \2147 , \2283_nR101a );
and \U$2794 ( \3497 , \2407_nRf3e , \1972 );
nor \U$2795 ( \3498 , \3495 , \3496 , \3497 );
and \U$2796 ( \3499 , \3491 , \3498 );
and \U$2797 ( \3500 , \3485 , \3490 );
or \U$2798 ( \3501 , \3499 , \3500 );
xor \U$2799 ( \3502 , \3478 , \3501 );
not \U$2800 ( \3503 , \3420 );
not \U$2801 ( \3504 , \3382 );
and \U$2802 ( \3505 , \3503 , \3504 );
and \U$2803 ( \3506 , \3420 , \3382 );
nor \U$2804 ( \3507 , \3505 , \3506 );
not \U$2805 ( \3508 , \3507 );
not \U$2806 ( \3509 , \3412 );
and \U$2807 ( \3510 , \3508 , \3509 );
and \U$2808 ( \3511 , \3507 , \3412 );
nor \U$2809 ( \3512 , \3510 , \3511 );
and \U$2810 ( \3513 , \3502 , \3512 );
and \U$2811 ( \3514 , \3478 , \3501 );
or \U$2812 ( \3515 , \3513 , \3514 );
xor \U$2813 ( \3516 , \3343 , \3350 );
xor \U$2814 ( \3517 , \3516 , \3358 );
not \U$2815 ( \3518 , \3517 );
not \U$2816 ( \3519 , \3373 );
not \U$2817 ( \3520 , \3368 );
or \U$2818 ( \3521 , \3519 , \3520 );
or \U$2819 ( \3522 , \3368 , \3373 );
nand \U$2820 ( \3523 , \3521 , \3522 );
nand \U$2821 ( \3524 , \3518 , \3523 );
xor \U$2822 ( \3525 , \3515 , \3524 );
xor \U$2823 ( \3526 , \3323 , \3325 );
xor \U$2824 ( \3527 , \3526 , \3327 );
and \U$2825 ( \3528 , \3525 , \3527 );
and \U$2826 ( \3529 , \3515 , \3524 );
or \U$2827 ( \3530 , \3528 , \3529 );
and \U$2828 ( \3531 , \3453 , \3530 );
and \U$2829 ( \3532 , \3447 , \3452 );
or \U$2830 ( \3533 , \3531 , \3532 );
not \U$2831 ( \3534 , \3533 );
xor \U$2832 ( \3535 , \3445 , \3534 );
nand \U$2833 ( \3536 , \2283_nR101a , \2209 );
or \U$2834 ( \3537 , \2167 , \2132_nR10f9 );
nand \U$2835 ( \3538 , \3537 , \2350 );
and \U$2836 ( \3539 , \3536 , \3538 );
and \U$2837 ( \3540 , \2353 , \2132_nR10f9 );
and \U$2838 ( \3541 , \2283_nR101a , \2211 );
nor \U$2839 ( \3542 , \3539 , \3540 , \3541 );
and \U$2840 ( \3543 , \3487 , \2642 );
not \U$2841 ( \3544 , \1907_nR1200 );
and \U$2842 ( \3545 , \2529 , \3544 );
and \U$2843 ( \3546 , \1728_nR12de , \2646 );
nor \U$2844 ( \3547 , \3543 , \3545 , \3546 );
xor \U$2845 ( \3548 , \3542 , \3547 );
and \U$2846 ( \3549 , \3548 , \1334 );
and \U$2847 ( \3550 , \3542 , \3547 );
or \U$2848 ( \3551 , \3549 , \3550 );
and \U$2849 ( \3552 , \2764_nRd2b , \1686 );
or \U$2850 ( \3553 , \1676 , \2570_nRdbd );
nand \U$2851 ( \3554 , \3553 , \1843 );
nand \U$2852 ( \3555 , \2764_nRd2b , \1684 );
and \U$2853 ( \3556 , \3554 , \3555 );
and \U$2854 ( \3557 , \2570_nRdbd , \1847 );
nor \U$2855 ( \3558 , \3552 , \3556 , \3557 );
nand \U$2856 ( \3559 , \2480_nRe8d , \1970 );
or \U$2857 ( \3560 , \1856 , \2407_nRf3e );
nand \U$2858 ( \3561 , \3560 , \2144 );
and \U$2859 ( \3562 , \3559 , \3561 );
and \U$2860 ( \3563 , \2147 , \2407_nRf3e );
and \U$2861 ( \3564 , \2480_nRe8d , \1972 );
nor \U$2862 ( \3565 , \3562 , \3563 , \3564 );
xor \U$2863 ( \3566 , \3558 , \3565 );
nand \U$2864 ( \3567 , \2817_nRc84 , \1631 );
or \U$2865 ( \3568 , \1507 , \3010_nRc05 );
nand \U$2866 ( \3569 , \3568 , \1637 );
and \U$2867 ( \3570 , \3567 , \3569 );
and \U$2868 ( \3571 , \1633 , \3010_nRc05 );
and \U$2869 ( \3572 , \2817_nRc84 , \1660 );
nor \U$2870 ( \3573 , \3570 , \3571 , \3572 );
and \U$2871 ( \3574 , \3566 , \3573 );
and \U$2872 ( \3575 , \3558 , \3565 );
or \U$2873 ( \3576 , \3574 , \3575 );
xor \U$2874 ( \3577 , \3551 , \3576 );
and \U$2875 ( \3578 , \3306_nRb1a , \1378 );
and \U$2876 ( \3579 , \1371 , \3411_nR9e2 );
nand \U$2877 ( \3580 , \3306_nRb1a , \1369 );
or \U$2878 ( \3581 , \1334 , \3411_nR9e2 );
nand \U$2879 ( \3582 , \3581 , \1374 );
and \U$2880 ( \3583 , \3580 , \3582 );
nor \U$2881 ( \3584 , \3578 , \3579 , \3583 );
and \U$2882 ( \3585 , \3577 , \3584 );
and \U$2883 ( \3586 , \3551 , \3576 );
or \U$2884 ( \3587 , \3585 , \3586 );
not \U$2885 ( \3588 , \3517 );
not \U$2886 ( \3589 , \3523 );
and \U$2887 ( \3590 , \3588 , \3589 );
and \U$2888 ( \3591 , \3517 , \3523 );
nor \U$2889 ( \3592 , \3590 , \3591 );
xor \U$2890 ( \3593 , \3587 , \3592 );
xor \U$2891 ( \3594 , \3478 , \3501 );
xor \U$2892 ( \3595 , \3594 , \3512 );
and \U$2893 ( \3596 , \3593 , \3595 );
and \U$2894 ( \3597 , \3587 , \3592 );
or \U$2895 ( \3598 , \3596 , \3597 );
xor \U$2896 ( \3599 , \3361 , \3374 );
xor \U$2897 ( \3600 , \3599 , \3422 );
xor \U$2898 ( \3601 , \3598 , \3600 );
xor \U$2899 ( \3602 , \3515 , \3524 );
xor \U$2900 ( \3603 , \3602 , \3527 );
and \U$2901 ( \3604 , \3601 , \3603 );
and \U$2902 ( \3605 , \3598 , \3600 );
or \U$2903 ( \3606 , \3604 , \3605 );
xor \U$2904 ( \3607 , \3447 , \3452 );
xor \U$2905 ( \3608 , \3607 , \3530 );
and \U$2906 ( \3609 , \3606 , \3608 );
xor \U$2907 ( \3610 , \3551 , \3576 );
xor \U$2908 ( \3611 , \3610 , \3584 );
xor \U$2909 ( \3612 , \3485 , \3490 );
xor \U$2910 ( \3613 , \3612 , \3498 );
or \U$2911 ( \3614 , \3611 , \3613 );
nand \U$2912 ( \3615 , \3127_nRb78 , \1432 );
or \U$2913 ( \3616 , \1392 , \3306_nRb1a );
nand \U$2914 ( \3617 , \3616 , \1437 );
and \U$2915 ( \3618 , \3615 , \3617 );
and \U$2916 ( \3619 , \1434 , \3306_nRb1a );
and \U$2917 ( \3620 , \3127_nRb78 , \1461 );
nor \U$2918 ( \3621 , \3618 , \3619 , \3620 );
nand \U$2919 ( \3622 , \2407_nRf3e , \2209 );
or \U$2920 ( \3623 , \2167 , \2283_nR101a );
nand \U$2921 ( \3624 , \3623 , \2350 );
and \U$2922 ( \3625 , \3622 , \3624 );
and \U$2923 ( \3626 , \2353 , \2283_nR101a );
and \U$2924 ( \3627 , \2407_nRf3e , \2211 );
nor \U$2925 ( \3628 , \3625 , \3626 , \3627 );
and \U$2926 ( \3629 , \3544 , \2642 );
and \U$2927 ( \3630 , \2529 , \2196 );
and \U$2928 ( \3631 , \1907_nR1200 , \2646 );
nor \U$2929 ( \3632 , \3629 , \3630 , \3631 );
xor \U$2930 ( \3633 , \3628 , \3632 );
nand \U$2931 ( \3634 , \2570_nRdbd , \1970 );
or \U$2932 ( \3635 , \1856 , \2480_nRe8d );
nand \U$2933 ( \3636 , \3635 , \2144 );
and \U$2934 ( \3637 , \3634 , \3636 );
and \U$2935 ( \3638 , \2147 , \2480_nRe8d );
and \U$2936 ( \3639 , \2570_nRdbd , \1972 );
nor \U$2937 ( \3640 , \3637 , \3638 , \3639 );
and \U$2938 ( \3641 , \3633 , \3640 );
and \U$2939 ( \3642 , \3628 , \3632 );
or \U$2940 ( \3643 , \3641 , \3642 );
xor \U$2941 ( \3644 , \3621 , \3643 );
nand \U$2942 ( \3645 , \3010_nRc05 , \1631 );
or \U$2943 ( \3646 , \1507 , \3127_nRb78 );
nand \U$2944 ( \3647 , \3646 , \1637 );
and \U$2945 ( \3648 , \3645 , \3647 );
and \U$2946 ( \3649 , \1633 , \3127_nRb78 );
and \U$2947 ( \3650 , \3010_nRc05 , \1660 );
nor \U$2948 ( \3651 , \3648 , \3649 , \3650 );
and \U$2949 ( \3652 , \2817_nRc84 , \1686 );
or \U$2950 ( \3653 , \1676 , \2764_nRd2b );
nand \U$2951 ( \3654 , \3653 , \1843 );
nand \U$2952 ( \3655 , \2817_nRc84 , \1684 );
and \U$2953 ( \3656 , \3654 , \3655 );
and \U$2954 ( \3657 , \2764_nRd2b , \1847 );
nor \U$2955 ( \3658 , \3652 , \3656 , \3657 );
xor \U$2956 ( \3659 , \3651 , \3658 );
nand \U$2957 ( \3660 , \3306_nRb1a , \1432 );
or \U$2958 ( \3661 , \1392 , \3411_nR9e2 );
nand \U$2959 ( \3662 , \3661 , \1437 );
and \U$2960 ( \3663 , \3660 , \3662 );
and \U$2961 ( \3664 , \1434 , \3411_nR9e2 );
and \U$2962 ( \3665 , \3306_nRb1a , \1461 );
nor \U$2963 ( \3666 , \3663 , \3664 , \3665 );
and \U$2964 ( \3667 , \3659 , \3666 );
and \U$2965 ( \3668 , \3651 , \3658 );
or \U$2966 ( \3669 , \3667 , \3668 );
and \U$2967 ( \3670 , \3644 , \3669 );
and \U$2968 ( \3671 , \3621 , \3643 );
or \U$2969 ( \3672 , \3670 , \3671 );
xor \U$2970 ( \3673 , \3460 , \3467 );
xor \U$2971 ( \3674 , \3673 , \3475 );
xor \U$2972 ( \3675 , \3672 , \3674 );
xor \U$2973 ( \3676 , \3558 , \3565 );
xor \U$2974 ( \3677 , \3676 , \3573 );
xor \U$2975 ( \3678 , \3542 , \3547 );
xor \U$2976 ( \3679 , \3678 , \1334 );
and \U$2977 ( \3680 , \3677 , \3679 );
and \U$2978 ( \3681 , \1378 , \3411_nR9e2 );
nand \U$2979 ( \3682 , \3411_nR9e2 , \1369 );
and \U$2980 ( \3683 , \3682 , \1333 );
nor \U$2981 ( \3684 , \3681 , \3683 );
xor \U$2982 ( \3685 , \3542 , \3547 );
xor \U$2983 ( \3686 , \3685 , \1334 );
and \U$2984 ( \3687 , \3684 , \3686 );
and \U$2985 ( \3688 , \3677 , \3684 );
or \U$2986 ( \3689 , \3680 , \3687 , \3688 );
and \U$2987 ( \3690 , \3675 , \3689 );
and \U$2988 ( \3691 , \3672 , \3674 );
or \U$2989 ( \3692 , \3690 , \3691 );
xor \U$2990 ( \3693 , \3614 , \3692 );
xor \U$2991 ( \3694 , \3587 , \3592 );
xor \U$2992 ( \3695 , \3694 , \3595 );
and \U$2993 ( \3696 , \3693 , \3695 );
and \U$2994 ( \3697 , \3614 , \3692 );
or \U$2995 ( \3698 , \3696 , \3697 );
xor \U$2996 ( \3699 , \3598 , \3600 );
xor \U$2997 ( \3700 , \3699 , \3603 );
and \U$2998 ( \3701 , \3698 , \3700 );
xor \U$2999 ( \3702 , \3672 , \3674 );
xor \U$3000 ( \3703 , \3702 , \3689 );
and \U$3001 ( \3704 , \3010_nRc05 , \1686 );
or \U$3002 ( \3705 , \1676 , \2817_nRc84 );
nand \U$3003 ( \3706 , \3705 , \1843 );
nand \U$3004 ( \3707 , \3010_nRc05 , \1684 );
and \U$3005 ( \3708 , \3706 , \3707 );
and \U$3006 ( \3709 , \2817_nRc84 , \1847 );
nor \U$3007 ( \3710 , \3704 , \3708 , \3709 );
nand \U$3008 ( \3711 , \2764_nRd2b , \1970 );
or \U$3009 ( \3712 , \1856 , \2570_nRdbd );
nand \U$3010 ( \3713 , \3712 , \2144 );
and \U$3011 ( \3714 , \3711 , \3713 );
and \U$3012 ( \3715 , \2147 , \2570_nRdbd );
and \U$3013 ( \3716 , \2764_nRd2b , \1972 );
nor \U$3014 ( \3717 , \3714 , \3715 , \3716 );
xor \U$3015 ( \3718 , \3710 , \3717 );
nand \U$3016 ( \3719 , \3127_nRb78 , \1631 );
or \U$3017 ( \3720 , \1507 , \3306_nRb1a );
nand \U$3018 ( \3721 , \3720 , \1637 );
and \U$3019 ( \3722 , \3719 , \3721 );
and \U$3020 ( \3723 , \1633 , \3306_nRb1a );
and \U$3021 ( \3724 , \3127_nRb78 , \1660 );
nor \U$3022 ( \3725 , \3722 , \3723 , \3724 );
and \U$3023 ( \3726 , \3718 , \3725 );
and \U$3024 ( \3727 , \3710 , \3717 );
or \U$3025 ( \3728 , \3726 , \3727 );
nand \U$3026 ( \3729 , \2480_nRe8d , \2209 );
or \U$3027 ( \3730 , \2167 , \2407_nRf3e );
nand \U$3028 ( \3731 , \3730 , \2350 );
and \U$3029 ( \3732 , \3729 , \3731 );
and \U$3030 ( \3733 , \2353 , \2407_nRf3e );
and \U$3031 ( \3734 , \2480_nRe8d , \2211 );
nor \U$3032 ( \3735 , \3732 , \3733 , \3734 );
and \U$3033 ( \3736 , \2196 , \2642 );
not \U$3034 ( \3737 , \2283_nR101a );
and \U$3035 ( \3738 , \2529 , \3737 );
and \U$3036 ( \3739 , \2132_nR10f9 , \2646 );
nor \U$3037 ( \3740 , \3736 , \3738 , \3739 );
xor \U$3038 ( \3741 , \3735 , \3740 );
and \U$3039 ( \3742 , \3741 , \1392 );
and \U$3040 ( \3743 , \3735 , \3740 );
or \U$3041 ( \3744 , \3742 , \3743 );
xor \U$3042 ( \3745 , \3728 , \3744 );
xor \U$3043 ( \3746 , \3651 , \3658 );
xor \U$3044 ( \3747 , \3746 , \3666 );
and \U$3045 ( \3748 , \3745 , \3747 );
and \U$3046 ( \3749 , \3728 , \3744 );
or \U$3047 ( \3750 , \3748 , \3749 );
xor \U$3048 ( \3751 , \3621 , \3643 );
xor \U$3049 ( \3752 , \3751 , \3669 );
xor \U$3050 ( \3753 , \3750 , \3752 );
xor \U$3051 ( \3754 , \3542 , \3547 );
xor \U$3052 ( \3755 , \3754 , \1334 );
xor \U$3053 ( \3756 , \3677 , \3684 );
xor \U$3054 ( \3757 , \3755 , \3756 );
and \U$3055 ( \3758 , \3753 , \3757 );
and \U$3056 ( \3759 , \3750 , \3752 );
or \U$3057 ( \3760 , \3758 , \3759 );
xnor \U$3058 ( \3761 , \3613 , \3611 );
xor \U$3059 ( \3762 , \3760 , \3761 );
xor \U$3060 ( \3763 , \3703 , \3762 );
not \U$3061 ( \3764 , \3763 );
xor \U$3062 ( \3765 , \3750 , \3752 );
xor \U$3063 ( \3766 , \3765 , \3757 );
and \U$3064 ( \3767 , \1461 , \3411_nR9e2 );
nand \U$3065 ( \3768 , \3411_nR9e2 , \1432 );
and \U$3066 ( \3769 , \3768 , \1449 );
nor \U$3067 ( \3770 , \3767 , \3769 );
nand \U$3068 ( \3771 , \2570_nRdbd , \2209 );
or \U$3069 ( \3772 , \2167 , \2480_nRe8d );
nand \U$3070 ( \3773 , \3772 , \2350 );
and \U$3071 ( \3774 , \3771 , \3773 );
and \U$3072 ( \3775 , \2353 , \2480_nRe8d );
and \U$3073 ( \3776 , \2570_nRdbd , \2211 );
nor \U$3074 ( \3777 , \3774 , \3775 , \3776 );
and \U$3075 ( \3778 , \3737 , \2642 );
not \U$3076 ( \3779 , \2407_nRf3e );
and \U$3077 ( \3780 , \2529 , \3779 );
and \U$3078 ( \3781 , \2283_nR101a , \2646 );
nor \U$3079 ( \3782 , \3778 , \3780 , \3781 );
xor \U$3080 ( \3783 , \3777 , \3782 );
nand \U$3081 ( \3784 , \2817_nRc84 , \1970 );
or \U$3082 ( \3785 , \1856 , \2764_nRd2b );
nand \U$3083 ( \3786 , \3785 , \2144 );
and \U$3084 ( \3787 , \3784 , \3786 );
and \U$3085 ( \3788 , \2147 , \2764_nRd2b );
and \U$3086 ( \3789 , \2817_nRc84 , \1972 );
nor \U$3087 ( \3790 , \3787 , \3788 , \3789 );
and \U$3088 ( \3791 , \3783 , \3790 );
and \U$3089 ( \3792 , \3777 , \3782 );
or \U$3090 ( \3793 , \3791 , \3792 );
xor \U$3091 ( \3794 , \3770 , \3793 );
xor \U$3092 ( \3795 , \3710 , \3717 );
xor \U$3093 ( \3796 , \3795 , \3725 );
and \U$3094 ( \3797 , \3794 , \3796 );
and \U$3095 ( \3798 , \3770 , \3793 );
or \U$3096 ( \3799 , \3797 , \3798 );
xor \U$3097 ( \3800 , \3628 , \3632 );
xor \U$3098 ( \3801 , \3800 , \3640 );
xor \U$3099 ( \3802 , \3799 , \3801 );
xor \U$3100 ( \3803 , \3728 , \3744 );
xor \U$3101 ( \3804 , \3803 , \3747 );
and \U$3102 ( \3805 , \3802 , \3804 );
and \U$3103 ( \3806 , \3799 , \3801 );
or \U$3104 ( \3807 , \3805 , \3806 );
nor \U$3105 ( \3808 , \3766 , \3807 );
xor \U$3106 ( \3809 , \3764 , \3808 );
and \U$3107 ( \3810 , \3766 , \3807 );
nor \U$3108 ( \3811 , \3810 , \3808 );
xor \U$3109 ( \3812 , \3799 , \3801 );
xor \U$3110 ( \3813 , \3812 , \3804 );
xor \U$3111 ( \3814 , \3735 , \3740 );
xor \U$3112 ( \3815 , \3814 , \1392 );
nand \U$3113 ( \3816 , \2764_nRd2b , \2209 );
or \U$3114 ( \3817 , \2167 , \2570_nRdbd );
nand \U$3115 ( \3818 , \3817 , \2350 );
and \U$3116 ( \3819 , \3816 , \3818 );
and \U$3117 ( \3820 , \2353 , \2570_nRdbd );
and \U$3118 ( \3821 , \2764_nRd2b , \2211 );
nor \U$3119 ( \3822 , \3819 , \3820 , \3821 );
and \U$3120 ( \3823 , \3779 , \2642 );
not \U$3121 ( \3824 , \2480_nRe8d );
and \U$3122 ( \3825 , \2529 , \3824 );
and \U$3123 ( \3826 , \2407_nRf3e , \2646 );
nor \U$3124 ( \3827 , \3823 , \3825 , \3826 );
xor \U$3125 ( \3828 , \3822 , \3827 );
and \U$3126 ( \3829 , \3828 , \1507 );
and \U$3127 ( \3830 , \3822 , \3827 );
or \U$3128 ( \3831 , \3829 , \3830 );
and \U$3129 ( \3832 , \3127_nRb78 , \1686 );
or \U$3130 ( \3833 , \1676 , \3010_nRc05 );
nand \U$3131 ( \3834 , \3833 , \1843 );
nand \U$3132 ( \3835 , \3127_nRb78 , \1684 );
and \U$3133 ( \3836 , \3834 , \3835 );
and \U$3134 ( \3837 , \3010_nRc05 , \1847 );
nor \U$3135 ( \3838 , \3832 , \3836 , \3837 );
xor \U$3136 ( \3839 , \3831 , \3838 );
and \U$3137 ( \3840 , \3306_nRb1a , \1686 );
or \U$3138 ( \3841 , \1676 , \3127_nRb78 );
nand \U$3139 ( \3842 , \3841 , \1843 );
nand \U$3140 ( \3843 , \3306_nRb1a , \1684 );
and \U$3141 ( \3844 , \3842 , \3843 );
and \U$3142 ( \3845 , \3127_nRb78 , \1847 );
nor \U$3143 ( \3846 , \3840 , \3844 , \3845 );
nand \U$3144 ( \3847 , \3010_nRc05 , \1970 );
or \U$3145 ( \3848 , \1856 , \2817_nRc84 );
nand \U$3146 ( \3849 , \3848 , \2144 );
and \U$3147 ( \3850 , \3847 , \3849 );
and \U$3148 ( \3851 , \2147 , \2817_nRc84 );
and \U$3149 ( \3852 , \3010_nRc05 , \1972 );
nor \U$3150 ( \3853 , \3850 , \3851 , \3852 );
xor \U$3151 ( \3854 , \3846 , \3853 );
and \U$3152 ( \3855 , \1660 , \3411_nR9e2 );
nand \U$3153 ( \3856 , \3411_nR9e2 , \1631 );
and \U$3154 ( \3857 , \3856 , \1635 );
nor \U$3155 ( \3858 , \3855 , \3857 );
and \U$3156 ( \3859 , \3854 , \3858 );
and \U$3157 ( \3860 , \3846 , \3853 );
or \U$3158 ( \3861 , \3859 , \3860 );
and \U$3159 ( \3862 , \3839 , \3861 );
and \U$3160 ( \3863 , \3831 , \3838 );
or \U$3161 ( \3864 , \3862 , \3863 );
nand \U$3162 ( \3865 , \3815 , \3864 );
not \U$3163 ( \3866 , \3306_nRb1a );
or \U$3164 ( \3867 , \1661 , \3866 );
not \U$3165 ( \3868 , \3411_nR9e2 );
or \U$3166 ( \3869 , \3868 , \1663 );
or \U$3167 ( \3870 , \1659 , \3866 );
or \U$3168 ( \3871 , \1507 , \3411_nR9e2 );
nand \U$3169 ( \3872 , \3871 , \1637 );
nand \U$3170 ( \3873 , \3870 , \3872 );
nand \U$3171 ( \3874 , \3867 , \3869 , \3873 );
not \U$3172 ( \3875 , \3874 );
xor \U$3173 ( \3876 , \3777 , \3782 );
xor \U$3174 ( \3877 , \3876 , \3790 );
nor \U$3175 ( \3878 , \3875 , \3877 );
and \U$3176 ( \3879 , \3865 , \3878 );
nor \U$3177 ( \3880 , \3864 , \3815 );
nor \U$3178 ( \3881 , \3879 , \3880 );
nor \U$3179 ( \3882 , \3813 , \3881 );
xor \U$3180 ( \3883 , \3811 , \3882 );
not \U$3181 ( \3884 , \3878 );
not \U$3182 ( \3885 , \3880 );
nand \U$3183 ( \3886 , \3885 , \3865 );
not \U$3184 ( \3887 , \3886 );
or \U$3185 ( \3888 , \3884 , \3887 );
or \U$3186 ( \3889 , \3886 , \3878 );
nand \U$3187 ( \3890 , \3888 , \3889 );
xor \U$3188 ( \3891 , \3770 , \3793 );
xor \U$3189 ( \3892 , \3891 , \3796 );
not \U$3190 ( \3893 , \3892 );
xor \U$3191 ( \3894 , \3890 , \3893 );
not \U$3192 ( \3895 , \3874 );
not \U$3193 ( \3896 , \3877 );
and \U$3194 ( \3897 , \3895 , \3896 );
and \U$3195 ( \3898 , \3874 , \3877 );
nor \U$3196 ( \3899 , \3897 , \3898 );
not \U$3197 ( \3900 , \3899 );
xor \U$3198 ( \3901 , \3831 , \3838 );
xor \U$3199 ( \3902 , \3901 , \3861 );
nand \U$3200 ( \3903 , \2817_nRc84 , \2209 );
or \U$3201 ( \3904 , \2167 , \2764_nRd2b );
nand \U$3202 ( \3905 , \3904 , \2350 );
and \U$3203 ( \3906 , \3903 , \3905 );
and \U$3204 ( \3907 , \2353 , \2764_nRd2b );
and \U$3205 ( \3908 , \2817_nRc84 , \2211 );
nor \U$3206 ( \3909 , \3906 , \3907 , \3908 );
and \U$3207 ( \3910 , \3824 , \2642 );
not \U$3208 ( \3911 , \2570_nRdbd );
and \U$3209 ( \3912 , \2529 , \3911 );
and \U$3210 ( \3913 , \2480_nRe8d , \2646 );
nor \U$3211 ( \3914 , \3910 , \3912 , \3913 );
xor \U$3212 ( \3915 , \3909 , \3914 );
nand \U$3213 ( \3916 , \3127_nRb78 , \1970 );
or \U$3214 ( \3917 , \1856 , \3010_nRc05 );
nand \U$3215 ( \3918 , \3917 , \2144 );
and \U$3216 ( \3919 , \3916 , \3918 );
and \U$3217 ( \3920 , \2147 , \3010_nRc05 );
and \U$3218 ( \3921 , \3127_nRb78 , \1972 );
nor \U$3219 ( \3922 , \3919 , \3920 , \3921 );
and \U$3220 ( \3923 , \3915 , \3922 );
and \U$3221 ( \3924 , \3909 , \3914 );
or \U$3222 ( \3925 , \3923 , \3924 );
xor \U$3223 ( \3926 , \3822 , \3827 );
xor \U$3224 ( \3927 , \3926 , \1507 );
and \U$3225 ( \3928 , \3925 , \3927 );
xor \U$3226 ( \3929 , \3846 , \3853 );
xor \U$3227 ( \3930 , \3929 , \3858 );
xor \U$3228 ( \3931 , \3822 , \3827 );
xor \U$3229 ( \3932 , \3931 , \1507 );
and \U$3230 ( \3933 , \3930 , \3932 );
and \U$3231 ( \3934 , \3925 , \3930 );
or \U$3232 ( \3935 , \3928 , \3933 , \3934 );
or \U$3233 ( \3936 , \3902 , \3935 );
not \U$3234 ( \3937 , \3936 );
or \U$3235 ( \3938 , \3900 , \3937 );
nand \U$3236 ( \3939 , \3935 , \3902 );
nand \U$3237 ( \3940 , \3938 , \3939 );
not \U$3238 ( \3941 , \3940 );
xor \U$3239 ( \3942 , \3894 , \3941 );
nand \U$3240 ( \3943 , \3939 , \3936 );
not \U$3241 ( \3944 , \3943 );
not \U$3242 ( \3945 , \3899 );
and \U$3243 ( \3946 , \3944 , \3945 );
and \U$3244 ( \3947 , \3943 , \3899 );
nor \U$3245 ( \3948 , \3946 , \3947 );
xor \U$3246 ( \3949 , \3822 , \3827 );
xor \U$3247 ( \3950 , \3949 , \1507 );
xor \U$3248 ( \3951 , \3925 , \3930 );
xor \U$3249 ( \3952 , \3950 , \3951 );
and \U$3250 ( \3953 , \3411_nR9e2 , \1686 );
or \U$3251 ( \3954 , \1676 , \3306_nRb1a );
nand \U$3252 ( \3955 , \3954 , \1843 );
nand \U$3253 ( \3956 , \3411_nR9e2 , \1684 );
and \U$3254 ( \3957 , \3955 , \3956 );
and \U$3255 ( \3958 , \3306_nRb1a , \1847 );
nor \U$3256 ( \3959 , \3953 , \3957 , \3958 );
nand \U$3257 ( \3960 , \3010_nRc05 , \2209 );
or \U$3258 ( \3961 , \2167 , \2817_nRc84 );
nand \U$3259 ( \3962 , \3961 , \2350 );
and \U$3260 ( \3963 , \3960 , \3962 );
and \U$3261 ( \3964 , \2353 , \2817_nRc84 );
and \U$3262 ( \3965 , \3010_nRc05 , \2211 );
nor \U$3263 ( \3966 , \3963 , \3964 , \3965 );
and \U$3264 ( \3967 , \3911 , \2642 );
not \U$3265 ( \3968 , \2764_nRd2b );
and \U$3266 ( \3969 , \2529 , \3968 );
and \U$3267 ( \3970 , \2570_nRdbd , \2646 );
nor \U$3268 ( \3971 , \3967 , \3969 , \3970 );
xor \U$3269 ( \3972 , \3966 , \3971 );
and \U$3270 ( \3973 , \3972 , \1676 );
and \U$3271 ( \3974 , \3966 , \3971 );
or \U$3272 ( \3975 , \3973 , \3974 );
xor \U$3273 ( \3976 , \3959 , \3975 );
nand \U$3274 ( \3977 , \3306_nRb1a , \1970 );
or \U$3275 ( \3978 , \1856 , \3127_nRb78 );
nand \U$3276 ( \3979 , \3978 , \2144 );
and \U$3277 ( \3980 , \3977 , \3979 );
and \U$3278 ( \3981 , \2147 , \3127_nRb78 );
and \U$3279 ( \3982 , \3306_nRb1a , \1972 );
nor \U$3280 ( \3983 , \3980 , \3981 , \3982 );
not \U$3281 ( \3984 , \3983 );
or \U$3282 ( \3985 , \1980 , \3868 );
or \U$3283 ( \3986 , \3411_nR9e2 , \1676 );
nand \U$3284 ( \3987 , \3985 , \3986 , \1843 );
nand \U$3285 ( \3988 , \3984 , \3987 );
and \U$3286 ( \3989 , \3976 , \3988 );
and \U$3287 ( \3990 , \3959 , \3975 );
or \U$3288 ( \3991 , \3989 , \3990 );
nor \U$3289 ( \3992 , \3952 , \3991 );
xor \U$3290 ( \3993 , \3948 , \3992 );
not \U$3291 ( \3994 , \3983 );
not \U$3292 ( \3995 , \3987 );
or \U$3293 ( \3996 , \3994 , \3995 );
or \U$3294 ( \3997 , \3987 , \3983 );
nand \U$3295 ( \3998 , \3996 , \3997 );
not \U$3296 ( \3999 , \3998 );
nand \U$3297 ( \4000 , \3127_nRb78 , \2209 );
or \U$3298 ( \4001 , \2167 , \3010_nRc05 );
nand \U$3299 ( \4002 , \4001 , \2350 );
and \U$3300 ( \4003 , \4000 , \4002 );
and \U$3301 ( \4004 , \2353 , \3010_nRc05 );
and \U$3302 ( \4005 , \3127_nRb78 , \2211 );
nor \U$3303 ( \4006 , \4003 , \4004 , \4005 );
and \U$3304 ( \4007 , \3968 , \2642 );
not \U$3305 ( \4008 , \2817_nRc84 );
and \U$3306 ( \4009 , \2529 , \4008 );
and \U$3307 ( \4010 , \2764_nRd2b , \2646 );
nor \U$3308 ( \4011 , \4007 , \4009 , \4010 );
xor \U$3309 ( \4012 , \4006 , \4011 );
nand \U$3310 ( \4013 , \3411_nR9e2 , \1970 );
or \U$3311 ( \4014 , \1856 , \3306_nRb1a );
nand \U$3312 ( \4015 , \4014 , \2144 );
and \U$3313 ( \4016 , \4013 , \4015 );
and \U$3314 ( \4017 , \2147 , \3306_nRb1a );
and \U$3315 ( \4018 , \3411_nR9e2 , \1972 );
nor \U$3316 ( \4019 , \4016 , \4017 , \4018 );
and \U$3317 ( \4020 , \4012 , \4019 );
and \U$3318 ( \4021 , \4006 , \4011 );
or \U$3319 ( \4022 , \4020 , \4021 );
xor \U$3320 ( \4023 , \3966 , \3971 );
xor \U$3321 ( \4024 , \4023 , \1676 );
nand \U$3322 ( \4025 , \4022 , \4024 );
not \U$3323 ( \4026 , \4025 );
nor \U$3324 ( \4027 , \4024 , \4022 );
nor \U$3325 ( \4028 , \4026 , \4027 );
not \U$3326 ( \4029 , \4028 );
and \U$3327 ( \4030 , \3999 , \4029 );
and \U$3328 ( \4031 , \3998 , \4028 );
nor \U$3329 ( \4032 , \4030 , \4031 );
xor \U$3330 ( \4033 , \4006 , \4011 );
xor \U$3331 ( \4034 , \4033 , \4019 );
and \U$3332 ( \4035 , \4008 , \2642 );
not \U$3333 ( \4036 , \3010_nRc05 );
and \U$3334 ( \4037 , \2529 , \4036 );
and \U$3335 ( \4038 , \2817_nRc84 , \2646 );
nor \U$3336 ( \4039 , \4035 , \4037 , \4038 );
xor \U$3337 ( \4040 , \1856 , \4039 );
nand \U$3338 ( \4041 , \3306_nRb1a , \2209 );
or \U$3339 ( \4042 , \2167 , \3127_nRb78 );
nand \U$3340 ( \4043 , \4042 , \2350 );
and \U$3341 ( \4044 , \4041 , \4043 );
and \U$3342 ( \4045 , \2353 , \3127_nRb78 );
and \U$3343 ( \4046 , \3306_nRb1a , \2211 );
nor \U$3344 ( \4047 , \4044 , \4045 , \4046 );
and \U$3345 ( \4048 , \4040 , \4047 );
and \U$3346 ( \4049 , \1856 , \4039 );
or \U$3347 ( \4050 , \4048 , \4049 );
nor \U$3348 ( \4051 , \4034 , \4050 );
xor \U$3349 ( \4052 , \4032 , \4051 );
not \U$3350 ( \4053 , \3127_nRb78 );
or \U$3351 ( \4054 , \2645 , \4053 );
or \U$3352 ( \4055 , \3127_nRb78 , \2531 );
or \U$3353 ( \4056 , \3306_nRb1a , \2530 );
nand \U$3354 ( \4057 , \4054 , \4055 , \4056 );
xor \U$3355 ( \4058 , \4057 , \2166 );
or \U$3356 ( \4059 , \2645 , \3866 );
or \U$3357 ( \4060 , \3306_nRb1a , \2531 );
or \U$3358 ( \4061 , \3411_nR9e2 , \2530 );
nand \U$3359 ( \4062 , \4059 , \4060 , \4061 );
nand \U$3360 ( \4063 , \3411_nR9e2 , \2528 );
and \U$3361 ( \4064 , \4062 , \2164 , \4063 );
xor \U$3362 ( \4065 , \4058 , \4064 );
not \U$3363 ( \4066 , \2353 );
or \U$3364 ( \4067 , \4066 , \3868 );
or \U$3365 ( \4068 , \3411_nR9e2 , \2167 );
nand \U$3366 ( \4069 , \4067 , \4068 , \2350 );
and \U$3367 ( \4070 , \4065 , \4069 );
and \U$3368 ( \4071 , \4058 , \4064 );
or \U$3369 ( \4072 , \4070 , \4071 );
and \U$3370 ( \4073 , \4057 , \2166 );
xor \U$3371 ( \4074 , \4072 , \4073 );
nand \U$3372 ( \4075 , \3411_nR9e2 , \2209 );
or \U$3373 ( \4076 , \2167 , \3306_nRb1a );
nand \U$3374 ( \4077 , \4076 , \2350 );
and \U$3375 ( \4078 , \4075 , \4077 );
and \U$3376 ( \4079 , \2353 , \3306_nRb1a );
and \U$3377 ( \4080 , \3411_nR9e2 , \2211 );
nor \U$3378 ( \4081 , \4078 , \4079 , \4080 );
and \U$3379 ( \4082 , \4036 , \2642 );
and \U$3380 ( \4083 , \2529 , \4053 );
and \U$3381 ( \4084 , \3010_nRc05 , \2646 );
nor \U$3382 ( \4085 , \4082 , \4083 , \4084 );
and \U$3383 ( \4086 , \4081 , \4085 );
nor \U$3384 ( \4087 , \4081 , \4085 );
nor \U$3385 ( \4088 , \4086 , \4087 );
and \U$3386 ( \4089 , \4074 , \4088 );
and \U$3387 ( \4090 , \4072 , \4073 );
or \U$3388 ( \4091 , \4089 , \4090 );
xor \U$3389 ( \4092 , \4091 , \4087 );
and \U$3390 ( \4093 , \3411_nR9e2 , \2147 );
and \U$3391 ( \4094 , \3868 , \1857 );
not \U$3392 ( \4095 , \2144 );
nor \U$3393 ( \4096 , \4093 , \4094 , \4095 );
xor \U$3394 ( \4097 , \1856 , \4039 );
xor \U$3395 ( \4098 , \4097 , \4047 );
and \U$3396 ( \4099 , \4096 , \4098 );
nor \U$3397 ( \4100 , \4096 , \4098 );
nor \U$3398 ( \4101 , \4099 , \4100 );
and \U$3399 ( \4102 , \4092 , \4101 );
and \U$3400 ( \4103 , \4091 , \4087 );
or \U$3401 ( \4104 , \4102 , \4103 );
xor \U$3402 ( \4105 , \4104 , \4100 );
and \U$3403 ( \4106 , \4034 , \4050 );
nor \U$3404 ( \4107 , \4106 , \4051 );
and \U$3405 ( \4108 , \4105 , \4107 );
and \U$3406 ( \4109 , \4104 , \4100 );
or \U$3407 ( \4110 , \4108 , \4109 );
and \U$3408 ( \4111 , \4052 , \4110 );
and \U$3409 ( \4112 , \4032 , \4051 );
or \U$3410 ( \4113 , \4111 , \4112 );
or \U$3411 ( \4114 , \3998 , \4027 );
nand \U$3412 ( \4115 , \4114 , \4025 );
not \U$3413 ( \4116 , \4115 );
xor \U$3414 ( \4117 , \4113 , \4116 );
xor \U$3415 ( \4118 , \3959 , \3975 );
xor \U$3416 ( \4119 , \4118 , \3988 );
xor \U$3417 ( \4120 , \3909 , \3914 );
xor \U$3418 ( \4121 , \4120 , \3922 );
and \U$3419 ( \4122 , \4119 , \4121 );
nor \U$3420 ( \4123 , \4119 , \4121 );
nor \U$3421 ( \4124 , \4122 , \4123 );
and \U$3422 ( \4125 , \4117 , \4124 );
and \U$3423 ( \4126 , \4113 , \4116 );
or \U$3424 ( \4127 , \4125 , \4126 );
xor \U$3425 ( \4128 , \4127 , \4123 );
and \U$3426 ( \4129 , \3952 , \3991 );
nor \U$3427 ( \4130 , \4129 , \3992 );
and \U$3428 ( \4131 , \4128 , \4130 );
and \U$3429 ( \4132 , \4127 , \4123 );
or \U$3430 ( \4133 , \4131 , \4132 );
and \U$3431 ( \4134 , \3993 , \4133 );
and \U$3432 ( \4135 , \3948 , \3992 );
or \U$3433 ( \4136 , \4134 , \4135 );
and \U$3434 ( \4137 , \3942 , \4136 );
and \U$3435 ( \4138 , \3894 , \3941 );
or \U$3436 ( \4139 , \4137 , \4138 );
and \U$3437 ( \4140 , \3890 , \3893 );
xor \U$3438 ( \4141 , \4139 , \4140 );
and \U$3439 ( \4142 , \3813 , \3881 );
nor \U$3440 ( \4143 , \4142 , \3882 );
and \U$3441 ( \4144 , \4141 , \4143 );
and \U$3442 ( \4145 , \4139 , \4140 );
or \U$3443 ( \4146 , \4144 , \4145 );
and \U$3444 ( \4147 , \3883 , \4146 );
and \U$3445 ( \4148 , \3811 , \3882 );
or \U$3446 ( \4149 , \4147 , \4148 );
and \U$3447 ( \4150 , \3809 , \4149 );
and \U$3448 ( \4151 , \3764 , \3808 );
or \U$3449 ( \4152 , \4150 , \4151 );
xor \U$3450 ( \4153 , \3672 , \3674 );
xor \U$3451 ( \4154 , \4153 , \3689 );
and \U$3452 ( \4155 , \3760 , \4154 );
xor \U$3453 ( \4156 , \3672 , \3674 );
xor \U$3454 ( \4157 , \4156 , \3689 );
and \U$3455 ( \4158 , \3761 , \4157 );
and \U$3456 ( \4159 , \3760 , \3761 );
or \U$3457 ( \4160 , \4155 , \4158 , \4159 );
xor \U$3458 ( \4161 , \3614 , \3692 );
xor \U$3459 ( \4162 , \4161 , \3695 );
nand \U$3460 ( \4163 , \4160 , \4162 );
and \U$3461 ( \4164 , \4152 , \4163 );
nor \U$3462 ( \4165 , \4162 , \4160 );
nor \U$3463 ( \4166 , \4164 , \4165 );
xor \U$3464 ( \4167 , \3598 , \3600 );
xor \U$3465 ( \4168 , \4167 , \3603 );
and \U$3466 ( \4169 , \4166 , \4168 );
and \U$3467 ( \4170 , \3698 , \4166 );
or \U$3468 ( \4171 , \3701 , \4169 , \4170 );
xor \U$3469 ( \4172 , \3447 , \3452 );
xor \U$3470 ( \4173 , \4172 , \3530 );
and \U$3471 ( \4174 , \4171 , \4173 );
and \U$3472 ( \4175 , \3606 , \4171 );
or \U$3473 ( \4176 , \3609 , \4174 , \4175 );
not \U$3474 ( \4177 , \4176 );
and \U$3475 ( \4178 , \3535 , \4177 );
and \U$3476 ( \4179 , \3445 , \3534 );
or \U$3477 ( \4180 , \4178 , \4179 );
and \U$3478 ( \4181 , \3443 , \4180 );
and \U$3479 ( \4182 , \3435 , \3442 );
or \U$3480 ( \4183 , \4181 , \4182 );
and \U$3481 ( \4184 , \3433 , \4183 );
and \U$3482 ( \4185 , \3268 , \3432 );
or \U$3483 ( \4186 , \4184 , \4185 );
not \U$3484 ( \4187 , \3264 );
not \U$3485 ( \4188 , \3260 );
or \U$3486 ( \4189 , \4187 , \4188 );
nand \U$3487 ( \4190 , \4189 , \3258 );
xor \U$3488 ( \4191 , \3147 , \3161 );
xor \U$3489 ( \4192 , \4191 , \3164 );
nand \U$3490 ( \4193 , \4190 , \4192 );
and \U$3491 ( \4194 , \4186 , \4193 );
nor \U$3492 ( \4195 , \4192 , \4190 );
nor \U$3493 ( \4196 , \4194 , \4195 );
xor \U$3494 ( \4197 , \2961 , \2963 );
xor \U$3495 ( \4198 , \4197 , \2966 );
and \U$3496 ( \4199 , \4196 , \4198 );
and \U$3497 ( \4200 , \3167 , \4196 );
or \U$3498 ( \4201 , \3170 , \4199 , \4200 );
xor \U$3499 ( \4202 , \2730 , \2731 );
xor \U$3500 ( \4203 , \4202 , \2891 );
and \U$3501 ( \4204 , \4201 , \4203 );
and \U$3502 ( \4205 , \2969 , \4201 );
or \U$3503 ( \4206 , \2972 , \4204 , \4205 );
and \U$3504 ( \4207 , \2897 , \4206 );
and \U$3505 ( \4208 , \2894 , \2896 );
or \U$3506 ( \4209 , \4207 , \4208 );
not \U$3507 ( \4210 , \4209 );
and \U$3508 ( \4211 , \2725 , \4210 );
and \U$3509 ( \4212 , \2623 , \2724 );
or \U$3510 ( \4213 , \4211 , \4212 );
not \U$3511 ( \4214 , \2619 );
not \U$3512 ( \4215 , \2610 );
and \U$3513 ( \4216 , \4214 , \4215 );
nor \U$3514 ( \4217 , \4216 , \2609 );
not \U$3515 ( \4218 , \2315 );
and \U$3516 ( \4219 , \2443 , \2446 );
not \U$3517 ( \4220 , \4219 );
or \U$3518 ( \4221 , \4218 , \4220 );
or \U$3519 ( \4222 , \4219 , \2315 );
nand \U$3520 ( \4223 , \4221 , \4222 );
nand \U$3521 ( \4224 , \4217 , \4223 );
and \U$3522 ( \4225 , \4213 , \4224 );
nor \U$3523 ( \4226 , \4223 , \4217 );
nor \U$3524 ( \4227 , \4225 , \4226 );
nor \U$3525 ( \4228 , \2451 , \4227 );
nor \U$3526 ( \4229 , \2448 , \4228 );
not \U$3527 ( \4230 , \4229 );
and \U$3528 ( \4231 , \2311 , \4230 );
and \U$3529 ( \4232 , \2190 , \2310 );
or \U$3530 ( \4233 , \4231 , \4232 );
and \U$3531 ( \4234 , \2186 , \4233 );
and \U$3532 ( \4235 , \2183 , \2185 );
or \U$3533 ( \4236 , \4234 , \4235 );
and \U$3534 ( \4237 , \2070 , \4236 );
and \U$3535 ( \4238 , \1963 , \2069 );
or \U$3536 ( \4239 , \4237 , \4238 );
and \U$3537 ( \4240 , \1961 , \4239 );
and \U$3538 ( \4241 , \1840 , \1960 );
or \U$3539 ( \4242 , \4240 , \4241 );
and \U$3540 ( \4243 , \1838 , \4242 );
and \U$3541 ( \4244 , \1657 , \1837 );
or \U$3542 ( \4245 , \4243 , \4244 );
and \U$3543 ( \4246 , \1655 , \4245 );
and \U$3544 ( \4247 , \1653 , \1654 );
or \U$3545 ( \4248 , \4246 , \4247 );
not \U$3546 ( \4249 , \4248 );
or \U$3547 ( \4250 , \1541 , \4249 );
or \U$3548 ( \4251 , \4248 , \1540 );
nand \U$3549 ( \4252 , \4250 , \4251 );
not \U$3550 ( \4253 , \1238 );
and \U$3551 ( \4254 , \4253 , RIb54aa68_14);
nor \U$3552 ( \4255 , \4254 , \1255 , \1258 );
and \U$3553 ( \4256 , \4253 , RIb54a9f0_13);
and \U$3554 ( \4257 , \703 , \1240 );
nor \U$3555 ( \4258 , \4256 , \4257 );
nor \U$3556 ( \4259 , \4255 , \4258 );
not \U$3557 ( \4260 , \1247 );
or \U$3558 ( \4261 , \4253 , \729 );
nand \U$3559 ( \4262 , \4261 , RIb54aae0_15);
nand \U$3560 ( \4263 , \4260 , \4262 );
nand \U$3561 ( \4264 , \730 , \1238 );
nand \U$3562 ( \4265 , \741 , \4264 );
and \U$3563 ( \4266 , \4259 , \4263 , \4265 , \695 );
and \U$3564 ( \4267 , RIb551890_249, \4266 );
and \U$3565 ( \4268 , RIb551ea8_262, \1308 );
and \U$3566 ( \4269 , \1269 , RIb551f98_264);
and \U$3567 ( \4270 , RIb551f20_263, \1280 );
nor \U$3568 ( \4271 , \4269 , \4270 );
and \U$3569 ( \4272 , \1297 , RIb551bd8_256);
and \U$3570 ( \4273 , RIb551b60_255, \1299 );
nor \U$3571 ( \4274 , \4272 , \4273 );
and \U$3572 ( \4275 , \1274 , RIb551cc8_258);
and \U$3573 ( \4276 , RIb551c50_257, \1276 );
nor \U$3574 ( \4277 , \4275 , \4276 );
and \U$3575 ( \4278 , \1312 , RIb551ae8_254);
and \U$3576 ( \4279 , RIb551a70_253, \1292 );
nor \U$3577 ( \4280 , \4278 , \4279 );
nand \U$3578 ( \4281 , \4271 , \4274 , \4277 , \4280 );
nor \U$3579 ( \4282 , \4267 , \4268 , \4281 );
and \U$3580 ( \4283 , \1283 , RIb551db8_260);
and \U$3581 ( \4284 , RIb551e30_261, \1265 );
nor \U$3582 ( \4285 , \4283 , \4284 );
and \U$3583 ( \4286 , RIb551980_251, \1305 );
and \U$3584 ( \4287 , RIb551908_250, \1314 );
and \U$3585 ( \4288 , \1285 , RIb551d40_259);
and \U$3586 ( \4289 , RIb5519f8_252, \1303 );
nor \U$3587 ( \4290 , \4288 , \4289 );
not \U$3588 ( \4291 , \4290 );
nor \U$3589 ( \4292 , \4286 , \4287 , \4291 );
nand \U$3590 ( \4293 , \4282 , \4285 , \744 , \4292 );
buf \U$3591 ( \4294 , \4293 );
buf \U$3592 ( \4295 , \766 );
_DC r12e0 ( \4296_nR12e0 , \4294 , \4295 );
xor \U$3593 ( \4297 , \694 , \4296_nR12e0 );
and \U$3594 ( \4298 , RIb54ac48_18, \4266 );
and \U$3595 ( \4299 , RIb54b260_31, \1308 );
and \U$3596 ( \4300 , \1269 , RIb54b350_33);
and \U$3597 ( \4301 , RIb54b2d8_32, \1280 );
nor \U$3598 ( \4302 , \4300 , \4301 );
and \U$3599 ( \4303 , \1297 , RIb54af90_25);
and \U$3600 ( \4304 , RIb54af18_24, \1299 );
nor \U$3601 ( \4305 , \4303 , \4304 );
and \U$3602 ( \4306 , \1274 , RIb54b080_27);
and \U$3603 ( \4307 , RIb54b008_26, \1276 );
nor \U$3604 ( \4308 , \4306 , \4307 );
and \U$3605 ( \4309 , \1312 , RIb54aea0_23);
and \U$3606 ( \4310 , RIb54ae28_22, \1292 );
nor \U$3607 ( \4311 , \4309 , \4310 );
nand \U$3608 ( \4312 , \4302 , \4305 , \4308 , \4311 );
nor \U$3609 ( \4313 , \4298 , \4299 , \4312 );
and \U$3610 ( \4314 , \1283 , RIb54b170_29);
and \U$3611 ( \4315 , RIb54b1e8_30, \1265 );
nor \U$3612 ( \4316 , \4314 , \4315 );
and \U$3613 ( \4317 , RIb54ad38_20, \1305 );
and \U$3614 ( \4318 , RIb54acc0_19, \1314 );
and \U$3615 ( \4319 , \1285 , RIb54b0f8_28);
and \U$3616 ( \4320 , RIb54adb0_21, \1303 );
nor \U$3617 ( \4321 , \4319 , \4320 );
not \U$3618 ( \4322 , \4321 );
nor \U$3619 ( \4323 , \4317 , \4318 , \4322 );
nand \U$3620 ( \4324 , \4313 , \4316 , \790 , \4323 );
buf \U$3621 ( \4325 , \4324 );
_DC r10fd ( \4326_nR10fd , \4325 , \4295 );
xor \U$3622 ( \4327 , \774 , \4326_nR10fd );
and \U$3623 ( \4328 , RIb54b440_35, \4266 );
and \U$3624 ( \4329 , RIb54ba58_48, \1308 );
and \U$3625 ( \4330 , \1269 , RIb54bb48_50);
and \U$3626 ( \4331 , RIb54bad0_49, \1280 );
nor \U$3627 ( \4332 , \4330 , \4331 );
and \U$3628 ( \4333 , \1312 , RIb54b698_40);
and \U$3629 ( \4334 , RIb54b620_39, \1292 );
nor \U$3630 ( \4335 , \4333 , \4334 );
and \U$3631 ( \4336 , \1274 , RIb54b878_44);
and \U$3632 ( \4337 , RIb54b800_43, \1276 );
nor \U$3633 ( \4338 , \4336 , \4337 );
and \U$3634 ( \4339 , \1297 , RIb54b788_42);
and \U$3635 ( \4340 , RIb54b710_41, \1299 );
nor \U$3636 ( \4341 , \4339 , \4340 );
nand \U$3637 ( \4342 , \4332 , \4335 , \4338 , \4341 );
nor \U$3638 ( \4343 , \4328 , \4329 , \4342 );
and \U$3639 ( \4344 , \1283 , RIb54b968_46);
and \U$3640 ( \4345 , RIb54b9e0_47, \1265 );
nor \U$3641 ( \4346 , \4344 , \4345 );
and \U$3642 ( \4347 , RIb54b530_37, \1305 );
and \U$3643 ( \4348 , RIb54b4b8_36, \1314 );
and \U$3644 ( \4349 , \1285 , RIb54b8f0_45);
and \U$3645 ( \4350 , RIb54b5a8_38, \1303 );
nor \U$3646 ( \4351 , \4349 , \4350 );
not \U$3647 ( \4352 , \4351 );
nor \U$3648 ( \4353 , \4347 , \4348 , \4352 );
nand \U$3649 ( \4354 , \4343 , \4346 , \826 , \4353 );
buf \U$3650 ( \4355 , \4354 );
_DC r10fb ( \4356_nR10fb , \4355 , \4295 );
xor \U$3651 ( \4357 , \810 , \4356_nR10fb );
and \U$3652 ( \4358 , RIb54bc38_52, \4266 );
and \U$3653 ( \4359 , RIb54c250_65, \1308 );
and \U$3654 ( \4360 , \1269 , RIb54c340_67);
and \U$3655 ( \4361 , RIb54c2c8_66, \1280 );
nor \U$3656 ( \4362 , \4360 , \4361 );
and \U$3657 ( \4363 , \1312 , RIb54be90_57);
and \U$3658 ( \4364 , RIb54be18_56, \1292 );
nor \U$3659 ( \4365 , \4363 , \4364 );
and \U$3660 ( \4366 , \1274 , RIb54c070_61);
and \U$3661 ( \4367 , RIb54bff8_60, \1276 );
nor \U$3662 ( \4368 , \4366 , \4367 );
and \U$3663 ( \4369 , \1297 , RIb54bf80_59);
and \U$3664 ( \4370 , RIb54bf08_58, \1299 );
nor \U$3665 ( \4371 , \4369 , \4370 );
nand \U$3666 ( \4372 , \4362 , \4365 , \4368 , \4371 );
nor \U$3667 ( \4373 , \4358 , \4359 , \4372 );
and \U$3668 ( \4374 , \1283 , RIb54c160_63);
and \U$3669 ( \4375 , RIb54c1d8_64, \1265 );
nor \U$3670 ( \4376 , \4374 , \4375 );
and \U$3671 ( \4377 , RIb54bd28_54, \1305 );
and \U$3672 ( \4378 , RIb54bcb0_53, \1314 );
and \U$3673 ( \4379 , \1285 , RIb54c0e8_62);
and \U$3674 ( \4380 , RIb54bda0_55, \1303 );
nor \U$3675 ( \4381 , \4379 , \4380 );
not \U$3676 ( \4382 , \4381 );
nor \U$3677 ( \4383 , \4377 , \4378 , \4382 );
nand \U$3678 ( \4384 , \4373 , \4376 , \862 , \4383 );
buf \U$3679 ( \4385 , \4384 );
_DC rf42 ( \4386_nRf42 , \4385 , \4295 );
xor \U$3680 ( \4387 , \846 , \4386_nRf42 );
and \U$3681 ( \4388 , RIb54cb38_84, \1269 );
and \U$3682 ( \4389 , RIb54c610_73, \1292 );
and \U$3683 ( \4390 , \1308 , RIb54ca48_82);
and \U$3684 ( \4391 , RIb54c9d0_81, \1265 );
nor \U$3685 ( \4392 , \4390 , \4391 );
and \U$3686 ( \4393 , \1314 , RIb54c4a8_70);
and \U$3687 ( \4394 , RIb54c430_69, \4266 );
nor \U$3688 ( \4395 , \4393 , \4394 );
and \U$3689 ( \4396 , \1283 , RIb54c958_80);
and \U$3690 ( \4397 , RIb54c8e0_79, \1285 );
nor \U$3691 ( \4398 , \4396 , \4397 );
and \U$3692 ( \4399 , \1303 , RIb54c598_72);
and \U$3693 ( \4400 , RIb54c520_71, \1305 );
nor \U$3694 ( \4401 , \4399 , \4400 );
nand \U$3695 ( \4402 , \4392 , \4395 , \4398 , \4401 );
nor \U$3696 ( \4403 , \4388 , \4389 , \4402 );
and \U$3697 ( \4404 , \1280 , RIb54cac0_83);
and \U$3698 ( \4405 , RIb54c868_78, \1274 );
nor \U$3699 ( \4406 , \4404 , \4405 );
and \U$3700 ( \4407 , RIb54c700_75, \1299 );
and \U$3701 ( \4408 , RIb54c688_74, \1312 );
and \U$3702 ( \4409 , \1297 , RIb54c778_76);
and \U$3703 ( \4410 , RIb54c7f0_77, \1276 );
nor \U$3704 ( \4411 , \4409 , \4410 );
not \U$3705 ( \4412 , \4411 );
nor \U$3706 ( \4413 , \4407 , \4408 , \4412 );
nand \U$3707 ( \4414 , \4403 , \4406 , \898 , \4413 );
buf \U$3708 ( \4415 , \4414 );
_DC rf40 ( \4416_nRf40 , \4415 , \4295 );
xor \U$3709 ( \4417 , \882 , \4416_nRf40 );
and \U$3710 ( \4418 , RIb54cc28_86, \4266 );
and \U$3711 ( \4419 , RIb54d240_99, \1308 );
and \U$3712 ( \4420 , \1269 , RIb54d330_101);
and \U$3713 ( \4421 , RIb54d2b8_100, \1280 );
nor \U$3714 ( \4422 , \4420 , \4421 );
and \U$3715 ( \4423 , \1299 , RIb54cef8_92);
and \U$3716 ( \4424 , RIb54cd90_89, \1303 );
nor \U$3717 ( \4425 , \4423 , \4424 );
and \U$3718 ( \4426 , \1297 , RIb54cf70_93);
and \U$3719 ( \4427 , RIb54cfe8_94, \1276 );
nor \U$3720 ( \4428 , \4426 , \4427 );
and \U$3721 ( \4429 , \1265 , RIb54d1c8_98);
and \U$3722 ( \4430 , RIb54d060_95, \1274 );
nor \U$3723 ( \4431 , \4429 , \4430 );
nand \U$3724 ( \4432 , \4422 , \4425 , \4428 , \4431 );
nor \U$3725 ( \4433 , \4418 , \4419 , \4432 );
and \U$3726 ( \4434 , \1283 , RIb54d150_97);
and \U$3727 ( \4435 , RIb54d0d8_96, \1285 );
nor \U$3728 ( \4436 , \4434 , \4435 );
and \U$3729 ( \4437 , RIb54cd18_88, \1305 );
and \U$3730 ( \4438 , RIb54cca0_87, \1314 );
and \U$3731 ( \4439 , \1312 , RIb54ce80_91);
and \U$3732 ( \4440 , RIb54ce08_90, \1292 );
nor \U$3733 ( \4441 , \4439 , \4440 );
not \U$3734 ( \4442 , \4441 );
nor \U$3735 ( \4443 , \4437 , \4438 , \4442 );
nand \U$3736 ( \4444 , \4433 , \4436 , \934 , \4443 );
buf \U$3737 ( \4445 , \4444 );
_DC rdc1 ( \4446_nRdc1 , \4445 , \4295 );
xor \U$3738 ( \4447 , \918 , \4446_nRdc1 );
and \U$3739 ( \4448 , RIb54d420_103, \4266 );
and \U$3740 ( \4449 , RIb54da38_116, \1308 );
and \U$3741 ( \4450 , \1269 , RIb54db28_118);
and \U$3742 ( \4451 , RIb54dab0_117, \1280 );
nor \U$3743 ( \4452 , \4450 , \4451 );
and \U$3744 ( \4453 , \1297 , RIb54d768_110);
and \U$3745 ( \4454 , RIb54d6f0_109, \1299 );
nor \U$3746 ( \4455 , \4453 , \4454 );
and \U$3747 ( \4456 , \1312 , RIb54d678_108);
and \U$3748 ( \4457 , RIb54d600_107, \1292 );
nor \U$3749 ( \4458 , \4456 , \4457 );
and \U$3750 ( \4459 , \1265 , RIb54d9c0_115);
and \U$3751 ( \4460 , RIb54d858_112, \1274 );
nor \U$3752 ( \4461 , \4459 , \4460 );
nand \U$3753 ( \4462 , \4452 , \4455 , \4458 , \4461 );
nor \U$3754 ( \4463 , \4448 , \4449 , \4462 );
and \U$3755 ( \4464 , \1283 , RIb54d948_114);
and \U$3756 ( \4465 , RIb54d8d0_113, \1285 );
nor \U$3757 ( \4466 , \4464 , \4465 );
and \U$3758 ( \4467 , RIb54d510_105, \1305 );
and \U$3759 ( \4468 , RIb54d498_104, \1314 );
and \U$3760 ( \4469 , \1303 , RIb54d588_106);
and \U$3761 ( \4470 , RIb54d7e0_111, \1276 );
nor \U$3762 ( \4471 , \4469 , \4470 );
not \U$3763 ( \4472 , \4471 );
nor \U$3764 ( \4473 , \4467 , \4468 , \4472 );
nand \U$3765 ( \4474 , \4463 , \4466 , \970 , \4473 );
buf \U$3766 ( \4475 , \4474 );
_DC rdbf ( \4476_nRdbf , \4475 , \4295 );
xor \U$3767 ( \4477 , \954 , \4476_nRdbf );
and \U$3768 ( \4478 , RIb54dc18_120, \4266 );
and \U$3769 ( \4479 , RIb54e230_133, \1308 );
and \U$3770 ( \4480 , \1269 , RIb54e320_135);
and \U$3771 ( \4481 , RIb54e2a8_134, \1280 );
nor \U$3772 ( \4482 , \4480 , \4481 );
and \U$3773 ( \4483 , \1312 , RIb54de70_125);
and \U$3774 ( \4484 , RIb54ddf8_124, \1292 );
nor \U$3775 ( \4485 , \4483 , \4484 );
and \U$3776 ( \4486 , \1274 , RIb54e050_129);
and \U$3777 ( \4487 , RIb54dfd8_128, \1276 );
nor \U$3778 ( \4488 , \4486 , \4487 );
and \U$3779 ( \4489 , \1297 , RIb54df60_127);
and \U$3780 ( \4490 , RIb54dee8_126, \1299 );
nor \U$3781 ( \4491 , \4489 , \4490 );
nand \U$3782 ( \4492 , \4482 , \4485 , \4488 , \4491 );
nor \U$3783 ( \4493 , \4478 , \4479 , \4492 );
and \U$3784 ( \4494 , \1283 , RIb54e140_131);
and \U$3785 ( \4495 , RIb54e1b8_132, \1265 );
nor \U$3786 ( \4496 , \4494 , \4495 );
and \U$3787 ( \4497 , RIb54dd08_122, \1305 );
and \U$3788 ( \4498 , RIb54dc90_121, \1314 );
and \U$3789 ( \4499 , \1285 , RIb54e0c8_130);
and \U$3790 ( \4500 , RIb54dd80_123, \1303 );
nor \U$3791 ( \4501 , \4499 , \4500 );
not \U$3792 ( \4502 , \4501 );
nor \U$3793 ( \4503 , \4497 , \4498 , \4502 );
nand \U$3794 ( \4504 , \4493 , \4496 , \1006 , \4503 );
buf \U$3795 ( \4505 , \4504 );
_DC rc88 ( \4506_nRc88 , \4505 , \4295 );
xor \U$3796 ( \4507 , \990 , \4506_nRc88 );
and \U$3797 ( \4508 , RIb54eb18_152, \1269 );
and \U$3798 ( \4509 , RIb54e5f0_141, \1292 );
and \U$3799 ( \4510 , \1308 , RIb54ea28_150);
and \U$3800 ( \4511 , RIb54e9b0_149, \1265 );
nor \U$3801 ( \4512 , \4510 , \4511 );
and \U$3802 ( \4513 , \1283 , RIb54e938_148);
and \U$3803 ( \4514 , RIb54e758_144, \1297 );
nor \U$3804 ( \4515 , \4513 , \4514 );
and \U$3805 ( \4516 , \1314 , RIb54e488_138);
and \U$3806 ( \4517 , RIb54e410_137, \4266 );
nor \U$3807 ( \4518 , \4516 , \4517 );
and \U$3808 ( \4519 , \1303 , RIb54e578_140);
and \U$3809 ( \4520 , RIb54e500_139, \1305 );
nor \U$3810 ( \4521 , \4519 , \4520 );
nand \U$3811 ( \4522 , \4512 , \4515 , \4518 , \4521 );
nor \U$3812 ( \4523 , \4508 , \4509 , \4522 );
and \U$3813 ( \4524 , \1280 , RIb54eaa0_151);
and \U$3814 ( \4525 , RIb54e8c0_147, \1285 );
nor \U$3815 ( \4526 , \4524 , \4525 );
and \U$3816 ( \4527 , RIb54e6e0_143, \1299 );
and \U$3817 ( \4528 , RIb54e668_142, \1312 );
and \U$3818 ( \4529 , \1274 , RIb54e848_146);
and \U$3819 ( \4530 , RIb54e7d0_145, \1276 );
nor \U$3820 ( \4531 , \4529 , \4530 );
not \U$3821 ( \4532 , \4531 );
nor \U$3822 ( \4533 , \4527 , \4528 , \4532 );
nand \U$3823 ( \4534 , \4523 , \4526 , \1042 , \4533 );
buf \U$3824 ( \4535 , \4534 );
_DC rc86 ( \4536_nRc86 , \4535 , \4295 );
xor \U$3825 ( \4537 , \1026 , \4536_nRc86 );
and \U$3826 ( \4538 , RIb54f310_169, \1269 );
and \U$3827 ( \4539 , RIb54ede8_158, \1292 );
and \U$3828 ( \4540 , \1308 , RIb54f220_167);
and \U$3829 ( \4541 , RIb54f1a8_166, \1265 );
nor \U$3830 ( \4542 , \4540 , \4541 );
and \U$3831 ( \4543 , \1314 , RIb54ec80_155);
and \U$3832 ( \4544 , RIb54ec08_154, \4266 );
nor \U$3833 ( \4545 , \4543 , \4544 );
and \U$3834 ( \4546 , \1283 , RIb54f130_165);
and \U$3835 ( \4547 , RIb54f0b8_164, \1285 );
nor \U$3836 ( \4548 , \4546 , \4547 );
and \U$3837 ( \4549 , \1303 , RIb54ed70_157);
and \U$3838 ( \4550 , RIb54ecf8_156, \1305 );
nor \U$3839 ( \4551 , \4549 , \4550 );
nand \U$3840 ( \4552 , \4542 , \4545 , \4548 , \4551 );
nor \U$3841 ( \4553 , \4538 , \4539 , \4552 );
and \U$3842 ( \4554 , \1280 , RIb54f298_168);
and \U$3843 ( \4555 , RIb54f040_163, \1274 );
nor \U$3844 ( \4556 , \4554 , \4555 );
and \U$3845 ( \4557 , RIb54eed8_160, \1299 );
and \U$3846 ( \4558 , RIb54ee60_159, \1312 );
and \U$3847 ( \4559 , \1297 , RIb54ef50_161);
and \U$3848 ( \4560 , RIb54efc8_162, \1276 );
nor \U$3849 ( \4561 , \4559 , \4560 );
not \U$3850 ( \4562 , \4561 );
nor \U$3851 ( \4563 , \4557 , \4558 , \4562 );
nand \U$3852 ( \4564 , \4553 , \4556 , \1078 , \4563 );
buf \U$3853 ( \4565 , \4564 );
_DC rb9a ( \4566_nRb9a , \4565 , \4295 );
xor \U$3854 ( \4567 , \1062 , \4566_nRb9a );
and \U$3855 ( \4568 , RIb54f400_171, \4266 );
and \U$3856 ( \4569 , RIb54fa18_184, \1308 );
and \U$3857 ( \4570 , \1269 , RIb54fb08_186);
and \U$3858 ( \4571 , RIb54fa90_185, \1280 );
nor \U$3859 ( \4572 , \4570 , \4571 );
and \U$3860 ( \4573 , \1297 , RIb54f748_178);
and \U$3861 ( \4574 , RIb54f6d0_177, \1299 );
nor \U$3862 ( \4575 , \4573 , \4574 );
and \U$3863 ( \4576 , \1274 , RIb54f838_180);
and \U$3864 ( \4577 , RIb54f7c0_179, \1276 );
nor \U$3865 ( \4578 , \4576 , \4577 );
and \U$3866 ( \4579 , \1312 , RIb54f658_176);
and \U$3867 ( \4580 , RIb54f5e0_175, \1292 );
nor \U$3868 ( \4581 , \4579 , \4580 );
nand \U$3869 ( \4582 , \4572 , \4575 , \4578 , \4581 );
nor \U$3870 ( \4583 , \4568 , \4569 , \4582 );
and \U$3871 ( \4584 , \1283 , RIb54f928_182);
and \U$3872 ( \4585 , RIb54f9a0_183, \1265 );
nor \U$3873 ( \4586 , \4584 , \4585 );
and \U$3874 ( \4587 , RIb54f4f0_173, \1305 );
and \U$3875 ( \4588 , RIb54f478_172, \1314 );
and \U$3876 ( \4589 , \1285 , RIb54f8b0_181);
and \U$3877 ( \4590 , RIb54f568_174, \1303 );
nor \U$3878 ( \4591 , \4589 , \4590 );
not \U$3879 ( \4592 , \4591 );
nor \U$3880 ( \4593 , \4587 , \4588 , \4592 );
nand \U$3881 ( \4594 , \4583 , \4586 , \1114 , \4593 );
buf \U$3882 ( \4595 , \4594 );
_DC rb9c ( \4596_nRb9c , \4595 , \4295 );
xor \U$3883 ( \4597 , \1098 , \4596_nRb9c );
and \U$3884 ( \4598 , RIb54fbf8_188, \4266 );
and \U$3885 ( \4599 , RIb550210_201, \1308 );
and \U$3886 ( \4600 , \1269 , RIb550300_203);
and \U$3887 ( \4601 , RIb550288_202, \1280 );
nor \U$3888 ( \4602 , \4600 , \4601 );
and \U$3889 ( \4603 , \1312 , RIb54fe50_193);
and \U$3890 ( \4604 , RIb54fdd8_192, \1292 );
nor \U$3891 ( \4605 , \4603 , \4604 );
and \U$3892 ( \4606 , \1274 , RIb550030_197);
and \U$3893 ( \4607 , RIb54ffb8_196, \1276 );
nor \U$3894 ( \4608 , \4606 , \4607 );
and \U$3895 ( \4609 , \1297 , RIb54ff40_195);
and \U$3896 ( \4610 , RIb54fec8_194, \1299 );
nor \U$3897 ( \4611 , \4609 , \4610 );
nand \U$3898 ( \4612 , \4602 , \4605 , \4608 , \4611 );
nor \U$3899 ( \4613 , \4598 , \4599 , \4612 );
and \U$3900 ( \4614 , \1283 , RIb550120_199);
and \U$3901 ( \4615 , RIb550198_200, \1265 );
nor \U$3902 ( \4616 , \4614 , \4615 );
and \U$3903 ( \4617 , RIb54fce8_190, \1305 );
and \U$3904 ( \4618 , RIb54fc70_189, \1314 );
and \U$3905 ( \4619 , \1285 , RIb5500a8_198);
and \U$3906 ( \4620 , RIb54fd60_191, \1303 );
nor \U$3907 ( \4621 , \4619 , \4620 );
not \U$3908 ( \4622 , \4621 );
nor \U$3909 ( \4623 , \4617 , \4618 , \4622 );
nand \U$3910 ( \4624 , \4613 , \4616 , \1145 , \4623 );
buf \U$3911 ( \4625 , \4624 );
_DC ra38 ( \4626_nRa38 , \4625 , \4295 );
xor \U$3912 ( \4627 , RIb54a900_11, \4626_nRa38 );
and \U$3913 ( \4628 , RIb550468_206, \4266 );
and \U$3914 ( \4629 , RIb550a08_218, \1265 );
and \U$3915 ( \4630 , \1280 , RIb550af8_220);
and \U$3916 ( \4631 , RIb550a80_219, \1308 );
nor \U$3917 ( \4632 , \4630 , \4631 );
and \U$3918 ( \4633 , \1297 , RIb5507b0_213);
and \U$3919 ( \4634 , RIb550738_212, \1299 );
nor \U$3920 ( \4635 , \4633 , \4634 );
and \U$3921 ( \4636 , \1312 , RIb5506c0_211);
and \U$3922 ( \4637 , RIb550648_210, \1292 );
nor \U$3923 ( \4638 , \4636 , \4637 );
and \U$3924 ( \4639 , \1269 , RIb550b70_221);
and \U$3925 ( \4640 , RIb550828_214, \1276 );
nor \U$3926 ( \4641 , \4639 , \4640 );
nand \U$3927 ( \4642 , \4632 , \4635 , \4638 , \4641 );
nor \U$3928 ( \4643 , \4628 , \4629 , \4642 );
and \U$3929 ( \4644 , \1283 , RIb550990_217);
and \U$3930 ( \4645 , RIb550918_216, \1285 );
nor \U$3931 ( \4646 , \4644 , \4645 );
and \U$3932 ( \4647 , RIb550558_208, \1305 );
and \U$3933 ( \4648 , RIb5504e0_207, \1314 );
and \U$3934 ( \4649 , \1274 , RIb5508a0_215);
and \U$3935 ( \4650 , RIb5505d0_209, \1303 );
nor \U$3936 ( \4651 , \4649 , \4650 );
not \U$3937 ( \4652 , \4651 );
nor \U$3938 ( \4653 , \4647 , \4648 , \4652 );
nand \U$3939 ( \4654 , \4643 , \4646 , \1176 , \4653 );
buf \U$3940 ( \4655 , \4654 );
_DC ra36 ( \4656_nRa36 , \4655 , \4295 );
nand \U$3941 ( \4657 , \4656_nRa36 , \1191 );
not \U$3942 ( \4658 , \4657 );
and \U$3943 ( \4659 , \4627 , \4658 );
and \U$3944 ( \4660 , RIb54a900_11, \4626_nRa38 );
or \U$3945 ( \4661 , \4659 , \4660 );
and \U$3946 ( \4662 , \4597 , \4661 );
and \U$3947 ( \4663 , \1098 , \4596_nRb9c );
or \U$3948 ( \4664 , \4662 , \4663 );
and \U$3949 ( \4665 , \4567 , \4664 );
and \U$3950 ( \4666 , \1062 , \4566_nRb9a );
or \U$3951 ( \4667 , \4665 , \4666 );
and \U$3952 ( \4668 , \4537 , \4667 );
and \U$3953 ( \4669 , \1026 , \4536_nRc86 );
or \U$3954 ( \4670 , \4668 , \4669 );
and \U$3955 ( \4671 , \4507 , \4670 );
and \U$3956 ( \4672 , \990 , \4506_nRc88 );
or \U$3957 ( \4673 , \4671 , \4672 );
and \U$3958 ( \4674 , \4477 , \4673 );
and \U$3959 ( \4675 , \954 , \4476_nRdbf );
or \U$3960 ( \4676 , \4674 , \4675 );
and \U$3961 ( \4677 , \4447 , \4676 );
and \U$3962 ( \4678 , \918 , \4446_nRdc1 );
or \U$3963 ( \4679 , \4677 , \4678 );
and \U$3964 ( \4680 , \4417 , \4679 );
and \U$3965 ( \4681 , \882 , \4416_nRf40 );
or \U$3966 ( \4682 , \4680 , \4681 );
and \U$3967 ( \4683 , \4387 , \4682 );
and \U$3968 ( \4684 , \846 , \4386_nRf42 );
or \U$3969 ( \4685 , \4683 , \4684 );
and \U$3970 ( \4686 , \4357 , \4685 );
and \U$3971 ( \4687 , \810 , \4356_nR10fb );
or \U$3972 ( \4688 , \4686 , \4687 );
and \U$3973 ( \4689 , \4327 , \4688 );
and \U$3974 ( \4690 , \774 , \4326_nR10fd );
or \U$3975 ( \4691 , \4689 , \4690 );
and \U$3976 ( \4692 , \4297 , \4691 );
and \U$3977 ( \4693 , \694 , \4296_nR12e0 );
or \U$3978 ( \4694 , \4692 , \4693 );
nor \U$3979 ( \4695 , \4694 , \1231 );
not \U$3980 ( \4696 , \4695 );
and \U$3981 ( \4697 , \4259 , \1240 );
and \U$3982 ( \4698 , \4263 , \4697 );
xnor \U$3983 ( \4699 , \4265 , \4698 );
not \U$3984 ( \4700 , \4699 );
xor \U$3985 ( \4701 , \4263 , \4697 );
not \U$3986 ( \4702 , \4701 );
and \U$3987 ( \4703 , \4698 , \4265 );
nor \U$3988 ( \4704 , \4703 , RIb54abd0_17);
nand \U$3989 ( \4705 , \4702 , \4704 );
nor \U$3990 ( \4706 , \4700 , \4705 );
not \U$3991 ( \4707 , \4258 );
and \U$3992 ( \4708 , \4255 , \1240 , \4707 );
nor \U$3993 ( \4709 , \4708 , \1257 );
and \U$3994 ( \4710 , \4258 , \1240 );
and \U$3995 ( \4711 , RIb54a9f0_13, \1237 );
nor \U$3996 ( \4712 , \4710 , \4711 );
nor \U$3997 ( \4713 , \4709 , \4712 );
and \U$3998 ( \4714 , \4706 , \4713 );
and \U$3999 ( \4715 , RIb5515c0_243, \4714 );
nand \U$4000 ( \4716 , \4712 , \4709 );
nor \U$4001 ( \4717 , \4704 , \4716 , \4701 );
and \U$4002 ( \4718 , \4717 , \4699 );
and \U$4003 ( \4719 , RIb550be8_222, \4718 );
not \U$4004 ( \4720 , \4709 );
nor \U$4005 ( \4721 , \4720 , \4712 );
and \U$4006 ( \4722 , \4706 , \4721 );
and \U$4007 ( \4723 , \4722 , RIb5516b0_245);
not \U$4008 ( \4724 , \4712 );
nor \U$4009 ( \4725 , \4724 , \4709 );
and \U$4010 ( \4726 , \4706 , \4725 );
and \U$4011 ( \4727 , RIb551638_244, \4726 );
nor \U$4012 ( \4728 , \4723 , \4727 );
nor \U$4013 ( \4729 , \4705 , \4699 );
and \U$4014 ( \4730 , \4729 , \4725 );
and \U$4015 ( \4731 , \4730 , RIb551278_236);
and \U$4016 ( \4732 , \4729 , \4713 );
and \U$4017 ( \4733 , RIb551200_235, \4732 );
nor \U$4018 ( \4734 , \4731 , \4733 );
nand \U$4019 ( \4735 , \4701 , \4704 );
nor \U$4020 ( \4736 , \4735 , \4699 );
not \U$4021 ( \4737 , \4736 );
nor \U$4022 ( \4738 , \4737 , \4716 );
and \U$4023 ( \4739 , \4738 , RIb551188_234);
and \U$4024 ( \4740 , \4736 , \4721 );
and \U$4025 ( \4741 , RIb551110_233, \4740 );
nor \U$4026 ( \4742 , \4739 , \4741 );
not \U$4027 ( \4743 , \4729 );
nor \U$4028 ( \4744 , \4743 , \4716 );
and \U$4029 ( \4745 , \4744 , RIb551368_238);
and \U$4030 ( \4746 , \4729 , \4721 );
and \U$4031 ( \4747 , RIb5512f0_237, \4746 );
nor \U$4032 ( \4748 , \4745 , \4747 );
nand \U$4033 ( \4749 , \4728 , \4734 , \4742 , \4748 );
nor \U$4034 ( \4750 , \4715 , \4719 , \4749 );
not \U$4035 ( \4751 , \4699 );
nor \U$4036 ( \4752 , \4751 , \4735 );
not \U$4037 ( \4753 , \4752 );
nor \U$4038 ( \4754 , \4753 , \4716 );
and \U$4039 ( \4755 , \4754 , RIb551548_242);
and \U$4040 ( \4756 , \4752 , \4721 );
and \U$4041 ( \4757 , RIb5514d0_241, \4756 );
nor \U$4042 ( \4758 , \4755 , \4757 );
and \U$4043 ( \4759 , \4736 , \4725 );
and \U$4044 ( \4760 , RIb551098_232, \4759 );
and \U$4045 ( \4761 , \4736 , \4713 );
and \U$4046 ( \4762 , RIb551020_231, \4761 );
and \U$4047 ( \4763 , \4752 , \4725 );
and \U$4048 ( \4764 , \4763 , RIb551458_240);
and \U$4049 ( \4765 , \4752 , \4713 );
and \U$4050 ( \4766 , RIb5513e0_239, \4765 );
nor \U$4051 ( \4767 , \4764 , \4766 );
not \U$4052 ( \4768 , \4767 );
nor \U$4053 ( \4769 , \4760 , \4762 , \4768 );
nand \U$4054 ( \4770 , \4750 , \4758 , \1270 , \4769 );
buf \U$4055 ( \4771 , \766 );
_DC r194f ( \4772_nR194f , \4770 , \4771 );
not \U$4056 ( \4773 , \4772_nR194f );
nor \U$4057 ( \4774 , \4696 , \4773 );
xor \U$4058 ( \4775 , \694 , \4296_nR12e0 );
xor \U$4059 ( \4776 , \4775 , \4691 );
not \U$4060 ( \4777 , \4776 );
xor \U$4061 ( \4778 , \774 , \4326_nR10fd );
xor \U$4062 ( \4779 , \4778 , \4688 );
not \U$4063 ( \4780 , \4779 );
and \U$4064 ( \4781 , \4777 , \4780 );
and \U$4065 ( \4782 , \4694 , \1231 );
nor \U$4066 ( \4783 , \4782 , \4695 );
nor \U$4067 ( \4784 , \4781 , \4783 );
not \U$4068 ( \4785 , \4784 );
and \U$4069 ( \4786 , RIb552178_268, \4740 );
and \U$4070 ( \4787 , RIb552718_280, \4722 );
and \U$4071 ( \4788 , \4714 , RIb552628_278);
and \U$4072 ( \4789 , RIb5524c0_275, \4763 );
nor \U$4073 ( \4790 , \4788 , \4789 );
and \U$4074 ( \4791 , \4759 , RIb552100_267);
and \U$4075 ( \4792 , RIb552088_266, \4761 );
nor \U$4076 ( \4793 , \4791 , \4792 );
and \U$4077 ( \4794 , \4718 , RIb552010_265);
and \U$4078 ( \4795 , RIb552448_274, \4765 );
nor \U$4079 ( \4796 , \4794 , \4795 );
and \U$4080 ( \4797 , \4754 , RIb5525b0_277);
and \U$4081 ( \4798 , RIb552538_276, \4756 );
nor \U$4082 ( \4799 , \4797 , \4798 );
nand \U$4083 ( \4800 , \4790 , \4793 , \4796 , \4799 );
nor \U$4084 ( \4801 , \4786 , \4787 , \4800 );
and \U$4085 ( \4802 , \4726 , RIb5526a0_279);
and \U$4086 ( \4803 , RIb5523d0_273, \4744 );
nor \U$4087 ( \4804 , \4802 , \4803 );
nand \U$4088 ( \4805 , RIb552790_281, \1269 );
and \U$4089 ( \4806 , RIb552358_272, \4746 );
and \U$4090 ( \4807 , RIb5522e0_271, \4730 );
and \U$4091 ( \4808 , \4738 , RIb5521f0_269);
and \U$4092 ( \4809 , RIb552268_270, \4732 );
nor \U$4093 ( \4810 , \4808 , \4809 );
not \U$4094 ( \4811 , \4810 );
nor \U$4095 ( \4812 , \4806 , \4807 , \4811 );
nand \U$4096 ( \4813 , \4801 , \4804 , \4805 , \4812 );
_DC r1a6c ( \4814_nR1a6c , \4813 , \4771 );
or \U$4097 ( \4815 , \4785 , \4814_nR1a6c );
not \U$4098 ( \4816 , \4814_nR1a6c );
and \U$4099 ( \4817 , \4783 , \4776 );
nor \U$4100 ( \4818 , \4783 , \4776 );
xnor \U$4101 ( \4819 , \4779 , \4776 );
not \U$4102 ( \4820 , \4819 );
nor \U$4103 ( \4821 , \4817 , \4818 , \4820 );
nand \U$4104 ( \4822 , \4821 , \4785 );
or \U$4105 ( \4823 , \4816 , \4822 );
or \U$4106 ( \4824 , \4821 , \4785 );
nand \U$4107 ( \4825 , \4815 , \4823 , \4824 );
xnor \U$4108 ( \4826 , \4774 , \4825 );
nand \U$4109 ( \4827 , \4820 , \4785 );
or \U$4110 ( \4828 , \4827 , \4816 );
or \U$4111 ( \4829 , \4773 , \4822 );
or \U$4112 ( \4830 , \4819 , \4816 );
or \U$4113 ( \4831 , \4785 , \4772_nR194f );
nand \U$4114 ( \4832 , \4831 , \4824 );
nand \U$4115 ( \4833 , \4830 , \4832 );
nand \U$4116 ( \4834 , \4828 , \4829 , \4833 );
xor \U$4117 ( \4835 , \810 , \4356_nR10fb );
xor \U$4118 ( \4836 , \4835 , \4685 );
xor \U$4119 ( \4837 , \846 , \4386_nRf42 );
xor \U$4120 ( \4838 , \4837 , \4682 );
nor \U$4121 ( \4839 , \4836 , \4838 );
or \U$4122 ( \4840 , \4779 , \4839 );
and \U$4123 ( \4841 , \4834 , \4840 );
and \U$4124 ( \4842 , RIb552970_285, \4740 );
and \U$4125 ( \4843 , RIb552e20_295, \4714 );
and \U$4126 ( \4844 , \4763 , RIb552cb8_292);
and \U$4127 ( \4845 , RIb552c40_291, \4765 );
nor \U$4128 ( \4846 , \4844 , \4845 );
and \U$4129 ( \4847 , \4722 , RIb552f10_297);
and \U$4130 ( \4848 , RIb5528f8_284, \4759 );
nor \U$4131 ( \4849 , \4847 , \4848 );
and \U$4132 ( \4850 , \4718 , RIb552808_282);
and \U$4133 ( \4851 , RIb552880_283, \4761 );
nor \U$4134 ( \4852 , \4850 , \4851 );
and \U$4135 ( \4853 , \4726 , RIb552e98_296);
and \U$4136 ( \4854 , RIb552d30_293, \4756 );
nor \U$4137 ( \4855 , \4853 , \4854 );
nand \U$4138 ( \4856 , \4846 , \4849 , \4852 , \4855 );
nor \U$4139 ( \4857 , \4842 , \4843 , \4856 );
and \U$4140 ( \4858 , \4744 , RIb552bc8_290);
and \U$4141 ( \4859 , RIb552da8_294, \4754 );
nor \U$4142 ( \4860 , \4858 , \4859 );
nand \U$4143 ( \4861 , RIb552f88_298, \1269 );
and \U$4144 ( \4862 , RIb552b50_289, \4746 );
and \U$4145 ( \4863 , RIb552ad8_288, \4730 );
and \U$4146 ( \4864 , \4738 , RIb5529e8_286);
and \U$4147 ( \4865 , RIb552a60_287, \4732 );
nor \U$4148 ( \4866 , \4864 , \4865 );
not \U$4149 ( \4867 , \4866 );
nor \U$4150 ( \4868 , \4862 , \4863 , \4867 );
nand \U$4151 ( \4869 , \4857 , \4860 , \4861 , \4868 );
_DC r1859 ( \4870_nR1859 , \4869 , \4771 );
not \U$4152 ( \4871 , \4870_nR1859 );
nor \U$4153 ( \4872 , \4696 , \4871 );
nor \U$4154 ( \4873 , \4841 , \4872 );
xor \U$4155 ( \4874 , \4826 , \4873 );
not \U$4156 ( \4875 , \4874 );
not \U$4157 ( \4876 , \4836 );
not \U$4158 ( \4877 , \4779 );
or \U$4159 ( \4878 , \4876 , \4877 );
or \U$4160 ( \4879 , \4779 , \4836 );
nand \U$4161 ( \4880 , \4878 , \4879 );
xor \U$4162 ( \4881 , \4838 , \4836 );
nor \U$4163 ( \4882 , \4880 , \4881 );
not \U$4164 ( \4883 , \4882 );
not \U$4165 ( \4884 , \4840 );
nor \U$4166 ( \4885 , \4883 , \4884 );
not \U$4167 ( \4886 , \4885 );
or \U$4168 ( \4887 , \4886 , \4816 );
or \U$4169 ( \4888 , \4883 , \4816 );
nand \U$4170 ( \4889 , \4888 , \4884 );
nand \U$4171 ( \4890 , \4887 , \4889 );
or \U$4172 ( \4891 , \4827 , \4773 );
or \U$4173 ( \4892 , \4871 , \4822 );
or \U$4174 ( \4893 , \4819 , \4773 );
or \U$4175 ( \4894 , \4785 , \4870_nR1859 );
nand \U$4176 ( \4895 , \4894 , \4824 );
nand \U$4177 ( \4896 , \4893 , \4895 );
nand \U$4178 ( \4897 , \4891 , \4892 , \4896 );
and \U$4179 ( \4898 , \4890 , \4897 );
and \U$4180 ( \4899 , \4834 , \4840 );
not \U$4181 ( \4900 , \4834 );
and \U$4182 ( \4901 , \4900 , \4884 );
nor \U$4183 ( \4902 , \4899 , \4901 );
xor \U$4184 ( \4903 , \4872 , \4902 );
and \U$4185 ( \4904 , \4898 , \4903 );
and \U$4186 ( \4905 , \4875 , \4904 );
or \U$4187 ( \4906 , \4905 , \4784 );
and \U$4188 ( \4907 , \4905 , \4784 );
and \U$4189 ( \4908 , \4774 , \4825 );
nor \U$4190 ( \4909 , \4907 , \4908 );
nand \U$4191 ( \4910 , \4906 , \4909 );
not \U$4192 ( \4911 , \4910 );
and \U$4193 ( \4912 , \4695 , \4814_nR1a6c );
and \U$4194 ( \4913 , \4826 , \4873 );
nor \U$4195 ( \4914 , \4912 , \4913 );
not \U$4196 ( \4915 , \4914 );
and \U$4197 ( \4916 , \4911 , \4915 );
and \U$4198 ( \4917 , \4910 , \4914 );
nor \U$4199 ( \4918 , \4916 , \4917 );
not \U$4200 ( \4919 , \4918 );
and \U$4201 ( \4920 , \4772_nR194f , \4885 );
and \U$4202 ( \4921 , \4840 , \4881 );
and \U$4203 ( \4922 , \4921 , \4814_nR1a6c );
nand \U$4204 ( \4923 , \4772_nR194f , \4882 );
or \U$4205 ( \4924 , \4840 , \4814_nR1a6c );
or \U$4206 ( \4925 , \4840 , \4881 );
nand \U$4207 ( \4926 , \4924 , \4925 );
and \U$4208 ( \4927 , \4923 , \4926 );
nor \U$4209 ( \4928 , \4920 , \4922 , \4927 );
xor \U$4210 ( \4929 , \882 , \4416_nRf40 );
xor \U$4211 ( \4930 , \4929 , \4679 );
xor \U$4212 ( \4931 , \918 , \4446_nRdc1 );
xor \U$4213 ( \4932 , \4931 , \4676 );
nor \U$4214 ( \4933 , \4930 , \4932 );
or \U$4215 ( \4934 , \4838 , \4933 );
not \U$4216 ( \4935 , \4934 );
xor \U$4217 ( \4936 , \4928 , \4935 );
not \U$4218 ( \4937 , \4827 );
and \U$4219 ( \4938 , \4870_nR1859 , \4937 );
not \U$4220 ( \4939 , \4822 );
and \U$4221 ( \4940 , RIb553960_319, \4740 );
and \U$4222 ( \4941 , RIb553e10_329, \4714 );
and \U$4223 ( \4942 , \4756 , RIb553d20_327);
and \U$4224 ( \4943 , RIb553ca8_326, \4763 );
nor \U$4225 ( \4944 , \4942 , \4943 );
and \U$4226 ( \4945 , \4722 , RIb553f00_331);
and \U$4227 ( \4946 , RIb5538e8_318, \4759 );
nor \U$4228 ( \4947 , \4945 , \4946 );
and \U$4229 ( \4948 , \4718 , RIb5537f8_316);
and \U$4230 ( \4949 , RIb553870_317, \4761 );
nor \U$4231 ( \4950 , \4948 , \4949 );
and \U$4232 ( \4951 , \4726 , RIb553e88_330);
and \U$4233 ( \4952 , RIb553d98_328, \4754 );
nor \U$4234 ( \4953 , \4951 , \4952 );
nand \U$4235 ( \4954 , \4944 , \4947 , \4950 , \4953 );
nor \U$4236 ( \4955 , \4940 , \4941 , \4954 );
and \U$4237 ( \4956 , \4744 , RIb553bb8_324);
and \U$4238 ( \4957 , RIb553c30_325, \4765 );
nor \U$4239 ( \4958 , \4956 , \4957 );
nand \U$4240 ( \4959 , RIb553f78_332, \1269 );
and \U$4241 ( \4960 , RIb553b40_323, \4746 );
and \U$4242 ( \4961 , RIb553ac8_322, \4730 );
and \U$4243 ( \4962 , \4738 , RIb5539d8_320);
and \U$4244 ( \4963 , RIb553a50_321, \4732 );
nor \U$4245 ( \4964 , \4962 , \4963 );
not \U$4246 ( \4965 , \4964 );
nor \U$4247 ( \4966 , \4960 , \4961 , \4965 );
nand \U$4248 ( \4967 , \4955 , \4958 , \4959 , \4966 );
_DC r171b ( \4968_nR171b , \4967 , \4771 );
and \U$4249 ( \4969 , \4939 , \4968_nR171b );
nand \U$4250 ( \4970 , \4870_nR1859 , \4820 );
or \U$4251 ( \4971 , \4785 , \4968_nR171b );
nand \U$4252 ( \4972 , \4971 , \4824 );
and \U$4253 ( \4973 , \4970 , \4972 );
nor \U$4254 ( \4974 , \4938 , \4969 , \4973 );
and \U$4255 ( \4975 , \4936 , \4974 );
and \U$4256 ( \4976 , \4928 , \4935 );
or \U$4257 ( \4977 , \4975 , \4976 );
xor \U$4258 ( \4978 , \4890 , \4897 );
not \U$4259 ( \4979 , \4978 );
nand \U$4260 ( \4980 , \4968_nR171b , \4695 );
not \U$4261 ( \4981 , \4980 );
and \U$4262 ( \4982 , \4979 , \4981 );
and \U$4263 ( \4983 , \4978 , \4980 );
nor \U$4264 ( \4984 , \4982 , \4983 );
nand \U$4265 ( \4985 , \4977 , \4984 );
xor \U$4266 ( \4986 , \4898 , \4903 );
and \U$4267 ( \4987 , \4985 , \4986 );
xor \U$4268 ( \4988 , \4875 , \4904 );
and \U$4269 ( \4989 , \4987 , \4988 );
not \U$4270 ( \4990 , \4989 );
and \U$4271 ( \4991 , \4919 , \4990 );
and \U$4272 ( \4992 , \4918 , \4989 );
nor \U$4273 ( \4993 , \4991 , \4992 );
not \U$4274 ( \4994 , \4993 );
not \U$4275 ( \4995 , \4978 );
nor \U$4276 ( \4996 , \4995 , \4980 );
not \U$4277 ( \4997 , \4996 );
or \U$4278 ( \4998 , \4984 , \4977 );
nand \U$4279 ( \4999 , \4998 , \4985 );
and \U$4280 ( \5000 , \4968_nR171b , \4937 );
and \U$4281 ( \5001 , RIb553708_314, \4722 );
and \U$4282 ( \5002 , RIb553000_299, \4718 );
and \U$4283 ( \5003 , \4730 , RIb5532d0_305);
and \U$4284 ( \5004 , RIb553258_304, \4732 );
nor \U$4285 ( \5005 , \5003 , \5004 );
and \U$4286 ( \5006 , \4744 , RIb5533c0_307);
and \U$4287 ( \5007 , RIb553348_306, \4746 );
nor \U$4288 ( \5008 , \5006 , \5007 );
and \U$4289 ( \5009 , \4738 , RIb5531e0_303);
and \U$4290 ( \5010 , RIb553168_302, \4740 );
nor \U$4291 ( \5011 , \5009 , \5010 );
and \U$4292 ( \5012 , \4763 , RIb5534b0_309);
and \U$4293 ( \5013 , RIb553438_308, \4765 );
nor \U$4294 ( \5014 , \5012 , \5013 );
nand \U$4295 ( \5015 , \5005 , \5008 , \5011 , \5014 );
nor \U$4296 ( \5016 , \5001 , \5002 , \5015 );
and \U$4297 ( \5017 , \4726 , RIb553690_313);
and \U$4298 ( \5018 , RIb553618_312, \4714 );
nor \U$4299 ( \5019 , \5017 , \5018 );
and \U$4300 ( \5020 , RIb5530f0_301, \4759 );
and \U$4301 ( \5021 , RIb553078_300, \4761 );
and \U$4302 ( \5022 , \4754 , RIb5535a0_311);
and \U$4303 ( \5023 , RIb553528_310, \4756 );
nor \U$4304 ( \5024 , \5022 , \5023 );
not \U$4305 ( \5025 , \5024 );
nor \U$4306 ( \5026 , \5020 , \5021 , \5025 );
nand \U$4307 ( \5027 , \5016 , \5019 , \1550 , \5026 );
_DC r162d ( \5028_nR162d , \5027 , \4771 );
and \U$4308 ( \5029 , \4939 , \5028_nR162d );
nand \U$4309 ( \5030 , \4968_nR171b , \4820 );
or \U$4310 ( \5031 , \4785 , \5028_nR162d );
nand \U$4311 ( \5032 , \5031 , \4824 );
and \U$4312 ( \5033 , \5030 , \5032 );
nor \U$4313 ( \5034 , \5000 , \5029 , \5033 );
and \U$4314 ( \5035 , RIb5546f8_348, \4722 );
and \U$4315 ( \5036 , RIb553ff0_333, \4718 );
and \U$4316 ( \5037 , \4754 , RIb554590_345);
and \U$4317 ( \5038 , RIb554518_344, \4756 );
nor \U$4318 ( \5039 , \5037 , \5038 );
and \U$4319 ( \5040 , \4730 , RIb5542c0_339);
and \U$4320 ( \5041 , RIb554248_338, \4732 );
nor \U$4321 ( \5042 , \5040 , \5041 );
and \U$4322 ( \5043 , \4738 , RIb5541d0_337);
and \U$4323 ( \5044 , RIb554158_336, \4740 );
nor \U$4324 ( \5045 , \5043 , \5044 );
and \U$4325 ( \5046 , \4744 , RIb5543b0_341);
and \U$4326 ( \5047 , RIb554338_340, \4746 );
nor \U$4327 ( \5048 , \5046 , \5047 );
nand \U$4328 ( \5049 , \5039 , \5042 , \5045 , \5048 );
nor \U$4329 ( \5050 , \5035 , \5036 , \5049 );
and \U$4330 ( \5051 , \4726 , RIb554680_347);
and \U$4331 ( \5052 , RIb554608_346, \4714 );
nor \U$4332 ( \5053 , \5051 , \5052 );
nand \U$4333 ( \5054 , RIb554770_349, \1269 );
and \U$4334 ( \5055 , RIb5540e0_335, \4759 );
and \U$4335 ( \5056 , RIb554068_334, \4761 );
and \U$4336 ( \5057 , \4763 , RIb5544a0_343);
and \U$4337 ( \5058 , RIb554428_342, \4765 );
nor \U$4338 ( \5059 , \5057 , \5058 );
not \U$4339 ( \5060 , \5059 );
nor \U$4340 ( \5061 , \5055 , \5056 , \5060 );
nand \U$4341 ( \5062 , \5050 , \5053 , \5054 , \5061 );
_DC r150e ( \5063_nR150e , \5062 , \4771 );
nand \U$4342 ( \5064 , \5063_nR150e , \4695 );
or \U$4343 ( \5065 , \5034 , \5064 );
and \U$4344 ( \5066 , \4838 , \4930 );
nor \U$4345 ( \5067 , \4838 , \4930 );
xor \U$4346 ( \5068 , \4930 , \4932 );
nor \U$4347 ( \5069 , \5066 , \5067 , \5068 );
and \U$4348 ( \5070 , \5069 , \4934 );
and \U$4349 ( \5071 , \4814_nR1a6c , \5070 );
and \U$4350 ( \5072 , \4816 , \4935 );
or \U$4351 ( \5073 , \5069 , \4934 );
not \U$4352 ( \5074 , \5073 );
nor \U$4353 ( \5075 , \5071 , \5072 , \5074 );
and \U$4354 ( \5076 , \4870_nR1859 , \4885 );
and \U$4355 ( \5077 , \4921 , \4772_nR194f );
nand \U$4356 ( \5078 , \4870_nR1859 , \4882 );
or \U$4357 ( \5079 , \4840 , \4772_nR194f );
nand \U$4358 ( \5080 , \5079 , \4925 );
and \U$4359 ( \5081 , \5078 , \5080 );
nor \U$4360 ( \5082 , \5076 , \5077 , \5081 );
or \U$4361 ( \5083 , \5075 , \5082 );
nand \U$4362 ( \5084 , \5065 , \5083 );
not \U$4363 ( \5085 , \5084 );
nand \U$4364 ( \5086 , \5028_nR162d , \4695 );
xor \U$4365 ( \5087 , \4928 , \4935 );
xor \U$4366 ( \5088 , \5087 , \4974 );
xnor \U$4367 ( \5089 , \5086 , \5088 );
nor \U$4368 ( \5090 , \5085 , \5089 );
and \U$4369 ( \5091 , \4999 , \5090 );
xor \U$4370 ( \5092 , \4985 , \4986 );
or \U$4371 ( \5093 , \5091 , \5092 );
not \U$4372 ( \5094 , \5093 );
or \U$4373 ( \5095 , \4997 , \5094 );
nand \U$4374 ( \5096 , \5092 , \5091 );
nand \U$4375 ( \5097 , \5095 , \5096 );
xor \U$4376 ( \5098 , \4987 , \4988 );
and \U$4377 ( \5099 , \5097 , \5098 );
not \U$4378 ( \5100 , \5097 );
not \U$4379 ( \5101 , \5098 );
and \U$4380 ( \5102 , \5100 , \5101 );
not \U$4381 ( \5103 , \4996 );
and \U$4382 ( \5104 , \5096 , \5093 );
not \U$4383 ( \5105 , \5104 );
or \U$4384 ( \5106 , \5103 , \5105 );
or \U$4385 ( \5107 , \5104 , \4996 );
nand \U$4386 ( \5108 , \5106 , \5107 );
xor \U$4387 ( \5109 , \4999 , \5090 );
not \U$4388 ( \5110 , \5089 );
not \U$4389 ( \5111 , \5084 );
and \U$4390 ( \5112 , \5110 , \5111 );
and \U$4391 ( \5113 , \5089 , \5084 );
nor \U$4392 ( \5114 , \5112 , \5113 );
not \U$4393 ( \5115 , \5068 );
nor \U$4394 ( \5116 , \4935 , \5115 );
and \U$4395 ( \5117 , \4814_nR1a6c , \5116 );
or \U$4396 ( \5118 , \4934 , \4772_nR194f );
nand \U$4397 ( \5119 , \5118 , \5073 );
nand \U$4398 ( \5120 , \4814_nR1a6c , \5068 );
and \U$4399 ( \5121 , \5119 , \5120 );
and \U$4400 ( \5122 , \4772_nR194f , \5070 );
nor \U$4401 ( \5123 , \5117 , \5121 , \5122 );
and \U$4402 ( \5124 , \4968_nR171b , \4885 );
and \U$4403 ( \5125 , \4921 , \4870_nR1859 );
nand \U$4404 ( \5126 , \4968_nR171b , \4882 );
or \U$4405 ( \5127 , \4840 , \4870_nR1859 );
nand \U$4406 ( \5128 , \5127 , \4925 );
and \U$4407 ( \5129 , \5126 , \5128 );
nor \U$4408 ( \5130 , \5124 , \5125 , \5129 );
nand \U$4409 ( \5131 , \5123 , \5130 );
xor \U$4410 ( \5132 , \954 , \4476_nRdbf );
xor \U$4411 ( \5133 , \5132 , \4673 );
xor \U$4412 ( \5134 , \990 , \4506_nRc88 );
xor \U$4413 ( \5135 , \5134 , \4670 );
nor \U$4414 ( \5136 , \5133 , \5135 );
or \U$4415 ( \5137 , \4932 , \5136 );
and \U$4416 ( \5138 , \5131 , \5137 );
and \U$4417 ( \5139 , RIb5556e8_382, \4722 );
and \U$4418 ( \5140 , RIb554fe0_367, \4718 );
and \U$4419 ( \5141 , \4726 , RIb555670_381);
and \U$4420 ( \5142 , RIb555580_379, \4754 );
nor \U$4421 ( \5143 , \5141 , \5142 );
and \U$4422 ( \5144 , \4744 , RIb5553a0_375);
and \U$4423 ( \5145 , RIb555328_374, \4746 );
nor \U$4424 ( \5146 , \5144 , \5145 );
and \U$4425 ( \5147 , \4738 , RIb5551c0_371);
and \U$4426 ( \5148 , RIb555148_370, \4740 );
nor \U$4427 ( \5149 , \5147 , \5148 );
and \U$4428 ( \5150 , \4730 , RIb5552b0_373);
and \U$4429 ( \5151 , RIb555238_372, \4732 );
nor \U$4430 ( \5152 , \5150 , \5151 );
nand \U$4431 ( \5153 , \5143 , \5146 , \5149 , \5152 );
nor \U$4432 ( \5154 , \5139 , \5140 , \5153 );
and \U$4433 ( \5155 , \4714 , RIb5555f8_380);
and \U$4434 ( \5156 , RIb555508_378, \4756 );
nor \U$4435 ( \5157 , \5155 , \5156 );
nand \U$4436 ( \5158 , RIb555760_383, \1269 );
and \U$4437 ( \5159 , RIb5550d0_369, \4759 );
and \U$4438 ( \5160 , RIb555058_368, \4761 );
and \U$4439 ( \5161 , \4763 , RIb555490_377);
and \U$4440 ( \5162 , RIb555418_376, \4765 );
nor \U$4441 ( \5163 , \5161 , \5162 );
not \U$4442 ( \5164 , \5163 );
nor \U$4443 ( \5165 , \5159 , \5160 , \5164 );
nand \U$4444 ( \5166 , \5154 , \5157 , \5158 , \5165 );
_DC r140b ( \5167_nR140b , \5166 , \4771 );
not \U$4445 ( \5168 , \5167_nR140b );
nor \U$4446 ( \5169 , \4696 , \5168 );
not \U$4447 ( \5170 , \5028_nR162d );
or \U$4448 ( \5171 , \4827 , \5170 );
not \U$4449 ( \5172 , \5063_nR150e );
or \U$4450 ( \5173 , \5172 , \4822 );
or \U$4451 ( \5174 , \4819 , \5170 );
or \U$4452 ( \5175 , \4785 , \5063_nR150e );
nand \U$4453 ( \5176 , \5175 , \4824 );
nand \U$4454 ( \5177 , \5174 , \5176 );
nand \U$4455 ( \5178 , \5171 , \5173 , \5177 );
and \U$4456 ( \5179 , \5169 , \5178 );
nor \U$4457 ( \5180 , \5130 , \5123 );
nor \U$4458 ( \5181 , \5138 , \5179 , \5180 );
xnor \U$4459 ( \5182 , \5064 , \5034 );
not \U$4460 ( \5183 , \5182 );
xor \U$4461 ( \5184 , \5075 , \5082 );
not \U$4462 ( \5185 , \5184 );
and \U$4463 ( \5186 , \5183 , \5185 );
and \U$4464 ( \5187 , \5182 , \5184 );
nor \U$4465 ( \5188 , \5186 , \5187 );
nand \U$4466 ( \5189 , \5181 , \5188 );
xor \U$4467 ( \5190 , \5169 , \5178 );
not \U$4468 ( \5191 , \5190 );
not \U$4469 ( \5192 , \5180 );
nand \U$4470 ( \5193 , \5192 , \5131 );
not \U$4471 ( \5194 , \5193 );
not \U$4472 ( \5195 , \5137 );
and \U$4473 ( \5196 , \5194 , \5195 );
and \U$4474 ( \5197 , \5193 , \5137 );
nor \U$4475 ( \5198 , \5196 , \5197 );
nor \U$4476 ( \5199 , \5191 , \5198 );
not \U$4477 ( \5200 , \5199 );
not \U$4478 ( \5201 , \5133 );
not \U$4479 ( \5202 , \4932 );
or \U$4480 ( \5203 , \5201 , \5202 );
or \U$4481 ( \5204 , \4932 , \5133 );
nand \U$4482 ( \5205 , \5203 , \5204 );
xor \U$4483 ( \5206 , \5135 , \5133 );
nor \U$4484 ( \5207 , \5205 , \5206 );
not \U$4485 ( \5208 , \5207 );
not \U$4486 ( \5209 , \5137 );
nor \U$4487 ( \5210 , \5208 , \5209 );
not \U$4488 ( \5211 , \5210 );
or \U$4489 ( \5212 , \5211 , \4816 );
or \U$4490 ( \5213 , \5208 , \4816 );
nand \U$4491 ( \5214 , \5213 , \5209 );
nand \U$4492 ( \5215 , \5212 , \5214 );
not \U$4493 ( \5216 , \5116 );
or \U$4494 ( \5217 , \5216 , \4773 );
not \U$4495 ( \5218 , \5070 );
or \U$4496 ( \5219 , \4871 , \5218 );
or \U$4497 ( \5220 , \5115 , \4773 );
or \U$4498 ( \5221 , \4934 , \4870_nR1859 );
nand \U$4499 ( \5222 , \5221 , \5073 );
nand \U$4500 ( \5223 , \5220 , \5222 );
nand \U$4501 ( \5224 , \5217 , \5219 , \5223 );
and \U$4502 ( \5225 , \5215 , \5224 );
and \U$4503 ( \5226 , \5028_nR162d , \4885 );
and \U$4504 ( \5227 , \4921 , \4968_nR171b );
nand \U$4505 ( \5228 , \5028_nR162d , \4882 );
or \U$4506 ( \5229 , \4840 , \4968_nR171b );
nand \U$4507 ( \5230 , \5229 , \4925 );
and \U$4508 ( \5231 , \5228 , \5230 );
nor \U$4509 ( \5232 , \5226 , \5227 , \5231 );
and \U$4510 ( \5233 , RIb554950_353, \4740 );
and \U$4511 ( \5234 , RIb554ef0_365, \4722 );
and \U$4512 ( \5235 , \4754 , RIb554d88_362);
and \U$4513 ( \5236 , RIb554e00_363, \4714 );
nor \U$4514 ( \5237 , \5235 , \5236 );
and \U$4515 ( \5238 , \4759 , RIb5548d8_352);
and \U$4516 ( \5239 , RIb554860_351, \4761 );
nor \U$4517 ( \5240 , \5238 , \5239 );
and \U$4518 ( \5241 , \4726 , RIb554e78_364);
and \U$4519 ( \5242 , RIb5547e8_350, \4718 );
nor \U$4520 ( \5243 , \5241 , \5242 );
and \U$4521 ( \5244 , \4756 , RIb554d10_361);
and \U$4522 ( \5245 , RIb554c98_360, \4763 );
nor \U$4523 ( \5246 , \5244 , \5245 );
nand \U$4524 ( \5247 , \5237 , \5240 , \5243 , \5246 );
nor \U$4525 ( \5248 , \5233 , \5234 , \5247 );
and \U$4526 ( \5249 , \4744 , RIb554ba8_358);
and \U$4527 ( \5250 , RIb554c20_359, \4765 );
nor \U$4528 ( \5251 , \5249 , \5250 );
nand \U$4529 ( \5252 , RIb554f68_366, \1269 );
and \U$4530 ( \5253 , RIb554b30_357, \4746 );
and \U$4531 ( \5254 , RIb554ab8_356, \4730 );
and \U$4532 ( \5255 , \4738 , RIb5549c8_354);
and \U$4533 ( \5256 , RIb554a40_355, \4732 );
nor \U$4534 ( \5257 , \5255 , \5256 );
not \U$4535 ( \5258 , \5257 );
nor \U$4536 ( \5259 , \5253 , \5254 , \5258 );
nand \U$4537 ( \5260 , \5248 , \5251 , \5252 , \5259 );
_DC r12fd ( \5261_nR12fd , \5260 , \4771 );
nand \U$4538 ( \5262 , \5261_nR12fd , \4695 );
and \U$4539 ( \5263 , \5232 , \5262 );
and \U$4540 ( \5264 , \5063_nR150e , \4937 );
and \U$4541 ( \5265 , \4939 , \5167_nR140b );
nand \U$4542 ( \5266 , \5063_nR150e , \4820 );
or \U$4543 ( \5267 , \4785 , \5167_nR140b );
nand \U$4544 ( \5268 , \5267 , \4824 );
and \U$4545 ( \5269 , \5266 , \5268 );
nor \U$4546 ( \5270 , \5264 , \5265 , \5269 );
nor \U$4547 ( \5271 , \5263 , \5270 );
nand \U$4548 ( \5272 , \5225 , \5271 );
nor \U$4549 ( \5273 , \5200 , \5272 );
nor \U$4550 ( \5274 , \5189 , \5273 );
or \U$4551 ( \5275 , \5114 , \5274 );
or \U$4552 ( \5276 , \5086 , \5088 );
nand \U$4553 ( \5277 , \5273 , \5189 );
nand \U$4554 ( \5278 , \5275 , \5276 , \5277 );
nand \U$4555 ( \5279 , \5109 , \5278 );
xor \U$4556 ( \5280 , \5108 , \5279 );
or \U$4557 ( \5281 , \5278 , \5109 );
nand \U$4558 ( \5282 , \5281 , \5279 );
not \U$4559 ( \5283 , \5190 );
not \U$4560 ( \5284 , \5198 );
and \U$4561 ( \5285 , \5283 , \5284 );
and \U$4562 ( \5286 , \5190 , \5198 );
nor \U$4563 ( \5287 , \5285 , \5286 );
not \U$4564 ( \5288 , \5287 );
xor \U$4565 ( \5289 , \5225 , \5271 );
nand \U$4566 ( \5290 , \5288 , \5289 );
not \U$4567 ( \5291 , \5290 );
nand \U$4568 ( \5292 , \4772_nR194f , \5207 );
or \U$4569 ( \5293 , \5137 , \4814_nR1a6c );
or \U$4570 ( \5294 , \5137 , \5206 );
nand \U$4571 ( \5295 , \5293 , \5294 );
and \U$4572 ( \5296 , \5292 , \5295 );
and \U$4573 ( \5297 , \5137 , \5206 );
and \U$4574 ( \5298 , \5297 , \4814_nR1a6c );
and \U$4575 ( \5299 , \4772_nR194f , \5210 );
nor \U$4576 ( \5300 , \5296 , \5298 , \5299 );
not \U$4577 ( \5301 , \5300 );
xor \U$4578 ( \5302 , \1026 , \4536_nRc86 );
xor \U$4579 ( \5303 , \5302 , \4667 );
xor \U$4580 ( \5304 , \1062 , \4566_nRb9a );
xor \U$4581 ( \5305 , \5304 , \4664 );
nor \U$4582 ( \5306 , \5303 , \5305 );
or \U$4583 ( \5307 , \5135 , \5306 );
not \U$4584 ( \5308 , \5307 );
not \U$4585 ( \5309 , \5308 );
and \U$4586 ( \5310 , \5301 , \5309 );
and \U$4587 ( \5311 , \5300 , \5308 );
and \U$4588 ( \5312 , \4870_nR1859 , \5116 );
or \U$4589 ( \5313 , \4934 , \4968_nR171b );
nand \U$4590 ( \5314 , \5313 , \5073 );
nand \U$4591 ( \5315 , \4870_nR1859 , \5068 );
and \U$4592 ( \5316 , \5314 , \5315 );
and \U$4593 ( \5317 , \4968_nR171b , \5070 );
nor \U$4594 ( \5318 , \5312 , \5316 , \5317 );
nor \U$4595 ( \5319 , \5311 , \5318 );
nor \U$4596 ( \5320 , \5310 , \5319 );
not \U$4597 ( \5321 , \5320 );
and \U$4598 ( \5322 , \5063_nR150e , \4885 );
and \U$4599 ( \5323 , \4921 , \5028_nR162d );
nand \U$4600 ( \5324 , \5063_nR150e , \4882 );
or \U$4601 ( \5325 , \4840 , \5028_nR162d );
nand \U$4602 ( \5326 , \5325 , \4925 );
and \U$4603 ( \5327 , \5324 , \5326 );
nor \U$4604 ( \5328 , \5322 , \5323 , \5327 );
and \U$4605 ( \5329 , RIb556138_404, \4740 );
and \U$4606 ( \5330 , RIb5564f8_412, \4756 );
and \U$4607 ( \5331 , \4722 , RIb5566d8_416);
and \U$4608 ( \5332 , RIb556660_415, \4726 );
nor \U$4609 ( \5333 , \5331 , \5332 );
and \U$4610 ( \5334 , \4759 , RIb5560c0_403);
and \U$4611 ( \5335 , RIb556048_402, \4761 );
nor \U$4612 ( \5336 , \5334 , \5335 );
and \U$4613 ( \5337 , \4718 , RIb555fd0_401);
and \U$4614 ( \5338 , RIb5565e8_414, \4714 );
nor \U$4615 ( \5339 , \5337 , \5338 );
and \U$4616 ( \5340 , \4754 , RIb556570_413);
and \U$4617 ( \5341 , RIb556408_410, \4765 );
nor \U$4618 ( \5342 , \5340 , \5341 );
nand \U$4619 ( \5343 , \5333 , \5336 , \5339 , \5342 );
nor \U$4620 ( \5344 , \5329 , \5330 , \5343 );
and \U$4621 ( \5345 , \4744 , RIb556390_409);
and \U$4622 ( \5346 , RIb556480_411, \4763 );
nor \U$4623 ( \5347 , \5345 , \5346 );
and \U$4624 ( \5348 , RIb556318_408, \4746 );
and \U$4625 ( \5349 , RIb5562a0_407, \4730 );
and \U$4626 ( \5350 , \4738 , RIb5561b0_405);
and \U$4627 ( \5351 , RIb556228_406, \4732 );
nor \U$4628 ( \5352 , \5350 , \5351 );
not \U$4629 ( \5353 , \5352 );
nor \U$4630 ( \5354 , \5348 , \5349 , \5353 );
nand \U$4631 ( \5355 , \5344 , \5347 , \1879 , \5354 );
_DC r121c ( \5356_nR121c , \5355 , \4771 );
nand \U$4632 ( \5357 , \5356_nR121c , \4695 );
and \U$4633 ( \5358 , \5328 , \5357 );
and \U$4634 ( \5359 , \5167_nR140b , \4937 );
and \U$4635 ( \5360 , \4939 , \5261_nR12fd );
nand \U$4636 ( \5361 , \5167_nR140b , \4820 );
or \U$4637 ( \5362 , \4785 , \5261_nR12fd );
nand \U$4638 ( \5363 , \5362 , \4824 );
and \U$4639 ( \5364 , \5361 , \5363 );
nor \U$4640 ( \5365 , \5359 , \5360 , \5364 );
nor \U$4641 ( \5366 , \5358 , \5365 );
nand \U$4642 ( \5367 , \5321 , \5366 );
not \U$4643 ( \5368 , \5367 );
xor \U$4644 ( \5369 , \5215 , \5224 );
not \U$4645 ( \5370 , \5369 );
not \U$4646 ( \5371 , \5270 );
not \U$4647 ( \5372 , \5232 );
and \U$4648 ( \5373 , \5371 , \5372 );
and \U$4649 ( \5374 , \5270 , \5232 );
nor \U$4650 ( \5375 , \5373 , \5374 );
not \U$4651 ( \5376 , \5375 );
not \U$4652 ( \5377 , \5262 );
and \U$4653 ( \5378 , \5376 , \5377 );
and \U$4654 ( \5379 , \5375 , \5262 );
nor \U$4655 ( \5380 , \5378 , \5379 );
nor \U$4656 ( \5381 , \5370 , \5380 );
nand \U$4657 ( \5382 , \5368 , \5381 );
not \U$4658 ( \5383 , \5382 );
or \U$4659 ( \5384 , \5291 , \5383 );
or \U$4660 ( \5385 , \5188 , \5181 );
nand \U$4661 ( \5386 , \5385 , \5189 );
nand \U$4662 ( \5387 , \5384 , \5386 );
not \U$4663 ( \5388 , \5182 );
nand \U$4664 ( \5389 , \5388 , \5184 );
xor \U$4665 ( \5390 , \5387 , \5389 );
not \U$4666 ( \5391 , \5277 );
nor \U$4667 ( \5392 , \5391 , \5274 );
not \U$4668 ( \5393 , \5392 );
not \U$4669 ( \5394 , \5114 );
and \U$4670 ( \5395 , \5393 , \5394 );
and \U$4671 ( \5396 , \5392 , \5114 );
nor \U$4672 ( \5397 , \5395 , \5396 );
and \U$4673 ( \5398 , \5390 , \5397 );
and \U$4674 ( \5399 , \5387 , \5389 );
or \U$4675 ( \5400 , \5398 , \5399 );
xor \U$4676 ( \5401 , \5282 , \5400 );
not \U$4677 ( \5402 , \5261_nR12fd );
or \U$4678 ( \5403 , \4827 , \5402 );
not \U$4679 ( \5404 , \5356_nR121c );
or \U$4680 ( \5405 , \5404 , \4822 );
or \U$4681 ( \5406 , \4819 , \5402 );
or \U$4682 ( \5407 , \4785 , \5356_nR121c );
nand \U$4683 ( \5408 , \5407 , \4824 );
nand \U$4684 ( \5409 , \5406 , \5408 );
nand \U$4685 ( \5410 , \5403 , \5405 , \5409 );
and \U$4686 ( \5411 , \4968_nR171b , \5116 );
or \U$4687 ( \5412 , \4934 , \5028_nR162d );
nand \U$4688 ( \5413 , \5412 , \5073 );
nand \U$4689 ( \5414 , \4968_nR171b , \5068 );
and \U$4690 ( \5415 , \5413 , \5414 );
and \U$4691 ( \5416 , \5028_nR162d , \5070 );
nor \U$4692 ( \5417 , \5411 , \5415 , \5416 );
and \U$4693 ( \5418 , \5167_nR140b , \4885 );
and \U$4694 ( \5419 , \4921 , \5063_nR150e );
nand \U$4695 ( \5420 , \5167_nR140b , \4882 );
or \U$4696 ( \5421 , \4840 , \5063_nR150e );
nand \U$4697 ( \5422 , \5421 , \4925 );
and \U$4698 ( \5423 , \5420 , \5422 );
nor \U$4699 ( \5424 , \5418 , \5419 , \5423 );
nand \U$4700 ( \5425 , \5417 , \5424 );
and \U$4701 ( \5426 , \5410 , \5425 );
nor \U$4702 ( \5427 , \5424 , \5417 );
nor \U$4703 ( \5428 , \5426 , \5427 );
not \U$4704 ( \5429 , \5428 );
not \U$4705 ( \5430 , \5303 );
not \U$4706 ( \5431 , \5135 );
or \U$4707 ( \5432 , \5430 , \5431 );
or \U$4708 ( \5433 , \5135 , \5303 );
nand \U$4709 ( \5434 , \5432 , \5433 );
xor \U$4710 ( \5435 , \5305 , \5303 );
nor \U$4711 ( \5436 , \5434 , \5435 );
not \U$4712 ( \5437 , \5436 );
nor \U$4713 ( \5438 , \5437 , \5308 );
not \U$4714 ( \5439 , \5438 );
or \U$4715 ( \5440 , \5439 , \4816 );
or \U$4716 ( \5441 , \5437 , \4816 );
nand \U$4717 ( \5442 , \5441 , \5308 );
nand \U$4718 ( \5443 , \5440 , \5442 );
or \U$4719 ( \5444 , \5211 , \4871 );
not \U$4720 ( \5445 , \5297 );
or \U$4721 ( \5446 , \4773 , \5445 );
or \U$4722 ( \5447 , \5208 , \4871 );
or \U$4723 ( \5448 , \5137 , \4772_nR194f );
nand \U$4724 ( \5449 , \5448 , \5294 );
nand \U$4725 ( \5450 , \5447 , \5449 );
nand \U$4726 ( \5451 , \5444 , \5446 , \5450 );
and \U$4727 ( \5452 , \5443 , \5451 );
nand \U$4728 ( \5453 , \5429 , \5452 );
not \U$4729 ( \5454 , \5453 );
not \U$4730 ( \5455 , \5300 );
or \U$4731 ( \5456 , \5318 , \5307 );
nand \U$4732 ( \5457 , \5307 , \5318 );
nand \U$4733 ( \5458 , \5456 , \5457 );
not \U$4734 ( \5459 , \5458 );
or \U$4735 ( \5460 , \5455 , \5459 );
or \U$4736 ( \5461 , \5458 , \5300 );
nand \U$4737 ( \5462 , \5460 , \5461 );
not \U$4738 ( \5463 , \5357 );
not \U$4739 ( \5464 , \5365 );
not \U$4740 ( \5465 , \5328 );
and \U$4741 ( \5466 , \5464 , \5465 );
and \U$4742 ( \5467 , \5365 , \5328 );
nor \U$4743 ( \5468 , \5466 , \5467 );
not \U$4744 ( \5469 , \5468 );
or \U$4745 ( \5470 , \5463 , \5469 );
or \U$4746 ( \5471 , \5468 , \5357 );
nand \U$4747 ( \5472 , \5470 , \5471 );
and \U$4748 ( \5473 , \5462 , \5472 );
nand \U$4749 ( \5474 , \5454 , \5473 );
not \U$4750 ( \5475 , \5474 );
not \U$4751 ( \5476 , \5289 );
not \U$4752 ( \5477 , \5287 );
or \U$4753 ( \5478 , \5476 , \5477 );
or \U$4754 ( \5479 , \5287 , \5289 );
nand \U$4755 ( \5480 , \5478 , \5479 );
not \U$4756 ( \5481 , \5366 );
not \U$4757 ( \5482 , \5320 );
and \U$4758 ( \5483 , \5481 , \5482 );
and \U$4759 ( \5484 , \5366 , \5320 );
nor \U$4760 ( \5485 , \5483 , \5484 );
not \U$4761 ( \5486 , \5380 );
not \U$4762 ( \5487 , \5369 );
and \U$4763 ( \5488 , \5486 , \5487 );
and \U$4764 ( \5489 , \5380 , \5369 );
nor \U$4765 ( \5490 , \5488 , \5489 );
nand \U$4766 ( \5491 , \5485 , \5490 );
xor \U$4767 ( \5492 , \5480 , \5491 );
not \U$4768 ( \5493 , \5492 );
or \U$4769 ( \5494 , \5475 , \5493 );
or \U$4770 ( \5495 , \5492 , \5474 );
nand \U$4771 ( \5496 , \5494 , \5495 );
not \U$4772 ( \5497 , \5367 );
not \U$4773 ( \5498 , \5381 );
or \U$4774 ( \5499 , \5497 , \5498 );
or \U$4775 ( \5500 , \5381 , \5367 );
nand \U$4776 ( \5501 , \5499 , \5500 );
xor \U$4777 ( \5502 , \5496 , \5501 );
xor \U$4778 ( \5503 , \5462 , \5472 );
not \U$4779 ( \5504 , \5503 );
not \U$4780 ( \5505 , \5428 );
not \U$4781 ( \5506 , \5452 );
and \U$4782 ( \5507 , \5505 , \5506 );
and \U$4783 ( \5508 , \5428 , \5452 );
nor \U$4784 ( \5509 , \5507 , \5508 );
nor \U$4785 ( \5510 , \5504 , \5509 );
xor \U$4786 ( \5511 , \5443 , \5451 );
not \U$4787 ( \5512 , \5427 );
nand \U$4788 ( \5513 , \5512 , \5425 );
not \U$4789 ( \5514 , \5513 );
not \U$4790 ( \5515 , \5410 );
or \U$4791 ( \5516 , \5514 , \5515 );
or \U$4792 ( \5517 , \5410 , \5513 );
nand \U$4793 ( \5518 , \5516 , \5517 );
and \U$4794 ( \5519 , \5511 , \5518 );
and \U$4795 ( \5520 , \5307 , \5435 );
not \U$4796 ( \5521 , \5520 );
or \U$4797 ( \5522 , \5521 , \4816 );
or \U$4798 ( \5523 , \4773 , \5439 );
or \U$4799 ( \5524 , \5437 , \4773 );
or \U$4800 ( \5525 , \5307 , \4814_nR1a6c );
or \U$4801 ( \5526 , \5307 , \5435 );
nand \U$4802 ( \5527 , \5525 , \5526 );
nand \U$4803 ( \5528 , \5524 , \5527 );
nand \U$4804 ( \5529 , \5522 , \5523 , \5528 );
xor \U$4805 ( \5530 , \1098 , \4596_nRb9c );
xor \U$4806 ( \5531 , \5530 , \4661 );
not \U$4807 ( \5532 , \5531 );
xor \U$4808 ( \5533 , RIb54a900_11, \4626_nRa38 );
xor \U$4809 ( \5534 , \5533 , \4658 );
not \U$4810 ( \5535 , \5534 );
and \U$4811 ( \5536 , \5532 , \5535 );
nor \U$4812 ( \5537 , \5536 , \5305 );
not \U$4813 ( \5538 , \5537 );
xor \U$4814 ( \5539 , \5529 , \5538 );
not \U$4815 ( \5540 , \4968_nR171b );
or \U$4816 ( \5541 , \5211 , \5540 );
or \U$4817 ( \5542 , \4871 , \5445 );
or \U$4818 ( \5543 , \5208 , \5540 );
or \U$4819 ( \5544 , \5137 , \4870_nR1859 );
nand \U$4820 ( \5545 , \5544 , \5294 );
nand \U$4821 ( \5546 , \5543 , \5545 );
nand \U$4822 ( \5547 , \5541 , \5542 , \5546 );
and \U$4823 ( \5548 , \5539 , \5547 );
and \U$4824 ( \5549 , \5529 , \5538 );
or \U$4825 ( \5550 , \5548 , \5549 );
and \U$4826 ( \5551 , \5261_nR12fd , \4885 );
and \U$4827 ( \5552 , \4921 , \5167_nR140b );
nand \U$4828 ( \5553 , \5261_nR12fd , \4882 );
or \U$4829 ( \5554 , \4840 , \5167_nR140b );
nand \U$4830 ( \5555 , \5554 , \4925 );
and \U$4831 ( \5556 , \5553 , \5555 );
nor \U$4832 ( \5557 , \5551 , \5552 , \5556 );
and \U$4833 ( \5558 , \5028_nR162d , \5116 );
or \U$4834 ( \5559 , \4934 , \5063_nR150e );
nand \U$4835 ( \5560 , \5559 , \5073 );
nand \U$4836 ( \5561 , \5028_nR162d , \5068 );
and \U$4837 ( \5562 , \5560 , \5561 );
and \U$4838 ( \5563 , \5063_nR150e , \5070 );
nor \U$4839 ( \5564 , \5558 , \5562 , \5563 );
xor \U$4840 ( \5565 , \5557 , \5564 );
and \U$4841 ( \5566 , \5356_nR121c , \4937 );
and \U$4842 ( \5567 , RIb555e68_398, \4726 );
and \U$4843 ( \5568 , RIb5557d8_384, \4718 );
and \U$4844 ( \5569 , \4722 , RIb555ee0_399);
and \U$4845 ( \5570 , RIb555d00_395, \4756 );
nor \U$4846 ( \5571 , \5569 , \5570 );
and \U$4847 ( \5572 , \4744 , RIb555b98_392);
and \U$4848 ( \5573 , RIb555b20_391, \4746 );
nor \U$4849 ( \5574 , \5572 , \5573 );
and \U$4850 ( \5575 , \4738 , RIb5559b8_388);
and \U$4851 ( \5576 , RIb555940_387, \4740 );
nor \U$4852 ( \5577 , \5575 , \5576 );
and \U$4853 ( \5578 , \4730 , RIb555aa8_390);
and \U$4854 ( \5579 , RIb555a30_389, \4732 );
nor \U$4855 ( \5580 , \5578 , \5579 );
nand \U$4856 ( \5581 , \5571 , \5574 , \5577 , \5580 );
nor \U$4857 ( \5582 , \5567 , \5568 , \5581 );
and \U$4858 ( \5583 , \4754 , RIb555d78_396);
and \U$4859 ( \5584 , RIb555df0_397, \4714 );
nor \U$4860 ( \5585 , \5583 , \5584 );
nand \U$4861 ( \5586 , RIb555f58_400, \1269 );
and \U$4862 ( \5587 , RIb5558c8_386, \4759 );
and \U$4863 ( \5588 , RIb555850_385, \4761 );
and \U$4864 ( \5589 , \4763 , RIb555c88_394);
and \U$4865 ( \5590 , RIb555c10_393, \4765 );
nor \U$4866 ( \5591 , \5589 , \5590 );
not \U$4867 ( \5592 , \5591 );
nor \U$4868 ( \5593 , \5587 , \5588 , \5592 );
nand \U$4869 ( \5594 , \5582 , \5585 , \5586 , \5593 );
_DC r111a ( \5595_nR111a , \5594 , \4771 );
and \U$4870 ( \5596 , \4939 , \5595_nR111a );
nand \U$4871 ( \5597 , \5356_nR121c , \4820 );
or \U$4872 ( \5598 , \4785 , \5595_nR111a );
nand \U$4873 ( \5599 , \5598 , \4824 );
and \U$4874 ( \5600 , \5597 , \5599 );
nor \U$4875 ( \5601 , \5566 , \5596 , \5600 );
and \U$4876 ( \5602 , \5565 , \5601 );
and \U$4877 ( \5603 , \5557 , \5564 );
or \U$4878 ( \5604 , \5602 , \5603 );
not \U$4879 ( \5605 , \5604 );
and \U$4880 ( \5606 , \5550 , \5605 );
and \U$4881 ( \5607 , \5519 , \5606 );
xor \U$4882 ( \5608 , \5510 , \5607 );
or \U$4883 ( \5609 , \5490 , \5485 );
nand \U$4884 ( \5610 , \5609 , \5491 );
and \U$4885 ( \5611 , \5608 , \5610 );
and \U$4886 ( \5612 , \5510 , \5607 );
or \U$4887 ( \5613 , \5611 , \5612 );
and \U$4888 ( \5614 , \5502 , \5613 );
and \U$4889 ( \5615 , \5496 , \5501 );
or \U$4890 ( \5616 , \5614 , \5615 );
not \U$4891 ( \5617 , \5199 );
not \U$4892 ( \5618 , \5272 );
and \U$4893 ( \5619 , \5617 , \5618 );
and \U$4894 ( \5620 , \5199 , \5272 );
nor \U$4895 ( \5621 , \5619 , \5620 );
and \U$4896 ( \5622 , \5491 , \5480 );
not \U$4897 ( \5623 , \5491 );
not \U$4898 ( \5624 , \5480 );
and \U$4899 ( \5625 , \5623 , \5624 );
nor \U$4900 ( \5626 , \5625 , \5474 );
nor \U$4901 ( \5627 , \5622 , \5626 );
nand \U$4902 ( \5628 , \5621 , \5627 );
not \U$4903 ( \5629 , \5628 );
nor \U$4904 ( \5630 , \5627 , \5621 );
nor \U$4905 ( \5631 , \5629 , \5630 );
not \U$4906 ( \5632 , \5631 );
not \U$4907 ( \5633 , \5290 );
xnor \U$4908 ( \5634 , \5382 , \5386 );
not \U$4909 ( \5635 , \5634 );
or \U$4910 ( \5636 , \5633 , \5635 );
or \U$4911 ( \5637 , \5634 , \5290 );
nand \U$4912 ( \5638 , \5636 , \5637 );
not \U$4913 ( \5639 , \5638 );
and \U$4914 ( \5640 , \5632 , \5639 );
and \U$4915 ( \5641 , \5631 , \5638 );
nor \U$4916 ( \5642 , \5640 , \5641 );
xor \U$4917 ( \5643 , \5616 , \5642 );
not \U$4918 ( \5644 , \5453 );
not \U$4919 ( \5645 , \5473 );
or \U$4920 ( \5646 , \5644 , \5645 );
or \U$4921 ( \5647 , \5473 , \5453 );
nand \U$4922 ( \5648 , \5646 , \5647 );
not \U$4923 ( \5649 , \5648 );
xor \U$4924 ( \5650 , \5510 , \5607 );
xor \U$4925 ( \5651 , \5650 , \5610 );
not \U$4926 ( \5652 , \5503 );
not \U$4927 ( \5653 , \5509 );
and \U$4928 ( \5654 , \5652 , \5653 );
and \U$4929 ( \5655 , \5503 , \5509 );
nor \U$4930 ( \5656 , \5654 , \5655 );
xor \U$4931 ( \5657 , \5511 , \5518 );
nand \U$4932 ( \5658 , \5595_nR111a , \4695 );
and \U$4933 ( \5659 , \5657 , \5658 );
xor \U$4934 ( \5660 , \5550 , \5605 );
nor \U$4935 ( \5661 , \5659 , \5660 );
or \U$4936 ( \5662 , \5656 , \5661 );
not \U$4937 ( \5663 , \5661 );
not \U$4938 ( \5664 , \5656 );
or \U$4939 ( \5665 , \5663 , \5664 );
not \U$4940 ( \5666 , \5531 );
not \U$4941 ( \5667 , \5305 );
or \U$4942 ( \5668 , \5666 , \5667 );
or \U$4943 ( \5669 , \5305 , \5531 );
nand \U$4944 ( \5670 , \5668 , \5669 );
or \U$4945 ( \5671 , \5532 , \5534 );
or \U$4946 ( \5672 , \5535 , \5531 );
nand \U$4947 ( \5673 , \5671 , \5672 );
nor \U$4948 ( \5674 , \5670 , \5673 );
not \U$4949 ( \5675 , \5674 );
nor \U$4950 ( \5676 , \5675 , \5537 );
not \U$4951 ( \5677 , \5676 );
or \U$4952 ( \5678 , \5677 , \4816 );
or \U$4953 ( \5679 , \5675 , \4816 );
nand \U$4954 ( \5680 , \5679 , \5537 );
nand \U$4955 ( \5681 , \5678 , \5680 );
not \U$4956 ( \5682 , \5681 );
and \U$4957 ( \5683 , \4772_nR194f , \5520 );
or \U$4958 ( \5684 , \5307 , \4772_nR194f );
nand \U$4959 ( \5685 , \5684 , \5526 );
nand \U$4960 ( \5686 , \4870_nR1859 , \5436 );
and \U$4961 ( \5687 , \5685 , \5686 );
and \U$4962 ( \5688 , \4870_nR1859 , \5438 );
nor \U$4963 ( \5689 , \5683 , \5687 , \5688 );
nor \U$4964 ( \5690 , \5682 , \5689 );
not \U$4965 ( \5691 , \5690 );
and \U$4966 ( \5692 , \5063_nR150e , \5116 );
or \U$4967 ( \5693 , \4934 , \5167_nR140b );
nand \U$4968 ( \5694 , \5693 , \5073 );
nand \U$4969 ( \5695 , \5063_nR150e , \5068 );
and \U$4970 ( \5696 , \5694 , \5695 );
and \U$4971 ( \5697 , \5167_nR140b , \5070 );
nor \U$4972 ( \5698 , \5692 , \5696 , \5697 );
nand \U$4973 ( \5699 , \5028_nR162d , \5207 );
or \U$4974 ( \5700 , \5137 , \4968_nR171b );
nand \U$4975 ( \5701 , \5700 , \5294 );
and \U$4976 ( \5702 , \5699 , \5701 );
and \U$4977 ( \5703 , \5297 , \4968_nR171b );
and \U$4978 ( \5704 , \5028_nR162d , \5210 );
nor \U$4979 ( \5705 , \5702 , \5703 , \5704 );
xor \U$4980 ( \5706 , \5698 , \5705 );
and \U$4981 ( \5707 , \5356_nR121c , \4885 );
and \U$4982 ( \5708 , \4921 , \5261_nR12fd );
nand \U$4983 ( \5709 , \5356_nR121c , \4882 );
or \U$4984 ( \5710 , \4840 , \5261_nR12fd );
nand \U$4985 ( \5711 , \5710 , \4925 );
and \U$4986 ( \5712 , \5709 , \5711 );
nor \U$4987 ( \5713 , \5707 , \5708 , \5712 );
and \U$4988 ( \5714 , \5706 , \5713 );
and \U$4989 ( \5715 , \5698 , \5705 );
or \U$4990 ( \5716 , \5714 , \5715 );
nor \U$4991 ( \5717 , \5691 , \5716 );
not \U$4992 ( \5718 , \5717 );
and \U$4993 ( \5719 , RIb557128_438, \4740 );
and \U$4994 ( \5720 , RIb557650_449, \4726 );
and \U$4995 ( \5721 , \4754 , RIb557560_447);
and \U$4996 ( \5722 , RIb5574e8_446, \4756 );
nor \U$4997 ( \5723 , \5721 , \5722 );
and \U$4998 ( \5724 , \4759 , RIb5570b0_437);
and \U$4999 ( \5725 , RIb557038_436, \4761 );
nor \U$5000 ( \5726 , \5724 , \5725 );
and \U$5001 ( \5727 , \4722 , RIb5576c8_450);
and \U$5002 ( \5728 , RIb556fc0_435, \4718 );
nor \U$5003 ( \5729 , \5727 , \5728 );
and \U$5004 ( \5730 , \4763 , RIb557470_445);
and \U$5005 ( \5731 , RIb5573f8_444, \4765 );
nor \U$5006 ( \5732 , \5730 , \5731 );
nand \U$5007 ( \5733 , \5723 , \5726 , \5729 , \5732 );
nor \U$5008 ( \5734 , \5719 , \5720 , \5733 );
and \U$5009 ( \5735 , \4744 , RIb557380_443);
and \U$5010 ( \5736 , RIb5575d8_448, \4714 );
nor \U$5011 ( \5737 , \5735 , \5736 );
nand \U$5012 ( \5738 , RIb557740_451, \1269 );
and \U$5013 ( \5739 , RIb557308_442, \4746 );
and \U$5014 ( \5740 , RIb557290_441, \4730 );
and \U$5015 ( \5741 , \4738 , RIb5571a0_439);
and \U$5016 ( \5742 , RIb557218_440, \4732 );
nor \U$5017 ( \5743 , \5741 , \5742 );
not \U$5018 ( \5744 , \5743 );
nor \U$5019 ( \5745 , \5739 , \5740 , \5744 );
nand \U$5020 ( \5746 , \5734 , \5737 , \5738 , \5745 );
_DC r1037 ( \5747_nR1037 , \5746 , \4771 );
nand \U$5021 ( \5748 , \5747_nR1037 , \4695 );
not \U$5022 ( \5749 , \5748 );
xor \U$5023 ( \5750 , \5529 , \5538 );
xor \U$5024 ( \5751 , \5750 , \5547 );
xor \U$5025 ( \5752 , \5557 , \5564 );
xor \U$5026 ( \5753 , \5752 , \5601 );
not \U$5027 ( \5754 , \5753 );
and \U$5028 ( \5755 , \5751 , \5754 );
nor \U$5029 ( \5756 , \5749 , \5755 );
nor \U$5030 ( \5757 , \5718 , \5756 );
nand \U$5031 ( \5758 , \5665 , \5757 );
nand \U$5032 ( \5759 , \5662 , \5758 );
or \U$5033 ( \5760 , \5651 , \5759 );
not \U$5034 ( \5761 , \5760 );
or \U$5035 ( \5762 , \5649 , \5761 );
nand \U$5036 ( \5763 , \5759 , \5651 );
nand \U$5037 ( \5764 , \5762 , \5763 );
xor \U$5038 ( \5765 , \5496 , \5501 );
xor \U$5039 ( \5766 , \5765 , \5613 );
xor \U$5040 ( \5767 , \5764 , \5766 );
not \U$5041 ( \5768 , \5648 );
and \U$5042 ( \5769 , \5763 , \5760 );
not \U$5043 ( \5770 , \5769 );
or \U$5044 ( \5771 , \5768 , \5770 );
or \U$5045 ( \5772 , \5769 , \5648 );
nand \U$5046 ( \5773 , \5771 , \5772 );
not \U$5047 ( \5774 , \5757 );
not \U$5048 ( \5775 , \5661 );
and \U$5049 ( \5776 , \5774 , \5775 );
and \U$5050 ( \5777 , \5757 , \5661 );
nor \U$5051 ( \5778 , \5776 , \5777 );
xnor \U$5052 ( \5779 , \5778 , \5656 );
not \U$5053 ( \5780 , \5658 );
nor \U$5054 ( \5781 , \5780 , \5606 );
not \U$5055 ( \5782 , \5781 );
not \U$5056 ( \5783 , \5519 );
and \U$5057 ( \5784 , \5782 , \5783 );
and \U$5058 ( \5785 , \5781 , \5519 );
nor \U$5059 ( \5786 , \5784 , \5785 );
xor \U$5060 ( \5787 , \5779 , \5786 );
xor \U$5061 ( \5788 , \5751 , \5754 );
not \U$5062 ( \5789 , \5788 );
not \U$5063 ( \5790 , \5748 );
and \U$5064 ( \5791 , \5789 , \5790 );
and \U$5065 ( \5792 , \5788 , \5748 );
nor \U$5066 ( \5793 , \5791 , \5792 );
not \U$5067 ( \5794 , \5793 );
or \U$5068 ( \5795 , \5716 , \5690 );
and \U$5069 ( \5796 , RIb556930_421, \4740 );
and \U$5070 ( \5797 , RIb556ed0_433, \4722 );
and \U$5071 ( \5798 , \4754 , RIb556d68_430);
and \U$5072 ( \5799 , RIb556de0_431, \4714 );
nor \U$5073 ( \5800 , \5798 , \5799 );
and \U$5074 ( \5801 , \4759 , RIb5568b8_420);
and \U$5075 ( \5802 , RIb556840_419, \4761 );
nor \U$5076 ( \5803 , \5801 , \5802 );
and \U$5077 ( \5804 , \4726 , RIb556e58_432);
and \U$5078 ( \5805 , RIb5567c8_418, \4718 );
nor \U$5079 ( \5806 , \5804 , \5805 );
and \U$5080 ( \5807 , \4756 , RIb556cf0_429);
and \U$5081 ( \5808 , RIb556c78_428, \4763 );
nor \U$5082 ( \5809 , \5807 , \5808 );
nand \U$5083 ( \5810 , \5800 , \5803 , \5806 , \5809 );
nor \U$5084 ( \5811 , \5796 , \5797 , \5810 );
and \U$5085 ( \5812 , \4744 , RIb556b88_426);
and \U$5086 ( \5813 , RIb556c00_427, \4765 );
nor \U$5087 ( \5814 , \5812 , \5813 );
nand \U$5088 ( \5815 , RIb556f48_434, \1269 );
and \U$5089 ( \5816 , RIb556b10_425, \4746 );
and \U$5090 ( \5817 , RIb556a98_424, \4730 );
and \U$5091 ( \5818 , \4738 , RIb5569a8_422);
and \U$5092 ( \5819 , RIb556a20_423, \4732 );
nor \U$5093 ( \5820 , \5818 , \5819 );
not \U$5094 ( \5821 , \5820 );
nor \U$5095 ( \5822 , \5816 , \5817 , \5821 );
nand \U$5096 ( \5823 , \5811 , \5814 , \5815 , \5822 );
_DC rf5f ( \5824_nRf5f , \5823 , \4771 );
nand \U$5097 ( \5825 , \5824_nRf5f , \4695 );
and \U$5098 ( \5826 , \5595_nR111a , \4937 );
and \U$5099 ( \5827 , \4939 , \5747_nR1037 );
nand \U$5100 ( \5828 , \5595_nR111a , \4820 );
or \U$5101 ( \5829 , \4785 , \5747_nR1037 );
nand \U$5102 ( \5830 , \5829 , \4824 );
and \U$5103 ( \5831 , \5828 , \5830 );
nor \U$5104 ( \5832 , \5826 , \5827 , \5831 );
or \U$5105 ( \5833 , \5825 , \5832 );
nand \U$5106 ( \5834 , \5690 , \5716 );
nand \U$5107 ( \5835 , \5795 , \5833 , \5834 );
nand \U$5108 ( \5836 , \5794 , \5835 );
not \U$5109 ( \5837 , \5689 );
not \U$5110 ( \5838 , \5681 );
and \U$5111 ( \5839 , \5837 , \5838 );
and \U$5112 ( \5840 , \5689 , \5681 );
nor \U$5113 ( \5841 , \5839 , \5840 );
xor \U$5114 ( \5842 , \5698 , \5705 );
xor \U$5115 ( \5843 , \5842 , \5713 );
and \U$5116 ( \5844 , \5841 , \5843 );
xnor \U$5117 ( \5845 , \5825 , \5832 );
xor \U$5118 ( \5846 , \5698 , \5705 );
xor \U$5119 ( \5847 , \5846 , \5713 );
and \U$5120 ( \5848 , \5845 , \5847 );
and \U$5121 ( \5849 , \5841 , \5845 );
or \U$5122 ( \5850 , \5844 , \5848 , \5849 );
not \U$5123 ( \5851 , \5850 );
and \U$5124 ( \5852 , \5167_nR140b , \5116 );
or \U$5125 ( \5853 , \4934 , \5261_nR12fd );
nand \U$5126 ( \5854 , \5853 , \5073 );
nand \U$5127 ( \5855 , \5167_nR140b , \5068 );
and \U$5128 ( \5856 , \5854 , \5855 );
and \U$5129 ( \5857 , \5261_nR12fd , \5070 );
nor \U$5130 ( \5858 , \5852 , \5856 , \5857 );
nand \U$5131 ( \5859 , \5063_nR150e , \5207 );
or \U$5132 ( \5860 , \5137 , \5028_nR162d );
nand \U$5133 ( \5861 , \5860 , \5294 );
and \U$5134 ( \5862 , \5859 , \5861 );
and \U$5135 ( \5863 , \5297 , \5028_nR162d );
and \U$5136 ( \5864 , \5063_nR150e , \5210 );
nor \U$5137 ( \5865 , \5862 , \5863 , \5864 );
xor \U$5138 ( \5866 , \5858 , \5865 );
and \U$5139 ( \5867 , \5595_nR111a , \4885 );
and \U$5140 ( \5868 , \4921 , \5356_nR121c );
nand \U$5141 ( \5869 , \5595_nR111a , \4882 );
or \U$5142 ( \5870 , \4840 , \5356_nR121c );
nand \U$5143 ( \5871 , \5870 , \4925 );
and \U$5144 ( \5872 , \5869 , \5871 );
nor \U$5145 ( \5873 , \5867 , \5868 , \5872 );
and \U$5146 ( \5874 , \5866 , \5873 );
and \U$5147 ( \5875 , \5858 , \5865 );
or \U$5148 ( \5876 , \5874 , \5875 );
nand \U$5149 ( \5877 , \4772_nR194f , \5674 );
or \U$5150 ( \5878 , \5538 , \4814_nR1a6c );
or \U$5151 ( \5879 , \5538 , \5673 );
nand \U$5152 ( \5880 , \5878 , \5879 );
and \U$5153 ( \5881 , \5877 , \5880 );
and \U$5154 ( \5882 , \5538 , \5673 );
and \U$5155 ( \5883 , \5882 , \4814_nR1a6c );
and \U$5156 ( \5884 , \4772_nR194f , \5676 );
nor \U$5157 ( \5885 , \5881 , \5883 , \5884 );
xor \U$5158 ( \5886 , \5885 , \5535 );
and \U$5159 ( \5887 , \4870_nR1859 , \5520 );
or \U$5160 ( \5888 , \5307 , \4870_nR1859 );
nand \U$5161 ( \5889 , \5888 , \5526 );
nand \U$5162 ( \5890 , \4968_nR171b , \5436 );
and \U$5163 ( \5891 , \5889 , \5890 );
and \U$5164 ( \5892 , \4968_nR171b , \5438 );
nor \U$5165 ( \5893 , \5887 , \5891 , \5892 );
and \U$5166 ( \5894 , \5886 , \5893 );
and \U$5167 ( \5895 , \5885 , \5535 );
or \U$5168 ( \5896 , \5894 , \5895 );
nor \U$5169 ( \5897 , \5876 , \5896 );
nand \U$5170 ( \5898 , \5851 , \5897 );
xor \U$5171 ( \5899 , \5836 , \5898 );
xnor \U$5172 ( \5900 , \5658 , \5657 );
not \U$5173 ( \5901 , \5900 );
not \U$5174 ( \5902 , \5660 );
and \U$5175 ( \5903 , \5901 , \5902 );
and \U$5176 ( \5904 , \5900 , \5660 );
nor \U$5177 ( \5905 , \5903 , \5904 );
and \U$5178 ( \5906 , \5899 , \5905 );
and \U$5179 ( \5907 , \5836 , \5898 );
or \U$5180 ( \5908 , \5906 , \5907 );
and \U$5181 ( \5909 , \5787 , \5908 );
and \U$5182 ( \5910 , \5779 , \5786 );
or \U$5183 ( \5911 , \5909 , \5910 );
xor \U$5184 ( \5912 , \5773 , \5911 );
nand \U$5185 ( \5913 , \5167_nR140b , \5207 );
or \U$5186 ( \5914 , \5137 , \5063_nR150e );
nand \U$5187 ( \5915 , \5914 , \5294 );
and \U$5188 ( \5916 , \5913 , \5915 );
and \U$5189 ( \5917 , \5297 , \5063_nR150e );
and \U$5190 ( \5918 , \5167_nR140b , \5210 );
nor \U$5191 ( \5919 , \5916 , \5917 , \5918 );
and \U$5192 ( \5920 , \4968_nR171b , \5520 );
or \U$5193 ( \5921 , \5307 , \4968_nR171b );
nand \U$5194 ( \5922 , \5921 , \5526 );
nand \U$5195 ( \5923 , \5028_nR162d , \5436 );
and \U$5196 ( \5924 , \5922 , \5923 );
and \U$5197 ( \5925 , \5028_nR162d , \5438 );
nor \U$5198 ( \5926 , \5920 , \5924 , \5925 );
xor \U$5199 ( \5927 , \5919 , \5926 );
and \U$5200 ( \5928 , \5261_nR12fd , \5116 );
or \U$5201 ( \5929 , \4934 , \5356_nR121c );
nand \U$5202 ( \5930 , \5929 , \5073 );
nand \U$5203 ( \5931 , \5261_nR12fd , \5068 );
and \U$5204 ( \5932 , \5930 , \5931 );
and \U$5205 ( \5933 , \5356_nR121c , \5070 );
nor \U$5206 ( \5934 , \5928 , \5932 , \5933 );
and \U$5207 ( \5935 , \5927 , \5934 );
and \U$5208 ( \5936 , \5919 , \5926 );
or \U$5209 ( \5937 , \5935 , \5936 );
nand \U$5210 ( \5938 , \4870_nR1859 , \5674 );
or \U$5211 ( \5939 , \5538 , \4772_nR194f );
nand \U$5212 ( \5940 , \5939 , \5879 );
and \U$5213 ( \5941 , \5938 , \5940 );
and \U$5214 ( \5942 , \5882 , \4772_nR194f );
and \U$5215 ( \5943 , \4870_nR1859 , \5676 );
nor \U$5216 ( \5944 , \5941 , \5942 , \5943 );
not \U$5217 ( \5945 , \5944 );
or \U$5218 ( \5946 , \5534 , \4814_nR1a6c );
or \U$5219 ( \5947 , \1191 , \4656_nRa36 );
nand \U$5220 ( \5948 , \5947 , \4657 );
nor \U$5221 ( \5949 , \5534 , \5948 );
not \U$5222 ( \5950 , \5949 );
nand \U$5223 ( \5951 , \5535 , \5950 );
nand \U$5224 ( \5952 , \5946 , \5951 );
nand \U$5225 ( \5953 , \5945 , \5952 );
xor \U$5226 ( \5954 , \5937 , \5953 );
and \U$5227 ( \5955 , \5747_nR1037 , \4885 );
and \U$5228 ( \5956 , \4921 , \5595_nR111a );
nand \U$5229 ( \5957 , \5747_nR1037 , \4882 );
or \U$5230 ( \5958 , \4840 , \5595_nR111a );
nand \U$5231 ( \5959 , \5958 , \4925 );
and \U$5232 ( \5960 , \5957 , \5959 );
nor \U$5233 ( \5961 , \5955 , \5956 , \5960 );
and \U$5234 ( \5962 , RIb557998_456, \4738 );
and \U$5235 ( \5963 , RIb557ec0_467, \4722 );
and \U$5236 ( \5964 , \4714 , RIb557dd0_465);
and \U$5237 ( \5965 , RIb557ce0_463, \4756 );
nor \U$5238 ( \5966 , \5964 , \5965 );
and \U$5239 ( \5967 , \4740 , RIb557920_455);
and \U$5240 ( \5968 , RIb5578a8_454, \4759 );
nor \U$5241 ( \5969 , \5967 , \5968 );
and \U$5242 ( \5970 , \4718 , RIb5577b8_452);
and \U$5243 ( \5971 , RIb557830_453, \4761 );
nor \U$5244 ( \5972 , \5970 , \5971 );
and \U$5245 ( \5973 , \4763 , RIb557c68_462);
and \U$5246 ( \5974 , RIb557bf0_461, \4765 );
nor \U$5247 ( \5975 , \5973 , \5974 );
nand \U$5248 ( \5976 , \5966 , \5969 , \5972 , \5975 );
nor \U$5249 ( \5977 , \5962 , \5963 , \5976 );
and \U$5250 ( \5978 , \4726 , RIb557e48_466);
and \U$5251 ( \5979 , RIb557d58_464, \4754 );
nor \U$5252 ( \5980 , \5978 , \5979 );
and \U$5253 ( \5981 , RIb557b78_460, \4744 );
and \U$5254 ( \5982 , RIb557b00_459, \4746 );
and \U$5255 ( \5983 , \4730 , RIb557a88_458);
and \U$5256 ( \5984 , RIb557a10_457, \4732 );
nor \U$5257 ( \5985 , \5983 , \5984 );
not \U$5258 ( \5986 , \5985 );
nor \U$5259 ( \5987 , \5981 , \5982 , \5986 );
nand \U$5260 ( \5988 , \5977 , \5980 , \2554 , \5987 );
_DC rddd ( \5989_nRddd , \5988 , \4771 );
nand \U$5261 ( \5990 , \5989_nRddd , \4695 );
and \U$5262 ( \5991 , \5961 , \5990 );
and \U$5263 ( \5992 , \5824_nRf5f , \4937 );
and \U$5264 ( \5993 , RIb558118_472, \4740 );
and \U$5265 ( \5994 , RIb5585c8_482, \4714 );
and \U$5266 ( \5995 , \4722 , RIb5586b8_484);
and \U$5267 ( \5996 , RIb558640_483, \4726 );
nor \U$5268 ( \5997 , \5995 , \5996 );
and \U$5269 ( \5998 , \4738 , RIb558190_473);
and \U$5270 ( \5999 , RIb5580a0_471, \4759 );
nor \U$5271 ( \6000 , \5998 , \5999 );
and \U$5272 ( \6001 , \4718 , RIb557fb0_469);
and \U$5273 ( \6002 , RIb558028_470, \4761 );
nor \U$5274 ( \6003 , \6001 , \6002 );
and \U$5275 ( \6004 , \4756 , RIb5584d8_480);
and \U$5276 ( \6005 , RIb5583e8_478, \4765 );
nor \U$5277 ( \6006 , \6004 , \6005 );
nand \U$5278 ( \6007 , \5997 , \6000 , \6003 , \6006 );
nor \U$5279 ( \6008 , \5993 , \5994 , \6007 );
and \U$5280 ( \6009 , \4754 , RIb558550_481);
and \U$5281 ( \6010 , RIb558460_479, \4763 );
nor \U$5282 ( \6011 , \6009 , \6010 );
and \U$5283 ( \6012 , RIb558370_477, \4744 );
and \U$5284 ( \6013 , RIb5582f8_476, \4746 );
and \U$5285 ( \6014 , \4730 , RIb558280_475);
and \U$5286 ( \6015 , RIb558208_474, \4732 );
nor \U$5287 ( \6016 , \6014 , \6015 );
not \U$5288 ( \6017 , \6016 );
nor \U$5289 ( \6018 , \6012 , \6013 , \6017 );
nand \U$5290 ( \6019 , \6008 , \6011 , \2464 , \6018 );
_DC rea9 ( \6020_nRea9 , \6019 , \4771 );
and \U$5291 ( \6021 , \4939 , \6020_nRea9 );
nand \U$5292 ( \6022 , \5824_nRf5f , \4820 );
or \U$5293 ( \6023 , \4785 , \6020_nRea9 );
nand \U$5294 ( \6024 , \6023 , \4824 );
and \U$5295 ( \6025 , \6022 , \6024 );
nor \U$5296 ( \6026 , \5992 , \6021 , \6025 );
nor \U$5297 ( \6027 , \5991 , \6026 );
not \U$5298 ( \6028 , \6027 );
and \U$5299 ( \6029 , \5954 , \6028 );
and \U$5300 ( \6030 , \5937 , \5953 );
or \U$5301 ( \6031 , \6029 , \6030 );
nand \U$5302 ( \6032 , \6020_nRea9 , \4695 );
and \U$5303 ( \6033 , \5747_nR1037 , \4937 );
and \U$5304 ( \6034 , \4939 , \5824_nRf5f );
nand \U$5305 ( \6035 , \5747_nR1037 , \4820 );
or \U$5306 ( \6036 , \4785 , \5824_nRf5f );
nand \U$5307 ( \6037 , \6036 , \4824 );
and \U$5308 ( \6038 , \6035 , \6037 );
nor \U$5309 ( \6039 , \6033 , \6034 , \6038 );
xnor \U$5310 ( \6040 , \6032 , \6039 );
xor \U$5311 ( \6041 , \6031 , \6040 );
xor \U$5312 ( \6042 , \5698 , \5705 );
xor \U$5313 ( \6043 , \6042 , \5713 );
xor \U$5314 ( \6044 , \5841 , \5845 );
xor \U$5315 ( \6045 , \6043 , \6044 );
xor \U$5316 ( \6046 , \6041 , \6045 );
not \U$5317 ( \6047 , \6046 );
not \U$5318 ( \6048 , \5896 );
or \U$5319 ( \6049 , \5876 , \6048 );
or \U$5320 ( \6050 , \6032 , \6039 );
not \U$5321 ( \6051 , \5876 );
or \U$5322 ( \6052 , \5896 , \6051 );
nand \U$5323 ( \6053 , \6049 , \6050 , \6052 );
nand \U$5324 ( \6054 , \6047 , \6053 );
not \U$5325 ( \6055 , \6040 );
xor \U$5326 ( \6056 , \5885 , \5535 );
xor \U$5327 ( \6057 , \6056 , \5893 );
xor \U$5328 ( \6058 , \6055 , \6057 );
xor \U$5329 ( \6059 , \5937 , \5953 );
xor \U$5330 ( \6060 , \6059 , \6028 );
and \U$5331 ( \6061 , \6058 , \6060 );
and \U$5332 ( \6062 , \6055 , \6057 );
or \U$5333 ( \6063 , \6061 , \6062 );
xor \U$5334 ( \6064 , \5858 , \5865 );
xor \U$5335 ( \6065 , \6064 , \5873 );
nand \U$5336 ( \6066 , \4968_nR171b , \5674 );
or \U$5337 ( \6067 , \5538 , \4870_nR1859 );
nand \U$5338 ( \6068 , \6067 , \5879 );
and \U$5339 ( \6069 , \6066 , \6068 );
and \U$5340 ( \6070 , \5882 , \4870_nR1859 );
and \U$5341 ( \6071 , \4968_nR171b , \5676 );
nor \U$5342 ( \6072 , \6069 , \6070 , \6071 );
not \U$5343 ( \6073 , \5951 );
and \U$5344 ( \6074 , \4816 , \6073 );
and \U$5345 ( \6075 , \5949 , \4773 );
nand \U$5346 ( \6076 , \5948 , \5534 );
not \U$5347 ( \6077 , \6076 );
and \U$5348 ( \6078 , \4814_nR1a6c , \6077 );
nor \U$5349 ( \6079 , \6074 , \6075 , \6078 );
xor \U$5350 ( \6080 , \6072 , \6079 );
and \U$5351 ( \6081 , \5028_nR162d , \5520 );
or \U$5352 ( \6082 , \5307 , \5028_nR162d );
nand \U$5353 ( \6083 , \6082 , \5526 );
nand \U$5354 ( \6084 , \5063_nR150e , \5436 );
and \U$5355 ( \6085 , \6083 , \6084 );
and \U$5356 ( \6086 , \5063_nR150e , \5438 );
nor \U$5357 ( \6087 , \6081 , \6085 , \6086 );
and \U$5358 ( \6088 , \6080 , \6087 );
and \U$5359 ( \6089 , \6072 , \6079 );
or \U$5360 ( \6090 , \6088 , \6089 );
not \U$5361 ( \6091 , \6090 );
and \U$5362 ( \6092 , \5356_nR121c , \5116 );
or \U$5363 ( \6093 , \4934 , \5595_nR111a );
nand \U$5364 ( \6094 , \6093 , \5073 );
nand \U$5365 ( \6095 , \5356_nR121c , \5068 );
and \U$5366 ( \6096 , \6094 , \6095 );
and \U$5367 ( \6097 , \5595_nR111a , \5070 );
nor \U$5368 ( \6098 , \6092 , \6096 , \6097 );
nand \U$5369 ( \6099 , \5261_nR12fd , \5207 );
or \U$5370 ( \6100 , \5137 , \5167_nR140b );
nand \U$5371 ( \6101 , \6100 , \5294 );
and \U$5372 ( \6102 , \6099 , \6101 );
and \U$5373 ( \6103 , \5297 , \5167_nR140b );
and \U$5374 ( \6104 , \5261_nR12fd , \5210 );
nor \U$5375 ( \6105 , \6102 , \6103 , \6104 );
xor \U$5376 ( \6106 , \6098 , \6105 );
and \U$5377 ( \6107 , \5824_nRf5f , \4885 );
and \U$5378 ( \6108 , \4921 , \5747_nR1037 );
nand \U$5379 ( \6109 , \5824_nRf5f , \4882 );
or \U$5380 ( \6110 , \4840 , \5747_nR1037 );
nand \U$5381 ( \6111 , \6110 , \4925 );
and \U$5382 ( \6112 , \6109 , \6111 );
nor \U$5383 ( \6113 , \6107 , \6108 , \6112 );
and \U$5384 ( \6114 , \6106 , \6113 );
and \U$5385 ( \6115 , \6098 , \6105 );
or \U$5386 ( \6116 , \6114 , \6115 );
not \U$5387 ( \6117 , \6116 );
nand \U$5388 ( \6118 , \6091 , \6117 );
xor \U$5389 ( \6119 , \6065 , \6118 );
xor \U$5390 ( \6120 , \5919 , \5926 );
xor \U$5391 ( \6121 , \6120 , \5934 );
not \U$5392 ( \6122 , \6121 );
not \U$5393 ( \6123 , \5990 );
not \U$5394 ( \6124 , \6026 );
not \U$5395 ( \6125 , \5961 );
and \U$5396 ( \6126 , \6124 , \6125 );
and \U$5397 ( \6127 , \6026 , \5961 );
nor \U$5398 ( \6128 , \6126 , \6127 );
not \U$5399 ( \6129 , \6128 );
or \U$5400 ( \6130 , \6123 , \6129 );
or \U$5401 ( \6131 , \6128 , \5990 );
nand \U$5402 ( \6132 , \6130 , \6131 );
nand \U$5403 ( \6133 , \6122 , \6132 );
and \U$5404 ( \6134 , \6119 , \6133 );
and \U$5405 ( \6135 , \6065 , \6118 );
or \U$5406 ( \6136 , \6134 , \6135 );
and \U$5407 ( \6137 , \6063 , \6136 );
xor \U$5408 ( \6138 , \6054 , \6137 );
xor \U$5409 ( \6139 , \6031 , \6040 );
and \U$5410 ( \6140 , \6139 , \6045 );
and \U$5411 ( \6141 , \6031 , \6040 );
or \U$5412 ( \6142 , \6140 , \6141 );
not \U$5413 ( \6143 , \5850 );
not \U$5414 ( \6144 , \5897 );
and \U$5415 ( \6145 , \6143 , \6144 );
and \U$5416 ( \6146 , \5850 , \5897 );
nor \U$5417 ( \6147 , \6145 , \6146 );
xor \U$5418 ( \6148 , \6142 , \6147 );
not \U$5419 ( \6149 , \5793 );
not \U$5420 ( \6150 , \5835 );
and \U$5421 ( \6151 , \6149 , \6150 );
and \U$5422 ( \6152 , \5793 , \5835 );
nor \U$5423 ( \6153 , \6151 , \6152 );
xor \U$5424 ( \6154 , \6148 , \6153 );
and \U$5425 ( \6155 , \6138 , \6154 );
and \U$5426 ( \6156 , \6054 , \6137 );
or \U$5427 ( \6157 , \6155 , \6156 );
xor \U$5428 ( \6158 , \6142 , \6147 );
and \U$5429 ( \6159 , \6158 , \6153 );
and \U$5430 ( \6160 , \6142 , \6147 );
or \U$5431 ( \6161 , \6159 , \6160 );
not \U$5432 ( \6162 , \5756 );
not \U$5433 ( \6163 , \5717 );
and \U$5434 ( \6164 , \6162 , \6163 );
and \U$5435 ( \6165 , \5756 , \5717 );
nor \U$5436 ( \6166 , \6164 , \6165 );
xor \U$5437 ( \6167 , \6161 , \6166 );
xor \U$5438 ( \6168 , \5836 , \5898 );
xor \U$5439 ( \6169 , \6168 , \5905 );
xor \U$5440 ( \6170 , \6167 , \6169 );
and \U$5441 ( \6171 , \6157 , \6170 );
xor \U$5442 ( \6172 , \6063 , \6136 );
not \U$5443 ( \6173 , \6172 );
not \U$5444 ( \6174 , \5944 );
not \U$5445 ( \6175 , \5952 );
and \U$5446 ( \6176 , \6174 , \6175 );
and \U$5447 ( \6177 , \5944 , \5952 );
nor \U$5448 ( \6178 , \6176 , \6177 );
and \U$5449 ( \6179 , \6020_nRea9 , \4885 );
and \U$5450 ( \6180 , \4921 , \5824_nRf5f );
nand \U$5451 ( \6181 , \6020_nRea9 , \4882 );
or \U$5452 ( \6182 , \4840 , \5824_nRf5f );
nand \U$5453 ( \6183 , \6182 , \4925 );
and \U$5454 ( \6184 , \6181 , \6183 );
nor \U$5455 ( \6185 , \6179 , \6180 , \6184 );
and \U$5456 ( \6186 , RIb558910_489, \4740 );
and \U$5457 ( \6187 , RIb558eb0_501, \4722 );
and \U$5458 ( \6188 , \4754 , RIb558d48_498);
and \U$5459 ( \6189 , RIb558dc0_499, \4714 );
nor \U$5460 ( \6190 , \6188 , \6189 );
and \U$5461 ( \6191 , \4759 , RIb558898_488);
and \U$5462 ( \6192 , RIb558820_487, \4761 );
nor \U$5463 ( \6193 , \6191 , \6192 );
and \U$5464 ( \6194 , \4726 , RIb558e38_500);
and \U$5465 ( \6195 , RIb5587a8_486, \4718 );
nor \U$5466 ( \6196 , \6194 , \6195 );
and \U$5467 ( \6197 , \4763 , RIb558c58_496);
and \U$5468 ( \6198 , RIb558be0_495, \4765 );
nor \U$5469 ( \6199 , \6197 , \6198 );
nand \U$5470 ( \6200 , \6190 , \6193 , \6196 , \6199 );
nor \U$5471 ( \6201 , \6186 , \6187 , \6200 );
and \U$5472 ( \6202 , \4744 , RIb558b68_494);
and \U$5473 ( \6203 , RIb558cd0_497, \4756 );
nor \U$5474 ( \6204 , \6202 , \6203 );
nand \U$5475 ( \6205 , RIb558f28_502, \1269 );
and \U$5476 ( \6206 , RIb558af0_493, \4746 );
and \U$5477 ( \6207 , RIb558a78_492, \4730 );
and \U$5478 ( \6208 , \4738 , RIb558988_490);
and \U$5479 ( \6209 , RIb558a00_491, \4732 );
nor \U$5480 ( \6210 , \6208 , \6209 );
not \U$5481 ( \6211 , \6210 );
nor \U$5482 ( \6212 , \6206 , \6207 , \6211 );
nand \U$5483 ( \6213 , \6201 , \6204 , \6205 , \6212 );
_DC rca5 ( \6214_nRca5 , \6213 , \4771 );
nand \U$5484 ( \6215 , \6214_nRca5 , \4695 );
and \U$5485 ( \6216 , \6185 , \6215 );
and \U$5486 ( \6217 , \5989_nRddd , \4937 );
and \U$5487 ( \6218 , RIb5595b8_516, \4714 );
and \U$5488 ( \6219 , RIb558fa0_503, \4718 );
and \U$5489 ( \6220 , \4738 , RIb559180_507);
and \U$5490 ( \6221 , RIb5591f8_508, \4732 );
nor \U$5491 ( \6222 , \6220 , \6221 );
and \U$5492 ( \6223 , \4726 , RIb559630_517);
and \U$5493 ( \6224 , RIb559360_511, \4744 );
nor \U$5494 ( \6225 , \6223 , \6224 );
and \U$5495 ( \6226 , \4746 , RIb5592e8_510);
and \U$5496 ( \6227 , RIb559270_509, \4730 );
nor \U$5497 ( \6228 , \6226 , \6227 );
and \U$5498 ( \6229 , \4722 , RIb5596a8_518);
and \U$5499 ( \6230 , RIb5594c8_514, \4756 );
nor \U$5500 ( \6231 , \6229 , \6230 );
nand \U$5501 ( \6232 , \6222 , \6225 , \6228 , \6231 );
nor \U$5502 ( \6233 , \6218 , \6219 , \6232 );
and \U$5503 ( \6234 , \4754 , RIb559540_515);
and \U$5504 ( \6235 , RIb559450_513, \4763 );
nor \U$5505 ( \6236 , \6234 , \6235 );
and \U$5506 ( \6237 , RIb559090_505, \4759 );
and \U$5507 ( \6238 , RIb559018_504, \4761 );
and \U$5508 ( \6239 , \4765 , RIb5593d8_512);
and \U$5509 ( \6240 , RIb559108_506, \4740 );
nor \U$5510 ( \6241 , \6239 , \6240 );
not \U$5511 ( \6242 , \6241 );
nor \U$5512 ( \6243 , \6237 , \6238 , \6242 );
nand \U$5513 ( \6244 , \6233 , \6236 , \2748 , \6243 );
_DC rd47 ( \6245_nRd47 , \6244 , \4771 );
and \U$5514 ( \6246 , \4939 , \6245_nRd47 );
nand \U$5515 ( \6247 , \5989_nRddd , \4820 );
or \U$5516 ( \6248 , \4785 , \6245_nRd47 );
nand \U$5517 ( \6249 , \6248 , \4824 );
and \U$5518 ( \6250 , \6247 , \6249 );
nor \U$5519 ( \6251 , \6217 , \6246 , \6250 );
nor \U$5520 ( \6252 , \6216 , \6251 );
not \U$5521 ( \6253 , \6252 );
nand \U$5522 ( \6254 , \5356_nR121c , \5207 );
or \U$5523 ( \6255 , \5137 , \5261_nR12fd );
nand \U$5524 ( \6256 , \6255 , \5294 );
and \U$5525 ( \6257 , \6254 , \6256 );
and \U$5526 ( \6258 , \5297 , \5261_nR12fd );
and \U$5527 ( \6259 , \5356_nR121c , \5210 );
nor \U$5528 ( \6260 , \6257 , \6258 , \6259 );
and \U$5529 ( \6261 , \5063_nR150e , \5520 );
or \U$5530 ( \6262 , \5307 , \5063_nR150e );
nand \U$5531 ( \6263 , \6262 , \5526 );
nand \U$5532 ( \6264 , \5167_nR140b , \5436 );
and \U$5533 ( \6265 , \6263 , \6264 );
and \U$5534 ( \6266 , \5167_nR140b , \5438 );
nor \U$5535 ( \6267 , \6261 , \6265 , \6266 );
xor \U$5536 ( \6268 , \6260 , \6267 );
and \U$5537 ( \6269 , \5595_nR111a , \5116 );
or \U$5538 ( \6270 , \4934 , \5747_nR1037 );
nand \U$5539 ( \6271 , \6270 , \5073 );
nand \U$5540 ( \6272 , \5595_nR111a , \5068 );
and \U$5541 ( \6273 , \6271 , \6272 );
and \U$5542 ( \6274 , \5747_nR1037 , \5070 );
nor \U$5543 ( \6275 , \6269 , \6273 , \6274 );
and \U$5544 ( \6276 , \6268 , \6275 );
and \U$5545 ( \6277 , \6260 , \6267 );
or \U$5546 ( \6278 , \6276 , \6277 );
nand \U$5547 ( \6279 , \6253 , \6278 );
or \U$5548 ( \6280 , \6076 , \4773 );
or \U$5549 ( \6281 , \4772_nR194f , \5951 );
or \U$5550 ( \6282 , \4870_nR1859 , \5950 );
nand \U$5551 ( \6283 , \6280 , \6281 , \6282 );
or \U$5552 ( \6284 , \5677 , \5170 );
not \U$5553 ( \6285 , \5882 );
or \U$5554 ( \6286 , \5540 , \6285 );
or \U$5555 ( \6287 , \5675 , \5170 );
or \U$5556 ( \6288 , \5538 , \4968_nR171b );
nand \U$5557 ( \6289 , \6288 , \5879 );
nand \U$5558 ( \6290 , \6287 , \6289 );
nand \U$5559 ( \6291 , \6284 , \6286 , \6290 );
and \U$5560 ( \6292 , \6283 , \6291 );
and \U$5561 ( \6293 , \6279 , \6292 );
not \U$5562 ( \6294 , \6252 );
nor \U$5563 ( \6295 , \6294 , \6278 );
nor \U$5564 ( \6296 , \6293 , \6295 );
nand \U$5565 ( \6297 , \6178 , \6296 );
xor \U$5566 ( \6298 , \6098 , \6105 );
xor \U$5567 ( \6299 , \6298 , \6113 );
not \U$5568 ( \6300 , \6299 );
nand \U$5569 ( \6301 , \6245_nRd47 , \4695 );
and \U$5570 ( \6302 , \6020_nRea9 , \4937 );
and \U$5571 ( \6303 , \4939 , \5989_nRddd );
nand \U$5572 ( \6304 , \6020_nRea9 , \4820 );
or \U$5573 ( \6305 , \4785 , \5989_nRddd );
nand \U$5574 ( \6306 , \6305 , \4824 );
and \U$5575 ( \6307 , \6304 , \6306 );
nor \U$5576 ( \6308 , \6302 , \6303 , \6307 );
xor \U$5577 ( \6309 , \6301 , \6308 );
and \U$5578 ( \6310 , \6300 , \6309 );
and \U$5579 ( \6311 , \6297 , \6310 );
nor \U$5580 ( \6312 , \6296 , \6178 );
nor \U$5581 ( \6313 , \6311 , \6312 );
not \U$5582 ( \6314 , \6132 );
not \U$5583 ( \6315 , \6121 );
and \U$5584 ( \6316 , \6314 , \6315 );
and \U$5585 ( \6317 , \6132 , \6121 );
nor \U$5586 ( \6318 , \6316 , \6317 );
not \U$5587 ( \6319 , \6318 );
or \U$5588 ( \6320 , \6116 , \6091 );
or \U$5589 ( \6321 , \6301 , \6308 );
or \U$5590 ( \6322 , \6090 , \6117 );
nand \U$5591 ( \6323 , \6320 , \6321 , \6322 );
nand \U$5592 ( \6324 , \6319 , \6323 );
xor \U$5593 ( \6325 , \6313 , \6324 );
xor \U$5594 ( \6326 , \6055 , \6057 );
xor \U$5595 ( \6327 , \6326 , \6060 );
and \U$5596 ( \6328 , \6325 , \6327 );
and \U$5597 ( \6329 , \6313 , \6324 );
or \U$5598 ( \6330 , \6328 , \6329 );
not \U$5599 ( \6331 , \6330 );
not \U$5600 ( \6332 , \6053 );
not \U$5601 ( \6333 , \6046 );
or \U$5602 ( \6334 , \6332 , \6333 );
or \U$5603 ( \6335 , \6046 , \6053 );
nand \U$5604 ( \6336 , \6334 , \6335 );
nand \U$5605 ( \6337 , \6331 , \6336 );
not \U$5606 ( \6338 , \6337 );
or \U$5607 ( \6339 , \6173 , \6338 );
not \U$5608 ( \6340 , \6336 );
nand \U$5609 ( \6341 , \6340 , \6330 );
nand \U$5610 ( \6342 , \6339 , \6341 );
xor \U$5611 ( \6343 , \6054 , \6137 );
xor \U$5612 ( \6344 , \6343 , \6154 );
and \U$5613 ( \6345 , \6342 , \6344 );
nand \U$5614 ( \6346 , \6337 , \6341 );
not \U$5615 ( \6347 , \6346 );
not \U$5616 ( \6348 , \6172 );
and \U$5617 ( \6349 , \6347 , \6348 );
and \U$5618 ( \6350 , \6346 , \6172 );
nor \U$5619 ( \6351 , \6349 , \6350 );
xor \U$5620 ( \6352 , \6072 , \6079 );
xor \U$5621 ( \6353 , \6352 , \6087 );
not \U$5622 ( \6354 , \6353 );
and \U$5623 ( \6355 , \5747_nR1037 , \5116 );
or \U$5624 ( \6356 , \4934 , \5824_nRf5f );
nand \U$5625 ( \6357 , \6356 , \5073 );
nand \U$5626 ( \6358 , \5747_nR1037 , \5068 );
and \U$5627 ( \6359 , \6357 , \6358 );
and \U$5628 ( \6360 , \5824_nRf5f , \5070 );
nor \U$5629 ( \6361 , \6355 , \6359 , \6360 );
nand \U$5630 ( \6362 , \5595_nR111a , \5207 );
or \U$5631 ( \6363 , \5137 , \5356_nR121c );
nand \U$5632 ( \6364 , \6363 , \5294 );
and \U$5633 ( \6365 , \6362 , \6364 );
and \U$5634 ( \6366 , \5297 , \5356_nR121c );
and \U$5635 ( \6367 , \5595_nR111a , \5210 );
nor \U$5636 ( \6368 , \6365 , \6366 , \6367 );
xor \U$5637 ( \6369 , \6361 , \6368 );
and \U$5638 ( \6370 , \5989_nRddd , \4885 );
and \U$5639 ( \6371 , \4921 , \6020_nRea9 );
nand \U$5640 ( \6372 , \5989_nRddd , \4882 );
or \U$5641 ( \6373 , \4840 , \6020_nRea9 );
nand \U$5642 ( \6374 , \6373 , \4925 );
and \U$5643 ( \6375 , \6372 , \6374 );
nor \U$5644 ( \6376 , \6370 , \6371 , \6375 );
and \U$5645 ( \6377 , \6369 , \6376 );
and \U$5646 ( \6378 , \6361 , \6368 );
or \U$5647 ( \6379 , \6377 , \6378 );
nand \U$5648 ( \6380 , \5063_nR150e , \5674 );
or \U$5649 ( \6381 , \5538 , \5028_nR162d );
nand \U$5650 ( \6382 , \6381 , \5879 );
and \U$5651 ( \6383 , \6380 , \6382 );
and \U$5652 ( \6384 , \5882 , \5028_nR162d );
and \U$5653 ( \6385 , \5063_nR150e , \5676 );
nor \U$5654 ( \6386 , \6383 , \6384 , \6385 );
and \U$5655 ( \6387 , \4871 , \6073 );
and \U$5656 ( \6388 , \5949 , \5540 );
and \U$5657 ( \6389 , \4870_nR1859 , \6077 );
nor \U$5658 ( \6390 , \6387 , \6388 , \6389 );
xor \U$5659 ( \6391 , \6386 , \6390 );
and \U$5660 ( \6392 , \5167_nR140b , \5520 );
or \U$5661 ( \6393 , \5307 , \5167_nR140b );
nand \U$5662 ( \6394 , \6393 , \5526 );
nand \U$5663 ( \6395 , \5261_nR12fd , \5436 );
and \U$5664 ( \6396 , \6394 , \6395 );
and \U$5665 ( \6397 , \5261_nR12fd , \5438 );
nor \U$5666 ( \6398 , \6392 , \6396 , \6397 );
and \U$5667 ( \6399 , \6391 , \6398 );
and \U$5668 ( \6400 , \6386 , \6390 );
or \U$5669 ( \6401 , \6399 , \6400 );
nor \U$5670 ( \6402 , \6379 , \6401 );
nand \U$5671 ( \6403 , \6354 , \6402 );
not \U$5672 ( \6404 , \6318 );
not \U$5673 ( \6405 , \6323 );
and \U$5674 ( \6406 , \6404 , \6405 );
and \U$5675 ( \6407 , \6318 , \6323 );
nor \U$5676 ( \6408 , \6406 , \6407 );
nand \U$5677 ( \6409 , \6403 , \6408 );
not \U$5678 ( \6410 , \6310 );
not \U$5679 ( \6411 , \6312 );
nand \U$5680 ( \6412 , \6411 , \6297 );
not \U$5681 ( \6413 , \6412 );
or \U$5682 ( \6414 , \6410 , \6413 );
or \U$5683 ( \6415 , \6412 , \6310 );
nand \U$5684 ( \6416 , \6414 , \6415 );
and \U$5685 ( \6417 , \6409 , \6416 );
nor \U$5686 ( \6418 , \6408 , \6403 );
nor \U$5687 ( \6419 , \6417 , \6418 );
xor \U$5688 ( \6420 , \6065 , \6118 );
xor \U$5689 ( \6421 , \6420 , \6133 );
xor \U$5690 ( \6422 , \6419 , \6421 );
xor \U$5691 ( \6423 , \6313 , \6324 );
xor \U$5692 ( \6424 , \6423 , \6327 );
and \U$5693 ( \6425 , \6422 , \6424 );
and \U$5694 ( \6426 , \6419 , \6421 );
or \U$5695 ( \6427 , \6425 , \6426 );
not \U$5696 ( \6428 , \6427 );
and \U$5697 ( \6429 , \6351 , \6428 );
not \U$5698 ( \6430 , \6351 );
not \U$5699 ( \6431 , \6428 );
and \U$5700 ( \6432 , \6430 , \6431 );
xor \U$5701 ( \6433 , \6283 , \6291 );
not \U$5702 ( \6434 , \6401 );
or \U$5703 ( \6435 , \6379 , \6434 );
and \U$5704 ( \6436 , RIb55a620_551, \4726 );
and \U$5705 ( \6437 , RIb559f90_537, \4718 );
and \U$5706 ( \6438 , \4744 , RIb55a350_545);
and \U$5707 ( \6439 , RIb55a440_547, \4763 );
nor \U$5708 ( \6440 , \6438 , \6439 );
and \U$5709 ( \6441 , \4746 , RIb55a2d8_544);
and \U$5710 ( \6442 , RIb55a260_543, \4730 );
nor \U$5711 ( \6443 , \6441 , \6442 );
and \U$5712 ( \6444 , \4738 , RIb55a170_541);
and \U$5713 ( \6445 , RIb55a1e8_542, \4732 );
nor \U$5714 ( \6446 , \6444 , \6445 );
and \U$5715 ( \6447 , \4722 , RIb55a698_552);
and \U$5716 ( \6448 , RIb55a4b8_548, \4756 );
nor \U$5717 ( \6449 , \6447 , \6448 );
nand \U$5718 ( \6450 , \6440 , \6443 , \6446 , \6449 );
nor \U$5719 ( \6451 , \6436 , \6437 , \6450 );
and \U$5720 ( \6452 , \4754 , RIb55a530_549);
and \U$5721 ( \6453 , RIb55a5a8_550, \4714 );
nor \U$5722 ( \6454 , \6452 , \6453 );
and \U$5723 ( \6455 , RIb55a080_539, \4759 );
and \U$5724 ( \6456 , RIb55a008_538, \4761 );
and \U$5725 ( \6457 , \4765 , RIb55a3c8_546);
and \U$5726 ( \6458 , RIb55a0f8_540, \4740 );
nor \U$5727 ( \6459 , \6457 , \6458 );
not \U$5728 ( \6460 , \6459 );
nor \U$5729 ( \6461 , \6455 , \6456 , \6460 );
nand \U$5730 ( \6462 , \6451 , \6454 , \2994 , \6461 );
_DC rc21 ( \6463_nRc21 , \6462 , \4771 );
nand \U$5731 ( \6464 , \6463_nRc21 , \4695 );
and \U$5732 ( \6465 , \6245_nRd47 , \4937 );
and \U$5733 ( \6466 , \4939 , \6214_nRca5 );
nand \U$5734 ( \6467 , \6245_nRd47 , \4820 );
or \U$5735 ( \6468 , \4785 , \6214_nRca5 );
nand \U$5736 ( \6469 , \6468 , \4824 );
and \U$5737 ( \6470 , \6467 , \6469 );
nor \U$5738 ( \6471 , \6465 , \6466 , \6470 );
or \U$5739 ( \6472 , \6464 , \6471 );
not \U$5740 ( \6473 , \6379 );
or \U$5741 ( \6474 , \6401 , \6473 );
nand \U$5742 ( \6475 , \6435 , \6472 , \6474 );
xor \U$5743 ( \6476 , \6433 , \6475 );
not \U$5744 ( \6477 , \6215 );
not \U$5745 ( \6478 , \6251 );
not \U$5746 ( \6479 , \6185 );
and \U$5747 ( \6480 , \6478 , \6479 );
and \U$5748 ( \6481 , \6251 , \6185 );
nor \U$5749 ( \6482 , \6480 , \6481 );
not \U$5750 ( \6483 , \6482 );
or \U$5751 ( \6484 , \6477 , \6483 );
or \U$5752 ( \6485 , \6482 , \6215 );
nand \U$5753 ( \6486 , \6484 , \6485 );
xnor \U$5754 ( \6487 , \6476 , \6486 );
xor \U$5755 ( \6488 , \6361 , \6368 );
xor \U$5756 ( \6489 , \6488 , \6376 );
xor \U$5757 ( \6490 , \6386 , \6390 );
xor \U$5758 ( \6491 , \6490 , \6398 );
xor \U$5759 ( \6492 , \6489 , \6491 );
xnor \U$5760 ( \6493 , \6464 , \6471 );
and \U$5761 ( \6494 , \6492 , \6493 );
and \U$5762 ( \6495 , \6489 , \6491 );
or \U$5763 ( \6496 , \6494 , \6495 );
xor \U$5764 ( \6497 , \6260 , \6267 );
xor \U$5765 ( \6498 , \6497 , \6275 );
xor \U$5766 ( \6499 , \6496 , \6498 );
nand \U$5767 ( \6500 , \5747_nR1037 , \5207 );
or \U$5768 ( \6501 , \5137 , \5595_nR111a );
nand \U$5769 ( \6502 , \6501 , \5294 );
and \U$5770 ( \6503 , \6500 , \6502 );
and \U$5771 ( \6504 , \5297 , \5595_nR111a );
and \U$5772 ( \6505 , \5747_nR1037 , \5210 );
nor \U$5773 ( \6506 , \6503 , \6504 , \6505 );
and \U$5774 ( \6507 , \5261_nR12fd , \5520 );
or \U$5775 ( \6508 , \5307 , \5261_nR12fd );
nand \U$5776 ( \6509 , \6508 , \5526 );
nand \U$5777 ( \6510 , \5356_nR121c , \5436 );
and \U$5778 ( \6511 , \6509 , \6510 );
and \U$5779 ( \6512 , \5356_nR121c , \5438 );
nor \U$5780 ( \6513 , \6507 , \6511 , \6512 );
xor \U$5781 ( \6514 , \6506 , \6513 );
and \U$5782 ( \6515 , \5824_nRf5f , \5116 );
or \U$5783 ( \6516 , \4934 , \6020_nRea9 );
nand \U$5784 ( \6517 , \6516 , \5073 );
nand \U$5785 ( \6518 , \5824_nRf5f , \5068 );
and \U$5786 ( \6519 , \6517 , \6518 );
and \U$5787 ( \6520 , \6020_nRea9 , \5070 );
nor \U$5788 ( \6521 , \6515 , \6519 , \6520 );
and \U$5789 ( \6522 , \6514 , \6521 );
and \U$5790 ( \6523 , \6506 , \6513 );
or \U$5791 ( \6524 , \6522 , \6523 );
nand \U$5792 ( \6525 , \5167_nR140b , \5674 );
or \U$5793 ( \6526 , \5538 , \5063_nR150e );
nand \U$5794 ( \6527 , \6526 , \5879 );
and \U$5795 ( \6528 , \6525 , \6527 );
and \U$5796 ( \6529 , \5882 , \5063_nR150e );
and \U$5797 ( \6530 , \5167_nR140b , \5676 );
nor \U$5798 ( \6531 , \6528 , \6529 , \6530 );
not \U$5799 ( \6532 , \6531 );
or \U$5800 ( \6533 , \6076 , \5540 );
or \U$5801 ( \6534 , \4968_nR171b , \5951 );
or \U$5802 ( \6535 , \5028_nR162d , \5950 );
nand \U$5803 ( \6536 , \6533 , \6534 , \6535 );
nand \U$5804 ( \6537 , \6532 , \6536 );
xor \U$5805 ( \6538 , \6524 , \6537 );
and \U$5806 ( \6539 , \6245_nRd47 , \4885 );
and \U$5807 ( \6540 , \4921 , \5989_nRddd );
nand \U$5808 ( \6541 , \6245_nRd47 , \4882 );
or \U$5809 ( \6542 , \4840 , \5989_nRddd );
nand \U$5810 ( \6543 , \6542 , \4925 );
and \U$5811 ( \6544 , \6541 , \6543 );
nor \U$5812 ( \6545 , \6539 , \6540 , \6544 );
and \U$5813 ( \6546 , RIb559978_524, \4738 );
and \U$5814 ( \6547 , RIb559ea0_535, \4722 );
and \U$5815 ( \6548 , \4763 , RIb559c48_530);
and \U$5816 ( \6549 , RIb559bd0_529, \4765 );
nor \U$5817 ( \6550 , \6548 , \6549 );
and \U$5818 ( \6551 , \4740 , RIb559900_523);
and \U$5819 ( \6552 , RIb559888_522, \4759 );
nor \U$5820 ( \6553 , \6551 , \6552 );
and \U$5821 ( \6554 , \4718 , RIb559798_520);
and \U$5822 ( \6555 , RIb559810_521, \4761 );
nor \U$5823 ( \6556 , \6554 , \6555 );
and \U$5824 ( \6557 , \4754 , RIb559d38_532);
and \U$5825 ( \6558 , RIb559db0_533, \4714 );
nor \U$5826 ( \6559 , \6557 , \6558 );
nand \U$5827 ( \6560 , \6550 , \6553 , \6556 , \6559 );
nor \U$5828 ( \6561 , \6546 , \6547 , \6560 );
and \U$5829 ( \6562 , \4726 , RIb559e28_534);
and \U$5830 ( \6563 , RIb559cc0_531, \4756 );
nor \U$5831 ( \6564 , \6562 , \6563 );
and \U$5832 ( \6565 , RIb559b58_528, \4744 );
and \U$5833 ( \6566 , RIb559ae0_527, \4746 );
and \U$5834 ( \6567 , \4730 , RIb559a68_526);
and \U$5835 ( \6568 , RIb5599f0_525, \4732 );
nor \U$5836 ( \6569 , \6567 , \6568 );
not \U$5837 ( \6570 , \6569 );
nor \U$5838 ( \6571 , \6565 , \6566 , \6570 );
nand \U$5839 ( \6572 , \6561 , \6564 , \3111 , \6571 );
_DC rb98 ( \6573_nRb98 , \6572 , \4771 );
nand \U$5840 ( \6574 , \6573_nRb98 , \4695 );
and \U$5841 ( \6575 , \6545 , \6574 );
and \U$5842 ( \6576 , \6214_nRca5 , \4937 );
and \U$5843 ( \6577 , \4939 , \6463_nRc21 );
nand \U$5844 ( \6578 , \6214_nRca5 , \4820 );
or \U$5845 ( \6579 , \4785 , \6463_nRc21 );
nand \U$5846 ( \6580 , \6579 , \4824 );
and \U$5847 ( \6581 , \6578 , \6580 );
nor \U$5848 ( \6582 , \6576 , \6577 , \6581 );
nor \U$5849 ( \6583 , \6575 , \6582 );
not \U$5850 ( \6584 , \6583 );
and \U$5851 ( \6585 , \6538 , \6584 );
and \U$5852 ( \6586 , \6524 , \6537 );
or \U$5853 ( \6587 , \6585 , \6586 );
xor \U$5854 ( \6588 , \6499 , \6587 );
xor \U$5855 ( \6589 , \6487 , \6588 );
nand \U$5856 ( \6590 , \5261_nR12fd , \5674 );
or \U$5857 ( \6591 , \5538 , \5167_nR140b );
nand \U$5858 ( \6592 , \6591 , \5879 );
and \U$5859 ( \6593 , \6590 , \6592 );
and \U$5860 ( \6594 , \5882 , \5167_nR140b );
and \U$5861 ( \6595 , \5261_nR12fd , \5676 );
nor \U$5862 ( \6596 , \6593 , \6594 , \6595 );
and \U$5863 ( \6597 , \5170 , \6073 );
and \U$5864 ( \6598 , \5949 , \5172 );
and \U$5865 ( \6599 , \5028_nR162d , \6077 );
nor \U$5866 ( \6600 , \6597 , \6598 , \6599 );
xor \U$5867 ( \6601 , \6596 , \6600 );
and \U$5868 ( \6602 , \5356_nR121c , \5520 );
or \U$5869 ( \6603 , \5307 , \5356_nR121c );
nand \U$5870 ( \6604 , \6603 , \5526 );
nand \U$5871 ( \6605 , \5595_nR111a , \5436 );
and \U$5872 ( \6606 , \6604 , \6605 );
and \U$5873 ( \6607 , \5595_nR111a , \5438 );
nor \U$5874 ( \6608 , \6602 , \6606 , \6607 );
and \U$5875 ( \6609 , \6601 , \6608 );
and \U$5876 ( \6610 , \6596 , \6600 );
or \U$5877 ( \6611 , \6609 , \6610 );
not \U$5878 ( \6612 , \6611 );
and \U$5879 ( \6613 , \6020_nRea9 , \5116 );
or \U$5880 ( \6614 , \4934 , \5989_nRddd );
nand \U$5881 ( \6615 , \6614 , \5073 );
nand \U$5882 ( \6616 , \6020_nRea9 , \5068 );
and \U$5883 ( \6617 , \6615 , \6616 );
and \U$5884 ( \6618 , \5989_nRddd , \5070 );
nor \U$5885 ( \6619 , \6613 , \6617 , \6618 );
nand \U$5886 ( \6620 , \5824_nRf5f , \5207 );
or \U$5887 ( \6621 , \5137 , \5747_nR1037 );
nand \U$5888 ( \6622 , \6621 , \5294 );
and \U$5889 ( \6623 , \6620 , \6622 );
and \U$5890 ( \6624 , \5297 , \5747_nR1037 );
and \U$5891 ( \6625 , \5824_nRf5f , \5210 );
nor \U$5892 ( \6626 , \6623 , \6624 , \6625 );
xor \U$5893 ( \6627 , \6619 , \6626 );
and \U$5894 ( \6628 , \6214_nRca5 , \4885 );
and \U$5895 ( \6629 , \4921 , \6245_nRd47 );
nand \U$5896 ( \6630 , \6214_nRca5 , \4882 );
or \U$5897 ( \6631 , \4840 , \6245_nRd47 );
nand \U$5898 ( \6632 , \6631 , \4925 );
and \U$5899 ( \6633 , \6630 , \6632 );
nor \U$5900 ( \6634 , \6628 , \6629 , \6633 );
and \U$5901 ( \6635 , \6627 , \6634 );
and \U$5902 ( \6636 , \6619 , \6626 );
or \U$5903 ( \6637 , \6635 , \6636 );
not \U$5904 ( \6638 , \6637 );
nand \U$5905 ( \6639 , \6612 , \6638 );
xor \U$5906 ( \6640 , \6489 , \6491 );
xor \U$5907 ( \6641 , \6640 , \6493 );
and \U$5908 ( \6642 , \6639 , \6641 );
xor \U$5909 ( \6643 , \6506 , \6513 );
xor \U$5910 ( \6644 , \6643 , \6521 );
not \U$5911 ( \6645 , \6644 );
not \U$5912 ( \6646 , \6574 );
not \U$5913 ( \6647 , \6582 );
not \U$5914 ( \6648 , \6545 );
and \U$5915 ( \6649 , \6647 , \6648 );
and \U$5916 ( \6650 , \6582 , \6545 );
nor \U$5917 ( \6651 , \6649 , \6650 );
not \U$5918 ( \6652 , \6651 );
or \U$5919 ( \6653 , \6646 , \6652 );
or \U$5920 ( \6654 , \6651 , \6574 );
nand \U$5921 ( \6655 , \6653 , \6654 );
nand \U$5922 ( \6656 , \6645 , \6655 );
xor \U$5923 ( \6657 , \6489 , \6491 );
xor \U$5924 ( \6658 , \6657 , \6493 );
and \U$5925 ( \6659 , \6656 , \6658 );
and \U$5926 ( \6660 , \6639 , \6656 );
or \U$5927 ( \6661 , \6642 , \6659 , \6660 );
and \U$5928 ( \6662 , \6589 , \6661 );
and \U$5929 ( \6663 , \6487 , \6588 );
nor \U$5930 ( \6664 , \6662 , \6663 );
not \U$5931 ( \6665 , \6353 );
not \U$5932 ( \6666 , \6402 );
or \U$5933 ( \6667 , \6665 , \6666 );
or \U$5934 ( \6668 , \6402 , \6353 );
nand \U$5935 ( \6669 , \6667 , \6668 );
not \U$5936 ( \6670 , \6292 );
not \U$5937 ( \6671 , \6295 );
nand \U$5938 ( \6672 , \6671 , \6279 );
not \U$5939 ( \6673 , \6672 );
or \U$5940 ( \6674 , \6670 , \6673 );
or \U$5941 ( \6675 , \6672 , \6292 );
nand \U$5942 ( \6676 , \6674 , \6675 );
xor \U$5943 ( \6677 , \6669 , \6676 );
xor \U$5944 ( \6678 , \6664 , \6677 );
not \U$5945 ( \6679 , \6433 );
not \U$5946 ( \6680 , \6475 );
or \U$5947 ( \6681 , \6679 , \6680 );
or \U$5948 ( \6682 , \6475 , \6433 );
nand \U$5949 ( \6683 , \6682 , \6486 );
nand \U$5950 ( \6684 , \6681 , \6683 );
xor \U$5951 ( \6685 , \6300 , \6309 );
xor \U$5952 ( \6686 , \6684 , \6685 );
xor \U$5953 ( \6687 , \6496 , \6498 );
and \U$5954 ( \6688 , \6687 , \6587 );
and \U$5955 ( \6689 , \6496 , \6498 );
or \U$5956 ( \6690 , \6688 , \6689 );
not \U$5957 ( \6691 , \6690 );
xor \U$5958 ( \6692 , \6686 , \6691 );
and \U$5959 ( \6693 , \6678 , \6692 );
and \U$5960 ( \6694 , \6664 , \6677 );
or \U$5961 ( \6695 , \6693 , \6694 );
xor \U$5962 ( \6696 , \6684 , \6685 );
and \U$5963 ( \6697 , \6696 , \6691 );
and \U$5964 ( \6698 , \6684 , \6685 );
or \U$5965 ( \6699 , \6697 , \6698 );
and \U$5966 ( \6700 , \6669 , \6676 );
xor \U$5967 ( \6701 , \6699 , \6700 );
not \U$5968 ( \6702 , \6416 );
not \U$5969 ( \6703 , \6418 );
nand \U$5970 ( \6704 , \6703 , \6409 );
not \U$5971 ( \6705 , \6704 );
or \U$5972 ( \6706 , \6702 , \6705 );
or \U$5973 ( \6707 , \6704 , \6416 );
nand \U$5974 ( \6708 , \6706 , \6707 );
xor \U$5975 ( \6709 , \6701 , \6708 );
xor \U$5976 ( \6710 , \6695 , \6709 );
xor \U$5977 ( \6711 , \6664 , \6677 );
xor \U$5978 ( \6712 , \6711 , \6692 );
xor \U$5979 ( \6713 , \6487 , \6588 );
xor \U$5980 ( \6714 , \6713 , \6661 );
not \U$5981 ( \6715 , \6655 );
not \U$5982 ( \6716 , \6644 );
and \U$5983 ( \6717 , \6715 , \6716 );
and \U$5984 ( \6718 , \6655 , \6644 );
nor \U$5985 ( \6719 , \6717 , \6718 );
not \U$5986 ( \6720 , \6719 );
or \U$5987 ( \6721 , \6637 , \6612 );
and \U$5988 ( \6722 , RIb55a878_556, \4759 );
and \U$5989 ( \6723 , RIb55ae90_569, \4722 );
and \U$5990 ( \6724 , \4763 , RIb55ac38_564);
and \U$5991 ( \6725 , RIb55abc0_563, \4765 );
nor \U$5992 ( \6726 , \6724 , \6725 );
and \U$5993 ( \6727 , \4746 , RIb55aad0_561);
and \U$5994 ( \6728 , RIb55a8f0_557, \4740 );
nor \U$5995 ( \6729 , \6727 , \6728 );
and \U$5996 ( \6730 , \4718 , RIb55a788_554);
and \U$5997 ( \6731 , RIb55a800_555, \4761 );
nor \U$5998 ( \6732 , \6730 , \6731 );
and \U$5999 ( \6733 , \4726 , RIb55ae18_568);
and \U$6000 ( \6734 , RIb55ada0_567, \4714 );
nor \U$6001 ( \6735 , \6733 , \6734 );
nand \U$6002 ( \6736 , \6726 , \6729 , \6732 , \6735 );
nor \U$6003 ( \6737 , \6722 , \6723 , \6736 );
and \U$6004 ( \6738 , \4754 , RIb55ad28_566);
and \U$6005 ( \6739 , RIb55acb0_565, \4756 );
nor \U$6006 ( \6740 , \6738 , \6739 );
and \U$6007 ( \6741 , RIb55ab48_562, \4744 );
and \U$6008 ( \6742 , RIb55aa58_560, \4730 );
and \U$6009 ( \6743 , \4738 , RIb55a968_558);
and \U$6010 ( \6744 , RIb55a9e0_559, \4732 );
nor \U$6011 ( \6745 , \6743 , \6744 );
not \U$6012 ( \6746 , \6745 );
nor \U$6013 ( \6747 , \6741 , \6742 , \6746 );
nand \U$6014 ( \6748 , \6737 , \6740 , \3290 , \6747 );
_DC rb36 ( \6749_nRb36 , \6748 , \4771 );
nand \U$6015 ( \6750 , \6749_nRb36 , \4695 );
and \U$6016 ( \6751 , \6463_nRc21 , \4937 );
and \U$6017 ( \6752 , \4939 , \6573_nRb98 );
nand \U$6018 ( \6753 , \6463_nRc21 , \4820 );
or \U$6019 ( \6754 , \4785 , \6573_nRb98 );
nand \U$6020 ( \6755 , \6754 , \4824 );
and \U$6021 ( \6756 , \6753 , \6755 );
nor \U$6022 ( \6757 , \6751 , \6752 , \6756 );
or \U$6023 ( \6758 , \6750 , \6757 );
or \U$6024 ( \6759 , \6611 , \6638 );
nand \U$6025 ( \6760 , \6721 , \6758 , \6759 );
nand \U$6026 ( \6761 , \6720 , \6760 );
xor \U$6027 ( \6762 , \6524 , \6537 );
xor \U$6028 ( \6763 , \6762 , \6584 );
xor \U$6029 ( \6764 , \6761 , \6763 );
xor \U$6030 ( \6765 , \6619 , \6626 );
xor \U$6031 ( \6766 , \6765 , \6634 );
xor \U$6032 ( \6767 , \6596 , \6600 );
xor \U$6033 ( \6768 , \6767 , \6608 );
xor \U$6034 ( \6769 , \6766 , \6768 );
xnor \U$6035 ( \6770 , \6750 , \6757 );
and \U$6036 ( \6771 , \6769 , \6770 );
and \U$6037 ( \6772 , \6766 , \6768 );
or \U$6038 ( \6773 , \6771 , \6772 );
nand \U$6039 ( \6774 , \6020_nRea9 , \5207 );
or \U$6040 ( \6775 , \5137 , \5824_nRf5f );
nand \U$6041 ( \6776 , \6775 , \5294 );
and \U$6042 ( \6777 , \6774 , \6776 );
and \U$6043 ( \6778 , \5297 , \5824_nRf5f );
and \U$6044 ( \6779 , \6020_nRea9 , \5210 );
nor \U$6045 ( \6780 , \6777 , \6778 , \6779 );
and \U$6046 ( \6781 , \5595_nR111a , \5520 );
or \U$6047 ( \6782 , \5307 , \5595_nR111a );
nand \U$6048 ( \6783 , \6782 , \5526 );
nand \U$6049 ( \6784 , \5747_nR1037 , \5436 );
and \U$6050 ( \6785 , \6783 , \6784 );
and \U$6051 ( \6786 , \5747_nR1037 , \5438 );
nor \U$6052 ( \6787 , \6781 , \6785 , \6786 );
xor \U$6053 ( \6788 , \6780 , \6787 );
and \U$6054 ( \6789 , \5989_nRddd , \5116 );
or \U$6055 ( \6790 , \4934 , \6245_nRd47 );
nand \U$6056 ( \6791 , \6790 , \5073 );
nand \U$6057 ( \6792 , \5989_nRddd , \5068 );
and \U$6058 ( \6793 , \6791 , \6792 );
and \U$6059 ( \6794 , \6245_nRd47 , \5070 );
nor \U$6060 ( \6795 , \6789 , \6793 , \6794 );
and \U$6061 ( \6796 , \6788 , \6795 );
and \U$6062 ( \6797 , \6780 , \6787 );
or \U$6063 ( \6798 , \6796 , \6797 );
nand \U$6064 ( \6799 , \5356_nR121c , \5674 );
or \U$6065 ( \6800 , \5538 , \5261_nR12fd );
nand \U$6066 ( \6801 , \6800 , \5879 );
and \U$6067 ( \6802 , \6799 , \6801 );
and \U$6068 ( \6803 , \5882 , \5261_nR12fd );
and \U$6069 ( \6804 , \5356_nR121c , \5676 );
nor \U$6070 ( \6805 , \6802 , \6803 , \6804 );
not \U$6071 ( \6806 , \6805 );
or \U$6072 ( \6807 , \6076 , \5172 );
or \U$6073 ( \6808 , \5063_nR150e , \5951 );
or \U$6074 ( \6809 , \5167_nR140b , \5950 );
nand \U$6075 ( \6810 , \6807 , \6808 , \6809 );
nand \U$6076 ( \6811 , \6806 , \6810 );
xor \U$6077 ( \6812 , \6798 , \6811 );
and \U$6078 ( \6813 , \6463_nRc21 , \4885 );
and \U$6079 ( \6814 , \4921 , \6214_nRca5 );
nand \U$6080 ( \6815 , \6463_nRc21 , \4882 );
or \U$6081 ( \6816 , \4840 , \6214_nRca5 );
nand \U$6082 ( \6817 , \6816 , \4925 );
and \U$6083 ( \6818 , \6815 , \6817 );
nor \U$6084 ( \6819 , \6813 , \6814 , \6818 );
and \U$6085 ( \6820 , RIb55b160_575, \4738 );
and \U$6086 ( \6821 , RIb55b610_585, \4726 );
and \U$6087 ( \6822 , \4722 , RIb55b688_586);
and \U$6088 ( \6823 , RIb55b520_583, \4754 );
nor \U$6089 ( \6824 , \6822 , \6823 );
and \U$6090 ( \6825 , \4740 , RIb55b0e8_574);
and \U$6091 ( \6826 , RIb55b070_573, \4759 );
nor \U$6092 ( \6827 , \6825 , \6826 );
and \U$6093 ( \6828 , \4718 , RIb55af80_571);
and \U$6094 ( \6829 , RIb55aff8_572, \4761 );
nor \U$6095 ( \6830 , \6828 , \6829 );
and \U$6096 ( \6831 , \4756 , RIb55b4a8_582);
and \U$6097 ( \6832 , RIb55b430_581, \4763 );
nor \U$6098 ( \6833 , \6831 , \6832 );
nand \U$6099 ( \6834 , \6824 , \6827 , \6830 , \6833 );
nor \U$6100 ( \6835 , \6820 , \6821 , \6834 );
and \U$6101 ( \6836 , \4714 , RIb55b598_584);
and \U$6102 ( \6837 , RIb55b3b8_580, \4765 );
nor \U$6103 ( \6838 , \6836 , \6837 );
and \U$6104 ( \6839 , RIb55b340_579, \4744 );
and \U$6105 ( \6840 , RIb55b2c8_578, \4746 );
and \U$6106 ( \6841 , \4730 , RIb55b250_577);
and \U$6107 ( \6842 , RIb55b1d8_576, \4732 );
nor \U$6108 ( \6843 , \6841 , \6842 );
not \U$6109 ( \6844 , \6843 );
nor \U$6110 ( \6845 , \6839 , \6840 , \6844 );
nand \U$6111 ( \6846 , \6835 , \6838 , \3395 , \6845 );
_DC ra33 ( \6847_nRa33 , \6846 , \4771 );
nand \U$6112 ( \6848 , \6847_nRa33 , \4695 );
and \U$6113 ( \6849 , \6819 , \6848 );
and \U$6114 ( \6850 , \6573_nRb98 , \4937 );
and \U$6115 ( \6851 , \4939 , \6749_nRb36 );
nand \U$6116 ( \6852 , \6573_nRb98 , \4820 );
or \U$6117 ( \6853 , \4785 , \6749_nRb36 );
nand \U$6118 ( \6854 , \6853 , \4824 );
and \U$6119 ( \6855 , \6852 , \6854 );
nor \U$6120 ( \6856 , \6850 , \6851 , \6855 );
nor \U$6121 ( \6857 , \6849 , \6856 );
not \U$6122 ( \6858 , \6857 );
and \U$6123 ( \6859 , \6812 , \6858 );
and \U$6124 ( \6860 , \6798 , \6811 );
or \U$6125 ( \6861 , \6859 , \6860 );
nand \U$6126 ( \6862 , \6773 , \6861 );
not \U$6127 ( \6863 , \6536 );
not \U$6128 ( \6864 , \6531 );
or \U$6129 ( \6865 , \6863 , \6864 );
or \U$6130 ( \6866 , \6531 , \6536 );
nand \U$6131 ( \6867 , \6865 , \6866 );
and \U$6132 ( \6868 , \6862 , \6867 );
nor \U$6133 ( \6869 , \6861 , \6773 );
nor \U$6134 ( \6870 , \6868 , \6869 );
and \U$6135 ( \6871 , \6764 , \6870 );
and \U$6136 ( \6872 , \6761 , \6763 );
or \U$6137 ( \6873 , \6871 , \6872 );
nor \U$6138 ( \6874 , \6714 , \6873 );
xor \U$6139 ( \6875 , \6712 , \6874 );
and \U$6140 ( \6876 , \6714 , \6873 );
nor \U$6141 ( \6877 , \6876 , \6874 );
xor \U$6142 ( \6878 , \6761 , \6763 );
xor \U$6143 ( \6879 , \6878 , \6870 );
xor \U$6144 ( \6880 , \6489 , \6491 );
xor \U$6145 ( \6881 , \6880 , \6493 );
xor \U$6146 ( \6882 , \6639 , \6656 );
xor \U$6147 ( \6883 , \6881 , \6882 );
nor \U$6148 ( \6884 , \6879 , \6883 );
xor \U$6149 ( \6885 , \6877 , \6884 );
and \U$6150 ( \6886 , \6879 , \6883 );
nor \U$6151 ( \6887 , \6886 , \6884 );
not \U$6152 ( \6888 , \6760 );
not \U$6153 ( \6889 , \6719 );
or \U$6154 ( \6890 , \6888 , \6889 );
or \U$6155 ( \6891 , \6719 , \6760 );
nand \U$6156 ( \6892 , \6890 , \6891 );
not \U$6157 ( \6893 , \6867 );
not \U$6158 ( \6894 , \6869 );
nand \U$6159 ( \6895 , \6894 , \6862 );
not \U$6160 ( \6896 , \6895 );
or \U$6161 ( \6897 , \6893 , \6896 );
or \U$6162 ( \6898 , \6895 , \6867 );
nand \U$6163 ( \6899 , \6897 , \6898 );
nand \U$6164 ( \6900 , \6892 , \6899 );
xor \U$6165 ( \6901 , \6780 , \6787 );
xor \U$6166 ( \6902 , \6901 , \6795 );
not \U$6167 ( \6903 , \6902 );
not \U$6168 ( \6904 , \6810 );
not \U$6169 ( \6905 , \6805 );
or \U$6170 ( \6906 , \6904 , \6905 );
or \U$6171 ( \6907 , \6805 , \6810 );
nand \U$6172 ( \6908 , \6906 , \6907 );
nand \U$6173 ( \6909 , \6903 , \6908 );
xor \U$6174 ( \6910 , \6766 , \6768 );
xor \U$6175 ( \6911 , \6910 , \6770 );
and \U$6176 ( \6912 , \6909 , \6911 );
and \U$6177 ( \6913 , \6245_nRd47 , \5116 );
or \U$6178 ( \6914 , \4934 , \6214_nRca5 );
nand \U$6179 ( \6915 , \6914 , \5073 );
nand \U$6180 ( \6916 , \6245_nRd47 , \5068 );
and \U$6181 ( \6917 , \6915 , \6916 );
and \U$6182 ( \6918 , \6214_nRca5 , \5070 );
nor \U$6183 ( \6919 , \6913 , \6917 , \6918 );
nand \U$6184 ( \6920 , \5989_nRddd , \5207 );
or \U$6185 ( \6921 , \5137 , \6020_nRea9 );
nand \U$6186 ( \6922 , \6921 , \5294 );
and \U$6187 ( \6923 , \6920 , \6922 );
and \U$6188 ( \6924 , \5297 , \6020_nRea9 );
and \U$6189 ( \6925 , \5989_nRddd , \5210 );
nor \U$6190 ( \6926 , \6923 , \6924 , \6925 );
xor \U$6191 ( \6927 , \6919 , \6926 );
and \U$6192 ( \6928 , \6573_nRb98 , \4885 );
and \U$6193 ( \6929 , \4921 , \6463_nRc21 );
nand \U$6194 ( \6930 , \6573_nRb98 , \4882 );
or \U$6195 ( \6931 , \4840 , \6463_nRc21 );
nand \U$6196 ( \6932 , \6931 , \4925 );
and \U$6197 ( \6933 , \6930 , \6932 );
nor \U$6198 ( \6934 , \6928 , \6929 , \6933 );
and \U$6199 ( \6935 , \6927 , \6934 );
and \U$6200 ( \6936 , \6919 , \6926 );
or \U$6201 ( \6937 , \6935 , \6936 );
nand \U$6202 ( \6938 , \5595_nR111a , \5674 );
or \U$6203 ( \6939 , \5538 , \5356_nR121c );
nand \U$6204 ( \6940 , \6939 , \5879 );
and \U$6205 ( \6941 , \6938 , \6940 );
and \U$6206 ( \6942 , \5882 , \5356_nR121c );
and \U$6207 ( \6943 , \5595_nR111a , \5676 );
nor \U$6208 ( \6944 , \6941 , \6942 , \6943 );
and \U$6209 ( \6945 , \5168 , \6073 );
and \U$6210 ( \6946 , \5949 , \5402 );
and \U$6211 ( \6947 , \5167_nR140b , \6077 );
nor \U$6212 ( \6948 , \6945 , \6946 , \6947 );
xor \U$6213 ( \6949 , \6944 , \6948 );
and \U$6214 ( \6950 , \5747_nR1037 , \5520 );
or \U$6215 ( \6951 , \5307 , \5747_nR1037 );
nand \U$6216 ( \6952 , \6951 , \5526 );
nand \U$6217 ( \6953 , \5824_nRf5f , \5436 );
and \U$6218 ( \6954 , \6952 , \6953 );
and \U$6219 ( \6955 , \5824_nRf5f , \5438 );
nor \U$6220 ( \6956 , \6950 , \6954 , \6955 );
and \U$6221 ( \6957 , \6949 , \6956 );
and \U$6222 ( \6958 , \6944 , \6948 );
or \U$6223 ( \6959 , \6957 , \6958 );
xor \U$6224 ( \6960 , \6937 , \6959 );
not \U$6225 ( \6961 , \6856 );
not \U$6226 ( \6962 , \6819 );
and \U$6227 ( \6963 , \6961 , \6962 );
and \U$6228 ( \6964 , \6856 , \6819 );
nor \U$6229 ( \6965 , \6963 , \6964 );
not \U$6230 ( \6966 , \6965 );
not \U$6231 ( \6967 , \6848 );
and \U$6232 ( \6968 , \6966 , \6967 );
and \U$6233 ( \6969 , \6965 , \6848 );
nor \U$6234 ( \6970 , \6968 , \6969 );
and \U$6235 ( \6971 , \6960 , \6970 );
and \U$6236 ( \6972 , \6937 , \6959 );
or \U$6237 ( \6973 , \6971 , \6972 );
xor \U$6238 ( \6974 , \6766 , \6768 );
xor \U$6239 ( \6975 , \6974 , \6770 );
and \U$6240 ( \6976 , \6973 , \6975 );
and \U$6241 ( \6977 , \6909 , \6973 );
or \U$6242 ( \6978 , \6912 , \6976 , \6977 );
and \U$6243 ( \6979 , \6900 , \6978 );
nor \U$6244 ( \6980 , \6899 , \6892 );
nor \U$6245 ( \6981 , \6979 , \6980 );
xor \U$6246 ( \6982 , \6887 , \6981 );
not \U$6247 ( \6983 , \6978 );
not \U$6248 ( \6984 , \6980 );
nand \U$6249 ( \6985 , \6984 , \6900 );
not \U$6250 ( \6986 , \6985 );
or \U$6251 ( \6987 , \6983 , \6986 );
or \U$6252 ( \6988 , \6985 , \6978 );
nand \U$6253 ( \6989 , \6987 , \6988 );
not \U$6254 ( \6990 , \6749_nRb36 );
or \U$6255 ( \6991 , \4827 , \6990 );
not \U$6256 ( \6992 , \6847_nRa33 );
or \U$6257 ( \6993 , \6992 , \4822 );
or \U$6258 ( \6994 , \4819 , \6990 );
or \U$6259 ( \6995 , \4785 , \6847_nRa33 );
nand \U$6260 ( \6996 , \6995 , \4824 );
nand \U$6261 ( \6997 , \6994 , \6996 );
nand \U$6262 ( \6998 , \6991 , \6993 , \6997 );
nand \U$6263 ( \6999 , \6245_nRd47 , \5207 );
or \U$6264 ( \7000 , \5137 , \5989_nRddd );
nand \U$6265 ( \7001 , \7000 , \5294 );
and \U$6266 ( \7002 , \6999 , \7001 );
and \U$6267 ( \7003 , \5297 , \5989_nRddd );
and \U$6268 ( \7004 , \6245_nRd47 , \5210 );
nor \U$6269 ( \7005 , \7002 , \7003 , \7004 );
and \U$6270 ( \7006 , \5824_nRf5f , \5520 );
or \U$6271 ( \7007 , \5307 , \5824_nRf5f );
nand \U$6272 ( \7008 , \7007 , \5526 );
nand \U$6273 ( \7009 , \6020_nRea9 , \5436 );
and \U$6274 ( \7010 , \7008 , \7009 );
and \U$6275 ( \7011 , \6020_nRea9 , \5438 );
nor \U$6276 ( \7012 , \7006 , \7010 , \7011 );
xor \U$6277 ( \7013 , \7005 , \7012 );
and \U$6278 ( \7014 , \6214_nRca5 , \5116 );
or \U$6279 ( \7015 , \4934 , \6463_nRc21 );
nand \U$6280 ( \7016 , \7015 , \5073 );
nand \U$6281 ( \7017 , \6214_nRca5 , \5068 );
and \U$6282 ( \7018 , \7016 , \7017 );
and \U$6283 ( \7019 , \6463_nRc21 , \5070 );
nor \U$6284 ( \7020 , \7014 , \7018 , \7019 );
and \U$6285 ( \7021 , \7013 , \7020 );
and \U$6286 ( \7022 , \7005 , \7012 );
or \U$6287 ( \7023 , \7021 , \7022 );
nand \U$6288 ( \7024 , \5747_nR1037 , \5674 );
or \U$6289 ( \7025 , \5538 , \5595_nR111a );
nand \U$6290 ( \7026 , \7025 , \5879 );
and \U$6291 ( \7027 , \7024 , \7026 );
and \U$6292 ( \7028 , \5882 , \5595_nR111a );
and \U$6293 ( \7029 , \5747_nR1037 , \5676 );
nor \U$6294 ( \7030 , \7027 , \7028 , \7029 );
and \U$6295 ( \7031 , \5402 , \6073 );
and \U$6296 ( \7032 , \5949 , \5404 );
and \U$6297 ( \7033 , \5261_nR12fd , \6077 );
nor \U$6298 ( \7034 , \7031 , \7032 , \7033 );
xor \U$6299 ( \7035 , \7030 , \7034 );
and \U$6300 ( \7036 , \7035 , \4785 );
and \U$6301 ( \7037 , \7030 , \7034 );
or \U$6302 ( \7038 , \7036 , \7037 );
nand \U$6303 ( \7039 , \7023 , \7038 );
and \U$6304 ( \7040 , \6998 , \7039 );
nor \U$6305 ( \7041 , \7038 , \7023 );
nor \U$6306 ( \7042 , \7040 , \7041 );
not \U$6307 ( \7043 , \6902 );
not \U$6308 ( \7044 , \6908 );
and \U$6309 ( \7045 , \7043 , \7044 );
and \U$6310 ( \7046 , \6902 , \6908 );
nor \U$6311 ( \7047 , \7045 , \7046 );
xor \U$6312 ( \7048 , \7042 , \7047 );
xor \U$6313 ( \7049 , \6937 , \6959 );
xor \U$6314 ( \7050 , \7049 , \6970 );
and \U$6315 ( \7051 , \7048 , \7050 );
and \U$6316 ( \7052 , \7042 , \7047 );
or \U$6317 ( \7053 , \7051 , \7052 );
xor \U$6318 ( \7054 , \6798 , \6811 );
xor \U$6319 ( \7055 , \7054 , \6858 );
xor \U$6320 ( \7056 , \7053 , \7055 );
xor \U$6321 ( \7057 , \6766 , \6768 );
xor \U$6322 ( \7058 , \7057 , \6770 );
xor \U$6323 ( \7059 , \6909 , \6973 );
xor \U$6324 ( \7060 , \7058 , \7059 );
and \U$6325 ( \7061 , \7056 , \7060 );
and \U$6326 ( \7062 , \7053 , \7055 );
or \U$6327 ( \7063 , \7061 , \7062 );
xor \U$6328 ( \7064 , \6989 , \7063 );
xor \U$6329 ( \7065 , \6944 , \6948 );
xor \U$6330 ( \7066 , \7065 , \6956 );
not \U$6331 ( \7067 , \7066 );
not \U$6332 ( \7068 , \7041 );
nand \U$6333 ( \7069 , \7068 , \7039 );
not \U$6334 ( \7070 , \7069 );
not \U$6335 ( \7071 , \6998 );
or \U$6336 ( \7072 , \7070 , \7071 );
or \U$6337 ( \7073 , \6998 , \7069 );
nand \U$6338 ( \7074 , \7072 , \7073 );
nand \U$6339 ( \7075 , \7067 , \7074 );
and \U$6340 ( \7076 , \6749_nRb36 , \4885 );
and \U$6341 ( \7077 , \4921 , \6573_nRb98 );
nand \U$6342 ( \7078 , \6749_nRb36 , \4882 );
or \U$6343 ( \7079 , \4840 , \6573_nRb98 );
nand \U$6344 ( \7080 , \7079 , \4925 );
and \U$6345 ( \7081 , \7078 , \7080 );
nor \U$6346 ( \7082 , \7076 , \7077 , \7081 );
nand \U$6347 ( \7083 , \5824_nRf5f , \5674 );
or \U$6348 ( \7084 , \5538 , \5747_nR1037 );
nand \U$6349 ( \7085 , \7084 , \5879 );
and \U$6350 ( \7086 , \7083 , \7085 );
and \U$6351 ( \7087 , \5882 , \5747_nR1037 );
and \U$6352 ( \7088 , \5824_nRf5f , \5676 );
nor \U$6353 ( \7089 , \7086 , \7087 , \7088 );
and \U$6354 ( \7090 , \5404 , \6073 );
not \U$6355 ( \7091 , \5595_nR111a );
and \U$6356 ( \7092 , \5949 , \7091 );
and \U$6357 ( \7093 , \5356_nR121c , \6077 );
nor \U$6358 ( \7094 , \7090 , \7092 , \7093 );
xor \U$6359 ( \7095 , \7089 , \7094 );
and \U$6360 ( \7096 , \6020_nRea9 , \5520 );
or \U$6361 ( \7097 , \5307 , \6020_nRea9 );
nand \U$6362 ( \7098 , \7097 , \5526 );
nand \U$6363 ( \7099 , \5989_nRddd , \5436 );
and \U$6364 ( \7100 , \7098 , \7099 );
and \U$6365 ( \7101 , \5989_nRddd , \5438 );
nor \U$6366 ( \7102 , \7096 , \7100 , \7101 );
and \U$6367 ( \7103 , \7095 , \7102 );
and \U$6368 ( \7104 , \7089 , \7094 );
or \U$6369 ( \7105 , \7103 , \7104 );
xor \U$6370 ( \7106 , \7082 , \7105 );
and \U$6371 ( \7107 , \6463_nRc21 , \5116 );
or \U$6372 ( \7108 , \4934 , \6573_nRb98 );
nand \U$6373 ( \7109 , \7108 , \5073 );
nand \U$6374 ( \7110 , \6463_nRc21 , \5068 );
and \U$6375 ( \7111 , \7109 , \7110 );
and \U$6376 ( \7112 , \6573_nRb98 , \5070 );
nor \U$6377 ( \7113 , \7107 , \7111 , \7112 );
nand \U$6378 ( \7114 , \6214_nRca5 , \5207 );
or \U$6379 ( \7115 , \5137 , \6245_nRd47 );
nand \U$6380 ( \7116 , \7115 , \5294 );
and \U$6381 ( \7117 , \7114 , \7116 );
and \U$6382 ( \7118 , \5297 , \6245_nRd47 );
and \U$6383 ( \7119 , \6214_nRca5 , \5210 );
nor \U$6384 ( \7120 , \7117 , \7118 , \7119 );
xor \U$6385 ( \7121 , \7113 , \7120 );
and \U$6386 ( \7122 , \6847_nRa33 , \4885 );
and \U$6387 ( \7123 , \4921 , \6749_nRb36 );
nand \U$6388 ( \7124 , \6847_nRa33 , \4882 );
or \U$6389 ( \7125 , \4840 , \6749_nRb36 );
nand \U$6390 ( \7126 , \7125 , \4925 );
and \U$6391 ( \7127 , \7124 , \7126 );
nor \U$6392 ( \7128 , \7122 , \7123 , \7127 );
and \U$6393 ( \7129 , \7121 , \7128 );
and \U$6394 ( \7130 , \7113 , \7120 );
or \U$6395 ( \7131 , \7129 , \7130 );
and \U$6396 ( \7132 , \7106 , \7131 );
and \U$6397 ( \7133 , \7082 , \7105 );
or \U$6398 ( \7134 , \7132 , \7133 );
xor \U$6399 ( \7135 , \6919 , \6926 );
xor \U$6400 ( \7136 , \7135 , \6934 );
xor \U$6401 ( \7137 , \7134 , \7136 );
xor \U$6402 ( \7138 , \7005 , \7012 );
xor \U$6403 ( \7139 , \7138 , \7020 );
xor \U$6404 ( \7140 , \7030 , \7034 );
xor \U$6405 ( \7141 , \7140 , \4785 );
and \U$6406 ( \7142 , \7139 , \7141 );
nand \U$6407 ( \7143 , \6847_nRa33 , \4820 );
and \U$6408 ( \7144 , \4784 , \7143 );
and \U$6409 ( \7145 , \6847_nRa33 , \4937 );
nor \U$6410 ( \7146 , \7144 , \7145 );
xor \U$6411 ( \7147 , \7030 , \7034 );
xor \U$6412 ( \7148 , \7147 , \4785 );
and \U$6413 ( \7149 , \7146 , \7148 );
and \U$6414 ( \7150 , \7139 , \7146 );
or \U$6415 ( \7151 , \7142 , \7149 , \7150 );
and \U$6416 ( \7152 , \7137 , \7151 );
and \U$6417 ( \7153 , \7134 , \7136 );
or \U$6418 ( \7154 , \7152 , \7153 );
xor \U$6419 ( \7155 , \7075 , \7154 );
xor \U$6420 ( \7156 , \7042 , \7047 );
xor \U$6421 ( \7157 , \7156 , \7050 );
and \U$6422 ( \7158 , \7155 , \7157 );
and \U$6423 ( \7159 , \7075 , \7154 );
or \U$6424 ( \7160 , \7158 , \7159 );
xor \U$6425 ( \7161 , \7053 , \7055 );
xor \U$6426 ( \7162 , \7161 , \7060 );
and \U$6427 ( \7163 , \7160 , \7162 );
xor \U$6428 ( \7164 , \7134 , \7136 );
xor \U$6429 ( \7165 , \7164 , \7151 );
nand \U$6430 ( \7166 , \6463_nRc21 , \5207 );
or \U$6431 ( \7167 , \5137 , \6214_nRca5 );
nand \U$6432 ( \7168 , \7167 , \5294 );
and \U$6433 ( \7169 , \7166 , \7168 );
and \U$6434 ( \7170 , \5297 , \6214_nRca5 );
and \U$6435 ( \7171 , \6463_nRc21 , \5210 );
nor \U$6436 ( \7172 , \7169 , \7170 , \7171 );
and \U$6437 ( \7173 , \5989_nRddd , \5520 );
or \U$6438 ( \7174 , \5307 , \5989_nRddd );
nand \U$6439 ( \7175 , \7174 , \5526 );
nand \U$6440 ( \7176 , \6245_nRd47 , \5436 );
and \U$6441 ( \7177 , \7175 , \7176 );
and \U$6442 ( \7178 , \6245_nRd47 , \5438 );
nor \U$6443 ( \7179 , \7173 , \7177 , \7178 );
xor \U$6444 ( \7180 , \7172 , \7179 );
and \U$6445 ( \7181 , \6573_nRb98 , \5116 );
or \U$6446 ( \7182 , \4934 , \6749_nRb36 );
nand \U$6447 ( \7183 , \7182 , \5073 );
nand \U$6448 ( \7184 , \6573_nRb98 , \5068 );
and \U$6449 ( \7185 , \7183 , \7184 );
and \U$6450 ( \7186 , \6749_nRb36 , \5070 );
nor \U$6451 ( \7187 , \7181 , \7185 , \7186 );
and \U$6452 ( \7188 , \7180 , \7187 );
and \U$6453 ( \7189 , \7172 , \7179 );
or \U$6454 ( \7190 , \7188 , \7189 );
nand \U$6455 ( \7191 , \6020_nRea9 , \5674 );
or \U$6456 ( \7192 , \5538 , \5824_nRf5f );
nand \U$6457 ( \7193 , \7192 , \5879 );
and \U$6458 ( \7194 , \7191 , \7193 );
and \U$6459 ( \7195 , \5882 , \5824_nRf5f );
and \U$6460 ( \7196 , \6020_nRea9 , \5676 );
nor \U$6461 ( \7197 , \7194 , \7195 , \7196 );
and \U$6462 ( \7198 , \7091 , \6073 );
not \U$6463 ( \7199 , \5747_nR1037 );
and \U$6464 ( \7200 , \5949 , \7199 );
and \U$6465 ( \7201 , \5595_nR111a , \6077 );
nor \U$6466 ( \7202 , \7198 , \7200 , \7201 );
xor \U$6467 ( \7203 , \7197 , \7202 );
and \U$6468 ( \7204 , \7203 , \4840 );
and \U$6469 ( \7205 , \7197 , \7202 );
or \U$6470 ( \7206 , \7204 , \7205 );
xor \U$6471 ( \7207 , \7190 , \7206 );
xor \U$6472 ( \7208 , \7113 , \7120 );
xor \U$6473 ( \7209 , \7208 , \7128 );
and \U$6474 ( \7210 , \7207 , \7209 );
and \U$6475 ( \7211 , \7190 , \7206 );
or \U$6476 ( \7212 , \7210 , \7211 );
xor \U$6477 ( \7213 , \7082 , \7105 );
xor \U$6478 ( \7214 , \7213 , \7131 );
xor \U$6479 ( \7215 , \7212 , \7214 );
xor \U$6480 ( \7216 , \7030 , \7034 );
xor \U$6481 ( \7217 , \7216 , \4785 );
xor \U$6482 ( \7218 , \7139 , \7146 );
xor \U$6483 ( \7219 , \7217 , \7218 );
and \U$6484 ( \7220 , \7215 , \7219 );
and \U$6485 ( \7221 , \7212 , \7214 );
or \U$6486 ( \7222 , \7220 , \7221 );
not \U$6487 ( \7223 , \7074 );
not \U$6488 ( \7224 , \7066 );
and \U$6489 ( \7225 , \7223 , \7224 );
and \U$6490 ( \7226 , \7074 , \7066 );
nor \U$6491 ( \7227 , \7225 , \7226 );
xor \U$6492 ( \7228 , \7222 , \7227 );
xor \U$6493 ( \7229 , \7165 , \7228 );
not \U$6494 ( \7230 , \7229 );
xor \U$6495 ( \7231 , \7212 , \7214 );
xor \U$6496 ( \7232 , \7231 , \7219 );
nand \U$6497 ( \7233 , \5989_nRddd , \5674 );
or \U$6498 ( \7234 , \5538 , \6020_nRea9 );
nand \U$6499 ( \7235 , \7234 , \5879 );
and \U$6500 ( \7236 , \7233 , \7235 );
and \U$6501 ( \7237 , \5882 , \6020_nRea9 );
and \U$6502 ( \7238 , \5989_nRddd , \5676 );
nor \U$6503 ( \7239 , \7236 , \7237 , \7238 );
not \U$6504 ( \7240 , \7239 );
and \U$6505 ( \7241 , \7199 , \6073 );
not \U$6506 ( \7242 , \5824_nRf5f );
and \U$6507 ( \7243 , \5949 , \7242 );
and \U$6508 ( \7244 , \5747_nR1037 , \6077 );
nor \U$6509 ( \7245 , \7241 , \7243 , \7244 );
not \U$6510 ( \7246 , \7245 );
and \U$6511 ( \7247 , \7240 , \7246 );
and \U$6512 ( \7248 , \7239 , \7245 );
and \U$6513 ( \7249 , \6245_nRd47 , \5520 );
or \U$6514 ( \7250 , \5307 , \6245_nRd47 );
nand \U$6515 ( \7251 , \7250 , \5526 );
nand \U$6516 ( \7252 , \6214_nRca5 , \5436 );
and \U$6517 ( \7253 , \7251 , \7252 );
and \U$6518 ( \7254 , \6214_nRca5 , \5438 );
nor \U$6519 ( \7255 , \7249 , \7253 , \7254 );
nor \U$6520 ( \7256 , \7248 , \7255 );
nor \U$6521 ( \7257 , \7247 , \7256 );
xor \U$6522 ( \7258 , \7172 , \7179 );
xor \U$6523 ( \7259 , \7258 , \7187 );
and \U$6524 ( \7260 , \7257 , \7259 );
and \U$6525 ( \7261 , \6847_nRa33 , \4921 );
and \U$6526 ( \7262 , \6992 , \4884 );
not \U$6527 ( \7263 , \4925 );
nor \U$6528 ( \7264 , \7261 , \7262 , \7263 );
xor \U$6529 ( \7265 , \7172 , \7179 );
xor \U$6530 ( \7266 , \7265 , \7187 );
and \U$6531 ( \7267 , \7264 , \7266 );
and \U$6532 ( \7268 , \7257 , \7264 );
or \U$6533 ( \7269 , \7260 , \7267 , \7268 );
xor \U$6534 ( \7270 , \7089 , \7094 );
xor \U$6535 ( \7271 , \7270 , \7102 );
xor \U$6536 ( \7272 , \7269 , \7271 );
xor \U$6537 ( \7273 , \7190 , \7206 );
xor \U$6538 ( \7274 , \7273 , \7209 );
and \U$6539 ( \7275 , \7272 , \7274 );
and \U$6540 ( \7276 , \7269 , \7271 );
or \U$6541 ( \7277 , \7275 , \7276 );
nor \U$6542 ( \7278 , \7232 , \7277 );
xor \U$6543 ( \7279 , \7230 , \7278 );
and \U$6544 ( \7280 , \7232 , \7277 );
nor \U$6545 ( \7281 , \7280 , \7278 );
xor \U$6546 ( \7282 , \7269 , \7271 );
xor \U$6547 ( \7283 , \7282 , \7274 );
nand \U$6548 ( \7284 , \6245_nRd47 , \5674 );
or \U$6549 ( \7285 , \5538 , \5989_nRddd );
nand \U$6550 ( \7286 , \7285 , \5879 );
and \U$6551 ( \7287 , \7284 , \7286 );
and \U$6552 ( \7288 , \5882 , \5989_nRddd );
and \U$6553 ( \7289 , \6245_nRd47 , \5676 );
nor \U$6554 ( \7290 , \7287 , \7288 , \7289 );
and \U$6555 ( \7291 , \7242 , \6073 );
not \U$6556 ( \7292 , \6020_nRea9 );
and \U$6557 ( \7293 , \5949 , \7292 );
and \U$6558 ( \7294 , \5824_nRf5f , \6077 );
nor \U$6559 ( \7295 , \7291 , \7293 , \7294 );
xor \U$6560 ( \7296 , \7290 , \7295 );
and \U$6561 ( \7297 , \7296 , \4934 );
and \U$6562 ( \7298 , \7290 , \7295 );
or \U$6563 ( \7299 , \7297 , \7298 );
nand \U$6564 ( \7300 , \6573_nRb98 , \5207 );
or \U$6565 ( \7301 , \5137 , \6463_nRc21 );
nand \U$6566 ( \7302 , \7301 , \5294 );
and \U$6567 ( \7303 , \7300 , \7302 );
and \U$6568 ( \7304 , \5297 , \6463_nRc21 );
and \U$6569 ( \7305 , \6573_nRb98 , \5210 );
nor \U$6570 ( \7306 , \7303 , \7304 , \7305 );
xor \U$6571 ( \7307 , \7299 , \7306 );
nand \U$6572 ( \7308 , \6749_nRb36 , \5207 );
or \U$6573 ( \7309 , \5137 , \6573_nRb98 );
nand \U$6574 ( \7310 , \7309 , \5294 );
and \U$6575 ( \7311 , \7308 , \7310 );
and \U$6576 ( \7312 , \5297 , \6573_nRb98 );
and \U$6577 ( \7313 , \6749_nRb36 , \5210 );
nor \U$6578 ( \7314 , \7311 , \7312 , \7313 );
and \U$6579 ( \7315 , \6214_nRca5 , \5520 );
or \U$6580 ( \7316 , \5307 , \6214_nRca5 );
nand \U$6581 ( \7317 , \7316 , \5526 );
nand \U$6582 ( \7318 , \6463_nRc21 , \5436 );
and \U$6583 ( \7319 , \7317 , \7318 );
and \U$6584 ( \7320 , \6463_nRc21 , \5438 );
nor \U$6585 ( \7321 , \7315 , \7319 , \7320 );
xor \U$6586 ( \7322 , \7314 , \7321 );
and \U$6587 ( \7323 , \5116 , \6847_nRa33 );
nand \U$6588 ( \7324 , \6847_nRa33 , \5068 );
and \U$6589 ( \7325 , \7324 , \4935 );
nor \U$6590 ( \7326 , \7323 , \7325 );
and \U$6591 ( \7327 , \7322 , \7326 );
and \U$6592 ( \7328 , \7314 , \7321 );
or \U$6593 ( \7329 , \7327 , \7328 );
and \U$6594 ( \7330 , \7307 , \7329 );
and \U$6595 ( \7331 , \7299 , \7306 );
or \U$6596 ( \7332 , \7330 , \7331 );
xor \U$6597 ( \7333 , \7197 , \7202 );
xor \U$6598 ( \7334 , \7333 , \4840 );
nand \U$6599 ( \7335 , \7332 , \7334 );
not \U$6600 ( \7336 , \7239 );
xor \U$6601 ( \7337 , \7245 , \7255 );
not \U$6602 ( \7338 , \7337 );
or \U$6603 ( \7339 , \7336 , \7338 );
or \U$6604 ( \7340 , \7337 , \7239 );
nand \U$6605 ( \7341 , \7339 , \7340 );
or \U$6606 ( \7342 , \5216 , \6990 );
or \U$6607 ( \7343 , \6992 , \5218 );
or \U$6608 ( \7344 , \5115 , \6990 );
or \U$6609 ( \7345 , \4934 , \6847_nRa33 );
nand \U$6610 ( \7346 , \7345 , \5073 );
nand \U$6611 ( \7347 , \7344 , \7346 );
nand \U$6612 ( \7348 , \7342 , \7343 , \7347 );
and \U$6613 ( \7349 , \7341 , \7348 );
and \U$6614 ( \7350 , \7335 , \7349 );
nor \U$6615 ( \7351 , \7334 , \7332 );
nor \U$6616 ( \7352 , \7350 , \7351 );
nor \U$6617 ( \7353 , \7283 , \7352 );
xor \U$6618 ( \7354 , \7281 , \7353 );
not \U$6619 ( \7355 , \7349 );
not \U$6620 ( \7356 , \7351 );
nand \U$6621 ( \7357 , \7356 , \7335 );
not \U$6622 ( \7358 , \7357 );
or \U$6623 ( \7359 , \7355 , \7358 );
or \U$6624 ( \7360 , \7357 , \7349 );
nand \U$6625 ( \7361 , \7359 , \7360 );
xor \U$6626 ( \7362 , \7172 , \7179 );
xor \U$6627 ( \7363 , \7362 , \7187 );
xor \U$6628 ( \7364 , \7257 , \7264 );
xor \U$6629 ( \7365 , \7363 , \7364 );
not \U$6630 ( \7366 , \7365 );
xor \U$6631 ( \7367 , \7361 , \7366 );
xor \U$6632 ( \7368 , \7299 , \7306 );
xor \U$6633 ( \7369 , \7368 , \7329 );
nand \U$6634 ( \7370 , \6214_nRca5 , \5674 );
or \U$6635 ( \7371 , \5538 , \6245_nRd47 );
nand \U$6636 ( \7372 , \7371 , \5879 );
and \U$6637 ( \7373 , \7370 , \7372 );
and \U$6638 ( \7374 , \5882 , \6245_nRd47 );
and \U$6639 ( \7375 , \6214_nRca5 , \5676 );
nor \U$6640 ( \7376 , \7373 , \7374 , \7375 );
and \U$6641 ( \7377 , \7292 , \6073 );
not \U$6642 ( \7378 , \5989_nRddd );
and \U$6643 ( \7379 , \5949 , \7378 );
and \U$6644 ( \7380 , \6020_nRea9 , \6077 );
nor \U$6645 ( \7381 , \7377 , \7379 , \7380 );
xor \U$6646 ( \7382 , \7376 , \7381 );
and \U$6647 ( \7383 , \6463_nRc21 , \5520 );
or \U$6648 ( \7384 , \5307 , \6463_nRc21 );
nand \U$6649 ( \7385 , \7384 , \5526 );
nand \U$6650 ( \7386 , \6573_nRb98 , \5436 );
and \U$6651 ( \7387 , \7385 , \7386 );
and \U$6652 ( \7388 , \6573_nRb98 , \5438 );
nor \U$6653 ( \7389 , \7383 , \7387 , \7388 );
and \U$6654 ( \7390 , \7382 , \7389 );
and \U$6655 ( \7391 , \7376 , \7381 );
or \U$6656 ( \7392 , \7390 , \7391 );
xor \U$6657 ( \7393 , \7290 , \7295 );
xor \U$6658 ( \7394 , \7393 , \4934 );
and \U$6659 ( \7395 , \7392 , \7394 );
xor \U$6660 ( \7396 , \7314 , \7321 );
xor \U$6661 ( \7397 , \7396 , \7326 );
xor \U$6662 ( \7398 , \7290 , \7295 );
xor \U$6663 ( \7399 , \7398 , \4934 );
and \U$6664 ( \7400 , \7397 , \7399 );
and \U$6665 ( \7401 , \7392 , \7397 );
or \U$6666 ( \7402 , \7395 , \7400 , \7401 );
nand \U$6667 ( \7403 , \7369 , \7402 );
xor \U$6668 ( \7404 , \7341 , \7348 );
and \U$6669 ( \7405 , \7403 , \7404 );
nor \U$6670 ( \7406 , \7402 , \7369 );
nor \U$6671 ( \7407 , \7405 , \7406 );
not \U$6672 ( \7408 , \7407 );
xor \U$6673 ( \7409 , \7367 , \7408 );
not \U$6674 ( \7410 , \7403 );
nor \U$6675 ( \7411 , \7410 , \7406 );
not \U$6676 ( \7412 , \7411 );
not \U$6677 ( \7413 , \7404 );
and \U$6678 ( \7414 , \7412 , \7413 );
and \U$6679 ( \7415 , \7411 , \7404 );
nor \U$6680 ( \7416 , \7414 , \7415 );
xor \U$6681 ( \7417 , \7290 , \7295 );
xor \U$6682 ( \7418 , \7417 , \4934 );
xor \U$6683 ( \7419 , \7392 , \7397 );
xor \U$6684 ( \7420 , \7418 , \7419 );
nand \U$6685 ( \7421 , \6847_nRa33 , \5207 );
or \U$6686 ( \7422 , \5137 , \6749_nRb36 );
nand \U$6687 ( \7423 , \7422 , \5294 );
and \U$6688 ( \7424 , \7421 , \7423 );
and \U$6689 ( \7425 , \5297 , \6749_nRb36 );
and \U$6690 ( \7426 , \6847_nRa33 , \5210 );
nor \U$6691 ( \7427 , \7424 , \7425 , \7426 );
nand \U$6692 ( \7428 , \6463_nRc21 , \5674 );
or \U$6693 ( \7429 , \5538 , \6214_nRca5 );
nand \U$6694 ( \7430 , \7429 , \5879 );
and \U$6695 ( \7431 , \7428 , \7430 );
and \U$6696 ( \7432 , \5882 , \6214_nRca5 );
and \U$6697 ( \7433 , \6463_nRc21 , \5676 );
nor \U$6698 ( \7434 , \7431 , \7432 , \7433 );
and \U$6699 ( \7435 , \7378 , \6073 );
not \U$6700 ( \7436 , \6245_nRd47 );
and \U$6701 ( \7437 , \5949 , \7436 );
and \U$6702 ( \7438 , \5989_nRddd , \6077 );
nor \U$6703 ( \7439 , \7435 , \7437 , \7438 );
xor \U$6704 ( \7440 , \7434 , \7439 );
and \U$6705 ( \7441 , \7440 , \5137 );
and \U$6706 ( \7442 , \7434 , \7439 );
or \U$6707 ( \7443 , \7441 , \7442 );
xor \U$6708 ( \7444 , \7427 , \7443 );
and \U$6709 ( \7445 , \6573_nRb98 , \5520 );
or \U$6710 ( \7446 , \5307 , \6573_nRb98 );
nand \U$6711 ( \7447 , \7446 , \5526 );
nand \U$6712 ( \7448 , \6749_nRb36 , \5436 );
and \U$6713 ( \7449 , \7447 , \7448 );
and \U$6714 ( \7450 , \6749_nRb36 , \5438 );
nor \U$6715 ( \7451 , \7445 , \7449 , \7450 );
not \U$6716 ( \7452 , \7451 );
or \U$6717 ( \7453 , \5445 , \6992 );
or \U$6718 ( \7454 , \6847_nRa33 , \5137 );
nand \U$6719 ( \7455 , \7453 , \7454 , \5294 );
nand \U$6720 ( \7456 , \7452 , \7455 );
and \U$6721 ( \7457 , \7444 , \7456 );
and \U$6722 ( \7458 , \7427 , \7443 );
or \U$6723 ( \7459 , \7457 , \7458 );
nor \U$6724 ( \7460 , \7420 , \7459 );
xor \U$6725 ( \7461 , \7416 , \7460 );
not \U$6726 ( \7462 , \6573_nRb98 );
or \U$6727 ( \7463 , \6076 , \7462 );
or \U$6728 ( \7464 , \6573_nRb98 , \5951 );
or \U$6729 ( \7465 , \6749_nRb36 , \5950 );
nand \U$6730 ( \7466 , \7463 , \7464 , \7465 );
xor \U$6731 ( \7467 , \7466 , \5537 );
or \U$6732 ( \7468 , \6076 , \6990 );
or \U$6733 ( \7469 , \6749_nRb36 , \5951 );
or \U$6734 ( \7470 , \6847_nRa33 , \5950 );
nand \U$6735 ( \7471 , \7468 , \7469 , \7470 );
nand \U$6736 ( \7472 , \6847_nRa33 , \5948 );
and \U$6737 ( \7473 , \7471 , \5535 , \7472 );
xor \U$6738 ( \7474 , \7467 , \7473 );
or \U$6739 ( \7475 , \6285 , \6992 );
or \U$6740 ( \7476 , \6847_nRa33 , \5538 );
nand \U$6741 ( \7477 , \7475 , \7476 , \5879 );
and \U$6742 ( \7478 , \7474 , \7477 );
and \U$6743 ( \7479 , \7467 , \7473 );
or \U$6744 ( \7480 , \7478 , \7479 );
and \U$6745 ( \7481 , \7466 , \5537 );
xor \U$6746 ( \7482 , \7480 , \7481 );
nand \U$6747 ( \7483 , \6847_nRa33 , \5674 );
or \U$6748 ( \7484 , \5538 , \6749_nRb36 );
nand \U$6749 ( \7485 , \7484 , \5879 );
and \U$6750 ( \7486 , \7483 , \7485 );
and \U$6751 ( \7487 , \5882 , \6749_nRb36 );
and \U$6752 ( \7488 , \6847_nRa33 , \5676 );
nor \U$6753 ( \7489 , \7486 , \7487 , \7488 );
not \U$6754 ( \7490 , \6463_nRc21 );
and \U$6755 ( \7491 , \7490 , \6073 );
and \U$6756 ( \7492 , \5949 , \7462 );
and \U$6757 ( \7493 , \6463_nRc21 , \6077 );
nor \U$6758 ( \7494 , \7491 , \7492 , \7493 );
and \U$6759 ( \7495 , \7489 , \7494 );
nor \U$6760 ( \7496 , \7489 , \7494 );
nor \U$6761 ( \7497 , \7495 , \7496 );
and \U$6762 ( \7498 , \7482 , \7497 );
and \U$6763 ( \7499 , \7480 , \7481 );
or \U$6764 ( \7500 , \7498 , \7499 );
xor \U$6765 ( \7501 , \7500 , \7496 );
and \U$6766 ( \7502 , \6847_nRa33 , \5520 );
and \U$6767 ( \7503 , \6992 , \5308 );
not \U$6768 ( \7504 , \5526 );
nor \U$6769 ( \7505 , \7502 , \7503 , \7504 );
not \U$6770 ( \7506 , \6214_nRca5 );
and \U$6771 ( \7507 , \7506 , \6073 );
and \U$6772 ( \7508 , \5949 , \7490 );
and \U$6773 ( \7509 , \6214_nRca5 , \6077 );
nor \U$6774 ( \7510 , \7507 , \7508 , \7509 );
xor \U$6775 ( \7511 , \5307 , \7510 );
nand \U$6776 ( \7512 , \6749_nRb36 , \5674 );
or \U$6777 ( \7513 , \5538 , \6573_nRb98 );
nand \U$6778 ( \7514 , \7513 , \5879 );
and \U$6779 ( \7515 , \7512 , \7514 );
and \U$6780 ( \7516 , \5882 , \6573_nRb98 );
and \U$6781 ( \7517 , \6749_nRb36 , \5676 );
nor \U$6782 ( \7518 , \7515 , \7516 , \7517 );
xor \U$6783 ( \7519 , \7511 , \7518 );
and \U$6784 ( \7520 , \7505 , \7519 );
nor \U$6785 ( \7521 , \7505 , \7519 );
nor \U$6786 ( \7522 , \7520 , \7521 );
and \U$6787 ( \7523 , \7501 , \7522 );
and \U$6788 ( \7524 , \7500 , \7496 );
or \U$6789 ( \7525 , \7523 , \7524 );
xor \U$6790 ( \7526 , \7525 , \7521 );
nand \U$6791 ( \7527 , \6573_nRb98 , \5674 );
or \U$6792 ( \7528 , \5538 , \6463_nRc21 );
nand \U$6793 ( \7529 , \7528 , \5879 );
and \U$6794 ( \7530 , \7527 , \7529 );
and \U$6795 ( \7531 , \5882 , \6463_nRc21 );
and \U$6796 ( \7532 , \6573_nRb98 , \5676 );
nor \U$6797 ( \7533 , \7530 , \7531 , \7532 );
and \U$6798 ( \7534 , \7436 , \6073 );
and \U$6799 ( \7535 , \5949 , \7506 );
and \U$6800 ( \7536 , \6245_nRd47 , \6077 );
nor \U$6801 ( \7537 , \7534 , \7535 , \7536 );
xor \U$6802 ( \7538 , \7533 , \7537 );
and \U$6803 ( \7539 , \6749_nRb36 , \5520 );
or \U$6804 ( \7540 , \5307 , \6749_nRb36 );
nand \U$6805 ( \7541 , \7540 , \5526 );
nand \U$6806 ( \7542 , \6847_nRa33 , \5436 );
and \U$6807 ( \7543 , \7541 , \7542 );
and \U$6808 ( \7544 , \6847_nRa33 , \5438 );
nor \U$6809 ( \7545 , \7539 , \7543 , \7544 );
xor \U$6810 ( \7546 , \7538 , \7545 );
xor \U$6811 ( \7547 , \5307 , \7510 );
and \U$6812 ( \7548 , \7547 , \7518 );
and \U$6813 ( \7549 , \5307 , \7510 );
or \U$6814 ( \7550 , \7548 , \7549 );
and \U$6815 ( \7551 , \7546 , \7550 );
nor \U$6816 ( \7552 , \7546 , \7550 );
nor \U$6817 ( \7553 , \7551 , \7552 );
and \U$6818 ( \7554 , \7526 , \7553 );
and \U$6819 ( \7555 , \7525 , \7521 );
or \U$6820 ( \7556 , \7554 , \7555 );
xor \U$6821 ( \7557 , \7556 , \7552 );
not \U$6822 ( \7558 , \7451 );
not \U$6823 ( \7559 , \7455 );
or \U$6824 ( \7560 , \7558 , \7559 );
or \U$6825 ( \7561 , \7455 , \7451 );
nand \U$6826 ( \7562 , \7560 , \7561 );
not \U$6827 ( \7563 , \7562 );
xor \U$6828 ( \7564 , \7533 , \7537 );
and \U$6829 ( \7565 , \7564 , \7545 );
and \U$6830 ( \7566 , \7533 , \7537 );
or \U$6831 ( \7567 , \7565 , \7566 );
xor \U$6832 ( \7568 , \7434 , \7439 );
xor \U$6833 ( \7569 , \7568 , \5137 );
nand \U$6834 ( \7570 , \7567 , \7569 );
not \U$6835 ( \7571 , \7570 );
nor \U$6836 ( \7572 , \7569 , \7567 );
nor \U$6837 ( \7573 , \7571 , \7572 );
not \U$6838 ( \7574 , \7573 );
and \U$6839 ( \7575 , \7563 , \7574 );
and \U$6840 ( \7576 , \7562 , \7573 );
nor \U$6841 ( \7577 , \7575 , \7576 );
and \U$6842 ( \7578 , \7557 , \7577 );
and \U$6843 ( \7579 , \7556 , \7552 );
or \U$6844 ( \7580 , \7578 , \7579 );
and \U$6845 ( \7581 , \7562 , \7570 );
nor \U$6846 ( \7582 , \7581 , \7572 );
not \U$6847 ( \7583 , \7582 );
xor \U$6848 ( \7584 , \7580 , \7583 );
xor \U$6849 ( \7585 , \7427 , \7443 );
xor \U$6850 ( \7586 , \7585 , \7456 );
xor \U$6851 ( \7587 , \7376 , \7381 );
xor \U$6852 ( \7588 , \7587 , \7389 );
and \U$6853 ( \7589 , \7586 , \7588 );
nor \U$6854 ( \7590 , \7586 , \7588 );
nor \U$6855 ( \7591 , \7589 , \7590 );
and \U$6856 ( \7592 , \7584 , \7591 );
and \U$6857 ( \7593 , \7580 , \7583 );
or \U$6858 ( \7594 , \7592 , \7593 );
xor \U$6859 ( \7595 , \7594 , \7590 );
and \U$6860 ( \7596 , \7420 , \7459 );
nor \U$6861 ( \7597 , \7596 , \7460 );
and \U$6862 ( \7598 , \7595 , \7597 );
and \U$6863 ( \7599 , \7594 , \7590 );
or \U$6864 ( \7600 , \7598 , \7599 );
and \U$6865 ( \7601 , \7461 , \7600 );
and \U$6866 ( \7602 , \7416 , \7460 );
or \U$6867 ( \7603 , \7601 , \7602 );
and \U$6868 ( \7604 , \7409 , \7603 );
and \U$6869 ( \7605 , \7367 , \7408 );
or \U$6870 ( \7606 , \7604 , \7605 );
and \U$6871 ( \7607 , \7361 , \7366 );
xor \U$6872 ( \7608 , \7606 , \7607 );
and \U$6873 ( \7609 , \7283 , \7352 );
nor \U$6874 ( \7610 , \7609 , \7353 );
and \U$6875 ( \7611 , \7608 , \7610 );
and \U$6876 ( \7612 , \7606 , \7607 );
or \U$6877 ( \7613 , \7611 , \7612 );
and \U$6878 ( \7614 , \7354 , \7613 );
and \U$6879 ( \7615 , \7281 , \7353 );
or \U$6880 ( \7616 , \7614 , \7615 );
and \U$6881 ( \7617 , \7279 , \7616 );
and \U$6882 ( \7618 , \7230 , \7278 );
or \U$6883 ( \7619 , \7617 , \7618 );
xor \U$6884 ( \7620 , \7134 , \7136 );
xor \U$6885 ( \7621 , \7620 , \7151 );
and \U$6886 ( \7622 , \7222 , \7621 );
xor \U$6887 ( \7623 , \7134 , \7136 );
xor \U$6888 ( \7624 , \7623 , \7151 );
and \U$6889 ( \7625 , \7227 , \7624 );
and \U$6890 ( \7626 , \7222 , \7227 );
or \U$6891 ( \7627 , \7622 , \7625 , \7626 );
xor \U$6892 ( \7628 , \7075 , \7154 );
xor \U$6893 ( \7629 , \7628 , \7157 );
nand \U$6894 ( \7630 , \7627 , \7629 );
and \U$6895 ( \7631 , \7619 , \7630 );
nor \U$6896 ( \7632 , \7629 , \7627 );
nor \U$6897 ( \7633 , \7631 , \7632 );
xor \U$6898 ( \7634 , \7053 , \7055 );
xor \U$6899 ( \7635 , \7634 , \7060 );
and \U$6900 ( \7636 , \7633 , \7635 );
and \U$6901 ( \7637 , \7160 , \7633 );
or \U$6902 ( \7638 , \7163 , \7636 , \7637 );
and \U$6903 ( \7639 , \7064 , \7638 );
and \U$6904 ( \7640 , \6989 , \7063 );
or \U$6905 ( \7641 , \7639 , \7640 );
not \U$6906 ( \7642 , \7641 );
and \U$6907 ( \7643 , \6982 , \7642 );
and \U$6908 ( \7644 , \6887 , \6981 );
or \U$6909 ( \7645 , \7643 , \7644 );
and \U$6910 ( \7646 , \6885 , \7645 );
and \U$6911 ( \7647 , \6877 , \6884 );
or \U$6912 ( \7648 , \7646 , \7647 );
and \U$6913 ( \7649 , \6875 , \7648 );
and \U$6914 ( \7650 , \6712 , \6874 );
or \U$6915 ( \7651 , \7649 , \7650 );
and \U$6916 ( \7652 , \6710 , \7651 );
and \U$6917 ( \7653 , \6695 , \6709 );
or \U$6918 ( \7654 , \7652 , \7653 );
xor \U$6919 ( \7655 , \6699 , \6700 );
and \U$6920 ( \7656 , \7655 , \6708 );
and \U$6921 ( \7657 , \6699 , \6700 );
nor \U$6922 ( \7658 , \7656 , \7657 );
xor \U$6923 ( \7659 , \6419 , \6421 );
xor \U$6924 ( \7660 , \7659 , \6424 );
nand \U$6925 ( \7661 , \7658 , \7660 );
and \U$6926 ( \7662 , \7654 , \7661 );
nor \U$6927 ( \7663 , \7660 , \7658 );
nor \U$6928 ( \7664 , \7662 , \7663 );
nor \U$6929 ( \7665 , \6432 , \7664 );
nor \U$6930 ( \7666 , \6429 , \7665 );
xor \U$6931 ( \7667 , \6054 , \6137 );
xor \U$6932 ( \7668 , \7667 , \6154 );
and \U$6933 ( \7669 , \7666 , \7668 );
and \U$6934 ( \7670 , \6342 , \7666 );
or \U$6935 ( \7671 , \6345 , \7669 , \7670 );
xor \U$6936 ( \7672 , \6161 , \6166 );
xor \U$6937 ( \7673 , \7672 , \6169 );
and \U$6938 ( \7674 , \7671 , \7673 );
and \U$6939 ( \7675 , \6157 , \7671 );
or \U$6940 ( \7676 , \6171 , \7674 , \7675 );
not \U$6941 ( \7677 , \7676 );
xor \U$6942 ( \7678 , \5779 , \5786 );
xor \U$6943 ( \7679 , \7678 , \5908 );
xor \U$6944 ( \7680 , \6161 , \6166 );
and \U$6945 ( \7681 , \7680 , \6169 );
and \U$6946 ( \7682 , \6161 , \6166 );
or \U$6947 ( \7683 , \7681 , \7682 );
and \U$6948 ( \7684 , \7679 , \7683 );
not \U$6949 ( \7685 , \7684 );
and \U$6950 ( \7686 , \7677 , \7685 );
nor \U$6951 ( \7687 , \7679 , \7683 );
nor \U$6952 ( \7688 , \7686 , \7687 );
and \U$6953 ( \7689 , \5912 , \7688 );
and \U$6954 ( \7690 , \5773 , \5911 );
or \U$6955 ( \7691 , \7689 , \7690 );
not \U$6956 ( \7692 , \7691 );
and \U$6957 ( \7693 , \5767 , \7692 );
and \U$6958 ( \7694 , \5764 , \5766 );
or \U$6959 ( \7695 , \7693 , \7694 );
and \U$6960 ( \7696 , \5643 , \7695 );
and \U$6961 ( \7697 , \5616 , \5642 );
or \U$6962 ( \7698 , \7696 , \7697 );
or \U$6963 ( \7699 , \5630 , \5638 );
nand \U$6964 ( \7700 , \7699 , \5628 );
xor \U$6965 ( \7701 , \5387 , \5389 );
xor \U$6966 ( \7702 , \7701 , \5397 );
nand \U$6967 ( \7703 , \7700 , \7702 );
and \U$6968 ( \7704 , \7698 , \7703 );
nor \U$6969 ( \7705 , \7702 , \7700 );
nor \U$6970 ( \7706 , \7704 , \7705 );
and \U$6971 ( \7707 , \5401 , \7706 );
and \U$6972 ( \7708 , \5282 , \5400 );
or \U$6973 ( \7709 , \7707 , \7708 );
and \U$6974 ( \7710 , \5280 , \7709 );
and \U$6975 ( \7711 , \5108 , \5279 );
or \U$6976 ( \7712 , \7710 , \7711 );
nor \U$6977 ( \7713 , \5102 , \7712 );
nor \U$6978 ( \7714 , \5099 , \7713 );
not \U$6979 ( \7715 , \7714 );
or \U$6980 ( \7716 , \4994 , \7715 );
or \U$6981 ( \7717 , \7714 , \4993 );
nand \U$6982 ( \7718 , \7716 , \7717 );
buf \U$6983 ( \7719 , \4414 );
buf \U$6984 ( \7720 , \766 );
_DC r53c ( \7721_nR53c , \7719 , \7720 );
not \U$6985 ( \7722 , \7721_nR53c );
buf \U$6986 ( \7723 , \4444 );
_DC r55b ( \7724_nR55b , \7723 , \7720 );
not \U$6987 ( \7725 , \7724_nR55b );
buf \U$6988 ( \7726 , \1157 );
buf \U$6989 ( \7727 , \766 );
_DC r613 ( \7728_nR613 , \7726 , \7727 );
not \U$6990 ( \7729 , \7728_nR613 );
not \U$6991 ( \7730 , \7729 );
buf \U$6992 ( \7731 , \4624 );
_DC r615 ( \7732_nR615 , \7731 , \7720 );
not \U$6993 ( \7733 , \7732_nR615 );
and \U$6994 ( \7734 , \7730 , \7733 );
buf \U$6995 ( \7735 , \1188 );
_DC r632 ( \7736_nR632 , \7735 , \7727 );
nor \U$6996 ( \7737 , \7734 , \7736_nR632 );
buf \U$6997 ( \7738 , \4654 );
_DC r634 ( \7739_nR634 , \7738 , \7720 );
and \U$6998 ( \7740 , \7737 , \7739_nR634 );
and \U$6999 ( \7741 , \7732_nR615 , \7729 );
nor \U$7000 ( \7742 , \7740 , \7741 );
buf \U$7001 ( \7743 , \4594 );
_DC r5f6 ( \7744_nR5f6 , \7743 , \7720 );
not \U$7002 ( \7745 , \7744_nR5f6 );
and \U$7003 ( \7746 , \7742 , \7745 );
buf \U$7004 ( \7747 , \1126 );
_DC r5f4 ( \7748_nR5f4 , \7747 , \7727 );
or \U$7005 ( \7749 , \7746 , \7748_nR5f4 );
or \U$7006 ( \7750 , \7745 , \7742 );
nand \U$7007 ( \7751 , \7749 , \7750 );
buf \U$7008 ( \7752 , \4564 );
_DC r5d7 ( \7753_nR5d7 , \7752 , \7720 );
and \U$7009 ( \7754 , \7751 , \7753_nR5d7 );
not \U$7010 ( \7755 , \7751 );
not \U$7011 ( \7756 , \7753_nR5d7 );
and \U$7012 ( \7757 , \7755 , \7756 );
buf \U$7013 ( \7758 , \1090 );
_DC r5d5 ( \7759_nR5d5 , \7758 , \7727 );
nor \U$7014 ( \7760 , \7757 , \7759_nR5d5 );
nor \U$7015 ( \7761 , \7754 , \7760 );
buf \U$7016 ( \7762 , \4534 );
_DC r5b8 ( \7763_nR5b8 , \7762 , \7720 );
not \U$7017 ( \7764 , \7763_nR5b8 );
buf \U$7018 ( \7765 , \1054 );
_DC r5b6 ( \7766_nR5b6 , \7765 , \7727 );
and \U$7019 ( \7767 , \7764 , \7766_nR5b6 );
or \U$7020 ( \7768 , \7761 , \7767 );
or \U$7021 ( \7769 , \7766_nR5b6 , \7764 );
nand \U$7022 ( \7770 , \7768 , \7769 );
buf \U$7023 ( \7771 , \4504 );
_DC r599 ( \7772_nR599 , \7771 , \7720 );
and \U$7024 ( \7773 , \7770 , \7772_nR599 );
not \U$7025 ( \7774 , \7770 );
not \U$7026 ( \7775 , \7772_nR599 );
and \U$7027 ( \7776 , \7774 , \7775 );
buf \U$7028 ( \7777 , \1018 );
_DC r597 ( \7778_nR597 , \7777 , \7727 );
nor \U$7029 ( \7779 , \7776 , \7778_nR597 );
nor \U$7030 ( \7780 , \7773 , \7779 );
buf \U$7031 ( \7781 , \4474 );
_DC r57a ( \7782_nR57a , \7781 , \7720 );
not \U$7032 ( \7783 , \7782_nR57a );
buf \U$7033 ( \7784 , \982 );
_DC r578 ( \7785_nR578 , \7784 , \7727 );
and \U$7034 ( \7786 , \7783 , \7785_nR578 );
or \U$7035 ( \7787 , \7780 , \7786 );
or \U$7036 ( \7788 , \7785_nR578 , \7783 );
nand \U$7037 ( \7789 , \7787 , \7788 );
not \U$7038 ( \7790 , \7789 );
or \U$7039 ( \7791 , \7725 , \7790 );
nor \U$7040 ( \7792 , \7789 , \7724_nR55b );
buf \U$7041 ( \7793 , \946 );
_DC r559 ( \7794_nR559 , \7793 , \7727 );
or \U$7042 ( \7795 , \7792 , \7794_nR559 );
nand \U$7043 ( \7796 , \7791 , \7795 );
not \U$7044 ( \7797 , \7796 );
or \U$7045 ( \7798 , \7722 , \7797 );
nor \U$7046 ( \7799 , \7796 , \7721_nR53c );
buf \U$7047 ( \7800 , \910 );
_DC r53a ( \7801_nR53a , \7800 , \7727 );
or \U$7048 ( \7802 , \7799 , \7801_nR53a );
nand \U$7049 ( \7803 , \7798 , \7802 );
buf \U$7050 ( \7804 , \4384 );
_DC r51d ( \7805_nR51d , \7804 , \7720 );
and \U$7051 ( \7806 , \7803 , \7805_nR51d );
not \U$7052 ( \7807 , \7803 );
not \U$7053 ( \7808 , \7805_nR51d );
and \U$7054 ( \7809 , \7807 , \7808 );
buf \U$7055 ( \7810 , \874 );
_DC r51b ( \7811_nR51b , \7810 , \7727 );
nor \U$7056 ( \7812 , \7809 , \7811_nR51b );
nor \U$7057 ( \7813 , \7806 , \7812 );
buf \U$7058 ( \7814 , \4354 );
_DC r4fe ( \7815_nR4fe , \7814 , \7720 );
not \U$7059 ( \7816 , \7815_nR4fe );
buf \U$7060 ( \7817 , \838 );
_DC r4fc ( \7818_nR4fc , \7817 , \7727 );
and \U$7061 ( \7819 , \7816 , \7818_nR4fc );
or \U$7062 ( \7820 , \7813 , \7819 );
or \U$7063 ( \7821 , \7818_nR4fc , \7816 );
nand \U$7064 ( \7822 , \7820 , \7821 );
buf \U$7065 ( \7823 , \4324 );
_DC r4df ( \7824_nR4df , \7823 , \7720 );
and \U$7066 ( \7825 , \7822 , \7824_nR4df );
not \U$7067 ( \7826 , \7822 );
not \U$7068 ( \7827 , \7824_nR4df );
and \U$7069 ( \7828 , \7826 , \7827 );
buf \U$7070 ( \7829 , \802 );
_DC r4c2 ( \7830_nR4c2 , \7829 , \7727 );
nor \U$7071 ( \7831 , \7828 , \7830_nR4c2 );
nor \U$7072 ( \7832 , \7825 , \7831 );
buf \U$7073 ( \7833 , \4293 );
_DC r4a4 ( \7834_nR4a4 , \7833 , \7720 );
not \U$7074 ( \7835 , \7834_nR4a4 );
buf \U$7075 ( \7836 , \764 );
_DC r486 ( \7837_nR486 , \7836 , \7727 );
and \U$7076 ( \7838 , \7835 , \7837_nR486 );
or \U$7077 ( \7839 , \7832 , \7838 );
or \U$7078 ( \7840 , \7837_nR486 , \7835 );
nand \U$7079 ( \7841 , \7839 , \7840 );
nor \U$7080 ( \7842 , \671 , RIb55b778_588);
nand \U$7081 ( \7843 , RIb54a810_9, \7842 );
not \U$7082 ( \7844 , \7843 );
nand \U$7083 ( \7845 , RIb54a798_8, \7844 );
not \U$7084 ( \7846 , \7845 );
nand \U$7085 ( \7847 , RIb54a720_7, \7846 );
not \U$7086 ( \7848 , \7847 );
nand \U$7087 ( \7849 , RIb54a6a8_6, \7848 );
not \U$7088 ( \7850 , \7849 );
and \U$7089 ( \7851 , \7850 , RIb54a630_5);
nand \U$7090 ( \7852 , RIb54a5b8_4, \7851 );
not \U$7091 ( \7853 , \7852 );
and \U$7092 ( \7854 , \7853 , RIb54a540_3);
nand \U$7093 ( \7855 , RIb54a4c8_2, \7854 );
not \U$7094 ( \7856 , \7855 );
nand \U$7095 ( \7857 , RIb54a450_1, \7856 );
not \U$7096 ( \7858 , \7857 );
not \U$7097 ( \7859 , RIb5517a0_247);
and \U$7098 ( \7860 , \7858 , \7859 );
and \U$7099 ( \7861 , \7857 , RIb5517a0_247);
nor \U$7100 ( \7862 , \7860 , \7861 );
buf \U$7101 ( \7863 , \4293 );
buf \U$7102 ( \7864 , \766 );
_DC raa0 ( \7865_nRaa0 , \7863 , \7864 );
or \U$7103 ( \7866 , \7862 , \7865_nRaa0 );
buf \U$7104 ( \7867 , \4324 );
_DC raa3 ( \7868_nRaa3 , \7867 , \7864 );
or \U$7105 ( \7869 , \7856 , RIb54a450_1);
nand \U$7106 ( \7870 , \7869 , \7857 );
or \U$7107 ( \7871 , \7868_nRaa3 , \7870 );
not \U$7108 ( \7872 , \7868_nRaa3 );
not \U$7109 ( \7873 , \7870 );
or \U$7110 ( \7874 , \7872 , \7873 );
or \U$7111 ( \7875 , \7851 , RIb54a5b8_4);
nand \U$7112 ( \7876 , \7875 , \7852 );
buf \U$7113 ( \7877 , \4414 );
_DC r35b ( \7878_nR35b , \7877 , \7864 );
and \U$7114 ( \7879 , \7876 , \7878_nR35b );
not \U$7115 ( \7880 , \7876 );
not \U$7116 ( \7881 , \7878_nR35b );
and \U$7117 ( \7882 , \7880 , \7881 );
nor \U$7118 ( \7883 , \7850 , RIb54a630_5);
buf \U$7119 ( \7884 , \4444 );
_DC r379 ( \7885_nR379 , \7884 , \7864 );
or \U$7120 ( \7886 , \7851 , \7883 , \7885_nR379 );
buf \U$7121 ( \7887 , \4474 );
_DC r397 ( \7888_nR397 , \7887 , \7864 );
not \U$7122 ( \7889 , \7888_nR397 );
or \U$7123 ( \7890 , \7848 , RIb54a6a8_6);
nand \U$7124 ( \7891 , \7890 , \7849 );
not \U$7125 ( \7892 , \7891 );
or \U$7126 ( \7893 , \7889 , \7892 );
or \U$7127 ( \7894 , \7891 , \7888_nR397 );
buf \U$7128 ( \7895 , \4504 );
_DC r3b5 ( \7896_nR3b5 , \7895 , \7864 );
not \U$7129 ( \7897 , \7896_nR3b5 );
buf \U$7130 ( \7898 , \4534 );
_DC r3d3 ( \7899_nR3d3 , \7898 , \7864 );
not \U$7131 ( \7900 , \7899_nR3d3 );
or \U$7132 ( \7901 , \7844 , RIb54a798_8);
nand \U$7133 ( \7902 , \7901 , \7845 );
not \U$7134 ( \7903 , \7902 );
or \U$7135 ( \7904 , \7900 , \7903 );
or \U$7136 ( \7905 , \7902 , \7899_nR3d3 );
buf \U$7137 ( \7906 , \4564 );
_DC r3f1 ( \7907_nR3f1 , \7906 , \7864 );
not \U$7138 ( \7908 , \7907_nR3f1 );
buf \U$7139 ( \7909 , \4594 );
_DC r40f ( \7910_nR40f , \7909 , \7864 );
not \U$7140 ( \7911 , \7910_nR40f );
nor \U$7141 ( \7912 , \1094 , RIb55b778_588);
not \U$7142 ( \7913 , RIb55b778_588);
nor \U$7143 ( \7914 , \7913 , RIb54a900_11);
buf \U$7144 ( \7915 , \4624 );
_DC r42d ( \7916_nR42d , \7915 , \7864 );
or \U$7145 ( \7917 , \7912 , \7914 , \7916_nR42d );
buf \U$7146 ( \7918 , \4654 );
_DC r44b ( \7919_nR44b , \7918 , \7864 );
nand \U$7147 ( \7920 , \7917 , \7919_nR44b );
or \U$7148 ( \7921 , \7920 , RIb550378_204);
or \U$7149 ( \7922 , \7912 , \7914 );
nand \U$7150 ( \7923 , \7922 , \7916_nR42d );
nand \U$7151 ( \7924 , \7921 , \7923 );
not \U$7152 ( \7925 , \7924 );
or \U$7153 ( \7926 , \7911 , \7925 );
or \U$7154 ( \7927 , \7924 , \7910_nR40f );
not \U$7155 ( \7928 , RIb54a888_10);
not \U$7156 ( \7929 , \7912 );
or \U$7157 ( \7930 , \7928 , \7929 );
or \U$7158 ( \7931 , \7912 , RIb54a888_10);
nand \U$7159 ( \7932 , \7930 , \7931 );
nand \U$7160 ( \7933 , \7927 , \7932 );
nand \U$7161 ( \7934 , \7926 , \7933 );
not \U$7162 ( \7935 , \7934 );
or \U$7163 ( \7936 , \7908 , \7935 );
or \U$7164 ( \7937 , \7934 , \7907_nR3f1 );
or \U$7165 ( \7938 , \7842 , RIb54a810_9);
nand \U$7166 ( \7939 , \7938 , \7843 );
nand \U$7167 ( \7940 , \7937 , \7939 );
nand \U$7168 ( \7941 , \7936 , \7940 );
nand \U$7169 ( \7942 , \7905 , \7941 );
nand \U$7170 ( \7943 , \7904 , \7942 );
not \U$7171 ( \7944 , \7943 );
or \U$7172 ( \7945 , \7897 , \7944 );
or \U$7173 ( \7946 , \7943 , \7896_nR3b5 );
or \U$7174 ( \7947 , \7846 , RIb54a720_7);
nand \U$7175 ( \7948 , \7947 , \7847 );
nand \U$7176 ( \7949 , \7946 , \7948 );
nand \U$7177 ( \7950 , \7945 , \7949 );
nand \U$7178 ( \7951 , \7894 , \7950 );
nand \U$7179 ( \7952 , \7893 , \7951 );
nand \U$7180 ( \7953 , \7886 , \7952 );
or \U$7181 ( \7954 , \7851 , \7883 );
nand \U$7182 ( \7955 , \7954 , \7885_nR379 );
and \U$7183 ( \7956 , \7953 , \7955 );
nor \U$7184 ( \7957 , \7882 , \7956 );
nor \U$7185 ( \7958 , \7879 , \7957 );
nor \U$7186 ( \7959 , \7853 , RIb54a540_3);
buf \U$7187 ( \7960 , \4384 );
_DC r33d ( \7961_nR33d , \7960 , \7864 );
nor \U$7188 ( \7962 , \7854 , \7959 , \7961_nR33d );
or \U$7189 ( \7963 , \7958 , \7962 );
or \U$7190 ( \7964 , \7854 , \7959 );
nand \U$7191 ( \7965 , \7964 , \7961_nR33d );
nand \U$7192 ( \7966 , \7963 , \7965 );
or \U$7193 ( \7967 , \7854 , RIb54a4c8_2);
nand \U$7194 ( \7968 , \7967 , \7855 );
buf \U$7195 ( \7969 , \4354 );
_DC r31f ( \7970_nR31f , \7969 , \7864 );
or \U$7196 ( \7971 , \7968 , \7970_nR31f );
and \U$7197 ( \7972 , \7966 , \7971 );
and \U$7198 ( \7973 , \7970_nR31f , \7968 );
nor \U$7199 ( \7974 , \7972 , \7973 );
nand \U$7200 ( \7975 , \7874 , \7974 );
nand \U$7201 ( \7976 , \7866 , \7871 , \7975 );
nand \U$7202 ( \7977 , \7865_nRaa0 , \7862 );
and \U$7203 ( \7978 , \7841 , \7976 , \1238 , \7977 );
_HMUX r23b8 ( \7979_nR23b8 , \4252 , \7718 , \7978 );
buf \U$7204 ( \7980 , \7979_nR23b8 );
xor \U$7205 ( \7981 , \1653 , \1654 );
xor \U$7206 ( \7982 , \7981 , \4245 );
xor \U$7207 ( \7983 , \5098 , \5097 );
not \U$7208 ( \7984 , \7983 );
not \U$7209 ( \7985 , \7712 );
or \U$7210 ( \7986 , \7984 , \7985 );
or \U$7211 ( \7987 , \7712 , \7983 );
nand \U$7212 ( \7988 , \7986 , \7987 );
_HMUX r237b ( \7989_nR237b , \7982 , \7988 , \7978 );
buf \U$7213 ( \7990 , \7989_nR237b );
xor \U$7214 ( \7991 , \1657 , \1837 );
xor \U$7215 ( \7992 , \7991 , \4242 );
xor \U$7216 ( \7993 , \5108 , \5279 );
xor \U$7217 ( \7994 , \7993 , \7709 );
not \U$7218 ( \7995 , \7994 );
_HMUX r2348 ( \7996_nR2348 , \7992 , \7995 , \7978 );
buf \U$7219 ( \7997 , \7996_nR2348 );
xor \U$7220 ( \7998 , \1840 , \1960 );
xor \U$7221 ( \7999 , \7998 , \4239 );
xor \U$7222 ( \8000 , \5282 , \5400 );
xor \U$7223 ( \8001 , \8000 , \7706 );
not \U$7224 ( \8002 , \8001 );
_HMUX r2309 ( \8003_nR2309 , \7999 , \8002 , \7978 );
buf \U$7225 ( \8004 , \8003_nR2309 );
xor \U$7226 ( \8005 , \1963 , \2069 );
xor \U$7227 ( \8006 , \8005 , \4236 );
not \U$7228 ( \8007 , \7705 );
nand \U$7229 ( \8008 , \8007 , \7703 );
not \U$7230 ( \8009 , \8008 );
not \U$7231 ( \8010 , \7698 );
or \U$7232 ( \8011 , \8009 , \8010 );
or \U$7233 ( \8012 , \7698 , \8008 );
nand \U$7234 ( \8013 , \8011 , \8012 );
_HMUX r22a9 ( \8014_nR22a9 , \8006 , \8013 , \7978 );
buf \U$7235 ( \8015 , \8014_nR22a9 );
xor \U$7236 ( \8016 , \2183 , \2185 );
xor \U$7237 ( \8017 , \8016 , \4233 );
xor \U$7238 ( \8018 , \5616 , \5642 );
xor \U$7239 ( \8019 , \8018 , \7695 );
_HMUX r2238 ( \8020_nR2238 , \8017 , \8019 , \7978 );
buf \U$7240 ( \8021 , \8020_nR2238 );
xor \U$7241 ( \8022 , \2190 , \2310 );
xor \U$7242 ( \8023 , \8022 , \4230 );
xor \U$7243 ( \8024 , \5764 , \5766 );
xor \U$7244 ( \8025 , \8024 , \7692 );
_HMUX r21a2 ( \8026_nR21a2 , \8023 , \8025 , \7978 );
buf \U$7245 ( \8027 , \8026_nR21a2 );
xor \U$7246 ( \8028 , \2447 , \2313 );
not \U$7247 ( \8029 , \8028 );
not \U$7248 ( \8030 , \4227 );
or \U$7249 ( \8031 , \8029 , \8030 );
or \U$7250 ( \8032 , \4227 , \8028 );
nand \U$7251 ( \8033 , \8031 , \8032 );
xor \U$7252 ( \8034 , \5773 , \5911 );
xor \U$7253 ( \8035 , \8034 , \7688 );
not \U$7254 ( \8036 , \8035 );
_HMUX r20fe ( \8037_nR20fe , \8033 , \8036 , \7978 );
buf \U$7255 ( \8038 , \8037_nR20fe );
not \U$7256 ( \8039 , \4226 );
nand \U$7257 ( \8040 , \8039 , \4224 );
not \U$7258 ( \8041 , \8040 );
not \U$7259 ( \8042 , \4213 );
or \U$7260 ( \8043 , \8041 , \8042 );
or \U$7261 ( \8044 , \4213 , \8040 );
nand \U$7262 ( \8045 , \8043 , \8044 );
nor \U$7263 ( \8046 , \7687 , \7684 );
not \U$7264 ( \8047 , \8046 );
not \U$7265 ( \8048 , \7676 );
or \U$7266 ( \8049 , \8047 , \8048 );
or \U$7267 ( \8050 , \7676 , \8046 );
nand \U$7268 ( \8051 , \8049 , \8050 );
_HMUX r2046 ( \8052_nR2046 , \8045 , \8051 , \7978 );
buf \U$7269 ( \8053 , \8052_nR2046 );
xor \U$7270 ( \8054 , \2623 , \2724 );
xor \U$7271 ( \8055 , \8054 , \4210 );
xor \U$7272 ( \8056 , \6161 , \6166 );
xor \U$7273 ( \8057 , \8056 , \6169 );
xor \U$7274 ( \8058 , \6157 , \7671 );
xor \U$7275 ( \8059 , \8057 , \8058 );
not \U$7276 ( \8060 , \8059 );
_HMUX r1f79 ( \8061_nR1f79 , \8055 , \8060 , \7978 );
buf \U$7277 ( \8062 , \8061_nR1f79 );
xor \U$7278 ( \8063 , \2894 , \2896 );
xor \U$7279 ( \8064 , \8063 , \4206 );
not \U$7280 ( \8065 , \8064 );
xor \U$7281 ( \8066 , \6054 , \6137 );
xor \U$7282 ( \8067 , \8066 , \6154 );
xor \U$7283 ( \8068 , \6342 , \7666 );
xor \U$7284 ( \8069 , \8067 , \8068 );
not \U$7285 ( \8070 , \8069 );
_HMUX r1eb0 ( \8071_nR1eb0 , \8065 , \8070 , \7978 );
buf \U$7286 ( \8072 , \8071_nR1eb0 );
xor \U$7287 ( \8073 , \2730 , \2731 );
xor \U$7288 ( \8074 , \8073 , \2891 );
xor \U$7289 ( \8075 , \2969 , \4201 );
xor \U$7290 ( \8076 , \8074 , \8075 );
not \U$7291 ( \8077 , \8076 );
not \U$7292 ( \8078 , \6427 );
not \U$7293 ( \8079 , \6351 );
or \U$7294 ( \8080 , \8078 , \8079 );
or \U$7295 ( \8081 , \6351 , \6427 );
nand \U$7296 ( \8082 , \8080 , \8081 );
not \U$7297 ( \8083 , \8082 );
not \U$7298 ( \8084 , \7664 );
or \U$7299 ( \8085 , \8083 , \8084 );
or \U$7300 ( \8086 , \7664 , \8082 );
nand \U$7301 ( \8087 , \8085 , \8086 );
_HMUX r1dda ( \8088_nR1dda , \8077 , \8087 , \7978 );
buf \U$7302 ( \8089 , \8088_nR1dda );
xor \U$7303 ( \8090 , \2961 , \2963 );
xor \U$7304 ( \8091 , \8090 , \2966 );
xor \U$7305 ( \8092 , \3167 , \4196 );
xor \U$7306 ( \8093 , \8091 , \8092 );
not \U$7307 ( \8094 , \8093 );
not \U$7308 ( \8095 , \7663 );
nand \U$7309 ( \8096 , \8095 , \7661 );
not \U$7310 ( \8097 , \8096 );
not \U$7311 ( \8098 , \7654 );
or \U$7312 ( \8099 , \8097 , \8098 );
or \U$7313 ( \8100 , \7654 , \8096 );
nand \U$7314 ( \8101 , \8099 , \8100 );
_HMUX r1cfd ( \8102_nR1cfd , \8094 , \8101 , \7978 );
buf \U$7315 ( \8103 , \8102_nR1cfd );
not \U$7316 ( \8104 , \4195 );
nand \U$7317 ( \8105 , \8104 , \4193 );
not \U$7318 ( \8106 , \8105 );
not \U$7319 ( \8107 , \4186 );
or \U$7320 ( \8108 , \8106 , \8107 );
or \U$7321 ( \8109 , \4186 , \8105 );
nand \U$7322 ( \8110 , \8108 , \8109 );
xor \U$7323 ( \8111 , \6695 , \6709 );
xor \U$7324 ( \8112 , \8111 , \7651 );
_HMUX r1c44 ( \8113_nR1c44 , \8110 , \8112 , \7978 );
buf \U$7325 ( \8114 , \8113_nR1c44 );
xor \U$7326 ( \8115 , \3268 , \3432 );
xor \U$7327 ( \8116 , \8115 , \4183 );
xor \U$7328 ( \8117 , \6712 , \6874 );
xor \U$7329 ( \8118 , \8117 , \7648 );
_HMUX r1b4c ( \8119_nR1b4c , \8116 , \8118 , \7978 );
buf \U$7330 ( \8120 , \8119_nR1b4c );
xor \U$7331 ( \8121 , \3435 , \3442 );
xor \U$7332 ( \8122 , \8121 , \4180 );
xor \U$7333 ( \8123 , \6877 , \6884 );
xor \U$7334 ( \8124 , \8123 , \7645 );
_HMUX r1a31 ( \8125_nR1a31 , \8122 , \8124 , \7978 );
buf \U$7335 ( \8126 , \8125_nR1a31 );
xor \U$7336 ( \8127 , \3445 , \3534 );
xor \U$7337 ( \8128 , \8127 , \4177 );
xor \U$7338 ( \8129 , \6887 , \6981 );
xor \U$7339 ( \8130 , \8129 , \7642 );
_HMUX r1915 ( \8131_nR1915 , \8128 , \8130 , \7978 );
buf \U$7340 ( \8132 , \8131_nR1915 );
xor \U$7341 ( \8133 , \3447 , \3452 );
xor \U$7342 ( \8134 , \8133 , \3530 );
xor \U$7343 ( \8135 , \3606 , \4171 );
xor \U$7344 ( \8136 , \8134 , \8135 );
not \U$7345 ( \8137 , \8136 );
xor \U$7346 ( \8138 , \6989 , \7063 );
xor \U$7347 ( \8139 , \8138 , \7638 );
not \U$7348 ( \8140 , \8139 );
_HMUX r181e ( \8141_nR181e , \8137 , \8140 , \7978 );
buf \U$7349 ( \8142 , \8141_nR181e );
xor \U$7350 ( \8143 , \3598 , \3600 );
xor \U$7351 ( \8144 , \8143 , \3603 );
xor \U$7352 ( \8145 , \3698 , \4166 );
xor \U$7353 ( \8146 , \8144 , \8145 );
not \U$7354 ( \8147 , \8146 );
xor \U$7355 ( \8148 , \7053 , \7055 );
xor \U$7356 ( \8149 , \8148 , \7060 );
xor \U$7357 ( \8150 , \7160 , \7633 );
xor \U$7358 ( \8151 , \8149 , \8150 );
not \U$7359 ( \8152 , \8151 );
_HMUX r16e0 ( \8153_nR16e0 , \8147 , \8152 , \7978 );
buf \U$7360 ( \8154 , \8153_nR16e0 );
not \U$7361 ( \8155 , \4165 );
nand \U$7362 ( \8156 , \8155 , \4163 );
not \U$7363 ( \8157 , \8156 );
not \U$7364 ( \8158 , \4152 );
or \U$7365 ( \8159 , \8157 , \8158 );
or \U$7366 ( \8160 , \4152 , \8156 );
nand \U$7367 ( \8161 , \8159 , \8160 );
not \U$7368 ( \8162 , \7632 );
nand \U$7369 ( \8163 , \8162 , \7630 );
not \U$7370 ( \8164 , \8163 );
not \U$7371 ( \8165 , \7619 );
or \U$7372 ( \8166 , \8164 , \8165 );
or \U$7373 ( \8167 , \7619 , \8163 );
nand \U$7374 ( \8168 , \8166 , \8167 );
_HMUX r15f3 ( \8169_nR15f3 , \8161 , \8168 , \7978 );
buf \U$7375 ( \8170 , \8169_nR15f3 );
xor \U$7376 ( \8171 , \3764 , \3808 );
xor \U$7377 ( \8172 , \8171 , \4149 );
xor \U$7378 ( \8173 , \7230 , \7278 );
xor \U$7379 ( \8174 , \8173 , \7616 );
_HMUX r14d3 ( \8175_nR14d3 , \8172 , \8174 , \7978 );
buf \U$7380 ( \8176 , \8175_nR14d3 );
xor \U$7381 ( \8177 , \3811 , \3882 );
xor \U$7382 ( \8178 , \8177 , \4146 );
xor \U$7383 ( \8179 , \7281 , \7353 );
xor \U$7384 ( \8180 , \8179 , \7613 );
_HMUX r13d0 ( \8181_nR13d0 , \8178 , \8180 , \7978 );
buf \U$7385 ( \8182 , \8181_nR13d0 );
xor \U$7386 ( \8183 , \4139 , \4140 );
xor \U$7387 ( \8184 , \8183 , \4143 );
xor \U$7388 ( \8185 , \7606 , \7607 );
xor \U$7389 ( \8186 , \8185 , \7610 );
_HMUX r12be ( \8187_nR12be , \8184 , \8186 , \7978 );
buf \U$7390 ( \8188 , \8187_nR12be );
xor \U$7391 ( \8189 , \3894 , \3941 );
xor \U$7392 ( \8190 , \8189 , \4136 );
xor \U$7393 ( \8191 , \7367 , \7408 );
xor \U$7394 ( \8192 , \8191 , \7603 );
_HMUX r11e2 ( \8193_nR11e2 , \8190 , \8192 , \7978 );
buf \U$7395 ( \8194 , \8193_nR11e2 );
xor \U$7396 ( \8195 , \3948 , \3992 );
xor \U$7397 ( \8196 , \8195 , \4133 );
xor \U$7398 ( \8197 , \7416 , \7460 );
xor \U$7399 ( \8198 , \8197 , \7600 );
_HMUX r10d7 ( \8199_nR10d7 , \8196 , \8198 , \7978 );
buf \U$7400 ( \8200 , \8199_nR10d7 );
xor \U$7401 ( \8201 , \4127 , \4123 );
xor \U$7402 ( \8202 , \8201 , \4130 );
xor \U$7403 ( \8203 , \7594 , \7590 );
xor \U$7404 ( \8204 , \8203 , \7597 );
_HMUX rffc ( \8205_nRffc , \8202 , \8204 , \7978 );
buf \U$7405 ( \8206 , \8205_nRffc );
xor \U$7406 ( \8207 , \4113 , \4116 );
xor \U$7407 ( \8208 , \8207 , \4124 );
xor \U$7408 ( \8209 , \7580 , \7583 );
xor \U$7409 ( \8210 , \8209 , \7591 );
_HMUX rf1c ( \8211_nRf1c , \8208 , \8210 , \7978 );
buf \U$7410 ( \8212 , \8211_nRf1c );
nand \U$7411 ( \8213 , RIb55bca0_599, RIb55bc28_598);
not \U$7412 ( \8214 , \8213 );
nand \U$7413 ( \8215 , \8214 , RIb55bbb0_597);
not \U$7414 ( \8216 , \8215 );
nand \U$7415 ( \8217 , \8216 , RIb55bb38_596);
not \U$7416 ( \8218 , \8217 );
nand \U$7417 ( \8219 , \8218 , RIb55bac0_595);
not \U$7418 ( \8220 , \8219 );
nand \U$7419 ( \8221 , \8220 , RIb55ba48_594);
not \U$7420 ( \8222 , \8221 );
nand \U$7421 ( \8223 , \8222 , RIb55b9d0_593);
not \U$7422 ( \8224 , \8223 );
nand \U$7423 ( \8225 , \8224 , RIb55b958_592);
not \U$7424 ( \8226 , \8225 );
nand \U$7425 ( \8227 , \8226 , RIb55b8e0_591);
not \U$7426 ( \8228 , \8227 );
nand \U$7427 ( \8229 , \8228 , RIb55b868_590);
not \U$7428 ( \8230 , \8229 );
nand \U$7429 ( \8231 , \8230 , RIb55b7f0_589);
not \U$7430 ( \8232 , \8231 );
not \U$7431 ( \8233 , RIb55c3a8_614);
and \U$7432 ( \8234 , \8232 , \8233 );
and \U$7433 ( \8235 , \8231 , RIb55c3a8_614);
nor \U$7434 ( \8236 , \8234 , \8235 );
not \U$7435 ( \8237 , RIb55bef8_604);
nand \U$7436 ( \8238 , RIb55be80_603, \8237 );
not \U$7437 ( \8239 , \8238 );
nand \U$7438 ( \8240 , \8239 , RIb55be08_602);
not \U$7439 ( \8241 , RIb55bd18_600);
nand \U$7440 ( \8242 , RIb55bd90_601, \8241 );
nor \U$7441 ( \8243 , \8240 , \8242 );
and \U$7442 ( \8244 , RIb551908_250, \8243 );
nand \U$7443 ( \8245 , RIb55bd90_601, RIb55bd18_600);
not \U$7444 ( \8246 , RIb55be08_602);
nor \U$7445 ( \8247 , \8245 , \8246 );
not \U$7446 ( \8248 , \8247 );
nor \U$7447 ( \8249 , \8248 , \8238 );
and \U$7448 ( \8250 , RIb551890_249, \8249 );
not \U$7449 ( \8251 , RIb55be80_603);
nand \U$7450 ( \8252 , \8251 , \8237 );
not \U$7451 ( \8253 , \8252 );
nand \U$7452 ( \8254 , RIb55be08_602, \8253 );
nor \U$7453 ( \8255 , \8254 , \8242 );
and \U$7454 ( \8256 , RIb551cc8_258, \8255 );
and \U$7455 ( \8257 , \8247 , \8253 );
and \U$7456 ( \8258 , RIb551c50_257, \8257 );
not \U$7457 ( \8259 , RIb55bd90_601);
nand \U$7458 ( \8260 , \8259 , RIb55bd18_600);
nor \U$7459 ( \8261 , \8260 , \8252 , RIb55be08_602);
and \U$7460 ( \8262 , \8261 , RIb551f20_263);
nor \U$7461 ( \8263 , \8242 , \8238 , RIb55be08_602);
and \U$7462 ( \8264 , RIb551ae8_254, \8263 );
nor \U$7463 ( \8265 , \8262 , \8264 );
not \U$7464 ( \8266 , \8265 );
nor \U$7465 ( \8267 , \8256 , \8258 , \8266 );
nor \U$7466 ( \8268 , RIb55bd18_600, RIb55bd90_601);
and \U$7467 ( \8269 , \8268 , \8246 );
and \U$7468 ( \8270 , \8269 , \8253 );
and \U$7469 ( \8271 , \8270 , RIb551f98_264);
nor \U$7470 ( \8272 , \8242 , \8252 , RIb55be08_602);
and \U$7471 ( \8273 , RIb551ea8_262, \8272 );
nor \U$7472 ( \8274 , \8271 , \8273 );
nor \U$7473 ( \8275 , \8260 , \8238 , RIb55be08_602);
and \U$7474 ( \8276 , \8275 , RIb551b60_255);
nor \U$7475 ( \8277 , \8245 , RIb55be08_602);
and \U$7476 ( \8278 , \8277 , \8253 );
and \U$7477 ( \8279 , RIb551e30_261, \8278 );
nor \U$7478 ( \8280 , \8276 , \8279 );
nand \U$7479 ( \8281 , \8251 , \8269 );
nor \U$7480 ( \8282 , \8281 , \8237 );
nand \U$7481 ( \8283 , RIb551818_248, \8282 );
nand \U$7482 ( \8284 , \8267 , \8274 , \8280 , \8283 );
nor \U$7483 ( \8285 , \8244 , \8250 , \8284 );
not \U$7484 ( \8286 , \8269 );
nor \U$7485 ( \8287 , \8286 , \8238 );
and \U$7486 ( \8288 , \8287 , RIb551bd8_256);
not \U$7487 ( \8289 , \8268 );
nor \U$7488 ( \8290 , \8289 , \8240 );
and \U$7489 ( \8291 , RIb5519f8_252, \8290 );
nor \U$7490 ( \8292 , \8288 , \8291 );
nor \U$7491 ( \8293 , \8240 , \8260 );
and \U$7492 ( \8294 , \8293 , RIb551980_251);
not \U$7493 ( \8295 , \8277 );
nor \U$7494 ( \8296 , \8295 , \8238 );
and \U$7495 ( \8297 , RIb551a70_253, \8296 );
nor \U$7496 ( \8298 , \8294 , \8297 );
not \U$7497 ( \8299 , \8268 );
nor \U$7498 ( \8300 , \8299 , \8254 );
and \U$7499 ( \8301 , \8300 , RIb551db8_260);
nor \U$7500 ( \8302 , \8254 , \8260 );
and \U$7501 ( \8303 , RIb551d40_259, \8302 );
nor \U$7502 ( \8304 , \8301 , \8303 );
nand \U$7503 ( \8305 , \8285 , \8292 , \8298 , \8304 );
buf \U$7504 ( \8306 , \8305 );
and \U$7505 ( \8307 , \8281 , RIb55bef8_604);
buf \U$7506 ( \8308 , \8307 );
_DC r2ce1 ( \8309_nR2ce1 , \8306 , \8308 );
xor \U$7507 ( \8310 , \8236 , \8309_nR2ce1 );
not \U$7508 ( \8311 , \8229 );
not \U$7509 ( \8312 , RIb55b7f0_589);
and \U$7510 ( \8313 , \8311 , \8312 );
and \U$7511 ( \8314 , \8229 , RIb55b7f0_589);
nor \U$7512 ( \8315 , \8313 , \8314 );
and \U$7513 ( \8316 , RIb54adb0_21, \8290 );
and \U$7514 ( \8317 , RIb54ae28_22, \8296 );
and \U$7515 ( \8318 , \8302 , RIb54b0f8_28);
and \U$7516 ( \8319 , RIb54b080_27, \8255 );
nor \U$7517 ( \8320 , \8318 , \8319 );
and \U$7518 ( \8321 , RIb54b2d8_32, \8261 );
and \U$7519 ( \8322 , RIb54b260_31, \8272 );
and \U$7520 ( \8323 , \8275 , RIb54af18_24);
and \U$7521 ( \8324 , RIb54aea0_23, \8263 );
nor \U$7522 ( \8325 , \8323 , \8324 );
not \U$7523 ( \8326 , \8325 );
nor \U$7524 ( \8327 , \8321 , \8322 , \8326 );
and \U$7525 ( \8328 , \8287 , RIb54af90_25);
and \U$7526 ( \8329 , RIb54ac48_18, \8249 );
nor \U$7527 ( \8330 , \8328 , \8329 );
nand \U$7528 ( \8331 , RIb54a978_12, \8282 );
nand \U$7529 ( \8332 , \8320 , \8327 , \8330 , \8331 );
nor \U$7530 ( \8333 , \8316 , \8317 , \8332 );
and \U$7531 ( \8334 , \8300 , RIb54b170_29);
and \U$7532 ( \8335 , RIb54b008_26, \8257 );
nor \U$7533 ( \8336 , \8334 , \8335 );
and \U$7534 ( \8337 , \8270 , RIb54b350_33);
and \U$7535 ( \8338 , RIb54b1e8_30, \8278 );
nor \U$7536 ( \8339 , \8337 , \8338 );
and \U$7537 ( \8340 , \8293 , RIb54ad38_20);
and \U$7538 ( \8341 , RIb54acc0_19, \8243 );
nor \U$7539 ( \8342 , \8340 , \8341 );
nand \U$7540 ( \8343 , \8333 , \8336 , \8339 , \8342 );
buf \U$7541 ( \8344 , \8343 );
_DC r2af6 ( \8345_nR2af6 , \8344 , \8308 );
xor \U$7542 ( \8346 , \8315 , \8345_nR2af6 );
not \U$7543 ( \8347 , \8227 );
not \U$7544 ( \8348 , RIb55b868_590);
and \U$7545 ( \8349 , \8347 , \8348 );
and \U$7546 ( \8350 , \8227 , RIb55b868_590);
nor \U$7547 ( \8351 , \8349 , \8350 );
and \U$7548 ( \8352 , RIb54ba58_48, \8272 );
and \U$7549 ( \8353 , RIb54b710_41, \8275 );
and \U$7550 ( \8354 , RIb54b4b8_36, \8243 );
and \U$7551 ( \8355 , RIb54b440_35, \8249 );
and \U$7552 ( \8356 , \8302 , RIb54b8f0_45);
and \U$7553 ( \8357 , RIb54b878_44, \8255 );
nor \U$7554 ( \8358 , \8356 , \8357 );
not \U$7555 ( \8359 , \8358 );
nor \U$7556 ( \8360 , \8354 , \8355 , \8359 );
nand \U$7557 ( \8361 , RIb54b3c8_34, \8282 );
and \U$7558 ( \8362 , \8287 , RIb54b788_42);
and \U$7559 ( \8363 , RIb54b800_43, \8257 );
nor \U$7560 ( \8364 , \8362 , \8363 );
and \U$7561 ( \8365 , \8290 , RIb54b5a8_38);
and \U$7562 ( \8366 , RIb54b530_37, \8293 );
nor \U$7563 ( \8367 , \8365 , \8366 );
nand \U$7564 ( \8368 , \8360 , \8361 , \8364 , \8367 );
nor \U$7565 ( \8369 , \8352 , \8353 , \8368 );
and \U$7566 ( \8370 , \8270 , RIb54bb48_50);
and \U$7567 ( \8371 , RIb54bad0_49, \8261 );
nor \U$7568 ( \8372 , \8370 , \8371 );
and \U$7569 ( \8373 , \8263 , RIb54b698_40);
and \U$7570 ( \8374 , RIb54b620_39, \8296 );
nor \U$7571 ( \8375 , \8373 , \8374 );
and \U$7572 ( \8376 , \8300 , RIb54b968_46);
and \U$7573 ( \8377 , RIb54b9e0_47, \8278 );
nor \U$7574 ( \8378 , \8376 , \8377 );
nand \U$7575 ( \8379 , \8369 , \8372 , \8375 , \8378 );
buf \U$7576 ( \8380 , \8379 );
_DC r2af4 ( \8381_nR2af4 , \8380 , \8308 );
xor \U$7577 ( \8382 , \8351 , \8381_nR2af4 );
not \U$7578 ( \8383 , \8225 );
not \U$7579 ( \8384 , RIb55b8e0_591);
and \U$7580 ( \8385 , \8383 , \8384 );
and \U$7581 ( \8386 , \8225 , RIb55b8e0_591);
nor \U$7582 ( \8387 , \8385 , \8386 );
and \U$7583 ( \8388 , RIb54bf08_58, \8275 );
and \U$7584 ( \8389 , RIb54c1d8_64, \8278 );
and \U$7585 ( \8390 , RIb54c070_61, \8255 );
and \U$7586 ( \8391 , RIb54bff8_60, \8257 );
and \U$7587 ( \8392 , \8290 , RIb54bda0_55);
and \U$7588 ( \8393 , RIb54bd28_54, \8293 );
nor \U$7589 ( \8394 , \8392 , \8393 );
not \U$7590 ( \8395 , \8394 );
nor \U$7591 ( \8396 , \8390 , \8391 , \8395 );
nand \U$7592 ( \8397 , RIb54bbc0_51, \8282 );
and \U$7593 ( \8398 , \8243 , RIb54bcb0_53);
and \U$7594 ( \8399 , RIb54bc38_52, \8249 );
nor \U$7595 ( \8400 , \8398 , \8399 );
and \U$7596 ( \8401 , \8300 , RIb54c160_63);
and \U$7597 ( \8402 , RIb54c0e8_62, \8302 );
nor \U$7598 ( \8403 , \8401 , \8402 );
nand \U$7599 ( \8404 , \8396 , \8397 , \8400 , \8403 );
nor \U$7600 ( \8405 , \8388 , \8389 , \8404 );
and \U$7601 ( \8406 , \8287 , RIb54bf80_59);
and \U$7602 ( \8407 , RIb54be18_56, \8296 );
nor \U$7603 ( \8408 , \8406 , \8407 );
and \U$7604 ( \8409 , \8261 , RIb54c2c8_66);
and \U$7605 ( \8410 , RIb54c250_65, \8272 );
nor \U$7606 ( \8411 , \8409 , \8410 );
and \U$7607 ( \8412 , \8270 , RIb54c340_67);
and \U$7608 ( \8413 , RIb54be90_57, \8263 );
nor \U$7609 ( \8414 , \8412 , \8413 );
nand \U$7610 ( \8415 , \8405 , \8408 , \8411 , \8414 );
buf \U$7611 ( \8416 , \8415 );
_DC r293b ( \8417_nR293b , \8416 , \8308 );
xor \U$7612 ( \8418 , \8387 , \8417_nR293b );
and \U$7613 ( \8419 , \8223 , RIb55b958_592);
not \U$7614 ( \8420 , \8223 );
not \U$7615 ( \8421 , RIb55b958_592);
and \U$7616 ( \8422 , \8420 , \8421 );
nor \U$7617 ( \8423 , \8419 , \8422 );
and \U$7618 ( \8424 , RIb54ca48_82, \8272 );
and \U$7619 ( \8425 , RIb54c700_75, \8275 );
and \U$7620 ( \8426 , RIb54c778_76, \8287 );
and \U$7621 ( \8427 , RIb54c7f0_77, \8257 );
and \U$7622 ( \8428 , \8243 , RIb54c4a8_70);
and \U$7623 ( \8429 , RIb54c430_69, \8249 );
nor \U$7624 ( \8430 , \8428 , \8429 );
not \U$7625 ( \8431 , \8430 );
nor \U$7626 ( \8432 , \8426 , \8427 , \8431 );
and \U$7627 ( \8433 , \8302 , RIb54c8e0_79);
and \U$7628 ( \8434 , RIb54c868_78, \8255 );
nor \U$7629 ( \8435 , \8433 , \8434 );
nand \U$7630 ( \8436 , RIb54c3b8_68, \8282 );
and \U$7631 ( \8437 , \8290 , RIb54c598_72);
and \U$7632 ( \8438 , RIb54c520_71, \8293 );
nor \U$7633 ( \8439 , \8437 , \8438 );
nand \U$7634 ( \8440 , \8432 , \8435 , \8436 , \8439 );
nor \U$7635 ( \8441 , \8424 , \8425 , \8440 );
and \U$7636 ( \8442 , \8270 , RIb54cb38_84);
and \U$7637 ( \8443 , RIb54cac0_83, \8261 );
nor \U$7638 ( \8444 , \8442 , \8443 );
and \U$7639 ( \8445 , \8263 , RIb54c688_74);
and \U$7640 ( \8446 , RIb54c610_73, \8296 );
nor \U$7641 ( \8447 , \8445 , \8446 );
and \U$7642 ( \8448 , \8300 , RIb54c958_80);
and \U$7643 ( \8449 , RIb54c9d0_81, \8278 );
nor \U$7644 ( \8450 , \8448 , \8449 );
nand \U$7645 ( \8451 , \8441 , \8444 , \8447 , \8450 );
buf \U$7646 ( \8452 , \8451 );
_DC r2939 ( \8453_nR2939 , \8452 , \8308 );
xor \U$7647 ( \8454 , \8423 , \8453_nR2939 );
not \U$7648 ( \8455 , \8221 );
not \U$7649 ( \8456 , RIb55b9d0_593);
and \U$7650 ( \8457 , \8455 , \8456 );
and \U$7651 ( \8458 , \8221 , RIb55b9d0_593);
nor \U$7652 ( \8459 , \8457 , \8458 );
and \U$7653 ( \8460 , RIb54d240_99, \8272 );
and \U$7654 ( \8461 , RIb54cef8_92, \8275 );
and \U$7655 ( \8462 , RIb54d060_95, \8255 );
and \U$7656 ( \8463 , RIb54cfe8_94, \8257 );
and \U$7657 ( \8464 , \8243 , RIb54cca0_87);
and \U$7658 ( \8465 , RIb54cc28_86, \8249 );
nor \U$7659 ( \8466 , \8464 , \8465 );
not \U$7660 ( \8467 , \8466 );
nor \U$7661 ( \8468 , \8462 , \8463 , \8467 );
nand \U$7662 ( \8469 , RIb54cbb0_85, \8282 );
and \U$7663 ( \8470 , \8287 , RIb54cf70_93);
and \U$7664 ( \8471 , RIb54ce08_90, \8296 );
nor \U$7665 ( \8472 , \8470 , \8471 );
and \U$7666 ( \8473 , \8290 , RIb54cd90_89);
and \U$7667 ( \8474 , RIb54cd18_88, \8293 );
nor \U$7668 ( \8475 , \8473 , \8474 );
nand \U$7669 ( \8476 , \8468 , \8469 , \8472 , \8475 );
nor \U$7670 ( \8477 , \8460 , \8461 , \8476 );
and \U$7671 ( \8478 , \8270 , RIb54d330_101);
and \U$7672 ( \8479 , RIb54d2b8_100, \8261 );
nor \U$7673 ( \8480 , \8478 , \8479 );
and \U$7674 ( \8481 , \8263 , RIb54ce80_91);
and \U$7675 ( \8482 , RIb54d1c8_98, \8278 );
nor \U$7676 ( \8483 , \8481 , \8482 );
and \U$7677 ( \8484 , \8300 , RIb54d150_97);
and \U$7678 ( \8485 , RIb54d0d8_96, \8302 );
nor \U$7679 ( \8486 , \8484 , \8485 );
nand \U$7680 ( \8487 , \8477 , \8480 , \8483 , \8486 );
buf \U$7681 ( \8488 , \8487 );
_DC r27af ( \8489_nR27af , \8488 , \8308 );
xor \U$7682 ( \8490 , \8459 , \8489_nR27af );
not \U$7683 ( \8491 , \8219 );
not \U$7684 ( \8492 , RIb55ba48_594);
and \U$7685 ( \8493 , \8491 , \8492 );
and \U$7686 ( \8494 , \8219 , RIb55ba48_594);
nor \U$7687 ( \8495 , \8493 , \8494 );
and \U$7688 ( \8496 , RIb54da38_116, \8272 );
and \U$7689 ( \8497 , RIb54d9c0_115, \8278 );
and \U$7690 ( \8498 , RIb54d858_112, \8255 );
and \U$7691 ( \8499 , RIb54d7e0_111, \8257 );
and \U$7692 ( \8500 , \8243 , RIb54d498_104);
and \U$7693 ( \8501 , RIb54d420_103, \8249 );
nor \U$7694 ( \8502 , \8500 , \8501 );
not \U$7695 ( \8503 , \8502 );
nor \U$7696 ( \8504 , \8498 , \8499 , \8503 );
and \U$7697 ( \8505 , \8300 , RIb54d948_114);
and \U$7698 ( \8506 , RIb54d8d0_113, \8302 );
nor \U$7699 ( \8507 , \8505 , \8506 );
nand \U$7700 ( \8508 , RIb54d3a8_102, \8282 );
and \U$7701 ( \8509 , \8290 , RIb54d588_106);
and \U$7702 ( \8510 , RIb54d510_105, \8293 );
nor \U$7703 ( \8511 , \8509 , \8510 );
nand \U$7704 ( \8512 , \8504 , \8507 , \8508 , \8511 );
nor \U$7705 ( \8513 , \8496 , \8497 , \8512 );
and \U$7706 ( \8514 , \8270 , RIb54db28_118);
and \U$7707 ( \8515 , RIb54dab0_117, \8261 );
nor \U$7708 ( \8516 , \8514 , \8515 );
and \U$7709 ( \8517 , \8275 , RIb54d6f0_109);
and \U$7710 ( \8518 , RIb54d678_108, \8263 );
nor \U$7711 ( \8519 , \8517 , \8518 );
and \U$7712 ( \8520 , \8287 , RIb54d768_110);
and \U$7713 ( \8521 , RIb54d600_107, \8296 );
nor \U$7714 ( \8522 , \8520 , \8521 );
nand \U$7715 ( \8523 , \8513 , \8516 , \8519 , \8522 );
buf \U$7716 ( \8524 , \8523 );
_DC r27ad ( \8525_nR27ad , \8524 , \8308 );
xor \U$7717 ( \8526 , \8495 , \8525_nR27ad );
not \U$7718 ( \8527 , \8217 );
not \U$7719 ( \8528 , RIb55bac0_595);
and \U$7720 ( \8529 , \8527 , \8528 );
and \U$7721 ( \8530 , \8217 , RIb55bac0_595);
nor \U$7722 ( \8531 , \8529 , \8530 );
and \U$7723 ( \8532 , RIb54e140_131, \8300 );
and \U$7724 ( \8533 , RIb54e0c8_130, \8302 );
and \U$7725 ( \8534 , RIb54e320_135, \8270 );
and \U$7726 ( \8535 , RIb54e2a8_134, \8261 );
and \U$7727 ( \8536 , \8275 , RIb54dee8_126);
and \U$7728 ( \8537 , RIb54de70_125, \8263 );
nor \U$7729 ( \8538 , \8536 , \8537 );
not \U$7730 ( \8539 , \8538 );
nor \U$7731 ( \8540 , \8534 , \8535 , \8539 );
and \U$7732 ( \8541 , \8255 , RIb54e050_129);
and \U$7733 ( \8542 , RIb54dfd8_128, \8257 );
nor \U$7734 ( \8543 , \8541 , \8542 );
and \U$7735 ( \8544 , \8287 , RIb54df60_127);
and \U$7736 ( \8545 , RIb54ddf8_124, \8296 );
nor \U$7737 ( \8546 , \8544 , \8545 );
nand \U$7738 ( \8547 , RIb54dba0_119, \8282 );
nand \U$7739 ( \8548 , \8540 , \8543 , \8546 , \8547 );
nor \U$7740 ( \8549 , \8532 , \8533 , \8548 );
and \U$7741 ( \8550 , \8243 , RIb54dc90_121);
and \U$7742 ( \8551 , RIb54dc18_120, \8249 );
nor \U$7743 ( \8552 , \8550 , \8551 );
and \U$7744 ( \8553 , \8272 , RIb54e230_133);
and \U$7745 ( \8554 , RIb54e1b8_132, \8278 );
nor \U$7746 ( \8555 , \8553 , \8554 );
and \U$7747 ( \8556 , \8290 , RIb54dd80_123);
and \U$7748 ( \8557 , RIb54dd08_122, \8293 );
nor \U$7749 ( \8558 , \8556 , \8557 );
nand \U$7750 ( \8559 , \8549 , \8552 , \8555 , \8558 );
buf \U$7751 ( \8560 , \8559 );
_DC r2667 ( \8561_nR2667 , \8560 , \8308 );
xor \U$7752 ( \8562 , \8531 , \8561_nR2667 );
not \U$7753 ( \8563 , \8215 );
not \U$7754 ( \8564 , RIb55bb38_596);
and \U$7755 ( \8565 , \8563 , \8564 );
and \U$7756 ( \8566 , \8215 , RIb55bb38_596);
nor \U$7757 ( \8567 , \8565 , \8566 );
and \U$7758 ( \8568 , RIb54e938_148, \8300 );
and \U$7759 ( \8569 , RIb54e8c0_147, \8302 );
and \U$7760 ( \8570 , RIb54eb18_152, \8270 );
and \U$7761 ( \8571 , RIb54eaa0_151, \8261 );
and \U$7762 ( \8572 , \8275 , RIb54e6e0_143);
and \U$7763 ( \8573 , RIb54e668_142, \8263 );
nor \U$7764 ( \8574 , \8572 , \8573 );
not \U$7765 ( \8575 , \8574 );
nor \U$7766 ( \8576 , \8570 , \8571 , \8575 );
nand \U$7767 ( \8577 , RIb54e398_136, \8282 );
and \U$7768 ( \8578 , \8287 , RIb54e758_144);
and \U$7769 ( \8579 , RIb54e7d0_145, \8257 );
nor \U$7770 ( \8580 , \8578 , \8579 );
and \U$7771 ( \8581 , \8255 , RIb54e848_146);
and \U$7772 ( \8582 , RIb54e500_139, \8293 );
nor \U$7773 ( \8583 , \8581 , \8582 );
nand \U$7774 ( \8584 , \8576 , \8577 , \8580 , \8583 );
nor \U$7775 ( \8585 , \8568 , \8569 , \8584 );
and \U$7776 ( \8586 , \8243 , RIb54e488_138);
and \U$7777 ( \8587 , RIb54e410_137, \8249 );
nor \U$7778 ( \8588 , \8586 , \8587 );
and \U$7779 ( \8589 , \8272 , RIb54ea28_150);
and \U$7780 ( \8590 , RIb54e9b0_149, \8278 );
nor \U$7781 ( \8591 , \8589 , \8590 );
and \U$7782 ( \8592 , \8290 , RIb54e578_140);
and \U$7783 ( \8593 , RIb54e5f0_141, \8296 );
nor \U$7784 ( \8594 , \8592 , \8593 );
nand \U$7785 ( \8595 , \8585 , \8588 , \8591 , \8594 );
buf \U$7786 ( \8596 , \8595 );
_DC r2665 ( \8597_nR2665 , \8596 , \8308 );
xor \U$7787 ( \8598 , \8567 , \8597_nR2665 );
not \U$7788 ( \8599 , \8213 );
not \U$7789 ( \8600 , RIb55bbb0_597);
and \U$7790 ( \8601 , \8599 , \8600 );
and \U$7791 ( \8602 , \8213 , RIb55bbb0_597);
nor \U$7792 ( \8603 , \8601 , \8602 );
and \U$7793 ( \8604 , RIb54eed8_160, \8275 );
and \U$7794 ( \8605 , RIb54ee60_159, \8263 );
and \U$7795 ( \8606 , RIb54ed70_157, \8290 );
and \U$7796 ( \8607 , RIb54ecf8_156, \8293 );
and \U$7797 ( \8608 , \8243 , RIb54ec80_155);
and \U$7798 ( \8609 , RIb54ec08_154, \8249 );
nor \U$7799 ( \8610 , \8608 , \8609 );
not \U$7800 ( \8611 , \8610 );
nor \U$7801 ( \8612 , \8606 , \8607 , \8611 );
nand \U$7802 ( \8613 , RIb54eb90_153, \8282 );
and \U$7803 ( \8614 , \8272 , RIb54f220_167);
and \U$7804 ( \8615 , RIb54f1a8_166, \8278 );
nor \U$7805 ( \8616 , \8614 , \8615 );
and \U$7806 ( \8617 , \8300 , RIb54f130_165);
and \U$7807 ( \8618 , RIb54f0b8_164, \8302 );
nor \U$7808 ( \8619 , \8617 , \8618 );
nand \U$7809 ( \8620 , \8612 , \8613 , \8616 , \8619 );
nor \U$7810 ( \8621 , \8604 , \8605 , \8620 );
and \U$7811 ( \8622 , \8287 , RIb54ef50_161);
and \U$7812 ( \8623 , RIb54ede8_158, \8296 );
nor \U$7813 ( \8624 , \8622 , \8623 );
and \U$7814 ( \8625 , \8270 , RIb54f310_169);
and \U$7815 ( \8626 , RIb54f298_168, \8261 );
nor \U$7816 ( \8627 , \8625 , \8626 );
and \U$7817 ( \8628 , \8255 , RIb54f040_163);
and \U$7818 ( \8629 , RIb54efc8_162, \8257 );
nor \U$7819 ( \8630 , \8628 , \8629 );
nand \U$7820 ( \8631 , \8621 , \8624 , \8627 , \8630 );
buf \U$7821 ( \8632 , \8631 );
_DC r2589 ( \8633_nR2589 , \8632 , \8308 );
xor \U$7822 ( \8634 , \8603 , \8633_nR2589 );
xnor \U$7823 ( \8635 , RIb55bc28_598, RIb55bca0_599);
and \U$7824 ( \8636 , RIb54f6d0_177, \8275 );
and \U$7825 ( \8637 , RIb54f658_176, \8263 );
and \U$7826 ( \8638 , RIb54fa18_184, \8272 );
and \U$7827 ( \8639 , RIb54f9a0_183, \8278 );
and \U$7828 ( \8640 , \8243 , RIb54f478_172);
and \U$7829 ( \8641 , RIb54f400_171, \8249 );
nor \U$7830 ( \8642 , \8640 , \8641 );
not \U$7831 ( \8643 , \8642 );
nor \U$7832 ( \8644 , \8638 , \8639 , \8643 );
and \U$7833 ( \8645 , \8300 , RIb54f928_182);
and \U$7834 ( \8646 , RIb54f8b0_181, \8302 );
nor \U$7835 ( \8647 , \8645 , \8646 );
nand \U$7836 ( \8648 , RIb54f388_170, \8282 );
and \U$7837 ( \8649 , \8290 , RIb54f568_174);
and \U$7838 ( \8650 , RIb54f4f0_173, \8293 );
nor \U$7839 ( \8651 , \8649 , \8650 );
nand \U$7840 ( \8652 , \8644 , \8647 , \8648 , \8651 );
nor \U$7841 ( \8653 , \8636 , \8637 , \8652 );
and \U$7842 ( \8654 , \8287 , RIb54f748_178);
and \U$7843 ( \8655 , RIb54f5e0_175, \8296 );
nor \U$7844 ( \8656 , \8654 , \8655 );
and \U$7845 ( \8657 , \8270 , RIb54fb08_186);
and \U$7846 ( \8658 , RIb54fa90_185, \8261 );
nor \U$7847 ( \8659 , \8657 , \8658 );
and \U$7848 ( \8660 , \8255 , RIb54f838_180);
and \U$7849 ( \8661 , RIb54f7c0_179, \8257 );
nor \U$7850 ( \8662 , \8660 , \8661 );
nand \U$7851 ( \8663 , \8653 , \8656 , \8659 , \8662 );
buf \U$7852 ( \8664 , \8663 );
_DC r258b ( \8665_nR258b , \8664 , \8308 );
xor \U$7853 ( \8666 , \8635 , \8665_nR258b );
and \U$7854 ( \8667 , RIb550738_212, \8275 );
and \U$7855 ( \8668 , RIb5506c0_211, \8263 );
and \U$7856 ( \8669 , RIb5504e0_207, \8243 );
and \U$7857 ( \8670 , RIb550468_206, \8249 );
and \U$7858 ( \8671 , \8300 , RIb550990_217);
and \U$7859 ( \8672 , RIb550918_216, \8302 );
nor \U$7860 ( \8673 , \8671 , \8672 );
not \U$7861 ( \8674 , \8673 );
nor \U$7862 ( \8675 , \8669 , \8670 , \8674 );
nand \U$7863 ( \8676 , RIb5503f0_205, \8282 );
and \U$7864 ( \8677 , \8272 , RIb550a80_219);
and \U$7865 ( \8678 , RIb550a08_218, \8278 );
nor \U$7866 ( \8679 , \8677 , \8678 );
and \U$7867 ( \8680 , \8290 , RIb5505d0_209);
and \U$7868 ( \8681 , RIb550558_208, \8293 );
nor \U$7869 ( \8682 , \8680 , \8681 );
nand \U$7870 ( \8683 , \8675 , \8676 , \8679 , \8682 );
nor \U$7871 ( \8684 , \8667 , \8668 , \8683 );
and \U$7872 ( \8685 , \8287 , RIb5507b0_213);
and \U$7873 ( \8686 , RIb550648_210, \8296 );
nor \U$7874 ( \8687 , \8685 , \8686 );
and \U$7875 ( \8688 , \8270 , RIb550b70_221);
and \U$7876 ( \8689 , RIb550af8_220, \8261 );
nor \U$7877 ( \8690 , \8688 , \8689 );
and \U$7878 ( \8691 , \8255 , RIb5508a0_215);
and \U$7879 ( \8692 , RIb550828_214, \8257 );
nor \U$7880 ( \8693 , \8691 , \8692 );
nand \U$7881 ( \8694 , \8684 , \8687 , \8690 , \8693 );
buf \U$7882 ( \8695 , \8694 );
_DC r23dd ( \8696_nR23dd , \8695 , \8308 );
not \U$7883 ( \8697 , RIb55bf70_605);
nand \U$7884 ( \8698 , \8696_nR23dd , \8697 );
and \U$7885 ( \8699 , RIb54fc70_189, \8243 );
and \U$7886 ( \8700 , RIb54fbf8_188, \8249 );
and \U$7887 ( \8701 , RIb550030_197, \8255 );
and \U$7888 ( \8702 , RIb54ffb8_196, \8257 );
and \U$7889 ( \8703 , \8270 , RIb550300_203);
and \U$7890 ( \8704 , RIb550288_202, \8261 );
nor \U$7891 ( \8705 , \8703 , \8704 );
not \U$7892 ( \8706 , \8705 );
nor \U$7893 ( \8707 , \8701 , \8702 , \8706 );
and \U$7894 ( \8708 , \8287 , RIb54ff40_195);
and \U$7895 ( \8709 , RIb54fec8_194, \8275 );
nor \U$7896 ( \8710 , \8708 , \8709 );
and \U$7897 ( \8711 , \8263 , RIb54fe50_193);
and \U$7898 ( \8712 , RIb54fdd8_192, \8296 );
nor \U$7899 ( \8713 , \8711 , \8712 );
nand \U$7900 ( \8714 , RIb54fb80_187, \8282 );
nand \U$7901 ( \8715 , \8707 , \8710 , \8713 , \8714 );
nor \U$7902 ( \8716 , \8699 , \8700 , \8715 );
and \U$7903 ( \8717 , \8300 , RIb550120_199);
and \U$7904 ( \8718 , RIb5500a8_198, \8302 );
nor \U$7905 ( \8719 , \8717 , \8718 );
and \U$7906 ( \8720 , \8272 , RIb550210_201);
and \U$7907 ( \8721 , RIb550198_200, \8278 );
nor \U$7908 ( \8722 , \8720 , \8721 );
and \U$7909 ( \8723 , \8290 , RIb54fd60_191);
and \U$7910 ( \8724 , RIb54fce8_190, \8293 );
nor \U$7911 ( \8725 , \8723 , \8724 );
nand \U$7912 ( \8726 , \8716 , \8719 , \8722 , \8725 );
buf \U$7913 ( \8727 , \8726 );
_DC r23df ( \8728_nR23df , \8727 , \8308 );
nand \U$7914 ( \8729 , \8728_nR23df , RIb55bca0_599);
and \U$7915 ( \8730 , \8698 , \8729 );
nor \U$7916 ( \8731 , RIb55bca0_599, \8728_nR23df );
nor \U$7917 ( \8732 , \8730 , \8731 );
and \U$7918 ( \8733 , \8666 , \8732 );
and \U$7919 ( \8734 , \8635 , \8665_nR258b );
or \U$7920 ( \8735 , \8733 , \8734 );
and \U$7921 ( \8736 , \8634 , \8735 );
and \U$7922 ( \8737 , \8603 , \8633_nR2589 );
or \U$7923 ( \8738 , \8736 , \8737 );
and \U$7924 ( \8739 , \8598 , \8738 );
and \U$7925 ( \8740 , \8567 , \8597_nR2665 );
or \U$7926 ( \8741 , \8739 , \8740 );
and \U$7927 ( \8742 , \8562 , \8741 );
and \U$7928 ( \8743 , \8531 , \8561_nR2667 );
or \U$7929 ( \8744 , \8742 , \8743 );
and \U$7930 ( \8745 , \8526 , \8744 );
and \U$7931 ( \8746 , \8495 , \8525_nR27ad );
or \U$7932 ( \8747 , \8745 , \8746 );
and \U$7933 ( \8748 , \8490 , \8747 );
and \U$7934 ( \8749 , \8459 , \8489_nR27af );
or \U$7935 ( \8750 , \8748 , \8749 );
and \U$7936 ( \8751 , \8454 , \8750 );
and \U$7937 ( \8752 , \8423 , \8453_nR2939 );
or \U$7938 ( \8753 , \8751 , \8752 );
and \U$7939 ( \8754 , \8418 , \8753 );
and \U$7940 ( \8755 , \8387 , \8417_nR293b );
or \U$7941 ( \8756 , \8754 , \8755 );
and \U$7942 ( \8757 , \8382 , \8756 );
and \U$7943 ( \8758 , \8351 , \8381_nR2af4 );
or \U$7944 ( \8759 , \8757 , \8758 );
and \U$7945 ( \8760 , \8346 , \8759 );
and \U$7946 ( \8761 , \8315 , \8345_nR2af6 );
or \U$7947 ( \8762 , \8760 , \8761 );
and \U$7948 ( \8763 , \8310 , \8762 );
and \U$7949 ( \8764 , \8236 , \8309_nR2ce1 );
or \U$7950 ( \8765 , \8763 , \8764 );
not \U$7951 ( \8766 , \8231 );
nand \U$7952 ( \8767 , \8766 , RIb55c3a8_614);
nor \U$7953 ( \8768 , \8765 , \8767 );
not \U$7954 ( \8769 , \8768 );
or \U$7955 ( \8770 , RIb55bfe8_606, RIb55c060_607, RIb55c0d8_608, RIb55c150_609);
or \U$7956 ( \8771 , RIb55c1c8_610, RIb55c240_611, RIb55c2b8_612, RIb55c330_613);
nor \U$7957 ( \8772 , \8770 , \8771 , RIb55bef8_604);
or \U$7958 ( \8773 , \8772 , \8246 );
and \U$7959 ( \8774 , \8772 , \8277 );
and \U$7960 ( \8775 , RIb55be08_602, \8245 );
nor \U$7961 ( \8776 , \8774 , \8775 );
nand \U$7962 ( \8777 , \8773 , \8776 );
not \U$7963 ( \8778 , \8777 );
and \U$7964 ( \8779 , \8772 , \8247 );
or \U$7965 ( \8780 , \8779 , \8251 );
and \U$7966 ( \8781 , \8247 , RIb55be80_603);
not \U$7967 ( \8782 , \8772 );
nor \U$7968 ( \8783 , \8781 , \8782 );
nand \U$7969 ( \8784 , \8247 , \8783 );
nand \U$7970 ( \8785 , \8780 , \8784 );
and \U$7971 ( \8786 , \8249 , \8772 );
nor \U$7972 ( \8787 , \8786 , RIb55bef8_604);
not \U$7973 ( \8788 , \8787 );
nor \U$7974 ( \8789 , \8778 , \8785 , \8788 );
and \U$7975 ( \8790 , \8782 , RIb55bd90_601);
nor \U$7976 ( \8791 , \8782 , \8260 );
nor \U$7977 ( \8792 , \8790 , \8791 );
not \U$7978 ( \8793 , \8792 );
not \U$7979 ( \8794 , \8242 );
or \U$7980 ( \8795 , \8793 , \8794 );
and \U$7981 ( \8796 , \8772 , \8241 );
and \U$7982 ( \8797 , RIb55bd18_600, \8782 );
nor \U$7983 ( \8798 , \8796 , \8797 );
nor \U$7984 ( \8799 , \8795 , \8798 );
and \U$7985 ( \8800 , \8789 , \8799 );
and \U$7986 ( \8801 , \8800 , RIb5514d0_241);
nand \U$7987 ( \8802 , \8787 , \8785 , \8777 );
not \U$7988 ( \8803 , \8798 );
nor \U$7989 ( \8804 , \8803 , \8795 );
not \U$7990 ( \8805 , \8804 );
nor \U$7991 ( \8806 , \8802 , \8805 );
and \U$7992 ( \8807 , \8806 , RIb551188_234);
not \U$7993 ( \8808 , \8785 );
nor \U$7994 ( \8809 , \8808 , \8777 , \8788 );
not \U$7995 ( \8810 , \8795 );
nor \U$7996 ( \8811 , \8810 , \8798 );
and \U$7997 ( \8812 , \8809 , \8811 );
and \U$7998 ( \8813 , RIb551200_235, \8812 );
nor \U$7999 ( \8814 , \8807 , \8813 );
nor \U$8000 ( \8815 , \8785 , \8777 );
and \U$8001 ( \8816 , \8804 , \8815 , \8788 );
and \U$8002 ( \8817 , \8816 , RIb550be8_222);
and \U$8003 ( \8818 , \8809 , \8804 );
and \U$8004 ( \8819 , RIb551368_238, \8818 );
nor \U$8005 ( \8820 , \8817 , \8819 );
not \U$8006 ( \8821 , \8789 );
nand \U$8007 ( \8822 , \8798 , \8795 );
nor \U$8008 ( \8823 , \8821 , \8822 );
and \U$8009 ( \8824 , \8823 , RIb551458_240);
and \U$8010 ( \8825 , \8789 , \8811 );
and \U$8011 ( \8826 , RIb5513e0_239, \8825 );
nor \U$8012 ( \8827 , \8824 , \8826 );
not \U$8013 ( \8828 , \8799 );
nor \U$8014 ( \8829 , \8828 , \8802 );
and \U$8015 ( \8830 , \8829 , RIb551110_233);
nor \U$8016 ( \8831 , \8802 , \8822 );
and \U$8017 ( \8832 , RIb551098_232, \8831 );
nor \U$8018 ( \8833 , \8830 , \8832 );
nand \U$8019 ( \8834 , \8814 , \8820 , \8827 , \8833 );
and \U$8020 ( \8835 , \8789 , \8804 );
and \U$8021 ( \8836 , \8835 , RIb551548_242);
not \U$8022 ( \8837 , \8811 );
nand \U$8023 ( \8838 , \8787 , \8815 );
nor \U$8024 ( \8839 , \8837 , \8838 );
and \U$8025 ( \8840 , RIb5515c0_243, \8839 );
nor \U$8026 ( \8841 , \8836 , \8840 );
not \U$8027 ( \8842 , \8841 );
nor \U$8028 ( \8843 , \8801 , \8834 , \8842 );
nor \U$8029 ( \8844 , \8838 , \8822 );
and \U$8030 ( \8845 , \8844 , RIb551638_244);
not \U$8031 ( \8846 , \8809 );
nor \U$8032 ( \8847 , \8846 , \8822 );
and \U$8033 ( \8848 , RIb551278_236, \8847 );
nor \U$8034 ( \8849 , \8845 , \8848 );
and \U$8035 ( \8850 , \8809 , \8799 );
and \U$8036 ( \8851 , \8850 , RIb5512f0_237);
not \U$8037 ( \8852 , \8811 );
nor \U$8038 ( \8853 , \8852 , \8802 );
and \U$8039 ( \8854 , RIb551020_231, \8853 );
nor \U$8040 ( \8855 , \8851 , \8854 );
nor \U$8041 ( \8856 , \8838 , \8805 );
and \U$8042 ( \8857 , \8856 , RIb551728_246);
not \U$8043 ( \8858 , \8799 );
nor \U$8044 ( \8859 , \8858 , \8838 );
and \U$8045 ( \8860 , RIb5516b0_245, \8859 );
nor \U$8046 ( \8861 , \8857 , \8860 );
nand \U$8047 ( \8862 , \8843 , \8849 , \8855 , \8861 );
buf \U$8048 ( \8863 , \8307 );
_DC r335c ( \8864_nR335c , \8862 , \8863 );
not \U$8049 ( \8865 , \8864_nR335c );
nor \U$8050 ( \8866 , \8769 , \8865 );
xor \U$8051 ( \8867 , \8236 , \8309_nR2ce1 );
xor \U$8052 ( \8868 , \8867 , \8762 );
not \U$8053 ( \8869 , \8868 );
xor \U$8054 ( \8870 , \8315 , \8345_nR2af6 );
xor \U$8055 ( \8871 , \8870 , \8759 );
not \U$8056 ( \8872 , \8871 );
and \U$8057 ( \8873 , \8869 , \8872 );
and \U$8058 ( \8874 , \8765 , \8767 );
nor \U$8059 ( \8875 , \8874 , \8768 );
nor \U$8060 ( \8876 , \8873 , \8875 );
not \U$8061 ( \8877 , \8876 );
and \U$8062 ( \8878 , \8847 , RIb5522e0_271);
and \U$8063 ( \8879 , \8859 , RIb552718_280);
and \U$8064 ( \8880 , RIb5526a0_279, \8844 );
nor \U$8065 ( \8881 , \8879 , \8880 );
and \U$8066 ( \8882 , \8806 , RIb5521f0_269);
and \U$8067 ( \8883 , RIb552268_270, \8812 );
nor \U$8068 ( \8884 , \8882 , \8883 );
and \U$8069 ( \8885 , \8816 , RIb552010_265);
and \U$8070 ( \8886 , RIb552178_268, \8829 );
nor \U$8071 ( \8887 , \8885 , \8886 );
and \U$8072 ( \8888 , \8835 , RIb5525b0_277);
and \U$8073 ( \8889 , RIb552628_278, \8839 );
nor \U$8074 ( \8890 , \8888 , \8889 );
nand \U$8075 ( \8891 , \8881 , \8884 , \8887 , \8890 );
and \U$8076 ( \8892 , \8818 , RIb5523d0_273);
and \U$8077 ( \8893 , RIb552358_272, \8850 );
nor \U$8078 ( \8894 , \8892 , \8893 );
not \U$8079 ( \8895 , \8894 );
nor \U$8080 ( \8896 , \8878 , \8891 , \8895 );
and \U$8081 ( \8897 , \8831 , RIb552100_267);
and \U$8082 ( \8898 , RIb552088_266, \8853 );
nor \U$8083 ( \8899 , \8897 , \8898 );
and \U$8084 ( \8900 , \8823 , RIb5524c0_275);
and \U$8085 ( \8901 , RIb552448_274, \8825 );
nor \U$8086 ( \8902 , \8900 , \8901 );
and \U$8087 ( \8903 , \8856 , RIb552790_281);
and \U$8088 ( \8904 , RIb552538_276, \8800 );
nor \U$8089 ( \8905 , \8903 , \8904 );
nand \U$8090 ( \8906 , \8896 , \8899 , \8902 , \8905 );
_DC r3482 ( \8907_nR3482 , \8906 , \8863 );
or \U$8091 ( \8908 , \8877 , \8907_nR3482 );
not \U$8092 ( \8909 , \8907_nR3482 );
and \U$8093 ( \8910 , \8875 , \8868 );
nor \U$8094 ( \8911 , \8875 , \8868 );
xor \U$8095 ( \8912 , \8868 , \8871 );
nor \U$8096 ( \8913 , \8910 , \8911 , \8912 );
and \U$8097 ( \8914 , \8913 , \8877 );
not \U$8098 ( \8915 , \8914 );
or \U$8099 ( \8916 , \8909 , \8915 );
or \U$8100 ( \8917 , \8913 , \8877 );
nand \U$8101 ( \8918 , \8908 , \8916 , \8917 );
xnor \U$8102 ( \8919 , \8866 , \8918 );
not \U$8103 ( \8920 , \8912 );
nor \U$8104 ( \8921 , \8876 , \8920 );
not \U$8105 ( \8922 , \8921 );
or \U$8106 ( \8923 , \8922 , \8909 );
or \U$8107 ( \8924 , \8865 , \8915 );
or \U$8108 ( \8925 , \8920 , \8909 );
or \U$8109 ( \8926 , \8877 , \8864_nR335c );
nand \U$8110 ( \8927 , \8926 , \8917 );
nand \U$8111 ( \8928 , \8925 , \8927 );
nand \U$8112 ( \8929 , \8923 , \8924 , \8928 );
xor \U$8113 ( \8930 , \8351 , \8381_nR2af4 );
xor \U$8114 ( \8931 , \8930 , \8756 );
xor \U$8115 ( \8932 , \8387 , \8417_nR293b );
xor \U$8116 ( \8933 , \8932 , \8753 );
nor \U$8117 ( \8934 , \8931 , \8933 );
or \U$8118 ( \8935 , \8871 , \8934 );
and \U$8119 ( \8936 , \8929 , \8935 );
and \U$8120 ( \8937 , \8825 , RIb552c40_291);
and \U$8121 ( \8938 , \8859 , RIb552f10_297);
and \U$8122 ( \8939 , RIb552e98_296, \8844 );
nor \U$8123 ( \8940 , \8938 , \8939 );
and \U$8124 ( \8941 , \8806 , RIb5529e8_286);
and \U$8125 ( \8942 , RIb552970_285, \8829 );
nor \U$8126 ( \8943 , \8941 , \8942 );
and \U$8127 ( \8944 , \8816 , RIb552808_282);
and \U$8128 ( \8945 , RIb552a60_287, \8812 );
nor \U$8129 ( \8946 , \8944 , \8945 );
and \U$8130 ( \8947 , \8835 , RIb552da8_294);
and \U$8131 ( \8948 , RIb552e20_295, \8839 );
nor \U$8132 ( \8949 , \8947 , \8948 );
nand \U$8133 ( \8950 , \8940 , \8943 , \8946 , \8949 );
and \U$8134 ( \8951 , \8800 , RIb552d30_293);
and \U$8135 ( \8952 , RIb552cb8_292, \8823 );
nor \U$8136 ( \8953 , \8951 , \8952 );
not \U$8137 ( \8954 , \8953 );
nor \U$8138 ( \8955 , \8937 , \8950 , \8954 );
and \U$8139 ( \8956 , \8850 , RIb552b50_289);
and \U$8140 ( \8957 , RIb552ad8_288, \8847 );
nor \U$8141 ( \8958 , \8956 , \8957 );
and \U$8142 ( \8959 , \8831 , RIb5528f8_284);
and \U$8143 ( \8960 , RIb552880_283, \8853 );
nor \U$8144 ( \8961 , \8959 , \8960 );
and \U$8145 ( \8962 , \8856 , RIb552f88_298);
and \U$8146 ( \8963 , RIb552bc8_290, \8818 );
nor \U$8147 ( \8964 , \8962 , \8963 );
nand \U$8148 ( \8965 , \8955 , \8958 , \8961 , \8964 );
_DC r3254 ( \8966_nR3254 , \8965 , \8863 );
not \U$8149 ( \8967 , \8966_nR3254 );
nor \U$8150 ( \8968 , \8769 , \8967 );
nor \U$8151 ( \8969 , \8936 , \8968 );
xor \U$8152 ( \8970 , \8919 , \8969 );
not \U$8153 ( \8971 , \8970 );
not \U$8154 ( \8972 , \8931 );
not \U$8155 ( \8973 , \8871 );
or \U$8156 ( \8974 , \8972 , \8973 );
or \U$8157 ( \8975 , \8871 , \8931 );
nand \U$8158 ( \8976 , \8974 , \8975 );
xor \U$8159 ( \8977 , \8933 , \8931 );
nor \U$8160 ( \8978 , \8976 , \8977 );
not \U$8161 ( \8979 , \8978 );
not \U$8162 ( \8980 , \8935 );
nor \U$8163 ( \8981 , \8979 , \8980 );
not \U$8164 ( \8982 , \8981 );
or \U$8165 ( \8983 , \8982 , \8909 );
or \U$8166 ( \8984 , \8979 , \8909 );
nand \U$8167 ( \8985 , \8984 , \8980 );
nand \U$8168 ( \8986 , \8983 , \8985 );
or \U$8169 ( \8987 , \8922 , \8865 );
or \U$8170 ( \8988 , \8967 , \8915 );
or \U$8171 ( \8989 , \8920 , \8865 );
or \U$8172 ( \8990 , \8877 , \8966_nR3254 );
nand \U$8173 ( \8991 , \8990 , \8917 );
nand \U$8174 ( \8992 , \8989 , \8991 );
nand \U$8175 ( \8993 , \8987 , \8988 , \8992 );
and \U$8176 ( \8994 , \8986 , \8993 );
and \U$8177 ( \8995 , \8929 , \8935 );
not \U$8178 ( \8996 , \8929 );
and \U$8179 ( \8997 , \8996 , \8980 );
nor \U$8180 ( \8998 , \8995 , \8997 );
xor \U$8181 ( \8999 , \8968 , \8998 );
and \U$8182 ( \9000 , \8994 , \8999 );
and \U$8183 ( \9001 , \8971 , \9000 );
or \U$8184 ( \9002 , \9001 , \8876 );
and \U$8185 ( \9003 , \8918 , \8866 );
and \U$8186 ( \9004 , \8876 , \9001 );
nor \U$8187 ( \9005 , \9003 , \9004 );
nand \U$8188 ( \9006 , \9002 , \9005 );
not \U$8189 ( \9007 , \9006 );
and \U$8190 ( \9008 , \8768 , \8907_nR3482 );
and \U$8191 ( \9009 , \8919 , \8969 );
nor \U$8192 ( \9010 , \9008 , \9009 );
not \U$8193 ( \9011 , \9010 );
and \U$8194 ( \9012 , \9007 , \9011 );
and \U$8195 ( \9013 , \9006 , \9010 );
nor \U$8196 ( \9014 , \9012 , \9013 );
not \U$8197 ( \9015 , \9014 );
and \U$8198 ( \9016 , \8864_nR335c , \8981 );
or \U$8199 ( \9017 , \8935 , \8907_nR3482 );
or \U$8200 ( \9018 , \8935 , \8977 );
nand \U$8201 ( \9019 , \9017 , \9018 );
nand \U$8202 ( \9020 , \8864_nR335c , \8978 );
and \U$8203 ( \9021 , \9019 , \9020 );
and \U$8204 ( \9022 , \8935 , \8977 );
and \U$8205 ( \9023 , \8907_nR3482 , \9022 );
nor \U$8206 ( \9024 , \9016 , \9021 , \9023 );
xor \U$8207 ( \9025 , \8423 , \8453_nR2939 );
xor \U$8208 ( \9026 , \9025 , \8750 );
xor \U$8209 ( \9027 , \8459 , \8489_nR27af );
xor \U$8210 ( \9028 , \9027 , \8747 );
nor \U$8211 ( \9029 , \9026 , \9028 );
or \U$8212 ( \9030 , \8933 , \9029 );
not \U$8213 ( \9031 , \9030 );
xor \U$8214 ( \9032 , \9024 , \9031 );
and \U$8215 ( \9033 , \8966_nR3254 , \8921 );
and \U$8216 ( \9034 , \8853 , RIb553870_317);
and \U$8217 ( \9035 , \8844 , RIb553e88_330);
and \U$8218 ( \9036 , RIb553e10_329, \8839 );
nor \U$8219 ( \9037 , \9035 , \9036 );
and \U$8220 ( \9038 , \8816 , RIb5537f8_316);
and \U$8221 ( \9039 , RIb553a50_321, \8812 );
nor \U$8222 ( \9040 , \9038 , \9039 );
and \U$8223 ( \9041 , \8835 , RIb553d98_328);
and \U$8224 ( \9042 , RIb553d20_327, \8800 );
nor \U$8225 ( \9043 , \9041 , \9042 );
and \U$8226 ( \9044 , \8806 , RIb5539d8_320);
and \U$8227 ( \9045 , RIb553960_319, \8829 );
nor \U$8228 ( \9046 , \9044 , \9045 );
nand \U$8229 ( \9047 , \9037 , \9040 , \9043 , \9046 );
and \U$8230 ( \9048 , \8847 , RIb553ac8_322);
and \U$8231 ( \9049 , RIb5538e8_318, \8831 );
nor \U$8232 ( \9050 , \9048 , \9049 );
not \U$8233 ( \9051 , \9050 );
nor \U$8234 ( \9052 , \9034 , \9047 , \9051 );
and \U$8235 ( \9053 , \8818 , RIb553bb8_324);
and \U$8236 ( \9054 , RIb553b40_323, \8850 );
nor \U$8237 ( \9055 , \9053 , \9054 );
and \U$8238 ( \9056 , \8823 , RIb553ca8_326);
and \U$8239 ( \9057 , RIb553c30_325, \8825 );
nor \U$8240 ( \9058 , \9056 , \9057 );
and \U$8241 ( \9059 , \8856 , RIb553f78_332);
and \U$8242 ( \9060 , RIb553f00_331, \8859 );
nor \U$8243 ( \9061 , \9059 , \9060 );
nand \U$8244 ( \9062 , \9052 , \9055 , \9058 , \9061 );
_DC r3133 ( \9063_nR3133 , \9062 , \8863 );
or \U$8245 ( \9064 , \8877 , \9063_nR3133 );
nand \U$8246 ( \9065 , \9064 , \8917 );
nand \U$8247 ( \9066 , \8966_nR3254 , \8912 );
and \U$8248 ( \9067 , \9065 , \9066 );
and \U$8249 ( \9068 , \9063_nR3133 , \8914 );
nor \U$8250 ( \9069 , \9033 , \9067 , \9068 );
and \U$8251 ( \9070 , \9032 , \9069 );
and \U$8252 ( \9071 , \9024 , \9031 );
or \U$8253 ( \9072 , \9070 , \9071 );
xor \U$8254 ( \9073 , \8986 , \8993 );
not \U$8255 ( \9074 , \9073 );
nand \U$8256 ( \9075 , \9063_nR3133 , \8768 );
not \U$8257 ( \9076 , \9075 );
and \U$8258 ( \9077 , \9074 , \9076 );
and \U$8259 ( \9078 , \9073 , \9075 );
nor \U$8260 ( \9079 , \9077 , \9078 );
nand \U$8261 ( \9080 , \9072 , \9079 );
xor \U$8262 ( \9081 , \8994 , \8999 );
and \U$8263 ( \9082 , \9080 , \9081 );
xor \U$8264 ( \9083 , \8971 , \9000 );
and \U$8265 ( \9084 , \9082 , \9083 );
not \U$8266 ( \9085 , \9084 );
and \U$8267 ( \9086 , \9015 , \9085 );
and \U$8268 ( \9087 , \9014 , \9084 );
nor \U$8269 ( \9088 , \9086 , \9087 );
not \U$8270 ( \9089 , \9088 );
xor \U$8271 ( \9090 , \9024 , \9031 );
xor \U$8272 ( \9091 , \9090 , \9069 );
not \U$8273 ( \9092 , \9091 );
and \U$8274 ( \9093 , \8839 , RIb553618_312);
nand \U$8275 ( \9094 , RIb553780_315, \8856 );
and \U$8276 ( \9095 , \8823 , RIb5534b0_309);
and \U$8277 ( \9096 , RIb553438_308, \8825 );
nor \U$8278 ( \9097 , \9095 , \9096 );
nand \U$8279 ( \9098 , RIb553708_314, \8859 );
nand \U$8280 ( \9099 , \9094 , \9097 , \9098 );
and \U$8281 ( \9100 , \8835 , RIb5535a0_311);
and \U$8282 ( \9101 , RIb553528_310, \8800 );
nor \U$8283 ( \9102 , \9100 , \9101 );
and \U$8284 ( \9103 , \8816 , RIb553000_299);
and \U$8285 ( \9104 , RIb553258_304, \8812 );
nor \U$8286 ( \9105 , \9103 , \9104 );
nand \U$8287 ( \9106 , \9102 , \9105 );
nor \U$8288 ( \9107 , \9093 , \9099 , \9106 );
and \U$8289 ( \9108 , \8818 , RIb5533c0_307);
and \U$8290 ( \9109 , RIb553348_306, \8850 );
nor \U$8291 ( \9110 , \9108 , \9109 );
and \U$8292 ( \9111 , \8806 , RIb5531e0_303);
and \U$8293 ( \9112 , RIb553168_302, \8829 );
nor \U$8294 ( \9113 , \9111 , \9112 );
and \U$8295 ( \9114 , RIb553690_313, \8844 );
and \U$8296 ( \9115 , RIb553078_300, \8853 );
and \U$8297 ( \9116 , \8847 , RIb5532d0_305);
and \U$8298 ( \9117 , RIb5530f0_301, \8831 );
nor \U$8299 ( \9118 , \9116 , \9117 );
not \U$8300 ( \9119 , \9118 );
nor \U$8301 ( \9120 , \9114 , \9115 , \9119 );
nand \U$8302 ( \9121 , \9107 , \9110 , \9113 , \9120 );
_DC r301c ( \9122_nR301c , \9121 , \8863 );
not \U$8303 ( \9123 , \9122_nR301c );
nor \U$8304 ( \9124 , \8769 , \9123 );
not \U$8305 ( \9125 , \9124 );
and \U$8306 ( \9126 , \9092 , \9125 );
and \U$8307 ( \9127 , \9091 , \9124 );
nor \U$8308 ( \9128 , \9126 , \9127 );
not \U$8309 ( \9129 , \9128 );
and \U$8310 ( \9130 , \8966_nR3254 , \8981 );
or \U$8311 ( \9131 , \8935 , \8864_nR335c );
nand \U$8312 ( \9132 , \9131 , \9018 );
nand \U$8313 ( \9133 , \8966_nR3254 , \8978 );
and \U$8314 ( \9134 , \9132 , \9133 );
and \U$8315 ( \9135 , \8864_nR335c , \9022 );
nor \U$8316 ( \9136 , \9130 , \9134 , \9135 );
and \U$8317 ( \9137 , \8933 , \9026 );
nor \U$8318 ( \9138 , \8933 , \9026 );
xor \U$8319 ( \9139 , \9026 , \9028 );
nor \U$8320 ( \9140 , \9137 , \9138 , \9139 );
and \U$8321 ( \9141 , \9140 , \9030 );
and \U$8322 ( \9142 , \8907_nR3482 , \9141 );
and \U$8323 ( \9143 , \8909 , \9031 );
or \U$8324 ( \9144 , \9140 , \9030 );
not \U$8325 ( \9145 , \9144 );
nor \U$8326 ( \9146 , \9142 , \9143 , \9145 );
or \U$8327 ( \9147 , \9136 , \9146 );
and \U$8328 ( \9148 , \8825 , RIb554428_342);
and \U$8329 ( \9149 , \8844 , RIb554680_347);
and \U$8330 ( \9150 , RIb554608_346, \8839 );
nor \U$8331 ( \9151 , \9149 , \9150 );
and \U$8332 ( \9152 , \8816 , RIb553ff0_333);
and \U$8333 ( \9153 , RIb554248_338, \8812 );
nor \U$8334 ( \9154 , \9152 , \9153 );
and \U$8335 ( \9155 , \8835 , RIb554590_345);
and \U$8336 ( \9156 , RIb554518_344, \8800 );
nor \U$8337 ( \9157 , \9155 , \9156 );
and \U$8338 ( \9158 , \8806 , RIb5541d0_337);
and \U$8339 ( \9159 , RIb554158_336, \8829 );
nor \U$8340 ( \9160 , \9158 , \9159 );
nand \U$8341 ( \9161 , \9151 , \9154 , \9157 , \9160 );
and \U$8342 ( \9162 , \8859 , RIb5546f8_348);
and \U$8343 ( \9163 , RIb5544a0_343, \8823 );
nor \U$8344 ( \9164 , \9162 , \9163 );
not \U$8345 ( \9165 , \9164 );
nor \U$8346 ( \9166 , \9148 , \9161 , \9165 );
and \U$8347 ( \9167 , \8850 , RIb554338_340);
and \U$8348 ( \9168 , RIb5542c0_339, \8847 );
nor \U$8349 ( \9169 , \9167 , \9168 );
and \U$8350 ( \9170 , \8831 , RIb5540e0_335);
and \U$8351 ( \9171 , RIb554068_334, \8853 );
nor \U$8352 ( \9172 , \9170 , \9171 );
and \U$8353 ( \9173 , \8856 , RIb554770_349);
and \U$8354 ( \9174 , RIb5543b0_341, \8818 );
nor \U$8355 ( \9175 , \9173 , \9174 );
nand \U$8356 ( \9176 , \9166 , \9169 , \9172 , \9175 );
_DC r2f04 ( \9177_nR2f04 , \9176 , \8863 );
nand \U$8357 ( \9178 , \9177_nR2f04 , \8768 );
and \U$8358 ( \9179 , \9063_nR3133 , \8921 );
or \U$8359 ( \9180 , \8877 , \9122_nR301c );
nand \U$8360 ( \9181 , \9180 , \8917 );
nand \U$8361 ( \9182 , \9063_nR3133 , \8912 );
and \U$8362 ( \9183 , \9181 , \9182 );
and \U$8363 ( \9184 , \9122_nR301c , \8914 );
nor \U$8364 ( \9185 , \9179 , \9183 , \9184 );
or \U$8365 ( \9186 , \9178 , \9185 );
nand \U$8366 ( \9187 , \9147 , \9186 );
nand \U$8367 ( \9188 , \9129 , \9187 );
not \U$8368 ( \9189 , \9188 );
or \U$8369 ( \9190 , \9079 , \9072 );
nand \U$8370 ( \9191 , \9190 , \9080 );
nand \U$8371 ( \9192 , \9189 , \9191 );
xor \U$8372 ( \9193 , \9080 , \9081 );
not \U$8373 ( \9194 , \9073 );
nor \U$8374 ( \9195 , \9194 , \9075 );
nor \U$8375 ( \9196 , \9193 , \9195 );
or \U$8376 ( \9197 , \9192 , \9196 );
nand \U$8377 ( \9198 , \9195 , \9193 );
nand \U$8378 ( \9199 , \9197 , \9198 );
xor \U$8379 ( \9200 , \9082 , \9083 );
and \U$8380 ( \9201 , \9199 , \9200 );
not \U$8381 ( \9202 , \9199 );
not \U$8382 ( \9203 , \9200 );
and \U$8383 ( \9204 , \9202 , \9203 );
not \U$8384 ( \9205 , \9188 );
not \U$8385 ( \9206 , \9191 );
or \U$8386 ( \9207 , \9205 , \9206 );
or \U$8387 ( \9208 , \9191 , \9188 );
nand \U$8388 ( \9209 , \9207 , \9208 );
not \U$8389 ( \9210 , \9209 );
not \U$8390 ( \9211 , \9124 );
nor \U$8391 ( \9212 , \9211 , \9091 );
not \U$8392 ( \9213 , \9212 );
and \U$8393 ( \9214 , \9210 , \9213 );
and \U$8394 ( \9215 , \9209 , \9212 );
nor \U$8395 ( \9216 , \9214 , \9215 );
not \U$8396 ( \9217 , \9216 );
nand \U$8397 ( \9218 , \8907_nR3482 , \9139 );
or \U$8398 ( \9219 , \9030 , \8864_nR335c );
nand \U$8399 ( \9220 , \9219 , \9144 );
and \U$8400 ( \9221 , \9218 , \9220 );
and \U$8401 ( \9222 , \9141 , \8864_nR335c );
not \U$8402 ( \9223 , \9139 );
nor \U$8403 ( \9224 , \9031 , \9223 );
and \U$8404 ( \9225 , \8907_nR3482 , \9224 );
nor \U$8405 ( \9226 , \9221 , \9222 , \9225 );
and \U$8406 ( \9227 , \9063_nR3133 , \8981 );
or \U$8407 ( \9228 , \8935 , \8966_nR3254 );
nand \U$8408 ( \9229 , \9228 , \9018 );
nand \U$8409 ( \9230 , \9063_nR3133 , \8978 );
and \U$8410 ( \9231 , \9229 , \9230 );
and \U$8411 ( \9232 , \8966_nR3254 , \9022 );
nor \U$8412 ( \9233 , \9227 , \9231 , \9232 );
nand \U$8413 ( \9234 , \9226 , \9233 );
xor \U$8414 ( \9235 , \8495 , \8525_nR27ad );
xor \U$8415 ( \9236 , \9235 , \8744 );
xor \U$8416 ( \9237 , \8531 , \8561_nR2667 );
xor \U$8417 ( \9238 , \9237 , \8741 );
nor \U$8418 ( \9239 , \9236 , \9238 );
or \U$8419 ( \9240 , \9028 , \9239 );
and \U$8420 ( \9241 , \9234 , \9240 );
and \U$8421 ( \9242 , \8844 , RIb555670_381);
nand \U$8422 ( \9243 , RIb555760_383, \8856 );
and \U$8423 ( \9244 , \8818 , RIb5553a0_375);
and \U$8424 ( \9245 , RIb555418_376, \8825 );
nor \U$8425 ( \9246 , \9244 , \9245 );
nand \U$8426 ( \9247 , RIb555490_377, \8823 );
nand \U$8427 ( \9248 , \9243 , \9246 , \9247 );
and \U$8428 ( \9249 , \8816 , RIb554fe0_367);
and \U$8429 ( \9250 , RIb555508_378, \8800 );
nor \U$8430 ( \9251 , \9249 , \9250 );
and \U$8431 ( \9252 , \8835 , RIb555580_379);
and \U$8432 ( \9253 , RIb5555f8_380, \8839 );
nor \U$8433 ( \9254 , \9252 , \9253 );
nand \U$8434 ( \9255 , \9251 , \9254 );
nor \U$8435 ( \9256 , \9242 , \9248 , \9255 );
and \U$8436 ( \9257 , \8850 , RIb555328_374);
and \U$8437 ( \9258 , RIb5552b0_373, \8847 );
nor \U$8438 ( \9259 , \9257 , \9258 );
and \U$8439 ( \9260 , \8806 , RIb5551c0_371);
and \U$8440 ( \9261 , RIb555148_370, \8829 );
nor \U$8441 ( \9262 , \9260 , \9261 );
and \U$8442 ( \9263 , RIb5556e8_382, \8859 );
and \U$8443 ( \9264 , RIb555058_368, \8853 );
and \U$8444 ( \9265 , \8812 , RIb555238_372);
and \U$8445 ( \9266 , RIb5550d0_369, \8831 );
nor \U$8446 ( \9267 , \9265 , \9266 );
not \U$8447 ( \9268 , \9267 );
nor \U$8448 ( \9269 , \9263 , \9264 , \9268 );
nand \U$8449 ( \9270 , \9256 , \9259 , \9262 , \9269 );
_DC r2e0d ( \9271_nR2e0d , \9270 , \8863 );
not \U$8450 ( \9272 , \9271_nR2e0d );
nor \U$8451 ( \9273 , \8769 , \9272 );
not \U$8452 ( \9274 , \9273 );
and \U$8453 ( \9275 , \9122_nR301c , \8921 );
or \U$8454 ( \9276 , \8877 , \9177_nR2f04 );
nand \U$8455 ( \9277 , \9276 , \8917 );
nand \U$8456 ( \9278 , \9122_nR301c , \8912 );
and \U$8457 ( \9279 , \9277 , \9278 );
and \U$8458 ( \9280 , \9177_nR2f04 , \8914 );
nor \U$8459 ( \9281 , \9275 , \9279 , \9280 );
nor \U$8460 ( \9282 , \9274 , \9281 );
nor \U$8461 ( \9283 , \9233 , \9226 );
nor \U$8462 ( \9284 , \9241 , \9282 , \9283 );
xnor \U$8463 ( \9285 , \9178 , \9185 );
not \U$8464 ( \9286 , \9285 );
xor \U$8465 ( \9287 , \9146 , \9136 );
not \U$8466 ( \9288 , \9287 );
and \U$8467 ( \9289 , \9286 , \9288 );
and \U$8468 ( \9290 , \9285 , \9287 );
nor \U$8469 ( \9291 , \9289 , \9290 );
nand \U$8470 ( \9292 , \9284 , \9291 );
not \U$8471 ( \9293 , \9224 );
or \U$8472 ( \9294 , \9293 , \8865 );
not \U$8473 ( \9295 , \9141 );
or \U$8474 ( \9296 , \8967 , \9295 );
or \U$8475 ( \9297 , \9223 , \8865 );
or \U$8476 ( \9298 , \9030 , \8966_nR3254 );
nand \U$8477 ( \9299 , \9298 , \9144 );
nand \U$8478 ( \9300 , \9297 , \9299 );
nand \U$8479 ( \9301 , \9294 , \9296 , \9300 );
not \U$8480 ( \9302 , \9301 );
not \U$8481 ( \9303 , \9240 );
not \U$8482 ( \9304 , \9236 );
not \U$8483 ( \9305 , \9028 );
or \U$8484 ( \9306 , \9304 , \9305 );
or \U$8485 ( \9307 , \9028 , \9236 );
nand \U$8486 ( \9308 , \9306 , \9307 );
xor \U$8487 ( \9309 , \9238 , \9236 );
nor \U$8488 ( \9310 , \9308 , \9309 );
not \U$8489 ( \9311 , \9310 );
nor \U$8490 ( \9312 , \9303 , \9311 );
and \U$8491 ( \9313 , \9312 , \8907_nR3482 );
and \U$8492 ( \9314 , \9310 , \8907_nR3482 );
nor \U$8493 ( \9315 , \9314 , \9240 );
nor \U$8494 ( \9316 , \9313 , \9315 );
nor \U$8495 ( \9317 , \9302 , \9316 );
and \U$8496 ( \9318 , \9122_nR301c , \8981 );
or \U$8497 ( \9319 , \8935 , \9063_nR3133 );
nand \U$8498 ( \9320 , \9319 , \9018 );
nand \U$8499 ( \9321 , \9122_nR301c , \8978 );
and \U$8500 ( \9322 , \9320 , \9321 );
and \U$8501 ( \9323 , \9063_nR3133 , \9022 );
nor \U$8502 ( \9324 , \9318 , \9322 , \9323 );
and \U$8503 ( \9325 , \8844 , RIb554e78_364);
nand \U$8504 ( \9326 , RIb554f68_366, \8856 );
and \U$8505 ( \9327 , \8823 , RIb554c98_360);
and \U$8506 ( \9328 , RIb554c20_359, \8825 );
nor \U$8507 ( \9329 , \9327 , \9328 );
nand \U$8508 ( \9330 , RIb554d10_361, \8800 );
nand \U$8509 ( \9331 , \9326 , \9329 , \9330 );
and \U$8510 ( \9332 , \8816 , RIb5547e8_350);
and \U$8511 ( \9333 , RIb554a40_355, \8812 );
nor \U$8512 ( \9334 , \9332 , \9333 );
and \U$8513 ( \9335 , \8835 , RIb554d88_362);
and \U$8514 ( \9336 , RIb554e00_363, \8839 );
nor \U$8515 ( \9337 , \9335 , \9336 );
nand \U$8516 ( \9338 , \9334 , \9337 );
nor \U$8517 ( \9339 , \9325 , \9331 , \9338 );
and \U$8518 ( \9340 , \8818 , RIb554ba8_358);
and \U$8519 ( \9341 , RIb554b30_357, \8850 );
nor \U$8520 ( \9342 , \9340 , \9341 );
and \U$8521 ( \9343 , \8806 , RIb5549c8_354);
and \U$8522 ( \9344 , RIb554950_353, \8829 );
nor \U$8523 ( \9345 , \9343 , \9344 );
and \U$8524 ( \9346 , RIb554ef0_365, \8859 );
and \U$8525 ( \9347 , RIb554860_351, \8853 );
and \U$8526 ( \9348 , \8847 , RIb554ab8_356);
and \U$8527 ( \9349 , RIb5548d8_352, \8831 );
nor \U$8528 ( \9350 , \9348 , \9349 );
not \U$8529 ( \9351 , \9350 );
nor \U$8530 ( \9352 , \9346 , \9347 , \9351 );
nand \U$8531 ( \9353 , \9339 , \9342 , \9345 , \9352 );
_DC r2cff ( \9354_nR2cff , \9353 , \8863 );
nand \U$8532 ( \9355 , \9354_nR2cff , \8768 );
and \U$8533 ( \9356 , \9324 , \9355 );
and \U$8534 ( \9357 , \9177_nR2f04 , \8921 );
or \U$8535 ( \9358 , \8877 , \9271_nR2e0d );
nand \U$8536 ( \9359 , \9358 , \8917 );
nand \U$8537 ( \9360 , \9177_nR2f04 , \8912 );
and \U$8538 ( \9361 , \9359 , \9360 );
and \U$8539 ( \9362 , \9271_nR2e0d , \8914 );
nor \U$8540 ( \9363 , \9357 , \9361 , \9362 );
nor \U$8541 ( \9364 , \9356 , \9363 );
and \U$8542 ( \9365 , \9317 , \9364 );
not \U$8543 ( \9366 , \9240 );
not \U$8544 ( \9367 , \9283 );
nand \U$8545 ( \9368 , \9367 , \9234 );
not \U$8546 ( \9369 , \9368 );
or \U$8547 ( \9370 , \9366 , \9369 );
or \U$8548 ( \9371 , \9368 , \9240 );
nand \U$8549 ( \9372 , \9370 , \9371 );
not \U$8550 ( \9373 , \9372 );
not \U$8551 ( \9374 , \9281 );
not \U$8552 ( \9375 , \9273 );
and \U$8553 ( \9376 , \9374 , \9375 );
and \U$8554 ( \9377 , \9281 , \9273 );
nor \U$8555 ( \9378 , \9376 , \9377 );
nor \U$8556 ( \9379 , \9373 , \9378 );
and \U$8557 ( \9380 , \9365 , \9379 );
xor \U$8558 ( \9381 , \9292 , \9380 );
not \U$8559 ( \9382 , \9187 );
not \U$8560 ( \9383 , \9128 );
or \U$8561 ( \9384 , \9382 , \9383 );
or \U$8562 ( \9385 , \9128 , \9187 );
nand \U$8563 ( \9386 , \9384 , \9385 );
and \U$8564 ( \9387 , \9381 , \9386 );
and \U$8565 ( \9388 , \9292 , \9380 );
or \U$8566 ( \9389 , \9387 , \9388 );
not \U$8567 ( \9390 , \9389 );
and \U$8568 ( \9391 , \9217 , \9390 );
and \U$8569 ( \9392 , \9216 , \9389 );
nor \U$8570 ( \9393 , \9391 , \9392 );
nand \U$8571 ( \9394 , \8864_nR335c , \9310 );
or \U$8572 ( \9395 , \9240 , \8907_nR3482 );
or \U$8573 ( \9396 , \9240 , \9309 );
nand \U$8574 ( \9397 , \9395 , \9396 );
and \U$8575 ( \9398 , \9394 , \9397 );
and \U$8576 ( \9399 , \9240 , \9309 );
and \U$8577 ( \9400 , \9399 , \8907_nR3482 );
and \U$8578 ( \9401 , \8864_nR335c , \9312 );
nor \U$8579 ( \9402 , \9398 , \9400 , \9401 );
not \U$8580 ( \9403 , \9402 );
xor \U$8581 ( \9404 , \8603 , \8633_nR2589 );
xor \U$8582 ( \9405 , \9404 , \8735 );
not \U$8583 ( \9406 , \9405 );
xor \U$8584 ( \9407 , \8567 , \8597_nR2665 );
xor \U$8585 ( \9408 , \9407 , \8738 );
not \U$8586 ( \9409 , \9408 );
and \U$8587 ( \9410 , \9406 , \9409 );
or \U$8588 ( \9411 , \9238 , \9410 );
not \U$8589 ( \9412 , \9411 );
not \U$8590 ( \9413 , \9412 );
and \U$8591 ( \9414 , \9403 , \9413 );
and \U$8592 ( \9415 , \9402 , \9412 );
nand \U$8593 ( \9416 , \8966_nR3254 , \9139 );
or \U$8594 ( \9417 , \9030 , \9063_nR3133 );
nand \U$8595 ( \9418 , \9417 , \9144 );
and \U$8596 ( \9419 , \9416 , \9418 );
and \U$8597 ( \9420 , \9141 , \9063_nR3133 );
and \U$8598 ( \9421 , \8966_nR3254 , \9224 );
nor \U$8599 ( \9422 , \9419 , \9420 , \9421 );
nor \U$8600 ( \9423 , \9415 , \9422 );
nor \U$8601 ( \9424 , \9414 , \9423 );
not \U$8602 ( \9425 , \9424 );
and \U$8603 ( \9426 , \9177_nR2f04 , \8981 );
or \U$8604 ( \9427 , \8935 , \9122_nR301c );
nand \U$8605 ( \9428 , \9427 , \9018 );
nand \U$8606 ( \9429 , \9177_nR2f04 , \8978 );
and \U$8607 ( \9430 , \9428 , \9429 );
and \U$8608 ( \9431 , \9122_nR301c , \9022 );
nor \U$8609 ( \9432 , \9426 , \9430 , \9431 );
and \U$8610 ( \9433 , \8835 , RIb556570_413);
nand \U$8611 ( \9434 , RIb556750_417, \8856 );
and \U$8612 ( \9435 , \8823 , RIb556480_411);
and \U$8613 ( \9436 , RIb5561b0_405, \8806 );
nor \U$8614 ( \9437 , \9435 , \9436 );
nand \U$8615 ( \9438 , RIb5564f8_412, \8800 );
nand \U$8616 ( \9439 , \9434 , \9437 , \9438 );
and \U$8617 ( \9440 , \8816 , RIb555fd0_401);
and \U$8618 ( \9441 , RIb5562a0_407, \8847 );
nor \U$8619 ( \9442 , \9440 , \9441 );
and \U$8620 ( \9443 , \8859 , RIb5566d8_416);
and \U$8621 ( \9444 , RIb556660_415, \8844 );
nor \U$8622 ( \9445 , \9443 , \9444 );
nand \U$8623 ( \9446 , \9442 , \9445 );
nor \U$8624 ( \9447 , \9433 , \9439 , \9446 );
and \U$8625 ( \9448 , \8839 , RIb5565e8_414);
and \U$8626 ( \9449 , RIb556048_402, \8853 );
nor \U$8627 ( \9450 , \9448 , \9449 );
and \U$8628 ( \9451 , \8850 , RIb556318_408);
and \U$8629 ( \9452 , RIb5560c0_403, \8831 );
nor \U$8630 ( \9453 , \9451 , \9452 );
and \U$8631 ( \9454 , RIb556228_406, \8812 );
and \U$8632 ( \9455 , RIb556138_404, \8829 );
and \U$8633 ( \9456 , \8818 , RIb556390_409);
and \U$8634 ( \9457 , RIb556408_410, \8825 );
nor \U$8635 ( \9458 , \9456 , \9457 );
not \U$8636 ( \9459 , \9458 );
nor \U$8637 ( \9460 , \9454 , \9455 , \9459 );
nand \U$8638 ( \9461 , \9447 , \9450 , \9453 , \9460 );
_DC r2c1e ( \9462_nR2c1e , \9461 , \8863 );
nand \U$8639 ( \9463 , \9462_nR2c1e , \8768 );
and \U$8640 ( \9464 , \9432 , \9463 );
and \U$8641 ( \9465 , \9271_nR2e0d , \8921 );
or \U$8642 ( \9466 , \8877 , \9354_nR2cff );
nand \U$8643 ( \9467 , \9466 , \8917 );
nand \U$8644 ( \9468 , \9271_nR2e0d , \8912 );
and \U$8645 ( \9469 , \9467 , \9468 );
and \U$8646 ( \9470 , \9354_nR2cff , \8914 );
nor \U$8647 ( \9471 , \9465 , \9469 , \9470 );
nor \U$8648 ( \9472 , \9464 , \9471 );
nand \U$8649 ( \9473 , \9425 , \9472 );
not \U$8650 ( \9474 , \9473 );
not \U$8651 ( \9475 , \9355 );
not \U$8652 ( \9476 , \9363 );
not \U$8653 ( \9477 , \9324 );
and \U$8654 ( \9478 , \9476 , \9477 );
and \U$8655 ( \9479 , \9363 , \9324 );
nor \U$8656 ( \9480 , \9478 , \9479 );
not \U$8657 ( \9481 , \9480 );
or \U$8658 ( \9482 , \9475 , \9481 );
or \U$8659 ( \9483 , \9480 , \9355 );
nand \U$8660 ( \9484 , \9482 , \9483 );
not \U$8661 ( \9485 , \9484 );
not \U$8662 ( \9486 , \9301 );
not \U$8663 ( \9487 , \9316 );
and \U$8664 ( \9488 , \9486 , \9487 );
and \U$8665 ( \9489 , \9301 , \9316 );
nor \U$8666 ( \9490 , \9488 , \9489 );
nor \U$8667 ( \9491 , \9485 , \9490 );
nand \U$8668 ( \9492 , \9474 , \9491 );
not \U$8669 ( \9493 , \9378 );
not \U$8670 ( \9494 , \9372 );
and \U$8671 ( \9495 , \9493 , \9494 );
and \U$8672 ( \9496 , \9378 , \9372 );
nor \U$8673 ( \9497 , \9495 , \9496 );
not \U$8674 ( \9498 , \9497 );
xor \U$8675 ( \9499 , \9317 , \9364 );
nand \U$8676 ( \9500 , \9498 , \9499 );
and \U$8677 ( \9501 , \9492 , \9500 );
not \U$8678 ( \9502 , \9291 );
not \U$8679 ( \9503 , \9284 );
and \U$8680 ( \9504 , \9502 , \9503 );
not \U$8681 ( \9505 , \9292 );
nor \U$8682 ( \9506 , \9504 , \9505 );
nor \U$8683 ( \9507 , \9501 , \9506 );
not \U$8684 ( \9508 , \9287 );
nor \U$8685 ( \9509 , \9508 , \9285 );
xor \U$8686 ( \9510 , \9507 , \9509 );
xor \U$8687 ( \9511 , \9292 , \9380 );
xor \U$8688 ( \9512 , \9511 , \9386 );
and \U$8689 ( \9513 , \9510 , \9512 );
and \U$8690 ( \9514 , \9507 , \9509 );
or \U$8691 ( \9515 , \9513 , \9514 );
xor \U$8692 ( \9516 , \9393 , \9515 );
xor \U$8693 ( \9517 , \9507 , \9509 );
xor \U$8694 ( \9518 , \9517 , \9512 );
not \U$8695 ( \9519 , \9472 );
not \U$8696 ( \9520 , \9424 );
and \U$8697 ( \9521 , \9519 , \9520 );
and \U$8698 ( \9522 , \9472 , \9424 );
nor \U$8699 ( \9523 , \9521 , \9522 );
not \U$8700 ( \9524 , \9484 );
not \U$8701 ( \9525 , \9490 );
and \U$8702 ( \9526 , \9524 , \9525 );
and \U$8703 ( \9527 , \9484 , \9490 );
nor \U$8704 ( \9528 , \9526 , \9527 );
nand \U$8705 ( \9529 , \9523 , \9528 );
not \U$8706 ( \9530 , \9499 );
not \U$8707 ( \9531 , \9497 );
or \U$8708 ( \9532 , \9530 , \9531 );
or \U$8709 ( \9533 , \9497 , \9499 );
nand \U$8710 ( \9534 , \9532 , \9533 );
xor \U$8711 ( \9535 , \9529 , \9534 );
not \U$8712 ( \9536 , \9408 );
not \U$8713 ( \9537 , \9238 );
or \U$8714 ( \9538 , \9536 , \9537 );
or \U$8715 ( \9539 , \9238 , \9408 );
nand \U$8716 ( \9540 , \9538 , \9539 );
xor \U$8717 ( \9541 , \9406 , \9409 );
nor \U$8718 ( \9542 , \9540 , \9541 );
not \U$8719 ( \9543 , \9542 );
nor \U$8720 ( \9544 , \9543 , \9412 );
not \U$8721 ( \9545 , \9544 );
or \U$8722 ( \9546 , \9545 , \8909 );
or \U$8723 ( \9547 , \9543 , \8909 );
nand \U$8724 ( \9548 , \9547 , \9412 );
nand \U$8725 ( \9549 , \9546 , \9548 );
not \U$8726 ( \9550 , \9312 );
or \U$8727 ( \9551 , \9550 , \8967 );
not \U$8728 ( \9552 , \9399 );
or \U$8729 ( \9553 , \8865 , \9552 );
or \U$8730 ( \9554 , \9311 , \8967 );
or \U$8731 ( \9555 , \9240 , \8864_nR335c );
nand \U$8732 ( \9556 , \9555 , \9396 );
nand \U$8733 ( \9557 , \9554 , \9556 );
nand \U$8734 ( \9558 , \9551 , \9553 , \9557 );
and \U$8735 ( \9559 , \9549 , \9558 );
and \U$8736 ( \9560 , \9271_nR2e0d , \8981 );
or \U$8737 ( \9561 , \8935 , \9177_nR2f04 );
nand \U$8738 ( \9562 , \9561 , \9018 );
nand \U$8739 ( \9563 , \9271_nR2e0d , \8978 );
and \U$8740 ( \9564 , \9562 , \9563 );
and \U$8741 ( \9565 , \9177_nR2f04 , \9022 );
nor \U$8742 ( \9566 , \9560 , \9564 , \9565 );
nand \U$8743 ( \9567 , \9063_nR3133 , \9139 );
or \U$8744 ( \9568 , \9030 , \9122_nR301c );
nand \U$8745 ( \9569 , \9568 , \9144 );
and \U$8746 ( \9570 , \9567 , \9569 );
and \U$8747 ( \9571 , \9141 , \9122_nR301c );
and \U$8748 ( \9572 , \9063_nR3133 , \9224 );
nor \U$8749 ( \9573 , \9570 , \9571 , \9572 );
xor \U$8750 ( \9574 , \9566 , \9573 );
and \U$8751 ( \9575 , \9354_nR2cff , \8921 );
or \U$8752 ( \9576 , \8877 , \9462_nR2c1e );
nand \U$8753 ( \9577 , \9576 , \8917 );
nand \U$8754 ( \9578 , \9354_nR2cff , \8912 );
and \U$8755 ( \9579 , \9577 , \9578 );
and \U$8756 ( \9580 , \9462_nR2c1e , \8914 );
nor \U$8757 ( \9581 , \9575 , \9579 , \9580 );
and \U$8758 ( \9582 , \9574 , \9581 );
and \U$8759 ( \9583 , \9566 , \9573 );
or \U$8760 ( \9584 , \9582 , \9583 );
not \U$8761 ( \9585 , \9584 );
and \U$8762 ( \9586 , \9559 , \9585 );
not \U$8763 ( \9587 , \9402 );
or \U$8764 ( \9588 , \9422 , \9411 );
nand \U$8765 ( \9589 , \9411 , \9422 );
nand \U$8766 ( \9590 , \9588 , \9589 );
not \U$8767 ( \9591 , \9590 );
or \U$8768 ( \9592 , \9587 , \9591 );
or \U$8769 ( \9593 , \9590 , \9402 );
nand \U$8770 ( \9594 , \9592 , \9593 );
not \U$8771 ( \9595 , \9463 );
not \U$8772 ( \9596 , \9471 );
not \U$8773 ( \9597 , \9432 );
and \U$8774 ( \9598 , \9596 , \9597 );
and \U$8775 ( \9599 , \9471 , \9432 );
nor \U$8776 ( \9600 , \9598 , \9599 );
not \U$8777 ( \9601 , \9600 );
or \U$8778 ( \9602 , \9595 , \9601 );
or \U$8779 ( \9603 , \9600 , \9463 );
nand \U$8780 ( \9604 , \9602 , \9603 );
and \U$8781 ( \9605 , \9594 , \9604 );
and \U$8782 ( \9606 , \9586 , \9605 );
and \U$8783 ( \9607 , \9535 , \9606 );
and \U$8784 ( \9608 , \9529 , \9534 );
or \U$8785 ( \9609 , \9607 , \9608 );
xor \U$8786 ( \9610 , \9365 , \9379 );
xor \U$8787 ( \9611 , \9609 , \9610 );
not \U$8788 ( \9612 , \9500 );
not \U$8789 ( \9613 , \9506 );
not \U$8790 ( \9614 , \9492 );
and \U$8791 ( \9615 , \9613 , \9614 );
and \U$8792 ( \9616 , \9506 , \9492 );
nor \U$8793 ( \9617 , \9615 , \9616 );
not \U$8794 ( \9618 , \9617 );
or \U$8795 ( \9619 , \9612 , \9618 );
or \U$8796 ( \9620 , \9617 , \9500 );
nand \U$8797 ( \9621 , \9619 , \9620 );
and \U$8798 ( \9622 , \9611 , \9621 );
and \U$8799 ( \9623 , \9609 , \9610 );
or \U$8800 ( \9624 , \9622 , \9623 );
xor \U$8801 ( \9625 , \9518 , \9624 );
not \U$8802 ( \9626 , \9473 );
not \U$8803 ( \9627 , \9491 );
or \U$8804 ( \9628 , \9626 , \9627 );
or \U$8805 ( \9629 , \9491 , \9473 );
nand \U$8806 ( \9630 , \9628 , \9629 );
xor \U$8807 ( \9631 , \9529 , \9534 );
xor \U$8808 ( \9632 , \9631 , \9606 );
and \U$8809 ( \9633 , \9630 , \9632 );
xor \U$8810 ( \9634 , \9559 , \9585 );
xor \U$8811 ( \9635 , \9594 , \9604 );
and \U$8812 ( \9636 , \9634 , \9635 );
xor \U$8813 ( \9637 , \9549 , \9558 );
not \U$8814 ( \9638 , \9637 );
xor \U$8815 ( \9639 , \9566 , \9573 );
xor \U$8816 ( \9640 , \9639 , \9581 );
nor \U$8817 ( \9641 , \9638 , \9640 );
and \U$8818 ( \9642 , \9354_nR2cff , \8981 );
or \U$8819 ( \9643 , \8935 , \9271_nR2e0d );
nand \U$8820 ( \9644 , \9643 , \9018 );
nand \U$8821 ( \9645 , \9354_nR2cff , \8978 );
and \U$8822 ( \9646 , \9644 , \9645 );
and \U$8823 ( \9647 , \9271_nR2e0d , \9022 );
nor \U$8824 ( \9648 , \9642 , \9646 , \9647 );
nand \U$8825 ( \9649 , \9122_nR301c , \9139 );
or \U$8826 ( \9650 , \9030 , \9177_nR2f04 );
nand \U$8827 ( \9651 , \9650 , \9144 );
and \U$8828 ( \9652 , \9649 , \9651 );
and \U$8829 ( \9653 , \9141 , \9177_nR2f04 );
and \U$8830 ( \9654 , \9122_nR301c , \9224 );
nor \U$8831 ( \9655 , \9652 , \9653 , \9654 );
xor \U$8832 ( \9656 , \9648 , \9655 );
and \U$8833 ( \9657 , \9462_nR2c1e , \8921 );
and \U$8834 ( \9658 , \8806 , RIb5559b8_388);
nand \U$8835 ( \9659 , RIb555f58_400, \8856 );
and \U$8836 ( \9660 , \8823 , RIb555c88_394);
and \U$8837 ( \9661 , RIb555940_387, \8829 );
nor \U$8838 ( \9662 , \9660 , \9661 );
nand \U$8839 ( \9663 , RIb555d00_395, \8800 );
nand \U$8840 ( \9664 , \9659 , \9662 , \9663 );
and \U$8841 ( \9665 , \8835 , RIb555d78_396);
and \U$8842 ( \9666 , RIb555df0_397, \8839 );
nor \U$8843 ( \9667 , \9665 , \9666 );
and \U$8844 ( \9668 , \8859 , RIb555ee0_399);
and \U$8845 ( \9669 , RIb555e68_398, \8844 );
nor \U$8846 ( \9670 , \9668 , \9669 );
nand \U$8847 ( \9671 , \9667 , \9670 );
nor \U$8848 ( \9672 , \9658 , \9664 , \9671 );
and \U$8849 ( \9673 , \8816 , RIb5557d8_384);
and \U$8850 ( \9674 , RIb555aa8_390, \8847 );
nor \U$8851 ( \9675 , \9673 , \9674 );
and \U$8852 ( \9676 , \8818 , RIb555b98_392);
and \U$8853 ( \9677 , RIb555c10_393, \8825 );
nor \U$8854 ( \9678 , \9676 , \9677 );
and \U$8855 ( \9679 , RIb555a30_389, \8812 );
and \U$8856 ( \9680 , RIb555850_385, \8853 );
and \U$8857 ( \9681 , \8850 , RIb555b20_391);
and \U$8858 ( \9682 , RIb5558c8_386, \8831 );
nor \U$8859 ( \9683 , \9681 , \9682 );
not \U$8860 ( \9684 , \9683 );
nor \U$8861 ( \9685 , \9679 , \9680 , \9684 );
nand \U$8862 ( \9686 , \9672 , \9675 , \9678 , \9685 );
_DC r2b14 ( \9687_nR2b14 , \9686 , \8863 );
or \U$8863 ( \9688 , \8877 , \9687_nR2b14 );
nand \U$8864 ( \9689 , \9688 , \8917 );
nand \U$8865 ( \9690 , \9462_nR2c1e , \8912 );
and \U$8866 ( \9691 , \9689 , \9690 );
and \U$8867 ( \9692 , \9687_nR2b14 , \8914 );
nor \U$8868 ( \9693 , \9657 , \9691 , \9692 );
and \U$8869 ( \9694 , \9656 , \9693 );
and \U$8870 ( \9695 , \9648 , \9655 );
or \U$8871 ( \9696 , \9694 , \9695 );
nand \U$8872 ( \9697 , \8864_nR335c , \9542 );
or \U$8873 ( \9698 , \9411 , \8907_nR3482 );
or \U$8874 ( \9699 , \9411 , \9541 );
nand \U$8875 ( \9700 , \9698 , \9699 );
and \U$8876 ( \9701 , \9697 , \9700 );
and \U$8877 ( \9702 , \9411 , \9541 );
and \U$8878 ( \9703 , \9702 , \8907_nR3482 );
and \U$8879 ( \9704 , \8864_nR335c , \9544 );
nor \U$8880 ( \9705 , \9701 , \9703 , \9704 );
not \U$8881 ( \9706 , \8698 );
not \U$8882 ( \9707 , \8731 );
nand \U$8883 ( \9708 , \9707 , \8729 );
not \U$8884 ( \9709 , \9708 );
or \U$8885 ( \9710 , \9706 , \9709 );
or \U$8886 ( \9711 , \9708 , \8698 );
nand \U$8887 ( \9712 , \9710 , \9711 );
xor \U$8888 ( \9713 , \8635 , \8665_nR258b );
xor \U$8889 ( \9714 , \9713 , \8732 );
not \U$8890 ( \9715 , \9714 );
and \U$8891 ( \9716 , \9712 , \9715 );
or \U$8892 ( \9717 , \9405 , \9716 );
not \U$8893 ( \9718 , \9717 );
xor \U$8894 ( \9719 , \9705 , \9718 );
nand \U$8895 ( \9720 , \9063_nR3133 , \9310 );
or \U$8896 ( \9721 , \9240 , \8966_nR3254 );
nand \U$8897 ( \9722 , \9721 , \9396 );
and \U$8898 ( \9723 , \9720 , \9722 );
and \U$8899 ( \9724 , \9399 , \8966_nR3254 );
and \U$8900 ( \9725 , \9063_nR3133 , \9312 );
nor \U$8901 ( \9726 , \9723 , \9724 , \9725 );
and \U$8902 ( \9727 , \9719 , \9726 );
and \U$8903 ( \9728 , \9705 , \9718 );
or \U$8904 ( \9729 , \9727 , \9728 );
nor \U$8905 ( \9730 , \9696 , \9729 );
and \U$8906 ( \9731 , \9641 , \9730 );
xor \U$8907 ( \9732 , \9636 , \9731 );
or \U$8908 ( \9733 , \9528 , \9523 );
nand \U$8909 ( \9734 , \9733 , \9529 );
and \U$8910 ( \9735 , \9732 , \9734 );
and \U$8911 ( \9736 , \9636 , \9731 );
or \U$8912 ( \9737 , \9735 , \9736 );
xor \U$8913 ( \9738 , \9529 , \9534 );
xor \U$8914 ( \9739 , \9738 , \9606 );
and \U$8915 ( \9740 , \9737 , \9739 );
and \U$8916 ( \9741 , \9630 , \9737 );
or \U$8917 ( \9742 , \9633 , \9740 , \9741 );
xor \U$8918 ( \9743 , \9609 , \9610 );
xor \U$8919 ( \9744 , \9743 , \9621 );
xor \U$8920 ( \9745 , \9742 , \9744 );
xor \U$8921 ( \9746 , \9529 , \9534 );
xor \U$8922 ( \9747 , \9746 , \9606 );
xor \U$8923 ( \9748 , \9630 , \9737 );
xor \U$8924 ( \9749 , \9747 , \9748 );
not \U$8925 ( \9750 , \9640 );
not \U$8926 ( \9751 , \9637 );
and \U$8927 ( \9752 , \9750 , \9751 );
and \U$8928 ( \9753 , \9640 , \9637 );
nor \U$8929 ( \9754 , \9752 , \9753 );
not \U$8930 ( \9755 , \9687_nR2b14 );
nor \U$8931 ( \9756 , \8769 , \9755 );
or \U$8932 ( \9757 , \9754 , \9756 );
xnor \U$8933 ( \9758 , \9729 , \9696 );
nand \U$8934 ( \9759 , \9757 , \9758 );
or \U$8935 ( \9760 , \9405 , \9714 );
nand \U$8936 ( \9761 , \9714 , \9405 );
nand \U$8937 ( \9762 , \9760 , \9761 );
xor \U$8938 ( \9763 , \9712 , \9715 );
nor \U$8939 ( \9764 , \9762 , \9763 );
not \U$8940 ( \9765 , \9764 );
nor \U$8941 ( \9766 , \9765 , \9718 );
not \U$8942 ( \9767 , \9766 );
or \U$8943 ( \9768 , \9767 , \8909 );
or \U$8944 ( \9769 , \9765 , \8909 );
nand \U$8945 ( \9770 , \9769 , \9718 );
nand \U$8946 ( \9771 , \9768 , \9770 );
not \U$8947 ( \9772 , \9771 );
nand \U$8948 ( \9773 , \8966_nR3254 , \9542 );
or \U$8949 ( \9774 , \9411 , \8864_nR335c );
nand \U$8950 ( \9775 , \9774 , \9699 );
and \U$8951 ( \9776 , \9773 , \9775 );
and \U$8952 ( \9777 , \9702 , \8864_nR335c );
and \U$8953 ( \9778 , \8966_nR3254 , \9544 );
nor \U$8954 ( \9779 , \9776 , \9777 , \9778 );
nor \U$8955 ( \9780 , \9772 , \9779 );
not \U$8956 ( \9781 , \9780 );
nand \U$8957 ( \9782 , \9177_nR2f04 , \9139 );
or \U$8958 ( \9783 , \9030 , \9271_nR2e0d );
nand \U$8959 ( \9784 , \9783 , \9144 );
and \U$8960 ( \9785 , \9782 , \9784 );
and \U$8961 ( \9786 , \9141 , \9271_nR2e0d );
and \U$8962 ( \9787 , \9177_nR2f04 , \9224 );
nor \U$8963 ( \9788 , \9785 , \9786 , \9787 );
nand \U$8964 ( \9789 , \9122_nR301c , \9310 );
or \U$8965 ( \9790 , \9240 , \9063_nR3133 );
nand \U$8966 ( \9791 , \9790 , \9396 );
and \U$8967 ( \9792 , \9789 , \9791 );
and \U$8968 ( \9793 , \9399 , \9063_nR3133 );
and \U$8969 ( \9794 , \9122_nR301c , \9312 );
nor \U$8970 ( \9795 , \9792 , \9793 , \9794 );
xor \U$8971 ( \9796 , \9788 , \9795 );
and \U$8972 ( \9797 , \9462_nR2c1e , \8981 );
or \U$8973 ( \9798 , \8935 , \9354_nR2cff );
nand \U$8974 ( \9799 , \9798 , \9018 );
nand \U$8975 ( \9800 , \9462_nR2c1e , \8978 );
and \U$8976 ( \9801 , \9799 , \9800 );
and \U$8977 ( \9802 , \9354_nR2cff , \9022 );
nor \U$8978 ( \9803 , \9797 , \9801 , \9802 );
and \U$8979 ( \9804 , \9796 , \9803 );
and \U$8980 ( \9805 , \9788 , \9795 );
or \U$8981 ( \9806 , \9804 , \9805 );
nor \U$8982 ( \9807 , \9781 , \9806 );
xor \U$8983 ( \9808 , \9648 , \9655 );
xor \U$8984 ( \9809 , \9808 , \9693 );
xor \U$8985 ( \9810 , \9705 , \9718 );
xor \U$8986 ( \9811 , \9810 , \9726 );
nor \U$8987 ( \9812 , \9809 , \9811 );
not \U$8988 ( \9813 , \9812 );
and \U$8989 ( \9814 , \8818 , RIb557380_443);
and \U$8990 ( \9815 , \8859 , RIb5576c8_450);
and \U$8991 ( \9816 , RIb557650_449, \8844 );
nor \U$8992 ( \9817 , \9815 , \9816 );
and \U$8993 ( \9818 , \8806 , RIb5571a0_439);
and \U$8994 ( \9819 , RIb557128_438, \8829 );
nor \U$8995 ( \9820 , \9818 , \9819 );
and \U$8996 ( \9821 , \8816 , RIb556fc0_435);
and \U$8997 ( \9822 , RIb557308_442, \8850 );
nor \U$8998 ( \9823 , \9821 , \9822 );
and \U$8999 ( \9824 , \8835 , RIb557560_447);
and \U$9000 ( \9825 , RIb5575d8_448, \8839 );
nor \U$9001 ( \9826 , \9824 , \9825 );
nand \U$9002 ( \9827 , \9817 , \9820 , \9823 , \9826 );
and \U$9003 ( \9828 , \8823 , RIb557470_445);
and \U$9004 ( \9829 , RIb5573f8_444, \8825 );
nor \U$9005 ( \9830 , \9828 , \9829 );
not \U$9006 ( \9831 , \9830 );
nor \U$9007 ( \9832 , \9814 , \9827 , \9831 );
and \U$9008 ( \9833 , \8847 , RIb557290_441);
and \U$9009 ( \9834 , RIb557218_440, \8812 );
nor \U$9010 ( \9835 , \9833 , \9834 );
and \U$9011 ( \9836 , \8831 , RIb5570b0_437);
and \U$9012 ( \9837 , RIb557038_436, \8853 );
nor \U$9013 ( \9838 , \9836 , \9837 );
and \U$9014 ( \9839 , \8856 , RIb557740_451);
and \U$9015 ( \9840 , RIb5574e8_446, \8800 );
nor \U$9016 ( \9841 , \9839 , \9840 );
nand \U$9017 ( \9842 , \9832 , \9835 , \9838 , \9841 );
_DC r2a34 ( \9843_nR2a34 , \9842 , \8863 );
nand \U$9018 ( \9844 , \9843_nR2a34 , \8768 );
nand \U$9019 ( \9845 , \9813 , \9844 );
and \U$9020 ( \9846 , \9807 , \9845 );
xor \U$9021 ( \9847 , \9759 , \9846 );
xor \U$9022 ( \9848 , \9634 , \9635 );
and \U$9023 ( \9849 , \9847 , \9848 );
and \U$9024 ( \9850 , \9759 , \9846 );
or \U$9025 ( \9851 , \9849 , \9850 );
xor \U$9026 ( \9852 , \9586 , \9605 );
xor \U$9027 ( \9853 , \9851 , \9852 );
xor \U$9028 ( \9854 , \9636 , \9731 );
xor \U$9029 ( \9855 , \9854 , \9734 );
and \U$9030 ( \9856 , \9853 , \9855 );
and \U$9031 ( \9857 , \9851 , \9852 );
or \U$9032 ( \9858 , \9856 , \9857 );
xor \U$9033 ( \9859 , \9749 , \9858 );
nor \U$9034 ( \9860 , \9730 , \9756 );
not \U$9035 ( \9861 , \9860 );
not \U$9036 ( \9862 , \9641 );
or \U$9037 ( \9863 , \9861 , \9862 );
or \U$9038 ( \9864 , \9641 , \9860 );
nand \U$9039 ( \9865 , \9863 , \9864 );
xor \U$9040 ( \9866 , \9759 , \9846 );
xor \U$9041 ( \9867 , \9866 , \9848 );
and \U$9042 ( \9868 , \9865 , \9867 );
or \U$9043 ( \9869 , \9806 , \9780 );
and \U$9044 ( \9870 , \8835 , RIb556d68_430);
nand \U$9045 ( \9871 , RIb556f48_434, \8856 );
and \U$9046 ( \9872 , \8818 , RIb556b88_426);
and \U$9047 ( \9873 , RIb556c00_427, \8825 );
nor \U$9048 ( \9874 , \9872 , \9873 );
nand \U$9049 ( \9875 , RIb556cf0_429, \8800 );
nand \U$9050 ( \9876 , \9871 , \9874 , \9875 );
and \U$9051 ( \9877 , \8816 , RIb5567c8_418);
and \U$9052 ( \9878 , RIb556c78_428, \8823 );
nor \U$9053 ( \9879 , \9877 , \9878 );
and \U$9054 ( \9880 , \8859 , RIb556ed0_433);
and \U$9055 ( \9881 , RIb556e58_432, \8844 );
nor \U$9056 ( \9882 , \9880 , \9881 );
nand \U$9057 ( \9883 , \9879 , \9882 );
nor \U$9058 ( \9884 , \9870 , \9876 , \9883 );
and \U$9059 ( \9885 , \8850 , RIb556b10_425);
and \U$9060 ( \9886 , RIb556a98_424, \8847 );
nor \U$9061 ( \9887 , \9885 , \9886 );
and \U$9062 ( \9888 , \8806 , RIb5569a8_422);
and \U$9063 ( \9889 , RIb556930_421, \8829 );
nor \U$9064 ( \9890 , \9888 , \9889 );
and \U$9065 ( \9891 , RIb556a20_423, \8812 );
and \U$9066 ( \9892 , RIb5568b8_420, \8831 );
and \U$9067 ( \9893 , \8839 , RIb556de0_431);
and \U$9068 ( \9894 , RIb556840_419, \8853 );
nor \U$9069 ( \9895 , \9893 , \9894 );
not \U$9070 ( \9896 , \9895 );
nor \U$9071 ( \9897 , \9891 , \9892 , \9896 );
nand \U$9072 ( \9898 , \9884 , \9887 , \9890 , \9897 );
_DC r2959 ( \9899_nR2959 , \9898 , \8863 );
nand \U$9073 ( \9900 , \9899_nR2959 , \8768 );
and \U$9074 ( \9901 , \9687_nR2b14 , \8921 );
or \U$9075 ( \9902 , \8877 , \9843_nR2a34 );
nand \U$9076 ( \9903 , \9902 , \8917 );
nand \U$9077 ( \9904 , \9687_nR2b14 , \8912 );
and \U$9078 ( \9905 , \9903 , \9904 );
and \U$9079 ( \9906 , \9843_nR2a34 , \8914 );
nor \U$9080 ( \9907 , \9901 , \9905 , \9906 );
or \U$9081 ( \9908 , \9900 , \9907 );
nand \U$9082 ( \9909 , \9780 , \9806 );
nand \U$9083 ( \9910 , \9869 , \9908 , \9909 );
not \U$9084 ( \9911 , \9844 );
and \U$9085 ( \9912 , \9809 , \9811 );
nor \U$9086 ( \9913 , \9912 , \9812 );
not \U$9087 ( \9914 , \9913 );
or \U$9088 ( \9915 , \9911 , \9914 );
or \U$9089 ( \9916 , \9913 , \9844 );
nand \U$9090 ( \9917 , \9915 , \9916 );
and \U$9091 ( \9918 , \9910 , \9917 );
nand \U$9092 ( \9919 , \9271_nR2e0d , \9139 );
or \U$9093 ( \9920 , \9030 , \9354_nR2cff );
nand \U$9094 ( \9921 , \9920 , \9144 );
and \U$9095 ( \9922 , \9919 , \9921 );
and \U$9096 ( \9923 , \9141 , \9354_nR2cff );
and \U$9097 ( \9924 , \9271_nR2e0d , \9224 );
nor \U$9098 ( \9925 , \9922 , \9923 , \9924 );
nand \U$9099 ( \9926 , \9177_nR2f04 , \9310 );
or \U$9100 ( \9927 , \9240 , \9122_nR301c );
nand \U$9101 ( \9928 , \9927 , \9396 );
and \U$9102 ( \9929 , \9926 , \9928 );
and \U$9103 ( \9930 , \9399 , \9122_nR301c );
and \U$9104 ( \9931 , \9177_nR2f04 , \9312 );
nor \U$9105 ( \9932 , \9929 , \9930 , \9931 );
xor \U$9106 ( \9933 , \9925 , \9932 );
and \U$9107 ( \9934 , \9687_nR2b14 , \8981 );
or \U$9108 ( \9935 , \8935 , \9462_nR2c1e );
nand \U$9109 ( \9936 , \9935 , \9018 );
nand \U$9110 ( \9937 , \9687_nR2b14 , \8978 );
and \U$9111 ( \9938 , \9936 , \9937 );
and \U$9112 ( \9939 , \9462_nR2c1e , \9022 );
nor \U$9113 ( \9940 , \9934 , \9938 , \9939 );
and \U$9114 ( \9941 , \9933 , \9940 );
and \U$9115 ( \9942 , \9925 , \9932 );
or \U$9116 ( \9943 , \9941 , \9942 );
nand \U$9117 ( \9944 , \8864_nR335c , \9764 );
or \U$9118 ( \9945 , \9717 , \8907_nR3482 );
or \U$9119 ( \9946 , \9717 , \9763 );
nand \U$9120 ( \9947 , \9945 , \9946 );
and \U$9121 ( \9948 , \9944 , \9947 );
and \U$9122 ( \9949 , \9717 , \9763 );
and \U$9123 ( \9950 , \9949 , \8907_nR3482 );
and \U$9124 ( \9951 , \8864_nR335c , \9766 );
nor \U$9125 ( \9952 , \9948 , \9950 , \9951 );
xor \U$9126 ( \9953 , \9952 , \9712 );
nand \U$9127 ( \9954 , \9063_nR3133 , \9542 );
or \U$9128 ( \9955 , \9411 , \8966_nR3254 );
nand \U$9129 ( \9956 , \9955 , \9699 );
and \U$9130 ( \9957 , \9954 , \9956 );
and \U$9131 ( \9958 , \9702 , \8966_nR3254 );
and \U$9132 ( \9959 , \9063_nR3133 , \9544 );
nor \U$9133 ( \9960 , \9957 , \9958 , \9959 );
and \U$9134 ( \9961 , \9953 , \9960 );
and \U$9135 ( \9962 , \9952 , \9712 );
or \U$9136 ( \9963 , \9961 , \9962 );
nor \U$9137 ( \9964 , \9943 , \9963 );
not \U$9138 ( \9965 , \9779 );
not \U$9139 ( \9966 , \9771 );
and \U$9140 ( \9967 , \9965 , \9966 );
and \U$9141 ( \9968 , \9779 , \9771 );
nor \U$9142 ( \9969 , \9967 , \9968 );
xor \U$9143 ( \9970 , \9788 , \9795 );
xor \U$9144 ( \9971 , \9970 , \9803 );
and \U$9145 ( \9972 , \9969 , \9971 );
xnor \U$9146 ( \9973 , \9900 , \9907 );
xor \U$9147 ( \9974 , \9788 , \9795 );
xor \U$9148 ( \9975 , \9974 , \9803 );
and \U$9149 ( \9976 , \9973 , \9975 );
and \U$9150 ( \9977 , \9969 , \9973 );
or \U$9151 ( \9978 , \9972 , \9976 , \9977 );
not \U$9152 ( \9979 , \9978 );
and \U$9153 ( \9980 , \9964 , \9979 );
xor \U$9154 ( \9981 , \9918 , \9980 );
not \U$9155 ( \9982 , \9758 );
xor \U$9156 ( \9983 , \9756 , \9754 );
not \U$9157 ( \9984 , \9983 );
or \U$9158 ( \9985 , \9982 , \9984 );
or \U$9159 ( \9986 , \9983 , \9758 );
nand \U$9160 ( \9987 , \9985 , \9986 );
and \U$9161 ( \9988 , \9981 , \9987 );
and \U$9162 ( \9989 , \9918 , \9980 );
or \U$9163 ( \9990 , \9988 , \9989 );
xor \U$9164 ( \9991 , \9759 , \9846 );
xor \U$9165 ( \9992 , \9991 , \9848 );
and \U$9166 ( \9993 , \9990 , \9992 );
and \U$9167 ( \9994 , \9865 , \9990 );
or \U$9168 ( \9995 , \9868 , \9993 , \9994 );
xor \U$9169 ( \9996 , \9851 , \9852 );
xor \U$9170 ( \9997 , \9996 , \9855 );
xor \U$9171 ( \9998 , \9995 , \9997 );
xor \U$9172 ( \9999 , \9759 , \9846 );
xor \U$9173 ( \10000 , \9999 , \9848 );
xor \U$9174 ( \10001 , \9865 , \9990 );
xor \U$9175 ( \10002 , \10000 , \10001 );
xor \U$9176 ( \10003 , \9788 , \9795 );
xor \U$9177 ( \10004 , \10003 , \9803 );
xor \U$9178 ( \10005 , \9969 , \9973 );
xor \U$9179 ( \10006 , \10004 , \10005 );
not \U$9180 ( \10007 , \9712 );
or \U$9181 ( \10008 , \10007 , \8907_nR3482 );
or \U$9182 ( \10009 , \8697 , \8696_nR23dd );
nand \U$9183 ( \10010 , \10009 , \8698 );
nor \U$9184 ( \10011 , \10007 , \10010 );
not \U$9185 ( \10012 , \10011 );
nand \U$9186 ( \10013 , \9712 , \10012 );
nand \U$9187 ( \10014 , \10008 , \10013 );
not \U$9188 ( \10015 , \10014 );
nand \U$9189 ( \10016 , \8966_nR3254 , \9764 );
or \U$9190 ( \10017 , \9717 , \8864_nR335c );
nand \U$9191 ( \10018 , \10017 , \9946 );
and \U$9192 ( \10019 , \10016 , \10018 );
and \U$9193 ( \10020 , \9949 , \8864_nR335c );
and \U$9194 ( \10021 , \8966_nR3254 , \9766 );
nor \U$9195 ( \10022 , \10019 , \10020 , \10021 );
nor \U$9196 ( \10023 , \10015 , \10022 );
not \U$9197 ( \10024 , \10023 );
and \U$9198 ( \10025 , \9843_nR2a34 , \8981 );
or \U$9199 ( \10026 , \8935 , \9687_nR2b14 );
nand \U$9200 ( \10027 , \10026 , \9018 );
nand \U$9201 ( \10028 , \9843_nR2a34 , \8978 );
and \U$9202 ( \10029 , \10027 , \10028 );
and \U$9203 ( \10030 , \9687_nR2b14 , \9022 );
nor \U$9204 ( \10031 , \10025 , \10029 , \10030 );
and \U$9205 ( \10032 , \8853 , RIb557830_453);
and \U$9206 ( \10033 , \8859 , RIb557ec0_467);
and \U$9207 ( \10034 , RIb557e48_466, \8844 );
nor \U$9208 ( \10035 , \10033 , \10034 );
and \U$9209 ( \10036 , \8806 , RIb557998_456);
and \U$9210 ( \10037 , RIb557920_455, \8829 );
nor \U$9211 ( \10038 , \10036 , \10037 );
and \U$9212 ( \10039 , \8816 , RIb5577b8_452);
and \U$9213 ( \10040 , RIb557a10_457, \8812 );
nor \U$9214 ( \10041 , \10039 , \10040 );
and \U$9215 ( \10042 , \8835 , RIb557d58_464);
and \U$9216 ( \10043 , RIb557dd0_465, \8839 );
nor \U$9217 ( \10044 , \10042 , \10043 );
nand \U$9218 ( \10045 , \10035 , \10038 , \10041 , \10044 );
and \U$9219 ( \10046 , \8825 , RIb557bf0_461);
and \U$9220 ( \10047 , RIb5578a8_454, \8831 );
nor \U$9221 ( \10048 , \10046 , \10047 );
not \U$9222 ( \10049 , \10048 );
nor \U$9223 ( \10050 , \10032 , \10045 , \10049 );
and \U$9224 ( \10051 , \8850 , RIb557b00_459);
and \U$9225 ( \10052 , RIb557a88_458, \8847 );
nor \U$9226 ( \10053 , \10051 , \10052 );
and \U$9227 ( \10054 , \8818 , RIb557b78_460);
and \U$9228 ( \10055 , RIb557c68_462, \8823 );
nor \U$9229 ( \10056 , \10054 , \10055 );
and \U$9230 ( \10057 , \8856 , RIb557f38_468);
and \U$9231 ( \10058 , RIb557ce0_463, \8800 );
nor \U$9232 ( \10059 , \10057 , \10058 );
nand \U$9233 ( \10060 , \10050 , \10053 , \10056 , \10059 );
_DC r27cd ( \10061_nR27cd , \10060 , \8863 );
nand \U$9234 ( \10062 , \10061_nR27cd , \8768 );
and \U$9235 ( \10063 , \10031 , \10062 );
and \U$9236 ( \10064 , \9899_nR2959 , \8921 );
and \U$9237 ( \10065 , \8825 , RIb5583e8_478);
and \U$9238 ( \10066 , \8844 , RIb558640_483);
and \U$9239 ( \10067 , RIb5585c8_482, \8839 );
nor \U$9240 ( \10068 , \10066 , \10067 );
and \U$9241 ( \10069 , \8816 , RIb557fb0_469);
and \U$9242 ( \10070 , RIb558208_474, \8812 );
nor \U$9243 ( \10071 , \10069 , \10070 );
and \U$9244 ( \10072 , \8835 , RIb558550_481);
and \U$9245 ( \10073 , RIb5584d8_480, \8800 );
nor \U$9246 ( \10074 , \10072 , \10073 );
and \U$9247 ( \10075 , \8806 , RIb558190_473);
and \U$9248 ( \10076 , RIb558118_472, \8829 );
nor \U$9249 ( \10077 , \10075 , \10076 );
nand \U$9250 ( \10078 , \10068 , \10071 , \10074 , \10077 );
and \U$9251 ( \10079 , \8859 , RIb5586b8_484);
and \U$9252 ( \10080 , RIb558460_479, \8823 );
nor \U$9253 ( \10081 , \10079 , \10080 );
not \U$9254 ( \10082 , \10081 );
nor \U$9255 ( \10083 , \10065 , \10078 , \10082 );
and \U$9256 ( \10084 , \8850 , RIb5582f8_476);
and \U$9257 ( \10085 , RIb558280_475, \8847 );
nor \U$9258 ( \10086 , \10084 , \10085 );
and \U$9259 ( \10087 , \8831 , RIb5580a0_471);
and \U$9260 ( \10088 , RIb558028_470, \8853 );
nor \U$9261 ( \10089 , \10087 , \10088 );
and \U$9262 ( \10090 , \8856 , RIb558730_485);
and \U$9263 ( \10091 , RIb558370_477, \8818 );
nor \U$9264 ( \10092 , \10090 , \10091 );
nand \U$9265 ( \10093 , \10083 , \10086 , \10089 , \10092 );
_DC r289e ( \10094_nR289e , \10093 , \8863 );
or \U$9266 ( \10095 , \8877 , \10094_nR289e );
nand \U$9267 ( \10096 , \10095 , \8917 );
nand \U$9268 ( \10097 , \9899_nR2959 , \8912 );
and \U$9269 ( \10098 , \10096 , \10097 );
and \U$9270 ( \10099 , \10094_nR289e , \8914 );
nor \U$9271 ( \10100 , \10064 , \10098 , \10099 );
nor \U$9272 ( \10101 , \10063 , \10100 );
not \U$9273 ( \10102 , \10101 );
nand \U$9274 ( \10103 , \9271_nR2e0d , \9310 );
or \U$9275 ( \10104 , \9240 , \9177_nR2f04 );
nand \U$9276 ( \10105 , \10104 , \9396 );
and \U$9277 ( \10106 , \10103 , \10105 );
and \U$9278 ( \10107 , \9399 , \9177_nR2f04 );
and \U$9279 ( \10108 , \9271_nR2e0d , \9312 );
nor \U$9280 ( \10109 , \10106 , \10107 , \10108 );
nand \U$9281 ( \10110 , \9122_nR301c , \9542 );
or \U$9282 ( \10111 , \9411 , \9063_nR3133 );
nand \U$9283 ( \10112 , \10111 , \9699 );
and \U$9284 ( \10113 , \10110 , \10112 );
and \U$9285 ( \10114 , \9702 , \9063_nR3133 );
and \U$9286 ( \10115 , \9122_nR301c , \9544 );
nor \U$9287 ( \10116 , \10113 , \10114 , \10115 );
xor \U$9288 ( \10117 , \10109 , \10116 );
nand \U$9289 ( \10118 , \9354_nR2cff , \9139 );
or \U$9290 ( \10119 , \9030 , \9462_nR2c1e );
nand \U$9291 ( \10120 , \10119 , \9144 );
and \U$9292 ( \10121 , \10118 , \10120 );
and \U$9293 ( \10122 , \9141 , \9462_nR2c1e );
and \U$9294 ( \10123 , \9354_nR2cff , \9224 );
nor \U$9295 ( \10124 , \10121 , \10122 , \10123 );
and \U$9296 ( \10125 , \10117 , \10124 );
and \U$9297 ( \10126 , \10109 , \10116 );
or \U$9298 ( \10127 , \10125 , \10126 );
nand \U$9299 ( \10128 , \10102 , \10127 );
not \U$9300 ( \10129 , \10128 );
or \U$9301 ( \10130 , \10024 , \10129 );
not \U$9302 ( \10131 , \10127 );
nand \U$9303 ( \10132 , \10131 , \10101 );
nand \U$9304 ( \10133 , \10130 , \10132 );
nand \U$9305 ( \10134 , \10094_nR289e , \8768 );
and \U$9306 ( \10135 , \9843_nR2a34 , \8921 );
or \U$9307 ( \10136 , \8877 , \9899_nR2959 );
nand \U$9308 ( \10137 , \10136 , \8917 );
nand \U$9309 ( \10138 , \9843_nR2a34 , \8912 );
and \U$9310 ( \10139 , \10137 , \10138 );
and \U$9311 ( \10140 , \9899_nR2959 , \8914 );
nor \U$9312 ( \10141 , \10135 , \10139 , \10140 );
xor \U$9313 ( \10142 , \10134 , \10141 );
nor \U$9314 ( \10143 , \10133 , \10142 );
or \U$9315 ( \10144 , \10006 , \10143 );
nand \U$9316 ( \10145 , \10142 , \10133 );
nand \U$9317 ( \10146 , \10144 , \10145 );
xor \U$9318 ( \10147 , \9964 , \9979 );
xor \U$9319 ( \10148 , \10146 , \10147 );
xor \U$9320 ( \10149 , \9910 , \9917 );
and \U$9321 ( \10150 , \10148 , \10149 );
and \U$9322 ( \10151 , \10146 , \10147 );
or \U$9323 ( \10152 , \10150 , \10151 );
xor \U$9324 ( \10153 , \9807 , \9845 );
xor \U$9325 ( \10154 , \10152 , \10153 );
xor \U$9326 ( \10155 , \9918 , \9980 );
xor \U$9327 ( \10156 , \10155 , \9987 );
and \U$9328 ( \10157 , \10154 , \10156 );
and \U$9329 ( \10158 , \10152 , \10153 );
or \U$9330 ( \10159 , \10157 , \10158 );
xor \U$9331 ( \10160 , \10002 , \10159 );
xor \U$9332 ( \10161 , \10152 , \10153 );
xor \U$9333 ( \10162 , \10161 , \10156 );
not \U$9334 ( \10163 , \9963 );
or \U$9335 ( \10164 , \9943 , \10163 );
not \U$9336 ( \10165 , \9943 );
or \U$9337 ( \10166 , \9963 , \10165 );
or \U$9338 ( \10167 , \10134 , \10141 );
nand \U$9339 ( \10168 , \10164 , \10166 , \10167 );
not \U$9340 ( \10169 , \10168 );
not \U$9341 ( \10170 , \10145 );
nor \U$9342 ( \10171 , \10170 , \10143 );
not \U$9343 ( \10172 , \10171 );
not \U$9344 ( \10173 , \10006 );
and \U$9345 ( \10174 , \10172 , \10173 );
and \U$9346 ( \10175 , \10171 , \10006 );
nor \U$9347 ( \10176 , \10174 , \10175 );
nor \U$9348 ( \10177 , \10169 , \10176 );
xor \U$9349 ( \10178 , \9952 , \9712 );
xor \U$9350 ( \10179 , \10178 , \9960 );
xor \U$9351 ( \10180 , \10142 , \10179 );
nand \U$9352 ( \10181 , \10132 , \10128 );
not \U$9353 ( \10182 , \10181 );
not \U$9354 ( \10183 , \10023 );
and \U$9355 ( \10184 , \10182 , \10183 );
and \U$9356 ( \10185 , \10181 , \10023 );
nor \U$9357 ( \10186 , \10184 , \10185 );
and \U$9358 ( \10187 , \10180 , \10186 );
and \U$9359 ( \10188 , \10142 , \10179 );
or \U$9360 ( \10189 , \10187 , \10188 );
xor \U$9361 ( \10190 , \9925 , \9932 );
xor \U$9362 ( \10191 , \10190 , \9940 );
nand \U$9363 ( \10192 , \9063_nR3133 , \9764 );
or \U$9364 ( \10193 , \9717 , \8966_nR3254 );
nand \U$9365 ( \10194 , \10193 , \9946 );
and \U$9366 ( \10195 , \10192 , \10194 );
and \U$9367 ( \10196 , \9949 , \8966_nR3254 );
and \U$9368 ( \10197 , \9063_nR3133 , \9766 );
nor \U$9369 ( \10198 , \10195 , \10196 , \10197 );
not \U$9370 ( \10199 , \10013 );
and \U$9371 ( \10200 , \8909 , \10199 );
and \U$9372 ( \10201 , \10011 , \8865 );
nand \U$9373 ( \10202 , \10010 , \10007 );
not \U$9374 ( \10203 , \10202 );
and \U$9375 ( \10204 , \8907_nR3482 , \10203 );
nor \U$9376 ( \10205 , \10200 , \10201 , \10204 );
xor \U$9377 ( \10206 , \10198 , \10205 );
nand \U$9378 ( \10207 , \9177_nR2f04 , \9542 );
or \U$9379 ( \10208 , \9411 , \9122_nR301c );
nand \U$9380 ( \10209 , \10208 , \9699 );
and \U$9381 ( \10210 , \10207 , \10209 );
and \U$9382 ( \10211 , \9702 , \9122_nR301c );
and \U$9383 ( \10212 , \9177_nR2f04 , \9544 );
nor \U$9384 ( \10213 , \10210 , \10211 , \10212 );
and \U$9385 ( \10214 , \10206 , \10213 );
and \U$9386 ( \10215 , \10198 , \10205 );
or \U$9387 ( \10216 , \10214 , \10215 );
not \U$9388 ( \10217 , \10216 );
nand \U$9389 ( \10218 , \9462_nR2c1e , \9139 );
or \U$9390 ( \10219 , \9030 , \9687_nR2b14 );
nand \U$9391 ( \10220 , \10219 , \9144 );
and \U$9392 ( \10221 , \10218 , \10220 );
and \U$9393 ( \10222 , \9141 , \9687_nR2b14 );
and \U$9394 ( \10223 , \9462_nR2c1e , \9224 );
nor \U$9395 ( \10224 , \10221 , \10222 , \10223 );
nand \U$9396 ( \10225 , \9354_nR2cff , \9310 );
or \U$9397 ( \10226 , \9240 , \9271_nR2e0d );
nand \U$9398 ( \10227 , \10226 , \9396 );
and \U$9399 ( \10228 , \10225 , \10227 );
and \U$9400 ( \10229 , \9399 , \9271_nR2e0d );
and \U$9401 ( \10230 , \9354_nR2cff , \9312 );
nor \U$9402 ( \10231 , \10228 , \10229 , \10230 );
xor \U$9403 ( \10232 , \10224 , \10231 );
and \U$9404 ( \10233 , \9899_nR2959 , \8981 );
or \U$9405 ( \10234 , \8935 , \9843_nR2a34 );
nand \U$9406 ( \10235 , \10234 , \9018 );
nand \U$9407 ( \10236 , \9899_nR2959 , \8978 );
and \U$9408 ( \10237 , \10235 , \10236 );
and \U$9409 ( \10238 , \9843_nR2a34 , \9022 );
nor \U$9410 ( \10239 , \10233 , \10237 , \10238 );
and \U$9411 ( \10240 , \10232 , \10239 );
and \U$9412 ( \10241 , \10224 , \10231 );
or \U$9413 ( \10242 , \10240 , \10241 );
not \U$9414 ( \10243 , \10242 );
nand \U$9415 ( \10244 , \10217 , \10243 );
xor \U$9416 ( \10245 , \10191 , \10244 );
xor \U$9417 ( \10246 , \10109 , \10116 );
xor \U$9418 ( \10247 , \10246 , \10124 );
not \U$9419 ( \10248 , \10247 );
not \U$9420 ( \10249 , \10062 );
not \U$9421 ( \10250 , \10100 );
not \U$9422 ( \10251 , \10031 );
and \U$9423 ( \10252 , \10250 , \10251 );
and \U$9424 ( \10253 , \10100 , \10031 );
nor \U$9425 ( \10254 , \10252 , \10253 );
not \U$9426 ( \10255 , \10254 );
or \U$9427 ( \10256 , \10249 , \10255 );
or \U$9428 ( \10257 , \10254 , \10062 );
nand \U$9429 ( \10258 , \10256 , \10257 );
nand \U$9430 ( \10259 , \10248 , \10258 );
and \U$9431 ( \10260 , \10245 , \10259 );
and \U$9432 ( \10261 , \10191 , \10244 );
or \U$9433 ( \10262 , \10260 , \10261 );
nand \U$9434 ( \10263 , \10189 , \10262 );
xor \U$9435 ( \10264 , \10177 , \10263 );
xor \U$9436 ( \10265 , \10146 , \10147 );
xor \U$9437 ( \10266 , \10265 , \10149 );
and \U$9438 ( \10267 , \10264 , \10266 );
and \U$9439 ( \10268 , \10177 , \10263 );
or \U$9440 ( \10269 , \10267 , \10268 );
xor \U$9441 ( \10270 , \10162 , \10269 );
xor \U$9442 ( \10271 , \10177 , \10263 );
xor \U$9443 ( \10272 , \10271 , \10266 );
not \U$9444 ( \10273 , \10022 );
not \U$9445 ( \10274 , \10014 );
and \U$9446 ( \10275 , \10273 , \10274 );
and \U$9447 ( \10276 , \10022 , \10014 );
nor \U$9448 ( \10277 , \10275 , \10276 );
and \U$9449 ( \10278 , \10094_nR289e , \8981 );
or \U$9450 ( \10279 , \8935 , \9899_nR2959 );
nand \U$9451 ( \10280 , \10279 , \9018 );
nand \U$9452 ( \10281 , \10094_nR289e , \8978 );
and \U$9453 ( \10282 , \10280 , \10281 );
and \U$9454 ( \10283 , \9899_nR2959 , \9022 );
nor \U$9455 ( \10284 , \10278 , \10282 , \10283 );
and \U$9456 ( \10285 , \8853 , RIb558820_487);
and \U$9457 ( \10286 , \8844 , RIb558e38_500);
and \U$9458 ( \10287 , RIb558dc0_499, \8839 );
nor \U$9459 ( \10288 , \10286 , \10287 );
and \U$9460 ( \10289 , \8816 , RIb5587a8_486);
and \U$9461 ( \10290 , RIb558a00_491, \8812 );
nor \U$9462 ( \10291 , \10289 , \10290 );
and \U$9463 ( \10292 , \8835 , RIb558d48_498);
and \U$9464 ( \10293 , RIb558cd0_497, \8800 );
nor \U$9465 ( \10294 , \10292 , \10293 );
and \U$9466 ( \10295 , \8806 , RIb558988_490);
and \U$9467 ( \10296 , RIb558910_489, \8829 );
nor \U$9468 ( \10297 , \10295 , \10296 );
nand \U$9469 ( \10298 , \10288 , \10291 , \10294 , \10297 );
and \U$9470 ( \10299 , \8847 , RIb558a78_492);
and \U$9471 ( \10300 , RIb558898_488, \8831 );
nor \U$9472 ( \10301 , \10299 , \10300 );
not \U$9473 ( \10302 , \10301 );
nor \U$9474 ( \10303 , \10285 , \10298 , \10302 );
and \U$9475 ( \10304 , \8818 , RIb558b68_494);
and \U$9476 ( \10305 , RIb558af0_493, \8850 );
nor \U$9477 ( \10306 , \10304 , \10305 );
and \U$9478 ( \10307 , \8823 , RIb558c58_496);
and \U$9479 ( \10308 , RIb558be0_495, \8825 );
nor \U$9480 ( \10309 , \10307 , \10308 );
and \U$9481 ( \10310 , \8856 , RIb558f28_502);
and \U$9482 ( \10311 , RIb558eb0_501, \8859 );
nor \U$9483 ( \10312 , \10310 , \10311 );
nand \U$9484 ( \10313 , \10303 , \10306 , \10309 , \10312 );
_DC r2685 ( \10314_nR2685 , \10313 , \8863 );
nand \U$9485 ( \10315 , \10314_nR2685 , \8768 );
and \U$9486 ( \10316 , \10284 , \10315 );
and \U$9487 ( \10317 , \10061_nR27cd , \8921 );
and \U$9488 ( \10318 , \8847 , RIb559270_509);
and \U$9489 ( \10319 , \8844 , RIb559630_517);
and \U$9490 ( \10320 , RIb5595b8_516, \8839 );
nor \U$9491 ( \10321 , \10319 , \10320 );
and \U$9492 ( \10322 , \8816 , RIb558fa0_503);
and \U$9493 ( \10323 , RIb559108_506, \8829 );
nor \U$9494 ( \10324 , \10322 , \10323 );
and \U$9495 ( \10325 , \8835 , RIb559540_515);
and \U$9496 ( \10326 , RIb5594c8_514, \8800 );
nor \U$9497 ( \10327 , \10325 , \10326 );
and \U$9498 ( \10328 , \8806 , RIb559180_507);
and \U$9499 ( \10329 , RIb5591f8_508, \8812 );
nor \U$9500 ( \10330 , \10328 , \10329 );
nand \U$9501 ( \10331 , \10321 , \10324 , \10327 , \10330 );
and \U$9502 ( \10332 , \8818 , RIb559360_511);
and \U$9503 ( \10333 , RIb5592e8_510, \8850 );
nor \U$9504 ( \10334 , \10332 , \10333 );
not \U$9505 ( \10335 , \10334 );
nor \U$9506 ( \10336 , \10318 , \10331 , \10335 );
and \U$9507 ( \10337 , \8831 , RIb559090_505);
and \U$9508 ( \10338 , RIb559018_504, \8853 );
nor \U$9509 ( \10339 , \10337 , \10338 );
and \U$9510 ( \10340 , \8823 , RIb559450_513);
and \U$9511 ( \10341 , RIb5593d8_512, \8825 );
nor \U$9512 ( \10342 , \10340 , \10341 );
and \U$9513 ( \10343 , \8856 , RIb559720_519);
and \U$9514 ( \10344 , RIb5596a8_518, \8859 );
nor \U$9515 ( \10345 , \10343 , \10344 );
nand \U$9516 ( \10346 , \10336 , \10339 , \10342 , \10345 );
_DC r272f ( \10347_nR272f , \10346 , \8863 );
or \U$9517 ( \10348 , \8877 , \10347_nR272f );
nand \U$9518 ( \10349 , \10348 , \8917 );
nand \U$9519 ( \10350 , \10061_nR27cd , \8912 );
and \U$9520 ( \10351 , \10349 , \10350 );
and \U$9521 ( \10352 , \10347_nR272f , \8914 );
nor \U$9522 ( \10353 , \10317 , \10351 , \10352 );
nor \U$9523 ( \10354 , \10316 , \10353 );
not \U$9524 ( \10355 , \10354 );
nand \U$9525 ( \10356 , \9462_nR2c1e , \9310 );
or \U$9526 ( \10357 , \9240 , \9354_nR2cff );
nand \U$9527 ( \10358 , \10357 , \9396 );
and \U$9528 ( \10359 , \10356 , \10358 );
and \U$9529 ( \10360 , \9399 , \9354_nR2cff );
and \U$9530 ( \10361 , \9462_nR2c1e , \9312 );
nor \U$9531 ( \10362 , \10359 , \10360 , \10361 );
nand \U$9532 ( \10363 , \9271_nR2e0d , \9542 );
or \U$9533 ( \10364 , \9411 , \9177_nR2f04 );
nand \U$9534 ( \10365 , \10364 , \9699 );
and \U$9535 ( \10366 , \10363 , \10365 );
and \U$9536 ( \10367 , \9702 , \9177_nR2f04 );
and \U$9537 ( \10368 , \9271_nR2e0d , \9544 );
nor \U$9538 ( \10369 , \10366 , \10367 , \10368 );
xor \U$9539 ( \10370 , \10362 , \10369 );
nand \U$9540 ( \10371 , \9687_nR2b14 , \9139 );
or \U$9541 ( \10372 , \9030 , \9843_nR2a34 );
nand \U$9542 ( \10373 , \10372 , \9144 );
and \U$9543 ( \10374 , \10371 , \10373 );
and \U$9544 ( \10375 , \9141 , \9843_nR2a34 );
and \U$9545 ( \10376 , \9687_nR2b14 , \9224 );
nor \U$9546 ( \10377 , \10374 , \10375 , \10376 );
and \U$9547 ( \10378 , \10370 , \10377 );
and \U$9548 ( \10379 , \10362 , \10369 );
or \U$9549 ( \10380 , \10378 , \10379 );
nand \U$9550 ( \10381 , \10355 , \10380 );
or \U$9551 ( \10382 , \10202 , \8865 );
or \U$9552 ( \10383 , \8864_nR335c , \10013 );
or \U$9553 ( \10384 , \8966_nR3254 , \10012 );
nand \U$9554 ( \10385 , \10382 , \10383 , \10384 );
or \U$9555 ( \10386 , \9767 , \9123 );
or \U$9556 ( \10387 , \9717 , \9063_nR3133 );
nand \U$9557 ( \10388 , \10387 , \9946 );
nand \U$9558 ( \10389 , \9122_nR301c , \9764 );
and \U$9559 ( \10390 , \10388 , \10389 );
and \U$9560 ( \10391 , \9063_nR3133 , \9949 );
nor \U$9561 ( \10392 , \10390 , \10391 );
nand \U$9562 ( \10393 , \10386 , \10392 );
and \U$9563 ( \10394 , \10385 , \10393 );
and \U$9564 ( \10395 , \10381 , \10394 );
not \U$9565 ( \10396 , \10354 );
nor \U$9566 ( \10397 , \10396 , \10380 );
nor \U$9567 ( \10398 , \10395 , \10397 );
nand \U$9568 ( \10399 , \10277 , \10398 );
xor \U$9569 ( \10400 , \10224 , \10231 );
xor \U$9570 ( \10401 , \10400 , \10239 );
not \U$9571 ( \10402 , \10401 );
nand \U$9572 ( \10403 , \10347_nR272f , \8768 );
and \U$9573 ( \10404 , \10094_nR289e , \8921 );
or \U$9574 ( \10405 , \8877 , \10061_nR27cd );
nand \U$9575 ( \10406 , \10405 , \8917 );
nand \U$9576 ( \10407 , \10094_nR289e , \8912 );
and \U$9577 ( \10408 , \10406 , \10407 );
and \U$9578 ( \10409 , \10061_nR27cd , \8914 );
nor \U$9579 ( \10410 , \10404 , \10408 , \10409 );
xor \U$9580 ( \10411 , \10403 , \10410 );
and \U$9581 ( \10412 , \10402 , \10411 );
and \U$9582 ( \10413 , \10399 , \10412 );
nor \U$9583 ( \10414 , \10398 , \10277 );
nor \U$9584 ( \10415 , \10413 , \10414 );
not \U$9585 ( \10416 , \10258 );
not \U$9586 ( \10417 , \10247 );
and \U$9587 ( \10418 , \10416 , \10417 );
and \U$9588 ( \10419 , \10258 , \10247 );
nor \U$9589 ( \10420 , \10418 , \10419 );
not \U$9590 ( \10421 , \10420 );
or \U$9591 ( \10422 , \10242 , \10217 );
or \U$9592 ( \10423 , \10216 , \10243 );
or \U$9593 ( \10424 , \10403 , \10410 );
nand \U$9594 ( \10425 , \10422 , \10423 , \10424 );
nand \U$9595 ( \10426 , \10421 , \10425 );
xor \U$9596 ( \10427 , \10415 , \10426 );
xor \U$9597 ( \10428 , \10142 , \10179 );
xor \U$9598 ( \10429 , \10428 , \10186 );
and \U$9599 ( \10430 , \10427 , \10429 );
and \U$9600 ( \10431 , \10415 , \10426 );
or \U$9601 ( \10432 , \10430 , \10431 );
xor \U$9602 ( \10433 , \10189 , \10262 );
xor \U$9603 ( \10434 , \10432 , \10433 );
not \U$9604 ( \10435 , \10176 );
not \U$9605 ( \10436 , \10168 );
and \U$9606 ( \10437 , \10435 , \10436 );
and \U$9607 ( \10438 , \10176 , \10168 );
nor \U$9608 ( \10439 , \10437 , \10438 );
and \U$9609 ( \10440 , \10434 , \10439 );
and \U$9610 ( \10441 , \10432 , \10433 );
or \U$9611 ( \10442 , \10440 , \10441 );
not \U$9612 ( \10443 , \10442 );
xor \U$9613 ( \10444 , \10272 , \10443 );
not \U$9614 ( \10445 , \10425 );
not \U$9615 ( \10446 , \10420 );
or \U$9616 ( \10447 , \10445 , \10446 );
or \U$9617 ( \10448 , \10420 , \10425 );
nand \U$9618 ( \10449 , \10447 , \10448 );
not \U$9619 ( \10450 , \10449 );
not \U$9620 ( \10451 , \10412 );
not \U$9621 ( \10452 , \10414 );
nand \U$9622 ( \10453 , \10452 , \10399 );
not \U$9623 ( \10454 , \10453 );
or \U$9624 ( \10455 , \10451 , \10454 );
or \U$9625 ( \10456 , \10453 , \10412 );
nand \U$9626 ( \10457 , \10455 , \10456 );
not \U$9627 ( \10458 , \10457 );
xor \U$9628 ( \10459 , \10198 , \10205 );
xor \U$9629 ( \10460 , \10459 , \10213 );
not \U$9630 ( \10461 , \10460 );
nand \U$9631 ( \10462 , \9843_nR2a34 , \9139 );
or \U$9632 ( \10463 , \9030 , \9899_nR2959 );
nand \U$9633 ( \10464 , \10463 , \9144 );
and \U$9634 ( \10465 , \10462 , \10464 );
and \U$9635 ( \10466 , \9141 , \9899_nR2959 );
and \U$9636 ( \10467 , \9843_nR2a34 , \9224 );
nor \U$9637 ( \10468 , \10465 , \10466 , \10467 );
nand \U$9638 ( \10469 , \9687_nR2b14 , \9310 );
or \U$9639 ( \10470 , \9240 , \9462_nR2c1e );
nand \U$9640 ( \10471 , \10470 , \9396 );
and \U$9641 ( \10472 , \10469 , \10471 );
and \U$9642 ( \10473 , \9399 , \9462_nR2c1e );
and \U$9643 ( \10474 , \9687_nR2b14 , \9312 );
nor \U$9644 ( \10475 , \10472 , \10473 , \10474 );
xor \U$9645 ( \10476 , \10468 , \10475 );
and \U$9646 ( \10477 , \10061_nR27cd , \8981 );
or \U$9647 ( \10478 , \8935 , \10094_nR289e );
nand \U$9648 ( \10479 , \10478 , \9018 );
nand \U$9649 ( \10480 , \10061_nR27cd , \8978 );
and \U$9650 ( \10481 , \10479 , \10480 );
and \U$9651 ( \10482 , \10094_nR289e , \9022 );
nor \U$9652 ( \10483 , \10477 , \10481 , \10482 );
and \U$9653 ( \10484 , \10476 , \10483 );
and \U$9654 ( \10485 , \10468 , \10475 );
or \U$9655 ( \10486 , \10484 , \10485 );
nand \U$9656 ( \10487 , \9177_nR2f04 , \9764 );
or \U$9657 ( \10488 , \9717 , \9122_nR301c );
nand \U$9658 ( \10489 , \10488 , \9946 );
and \U$9659 ( \10490 , \10487 , \10489 );
and \U$9660 ( \10491 , \9949 , \9122_nR301c );
and \U$9661 ( \10492 , \9177_nR2f04 , \9766 );
nor \U$9662 ( \10493 , \10490 , \10491 , \10492 );
and \U$9663 ( \10494 , \8967 , \10199 );
not \U$9664 ( \10495 , \9063_nR3133 );
and \U$9665 ( \10496 , \10011 , \10495 );
and \U$9666 ( \10497 , \8966_nR3254 , \10203 );
nor \U$9667 ( \10498 , \10494 , \10496 , \10497 );
xor \U$9668 ( \10499 , \10493 , \10498 );
nand \U$9669 ( \10500 , \9354_nR2cff , \9542 );
or \U$9670 ( \10501 , \9411 , \9271_nR2e0d );
nand \U$9671 ( \10502 , \10501 , \9699 );
and \U$9672 ( \10503 , \10500 , \10502 );
and \U$9673 ( \10504 , \9702 , \9271_nR2e0d );
and \U$9674 ( \10505 , \9354_nR2cff , \9544 );
nor \U$9675 ( \10506 , \10503 , \10504 , \10505 );
and \U$9676 ( \10507 , \10499 , \10506 );
and \U$9677 ( \10508 , \10493 , \10498 );
or \U$9678 ( \10509 , \10507 , \10508 );
nor \U$9679 ( \10510 , \10486 , \10509 );
nand \U$9680 ( \10511 , \10461 , \10510 );
not \U$9681 ( \10512 , \10511 );
and \U$9682 ( \10513 , \10458 , \10512 );
and \U$9683 ( \10514 , \10457 , \10511 );
nor \U$9684 ( \10515 , \10513 , \10514 );
not \U$9685 ( \10516 , \10515 );
or \U$9686 ( \10517 , \10450 , \10516 );
or \U$9687 ( \10518 , \10515 , \10449 );
nand \U$9688 ( \10519 , \10517 , \10518 );
not \U$9689 ( \10520 , \10519 );
not \U$9690 ( \10521 , \10460 );
not \U$9691 ( \10522 , \10510 );
or \U$9692 ( \10523 , \10521 , \10522 );
or \U$9693 ( \10524 , \10510 , \10460 );
nand \U$9694 ( \10525 , \10523 , \10524 );
not \U$9695 ( \10526 , \10394 );
not \U$9696 ( \10527 , \10397 );
nand \U$9697 ( \10528 , \10527 , \10381 );
not \U$9698 ( \10529 , \10528 );
or \U$9699 ( \10530 , \10526 , \10529 );
or \U$9700 ( \10531 , \10528 , \10394 );
nand \U$9701 ( \10532 , \10530 , \10531 );
and \U$9702 ( \10533 , \10525 , \10532 );
not \U$9703 ( \10534 , \10533 );
not \U$9704 ( \10535 , \10509 );
or \U$9705 ( \10536 , \10486 , \10535 );
not \U$9706 ( \10537 , \10486 );
or \U$9707 ( \10538 , \10509 , \10537 );
and \U$9708 ( \10539 , \8839 , RIb55a5a8_550);
nand \U$9709 ( \10540 , RIb55a710_553, \8856 );
and \U$9710 ( \10541 , \8823 , RIb55a440_547);
and \U$9711 ( \10542 , RIb55a3c8_546, \8825 );
nor \U$9712 ( \10543 , \10541 , \10542 );
nand \U$9713 ( \10544 , RIb55a698_552, \8859 );
nand \U$9714 ( \10545 , \10540 , \10543 , \10544 );
and \U$9715 ( \10546 , \8835 , RIb55a530_549);
and \U$9716 ( \10547 , RIb55a4b8_548, \8800 );
nor \U$9717 ( \10548 , \10546 , \10547 );
and \U$9718 ( \10549 , \8816 , RIb559f90_537);
and \U$9719 ( \10550 , RIb55a1e8_542, \8812 );
nor \U$9720 ( \10551 , \10549 , \10550 );
nand \U$9721 ( \10552 , \10548 , \10551 );
nor \U$9722 ( \10553 , \10539 , \10545 , \10552 );
and \U$9723 ( \10554 , \8818 , RIb55a350_545);
and \U$9724 ( \10555 , RIb55a2d8_544, \8850 );
nor \U$9725 ( \10556 , \10554 , \10555 );
and \U$9726 ( \10557 , \8806 , RIb55a170_541);
and \U$9727 ( \10558 , RIb55a0f8_540, \8829 );
nor \U$9728 ( \10559 , \10557 , \10558 );
and \U$9729 ( \10560 , RIb55a620_551, \8844 );
and \U$9730 ( \10561 , RIb55a008_538, \8853 );
and \U$9731 ( \10562 , \8847 , RIb55a260_543);
and \U$9732 ( \10563 , RIb55a080_539, \8831 );
nor \U$9733 ( \10564 , \10562 , \10563 );
not \U$9734 ( \10565 , \10564 );
nor \U$9735 ( \10566 , \10560 , \10561 , \10565 );
nand \U$9736 ( \10567 , \10553 , \10556 , \10559 , \10566 );
_DC r260a ( \10568_nR260a , \10567 , \8863 );
nand \U$9737 ( \10569 , \10568_nR260a , \8768 );
and \U$9738 ( \10570 , \10347_nR272f , \8921 );
or \U$9739 ( \10571 , \8877 , \10314_nR2685 );
nand \U$9740 ( \10572 , \10571 , \8917 );
nand \U$9741 ( \10573 , \10347_nR272f , \8912 );
and \U$9742 ( \10574 , \10572 , \10573 );
and \U$9743 ( \10575 , \10314_nR2685 , \8914 );
nor \U$9744 ( \10576 , \10570 , \10574 , \10575 );
or \U$9745 ( \10577 , \10569 , \10576 );
nand \U$9746 ( \10578 , \10536 , \10538 , \10577 );
xor \U$9747 ( \10579 , \10385 , \10393 );
xor \U$9748 ( \10580 , \10578 , \10579 );
not \U$9749 ( \10581 , \10315 );
not \U$9750 ( \10582 , \10353 );
not \U$9751 ( \10583 , \10284 );
and \U$9752 ( \10584 , \10582 , \10583 );
and \U$9753 ( \10585 , \10353 , \10284 );
nor \U$9754 ( \10586 , \10584 , \10585 );
not \U$9755 ( \10587 , \10586 );
or \U$9756 ( \10588 , \10581 , \10587 );
or \U$9757 ( \10589 , \10586 , \10315 );
nand \U$9758 ( \10590 , \10588 , \10589 );
and \U$9759 ( \10591 , \10580 , \10590 );
and \U$9760 ( \10592 , \10578 , \10579 );
or \U$9761 ( \10593 , \10591 , \10592 );
xor \U$9762 ( \10594 , \10402 , \10411 );
and \U$9763 ( \10595 , \10593 , \10594 );
not \U$9764 ( \10596 , \10593 );
not \U$9765 ( \10597 , \10594 );
and \U$9766 ( \10598 , \10596 , \10597 );
xor \U$9767 ( \10599 , \10468 , \10475 );
xor \U$9768 ( \10600 , \10599 , \10483 );
xor \U$9769 ( \10601 , \10493 , \10498 );
xor \U$9770 ( \10602 , \10601 , \10506 );
xor \U$9771 ( \10603 , \10600 , \10602 );
xnor \U$9772 ( \10604 , \10569 , \10576 );
and \U$9773 ( \10605 , \10603 , \10604 );
and \U$9774 ( \10606 , \10600 , \10602 );
or \U$9775 ( \10607 , \10605 , \10606 );
xor \U$9776 ( \10608 , \10362 , \10369 );
xor \U$9777 ( \10609 , \10608 , \10377 );
xor \U$9778 ( \10610 , \10607 , \10609 );
nand \U$9779 ( \10611 , \9843_nR2a34 , \9310 );
or \U$9780 ( \10612 , \9240 , \9687_nR2b14 );
nand \U$9781 ( \10613 , \10612 , \9396 );
and \U$9782 ( \10614 , \10611 , \10613 );
and \U$9783 ( \10615 , \9399 , \9687_nR2b14 );
and \U$9784 ( \10616 , \9843_nR2a34 , \9312 );
nor \U$9785 ( \10617 , \10614 , \10615 , \10616 );
nand \U$9786 ( \10618 , \9462_nR2c1e , \9542 );
or \U$9787 ( \10619 , \9411 , \9354_nR2cff );
nand \U$9788 ( \10620 , \10619 , \9699 );
and \U$9789 ( \10621 , \10618 , \10620 );
and \U$9790 ( \10622 , \9702 , \9354_nR2cff );
and \U$9791 ( \10623 , \9462_nR2c1e , \9544 );
nor \U$9792 ( \10624 , \10621 , \10622 , \10623 );
xor \U$9793 ( \10625 , \10617 , \10624 );
nand \U$9794 ( \10626 , \9899_nR2959 , \9139 );
or \U$9795 ( \10627 , \9030 , \10094_nR289e );
nand \U$9796 ( \10628 , \10627 , \9144 );
and \U$9797 ( \10629 , \10626 , \10628 );
and \U$9798 ( \10630 , \9141 , \10094_nR289e );
and \U$9799 ( \10631 , \9899_nR2959 , \9224 );
nor \U$9800 ( \10632 , \10629 , \10630 , \10631 );
and \U$9801 ( \10633 , \10625 , \10632 );
and \U$9802 ( \10634 , \10617 , \10624 );
or \U$9803 ( \10635 , \10633 , \10634 );
nand \U$9804 ( \10636 , \9271_nR2e0d , \9764 );
or \U$9805 ( \10637 , \9717 , \9177_nR2f04 );
nand \U$9806 ( \10638 , \10637 , \9946 );
and \U$9807 ( \10639 , \10636 , \10638 );
and \U$9808 ( \10640 , \9949 , \9177_nR2f04 );
and \U$9809 ( \10641 , \9271_nR2e0d , \9766 );
nor \U$9810 ( \10642 , \10639 , \10640 , \10641 );
not \U$9811 ( \10643 , \10642 );
or \U$9812 ( \10644 , \10202 , \10495 );
or \U$9813 ( \10645 , \9063_nR3133 , \10013 );
or \U$9814 ( \10646 , \9122_nR301c , \10012 );
nand \U$9815 ( \10647 , \10644 , \10645 , \10646 );
nand \U$9816 ( \10648 , \10643 , \10647 );
xor \U$9817 ( \10649 , \10635 , \10648 );
and \U$9818 ( \10650 , \10347_nR272f , \8981 );
or \U$9819 ( \10651 , \8935 , \10061_nR27cd );
nand \U$9820 ( \10652 , \10651 , \9018 );
nand \U$9821 ( \10653 , \10347_nR272f , \8978 );
and \U$9822 ( \10654 , \10652 , \10653 );
and \U$9823 ( \10655 , \10061_nR27cd , \9022 );
nor \U$9824 ( \10656 , \10650 , \10654 , \10655 );
and \U$9825 ( \10657 , \8839 , RIb559db0_533);
nand \U$9826 ( \10658 , RIb559f18_536, \8856 );
and \U$9827 ( \10659 , \8823 , RIb559c48_530);
and \U$9828 ( \10660 , RIb559bd0_529, \8825 );
nor \U$9829 ( \10661 , \10659 , \10660 );
nand \U$9830 ( \10662 , RIb559ea0_535, \8859 );
nand \U$9831 ( \10663 , \10658 , \10661 , \10662 );
and \U$9832 ( \10664 , \8835 , RIb559d38_532);
and \U$9833 ( \10665 , RIb559cc0_531, \8800 );
nor \U$9834 ( \10666 , \10664 , \10665 );
and \U$9835 ( \10667 , \8816 , RIb559798_520);
and \U$9836 ( \10668 , RIb5599f0_525, \8812 );
nor \U$9837 ( \10669 , \10667 , \10668 );
nand \U$9838 ( \10670 , \10666 , \10669 );
nor \U$9839 ( \10671 , \10657 , \10663 , \10670 );
and \U$9840 ( \10672 , \8818 , RIb559b58_528);
and \U$9841 ( \10673 , RIb559ae0_527, \8850 );
nor \U$9842 ( \10674 , \10672 , \10673 );
and \U$9843 ( \10675 , \8806 , RIb559978_524);
and \U$9844 ( \10676 , RIb559900_523, \8829 );
nor \U$9845 ( \10677 , \10675 , \10676 );
and \U$9846 ( \10678 , RIb559e28_534, \8844 );
and \U$9847 ( \10679 , RIb559810_521, \8853 );
and \U$9848 ( \10680 , \8847 , RIb559a68_526);
and \U$9849 ( \10681 , RIb559888_522, \8831 );
nor \U$9850 ( \10682 , \10680 , \10681 );
not \U$9851 ( \10683 , \10682 );
nor \U$9852 ( \10684 , \10678 , \10679 , \10683 );
nand \U$9853 ( \10685 , \10671 , \10674 , \10677 , \10684 );
_DC r2587 ( \10686_nR2587 , \10685 , \8863 );
nand \U$9854 ( \10687 , \10686_nR2587 , \8768 );
and \U$9855 ( \10688 , \10656 , \10687 );
and \U$9856 ( \10689 , \10314_nR2685 , \8921 );
or \U$9857 ( \10690 , \8877 , \10568_nR260a );
nand \U$9858 ( \10691 , \10690 , \8917 );
nand \U$9859 ( \10692 , \10314_nR2685 , \8912 );
and \U$9860 ( \10693 , \10691 , \10692 );
and \U$9861 ( \10694 , \10568_nR260a , \8914 );
nor \U$9862 ( \10695 , \10689 , \10693 , \10694 );
nor \U$9863 ( \10696 , \10688 , \10695 );
not \U$9864 ( \10697 , \10696 );
and \U$9865 ( \10698 , \10649 , \10697 );
and \U$9866 ( \10699 , \10635 , \10648 );
or \U$9867 ( \10700 , \10698 , \10699 );
and \U$9868 ( \10701 , \10610 , \10700 );
and \U$9869 ( \10702 , \10607 , \10609 );
or \U$9870 ( \10703 , \10701 , \10702 );
nor \U$9871 ( \10704 , \10598 , \10703 );
nor \U$9872 ( \10705 , \10595 , \10704 );
not \U$9873 ( \10706 , \10705 );
or \U$9874 ( \10707 , \10534 , \10706 );
or \U$9875 ( \10708 , \10705 , \10533 );
nand \U$9876 ( \10709 , \10707 , \10708 );
not \U$9877 ( \10710 , \10709 );
and \U$9878 ( \10711 , \10520 , \10710 );
and \U$9879 ( \10712 , \10519 , \10709 );
nor \U$9880 ( \10713 , \10711 , \10712 );
not \U$9881 ( \10714 , \10703 );
xor \U$9882 ( \10715 , \10594 , \10593 );
not \U$9883 ( \10716 , \10715 );
or \U$9884 ( \10717 , \10714 , \10716 );
or \U$9885 ( \10718 , \10715 , \10703 );
nand \U$9886 ( \10719 , \10717 , \10718 );
xor \U$9887 ( \10720 , \10525 , \10532 );
xor \U$9888 ( \10721 , \10719 , \10720 );
xor \U$9889 ( \10722 , \10578 , \10579 );
xor \U$9890 ( \10723 , \10722 , \10590 );
not \U$9891 ( \10724 , \10723 );
nand \U$9892 ( \10725 , \9354_nR2cff , \9764 );
or \U$9893 ( \10726 , \9717 , \9271_nR2e0d );
nand \U$9894 ( \10727 , \10726 , \9946 );
and \U$9895 ( \10728 , \10725 , \10727 );
and \U$9896 ( \10729 , \9949 , \9271_nR2e0d );
and \U$9897 ( \10730 , \9354_nR2cff , \9766 );
nor \U$9898 ( \10731 , \10728 , \10729 , \10730 );
and \U$9899 ( \10732 , \9123 , \10199 );
not \U$9900 ( \10733 , \9177_nR2f04 );
and \U$9901 ( \10734 , \10011 , \10733 );
and \U$9902 ( \10735 , \9122_nR301c , \10203 );
nor \U$9903 ( \10736 , \10732 , \10734 , \10735 );
xor \U$9904 ( \10737 , \10731 , \10736 );
nand \U$9905 ( \10738 , \9687_nR2b14 , \9542 );
or \U$9906 ( \10739 , \9411 , \9462_nR2c1e );
nand \U$9907 ( \10740 , \10739 , \9699 );
and \U$9908 ( \10741 , \10738 , \10740 );
and \U$9909 ( \10742 , \9702 , \9462_nR2c1e );
and \U$9910 ( \10743 , \9687_nR2b14 , \9544 );
nor \U$9911 ( \10744 , \10741 , \10742 , \10743 );
and \U$9912 ( \10745 , \10737 , \10744 );
and \U$9913 ( \10746 , \10731 , \10736 );
or \U$9914 ( \10747 , \10745 , \10746 );
not \U$9915 ( \10748 , \10747 );
nand \U$9916 ( \10749 , \10094_nR289e , \9139 );
or \U$9917 ( \10750 , \9030 , \10061_nR27cd );
nand \U$9918 ( \10751 , \10750 , \9144 );
and \U$9919 ( \10752 , \10749 , \10751 );
and \U$9920 ( \10753 , \9141 , \10061_nR27cd );
and \U$9921 ( \10754 , \10094_nR289e , \9224 );
nor \U$9922 ( \10755 , \10752 , \10753 , \10754 );
nand \U$9923 ( \10756 , \9899_nR2959 , \9310 );
or \U$9924 ( \10757 , \9240 , \9843_nR2a34 );
nand \U$9925 ( \10758 , \10757 , \9396 );
and \U$9926 ( \10759 , \10756 , \10758 );
and \U$9927 ( \10760 , \9399 , \9843_nR2a34 );
and \U$9928 ( \10761 , \9899_nR2959 , \9312 );
nor \U$9929 ( \10762 , \10759 , \10760 , \10761 );
xor \U$9930 ( \10763 , \10755 , \10762 );
and \U$9931 ( \10764 , \10314_nR2685 , \8981 );
or \U$9932 ( \10765 , \8935 , \10347_nR272f );
nand \U$9933 ( \10766 , \10765 , \9018 );
nand \U$9934 ( \10767 , \10314_nR2685 , \8978 );
and \U$9935 ( \10768 , \10766 , \10767 );
and \U$9936 ( \10769 , \10347_nR272f , \9022 );
nor \U$9937 ( \10770 , \10764 , \10768 , \10769 );
and \U$9938 ( \10771 , \10763 , \10770 );
and \U$9939 ( \10772 , \10755 , \10762 );
or \U$9940 ( \10773 , \10771 , \10772 );
not \U$9941 ( \10774 , \10773 );
nand \U$9942 ( \10775 , \10748 , \10774 );
not \U$9943 ( \10776 , \10775 );
not \U$9944 ( \10777 , \10776 );
not \U$9945 ( \10778 , \10687 );
not \U$9946 ( \10779 , \10695 );
not \U$9947 ( \10780 , \10656 );
and \U$9948 ( \10781 , \10779 , \10780 );
and \U$9949 ( \10782 , \10695 , \10656 );
nor \U$9950 ( \10783 , \10781 , \10782 );
not \U$9951 ( \10784 , \10783 );
or \U$9952 ( \10785 , \10778 , \10784 );
or \U$9953 ( \10786 , \10783 , \10687 );
nand \U$9954 ( \10787 , \10785 , \10786 );
not \U$9955 ( \10788 , \10787 );
xor \U$9956 ( \10789 , \10617 , \10624 );
xor \U$9957 ( \10790 , \10789 , \10632 );
nor \U$9958 ( \10791 , \10788 , \10790 );
not \U$9959 ( \10792 , \10791 );
or \U$9960 ( \10793 , \10777 , \10792 );
not \U$9961 ( \10794 , \10791 );
and \U$9962 ( \10795 , \10775 , \10794 );
xor \U$9963 ( \10796 , \10600 , \10602 );
xor \U$9964 ( \10797 , \10796 , \10604 );
or \U$9965 ( \10798 , \10795 , \10797 );
nand \U$9966 ( \10799 , \10793 , \10798 );
not \U$9967 ( \10800 , \10799 );
or \U$9968 ( \10801 , \10724 , \10800 );
nor \U$9969 ( \10802 , \10799 , \10723 );
xor \U$9970 ( \10803 , \10607 , \10609 );
xor \U$9971 ( \10804 , \10803 , \10700 );
or \U$9972 ( \10805 , \10802 , \10804 );
nand \U$9973 ( \10806 , \10801 , \10805 );
and \U$9974 ( \10807 , \10721 , \10806 );
and \U$9975 ( \10808 , \10719 , \10720 );
or \U$9976 ( \10809 , \10807 , \10808 );
xor \U$9977 ( \10810 , \10713 , \10809 );
xor \U$9978 ( \10811 , \10719 , \10720 );
xor \U$9979 ( \10812 , \10811 , \10806 );
not \U$9980 ( \10813 , \10804 );
not \U$9981 ( \10814 , \10799 );
and \U$9982 ( \10815 , \10813 , \10814 );
and \U$9983 ( \10816 , \10804 , \10799 );
nor \U$9984 ( \10817 , \10815 , \10816 );
not \U$9985 ( \10818 , \10817 );
not \U$9986 ( \10819 , \10723 );
and \U$9987 ( \10820 , \10818 , \10819 );
and \U$9988 ( \10821 , \10817 , \10723 );
nor \U$9989 ( \10822 , \10820 , \10821 );
not \U$9990 ( \10823 , \10787 );
not \U$9991 ( \10824 , \10790 );
and \U$9992 ( \10825 , \10823 , \10824 );
and \U$9993 ( \10826 , \10787 , \10790 );
nor \U$9994 ( \10827 , \10825 , \10826 );
not \U$9995 ( \10828 , \10827 );
or \U$9996 ( \10829 , \10773 , \10748 );
or \U$9997 ( \10830 , \10747 , \10774 );
and \U$9998 ( \10831 , \8825 , RIb55abc0_563);
and \U$9999 ( \10832 , \8847 , RIb55aa58_560);
and \U$10000 ( \10833 , RIb55a9e0_559, \8812 );
nor \U$10001 ( \10834 , \10832 , \10833 );
and \U$10002 ( \10835 , \8806 , RIb55a968_558);
and \U$10003 ( \10836 , RIb55a8f0_557, \8829 );
nor \U$10004 ( \10837 , \10835 , \10836 );
and \U$10005 ( \10838 , \8816 , RIb55a788_554);
and \U$10006 ( \10839 , RIb55ac38_564, \8823 );
nor \U$10007 ( \10840 , \10838 , \10839 );
and \U$10008 ( \10841 , \8818 , RIb55ab48_562);
and \U$10009 ( \10842 , RIb55aad0_561, \8850 );
nor \U$10010 ( \10843 , \10841 , \10842 );
nand \U$10011 ( \10844 , \10834 , \10837 , \10840 , \10843 );
and \U$10012 ( \10845 , \8859 , RIb55ae90_569);
and \U$10013 ( \10846 , RIb55ae18_568, \8844 );
nor \U$10014 ( \10847 , \10845 , \10846 );
not \U$10015 ( \10848 , \10847 );
nor \U$10016 ( \10849 , \10831 , \10844 , \10848 );
and \U$10017 ( \10850 , \8831 , RIb55a878_556);
and \U$10018 ( \10851 , RIb55a800_555, \8853 );
nor \U$10019 ( \10852 , \10850 , \10851 );
and \U$10020 ( \10853 , \8835 , RIb55ad28_566);
and \U$10021 ( \10854 , RIb55acb0_565, \8800 );
nor \U$10022 ( \10855 , \10853 , \10854 );
and \U$10023 ( \10856 , \8856 , RIb55af08_570);
and \U$10024 ( \10857 , RIb55ada0_567, \8839 );
nor \U$10025 ( \10858 , \10856 , \10857 );
nand \U$10026 ( \10859 , \10849 , \10852 , \10855 , \10858 );
_DC r251b ( \10860_nR251b , \10859 , \8863 );
nand \U$10027 ( \10861 , \10860_nR251b , \8768 );
and \U$10028 ( \10862 , \10568_nR260a , \8921 );
or \U$10029 ( \10863 , \8877 , \10686_nR2587 );
nand \U$10030 ( \10864 , \10863 , \8917 );
nand \U$10031 ( \10865 , \10568_nR260a , \8912 );
and \U$10032 ( \10866 , \10864 , \10865 );
and \U$10033 ( \10867 , \10686_nR2587 , \8914 );
nor \U$10034 ( \10868 , \10862 , \10866 , \10867 );
or \U$10035 ( \10869 , \10861 , \10868 );
nand \U$10036 ( \10870 , \10829 , \10830 , \10869 );
nand \U$10037 ( \10871 , \10828 , \10870 );
xor \U$10038 ( \10872 , \10635 , \10648 );
xor \U$10039 ( \10873 , \10872 , \10697 );
xor \U$10040 ( \10874 , \10871 , \10873 );
xor \U$10041 ( \10875 , \10755 , \10762 );
xor \U$10042 ( \10876 , \10875 , \10770 );
xor \U$10043 ( \10877 , \10731 , \10736 );
xor \U$10044 ( \10878 , \10877 , \10744 );
xor \U$10045 ( \10879 , \10876 , \10878 );
xnor \U$10046 ( \10880 , \10861 , \10868 );
and \U$10047 ( \10881 , \10879 , \10880 );
and \U$10048 ( \10882 , \10876 , \10878 );
or \U$10049 ( \10883 , \10881 , \10882 );
not \U$10050 ( \10884 , \10642 );
not \U$10051 ( \10885 , \10647 );
and \U$10052 ( \10886 , \10884 , \10885 );
and \U$10053 ( \10887 , \10642 , \10647 );
nor \U$10054 ( \10888 , \10886 , \10887 );
xor \U$10055 ( \10889 , \10883 , \10888 );
and \U$10056 ( \10890 , \10568_nR260a , \8981 );
or \U$10057 ( \10891 , \8935 , \10314_nR2685 );
nand \U$10058 ( \10892 , \10891 , \9018 );
nand \U$10059 ( \10893 , \10568_nR260a , \8978 );
and \U$10060 ( \10894 , \10892 , \10893 );
and \U$10061 ( \10895 , \10314_nR2685 , \9022 );
nor \U$10062 ( \10896 , \10890 , \10894 , \10895 );
and \U$10063 ( \10897 , \8825 , RIb55b3b8_580);
and \U$10064 ( \10898 , \8859 , RIb55b688_586);
and \U$10065 ( \10899 , RIb55b610_585, \8844 );
nor \U$10066 ( \10900 , \10898 , \10899 );
and \U$10067 ( \10901 , \8806 , RIb55b160_575);
and \U$10068 ( \10902 , RIb55b0e8_574, \8829 );
nor \U$10069 ( \10903 , \10901 , \10902 );
and \U$10070 ( \10904 , \8816 , RIb55af80_571);
and \U$10071 ( \10905 , RIb55b1d8_576, \8812 );
nor \U$10072 ( \10906 , \10904 , \10905 );
and \U$10073 ( \10907 , \8835 , RIb55b520_583);
and \U$10074 ( \10908 , RIb55b598_584, \8839 );
nor \U$10075 ( \10909 , \10907 , \10908 );
nand \U$10076 ( \10910 , \10900 , \10903 , \10906 , \10909 );
and \U$10077 ( \10911 , \8800 , RIb55b4a8_582);
and \U$10078 ( \10912 , RIb55b430_581, \8823 );
nor \U$10079 ( \10913 , \10911 , \10912 );
not \U$10080 ( \10914 , \10913 );
nor \U$10081 ( \10915 , \10897 , \10910 , \10914 );
and \U$10082 ( \10916 , \8850 , RIb55b2c8_578);
and \U$10083 ( \10917 , RIb55b250_577, \8847 );
nor \U$10084 ( \10918 , \10916 , \10917 );
and \U$10085 ( \10919 , \8831 , RIb55b070_573);
and \U$10086 ( \10920 , RIb55aff8_572, \8853 );
nor \U$10087 ( \10921 , \10919 , \10920 );
and \U$10088 ( \10922 , \8856 , RIb55b700_587);
and \U$10089 ( \10923 , RIb55b340_579, \8818 );
nor \U$10090 ( \10924 , \10922 , \10923 );
nand \U$10091 ( \10925 , \10915 , \10918 , \10921 , \10924 );
_DC r23da ( \10926_nR23da , \10925 , \8863 );
nand \U$10092 ( \10927 , \10926_nR23da , \8768 );
and \U$10093 ( \10928 , \10896 , \10927 );
and \U$10094 ( \10929 , \10686_nR2587 , \8921 );
or \U$10095 ( \10930 , \8877 , \10860_nR251b );
nand \U$10096 ( \10931 , \10930 , \8917 );
nand \U$10097 ( \10932 , \10686_nR2587 , \8912 );
and \U$10098 ( \10933 , \10931 , \10932 );
and \U$10099 ( \10934 , \10860_nR251b , \8914 );
nor \U$10100 ( \10935 , \10929 , \10933 , \10934 );
nor \U$10101 ( \10936 , \10928 , \10935 );
not \U$10102 ( \10937 , \10936 );
nand \U$10103 ( \10938 , \10094_nR289e , \9310 );
or \U$10104 ( \10939 , \9240 , \9899_nR2959 );
nand \U$10105 ( \10940 , \10939 , \9396 );
and \U$10106 ( \10941 , \10938 , \10940 );
and \U$10107 ( \10942 , \9399 , \9899_nR2959 );
and \U$10108 ( \10943 , \10094_nR289e , \9312 );
nor \U$10109 ( \10944 , \10941 , \10942 , \10943 );
nand \U$10110 ( \10945 , \9843_nR2a34 , \9542 );
or \U$10111 ( \10946 , \9411 , \9687_nR2b14 );
nand \U$10112 ( \10947 , \10946 , \9699 );
and \U$10113 ( \10948 , \10945 , \10947 );
and \U$10114 ( \10949 , \9702 , \9687_nR2b14 );
and \U$10115 ( \10950 , \9843_nR2a34 , \9544 );
nor \U$10116 ( \10951 , \10948 , \10949 , \10950 );
xor \U$10117 ( \10952 , \10944 , \10951 );
nand \U$10118 ( \10953 , \10061_nR27cd , \9139 );
or \U$10119 ( \10954 , \9030 , \10347_nR272f );
nand \U$10120 ( \10955 , \10954 , \9144 );
and \U$10121 ( \10956 , \10953 , \10955 );
and \U$10122 ( \10957 , \9141 , \10347_nR272f );
and \U$10123 ( \10958 , \10061_nR27cd , \9224 );
nor \U$10124 ( \10959 , \10956 , \10957 , \10958 );
and \U$10125 ( \10960 , \10952 , \10959 );
and \U$10126 ( \10961 , \10944 , \10951 );
or \U$10127 ( \10962 , \10960 , \10961 );
nand \U$10128 ( \10963 , \10937 , \10962 );
or \U$10129 ( \10964 , \10202 , \10733 );
or \U$10130 ( \10965 , \9177_nR2f04 , \10013 );
or \U$10131 ( \10966 , \9271_nR2e0d , \10012 );
nand \U$10132 ( \10967 , \10964 , \10965 , \10966 );
not \U$10133 ( \10968 , \9462_nR2c1e );
or \U$10134 ( \10969 , \9767 , \10968 );
or \U$10135 ( \10970 , \9717 , \9354_nR2cff );
nand \U$10136 ( \10971 , \10970 , \9946 );
nand \U$10137 ( \10972 , \9462_nR2c1e , \9764 );
and \U$10138 ( \10973 , \10971 , \10972 );
and \U$10139 ( \10974 , \9354_nR2cff , \9949 );
nor \U$10140 ( \10975 , \10973 , \10974 );
nand \U$10141 ( \10976 , \10969 , \10975 );
and \U$10142 ( \10977 , \10967 , \10976 );
and \U$10143 ( \10978 , \10963 , \10977 );
not \U$10144 ( \10979 , \10936 );
nor \U$10145 ( \10980 , \10979 , \10962 );
nor \U$10146 ( \10981 , \10978 , \10980 );
and \U$10147 ( \10982 , \10889 , \10981 );
and \U$10148 ( \10983 , \10883 , \10888 );
or \U$10149 ( \10984 , \10982 , \10983 );
and \U$10150 ( \10985 , \10874 , \10984 );
and \U$10151 ( \10986 , \10871 , \10873 );
or \U$10152 ( \10987 , \10985 , \10986 );
nor \U$10153 ( \10988 , \10822 , \10987 );
xor \U$10154 ( \10989 , \10812 , \10988 );
and \U$10155 ( \10990 , \10822 , \10987 );
nor \U$10156 ( \10991 , \10990 , \10988 );
xor \U$10157 ( \10992 , \10871 , \10873 );
xor \U$10158 ( \10993 , \10992 , \10984 );
xor \U$10159 ( \10994 , \10775 , \10794 );
not \U$10160 ( \10995 , \10994 );
not \U$10161 ( \10996 , \10797 );
and \U$10162 ( \10997 , \10995 , \10996 );
and \U$10163 ( \10998 , \10994 , \10797 );
nor \U$10164 ( \10999 , \10997 , \10998 );
nor \U$10165 ( \11000 , \10993 , \10999 );
xor \U$10166 ( \11001 , \10991 , \11000 );
and \U$10167 ( \11002 , \10993 , \10999 );
nor \U$10168 ( \11003 , \11002 , \11000 );
not \U$10169 ( \11004 , \10827 );
not \U$10170 ( \11005 , \10870 );
and \U$10171 ( \11006 , \11004 , \11005 );
and \U$10172 ( \11007 , \10827 , \10870 );
nor \U$10173 ( \11008 , \11006 , \11007 );
xor \U$10174 ( \11009 , \10883 , \10888 );
xor \U$10175 ( \11010 , \11009 , \10981 );
and \U$10176 ( \11011 , \11008 , \11010 );
xor \U$10177 ( \11012 , \10876 , \10878 );
xor \U$10178 ( \11013 , \11012 , \10880 );
nand \U$10179 ( \11014 , \10347_nR272f , \9139 );
or \U$10180 ( \11015 , \9030 , \10314_nR2685 );
nand \U$10181 ( \11016 , \11015 , \9144 );
and \U$10182 ( \11017 , \11014 , \11016 );
and \U$10183 ( \11018 , \9141 , \10314_nR2685 );
and \U$10184 ( \11019 , \10347_nR272f , \9224 );
nor \U$10185 ( \11020 , \11017 , \11018 , \11019 );
nand \U$10186 ( \11021 , \10061_nR27cd , \9310 );
or \U$10187 ( \11022 , \9240 , \10094_nR289e );
nand \U$10188 ( \11023 , \11022 , \9396 );
and \U$10189 ( \11024 , \11021 , \11023 );
and \U$10190 ( \11025 , \9399 , \10094_nR289e );
and \U$10191 ( \11026 , \10061_nR27cd , \9312 );
nor \U$10192 ( \11027 , \11024 , \11025 , \11026 );
xor \U$10193 ( \11028 , \11020 , \11027 );
and \U$10194 ( \11029 , \10686_nR2587 , \8981 );
or \U$10195 ( \11030 , \8935 , \10568_nR260a );
nand \U$10196 ( \11031 , \11030 , \9018 );
nand \U$10197 ( \11032 , \10686_nR2587 , \8978 );
and \U$10198 ( \11033 , \11031 , \11032 );
and \U$10199 ( \11034 , \10568_nR260a , \9022 );
nor \U$10200 ( \11035 , \11029 , \11033 , \11034 );
and \U$10201 ( \11036 , \11028 , \11035 );
and \U$10202 ( \11037 , \11020 , \11027 );
or \U$10203 ( \11038 , \11036 , \11037 );
nand \U$10204 ( \11039 , \9687_nR2b14 , \9764 );
or \U$10205 ( \11040 , \9717 , \9462_nR2c1e );
nand \U$10206 ( \11041 , \11040 , \9946 );
and \U$10207 ( \11042 , \11039 , \11041 );
and \U$10208 ( \11043 , \9949 , \9462_nR2c1e );
and \U$10209 ( \11044 , \9687_nR2b14 , \9766 );
nor \U$10210 ( \11045 , \11042 , \11043 , \11044 );
and \U$10211 ( \11046 , \9272 , \10199 );
not \U$10212 ( \11047 , \9354_nR2cff );
and \U$10213 ( \11048 , \10011 , \11047 );
and \U$10214 ( \11049 , \9271_nR2e0d , \10203 );
nor \U$10215 ( \11050 , \11046 , \11048 , \11049 );
xor \U$10216 ( \11051 , \11045 , \11050 );
nand \U$10217 ( \11052 , \9899_nR2959 , \9542 );
or \U$10218 ( \11053 , \9411 , \9843_nR2a34 );
nand \U$10219 ( \11054 , \11053 , \9699 );
and \U$10220 ( \11055 , \11052 , \11054 );
and \U$10221 ( \11056 , \9702 , \9843_nR2a34 );
and \U$10222 ( \11057 , \9899_nR2959 , \9544 );
nor \U$10223 ( \11058 , \11055 , \11056 , \11057 );
and \U$10224 ( \11059 , \11051 , \11058 );
and \U$10225 ( \11060 , \11045 , \11050 );
or \U$10226 ( \11061 , \11059 , \11060 );
xor \U$10227 ( \11062 , \11038 , \11061 );
not \U$10228 ( \11063 , \10935 );
not \U$10229 ( \11064 , \10896 );
and \U$10230 ( \11065 , \11063 , \11064 );
and \U$10231 ( \11066 , \10935 , \10896 );
nor \U$10232 ( \11067 , \11065 , \11066 );
not \U$10233 ( \11068 , \11067 );
not \U$10234 ( \11069 , \10927 );
and \U$10235 ( \11070 , \11068 , \11069 );
and \U$10236 ( \11071 , \11067 , \10927 );
nor \U$10237 ( \11072 , \11070 , \11071 );
and \U$10238 ( \11073 , \11062 , \11072 );
and \U$10239 ( \11074 , \11038 , \11061 );
or \U$10240 ( \11075 , \11073 , \11074 );
nand \U$10241 ( \11076 , \11013 , \11075 );
xor \U$10242 ( \11077 , \10967 , \10976 );
not \U$10243 ( \11078 , \11077 );
xor \U$10244 ( \11079 , \10944 , \10951 );
xor \U$10245 ( \11080 , \11079 , \10959 );
nor \U$10246 ( \11081 , \11078 , \11080 );
and \U$10247 ( \11082 , \11076 , \11081 );
nor \U$10248 ( \11083 , \11075 , \11013 );
nor \U$10249 ( \11084 , \11082 , \11083 );
xor \U$10250 ( \11085 , \10883 , \10888 );
xor \U$10251 ( \11086 , \11085 , \10981 );
and \U$10252 ( \11087 , \11084 , \11086 );
and \U$10253 ( \11088 , \11008 , \11084 );
or \U$10254 ( \11089 , \11011 , \11087 , \11088 );
not \U$10255 ( \11090 , \11089 );
xor \U$10256 ( \11091 , \11003 , \11090 );
not \U$10257 ( \11092 , \11081 );
not \U$10258 ( \11093 , \11083 );
nand \U$10259 ( \11094 , \11093 , \11076 );
not \U$10260 ( \11095 , \11094 );
or \U$10261 ( \11096 , \11092 , \11095 );
or \U$10262 ( \11097 , \11094 , \11081 );
nand \U$10263 ( \11098 , \11096 , \11097 );
not \U$10264 ( \11099 , \10977 );
not \U$10265 ( \11100 , \10980 );
nand \U$10266 ( \11101 , \11100 , \10963 );
not \U$10267 ( \11102 , \11101 );
or \U$10268 ( \11103 , \11099 , \11102 );
or \U$10269 ( \11104 , \11101 , \10977 );
nand \U$10270 ( \11105 , \11103 , \11104 );
nor \U$10271 ( \11106 , \11098 , \11105 );
nand \U$10272 ( \11107 , \9843_nR2a34 , \9764 );
or \U$10273 ( \11108 , \9717 , \9687_nR2b14 );
nand \U$10274 ( \11109 , \11108 , \9946 );
and \U$10275 ( \11110 , \11107 , \11109 );
and \U$10276 ( \11111 , \9949 , \9687_nR2b14 );
and \U$10277 ( \11112 , \9843_nR2a34 , \9766 );
nor \U$10278 ( \11113 , \11110 , \11111 , \11112 );
and \U$10279 ( \11114 , \11047 , \10199 );
and \U$10280 ( \11115 , \10011 , \10968 );
and \U$10281 ( \11116 , \9354_nR2cff , \10203 );
nor \U$10282 ( \11117 , \11114 , \11115 , \11116 );
xor \U$10283 ( \11118 , \11113 , \11117 );
and \U$10284 ( \11119 , \11118 , \8877 );
and \U$10285 ( \11120 , \11113 , \11117 );
or \U$10286 ( \11121 , \11119 , \11120 );
nand \U$10287 ( \11122 , \10347_nR272f , \9310 );
or \U$10288 ( \11123 , \9240 , \10061_nR27cd );
nand \U$10289 ( \11124 , \11123 , \9396 );
and \U$10290 ( \11125 , \11122 , \11124 );
and \U$10291 ( \11126 , \9399 , \10061_nR27cd );
and \U$10292 ( \11127 , \10347_nR272f , \9312 );
nor \U$10293 ( \11128 , \11125 , \11126 , \11127 );
nand \U$10294 ( \11129 , \10094_nR289e , \9542 );
or \U$10295 ( \11130 , \9411 , \9899_nR2959 );
nand \U$10296 ( \11131 , \11130 , \9699 );
and \U$10297 ( \11132 , \11129 , \11131 );
and \U$10298 ( \11133 , \9702 , \9899_nR2959 );
and \U$10299 ( \11134 , \10094_nR289e , \9544 );
nor \U$10300 ( \11135 , \11132 , \11133 , \11134 );
xor \U$10301 ( \11136 , \11128 , \11135 );
nand \U$10302 ( \11137 , \10314_nR2685 , \9139 );
or \U$10303 ( \11138 , \9030 , \10568_nR260a );
nand \U$10304 ( \11139 , \11138 , \9144 );
and \U$10305 ( \11140 , \11137 , \11139 );
and \U$10306 ( \11141 , \9141 , \10568_nR260a );
and \U$10307 ( \11142 , \10314_nR2685 , \9224 );
nor \U$10308 ( \11143 , \11140 , \11141 , \11142 );
and \U$10309 ( \11144 , \11136 , \11143 );
and \U$10310 ( \11145 , \11128 , \11135 );
or \U$10311 ( \11146 , \11144 , \11145 );
xor \U$10312 ( \11147 , \11121 , \11146 );
and \U$10313 ( \11148 , \10860_nR251b , \8921 );
or \U$10314 ( \11149 , \8877 , \10926_nR23da );
nand \U$10315 ( \11150 , \11149 , \8917 );
nand \U$10316 ( \11151 , \10860_nR251b , \8912 );
and \U$10317 ( \11152 , \11150 , \11151 );
and \U$10318 ( \11153 , \10926_nR23da , \8914 );
nor \U$10319 ( \11154 , \11148 , \11152 , \11153 );
and \U$10320 ( \11155 , \11147 , \11154 );
and \U$10321 ( \11156 , \11121 , \11146 );
or \U$10322 ( \11157 , \11155 , \11156 );
not \U$10323 ( \11158 , \11080 );
not \U$10324 ( \11159 , \11077 );
and \U$10325 ( \11160 , \11158 , \11159 );
and \U$10326 ( \11161 , \11080 , \11077 );
nor \U$10327 ( \11162 , \11160 , \11161 );
xor \U$10328 ( \11163 , \11157 , \11162 );
xor \U$10329 ( \11164 , \11038 , \11061 );
xor \U$10330 ( \11165 , \11164 , \11072 );
and \U$10331 ( \11166 , \11163 , \11165 );
and \U$10332 ( \11167 , \11157 , \11162 );
or \U$10333 ( \11168 , \11166 , \11167 );
or \U$10334 ( \11169 , \11106 , \11168 );
nand \U$10335 ( \11170 , \11105 , \11098 );
nand \U$10336 ( \11171 , \11169 , \11170 );
xor \U$10337 ( \11172 , \10883 , \10888 );
xor \U$10338 ( \11173 , \11172 , \10981 );
xor \U$10339 ( \11174 , \11008 , \11084 );
xor \U$10340 ( \11175 , \11173 , \11174 );
not \U$10341 ( \11176 , \11175 );
xor \U$10342 ( \11177 , \11171 , \11176 );
not \U$10343 ( \11178 , \11168 );
not \U$10344 ( \11179 , \11106 );
nand \U$10345 ( \11180 , \11179 , \11170 );
not \U$10346 ( \11181 , \11180 );
or \U$10347 ( \11182 , \11178 , \11181 );
or \U$10348 ( \11183 , \11180 , \11168 );
nand \U$10349 ( \11184 , \11182 , \11183 );
xor \U$10350 ( \11185 , \11121 , \11146 );
xor \U$10351 ( \11186 , \11185 , \11154 );
xor \U$10352 ( \11187 , \11045 , \11050 );
xor \U$10353 ( \11188 , \11187 , \11058 );
or \U$10354 ( \11189 , \11186 , \11188 );
and \U$10355 ( \11190 , \10860_nR251b , \8981 );
or \U$10356 ( \11191 , \8935 , \10686_nR2587 );
nand \U$10357 ( \11192 , \11191 , \9018 );
nand \U$10358 ( \11193 , \10860_nR251b , \8978 );
and \U$10359 ( \11194 , \11192 , \11193 );
and \U$10360 ( \11195 , \10686_nR2587 , \9022 );
nor \U$10361 ( \11196 , \11190 , \11194 , \11195 );
nand \U$10362 ( \11197 , \9899_nR2959 , \9764 );
or \U$10363 ( \11198 , \9717 , \9843_nR2a34 );
nand \U$10364 ( \11199 , \11198 , \9946 );
and \U$10365 ( \11200 , \11197 , \11199 );
and \U$10366 ( \11201 , \9949 , \9843_nR2a34 );
and \U$10367 ( \11202 , \9899_nR2959 , \9766 );
nor \U$10368 ( \11203 , \11200 , \11201 , \11202 );
and \U$10369 ( \11204 , \10968 , \10199 );
and \U$10370 ( \11205 , \10011 , \9755 );
and \U$10371 ( \11206 , \9462_nR2c1e , \10203 );
nor \U$10372 ( \11207 , \11204 , \11205 , \11206 );
xor \U$10373 ( \11208 , \11203 , \11207 );
nand \U$10374 ( \11209 , \10061_nR27cd , \9542 );
or \U$10375 ( \11210 , \9411 , \10094_nR289e );
nand \U$10376 ( \11211 , \11210 , \9699 );
and \U$10377 ( \11212 , \11209 , \11211 );
and \U$10378 ( \11213 , \9702 , \10094_nR289e );
and \U$10379 ( \11214 , \10061_nR27cd , \9544 );
nor \U$10380 ( \11215 , \11212 , \11213 , \11214 );
and \U$10381 ( \11216 , \11208 , \11215 );
and \U$10382 ( \11217 , \11203 , \11207 );
or \U$10383 ( \11218 , \11216 , \11217 );
xor \U$10384 ( \11219 , \11196 , \11218 );
nand \U$10385 ( \11220 , \10568_nR260a , \9139 );
or \U$10386 ( \11221 , \9030 , \10686_nR2587 );
nand \U$10387 ( \11222 , \11221 , \9144 );
and \U$10388 ( \11223 , \11220 , \11222 );
and \U$10389 ( \11224 , \9141 , \10686_nR2587 );
and \U$10390 ( \11225 , \10568_nR260a , \9224 );
nor \U$10391 ( \11226 , \11223 , \11224 , \11225 );
nand \U$10392 ( \11227 , \10314_nR2685 , \9310 );
or \U$10393 ( \11228 , \9240 , \10347_nR272f );
nand \U$10394 ( \11229 , \11228 , \9396 );
and \U$10395 ( \11230 , \11227 , \11229 );
and \U$10396 ( \11231 , \9399 , \10347_nR272f );
and \U$10397 ( \11232 , \10314_nR2685 , \9312 );
nor \U$10398 ( \11233 , \11230 , \11231 , \11232 );
xor \U$10399 ( \11234 , \11226 , \11233 );
and \U$10400 ( \11235 , \10926_nR23da , \8981 );
or \U$10401 ( \11236 , \8935 , \10860_nR251b );
nand \U$10402 ( \11237 , \11236 , \9018 );
nand \U$10403 ( \11238 , \10926_nR23da , \8978 );
and \U$10404 ( \11239 , \11237 , \11238 );
and \U$10405 ( \11240 , \10860_nR251b , \9022 );
nor \U$10406 ( \11241 , \11235 , \11239 , \11240 );
and \U$10407 ( \11242 , \11234 , \11241 );
and \U$10408 ( \11243 , \11226 , \11233 );
or \U$10409 ( \11244 , \11242 , \11243 );
and \U$10410 ( \11245 , \11219 , \11244 );
and \U$10411 ( \11246 , \11196 , \11218 );
or \U$10412 ( \11247 , \11245 , \11246 );
xor \U$10413 ( \11248 , \11020 , \11027 );
xor \U$10414 ( \11249 , \11248 , \11035 );
xor \U$10415 ( \11250 , \11247 , \11249 );
xor \U$10416 ( \11251 , \11113 , \11117 );
xor \U$10417 ( \11252 , \11251 , \8877 );
xor \U$10418 ( \11253 , \11128 , \11135 );
xor \U$10419 ( \11254 , \11253 , \11143 );
xor \U$10420 ( \11255 , \11252 , \11254 );
nand \U$10421 ( \11256 , \10926_nR23da , \8912 );
and \U$10422 ( \11257 , \8876 , \11256 );
and \U$10423 ( \11258 , \10926_nR23da , \8921 );
nor \U$10424 ( \11259 , \11257 , \11258 );
and \U$10425 ( \11260 , \11255 , \11259 );
and \U$10426 ( \11261 , \11252 , \11254 );
or \U$10427 ( \11262 , \11260 , \11261 );
and \U$10428 ( \11263 , \11250 , \11262 );
and \U$10429 ( \11264 , \11247 , \11249 );
or \U$10430 ( \11265 , \11263 , \11264 );
xor \U$10431 ( \11266 , \11189 , \11265 );
xor \U$10432 ( \11267 , \11157 , \11162 );
xor \U$10433 ( \11268 , \11267 , \11165 );
and \U$10434 ( \11269 , \11266 , \11268 );
and \U$10435 ( \11270 , \11189 , \11265 );
or \U$10436 ( \11271 , \11269 , \11270 );
xor \U$10437 ( \11272 , \11184 , \11271 );
xor \U$10438 ( \11273 , \11247 , \11249 );
xor \U$10439 ( \11274 , \11273 , \11262 );
xor \U$10440 ( \11275 , \11196 , \11218 );
xor \U$10441 ( \11276 , \11275 , \11244 );
xor \U$10442 ( \11277 , \11252 , \11254 );
xor \U$10443 ( \11278 , \11277 , \11259 );
and \U$10444 ( \11279 , \11276 , \11278 );
nand \U$10445 ( \11280 , \10568_nR260a , \9310 );
or \U$10446 ( \11281 , \9240 , \10314_nR2685 );
nand \U$10447 ( \11282 , \11281 , \9396 );
and \U$10448 ( \11283 , \11280 , \11282 );
and \U$10449 ( \11284 , \9399 , \10314_nR2685 );
and \U$10450 ( \11285 , \10568_nR260a , \9312 );
nor \U$10451 ( \11286 , \11283 , \11284 , \11285 );
nand \U$10452 ( \11287 , \10347_nR272f , \9542 );
or \U$10453 ( \11288 , \9411 , \10061_nR27cd );
nand \U$10454 ( \11289 , \11288 , \9699 );
and \U$10455 ( \11290 , \11287 , \11289 );
and \U$10456 ( \11291 , \9702 , \10061_nR27cd );
and \U$10457 ( \11292 , \10347_nR272f , \9544 );
nor \U$10458 ( \11293 , \11290 , \11291 , \11292 );
xor \U$10459 ( \11294 , \11286 , \11293 );
nand \U$10460 ( \11295 , \10686_nR2587 , \9139 );
or \U$10461 ( \11296 , \9030 , \10860_nR251b );
nand \U$10462 ( \11297 , \11296 , \9144 );
and \U$10463 ( \11298 , \11295 , \11297 );
and \U$10464 ( \11299 , \9141 , \10860_nR251b );
and \U$10465 ( \11300 , \10686_nR2587 , \9224 );
nor \U$10466 ( \11301 , \11298 , \11299 , \11300 );
and \U$10467 ( \11302 , \11294 , \11301 );
and \U$10468 ( \11303 , \11286 , \11293 );
or \U$10469 ( \11304 , \11302 , \11303 );
nand \U$10470 ( \11305 , \10094_nR289e , \9764 );
or \U$10471 ( \11306 , \9717 , \9899_nR2959 );
nand \U$10472 ( \11307 , \11306 , \9946 );
and \U$10473 ( \11308 , \11305 , \11307 );
and \U$10474 ( \11309 , \9949 , \9899_nR2959 );
and \U$10475 ( \11310 , \10094_nR289e , \9766 );
nor \U$10476 ( \11311 , \11308 , \11309 , \11310 );
and \U$10477 ( \11312 , \9755 , \10199 );
not \U$10478 ( \11313 , \9843_nR2a34 );
and \U$10479 ( \11314 , \10011 , \11313 );
and \U$10480 ( \11315 , \9687_nR2b14 , \10203 );
nor \U$10481 ( \11316 , \11312 , \11314 , \11315 );
xor \U$10482 ( \11317 , \11311 , \11316 );
and \U$10483 ( \11318 , \11317 , \8935 );
and \U$10484 ( \11319 , \11311 , \11316 );
or \U$10485 ( \11320 , \11318 , \11319 );
xor \U$10486 ( \11321 , \11304 , \11320 );
xor \U$10487 ( \11322 , \11226 , \11233 );
xor \U$10488 ( \11323 , \11322 , \11241 );
and \U$10489 ( \11324 , \11321 , \11323 );
and \U$10490 ( \11325 , \11304 , \11320 );
or \U$10491 ( \11326 , \11324 , \11325 );
xor \U$10492 ( \11327 , \11252 , \11254 );
xor \U$10493 ( \11328 , \11327 , \11259 );
and \U$10494 ( \11329 , \11326 , \11328 );
and \U$10495 ( \11330 , \11276 , \11326 );
or \U$10496 ( \11331 , \11279 , \11329 , \11330 );
xnor \U$10497 ( \11332 , \11188 , \11186 );
xor \U$10498 ( \11333 , \11331 , \11332 );
xor \U$10499 ( \11334 , \11274 , \11333 );
not \U$10500 ( \11335 , \11334 );
xor \U$10501 ( \11336 , \11252 , \11254 );
xor \U$10502 ( \11337 , \11336 , \11259 );
xor \U$10503 ( \11338 , \11276 , \11326 );
xor \U$10504 ( \11339 , \11337 , \11338 );
not \U$10505 ( \11340 , \10926_nR23da );
and \U$10506 ( \11341 , \11340 , \8980 );
and \U$10507 ( \11342 , \10926_nR23da , \9022 );
not \U$10508 ( \11343 , \9018 );
nor \U$10509 ( \11344 , \11341 , \11342 , \11343 );
nand \U$10510 ( \11345 , \10061_nR27cd , \9764 );
or \U$10511 ( \11346 , \9717 , \10094_nR289e );
nand \U$10512 ( \11347 , \11346 , \9946 );
and \U$10513 ( \11348 , \11345 , \11347 );
and \U$10514 ( \11349 , \9949 , \10094_nR289e );
and \U$10515 ( \11350 , \10061_nR27cd , \9766 );
nor \U$10516 ( \11351 , \11348 , \11349 , \11350 );
not \U$10517 ( \11352 , \11351 );
and \U$10518 ( \11353 , \11313 , \10199 );
not \U$10519 ( \11354 , \9899_nR2959 );
and \U$10520 ( \11355 , \10011 , \11354 );
and \U$10521 ( \11356 , \9843_nR2a34 , \10203 );
nor \U$10522 ( \11357 , \11353 , \11355 , \11356 );
not \U$10523 ( \11358 , \11357 );
and \U$10524 ( \11359 , \11352 , \11358 );
and \U$10525 ( \11360 , \11351 , \11357 );
nand \U$10526 ( \11361 , \10314_nR2685 , \9542 );
or \U$10527 ( \11362 , \9411 , \10347_nR272f );
nand \U$10528 ( \11363 , \11362 , \9699 );
and \U$10529 ( \11364 , \11361 , \11363 );
and \U$10530 ( \11365 , \9702 , \10347_nR272f );
and \U$10531 ( \11366 , \10314_nR2685 , \9544 );
nor \U$10532 ( \11367 , \11364 , \11365 , \11366 );
nor \U$10533 ( \11368 , \11360 , \11367 );
nor \U$10534 ( \11369 , \11359 , \11368 );
and \U$10535 ( \11370 , \11344 , \11369 );
not \U$10536 ( \11371 , \11370 );
xor \U$10537 ( \11372 , \11286 , \11293 );
xor \U$10538 ( \11373 , \11372 , \11301 );
not \U$10539 ( \11374 , \11373 );
and \U$10540 ( \11375 , \11371 , \11374 );
nor \U$10541 ( \11376 , \11344 , \11369 );
nor \U$10542 ( \11377 , \11375 , \11376 );
xor \U$10543 ( \11378 , \11203 , \11207 );
xor \U$10544 ( \11379 , \11378 , \11215 );
xor \U$10545 ( \11380 , \11377 , \11379 );
xor \U$10546 ( \11381 , \11304 , \11320 );
xor \U$10547 ( \11382 , \11381 , \11323 );
and \U$10548 ( \11383 , \11380 , \11382 );
and \U$10549 ( \11384 , \11377 , \11379 );
or \U$10550 ( \11385 , \11383 , \11384 );
nor \U$10551 ( \11386 , \11339 , \11385 );
xor \U$10552 ( \11387 , \11335 , \11386 );
and \U$10553 ( \11388 , \11339 , \11385 );
nor \U$10554 ( \11389 , \11388 , \11386 );
xor \U$10555 ( \11390 , \11377 , \11379 );
xor \U$10556 ( \11391 , \11390 , \11382 );
nand \U$10557 ( \11392 , \10347_nR272f , \9764 );
or \U$10558 ( \11393 , \9717 , \10061_nR27cd );
nand \U$10559 ( \11394 , \11393 , \9946 );
and \U$10560 ( \11395 , \11392 , \11394 );
and \U$10561 ( \11396 , \9949 , \10061_nR27cd );
and \U$10562 ( \11397 , \10347_nR272f , \9766 );
nor \U$10563 ( \11398 , \11395 , \11396 , \11397 );
and \U$10564 ( \11399 , \11354 , \10199 );
not \U$10565 ( \11400 , \10094_nR289e );
and \U$10566 ( \11401 , \10011 , \11400 );
and \U$10567 ( \11402 , \9899_nR2959 , \10203 );
nor \U$10568 ( \11403 , \11399 , \11401 , \11402 );
xor \U$10569 ( \11404 , \11398 , \11403 );
and \U$10570 ( \11405 , \11404 , \9030 );
and \U$10571 ( \11406 , \11398 , \11403 );
or \U$10572 ( \11407 , \11405 , \11406 );
nand \U$10573 ( \11408 , \10686_nR2587 , \9310 );
or \U$10574 ( \11409 , \9240 , \10568_nR260a );
nand \U$10575 ( \11410 , \11409 , \9396 );
and \U$10576 ( \11411 , \11408 , \11410 );
and \U$10577 ( \11412 , \9399 , \10568_nR260a );
and \U$10578 ( \11413 , \10686_nR2587 , \9312 );
nor \U$10579 ( \11414 , \11411 , \11412 , \11413 );
xor \U$10580 ( \11415 , \11407 , \11414 );
nand \U$10581 ( \11416 , \10860_nR251b , \9310 );
or \U$10582 ( \11417 , \9240 , \10686_nR2587 );
nand \U$10583 ( \11418 , \11417 , \9396 );
and \U$10584 ( \11419 , \11416 , \11418 );
and \U$10585 ( \11420 , \9399 , \10686_nR2587 );
and \U$10586 ( \11421 , \10860_nR251b , \9312 );
nor \U$10587 ( \11422 , \11419 , \11420 , \11421 );
nand \U$10588 ( \11423 , \10568_nR260a , \9542 );
or \U$10589 ( \11424 , \9411 , \10314_nR2685 );
nand \U$10590 ( \11425 , \11424 , \9699 );
and \U$10591 ( \11426 , \11423 , \11425 );
and \U$10592 ( \11427 , \9702 , \10314_nR2685 );
and \U$10593 ( \11428 , \10568_nR260a , \9544 );
nor \U$10594 ( \11429 , \11426 , \11427 , \11428 );
xor \U$10595 ( \11430 , \11422 , \11429 );
and \U$10596 ( \11431 , \9224 , \10926_nR23da );
nand \U$10597 ( \11432 , \10926_nR23da , \9139 );
and \U$10598 ( \11433 , \11432 , \9031 );
nor \U$10599 ( \11434 , \11431 , \11433 );
and \U$10600 ( \11435 , \11430 , \11434 );
and \U$10601 ( \11436 , \11422 , \11429 );
or \U$10602 ( \11437 , \11435 , \11436 );
and \U$10603 ( \11438 , \11415 , \11437 );
and \U$10604 ( \11439 , \11407 , \11414 );
or \U$10605 ( \11440 , \11438 , \11439 );
xor \U$10606 ( \11441 , \11311 , \11316 );
xor \U$10607 ( \11442 , \11441 , \8935 );
nand \U$10608 ( \11443 , \11440 , \11442 );
not \U$10609 ( \11444 , \11351 );
xor \U$10610 ( \11445 , \11357 , \11367 );
not \U$10611 ( \11446 , \11445 );
or \U$10612 ( \11447 , \11444 , \11446 );
or \U$10613 ( \11448 , \11445 , \11351 );
nand \U$10614 ( \11449 , \11447 , \11448 );
not \U$10615 ( \11450 , \10860_nR251b );
or \U$10616 ( \11451 , \9293 , \11450 );
or \U$10617 ( \11452 , \11340 , \9295 );
or \U$10618 ( \11453 , \9223 , \11450 );
or \U$10619 ( \11454 , \9030 , \10926_nR23da );
nand \U$10620 ( \11455 , \11454 , \9144 );
nand \U$10621 ( \11456 , \11453 , \11455 );
nand \U$10622 ( \11457 , \11451 , \11452 , \11456 );
and \U$10623 ( \11458 , \11449 , \11457 );
and \U$10624 ( \11459 , \11443 , \11458 );
nor \U$10625 ( \11460 , \11440 , \11442 );
nor \U$10626 ( \11461 , \11459 , \11460 );
nor \U$10627 ( \11462 , \11391 , \11461 );
xor \U$10628 ( \11463 , \11389 , \11462 );
not \U$10629 ( \11464 , \11458 );
not \U$10630 ( \11465 , \11460 );
nand \U$10631 ( \11466 , \11465 , \11443 );
not \U$10632 ( \11467 , \11466 );
or \U$10633 ( \11468 , \11464 , \11467 );
or \U$10634 ( \11469 , \11466 , \11458 );
nand \U$10635 ( \11470 , \11468 , \11469 );
not \U$10636 ( \11471 , \11373 );
nor \U$10637 ( \11472 , \11376 , \11370 );
not \U$10638 ( \11473 , \11472 );
or \U$10639 ( \11474 , \11471 , \11473 );
or \U$10640 ( \11475 , \11472 , \11373 );
nand \U$10641 ( \11476 , \11474 , \11475 );
xor \U$10642 ( \11477 , \11470 , \11476 );
xor \U$10643 ( \11478 , \11407 , \11414 );
xor \U$10644 ( \11479 , \11478 , \11437 );
nand \U$10645 ( \11480 , \10314_nR2685 , \9764 );
or \U$10646 ( \11481 , \9717 , \10347_nR272f );
nand \U$10647 ( \11482 , \11481 , \9946 );
and \U$10648 ( \11483 , \11480 , \11482 );
and \U$10649 ( \11484 , \9949 , \10347_nR272f );
and \U$10650 ( \11485 , \10314_nR2685 , \9766 );
nor \U$10651 ( \11486 , \11483 , \11484 , \11485 );
and \U$10652 ( \11487 , \11400 , \10199 );
not \U$10653 ( \11488 , \10061_nR27cd );
and \U$10654 ( \11489 , \10011 , \11488 );
and \U$10655 ( \11490 , \10094_nR289e , \10203 );
nor \U$10656 ( \11491 , \11487 , \11489 , \11490 );
xor \U$10657 ( \11492 , \11486 , \11491 );
nand \U$10658 ( \11493 , \10686_nR2587 , \9542 );
or \U$10659 ( \11494 , \9411 , \10568_nR260a );
nand \U$10660 ( \11495 , \11494 , \9699 );
and \U$10661 ( \11496 , \11493 , \11495 );
and \U$10662 ( \11497 , \9702 , \10568_nR260a );
and \U$10663 ( \11498 , \10686_nR2587 , \9544 );
nor \U$10664 ( \11499 , \11496 , \11497 , \11498 );
and \U$10665 ( \11500 , \11492 , \11499 );
and \U$10666 ( \11501 , \11486 , \11491 );
or \U$10667 ( \11502 , \11500 , \11501 );
xor \U$10668 ( \11503 , \11398 , \11403 );
xor \U$10669 ( \11504 , \11503 , \9030 );
and \U$10670 ( \11505 , \11502 , \11504 );
xor \U$10671 ( \11506 , \11422 , \11429 );
xor \U$10672 ( \11507 , \11506 , \11434 );
xor \U$10673 ( \11508 , \11398 , \11403 );
xor \U$10674 ( \11509 , \11508 , \9030 );
and \U$10675 ( \11510 , \11507 , \11509 );
and \U$10676 ( \11511 , \11502 , \11507 );
or \U$10677 ( \11512 , \11505 , \11510 , \11511 );
nand \U$10678 ( \11513 , \11479 , \11512 );
xor \U$10679 ( \11514 , \11449 , \11457 );
and \U$10680 ( \11515 , \11513 , \11514 );
nor \U$10681 ( \11516 , \11512 , \11479 );
nor \U$10682 ( \11517 , \11515 , \11516 );
not \U$10683 ( \11518 , \11517 );
xor \U$10684 ( \11519 , \11477 , \11518 );
not \U$10685 ( \11520 , \11513 );
nor \U$10686 ( \11521 , \11520 , \11516 );
not \U$10687 ( \11522 , \11521 );
not \U$10688 ( \11523 , \11514 );
and \U$10689 ( \11524 , \11522 , \11523 );
and \U$10690 ( \11525 , \11521 , \11514 );
nor \U$10691 ( \11526 , \11524 , \11525 );
xor \U$10692 ( \11527 , \11398 , \11403 );
xor \U$10693 ( \11528 , \11527 , \9030 );
xor \U$10694 ( \11529 , \11502 , \11507 );
xor \U$10695 ( \11530 , \11528 , \11529 );
nand \U$10696 ( \11531 , \10926_nR23da , \9310 );
or \U$10697 ( \11532 , \9240 , \10860_nR251b );
nand \U$10698 ( \11533 , \11532 , \9396 );
and \U$10699 ( \11534 , \11531 , \11533 );
and \U$10700 ( \11535 , \9399 , \10860_nR251b );
and \U$10701 ( \11536 , \10926_nR23da , \9312 );
nor \U$10702 ( \11537 , \11534 , \11535 , \11536 );
and \U$10703 ( \11538 , \11488 , \10199 );
not \U$10704 ( \11539 , \10347_nR272f );
and \U$10705 ( \11540 , \10011 , \11539 );
and \U$10706 ( \11541 , \10061_nR27cd , \10203 );
nor \U$10707 ( \11542 , \11538 , \11540 , \11541 );
and \U$10708 ( \11543 , \9240 , \11542 );
not \U$10709 ( \11544 , \11543 );
nand \U$10710 ( \11545 , \10568_nR260a , \9764 );
or \U$10711 ( \11546 , \9717 , \10314_nR2685 );
nand \U$10712 ( \11547 , \11546 , \9946 );
and \U$10713 ( \11548 , \11545 , \11547 );
and \U$10714 ( \11549 , \9949 , \10314_nR2685 );
and \U$10715 ( \11550 , \10568_nR260a , \9766 );
nor \U$10716 ( \11551 , \11548 , \11549 , \11550 );
not \U$10717 ( \11552 , \11551 );
and \U$10718 ( \11553 , \11544 , \11552 );
nor \U$10719 ( \11554 , \9240 , \11542 );
nor \U$10720 ( \11555 , \11553 , \11554 );
xor \U$10721 ( \11556 , \11537 , \11555 );
nand \U$10722 ( \11557 , \10860_nR251b , \9542 );
or \U$10723 ( \11558 , \9411 , \10686_nR2587 );
nand \U$10724 ( \11559 , \11558 , \9699 );
and \U$10725 ( \11560 , \11557 , \11559 );
and \U$10726 ( \11561 , \9702 , \10686_nR2587 );
and \U$10727 ( \11562 , \10860_nR251b , \9544 );
nor \U$10728 ( \11563 , \11560 , \11561 , \11562 );
not \U$10729 ( \11564 , \11563 );
or \U$10730 ( \11565 , \9552 , \11340 );
or \U$10731 ( \11566 , \10926_nR23da , \9240 );
nand \U$10732 ( \11567 , \11565 , \11566 , \9396 );
nand \U$10733 ( \11568 , \11564 , \11567 );
and \U$10734 ( \11569 , \11556 , \11568 );
and \U$10735 ( \11570 , \11537 , \11555 );
or \U$10736 ( \11571 , \11569 , \11570 );
nor \U$10737 ( \11572 , \11530 , \11571 );
xor \U$10738 ( \11573 , \11526 , \11572 );
xor \U$10739 ( \11574 , \11537 , \11555 );
xor \U$10740 ( \11575 , \11574 , \11568 );
xor \U$10741 ( \11576 , \11486 , \11491 );
xor \U$10742 ( \11577 , \11576 , \11499 );
and \U$10743 ( \11578 , \11575 , \11577 );
nor \U$10744 ( \11579 , \11575 , \11577 );
nor \U$10745 ( \11580 , \11578 , \11579 );
not \U$10746 ( \11581 , \11551 );
nor \U$10747 ( \11582 , \11543 , \11554 );
not \U$10748 ( \11583 , \11582 );
or \U$10749 ( \11584 , \11581 , \11583 );
or \U$10750 ( \11585 , \11582 , \11551 );
nand \U$10751 ( \11586 , \11584 , \11585 );
nand \U$10752 ( \11587 , \10686_nR2587 , \9764 );
or \U$10753 ( \11588 , \9717 , \10568_nR260a );
nand \U$10754 ( \11589 , \11588 , \9946 );
and \U$10755 ( \11590 , \11587 , \11589 );
and \U$10756 ( \11591 , \9949 , \10568_nR260a );
and \U$10757 ( \11592 , \10686_nR2587 , \9766 );
nor \U$10758 ( \11593 , \11590 , \11591 , \11592 );
and \U$10759 ( \11594 , \11539 , \10199 );
not \U$10760 ( \11595 , \10314_nR2685 );
and \U$10761 ( \11596 , \10011 , \11595 );
and \U$10762 ( \11597 , \10347_nR272f , \10203 );
nor \U$10763 ( \11598 , \11594 , \11596 , \11597 );
or \U$10764 ( \11599 , \11593 , \11598 );
not \U$10765 ( \11600 , \11598 );
not \U$10766 ( \11601 , \11593 );
or \U$10767 ( \11602 , \11600 , \11601 );
or \U$10768 ( \11603 , \9545 , \11340 );
not \U$10769 ( \11604 , \9702 );
or \U$10770 ( \11605 , \11450 , \11604 );
or \U$10771 ( \11606 , \9543 , \11340 );
or \U$10772 ( \11607 , \9411 , \10860_nR251b );
nand \U$10773 ( \11608 , \11607 , \9699 );
nand \U$10774 ( \11609 , \11606 , \11608 );
nand \U$10775 ( \11610 , \11603 , \11605 , \11609 );
nand \U$10776 ( \11611 , \11602 , \11610 );
nand \U$10777 ( \11612 , \11599 , \11611 );
xor \U$10778 ( \11613 , \11586 , \11612 );
not \U$10779 ( \11614 , \11563 );
not \U$10780 ( \11615 , \11567 );
or \U$10781 ( \11616 , \11614 , \11615 );
or \U$10782 ( \11617 , \11567 , \11563 );
nand \U$10783 ( \11618 , \11616 , \11617 );
and \U$10784 ( \11619 , \11613 , \11618 );
and \U$10785 ( \11620 , \11586 , \11612 );
or \U$10786 ( \11621 , \11619 , \11620 );
xor \U$10787 ( \11622 , \11580 , \11621 );
not \U$10788 ( \11623 , \10686_nR2587 );
or \U$10789 ( \11624 , \10202 , \11623 );
or \U$10790 ( \11625 , \10686_nR2587 , \10013 );
or \U$10791 ( \11626 , \10860_nR251b , \10012 );
nand \U$10792 ( \11627 , \11624 , \11625 , \11626 );
xor \U$10793 ( \11628 , \11627 , \9718 );
or \U$10794 ( \11629 , \10202 , \11450 );
or \U$10795 ( \11630 , \10860_nR251b , \10013 );
or \U$10796 ( \11631 , \10926_nR23da , \10012 );
nand \U$10797 ( \11632 , \11629 , \11630 , \11631 );
nand \U$10798 ( \11633 , \10926_nR23da , \10010 );
and \U$10799 ( \11634 , \11632 , \9712 , \11633 );
xor \U$10800 ( \11635 , \11628 , \11634 );
not \U$10801 ( \11636 , \9949 );
or \U$10802 ( \11637 , \11636 , \11340 );
or \U$10803 ( \11638 , \10926_nR23da , \9717 );
nand \U$10804 ( \11639 , \11637 , \11638 , \9946 );
and \U$10805 ( \11640 , \11635 , \11639 );
and \U$10806 ( \11641 , \11628 , \11634 );
or \U$10807 ( \11642 , \11640 , \11641 );
and \U$10808 ( \11643 , \11627 , \9718 );
xor \U$10809 ( \11644 , \11642 , \11643 );
nand \U$10810 ( \11645 , \10926_nR23da , \9764 );
or \U$10811 ( \11646 , \9717 , \10860_nR251b );
nand \U$10812 ( \11647 , \11646 , \9946 );
and \U$10813 ( \11648 , \11645 , \11647 );
and \U$10814 ( \11649 , \9949 , \10860_nR251b );
and \U$10815 ( \11650 , \10926_nR23da , \9766 );
nor \U$10816 ( \11651 , \11648 , \11649 , \11650 );
not \U$10817 ( \11652 , \10568_nR260a );
and \U$10818 ( \11653 , \11652 , \10199 );
and \U$10819 ( \11654 , \10011 , \11623 );
and \U$10820 ( \11655 , \10568_nR260a , \10203 );
nor \U$10821 ( \11656 , \11653 , \11654 , \11655 );
and \U$10822 ( \11657 , \11651 , \11656 );
nor \U$10823 ( \11658 , \11651 , \11656 );
nor \U$10824 ( \11659 , \11657 , \11658 );
and \U$10825 ( \11660 , \11644 , \11659 );
and \U$10826 ( \11661 , \11642 , \11643 );
or \U$10827 ( \11662 , \11660 , \11661 );
xor \U$10828 ( \11663 , \11662 , \11658 );
and \U$10829 ( \11664 , \10926_nR23da , \9702 );
and \U$10830 ( \11665 , \11340 , \9412 );
not \U$10831 ( \11666 , \9699 );
nor \U$10832 ( \11667 , \11664 , \11665 , \11666 );
and \U$10833 ( \11668 , \11595 , \10199 );
and \U$10834 ( \11669 , \10011 , \11652 );
and \U$10835 ( \11670 , \10314_nR2685 , \10203 );
nor \U$10836 ( \11671 , \11668 , \11669 , \11670 );
xor \U$10837 ( \11672 , \9411 , \11671 );
nand \U$10838 ( \11673 , \10860_nR251b , \9764 );
or \U$10839 ( \11674 , \9717 , \10686_nR2587 );
nand \U$10840 ( \11675 , \11674 , \9946 );
and \U$10841 ( \11676 , \11673 , \11675 );
and \U$10842 ( \11677 , \9949 , \10686_nR2587 );
and \U$10843 ( \11678 , \10860_nR251b , \9766 );
nor \U$10844 ( \11679 , \11676 , \11677 , \11678 );
xor \U$10845 ( \11680 , \11672 , \11679 );
and \U$10846 ( \11681 , \11667 , \11680 );
nor \U$10847 ( \11682 , \11667 , \11680 );
nor \U$10848 ( \11683 , \11681 , \11682 );
and \U$10849 ( \11684 , \11663 , \11683 );
and \U$10850 ( \11685 , \11662 , \11658 );
or \U$10851 ( \11686 , \11684 , \11685 );
xor \U$10852 ( \11687 , \11686 , \11682 );
not \U$10853 ( \11688 , \11598 );
not \U$10854 ( \11689 , \11610 );
or \U$10855 ( \11690 , \11688 , \11689 );
or \U$10856 ( \11691 , \11610 , \11598 );
nand \U$10857 ( \11692 , \11690 , \11691 );
not \U$10858 ( \11693 , \11692 );
not \U$10859 ( \11694 , \11593 );
and \U$10860 ( \11695 , \11693 , \11694 );
and \U$10861 ( \11696 , \11692 , \11593 );
nor \U$10862 ( \11697 , \11695 , \11696 );
xor \U$10863 ( \11698 , \9411 , \11671 );
and \U$10864 ( \11699 , \11698 , \11679 );
and \U$10865 ( \11700 , \9411 , \11671 );
or \U$10866 ( \11701 , \11699 , \11700 );
and \U$10867 ( \11702 , \11697 , \11701 );
nor \U$10868 ( \11703 , \11697 , \11701 );
nor \U$10869 ( \11704 , \11702 , \11703 );
and \U$10870 ( \11705 , \11687 , \11704 );
and \U$10871 ( \11706 , \11686 , \11682 );
or \U$10872 ( \11707 , \11705 , \11706 );
xor \U$10873 ( \11708 , \11707 , \11703 );
xor \U$10874 ( \11709 , \11586 , \11612 );
xor \U$10875 ( \11710 , \11709 , \11618 );
and \U$10876 ( \11711 , \11708 , \11710 );
and \U$10877 ( \11712 , \11707 , \11703 );
or \U$10878 ( \11713 , \11711 , \11712 );
and \U$10879 ( \11714 , \11622 , \11713 );
and \U$10880 ( \11715 , \11580 , \11621 );
or \U$10881 ( \11716 , \11714 , \11715 );
xor \U$10882 ( \11717 , \11716 , \11579 );
and \U$10883 ( \11718 , \11530 , \11571 );
nor \U$10884 ( \11719 , \11718 , \11572 );
and \U$10885 ( \11720 , \11717 , \11719 );
and \U$10886 ( \11721 , \11716 , \11579 );
or \U$10887 ( \11722 , \11720 , \11721 );
and \U$10888 ( \11723 , \11573 , \11722 );
and \U$10889 ( \11724 , \11526 , \11572 );
or \U$10890 ( \11725 , \11723 , \11724 );
and \U$10891 ( \11726 , \11519 , \11725 );
and \U$10892 ( \11727 , \11477 , \11518 );
or \U$10893 ( \11728 , \11726 , \11727 );
and \U$10894 ( \11729 , \11470 , \11476 );
xor \U$10895 ( \11730 , \11728 , \11729 );
and \U$10896 ( \11731 , \11391 , \11461 );
nor \U$10897 ( \11732 , \11731 , \11462 );
and \U$10898 ( \11733 , \11730 , \11732 );
and \U$10899 ( \11734 , \11728 , \11729 );
or \U$10900 ( \11735 , \11733 , \11734 );
and \U$10901 ( \11736 , \11463 , \11735 );
and \U$10902 ( \11737 , \11389 , \11462 );
or \U$10903 ( \11738 , \11736 , \11737 );
and \U$10904 ( \11739 , \11387 , \11738 );
and \U$10905 ( \11740 , \11335 , \11386 );
or \U$10906 ( \11741 , \11739 , \11740 );
xor \U$10907 ( \11742 , \11247 , \11249 );
xor \U$10908 ( \11743 , \11742 , \11262 );
and \U$10909 ( \11744 , \11331 , \11743 );
xor \U$10910 ( \11745 , \11247 , \11249 );
xor \U$10911 ( \11746 , \11745 , \11262 );
and \U$10912 ( \11747 , \11332 , \11746 );
and \U$10913 ( \11748 , \11331 , \11332 );
or \U$10914 ( \11749 , \11744 , \11747 , \11748 );
xor \U$10915 ( \11750 , \11189 , \11265 );
xor \U$10916 ( \11751 , \11750 , \11268 );
nand \U$10917 ( \11752 , \11749 , \11751 );
and \U$10918 ( \11753 , \11741 , \11752 );
nor \U$10919 ( \11754 , \11751 , \11749 );
nor \U$10920 ( \11755 , \11753 , \11754 );
and \U$10921 ( \11756 , \11272 , \11755 );
and \U$10922 ( \11757 , \11184 , \11271 );
or \U$10923 ( \11758 , \11756 , \11757 );
not \U$10924 ( \11759 , \11758 );
and \U$10925 ( \11760 , \11177 , \11759 );
and \U$10926 ( \11761 , \11171 , \11176 );
or \U$10927 ( \11762 , \11760 , \11761 );
and \U$10928 ( \11763 , \11091 , \11762 );
and \U$10929 ( \11764 , \11003 , \11090 );
or \U$10930 ( \11765 , \11763 , \11764 );
and \U$10931 ( \11766 , \11001 , \11765 );
and \U$10932 ( \11767 , \10991 , \11000 );
or \U$10933 ( \11768 , \11766 , \11767 );
and \U$10934 ( \11769 , \10989 , \11768 );
and \U$10935 ( \11770 , \10812 , \10988 );
or \U$10936 ( \11771 , \11769 , \11770 );
and \U$10937 ( \11772 , \10810 , \11771 );
and \U$10938 ( \11773 , \10713 , \10809 );
or \U$10939 ( \11774 , \11772 , \11773 );
not \U$10940 ( \11775 , \10705 );
and \U$10941 ( \11776 , \11775 , \10533 );
not \U$10942 ( \11777 , \10533 );
nand \U$10943 ( \11778 , \11777 , \10705 );
and \U$10944 ( \11779 , \11778 , \10519 );
nor \U$10945 ( \11780 , \11776 , \11779 );
not \U$10946 ( \11781 , \10511 );
and \U$10947 ( \11782 , \10449 , \11781 );
not \U$10948 ( \11783 , \10449 );
nand \U$10949 ( \11784 , \11783 , \10511 );
and \U$10950 ( \11785 , \10457 , \11784 );
nor \U$10951 ( \11786 , \11782 , \11785 );
xor \U$10952 ( \11787 , \10191 , \10244 );
xor \U$10953 ( \11788 , \11787 , \10259 );
xor \U$10954 ( \11789 , \11786 , \11788 );
xor \U$10955 ( \11790 , \10415 , \10426 );
xor \U$10956 ( \11791 , \11790 , \10429 );
xor \U$10957 ( \11792 , \11789 , \11791 );
nand \U$10958 ( \11793 , \11780 , \11792 );
and \U$10959 ( \11794 , \11774 , \11793 );
nor \U$10960 ( \11795 , \11792 , \11780 );
nor \U$10961 ( \11796 , \11794 , \11795 );
xor \U$10962 ( \11797 , \10432 , \10433 );
xor \U$10963 ( \11798 , \11797 , \10439 );
xor \U$10964 ( \11799 , \11786 , \11788 );
and \U$10965 ( \11800 , \11799 , \11791 );
and \U$10966 ( \11801 , \11786 , \11788 );
or \U$10967 ( \11802 , \11800 , \11801 );
and \U$10968 ( \11803 , \11798 , \11802 );
or \U$10969 ( \11804 , \11796 , \11803 );
or \U$10970 ( \11805 , \11802 , \11798 );
nand \U$10971 ( \11806 , \11804 , \11805 );
and \U$10972 ( \11807 , \10444 , \11806 );
and \U$10973 ( \11808 , \10272 , \10443 );
or \U$10974 ( \11809 , \11807 , \11808 );
and \U$10975 ( \11810 , \10270 , \11809 );
and \U$10976 ( \11811 , \10162 , \10269 );
or \U$10977 ( \11812 , \11810 , \11811 );
and \U$10978 ( \11813 , \10160 , \11812 );
and \U$10979 ( \11814 , \10002 , \10159 );
or \U$10980 ( \11815 , \11813 , \11814 );
and \U$10981 ( \11816 , \9998 , \11815 );
and \U$10982 ( \11817 , \9995 , \9997 );
or \U$10983 ( \11818 , \11816 , \11817 );
and \U$10984 ( \11819 , \9859 , \11818 );
and \U$10985 ( \11820 , \9749 , \9858 );
or \U$10986 ( \11821 , \11819 , \11820 );
and \U$10987 ( \11822 , \9745 , \11821 );
and \U$10988 ( \11823 , \9742 , \9744 );
or \U$10989 ( \11824 , \11822 , \11823 );
and \U$10990 ( \11825 , \9625 , \11824 );
and \U$10991 ( \11826 , \9518 , \9624 );
or \U$10992 ( \11827 , \11825 , \11826 );
and \U$10993 ( \11828 , \9516 , \11827 );
and \U$10994 ( \11829 , \9393 , \9515 );
or \U$10995 ( \11830 , \11828 , \11829 );
not \U$10996 ( \11831 , \9192 );
not \U$10997 ( \11832 , \9196 );
nand \U$10998 ( \11833 , \11832 , \9198 );
not \U$10999 ( \11834 , \11833 );
or \U$11000 ( \11835 , \11831 , \11834 );
or \U$11001 ( \11836 , \11833 , \9192 );
nand \U$11002 ( \11837 , \11835 , \11836 );
or \U$11003 ( \11838 , \9389 , \9212 );
nand \U$11004 ( \11839 , \11838 , \9209 );
nand \U$11005 ( \11840 , \11837 , \11839 );
and \U$11006 ( \11841 , \11830 , \11840 );
nor \U$11007 ( \11842 , \11839 , \11837 );
nor \U$11008 ( \11843 , \11841 , \11842 );
nor \U$11009 ( \11844 , \9204 , \11843 );
nor \U$11010 ( \11845 , \9201 , \11844 );
not \U$11011 ( \11846 , \11845 );
or \U$11012 ( \11847 , \9089 , \11846 );
or \U$11013 ( \11848 , \11845 , \9088 );
nand \U$11014 ( \11849 , \11847 , \11848 );
not \U$11015 ( \11850 , \8783 );
and \U$11016 ( \11851 , \11850 , RIb55bd90_601);
nor \U$11017 ( \11852 , \11851 , \8791 , \8794 );
and \U$11018 ( \11853 , \11850 , RIb55bd18_600);
and \U$11019 ( \11854 , \8241 , \8772 );
nor \U$11020 ( \11855 , \11853 , \11854 );
nor \U$11021 ( \11856 , \11852 , \11855 );
nand \U$11022 ( \11857 , \8251 , \8784 );
or \U$11023 ( \11858 , \8783 , \8246 );
nand \U$11024 ( \11859 , \11858 , \8776 );
and \U$11025 ( \11860 , \11856 , \11857 , \11859 , \8237 );
and \U$11026 ( \11861 , RIb551890_249, \11860 );
and \U$11027 ( \11862 , RIb551db8_260, \8835 );
and \U$11028 ( \11863 , \8844 , RIb551ea8_262);
and \U$11029 ( \11864 , RIb551e30_261, \8839 );
nor \U$11030 ( \11865 , \11863 , \11864 );
and \U$11031 ( \11866 , \8829 , RIb551980_251);
and \U$11032 ( \11867 , RIb551908_250, \8831 );
nor \U$11033 ( \11868 , \11866 , \11867 );
and \U$11034 ( \11869 , \8806 , RIb5519f8_252);
and \U$11035 ( \11870 , RIb551a70_253, \8812 );
nor \U$11036 ( \11871 , \11869 , \11870 );
and \U$11037 ( \11872 , \8856 , RIb551f98_264);
and \U$11038 ( \11873 , RIb551f20_263, \8859 );
nor \U$11039 ( \11874 , \11872 , \11873 );
nand \U$11040 ( \11875 , \11865 , \11868 , \11871 , \11874 );
nor \U$11041 ( \11876 , \11861 , \11862 , \11875 );
and \U$11042 ( \11877 , \8800 , RIb551d40_259);
and \U$11043 ( \11878 , RIb551cc8_258, \8823 );
nor \U$11044 ( \11879 , \11877 , \11878 );
and \U$11045 ( \11880 , RIb551bd8_256, \8818 );
and \U$11046 ( \11881 , RIb551c50_257, \8825 );
and \U$11047 ( \11882 , \8850 , RIb551b60_255);
and \U$11048 ( \11883 , RIb551ae8_254, \8847 );
nor \U$11049 ( \11884 , \11882 , \11883 );
not \U$11050 ( \11885 , \11884 );
nor \U$11051 ( \11886 , \11880 , \11881 , \11885 );
nand \U$11052 ( \11887 , \11876 , \11879 , \8283 , \11886 );
buf \U$11053 ( \11888 , \11887 );
buf \U$11054 ( \11889 , \8307 );
_DC r2d01 ( \11890_nR2d01 , \11888 , \11889 );
xor \U$11055 ( \11891 , \8236 , \11890_nR2d01 );
and \U$11056 ( \11892 , RIb54acc0_19, \8831 );
and \U$11057 ( \11893 , RIb54b350_33, \8856 );
and \U$11058 ( \11894 , \8850 , RIb54af18_24);
and \U$11059 ( \11895 , RIb54aea0_23, \8847 );
nor \U$11060 ( \11896 , \11894 , \11895 );
and \U$11061 ( \11897 , \8823 , RIb54b080_27);
and \U$11062 ( \11898 , RIb54b008_26, \8825 );
nor \U$11063 ( \11899 , \11897 , \11898 );
and \U$11064 ( \11900 , \8835 , RIb54b170_29);
and \U$11065 ( \11901 , RIb54b0f8_28, \8800 );
nor \U$11066 ( \11902 , \11900 , \11901 );
and \U$11067 ( \11903 , \8818 , RIb54af90_25);
and \U$11068 ( \11904 , RIb54ac48_18, \11860 );
nor \U$11069 ( \11905 , \11903 , \11904 );
nand \U$11070 ( \11906 , \11896 , \11899 , \11902 , \11905 );
nor \U$11071 ( \11907 , \11892 , \11893 , \11906 );
and \U$11072 ( \11908 , \8859 , RIb54b2d8_32);
and \U$11073 ( \11909 , RIb54b260_31, \8844 );
nor \U$11074 ( \11910 , \11908 , \11909 );
and \U$11075 ( \11911 , RIb54b1e8_30, \8839 );
and \U$11076 ( \11912 , RIb54ae28_22, \8812 );
and \U$11077 ( \11913 , \8806 , RIb54adb0_21);
and \U$11078 ( \11914 , RIb54ad38_20, \8829 );
nor \U$11079 ( \11915 , \11913 , \11914 );
not \U$11080 ( \11916 , \11915 );
nor \U$11081 ( \11917 , \11911 , \11912 , \11916 );
nand \U$11082 ( \11918 , \11907 , \11910 , \8331 , \11917 );
buf \U$11083 ( \11919 , \11918 );
_DC r2b18 ( \11920_nR2b18 , \11919 , \11889 );
xor \U$11084 ( \11921 , \8315 , \11920_nR2b18 );
and \U$11085 ( \11922 , RIb54b4b8_36, \8831 );
and \U$11086 ( \11923 , RIb54bb48_50, \8856 );
and \U$11087 ( \11924 , \8850 , RIb54b710_41);
and \U$11088 ( \11925 , RIb54b698_40, \8847 );
nor \U$11089 ( \11926 , \11924 , \11925 );
and \U$11090 ( \11927 , \8823 , RIb54b878_44);
and \U$11091 ( \11928 , RIb54b800_43, \8825 );
nor \U$11092 ( \11929 , \11927 , \11928 );
and \U$11093 ( \11930 , \8835 , RIb54b968_46);
and \U$11094 ( \11931 , RIb54b8f0_45, \8800 );
nor \U$11095 ( \11932 , \11930 , \11931 );
and \U$11096 ( \11933 , \8818 , RIb54b788_42);
and \U$11097 ( \11934 , RIb54b440_35, \11860 );
nor \U$11098 ( \11935 , \11933 , \11934 );
nand \U$11099 ( \11936 , \11926 , \11929 , \11932 , \11935 );
nor \U$11100 ( \11937 , \11922 , \11923 , \11936 );
and \U$11101 ( \11938 , \8859 , RIb54bad0_49);
and \U$11102 ( \11939 , RIb54ba58_48, \8844 );
nor \U$11103 ( \11940 , \11938 , \11939 );
and \U$11104 ( \11941 , RIb54b9e0_47, \8839 );
and \U$11105 ( \11942 , RIb54b620_39, \8812 );
and \U$11106 ( \11943 , \8806 , RIb54b5a8_38);
and \U$11107 ( \11944 , RIb54b530_37, \8829 );
nor \U$11108 ( \11945 , \11943 , \11944 );
not \U$11109 ( \11946 , \11945 );
nor \U$11110 ( \11947 , \11941 , \11942 , \11946 );
nand \U$11111 ( \11948 , \11937 , \11940 , \8361 , \11947 );
buf \U$11112 ( \11949 , \11948 );
_DC r2b16 ( \11950_nR2b16 , \11949 , \11889 );
xor \U$11113 ( \11951 , \8351 , \11950_nR2b16 );
and \U$11114 ( \11952 , RIb54bcb0_53, \8831 );
and \U$11115 ( \11953 , RIb54c340_67, \8856 );
and \U$11116 ( \11954 , \8850 , RIb54bf08_58);
and \U$11117 ( \11955 , RIb54be90_57, \8847 );
nor \U$11118 ( \11956 , \11954 , \11955 );
and \U$11119 ( \11957 , \8823 , RIb54c070_61);
and \U$11120 ( \11958 , RIb54bff8_60, \8825 );
nor \U$11121 ( \11959 , \11957 , \11958 );
and \U$11122 ( \11960 , \8835 , RIb54c160_63);
and \U$11123 ( \11961 , RIb54c0e8_62, \8800 );
nor \U$11124 ( \11962 , \11960 , \11961 );
and \U$11125 ( \11963 , \8818 , RIb54bf80_59);
and \U$11126 ( \11964 , RIb54bc38_52, \11860 );
nor \U$11127 ( \11965 , \11963 , \11964 );
nand \U$11128 ( \11966 , \11956 , \11959 , \11962 , \11965 );
nor \U$11129 ( \11967 , \11952 , \11953 , \11966 );
and \U$11130 ( \11968 , \8859 , RIb54c2c8_66);
and \U$11131 ( \11969 , RIb54c250_65, \8844 );
nor \U$11132 ( \11970 , \11968 , \11969 );
and \U$11133 ( \11971 , RIb54c1d8_64, \8839 );
and \U$11134 ( \11972 , RIb54be18_56, \8812 );
and \U$11135 ( \11973 , \8806 , RIb54bda0_55);
and \U$11136 ( \11974 , RIb54bd28_54, \8829 );
nor \U$11137 ( \11975 , \11973 , \11974 );
not \U$11138 ( \11976 , \11975 );
nor \U$11139 ( \11977 , \11971 , \11972 , \11976 );
nand \U$11140 ( \11978 , \11967 , \11970 , \8397 , \11977 );
buf \U$11141 ( \11979 , \11978 );
_DC r295d ( \11980_nR295d , \11979 , \11889 );
xor \U$11142 ( \11981 , \8387 , \11980_nR295d );
and \U$11143 ( \11982 , RIb54c4a8_70, \8831 );
and \U$11144 ( \11983 , RIb54cb38_84, \8856 );
and \U$11145 ( \11984 , \8850 , RIb54c700_75);
and \U$11146 ( \11985 , RIb54c688_74, \8847 );
nor \U$11147 ( \11986 , \11984 , \11985 );
and \U$11148 ( \11987 , \8823 , RIb54c868_78);
and \U$11149 ( \11988 , RIb54c7f0_77, \8825 );
nor \U$11150 ( \11989 , \11987 , \11988 );
and \U$11151 ( \11990 , \8835 , RIb54c958_80);
and \U$11152 ( \11991 , RIb54c8e0_79, \8800 );
nor \U$11153 ( \11992 , \11990 , \11991 );
and \U$11154 ( \11993 , \8818 , RIb54c778_76);
and \U$11155 ( \11994 , RIb54c430_69, \11860 );
nor \U$11156 ( \11995 , \11993 , \11994 );
nand \U$11157 ( \11996 , \11986 , \11989 , \11992 , \11995 );
nor \U$11158 ( \11997 , \11982 , \11983 , \11996 );
and \U$11159 ( \11998 , \8859 , RIb54cac0_83);
and \U$11160 ( \11999 , RIb54ca48_82, \8844 );
nor \U$11161 ( \12000 , \11998 , \11999 );
and \U$11162 ( \12001 , RIb54c9d0_81, \8839 );
and \U$11163 ( \12002 , RIb54c610_73, \8812 );
and \U$11164 ( \12003 , \8806 , RIb54c598_72);
and \U$11165 ( \12004 , RIb54c520_71, \8829 );
nor \U$11166 ( \12005 , \12003 , \12004 );
not \U$11167 ( \12006 , \12005 );
nor \U$11168 ( \12007 , \12001 , \12002 , \12006 );
nand \U$11169 ( \12008 , \11997 , \12000 , \8436 , \12007 );
buf \U$11170 ( \12009 , \12008 );
_DC r295b ( \12010_nR295b , \12009 , \11889 );
xor \U$11171 ( \12011 , \8423 , \12010_nR295b );
and \U$11172 ( \12012 , RIb54cca0_87, \8831 );
and \U$11173 ( \12013 , RIb54d330_101, \8856 );
and \U$11174 ( \12014 , \8850 , RIb54cef8_92);
and \U$11175 ( \12015 , RIb54ce80_91, \8847 );
nor \U$11176 ( \12016 , \12014 , \12015 );
and \U$11177 ( \12017 , \8823 , RIb54d060_95);
and \U$11178 ( \12018 , RIb54cfe8_94, \8825 );
nor \U$11179 ( \12019 , \12017 , \12018 );
and \U$11180 ( \12020 , \8835 , RIb54d150_97);
and \U$11181 ( \12021 , RIb54d0d8_96, \8800 );
nor \U$11182 ( \12022 , \12020 , \12021 );
and \U$11183 ( \12023 , \8818 , RIb54cf70_93);
and \U$11184 ( \12024 , RIb54cc28_86, \11860 );
nor \U$11185 ( \12025 , \12023 , \12024 );
nand \U$11186 ( \12026 , \12016 , \12019 , \12022 , \12025 );
nor \U$11187 ( \12027 , \12012 , \12013 , \12026 );
and \U$11188 ( \12028 , \8859 , RIb54d2b8_100);
and \U$11189 ( \12029 , RIb54d240_99, \8844 );
nor \U$11190 ( \12030 , \12028 , \12029 );
and \U$11191 ( \12031 , RIb54d1c8_98, \8839 );
and \U$11192 ( \12032 , RIb54ce08_90, \8812 );
and \U$11193 ( \12033 , \8806 , RIb54cd90_89);
and \U$11194 ( \12034 , RIb54cd18_88, \8829 );
nor \U$11195 ( \12035 , \12033 , \12034 );
not \U$11196 ( \12036 , \12035 );
nor \U$11197 ( \12037 , \12031 , \12032 , \12036 );
nand \U$11198 ( \12038 , \12027 , \12030 , \8469 , \12037 );
buf \U$11199 ( \12039 , \12038 );
_DC r27d1 ( \12040_nR27d1 , \12039 , \11889 );
xor \U$11200 ( \12041 , \8459 , \12040_nR27d1 );
and \U$11201 ( \12042 , RIb54d498_104, \8831 );
and \U$11202 ( \12043 , RIb54db28_118, \8856 );
and \U$11203 ( \12044 , \8850 , RIb54d6f0_109);
and \U$11204 ( \12045 , RIb54d678_108, \8847 );
nor \U$11205 ( \12046 , \12044 , \12045 );
and \U$11206 ( \12047 , \8823 , RIb54d858_112);
and \U$11207 ( \12048 , RIb54d7e0_111, \8825 );
nor \U$11208 ( \12049 , \12047 , \12048 );
and \U$11209 ( \12050 , \8835 , RIb54d948_114);
and \U$11210 ( \12051 , RIb54d8d0_113, \8800 );
nor \U$11211 ( \12052 , \12050 , \12051 );
and \U$11212 ( \12053 , \8818 , RIb54d768_110);
and \U$11213 ( \12054 , RIb54d420_103, \11860 );
nor \U$11214 ( \12055 , \12053 , \12054 );
nand \U$11215 ( \12056 , \12046 , \12049 , \12052 , \12055 );
nor \U$11216 ( \12057 , \12042 , \12043 , \12056 );
and \U$11217 ( \12058 , \8859 , RIb54dab0_117);
and \U$11218 ( \12059 , RIb54da38_116, \8844 );
nor \U$11219 ( \12060 , \12058 , \12059 );
and \U$11220 ( \12061 , RIb54d9c0_115, \8839 );
and \U$11221 ( \12062 , RIb54d600_107, \8812 );
and \U$11222 ( \12063 , \8806 , RIb54d588_106);
and \U$11223 ( \12064 , RIb54d510_105, \8829 );
nor \U$11224 ( \12065 , \12063 , \12064 );
not \U$11225 ( \12066 , \12065 );
nor \U$11226 ( \12067 , \12061 , \12062 , \12066 );
nand \U$11227 ( \12068 , \12057 , \12060 , \8508 , \12067 );
buf \U$11228 ( \12069 , \12068 );
_DC r27cf ( \12070_nR27cf , \12069 , \11889 );
xor \U$11229 ( \12071 , \8495 , \12070_nR27cf );
and \U$11230 ( \12072 , RIb54dc90_121, \8831 );
and \U$11231 ( \12073 , RIb54e320_135, \8856 );
and \U$11232 ( \12074 , \8850 , RIb54dee8_126);
and \U$11233 ( \12075 , RIb54de70_125, \8847 );
nor \U$11234 ( \12076 , \12074 , \12075 );
and \U$11235 ( \12077 , \8823 , RIb54e050_129);
and \U$11236 ( \12078 , RIb54dfd8_128, \8825 );
nor \U$11237 ( \12079 , \12077 , \12078 );
and \U$11238 ( \12080 , \8835 , RIb54e140_131);
and \U$11239 ( \12081 , RIb54e0c8_130, \8800 );
nor \U$11240 ( \12082 , \12080 , \12081 );
and \U$11241 ( \12083 , \8818 , RIb54df60_127);
and \U$11242 ( \12084 , RIb54dc18_120, \11860 );
nor \U$11243 ( \12085 , \12083 , \12084 );
nand \U$11244 ( \12086 , \12076 , \12079 , \12082 , \12085 );
nor \U$11245 ( \12087 , \12072 , \12073 , \12086 );
and \U$11246 ( \12088 , \8859 , RIb54e2a8_134);
and \U$11247 ( \12089 , RIb54e230_133, \8844 );
nor \U$11248 ( \12090 , \12088 , \12089 );
and \U$11249 ( \12091 , RIb54e1b8_132, \8839 );
and \U$11250 ( \12092 , RIb54ddf8_124, \8812 );
and \U$11251 ( \12093 , \8806 , RIb54dd80_123);
and \U$11252 ( \12094 , RIb54dd08_122, \8829 );
nor \U$11253 ( \12095 , \12093 , \12094 );
not \U$11254 ( \12096 , \12095 );
nor \U$11255 ( \12097 , \12091 , \12092 , \12096 );
nand \U$11256 ( \12098 , \12087 , \12090 , \8547 , \12097 );
buf \U$11257 ( \12099 , \12098 );
_DC r2689 ( \12100_nR2689 , \12099 , \11889 );
xor \U$11258 ( \12101 , \8531 , \12100_nR2689 );
and \U$11259 ( \12102 , RIb54e488_138, \8831 );
and \U$11260 ( \12103 , RIb54eb18_152, \8856 );
and \U$11261 ( \12104 , \8850 , RIb54e6e0_143);
and \U$11262 ( \12105 , RIb54e668_142, \8847 );
nor \U$11263 ( \12106 , \12104 , \12105 );
and \U$11264 ( \12107 , \8823 , RIb54e848_146);
and \U$11265 ( \12108 , RIb54e7d0_145, \8825 );
nor \U$11266 ( \12109 , \12107 , \12108 );
and \U$11267 ( \12110 , \8835 , RIb54e938_148);
and \U$11268 ( \12111 , RIb54e8c0_147, \8800 );
nor \U$11269 ( \12112 , \12110 , \12111 );
and \U$11270 ( \12113 , \8818 , RIb54e758_144);
and \U$11271 ( \12114 , RIb54e410_137, \11860 );
nor \U$11272 ( \12115 , \12113 , \12114 );
nand \U$11273 ( \12116 , \12106 , \12109 , \12112 , \12115 );
nor \U$11274 ( \12117 , \12102 , \12103 , \12116 );
and \U$11275 ( \12118 , \8859 , RIb54eaa0_151);
and \U$11276 ( \12119 , RIb54ea28_150, \8844 );
nor \U$11277 ( \12120 , \12118 , \12119 );
and \U$11278 ( \12121 , RIb54e9b0_149, \8839 );
and \U$11279 ( \12122 , RIb54e5f0_141, \8812 );
and \U$11280 ( \12123 , \8806 , RIb54e578_140);
and \U$11281 ( \12124 , RIb54e500_139, \8829 );
nor \U$11282 ( \12125 , \12123 , \12124 );
not \U$11283 ( \12126 , \12125 );
nor \U$11284 ( \12127 , \12121 , \12122 , \12126 );
nand \U$11285 ( \12128 , \12117 , \12120 , \8577 , \12127 );
buf \U$11286 ( \12129 , \12128 );
_DC r2687 ( \12130_nR2687 , \12129 , \11889 );
xor \U$11287 ( \12131 , \8567 , \12130_nR2687 );
and \U$11288 ( \12132 , RIb54ec08_154, \11860 );
and \U$11289 ( \12133 , RIb54f130_165, \8835 );
and \U$11290 ( \12134 , \8844 , RIb54f220_167);
and \U$11291 ( \12135 , RIb54f1a8_166, \8839 );
nor \U$11292 ( \12136 , \12134 , \12135 );
and \U$11293 ( \12137 , \8806 , RIb54ed70_157);
and \U$11294 ( \12138 , RIb54ede8_158, \8812 );
nor \U$11295 ( \12139 , \12137 , \12138 );
and \U$11296 ( \12140 , \8829 , RIb54ecf8_156);
and \U$11297 ( \12141 , RIb54ec80_155, \8831 );
nor \U$11298 ( \12142 , \12140 , \12141 );
and \U$11299 ( \12143 , \8856 , RIb54f310_169);
and \U$11300 ( \12144 , RIb54f298_168, \8859 );
nor \U$11301 ( \12145 , \12143 , \12144 );
nand \U$11302 ( \12146 , \12136 , \12139 , \12142 , \12145 );
nor \U$11303 ( \12147 , \12132 , \12133 , \12146 );
and \U$11304 ( \12148 , \8800 , RIb54f0b8_164);
and \U$11305 ( \12149 , RIb54f040_163, \8823 );
nor \U$11306 ( \12150 , \12148 , \12149 );
and \U$11307 ( \12151 , RIb54ef50_161, \8818 );
and \U$11308 ( \12152 , RIb54efc8_162, \8825 );
and \U$11309 ( \12153 , \8850 , RIb54eed8_160);
and \U$11310 ( \12154 , RIb54ee60_159, \8847 );
nor \U$11311 ( \12155 , \12153 , \12154 );
not \U$11312 ( \12156 , \12155 );
nor \U$11313 ( \12157 , \12151 , \12152 , \12156 );
nand \U$11314 ( \12158 , \12147 , \12150 , \8613 , \12157 );
buf \U$11315 ( \12159 , \12158 );
_DC r25a9 ( \12160_nR25a9 , \12159 , \11889 );
xor \U$11316 ( \12161 , \8603 , \12160_nR25a9 );
and \U$11317 ( \12162 , RIb54f478_172, \8831 );
and \U$11318 ( \12163 , RIb54fb08_186, \8856 );
and \U$11319 ( \12164 , \8818 , RIb54f748_178);
and \U$11320 ( \12165 , RIb54f6d0_177, \8850 );
nor \U$11321 ( \12166 , \12164 , \12165 );
and \U$11322 ( \12167 , \8823 , RIb54f838_180);
and \U$11323 ( \12168 , RIb54f7c0_179, \8825 );
nor \U$11324 ( \12169 , \12167 , \12168 );
and \U$11325 ( \12170 , \8835 , RIb54f928_182);
and \U$11326 ( \12171 , RIb54f8b0_181, \8800 );
nor \U$11327 ( \12172 , \12170 , \12171 );
and \U$11328 ( \12173 , \8847 , RIb54f658_176);
and \U$11329 ( \12174 , RIb54f400_171, \11860 );
nor \U$11330 ( \12175 , \12173 , \12174 );
nand \U$11331 ( \12176 , \12166 , \12169 , \12172 , \12175 );
nor \U$11332 ( \12177 , \12162 , \12163 , \12176 );
and \U$11333 ( \12178 , \8859 , RIb54fa90_185);
and \U$11334 ( \12179 , RIb54fa18_184, \8844 );
nor \U$11335 ( \12180 , \12178 , \12179 );
and \U$11336 ( \12181 , RIb54f9a0_183, \8839 );
and \U$11337 ( \12182 , RIb54f5e0_175, \8812 );
and \U$11338 ( \12183 , \8806 , RIb54f568_174);
and \U$11339 ( \12184 , RIb54f4f0_173, \8829 );
nor \U$11340 ( \12185 , \12183 , \12184 );
not \U$11341 ( \12186 , \12185 );
nor \U$11342 ( \12187 , \12181 , \12182 , \12186 );
nand \U$11343 ( \12188 , \12177 , \12180 , \8648 , \12187 );
buf \U$11344 ( \12189 , \12188 );
_DC r25ab ( \12190_nR25ab , \12189 , \11889 );
xor \U$11345 ( \12191 , \8635 , \12190_nR25ab );
and \U$11346 ( \12192 , RIb5504e0_207, \8831 );
and \U$11347 ( \12193 , RIb550b70_221, \8856 );
and \U$11348 ( \12194 , \8850 , RIb550738_212);
and \U$11349 ( \12195 , RIb5506c0_211, \8847 );
nor \U$11350 ( \12196 , \12194 , \12195 );
and \U$11351 ( \12197 , \8823 , RIb5508a0_215);
and \U$11352 ( \12198 , RIb550828_214, \8825 );
nor \U$11353 ( \12199 , \12197 , \12198 );
and \U$11354 ( \12200 , \8835 , RIb550990_217);
and \U$11355 ( \12201 , RIb550918_216, \8800 );
nor \U$11356 ( \12202 , \12200 , \12201 );
and \U$11357 ( \12203 , \8818 , RIb5507b0_213);
and \U$11358 ( \12204 , RIb550468_206, \11860 );
nor \U$11359 ( \12205 , \12203 , \12204 );
nand \U$11360 ( \12206 , \12196 , \12199 , \12202 , \12205 );
nor \U$11361 ( \12207 , \12192 , \12193 , \12206 );
and \U$11362 ( \12208 , \8859 , RIb550af8_220);
and \U$11363 ( \12209 , RIb550a80_219, \8844 );
nor \U$11364 ( \12210 , \12208 , \12209 );
and \U$11365 ( \12211 , RIb550a08_218, \8839 );
and \U$11366 ( \12212 , RIb550648_210, \8812 );
and \U$11367 ( \12213 , \8806 , RIb5505d0_209);
and \U$11368 ( \12214 , RIb550558_208, \8829 );
nor \U$11369 ( \12215 , \12213 , \12214 );
not \U$11370 ( \12216 , \12215 );
nor \U$11371 ( \12217 , \12211 , \12212 , \12216 );
nand \U$11372 ( \12218 , \12207 , \12210 , \8676 , \12217 );
buf \U$11373 ( \12219 , \12218 );
_DC r2433 ( \12220_nR2433 , \12219 , \11889 );
nand \U$11374 ( \12221 , \12220_nR2433 , \8697 );
and \U$11375 ( \12222 , RIb54fbf8_188, \11860 );
and \U$11376 ( \12223 , RIb550120_199, \8835 );
and \U$11377 ( \12224 , \8844 , RIb550210_201);
and \U$11378 ( \12225 , RIb550198_200, \8839 );
nor \U$11379 ( \12226 , \12224 , \12225 );
and \U$11380 ( \12227 , \8806 , RIb54fd60_191);
and \U$11381 ( \12228 , RIb54fdd8_192, \8812 );
nor \U$11382 ( \12229 , \12227 , \12228 );
and \U$11383 ( \12230 , \8829 , RIb54fce8_190);
and \U$11384 ( \12231 , RIb54fc70_189, \8831 );
nor \U$11385 ( \12232 , \12230 , \12231 );
and \U$11386 ( \12233 , \8856 , RIb550300_203);
and \U$11387 ( \12234 , RIb550288_202, \8859 );
nor \U$11388 ( \12235 , \12233 , \12234 );
nand \U$11389 ( \12236 , \12226 , \12229 , \12232 , \12235 );
nor \U$11390 ( \12237 , \12222 , \12223 , \12236 );
and \U$11391 ( \12238 , \8800 , RIb5500a8_198);
and \U$11392 ( \12239 , RIb550030_197, \8823 );
nor \U$11393 ( \12240 , \12238 , \12239 );
and \U$11394 ( \12241 , RIb54ff40_195, \8818 );
and \U$11395 ( \12242 , RIb54ffb8_196, \8825 );
and \U$11396 ( \12243 , \8850 , RIb54fec8_194);
and \U$11397 ( \12244 , RIb54fe50_193, \8847 );
nor \U$11398 ( \12245 , \12243 , \12244 );
not \U$11399 ( \12246 , \12245 );
nor \U$11400 ( \12247 , \12241 , \12242 , \12246 );
nand \U$11401 ( \12248 , \12237 , \12240 , \8714 , \12247 );
buf \U$11402 ( \12249 , \12248 );
_DC r2435 ( \12250_nR2435 , \12249 , \11889 );
nand \U$11403 ( \12251 , \12250_nR2435 , RIb55bca0_599);
and \U$11404 ( \12252 , \12221 , \12251 );
nor \U$11405 ( \12253 , RIb55bca0_599, \12250_nR2435 );
nor \U$11406 ( \12254 , \12252 , \12253 );
and \U$11407 ( \12255 , \12191 , \12254 );
and \U$11408 ( \12256 , \8635 , \12190_nR25ab );
or \U$11409 ( \12257 , \12255 , \12256 );
and \U$11410 ( \12258 , \12161 , \12257 );
and \U$11411 ( \12259 , \8603 , \12160_nR25a9 );
or \U$11412 ( \12260 , \12258 , \12259 );
and \U$11413 ( \12261 , \12131 , \12260 );
and \U$11414 ( \12262 , \8567 , \12130_nR2687 );
or \U$11415 ( \12263 , \12261 , \12262 );
and \U$11416 ( \12264 , \12101 , \12263 );
and \U$11417 ( \12265 , \8531 , \12100_nR2689 );
or \U$11418 ( \12266 , \12264 , \12265 );
and \U$11419 ( \12267 , \12071 , \12266 );
and \U$11420 ( \12268 , \8495 , \12070_nR27cf );
or \U$11421 ( \12269 , \12267 , \12268 );
and \U$11422 ( \12270 , \12041 , \12269 );
and \U$11423 ( \12271 , \8459 , \12040_nR27d1 );
or \U$11424 ( \12272 , \12270 , \12271 );
and \U$11425 ( \12273 , \12011 , \12272 );
and \U$11426 ( \12274 , \8423 , \12010_nR295b );
or \U$11427 ( \12275 , \12273 , \12274 );
and \U$11428 ( \12276 , \11981 , \12275 );
and \U$11429 ( \12277 , \8387 , \11980_nR295d );
or \U$11430 ( \12278 , \12276 , \12277 );
and \U$11431 ( \12279 , \11951 , \12278 );
and \U$11432 ( \12280 , \8351 , \11950_nR2b16 );
or \U$11433 ( \12281 , \12279 , \12280 );
and \U$11434 ( \12282 , \11921 , \12281 );
and \U$11435 ( \12283 , \8315 , \11920_nR2b18 );
or \U$11436 ( \12284 , \12282 , \12283 );
and \U$11437 ( \12285 , \11891 , \12284 );
and \U$11438 ( \12286 , \8236 , \11890_nR2d01 );
or \U$11439 ( \12287 , \12285 , \12286 );
nor \U$11440 ( \12288 , \12287 , \8767 );
not \U$11441 ( \12289 , \12288 );
and \U$11442 ( \12290 , \11856 , \8772 );
and \U$11443 ( \12291 , \11859 , \12290 );
xnor \U$11444 ( \12292 , \11857 , \12291 );
not \U$11445 ( \12293 , \12292 );
xor \U$11446 ( \12294 , \11859 , \12290 );
not \U$11447 ( \12295 , \12294 );
and \U$11448 ( \12296 , \12291 , \11857 );
nor \U$11449 ( \12297 , \12296 , RIb55bef8_604);
nand \U$11450 ( \12298 , \12295 , \12297 );
nor \U$11451 ( \12299 , \12293 , \12298 );
not \U$11452 ( \12300 , \12299 );
not \U$11453 ( \12301 , \11855 );
and \U$11454 ( \12302 , \11852 , \8772 , \12301 );
nor \U$11455 ( \12303 , \12302 , \8793 );
not \U$11456 ( \12304 , \12303 );
and \U$11457 ( \12305 , \11855 , \8772 );
and \U$11458 ( \12306 , RIb55bd18_600, \8782 );
nor \U$11459 ( \12307 , \12305 , \12306 );
nand \U$11460 ( \12308 , \12304 , \12307 );
nor \U$11461 ( \12309 , \12300 , \12308 );
and \U$11462 ( \12310 , RIb551638_244, \12309 );
nand \U$11463 ( \12311 , \12307 , \12303 );
nor \U$11464 ( \12312 , \12297 , \12311 , \12294 );
and \U$11465 ( \12313 , \12312 , \12292 );
and \U$11466 ( \12314 , RIb550be8_222, \12313 );
not \U$11467 ( \12315 , \12303 );
nor \U$11468 ( \12316 , \12315 , \12307 );
and \U$11469 ( \12317 , \12299 , \12316 );
and \U$11470 ( \12318 , \12317 , RIb5516b0_245);
nor \U$11471 ( \12319 , \12303 , \12307 );
and \U$11472 ( \12320 , \12299 , \12319 );
and \U$11473 ( \12321 , RIb5515c0_243, \12320 );
nor \U$11474 ( \12322 , \12318 , \12321 );
or \U$11475 ( \12323 , \12298 , \12292 );
nor \U$11476 ( \12324 , \12323 , \12311 );
and \U$11477 ( \12325 , \12324 , RIb551368_238);
not \U$11478 ( \12326 , \12316 );
nor \U$11479 ( \12327 , \12326 , \12323 );
and \U$11480 ( \12328 , RIb5512f0_237, \12327 );
nor \U$11481 ( \12329 , \12325 , \12328 );
nor \U$11482 ( \12330 , \12323 , \12308 );
and \U$11483 ( \12331 , \12330 , RIb551278_236);
not \U$11484 ( \12332 , \12319 );
nor \U$11485 ( \12333 , \12332 , \12323 );
and \U$11486 ( \12334 , RIb551200_235, \12333 );
nor \U$11487 ( \12335 , \12331 , \12334 );
nand \U$11488 ( \12336 , \12294 , \12297 );
or \U$11489 ( \12337 , \12336 , \12292 );
nor \U$11490 ( \12338 , \12337 , \12311 );
and \U$11491 ( \12339 , \12338 , RIb551188_234);
not \U$11492 ( \12340 , \12316 );
nor \U$11493 ( \12341 , \12340 , \12337 );
and \U$11494 ( \12342 , RIb551110_233, \12341 );
nor \U$11495 ( \12343 , \12339 , \12342 );
nand \U$11496 ( \12344 , \12322 , \12329 , \12335 , \12343 );
nor \U$11497 ( \12345 , \12310 , \12314 , \12344 );
not \U$11498 ( \12346 , \12292 );
nor \U$11499 ( \12347 , \12346 , \12336 );
not \U$11500 ( \12348 , \12347 );
nor \U$11501 ( \12349 , \12348 , \12311 );
and \U$11502 ( \12350 , \12349 , RIb551548_242);
and \U$11503 ( \12351 , \12347 , \12316 );
and \U$11504 ( \12352 , RIb5514d0_241, \12351 );
nor \U$11505 ( \12353 , \12350 , \12352 );
nand \U$11506 ( \12354 , RIb551728_246, \8856 );
not \U$11507 ( \12355 , \12347 );
nor \U$11508 ( \12356 , \12355 , \12308 );
and \U$11509 ( \12357 , RIb551458_240, \12356 );
and \U$11510 ( \12358 , \12347 , \12319 );
and \U$11511 ( \12359 , RIb5513e0_239, \12358 );
nor \U$11512 ( \12360 , \12337 , \12308 );
and \U$11513 ( \12361 , \12360 , RIb551098_232);
not \U$11514 ( \12362 , \12319 );
nor \U$11515 ( \12363 , \12362 , \12337 );
and \U$11516 ( \12364 , RIb551020_231, \12363 );
nor \U$11517 ( \12365 , \12361 , \12364 );
not \U$11518 ( \12366 , \12365 );
nor \U$11519 ( \12367 , \12357 , \12359 , \12366 );
nand \U$11520 ( \12368 , \12345 , \12353 , \12354 , \12367 );
buf \U$11521 ( \12369 , \8307 );
_DC r3379 ( \12370_nR3379 , \12368 , \12369 );
not \U$11522 ( \12371 , \12370_nR3379 );
nor \U$11523 ( \12372 , \12289 , \12371 );
and \U$11524 ( \12373 , \12287 , \8767 );
nor \U$11525 ( \12374 , \12373 , \12288 );
xor \U$11526 ( \12375 , \8236 , \11890_nR2d01 );
xor \U$11527 ( \12376 , \12375 , \12284 );
and \U$11528 ( \12377 , \12374 , \12376 );
nor \U$11529 ( \12378 , \12374 , \12376 );
xor \U$11530 ( \12379 , \8315 , \11920_nR2b18 );
xor \U$11531 ( \12380 , \12379 , \12281 );
xor \U$11532 ( \12381 , \12376 , \12380 );
nor \U$11533 ( \12382 , \12377 , \12378 , \12381 );
not \U$11534 ( \12383 , \12376 );
not \U$11535 ( \12384 , \12380 );
and \U$11536 ( \12385 , \12383 , \12384 );
nor \U$11537 ( \12386 , \12385 , \12374 );
not \U$11538 ( \12387 , \12386 );
and \U$11539 ( \12388 , \12382 , \12387 );
not \U$11540 ( \12389 , \12388 );
and \U$11541 ( \12390 , RIb552628_278, \12320 );
and \U$11542 ( \12391 , RIb552010_265, \12313 );
and \U$11543 ( \12392 , \12317 , RIb552718_280);
and \U$11544 ( \12393 , RIb5526a0_279, \12309 );
nor \U$11545 ( \12394 , \12392 , \12393 );
and \U$11546 ( \12395 , \12324 , RIb5523d0_273);
and \U$11547 ( \12396 , RIb552358_272, \12327 );
nor \U$11548 ( \12397 , \12395 , \12396 );
and \U$11549 ( \12398 , \12330 , RIb5522e0_271);
and \U$11550 ( \12399 , RIb552268_270, \12333 );
nor \U$11551 ( \12400 , \12398 , \12399 );
and \U$11552 ( \12401 , \12338 , RIb5521f0_269);
and \U$11553 ( \12402 , RIb552178_268, \12341 );
nor \U$11554 ( \12403 , \12401 , \12402 );
nand \U$11555 ( \12404 , \12394 , \12397 , \12400 , \12403 );
nor \U$11556 ( \12405 , \12390 , \12391 , \12404 );
and \U$11557 ( \12406 , \12349 , RIb5525b0_277);
and \U$11558 ( \12407 , RIb552538_276, \12351 );
nor \U$11559 ( \12408 , \12406 , \12407 );
nand \U$11560 ( \12409 , RIb552790_281, \8856 );
and \U$11561 ( \12410 , RIb5524c0_275, \12356 );
and \U$11562 ( \12411 , RIb552448_274, \12358 );
and \U$11563 ( \12412 , \12360 , RIb552100_267);
and \U$11564 ( \12413 , RIb552088_266, \12363 );
nor \U$11565 ( \12414 , \12412 , \12413 );
not \U$11566 ( \12415 , \12414 );
nor \U$11567 ( \12416 , \12410 , \12411 , \12415 );
nand \U$11568 ( \12417 , \12405 , \12408 , \12409 , \12416 );
_DC r349f ( \12418_nR349f , \12417 , \12369 );
not \U$11569 ( \12419 , \12418_nR349f );
or \U$11570 ( \12420 , \12389 , \12419 );
or \U$11571 ( \12421 , \12418_nR349f , \12387 );
or \U$11572 ( \12422 , \12382 , \12387 );
nand \U$11573 ( \12423 , \12420 , \12421 , \12422 );
xnor \U$11574 ( \12424 , \12372 , \12423 );
not \U$11575 ( \12425 , \12381 );
nor \U$11576 ( \12426 , \12386 , \12425 );
not \U$11577 ( \12427 , \12426 );
or \U$11578 ( \12428 , \12427 , \12419 );
or \U$11579 ( \12429 , \12371 , \12389 );
or \U$11580 ( \12430 , \12425 , \12419 );
or \U$11581 ( \12431 , \12387 , \12370_nR3379 );
nand \U$11582 ( \12432 , \12431 , \12422 );
nand \U$11583 ( \12433 , \12430 , \12432 );
nand \U$11584 ( \12434 , \12428 , \12429 , \12433 );
xor \U$11585 ( \12435 , \8351 , \11950_nR2b16 );
xor \U$11586 ( \12436 , \12435 , \12278 );
xor \U$11587 ( \12437 , \8387 , \11980_nR295d );
xor \U$11588 ( \12438 , \12437 , \12275 );
nor \U$11589 ( \12439 , \12436 , \12438 );
or \U$11590 ( \12440 , \12380 , \12439 );
and \U$11591 ( \12441 , \12434 , \12440 );
and \U$11592 ( \12442 , RIb552f10_297, \12317 );
and \U$11593 ( \12443 , RIb552808_282, \12313 );
and \U$11594 ( \12444 , \12330 , RIb552ad8_288);
and \U$11595 ( \12445 , RIb552a60_287, \12333 );
nor \U$11596 ( \12446 , \12444 , \12445 );
and \U$11597 ( \12447 , \12324 , RIb552bc8_290);
and \U$11598 ( \12448 , RIb552b50_289, \12327 );
nor \U$11599 ( \12449 , \12447 , \12448 );
and \U$11600 ( \12450 , \12338 , RIb5529e8_286);
and \U$11601 ( \12451 , RIb552970_285, \12341 );
nor \U$11602 ( \12452 , \12450 , \12451 );
and \U$11603 ( \12453 , \12356 , RIb552cb8_292);
and \U$11604 ( \12454 , RIb552c40_291, \12358 );
nor \U$11605 ( \12455 , \12453 , \12454 );
nand \U$11606 ( \12456 , \12446 , \12449 , \12452 , \12455 );
nor \U$11607 ( \12457 , \12442 , \12443 , \12456 );
and \U$11608 ( \12458 , \12309 , RIb552e98_296);
and \U$11609 ( \12459 , RIb552e20_295, \12320 );
nor \U$11610 ( \12460 , \12458 , \12459 );
nand \U$11611 ( \12461 , RIb552f88_298, \8856 );
and \U$11612 ( \12462 , RIb552da8_294, \12349 );
and \U$11613 ( \12463 , RIb552d30_293, \12351 );
and \U$11614 ( \12464 , \12360 , RIb5528f8_284);
and \U$11615 ( \12465 , RIb552880_283, \12363 );
nor \U$11616 ( \12466 , \12464 , \12465 );
not \U$11617 ( \12467 , \12466 );
nor \U$11618 ( \12468 , \12462 , \12463 , \12467 );
nand \U$11619 ( \12469 , \12457 , \12460 , \12461 , \12468 );
_DC r3271 ( \12470_nR3271 , \12469 , \12369 );
nand \U$11620 ( \12471 , \12470_nR3271 , \12288 );
not \U$11621 ( \12472 , \12471 );
nor \U$11622 ( \12473 , \12441 , \12472 );
xor \U$11623 ( \12474 , \12424 , \12473 );
not \U$11624 ( \12475 , \12474 );
not \U$11625 ( \12476 , \12436 );
not \U$11626 ( \12477 , \12380 );
or \U$11627 ( \12478 , \12476 , \12477 );
or \U$11628 ( \12479 , \12380 , \12436 );
nand \U$11629 ( \12480 , \12478 , \12479 );
xor \U$11630 ( \12481 , \12438 , \12436 );
nor \U$11631 ( \12482 , \12480 , \12481 );
not \U$11632 ( \12483 , \12482 );
not \U$11633 ( \12484 , \12440 );
nor \U$11634 ( \12485 , \12483 , \12484 );
not \U$11635 ( \12486 , \12485 );
or \U$11636 ( \12487 , \12486 , \12419 );
or \U$11637 ( \12488 , \12483 , \12419 );
nand \U$11638 ( \12489 , \12488 , \12484 );
nand \U$11639 ( \12490 , \12487 , \12489 );
or \U$11640 ( \12491 , \12427 , \12371 );
not \U$11641 ( \12492 , \12470_nR3271 );
or \U$11642 ( \12493 , \12492 , \12389 );
or \U$11643 ( \12494 , \12425 , \12371 );
or \U$11644 ( \12495 , \12387 , \12470_nR3271 );
nand \U$11645 ( \12496 , \12495 , \12422 );
nand \U$11646 ( \12497 , \12494 , \12496 );
nand \U$11647 ( \12498 , \12491 , \12493 , \12497 );
and \U$11648 ( \12499 , \12490 , \12498 );
not \U$11649 ( \12500 , \12471 );
and \U$11650 ( \12501 , \12434 , \12440 );
not \U$11651 ( \12502 , \12434 );
and \U$11652 ( \12503 , \12502 , \12484 );
nor \U$11653 ( \12504 , \12501 , \12503 );
not \U$11654 ( \12505 , \12504 );
or \U$11655 ( \12506 , \12500 , \12505 );
or \U$11656 ( \12507 , \12504 , \12471 );
nand \U$11657 ( \12508 , \12506 , \12507 );
and \U$11658 ( \12509 , \12499 , \12508 );
xor \U$11659 ( \12510 , \12475 , \12509 );
and \U$11660 ( \12511 , \12370_nR3379 , \12485 );
and \U$11661 ( \12512 , \12440 , \12481 );
and \U$11662 ( \12513 , \12512 , \12418_nR349f );
nand \U$11663 ( \12514 , \12370_nR3379 , \12482 );
or \U$11664 ( \12515 , \12440 , \12418_nR349f );
or \U$11665 ( \12516 , \12440 , \12481 );
nand \U$11666 ( \12517 , \12515 , \12516 );
and \U$11667 ( \12518 , \12514 , \12517 );
nor \U$11668 ( \12519 , \12511 , \12513 , \12518 );
and \U$11669 ( \12520 , \12470_nR3271 , \12426 );
and \U$11670 ( \12521 , RIb553f00_331, \12317 );
and \U$11671 ( \12522 , RIb5537f8_316, \12313 );
and \U$11672 ( \12523 , \12309 , RIb553e88_330);
and \U$11673 ( \12524 , RIb553e10_329, \12320 );
nor \U$11674 ( \12525 , \12523 , \12524 );
and \U$11675 ( \12526 , \12324 , RIb553bb8_324);
and \U$11676 ( \12527 , RIb553b40_323, \12327 );
nor \U$11677 ( \12528 , \12526 , \12527 );
and \U$11678 ( \12529 , \12330 , RIb553ac8_322);
and \U$11679 ( \12530 , RIb553a50_321, \12333 );
nor \U$11680 ( \12531 , \12529 , \12530 );
and \U$11681 ( \12532 , \12338 , RIb5539d8_320);
and \U$11682 ( \12533 , RIb553960_319, \12341 );
nor \U$11683 ( \12534 , \12532 , \12533 );
nand \U$11684 ( \12535 , \12525 , \12528 , \12531 , \12534 );
nor \U$11685 ( \12536 , \12521 , \12522 , \12535 );
and \U$11686 ( \12537 , \12349 , RIb553d98_328);
and \U$11687 ( \12538 , RIb553d20_327, \12351 );
nor \U$11688 ( \12539 , \12537 , \12538 );
nand \U$11689 ( \12540 , RIb553f78_332, \8856 );
and \U$11690 ( \12541 , RIb553ca8_326, \12356 );
and \U$11691 ( \12542 , RIb553c30_325, \12358 );
and \U$11692 ( \12543 , \12360 , RIb5538e8_318);
and \U$11693 ( \12544 , RIb553870_317, \12363 );
nor \U$11694 ( \12545 , \12543 , \12544 );
not \U$11695 ( \12546 , \12545 );
nor \U$11696 ( \12547 , \12541 , \12542 , \12546 );
nand \U$11697 ( \12548 , \12536 , \12539 , \12540 , \12547 );
_DC r3150 ( \12549_nR3150 , \12548 , \12369 );
and \U$11698 ( \12550 , \12388 , \12549_nR3150 );
nand \U$11699 ( \12551 , \12470_nR3271 , \12381 );
or \U$11700 ( \12552 , \12387 , \12549_nR3150 );
nand \U$11701 ( \12553 , \12552 , \12422 );
and \U$11702 ( \12554 , \12551 , \12553 );
nor \U$11703 ( \12555 , \12520 , \12550 , \12554 );
nand \U$11704 ( \12556 , \12519 , \12555 );
xor \U$11705 ( \12557 , \8423 , \12010_nR295b );
xor \U$11706 ( \12558 , \12557 , \12272 );
xor \U$11707 ( \12559 , \8459 , \12040_nR27d1 );
xor \U$11708 ( \12560 , \12559 , \12269 );
nor \U$11709 ( \12561 , \12558 , \12560 );
or \U$11710 ( \12562 , \12438 , \12561 );
and \U$11711 ( \12563 , \12556 , \12562 );
nor \U$11712 ( \12564 , \12555 , \12519 );
nor \U$11713 ( \12565 , \12563 , \12564 );
xor \U$11714 ( \12566 , \12490 , \12498 );
not \U$11715 ( \12567 , \12566 );
nand \U$11716 ( \12568 , \12549_nR3150 , \12288 );
not \U$11717 ( \12569 , \12568 );
and \U$11718 ( \12570 , \12567 , \12569 );
and \U$11719 ( \12571 , \12566 , \12568 );
nor \U$11720 ( \12572 , \12570 , \12571 );
nand \U$11721 ( \12573 , \12565 , \12572 );
xor \U$11722 ( \12574 , \12499 , \12508 );
and \U$11723 ( \12575 , \12573 , \12574 );
and \U$11724 ( \12576 , \12510 , \12575 );
not \U$11725 ( \12577 , \12576 );
and \U$11726 ( \12578 , \12475 , \12509 );
or \U$11727 ( \12579 , \12578 , \12386 );
and \U$11728 ( \12580 , \12578 , \12386 );
and \U$11729 ( \12581 , \12372 , \12423 );
nor \U$11730 ( \12582 , \12580 , \12581 );
nand \U$11731 ( \12583 , \12579 , \12582 );
not \U$11732 ( \12584 , \12583 );
and \U$11733 ( \12585 , \12288 , \12418_nR349f );
and \U$11734 ( \12586 , \12424 , \12473 );
nor \U$11735 ( \12587 , \12585 , \12586 );
not \U$11736 ( \12588 , \12587 );
and \U$11737 ( \12589 , \12584 , \12588 );
and \U$11738 ( \12590 , \12583 , \12587 );
nor \U$11739 ( \12591 , \12589 , \12590 );
not \U$11740 ( \12592 , \12591 );
or \U$11741 ( \12593 , \12577 , \12592 );
or \U$11742 ( \12594 , \12591 , \12576 );
nand \U$11743 ( \12595 , \12593 , \12594 );
not \U$11744 ( \12596 , \12595 );
xor \U$11745 ( \12597 , \12573 , \12574 );
not \U$11746 ( \12598 , \12566 );
nor \U$11747 ( \12599 , \12598 , \12568 );
xor \U$11748 ( \12600 , \12597 , \12599 );
or \U$11749 ( \12601 , \12572 , \12565 );
nand \U$11750 ( \12602 , \12601 , \12573 );
not \U$11751 ( \12603 , \12602 );
and \U$11752 ( \12604 , RIb553168_302, \12341 );
and \U$11753 ( \12605 , RIb5534b0_309, \12356 );
and \U$11754 ( \12606 , \12309 , RIb553690_313);
and \U$11755 ( \12607 , RIb553618_312, \12320 );
nor \U$11756 ( \12608 , \12606 , \12607 );
and \U$11757 ( \12609 , \12360 , RIb5530f0_301);
and \U$11758 ( \12610 , RIb553078_300, \12363 );
nor \U$11759 ( \12611 , \12609 , \12610 );
and \U$11760 ( \12612 , \12317 , RIb553708_314);
and \U$11761 ( \12613 , RIb553000_299, \12313 );
nor \U$11762 ( \12614 , \12612 , \12613 );
and \U$11763 ( \12615 , \12349 , RIb5535a0_311);
and \U$11764 ( \12616 , RIb553528_310, \12351 );
nor \U$11765 ( \12617 , \12615 , \12616 );
nand \U$11766 ( \12618 , \12608 , \12611 , \12614 , \12617 );
nor \U$11767 ( \12619 , \12604 , \12605 , \12618 );
and \U$11768 ( \12620 , \12324 , RIb5533c0_307);
and \U$11769 ( \12621 , RIb553438_308, \12358 );
nor \U$11770 ( \12622 , \12620 , \12621 );
and \U$11771 ( \12623 , RIb5531e0_303, \12338 );
and \U$11772 ( \12624 , RIb553258_304, \12333 );
and \U$11773 ( \12625 , \12327 , RIb553348_306);
and \U$11774 ( \12626 , RIb5532d0_305, \12330 );
nor \U$11775 ( \12627 , \12625 , \12626 );
not \U$11776 ( \12628 , \12627 );
nor \U$11777 ( \12629 , \12623 , \12624 , \12628 );
nand \U$11778 ( \12630 , \12619 , \12622 , \9094 , \12629 );
_DC r3038 ( \12631_nR3038 , \12630 , \12369 );
not \U$11779 ( \12632 , \12631_nR3038 );
nor \U$11780 ( \12633 , \12289 , \12632 );
not \U$11781 ( \12634 , \12562 );
not \U$11782 ( \12635 , \12564 );
nand \U$11783 ( \12636 , \12635 , \12556 );
not \U$11784 ( \12637 , \12636 );
or \U$11785 ( \12638 , \12634 , \12637 );
or \U$11786 ( \12639 , \12636 , \12562 );
nand \U$11787 ( \12640 , \12638 , \12639 );
xnor \U$11788 ( \12641 , \12633 , \12640 );
not \U$11789 ( \12642 , \12641 );
and \U$11790 ( \12643 , \12470_nR3271 , \12485 );
and \U$11791 ( \12644 , \12512 , \12370_nR3379 );
nand \U$11792 ( \12645 , \12470_nR3271 , \12482 );
or \U$11793 ( \12646 , \12440 , \12370_nR3379 );
nand \U$11794 ( \12647 , \12646 , \12516 );
and \U$11795 ( \12648 , \12645 , \12647 );
nor \U$11796 ( \12649 , \12643 , \12644 , \12648 );
and \U$11797 ( \12650 , \12438 , \12558 );
xor \U$11798 ( \12651 , \12558 , \12560 );
nor \U$11799 ( \12652 , \12438 , \12558 );
nor \U$11800 ( \12653 , \12650 , \12651 , \12652 );
and \U$11801 ( \12654 , \12653 , \12562 );
and \U$11802 ( \12655 , \12418_nR349f , \12654 );
not \U$11803 ( \12656 , \12562 );
and \U$11804 ( \12657 , \12419 , \12656 );
or \U$11805 ( \12658 , \12653 , \12562 );
not \U$11806 ( \12659 , \12658 );
nor \U$11807 ( \12660 , \12655 , \12657 , \12659 );
or \U$11808 ( \12661 , \12649 , \12660 );
and \U$11809 ( \12662 , RIb554608_346, \12320 );
and \U$11810 ( \12663 , RIb553ff0_333, \12313 );
and \U$11811 ( \12664 , \12317 , RIb5546f8_348);
and \U$11812 ( \12665 , RIb554680_347, \12309 );
nor \U$11813 ( \12666 , \12664 , \12665 );
and \U$11814 ( \12667 , \12324 , RIb5543b0_341);
and \U$11815 ( \12668 , RIb554338_340, \12327 );
nor \U$11816 ( \12669 , \12667 , \12668 );
and \U$11817 ( \12670 , \12330 , RIb5542c0_339);
and \U$11818 ( \12671 , RIb554248_338, \12333 );
nor \U$11819 ( \12672 , \12670 , \12671 );
and \U$11820 ( \12673 , \12338 , RIb5541d0_337);
and \U$11821 ( \12674 , RIb554158_336, \12341 );
nor \U$11822 ( \12675 , \12673 , \12674 );
nand \U$11823 ( \12676 , \12666 , \12669 , \12672 , \12675 );
nor \U$11824 ( \12677 , \12662 , \12663 , \12676 );
and \U$11825 ( \12678 , \12349 , RIb554590_345);
and \U$11826 ( \12679 , RIb554518_344, \12351 );
nor \U$11827 ( \12680 , \12678 , \12679 );
nand \U$11828 ( \12681 , RIb554770_349, \8856 );
and \U$11829 ( \12682 , RIb5544a0_343, \12356 );
and \U$11830 ( \12683 , RIb554428_342, \12358 );
and \U$11831 ( \12684 , \12360 , RIb5540e0_335);
and \U$11832 ( \12685 , RIb554068_334, \12363 );
nor \U$11833 ( \12686 , \12684 , \12685 );
not \U$11834 ( \12687 , \12686 );
nor \U$11835 ( \12688 , \12682 , \12683 , \12687 );
nand \U$11836 ( \12689 , \12677 , \12680 , \12681 , \12688 );
_DC r2f21 ( \12690_nR2f21 , \12689 , \12369 );
nand \U$11837 ( \12691 , \12690_nR2f21 , \12288 );
and \U$11838 ( \12692 , \12549_nR3150 , \12426 );
and \U$11839 ( \12693 , \12388 , \12631_nR3038 );
nand \U$11840 ( \12694 , \12549_nR3150 , \12381 );
or \U$11841 ( \12695 , \12387 , \12631_nR3038 );
nand \U$11842 ( \12696 , \12695 , \12422 );
and \U$11843 ( \12697 , \12694 , \12696 );
nor \U$11844 ( \12698 , \12692 , \12693 , \12697 );
or \U$11845 ( \12699 , \12691 , \12698 );
nand \U$11846 ( \12700 , \12661 , \12699 );
nand \U$11847 ( \12701 , \12642 , \12700 );
nor \U$11848 ( \12702 , \12603 , \12701 );
and \U$11849 ( \12703 , \12600 , \12702 );
and \U$11850 ( \12704 , \12597 , \12599 );
or \U$11851 ( \12705 , \12703 , \12704 );
xor \U$11852 ( \12706 , \12510 , \12575 );
xor \U$11853 ( \12707 , \12705 , \12706 );
xor \U$11854 ( \12708 , \12597 , \12599 );
xor \U$11855 ( \12709 , \12708 , \12702 );
and \U$11856 ( \12710 , \12640 , \12633 );
not \U$11857 ( \12711 , \12651 );
nor \U$11858 ( \12712 , \12656 , \12711 );
and \U$11859 ( \12713 , \12418_nR349f , \12712 );
or \U$11860 ( \12714 , \12562 , \12370_nR3379 );
nand \U$11861 ( \12715 , \12714 , \12658 );
nand \U$11862 ( \12716 , \12418_nR349f , \12651 );
and \U$11863 ( \12717 , \12715 , \12716 );
and \U$11864 ( \12718 , \12370_nR3379 , \12654 );
nor \U$11865 ( \12719 , \12713 , \12717 , \12718 );
and \U$11866 ( \12720 , \12549_nR3150 , \12485 );
and \U$11867 ( \12721 , \12512 , \12470_nR3271 );
nand \U$11868 ( \12722 , \12549_nR3150 , \12482 );
or \U$11869 ( \12723 , \12440 , \12470_nR3271 );
nand \U$11870 ( \12724 , \12723 , \12516 );
and \U$11871 ( \12725 , \12722 , \12724 );
nor \U$11872 ( \12726 , \12720 , \12721 , \12725 );
nand \U$11873 ( \12727 , \12719 , \12726 );
xor \U$11874 ( \12728 , \8495 , \12070_nR27cf );
xor \U$11875 ( \12729 , \12728 , \12266 );
xor \U$11876 ( \12730 , \8531 , \12100_nR2689 );
xor \U$11877 ( \12731 , \12730 , \12263 );
nor \U$11878 ( \12732 , \12729 , \12731 );
or \U$11879 ( \12733 , \12560 , \12732 );
and \U$11880 ( \12734 , \12727 , \12733 );
and \U$11881 ( \12735 , RIb555148_370, \12341 );
and \U$11882 ( \12736 , RIb555670_381, \12309 );
and \U$11883 ( \12737 , \12349 , RIb555580_379);
and \U$11884 ( \12738 , RIb5555f8_380, \12320 );
nor \U$11885 ( \12739 , \12737 , \12738 );
and \U$11886 ( \12740 , \12360 , RIb5550d0_369);
and \U$11887 ( \12741 , RIb555058_368, \12363 );
nor \U$11888 ( \12742 , \12740 , \12741 );
and \U$11889 ( \12743 , \12317 , RIb5556e8_382);
and \U$11890 ( \12744 , RIb554fe0_367, \12313 );
nor \U$11891 ( \12745 , \12743 , \12744 );
and \U$11892 ( \12746 , \12356 , RIb555490_377);
and \U$11893 ( \12747 , RIb555418_376, \12358 );
nor \U$11894 ( \12748 , \12746 , \12747 );
nand \U$11895 ( \12749 , \12739 , \12742 , \12745 , \12748 );
nor \U$11896 ( \12750 , \12735 , \12736 , \12749 );
and \U$11897 ( \12751 , \12324 , RIb5553a0_375);
and \U$11898 ( \12752 , RIb555508_378, \12351 );
nor \U$11899 ( \12753 , \12751 , \12752 );
and \U$11900 ( \12754 , RIb5551c0_371, \12338 );
and \U$11901 ( \12755 , RIb555238_372, \12333 );
and \U$11902 ( \12756 , \12327 , RIb555328_374);
and \U$11903 ( \12757 , RIb5552b0_373, \12330 );
nor \U$11904 ( \12758 , \12756 , \12757 );
not \U$11905 ( \12759 , \12758 );
nor \U$11906 ( \12760 , \12754 , \12755 , \12759 );
nand \U$11907 ( \12761 , \12750 , \12753 , \9243 , \12760 );
_DC r2e29 ( \12762_nR2e29 , \12761 , \12369 );
not \U$11908 ( \12763 , \12762_nR2e29 );
nor \U$11909 ( \12764 , \12289 , \12763 );
not \U$11910 ( \12765 , \12764 );
and \U$11911 ( \12766 , \12631_nR3038 , \12426 );
and \U$11912 ( \12767 , \12388 , \12690_nR2f21 );
nand \U$11913 ( \12768 , \12631_nR3038 , \12381 );
or \U$11914 ( \12769 , \12387 , \12690_nR2f21 );
nand \U$11915 ( \12770 , \12769 , \12422 );
and \U$11916 ( \12771 , \12768 , \12770 );
nor \U$11917 ( \12772 , \12766 , \12767 , \12771 );
nor \U$11918 ( \12773 , \12765 , \12772 );
nor \U$11919 ( \12774 , \12726 , \12719 );
nor \U$11920 ( \12775 , \12734 , \12773 , \12774 );
xnor \U$11921 ( \12776 , \12691 , \12698 );
not \U$11922 ( \12777 , \12776 );
xor \U$11923 ( \12778 , \12660 , \12649 );
not \U$11924 ( \12779 , \12778 );
and \U$11925 ( \12780 , \12777 , \12779 );
and \U$11926 ( \12781 , \12776 , \12778 );
nor \U$11927 ( \12782 , \12780 , \12781 );
nand \U$11928 ( \12783 , \12775 , \12782 );
not \U$11929 ( \12784 , \12712 );
or \U$11930 ( \12785 , \12784 , \12371 );
not \U$11931 ( \12786 , \12654 );
or \U$11932 ( \12787 , \12492 , \12786 );
or \U$11933 ( \12788 , \12711 , \12371 );
or \U$11934 ( \12789 , \12562 , \12470_nR3271 );
nand \U$11935 ( \12790 , \12789 , \12658 );
nand \U$11936 ( \12791 , \12788 , \12790 );
nand \U$11937 ( \12792 , \12785 , \12787 , \12791 );
not \U$11938 ( \12793 , \12792 );
not \U$11939 ( \12794 , \12733 );
not \U$11940 ( \12795 , \12729 );
not \U$11941 ( \12796 , \12560 );
or \U$11942 ( \12797 , \12795 , \12796 );
or \U$11943 ( \12798 , \12560 , \12729 );
nand \U$11944 ( \12799 , \12797 , \12798 );
xor \U$11945 ( \12800 , \12731 , \12729 );
nor \U$11946 ( \12801 , \12799 , \12800 );
not \U$11947 ( \12802 , \12801 );
nor \U$11948 ( \12803 , \12794 , \12802 );
and \U$11949 ( \12804 , \12803 , \12418_nR349f );
and \U$11950 ( \12805 , \12801 , \12418_nR349f );
nor \U$11951 ( \12806 , \12805 , \12733 );
nor \U$11952 ( \12807 , \12804 , \12806 );
nor \U$11953 ( \12808 , \12793 , \12807 );
and \U$11954 ( \12809 , \12631_nR3038 , \12485 );
and \U$11955 ( \12810 , \12512 , \12549_nR3150 );
nand \U$11956 ( \12811 , \12631_nR3038 , \12482 );
or \U$11957 ( \12812 , \12440 , \12549_nR3150 );
nand \U$11958 ( \12813 , \12812 , \12516 );
and \U$11959 ( \12814 , \12811 , \12813 );
nor \U$11960 ( \12815 , \12809 , \12810 , \12814 );
and \U$11961 ( \12816 , RIb554950_353, \12341 );
and \U$11962 ( \12817 , RIb554ef0_365, \12317 );
and \U$11963 ( \12818 , \12320 , RIb554e00_363);
and \U$11964 ( \12819 , RIb554c98_360, \12356 );
nor \U$11965 ( \12820 , \12818 , \12819 );
and \U$11966 ( \12821 , \12360 , RIb5548d8_352);
and \U$11967 ( \12822 , RIb554860_351, \12363 );
nor \U$11968 ( \12823 , \12821 , \12822 );
and \U$11969 ( \12824 , \12313 , RIb5547e8_350);
and \U$11970 ( \12825 , RIb554c20_359, \12358 );
nor \U$11971 ( \12826 , \12824 , \12825 );
and \U$11972 ( \12827 , \12349 , RIb554d88_362);
and \U$11973 ( \12828 , RIb554d10_361, \12351 );
nor \U$11974 ( \12829 , \12827 , \12828 );
nand \U$11975 ( \12830 , \12820 , \12823 , \12826 , \12829 );
nor \U$11976 ( \12831 , \12816 , \12817 , \12830 );
and \U$11977 ( \12832 , \12309 , RIb554e78_364);
and \U$11978 ( \12833 , RIb554ba8_358, \12324 );
nor \U$11979 ( \12834 , \12832 , \12833 );
and \U$11980 ( \12835 , RIb5549c8_354, \12338 );
and \U$11981 ( \12836 , RIb554a40_355, \12333 );
and \U$11982 ( \12837 , \12327 , RIb554b30_357);
and \U$11983 ( \12838 , RIb554ab8_356, \12330 );
nor \U$11984 ( \12839 , \12837 , \12838 );
not \U$11985 ( \12840 , \12839 );
nor \U$11986 ( \12841 , \12835 , \12836 , \12840 );
nand \U$11987 ( \12842 , \12831 , \12834 , \9326 , \12841 );
_DC r2d1d ( \12843_nR2d1d , \12842 , \12369 );
nand \U$11988 ( \12844 , \12843_nR2d1d , \12288 );
and \U$11989 ( \12845 , \12815 , \12844 );
and \U$11990 ( \12846 , \12690_nR2f21 , \12426 );
and \U$11991 ( \12847 , \12388 , \12762_nR2e29 );
nand \U$11992 ( \12848 , \12690_nR2f21 , \12381 );
or \U$11993 ( \12849 , \12387 , \12762_nR2e29 );
nand \U$11994 ( \12850 , \12849 , \12422 );
and \U$11995 ( \12851 , \12848 , \12850 );
nor \U$11996 ( \12852 , \12846 , \12847 , \12851 );
nor \U$11997 ( \12853 , \12845 , \12852 );
and \U$11998 ( \12854 , \12808 , \12853 );
not \U$11999 ( \12855 , \12733 );
not \U$12000 ( \12856 , \12774 );
nand \U$12001 ( \12857 , \12856 , \12727 );
not \U$12002 ( \12858 , \12857 );
or \U$12003 ( \12859 , \12855 , \12858 );
or \U$12004 ( \12860 , \12857 , \12733 );
nand \U$12005 ( \12861 , \12859 , \12860 );
not \U$12006 ( \12862 , \12861 );
not \U$12007 ( \12863 , \12772 );
not \U$12008 ( \12864 , \12764 );
and \U$12009 ( \12865 , \12863 , \12864 );
and \U$12010 ( \12866 , \12772 , \12764 );
nor \U$12011 ( \12867 , \12865 , \12866 );
nor \U$12012 ( \12868 , \12862 , \12867 );
and \U$12013 ( \12869 , \12854 , \12868 );
xor \U$12014 ( \12870 , \12783 , \12869 );
not \U$12015 ( \12871 , \12700 );
not \U$12016 ( \12872 , \12641 );
or \U$12017 ( \12873 , \12871 , \12872 );
or \U$12018 ( \12874 , \12641 , \12700 );
nand \U$12019 ( \12875 , \12873 , \12874 );
and \U$12020 ( \12876 , \12870 , \12875 );
and \U$12021 ( \12877 , \12783 , \12869 );
or \U$12022 ( \12878 , \12876 , \12877 );
nor \U$12023 ( \12879 , \12710 , \12878 );
not \U$12024 ( \12880 , \12701 );
not \U$12025 ( \12881 , \12602 );
and \U$12026 ( \12882 , \12880 , \12881 );
and \U$12027 ( \12883 , \12701 , \12602 );
nor \U$12028 ( \12884 , \12882 , \12883 );
nor \U$12029 ( \12885 , \12879 , \12884 );
xor \U$12030 ( \12886 , \12709 , \12885 );
and \U$12031 ( \12887 , \12879 , \12884 );
nor \U$12032 ( \12888 , \12887 , \12885 );
and \U$12033 ( \12889 , \12370_nR3379 , \12803 );
or \U$12034 ( \12890 , \12733 , \12418_nR349f );
or \U$12035 ( \12891 , \12733 , \12800 );
nand \U$12036 ( \12892 , \12890 , \12891 );
nand \U$12037 ( \12893 , \12370_nR3379 , \12801 );
and \U$12038 ( \12894 , \12892 , \12893 );
and \U$12039 ( \12895 , \12733 , \12800 );
and \U$12040 ( \12896 , \12418_nR349f , \12895 );
nor \U$12041 ( \12897 , \12889 , \12894 , \12896 );
and \U$12042 ( \12898 , \12470_nR3271 , \12712 );
or \U$12043 ( \12899 , \12562 , \12549_nR3150 );
nand \U$12044 ( \12900 , \12899 , \12658 );
nand \U$12045 ( \12901 , \12470_nR3271 , \12651 );
and \U$12046 ( \12902 , \12900 , \12901 );
and \U$12047 ( \12903 , \12549_nR3150 , \12654 );
nor \U$12048 ( \12904 , \12898 , \12902 , \12903 );
nand \U$12049 ( \12905 , \12897 , \12904 );
xor \U$12050 ( \12906 , \8603 , \12160_nR25a9 );
xor \U$12051 ( \12907 , \12906 , \12257 );
not \U$12052 ( \12908 , \12907 );
xor \U$12053 ( \12909 , \8567 , \12130_nR2687 );
xor \U$12054 ( \12910 , \12909 , \12260 );
not \U$12055 ( \12911 , \12910 );
and \U$12056 ( \12912 , \12908 , \12911 );
or \U$12057 ( \12913 , \12731 , \12912 );
and \U$12058 ( \12914 , \12905 , \12913 );
nor \U$12059 ( \12915 , \12904 , \12897 );
nor \U$12060 ( \12916 , \12914 , \12915 );
not \U$12061 ( \12917 , \12916 );
and \U$12062 ( \12918 , \12690_nR2f21 , \12485 );
and \U$12063 ( \12919 , \12512 , \12631_nR3038 );
nand \U$12064 ( \12920 , \12690_nR2f21 , \12482 );
or \U$12065 ( \12921 , \12440 , \12631_nR3038 );
nand \U$12066 ( \12922 , \12921 , \12516 );
and \U$12067 ( \12923 , \12920 , \12922 );
nor \U$12068 ( \12924 , \12918 , \12919 , \12923 );
and \U$12069 ( \12925 , RIb5566d8_416, \12317 );
and \U$12070 ( \12926 , RIb555fd0_401, \12313 );
and \U$12071 ( \12927 , \12330 , RIb5562a0_407);
and \U$12072 ( \12928 , RIb556228_406, \12333 );
nor \U$12073 ( \12929 , \12927 , \12928 );
and \U$12074 ( \12930 , \12324 , RIb556390_409);
and \U$12075 ( \12931 , RIb556318_408, \12327 );
nor \U$12076 ( \12932 , \12930 , \12931 );
and \U$12077 ( \12933 , \12338 , RIb5561b0_405);
and \U$12078 ( \12934 , RIb556138_404, \12341 );
nor \U$12079 ( \12935 , \12933 , \12934 );
and \U$12080 ( \12936 , \12349 , RIb556570_413);
and \U$12081 ( \12937 , RIb556480_411, \12356 );
nor \U$12082 ( \12938 , \12936 , \12937 );
nand \U$12083 ( \12939 , \12929 , \12932 , \12935 , \12938 );
nor \U$12084 ( \12940 , \12925 , \12926 , \12939 );
and \U$12085 ( \12941 , \12309 , RIb556660_415);
and \U$12086 ( \12942 , RIb5565e8_414, \12320 );
nor \U$12087 ( \12943 , \12941 , \12942 );
and \U$12088 ( \12944 , RIb5564f8_412, \12351 );
and \U$12089 ( \12945 , RIb556408_410, \12358 );
and \U$12090 ( \12946 , \12360 , RIb5560c0_403);
and \U$12091 ( \12947 , RIb556048_402, \12363 );
nor \U$12092 ( \12948 , \12946 , \12947 );
not \U$12093 ( \12949 , \12948 );
nor \U$12094 ( \12950 , \12944 , \12945 , \12949 );
nand \U$12095 ( \12951 , \12940 , \12943 , \9434 , \12950 );
_DC r2c3a ( \12952_nR2c3a , \12951 , \12369 );
nand \U$12096 ( \12953 , \12952_nR2c3a , \12288 );
and \U$12097 ( \12954 , \12924 , \12953 );
and \U$12098 ( \12955 , \12762_nR2e29 , \12426 );
and \U$12099 ( \12956 , \12388 , \12843_nR2d1d );
nand \U$12100 ( \12957 , \12762_nR2e29 , \12381 );
or \U$12101 ( \12958 , \12387 , \12843_nR2d1d );
nand \U$12102 ( \12959 , \12958 , \12422 );
and \U$12103 ( \12960 , \12957 , \12959 );
nor \U$12104 ( \12961 , \12955 , \12956 , \12960 );
nor \U$12105 ( \12962 , \12954 , \12961 );
nand \U$12106 ( \12963 , \12917 , \12962 );
not \U$12107 ( \12964 , \12963 );
not \U$12108 ( \12965 , \12844 );
not \U$12109 ( \12966 , \12852 );
not \U$12110 ( \12967 , \12815 );
and \U$12111 ( \12968 , \12966 , \12967 );
and \U$12112 ( \12969 , \12852 , \12815 );
nor \U$12113 ( \12970 , \12968 , \12969 );
not \U$12114 ( \12971 , \12970 );
or \U$12115 ( \12972 , \12965 , \12971 );
or \U$12116 ( \12973 , \12970 , \12844 );
nand \U$12117 ( \12974 , \12972 , \12973 );
not \U$12118 ( \12975 , \12974 );
not \U$12119 ( \12976 , \12792 );
not \U$12120 ( \12977 , \12807 );
and \U$12121 ( \12978 , \12976 , \12977 );
and \U$12122 ( \12979 , \12792 , \12807 );
nor \U$12123 ( \12980 , \12978 , \12979 );
nor \U$12124 ( \12981 , \12975 , \12980 );
nand \U$12125 ( \12982 , \12964 , \12981 );
not \U$12126 ( \12983 , \12867 );
not \U$12127 ( \12984 , \12861 );
and \U$12128 ( \12985 , \12983 , \12984 );
and \U$12129 ( \12986 , \12867 , \12861 );
nor \U$12130 ( \12987 , \12985 , \12986 );
not \U$12131 ( \12988 , \12987 );
xor \U$12132 ( \12989 , \12808 , \12853 );
nand \U$12133 ( \12990 , \12988 , \12989 );
and \U$12134 ( \12991 , \12982 , \12990 );
not \U$12135 ( \12992 , \12782 );
not \U$12136 ( \12993 , \12775 );
and \U$12137 ( \12994 , \12992 , \12993 );
not \U$12138 ( \12995 , \12783 );
nor \U$12139 ( \12996 , \12994 , \12995 );
nor \U$12140 ( \12997 , \12991 , \12996 );
not \U$12141 ( \12998 , \12778 );
nor \U$12142 ( \12999 , \12998 , \12776 );
xor \U$12143 ( \13000 , \12997 , \12999 );
xor \U$12144 ( \13001 , \12783 , \12869 );
xor \U$12145 ( \13002 , \13001 , \12875 );
and \U$12146 ( \13003 , \13000 , \13002 );
and \U$12147 ( \13004 , \12997 , \12999 );
or \U$12148 ( \13005 , \13003 , \13004 );
xor \U$12149 ( \13006 , \12888 , \13005 );
not \U$12150 ( \13007 , \12989 );
not \U$12151 ( \13008 , \12987 );
or \U$12152 ( \13009 , \13007 , \13008 );
or \U$12153 ( \13010 , \12987 , \12989 );
nand \U$12154 ( \13011 , \13009 , \13010 );
not \U$12155 ( \13012 , \12910 );
not \U$12156 ( \13013 , \12731 );
or \U$12157 ( \13014 , \13012 , \13013 );
or \U$12158 ( \13015 , \12731 , \12910 );
nand \U$12159 ( \13016 , \13014 , \13015 );
xor \U$12160 ( \13017 , \12908 , \12911 );
nor \U$12161 ( \13018 , \13016 , \13017 );
not \U$12162 ( \13019 , \13018 );
not \U$12163 ( \13020 , \12913 );
nor \U$12164 ( \13021 , \13019 , \13020 );
not \U$12165 ( \13022 , \13021 );
or \U$12166 ( \13023 , \13022 , \12419 );
or \U$12167 ( \13024 , \13019 , \12419 );
nand \U$12168 ( \13025 , \13024 , \13020 );
nand \U$12169 ( \13026 , \13023 , \13025 );
not \U$12170 ( \13027 , \12803 );
or \U$12171 ( \13028 , \13027 , \12492 );
not \U$12172 ( \13029 , \12895 );
or \U$12173 ( \13030 , \12371 , \13029 );
or \U$12174 ( \13031 , \12802 , \12492 );
or \U$12175 ( \13032 , \12733 , \12370_nR3379 );
nand \U$12176 ( \13033 , \13032 , \12891 );
nand \U$12177 ( \13034 , \13031 , \13033 );
nand \U$12178 ( \13035 , \13028 , \13030 , \13034 );
and \U$12179 ( \13036 , \13026 , \13035 );
and \U$12180 ( \13037 , \12762_nR2e29 , \12485 );
and \U$12181 ( \13038 , \12512 , \12690_nR2f21 );
nand \U$12182 ( \13039 , \12762_nR2e29 , \12482 );
or \U$12183 ( \13040 , \12440 , \12690_nR2f21 );
nand \U$12184 ( \13041 , \13040 , \12516 );
and \U$12185 ( \13042 , \13039 , \13041 );
nor \U$12186 ( \13043 , \13037 , \13038 , \13042 );
and \U$12187 ( \13044 , \12549_nR3150 , \12712 );
or \U$12188 ( \13045 , \12562 , \12631_nR3038 );
nand \U$12189 ( \13046 , \13045 , \12658 );
nand \U$12190 ( \13047 , \12549_nR3150 , \12651 );
and \U$12191 ( \13048 , \13046 , \13047 );
and \U$12192 ( \13049 , \12631_nR3038 , \12654 );
nor \U$12193 ( \13050 , \13044 , \13048 , \13049 );
xor \U$12194 ( \13051 , \13043 , \13050 );
and \U$12195 ( \13052 , \12843_nR2d1d , \12426 );
and \U$12196 ( \13053 , \12388 , \12952_nR2c3a );
nand \U$12197 ( \13054 , \12843_nR2d1d , \12381 );
or \U$12198 ( \13055 , \12387 , \12952_nR2c3a );
nand \U$12199 ( \13056 , \13055 , \12422 );
and \U$12200 ( \13057 , \13054 , \13056 );
nor \U$12201 ( \13058 , \13052 , \13053 , \13057 );
and \U$12202 ( \13059 , \13051 , \13058 );
and \U$12203 ( \13060 , \13043 , \13050 );
or \U$12204 ( \13061 , \13059 , \13060 );
not \U$12205 ( \13062 , \13061 );
and \U$12206 ( \13063 , \13036 , \13062 );
not \U$12207 ( \13064 , \12913 );
not \U$12208 ( \13065 , \12915 );
nand \U$12209 ( \13066 , \13065 , \12905 );
not \U$12210 ( \13067 , \13066 );
or \U$12211 ( \13068 , \13064 , \13067 );
or \U$12212 ( \13069 , \13066 , \12913 );
nand \U$12213 ( \13070 , \13068 , \13069 );
not \U$12214 ( \13071 , \12953 );
not \U$12215 ( \13072 , \12961 );
not \U$12216 ( \13073 , \12924 );
and \U$12217 ( \13074 , \13072 , \13073 );
and \U$12218 ( \13075 , \12961 , \12924 );
nor \U$12219 ( \13076 , \13074 , \13075 );
not \U$12220 ( \13077 , \13076 );
or \U$12221 ( \13078 , \13071 , \13077 );
or \U$12222 ( \13079 , \13076 , \12953 );
nand \U$12223 ( \13080 , \13078 , \13079 );
and \U$12224 ( \13081 , \13070 , \13080 );
and \U$12225 ( \13082 , \13063 , \13081 );
xor \U$12226 ( \13083 , \13011 , \13082 );
not \U$12227 ( \13084 , \12962 );
not \U$12228 ( \13085 , \12916 );
and \U$12229 ( \13086 , \13084 , \13085 );
and \U$12230 ( \13087 , \12962 , \12916 );
nor \U$12231 ( \13088 , \13086 , \13087 );
not \U$12232 ( \13089 , \12974 );
not \U$12233 ( \13090 , \12980 );
and \U$12234 ( \13091 , \13089 , \13090 );
and \U$12235 ( \13092 , \12974 , \12980 );
nor \U$12236 ( \13093 , \13091 , \13092 );
nand \U$12237 ( \13094 , \13088 , \13093 );
and \U$12238 ( \13095 , \13083 , \13094 );
and \U$12239 ( \13096 , \13011 , \13082 );
or \U$12240 ( \13097 , \13095 , \13096 );
xor \U$12241 ( \13098 , \12854 , \12868 );
xor \U$12242 ( \13099 , \13097 , \13098 );
not \U$12243 ( \13100 , \12990 );
not \U$12244 ( \13101 , \12996 );
not \U$12245 ( \13102 , \12982 );
and \U$12246 ( \13103 , \13101 , \13102 );
and \U$12247 ( \13104 , \12996 , \12982 );
nor \U$12248 ( \13105 , \13103 , \13104 );
not \U$12249 ( \13106 , \13105 );
or \U$12250 ( \13107 , \13100 , \13106 );
or \U$12251 ( \13108 , \13105 , \12990 );
nand \U$12252 ( \13109 , \13107 , \13108 );
and \U$12253 ( \13110 , \13099 , \13109 );
and \U$12254 ( \13111 , \13097 , \13098 );
or \U$12255 ( \13112 , \13110 , \13111 );
xor \U$12256 ( \13113 , \12997 , \12999 );
xor \U$12257 ( \13114 , \13113 , \13002 );
xor \U$12258 ( \13115 , \13112 , \13114 );
not \U$12259 ( \13116 , \12963 );
not \U$12260 ( \13117 , \12981 );
or \U$12261 ( \13118 , \13116 , \13117 );
or \U$12262 ( \13119 , \12981 , \12963 );
nand \U$12263 ( \13120 , \13118 , \13119 );
xor \U$12264 ( \13121 , \13011 , \13082 );
xor \U$12265 ( \13122 , \13121 , \13094 );
and \U$12266 ( \13123 , \13120 , \13122 );
xor \U$12267 ( \13124 , \13036 , \13062 );
xor \U$12268 ( \13125 , \13070 , \13080 );
and \U$12269 ( \13126 , \13124 , \13125 );
xor \U$12270 ( \13127 , \13026 , \13035 );
xor \U$12271 ( \13128 , \13043 , \13050 );
xor \U$12272 ( \13129 , \13128 , \13058 );
not \U$12273 ( \13130 , \13129 );
and \U$12274 ( \13131 , \13127 , \13130 );
and \U$12275 ( \13132 , \12843_nR2d1d , \12485 );
and \U$12276 ( \13133 , \12512 , \12762_nR2e29 );
nand \U$12277 ( \13134 , \12843_nR2d1d , \12482 );
or \U$12278 ( \13135 , \12440 , \12762_nR2e29 );
nand \U$12279 ( \13136 , \13135 , \12516 );
and \U$12280 ( \13137 , \13134 , \13136 );
nor \U$12281 ( \13138 , \13132 , \13133 , \13137 );
and \U$12282 ( \13139 , \12631_nR3038 , \12712 );
or \U$12283 ( \13140 , \12562 , \12690_nR2f21 );
nand \U$12284 ( \13141 , \13140 , \12658 );
nand \U$12285 ( \13142 , \12631_nR3038 , \12651 );
and \U$12286 ( \13143 , \13141 , \13142 );
and \U$12287 ( \13144 , \12690_nR2f21 , \12654 );
nor \U$12288 ( \13145 , \13139 , \13143 , \13144 );
xor \U$12289 ( \13146 , \13138 , \13145 );
and \U$12290 ( \13147 , \12952_nR2c3a , \12426 );
and \U$12291 ( \13148 , RIb555e68_398, \12309 );
and \U$12292 ( \13149 , RIb5557d8_384, \12313 );
and \U$12293 ( \13150 , \12338 , RIb5559b8_388);
and \U$12294 ( \13151 , RIb555940_387, \12341 );
nor \U$12295 ( \13152 , \13150 , \13151 );
and \U$12296 ( \13153 , \12324 , RIb555b98_392);
and \U$12297 ( \13154 , RIb555b20_391, \12327 );
nor \U$12298 ( \13155 , \13153 , \13154 );
and \U$12299 ( \13156 , \12330 , RIb555aa8_390);
and \U$12300 ( \13157 , RIb555a30_389, \12333 );
nor \U$12301 ( \13158 , \13156 , \13157 );
and \U$12302 ( \13159 , \12317 , RIb555ee0_399);
and \U$12303 ( \13160 , RIb555c10_393, \12358 );
nor \U$12304 ( \13161 , \13159 , \13160 );
nand \U$12305 ( \13162 , \13152 , \13155 , \13158 , \13161 );
nor \U$12306 ( \13163 , \13148 , \13149 , \13162 );
and \U$12307 ( \13164 , \12349 , RIb555d78_396);
and \U$12308 ( \13165 , RIb555df0_397, \12320 );
nor \U$12309 ( \13166 , \13164 , \13165 );
and \U$12310 ( \13167 , RIb555d00_395, \12351 );
and \U$12311 ( \13168 , RIb555c88_394, \12356 );
and \U$12312 ( \13169 , \12360 , RIb5558c8_386);
and \U$12313 ( \13170 , RIb555850_385, \12363 );
nor \U$12314 ( \13171 , \13169 , \13170 );
not \U$12315 ( \13172 , \13171 );
nor \U$12316 ( \13173 , \13167 , \13168 , \13172 );
nand \U$12317 ( \13174 , \13163 , \13166 , \9659 , \13173 );
_DC r2b34 ( \13175_nR2b34 , \13174 , \12369 );
and \U$12318 ( \13176 , \12388 , \13175_nR2b34 );
nand \U$12319 ( \13177 , \12952_nR2c3a , \12381 );
or \U$12320 ( \13178 , \12387 , \13175_nR2b34 );
nand \U$12321 ( \13179 , \13178 , \12422 );
and \U$12322 ( \13180 , \13177 , \13179 );
nor \U$12323 ( \13181 , \13147 , \13176 , \13180 );
and \U$12324 ( \13182 , \13146 , \13181 );
and \U$12325 ( \13183 , \13138 , \13145 );
or \U$12326 ( \13184 , \13182 , \13183 );
nand \U$12327 ( \13185 , \12370_nR3379 , \13018 );
or \U$12328 ( \13186 , \12913 , \12418_nR349f );
or \U$12329 ( \13187 , \12913 , \13017 );
nand \U$12330 ( \13188 , \13186 , \13187 );
and \U$12331 ( \13189 , \13185 , \13188 );
and \U$12332 ( \13190 , \12913 , \13017 );
and \U$12333 ( \13191 , \13190 , \12418_nR349f );
and \U$12334 ( \13192 , \12370_nR3379 , \13021 );
nor \U$12335 ( \13193 , \13189 , \13191 , \13192 );
and \U$12336 ( \13194 , \12549_nR3150 , \12803 );
or \U$12337 ( \13195 , \12733 , \12470_nR3271 );
nand \U$12338 ( \13196 , \13195 , \12891 );
nand \U$12339 ( \13197 , \12549_nR3150 , \12801 );
and \U$12340 ( \13198 , \13196 , \13197 );
and \U$12341 ( \13199 , \12470_nR3271 , \12895 );
nor \U$12342 ( \13200 , \13194 , \13198 , \13199 );
nand \U$12343 ( \13201 , \13193 , \13200 );
not \U$12344 ( \13202 , \12221 );
not \U$12345 ( \13203 , \12253 );
nand \U$12346 ( \13204 , \13203 , \12251 );
not \U$12347 ( \13205 , \13204 );
or \U$12348 ( \13206 , \13202 , \13205 );
or \U$12349 ( \13207 , \13204 , \12221 );
nand \U$12350 ( \13208 , \13206 , \13207 );
xor \U$12351 ( \13209 , \8635 , \12190_nR25ab );
xor \U$12352 ( \13210 , \13209 , \12254 );
not \U$12353 ( \13211 , \13210 );
and \U$12354 ( \13212 , \13208 , \13211 );
or \U$12355 ( \13213 , \12907 , \13212 );
and \U$12356 ( \13214 , \13201 , \13213 );
nor \U$12357 ( \13215 , \13200 , \13193 );
nor \U$12358 ( \13216 , \13214 , \13215 );
nor \U$12359 ( \13217 , \13184 , \13216 );
and \U$12360 ( \13218 , \13131 , \13217 );
xor \U$12361 ( \13219 , \13126 , \13218 );
or \U$12362 ( \13220 , \13093 , \13088 );
nand \U$12363 ( \13221 , \13220 , \13094 );
and \U$12364 ( \13222 , \13219 , \13221 );
and \U$12365 ( \13223 , \13126 , \13218 );
or \U$12366 ( \13224 , \13222 , \13223 );
xor \U$12367 ( \13225 , \13011 , \13082 );
xor \U$12368 ( \13226 , \13225 , \13094 );
and \U$12369 ( \13227 , \13224 , \13226 );
and \U$12370 ( \13228 , \13120 , \13224 );
or \U$12371 ( \13229 , \13123 , \13227 , \13228 );
xor \U$12372 ( \13230 , \13097 , \13098 );
xor \U$12373 ( \13231 , \13230 , \13109 );
xor \U$12374 ( \13232 , \13229 , \13231 );
xor \U$12375 ( \13233 , \13011 , \13082 );
xor \U$12376 ( \13234 , \13233 , \13094 );
xor \U$12377 ( \13235 , \13120 , \13224 );
xor \U$12378 ( \13236 , \13234 , \13235 );
nand \U$12379 ( \13237 , \13175_nR2b34 , \12288 );
not \U$12380 ( \13238 , \13237 );
xor \U$12381 ( \13239 , \13127 , \13130 );
not \U$12382 ( \13240 , \13239 );
or \U$12383 ( \13241 , \13238 , \13240 );
xnor \U$12384 ( \13242 , \13216 , \13184 );
nand \U$12385 ( \13243 , \13241 , \13242 );
or \U$12386 ( \13244 , \12907 , \13210 );
nand \U$12387 ( \13245 , \13210 , \12907 );
nand \U$12388 ( \13246 , \13244 , \13245 );
xor \U$12389 ( \13247 , \13208 , \13211 );
nor \U$12390 ( \13248 , \13246 , \13247 );
not \U$12391 ( \13249 , \13248 );
not \U$12392 ( \13250 , \13213 );
nor \U$12393 ( \13251 , \13249 , \13250 );
not \U$12394 ( \13252 , \13251 );
or \U$12395 ( \13253 , \13252 , \12419 );
or \U$12396 ( \13254 , \13249 , \12419 );
nand \U$12397 ( \13255 , \13254 , \13250 );
nand \U$12398 ( \13256 , \13253 , \13255 );
not \U$12399 ( \13257 , \13256 );
nand \U$12400 ( \13258 , \12470_nR3271 , \13018 );
or \U$12401 ( \13259 , \12913 , \12370_nR3379 );
nand \U$12402 ( \13260 , \13259 , \13187 );
and \U$12403 ( \13261 , \13258 , \13260 );
and \U$12404 ( \13262 , \13190 , \12370_nR3379 );
and \U$12405 ( \13263 , \12470_nR3271 , \13021 );
nor \U$12406 ( \13264 , \13261 , \13262 , \13263 );
nor \U$12407 ( \13265 , \13257 , \13264 );
not \U$12408 ( \13266 , \13265 );
and \U$12409 ( \13267 , \12690_nR2f21 , \12712 );
or \U$12410 ( \13268 , \12562 , \12762_nR2e29 );
nand \U$12411 ( \13269 , \13268 , \12658 );
nand \U$12412 ( \13270 , \12690_nR2f21 , \12651 );
and \U$12413 ( \13271 , \13269 , \13270 );
and \U$12414 ( \13272 , \12762_nR2e29 , \12654 );
nor \U$12415 ( \13273 , \13267 , \13271 , \13272 );
and \U$12416 ( \13274 , \12631_nR3038 , \12803 );
or \U$12417 ( \13275 , \12733 , \12549_nR3150 );
nand \U$12418 ( \13276 , \13275 , \12891 );
nand \U$12419 ( \13277 , \12631_nR3038 , \12801 );
and \U$12420 ( \13278 , \13276 , \13277 );
and \U$12421 ( \13279 , \12549_nR3150 , \12895 );
nor \U$12422 ( \13280 , \13274 , \13278 , \13279 );
xor \U$12423 ( \13281 , \13273 , \13280 );
and \U$12424 ( \13282 , \12952_nR2c3a , \12485 );
and \U$12425 ( \13283 , \12512 , \12843_nR2d1d );
nand \U$12426 ( \13284 , \12952_nR2c3a , \12482 );
or \U$12427 ( \13285 , \12440 , \12843_nR2d1d );
nand \U$12428 ( \13286 , \13285 , \12516 );
and \U$12429 ( \13287 , \13284 , \13286 );
nor \U$12430 ( \13288 , \13282 , \13283 , \13287 );
and \U$12431 ( \13289 , \13281 , \13288 );
and \U$12432 ( \13290 , \13273 , \13280 );
or \U$12433 ( \13291 , \13289 , \13290 );
nor \U$12434 ( \13292 , \13266 , \13291 );
not \U$12435 ( \13293 , \13292 );
and \U$12436 ( \13294 , RIb557128_438, \12341 );
and \U$12437 ( \13295 , RIb557560_447, \12349 );
and \U$12438 ( \13296 , \12356 , RIb557470_445);
and \U$12439 ( \13297 , RIb5573f8_444, \12358 );
nor \U$12440 ( \13298 , \13296 , \13297 );
and \U$12441 ( \13299 , \12317 , RIb5576c8_450);
and \U$12442 ( \13300 , RIb5570b0_437, \12360 );
nor \U$12443 ( \13301 , \13299 , \13300 );
and \U$12444 ( \13302 , \12313 , RIb556fc0_435);
and \U$12445 ( \13303 , RIb557038_436, \12363 );
nor \U$12446 ( \13304 , \13302 , \13303 );
and \U$12447 ( \13305 , \12309 , RIb557650_449);
and \U$12448 ( \13306 , RIb5575d8_448, \12320 );
nor \U$12449 ( \13307 , \13305 , \13306 );
nand \U$12450 ( \13308 , \13298 , \13301 , \13304 , \13307 );
nor \U$12451 ( \13309 , \13294 , \13295 , \13308 );
and \U$12452 ( \13310 , \12324 , RIb557380_443);
and \U$12453 ( \13311 , RIb5574e8_446, \12351 );
nor \U$12454 ( \13312 , \13310 , \13311 );
nand \U$12455 ( \13313 , RIb557740_451, \8856 );
and \U$12456 ( \13314 , RIb5571a0_439, \12338 );
and \U$12457 ( \13315 , RIb557218_440, \12333 );
and \U$12458 ( \13316 , \12327 , RIb557308_442);
and \U$12459 ( \13317 , RIb557290_441, \12330 );
nor \U$12460 ( \13318 , \13316 , \13317 );
not \U$12461 ( \13319 , \13318 );
nor \U$12462 ( \13320 , \13314 , \13315 , \13319 );
nand \U$12463 ( \13321 , \13309 , \13312 , \13313 , \13320 );
_DC r2a51 ( \13322_nR2a51 , \13321 , \12369 );
nand \U$12464 ( \13323 , \13322_nR2a51 , \12288 );
not \U$12465 ( \13324 , \13323 );
not \U$12466 ( \13325 , \13213 );
not \U$12467 ( \13326 , \13215 );
nand \U$12468 ( \13327 , \13326 , \13201 );
not \U$12469 ( \13328 , \13327 );
or \U$12470 ( \13329 , \13325 , \13328 );
or \U$12471 ( \13330 , \13327 , \13213 );
nand \U$12472 ( \13331 , \13329 , \13330 );
xor \U$12473 ( \13332 , \13138 , \13145 );
xor \U$12474 ( \13333 , \13332 , \13181 );
not \U$12475 ( \13334 , \13333 );
and \U$12476 ( \13335 , \13331 , \13334 );
nor \U$12477 ( \13336 , \13324 , \13335 );
nor \U$12478 ( \13337 , \13293 , \13336 );
xor \U$12479 ( \13338 , \13243 , \13337 );
xor \U$12480 ( \13339 , \13124 , \13125 );
and \U$12481 ( \13340 , \13338 , \13339 );
and \U$12482 ( \13341 , \13243 , \13337 );
or \U$12483 ( \13342 , \13340 , \13341 );
xor \U$12484 ( \13343 , \13063 , \13081 );
xor \U$12485 ( \13344 , \13342 , \13343 );
xor \U$12486 ( \13345 , \13126 , \13218 );
xor \U$12487 ( \13346 , \13345 , \13221 );
and \U$12488 ( \13347 , \13344 , \13346 );
and \U$12489 ( \13348 , \13342 , \13343 );
or \U$12490 ( \13349 , \13347 , \13348 );
xor \U$12491 ( \13350 , \13236 , \13349 );
xor \U$12492 ( \13351 , \13342 , \13343 );
xor \U$12493 ( \13352 , \13351 , \13346 );
xor \U$12494 ( \13353 , \13331 , \13334 );
not \U$12495 ( \13354 , \13353 );
not \U$12496 ( \13355 , \13323 );
and \U$12497 ( \13356 , \13354 , \13355 );
and \U$12498 ( \13357 , \13353 , \13323 );
nor \U$12499 ( \13358 , \13356 , \13357 );
not \U$12500 ( \13359 , \13358 );
or \U$12501 ( \13360 , \13291 , \13265 );
and \U$12502 ( \13361 , RIb556ed0_433, \12317 );
and \U$12503 ( \13362 , RIb5567c8_418, \12313 );
and \U$12504 ( \13363 , \12330 , RIb556a98_424);
and \U$12505 ( \13364 , RIb556a20_423, \12333 );
nor \U$12506 ( \13365 , \13363 , \13364 );
and \U$12507 ( \13366 , \12324 , RIb556b88_426);
and \U$12508 ( \13367 , RIb556b10_425, \12327 );
nor \U$12509 ( \13368 , \13366 , \13367 );
and \U$12510 ( \13369 , \12338 , RIb5569a8_422);
and \U$12511 ( \13370 , RIb556930_421, \12341 );
nor \U$12512 ( \13371 , \13369 , \13370 );
and \U$12513 ( \13372 , \12356 , RIb556c78_428);
and \U$12514 ( \13373 , RIb556c00_427, \12358 );
nor \U$12515 ( \13374 , \13372 , \13373 );
nand \U$12516 ( \13375 , \13365 , \13368 , \13371 , \13374 );
nor \U$12517 ( \13376 , \13361 , \13362 , \13375 );
and \U$12518 ( \13377 , \12309 , RIb556e58_432);
and \U$12519 ( \13378 , RIb556de0_431, \12320 );
nor \U$12520 ( \13379 , \13377 , \13378 );
and \U$12521 ( \13380 , RIb556d68_430, \12349 );
and \U$12522 ( \13381 , RIb556cf0_429, \12351 );
and \U$12523 ( \13382 , \12360 , RIb5568b8_420);
and \U$12524 ( \13383 , RIb556840_419, \12363 );
nor \U$12525 ( \13384 , \13382 , \13383 );
not \U$12526 ( \13385 , \13384 );
nor \U$12527 ( \13386 , \13380 , \13381 , \13385 );
nand \U$12528 ( \13387 , \13376 , \13379 , \9871 , \13386 );
_DC r2979 ( \13388_nR2979 , \13387 , \12369 );
nand \U$12529 ( \13389 , \13388_nR2979 , \12288 );
and \U$12530 ( \13390 , \13175_nR2b34 , \12426 );
and \U$12531 ( \13391 , \12388 , \13322_nR2a51 );
nand \U$12532 ( \13392 , \13175_nR2b34 , \12381 );
or \U$12533 ( \13393 , \12387 , \13322_nR2a51 );
nand \U$12534 ( \13394 , \13393 , \12422 );
and \U$12535 ( \13395 , \13392 , \13394 );
nor \U$12536 ( \13396 , \13390 , \13391 , \13395 );
or \U$12537 ( \13397 , \13389 , \13396 );
nand \U$12538 ( \13398 , \13265 , \13291 );
nand \U$12539 ( \13399 , \13360 , \13397 , \13398 );
nand \U$12540 ( \13400 , \13359 , \13399 );
not \U$12541 ( \13401 , \13264 );
not \U$12542 ( \13402 , \13256 );
and \U$12543 ( \13403 , \13401 , \13402 );
and \U$12544 ( \13404 , \13264 , \13256 );
nor \U$12545 ( \13405 , \13403 , \13404 );
xor \U$12546 ( \13406 , \13273 , \13280 );
xor \U$12547 ( \13407 , \13406 , \13288 );
and \U$12548 ( \13408 , \13405 , \13407 );
xnor \U$12549 ( \13409 , \13389 , \13396 );
xor \U$12550 ( \13410 , \13273 , \13280 );
xor \U$12551 ( \13411 , \13410 , \13288 );
and \U$12552 ( \13412 , \13409 , \13411 );
and \U$12553 ( \13413 , \13405 , \13409 );
or \U$12554 ( \13414 , \13408 , \13412 , \13413 );
not \U$12555 ( \13415 , \13414 );
not \U$12556 ( \13416 , \13175_nR2b34 );
or \U$12557 ( \13417 , \12486 , \13416 );
and \U$12558 ( \13418 , \12512 , \12952_nR2c3a );
nand \U$12559 ( \13419 , \13175_nR2b34 , \12482 );
or \U$12560 ( \13420 , \12440 , \12952_nR2c3a );
nand \U$12561 ( \13421 , \13420 , \12516 );
and \U$12562 ( \13422 , \13419 , \13421 );
nor \U$12563 ( \13423 , \13418 , \13422 );
nand \U$12564 ( \13424 , \13417 , \13423 );
and \U$12565 ( \13425 , \12690_nR2f21 , \12803 );
or \U$12566 ( \13426 , \12733 , \12631_nR3038 );
nand \U$12567 ( \13427 , \13426 , \12891 );
nand \U$12568 ( \13428 , \12690_nR2f21 , \12801 );
and \U$12569 ( \13429 , \13427 , \13428 );
and \U$12570 ( \13430 , \12631_nR3038 , \12895 );
nor \U$12571 ( \13431 , \13425 , \13429 , \13430 );
and \U$12572 ( \13432 , \12762_nR2e29 , \12712 );
or \U$12573 ( \13433 , \12562 , \12843_nR2d1d );
nand \U$12574 ( \13434 , \13433 , \12658 );
nand \U$12575 ( \13435 , \12762_nR2e29 , \12651 );
and \U$12576 ( \13436 , \13434 , \13435 );
and \U$12577 ( \13437 , \12843_nR2d1d , \12654 );
nor \U$12578 ( \13438 , \13432 , \13436 , \13437 );
nand \U$12579 ( \13439 , \13431 , \13438 );
and \U$12580 ( \13440 , \13424 , \13439 );
nor \U$12581 ( \13441 , \13438 , \13431 );
nor \U$12582 ( \13442 , \13440 , \13441 );
nand \U$12583 ( \13443 , \12370_nR3379 , \13248 );
or \U$12584 ( \13444 , \13213 , \12418_nR349f );
or \U$12585 ( \13445 , \13213 , \13247 );
nand \U$12586 ( \13446 , \13444 , \13445 );
and \U$12587 ( \13447 , \13443 , \13446 );
and \U$12588 ( \13448 , \13213 , \13247 );
and \U$12589 ( \13449 , \13448 , \12418_nR349f );
and \U$12590 ( \13450 , \12370_nR3379 , \13251 );
nor \U$12591 ( \13451 , \13447 , \13449 , \13450 );
xor \U$12592 ( \13452 , \13451 , \13208 );
nand \U$12593 ( \13453 , \12549_nR3150 , \13018 );
or \U$12594 ( \13454 , \12913 , \12470_nR3271 );
nand \U$12595 ( \13455 , \13454 , \13187 );
and \U$12596 ( \13456 , \13453 , \13455 );
and \U$12597 ( \13457 , \13190 , \12470_nR3271 );
and \U$12598 ( \13458 , \12549_nR3150 , \13021 );
nor \U$12599 ( \13459 , \13456 , \13457 , \13458 );
and \U$12600 ( \13460 , \13452 , \13459 );
and \U$12601 ( \13461 , \13451 , \13208 );
or \U$12602 ( \13462 , \13460 , \13461 );
nor \U$12603 ( \13463 , \13442 , \13462 );
nand \U$12604 ( \13464 , \13415 , \13463 );
xor \U$12605 ( \13465 , \13400 , \13464 );
xor \U$12606 ( \13466 , \13242 , \13239 );
not \U$12607 ( \13467 , \13466 );
not \U$12608 ( \13468 , \13237 );
and \U$12609 ( \13469 , \13467 , \13468 );
and \U$12610 ( \13470 , \13466 , \13237 );
nor \U$12611 ( \13471 , \13469 , \13470 );
and \U$12612 ( \13472 , \13465 , \13471 );
and \U$12613 ( \13473 , \13400 , \13464 );
or \U$12614 ( \13474 , \13472 , \13473 );
not \U$12615 ( \13475 , \13131 );
not \U$12616 ( \13476 , \13237 );
nor \U$12617 ( \13477 , \13476 , \13217 );
not \U$12618 ( \13478 , \13477 );
and \U$12619 ( \13479 , \13475 , \13478 );
and \U$12620 ( \13480 , \13131 , \13477 );
nor \U$12621 ( \13481 , \13479 , \13480 );
nor \U$12622 ( \13482 , \13474 , \13481 );
not \U$12623 ( \13483 , \13482 );
xor \U$12624 ( \13484 , \13243 , \13337 );
xor \U$12625 ( \13485 , \13484 , \13339 );
not \U$12626 ( \13486 , \13485 );
and \U$12627 ( \13487 , \13483 , \13486 );
and \U$12628 ( \13488 , \13474 , \13481 );
nor \U$12629 ( \13489 , \13487 , \13488 );
xor \U$12630 ( \13490 , \13352 , \13489 );
not \U$12631 ( \13491 , \13485 );
nor \U$12632 ( \13492 , \13482 , \13488 );
not \U$12633 ( \13493 , \13492 );
or \U$12634 ( \13494 , \13491 , \13493 );
or \U$12635 ( \13495 , \13492 , \13485 );
nand \U$12636 ( \13496 , \13494 , \13495 );
and \U$12637 ( \13497 , \12762_nR2e29 , \12803 );
or \U$12638 ( \13498 , \12733 , \12690_nR2f21 );
nand \U$12639 ( \13499 , \13498 , \12891 );
nand \U$12640 ( \13500 , \12762_nR2e29 , \12801 );
and \U$12641 ( \13501 , \13499 , \13500 );
and \U$12642 ( \13502 , \12690_nR2f21 , \12895 );
nor \U$12643 ( \13503 , \13497 , \13501 , \13502 );
nand \U$12644 ( \13504 , \12631_nR3038 , \13018 );
or \U$12645 ( \13505 , \12913 , \12549_nR3150 );
nand \U$12646 ( \13506 , \13505 , \13187 );
and \U$12647 ( \13507 , \13504 , \13506 );
and \U$12648 ( \13508 , \13190 , \12549_nR3150 );
and \U$12649 ( \13509 , \12631_nR3038 , \13021 );
nor \U$12650 ( \13510 , \13507 , \13508 , \13509 );
xor \U$12651 ( \13511 , \13503 , \13510 );
and \U$12652 ( \13512 , \12843_nR2d1d , \12712 );
or \U$12653 ( \13513 , \12562 , \12952_nR2c3a );
nand \U$12654 ( \13514 , \13513 , \12658 );
nand \U$12655 ( \13515 , \12843_nR2d1d , \12651 );
and \U$12656 ( \13516 , \13514 , \13515 );
and \U$12657 ( \13517 , \12952_nR2c3a , \12654 );
nor \U$12658 ( \13518 , \13512 , \13516 , \13517 );
and \U$12659 ( \13519 , \13511 , \13518 );
and \U$12660 ( \13520 , \13503 , \13510 );
or \U$12661 ( \13521 , \13519 , \13520 );
nand \U$12662 ( \13522 , \12470_nR3271 , \13248 );
or \U$12663 ( \13523 , \13213 , \12370_nR3379 );
nand \U$12664 ( \13524 , \13523 , \13445 );
and \U$12665 ( \13525 , \13522 , \13524 );
and \U$12666 ( \13526 , \13448 , \12370_nR3379 );
and \U$12667 ( \13527 , \12470_nR3271 , \13251 );
nor \U$12668 ( \13528 , \13525 , \13526 , \13527 );
not \U$12669 ( \13529 , \13528 );
not \U$12670 ( \13530 , \13208 );
or \U$12671 ( \13531 , \13530 , \12418_nR349f );
or \U$12672 ( \13532 , \8697 , \12220_nR2433 );
nand \U$12673 ( \13533 , \13532 , \12221 );
nor \U$12674 ( \13534 , \13530 , \13533 );
not \U$12675 ( \13535 , \13534 );
nand \U$12676 ( \13536 , \13208 , \13535 );
nand \U$12677 ( \13537 , \13531 , \13536 );
nand \U$12678 ( \13538 , \13529 , \13537 );
xor \U$12679 ( \13539 , \13521 , \13538 );
and \U$12680 ( \13540 , \13322_nR2a51 , \12485 );
and \U$12681 ( \13541 , \12512 , \13175_nR2b34 );
nand \U$12682 ( \13542 , \13322_nR2a51 , \12482 );
or \U$12683 ( \13543 , \12440 , \13175_nR2b34 );
nand \U$12684 ( \13544 , \13543 , \12516 );
and \U$12685 ( \13545 , \13542 , \13544 );
nor \U$12686 ( \13546 , \13540 , \13541 , \13545 );
and \U$12687 ( \13547 , RIb557920_455, \12341 );
and \U$12688 ( \13548 , RIb557e48_466, \12309 );
and \U$12689 ( \13549 , \12320 , RIb557dd0_465);
and \U$12690 ( \13550 , RIb557bf0_461, \12358 );
nor \U$12691 ( \13551 , \13549 , \13550 );
and \U$12692 ( \13552 , \12360 , RIb5578a8_454);
and \U$12693 ( \13553 , RIb557830_453, \12363 );
nor \U$12694 ( \13554 , \13552 , \13553 );
and \U$12695 ( \13555 , \12317 , RIb557ec0_467);
and \U$12696 ( \13556 , RIb5577b8_452, \12313 );
nor \U$12697 ( \13557 , \13555 , \13556 );
and \U$12698 ( \13558 , \12324 , RIb557b78_460);
and \U$12699 ( \13559 , RIb557b00_459, \12327 );
nor \U$12700 ( \13560 , \13558 , \13559 );
nand \U$12701 ( \13561 , \13551 , \13554 , \13557 , \13560 );
nor \U$12702 ( \13562 , \13547 , \13548 , \13561 );
and \U$12703 ( \13563 , \12349 , RIb557d58_464);
and \U$12704 ( \13564 , RIb557ce0_463, \12351 );
nor \U$12705 ( \13565 , \13563 , \13564 );
nand \U$12706 ( \13566 , RIb557f38_468, \8856 );
and \U$12707 ( \13567 , RIb557998_456, \12338 );
and \U$12708 ( \13568 , RIb557a10_457, \12333 );
and \U$12709 ( \13569 , \12330 , RIb557a88_458);
and \U$12710 ( \13570 , RIb557c68_462, \12356 );
nor \U$12711 ( \13571 , \13569 , \13570 );
not \U$12712 ( \13572 , \13571 );
nor \U$12713 ( \13573 , \13567 , \13568 , \13572 );
nand \U$12714 ( \13574 , \13562 , \13565 , \13566 , \13573 );
_DC r27ee ( \13575_nR27ee , \13574 , \12369 );
nand \U$12715 ( \13576 , \13575_nR27ee , \12288 );
and \U$12716 ( \13577 , \13546 , \13576 );
and \U$12717 ( \13578 , \13388_nR2979 , \12426 );
and \U$12718 ( \13579 , RIb5586b8_484, \12317 );
and \U$12719 ( \13580 , RIb557fb0_469, \12313 );
and \U$12720 ( \13581 , \12330 , RIb558280_475);
and \U$12721 ( \13582 , RIb558208_474, \12333 );
nor \U$12722 ( \13583 , \13581 , \13582 );
and \U$12723 ( \13584 , \12324 , RIb558370_477);
and \U$12724 ( \13585 , RIb5582f8_476, \12327 );
nor \U$12725 ( \13586 , \13584 , \13585 );
and \U$12726 ( \13587 , \12338 , RIb558190_473);
and \U$12727 ( \13588 , RIb558118_472, \12341 );
nor \U$12728 ( \13589 , \13587 , \13588 );
and \U$12729 ( \13590 , \12320 , RIb5585c8_482);
and \U$12730 ( \13591 , RIb5583e8_478, \12358 );
nor \U$12731 ( \13592 , \13590 , \13591 );
nand \U$12732 ( \13593 , \13583 , \13586 , \13589 , \13592 );
nor \U$12733 ( \13594 , \13579 , \13580 , \13593 );
and \U$12734 ( \13595 , \12309 , RIb558640_483);
and \U$12735 ( \13596 , RIb558550_481, \12349 );
nor \U$12736 ( \13597 , \13595 , \13596 );
nand \U$12737 ( \13598 , RIb558730_485, \8856 );
and \U$12738 ( \13599 , RIb5584d8_480, \12351 );
and \U$12739 ( \13600 , RIb558460_479, \12356 );
and \U$12740 ( \13601 , \12360 , RIb5580a0_471);
and \U$12741 ( \13602 , RIb558028_470, \12363 );
nor \U$12742 ( \13603 , \13601 , \13602 );
not \U$12743 ( \13604 , \13603 );
nor \U$12744 ( \13605 , \13599 , \13600 , \13604 );
nand \U$12745 ( \13606 , \13594 , \13597 , \13598 , \13605 );
_DC r28bb ( \13607_nR28bb , \13606 , \12369 );
and \U$12746 ( \13608 , \12388 , \13607_nR28bb );
nand \U$12747 ( \13609 , \13388_nR2979 , \12381 );
or \U$12748 ( \13610 , \12387 , \13607_nR28bb );
nand \U$12749 ( \13611 , \13610 , \12422 );
and \U$12750 ( \13612 , \13609 , \13611 );
nor \U$12751 ( \13613 , \13578 , \13608 , \13612 );
nor \U$12752 ( \13614 , \13577 , \13613 );
not \U$12753 ( \13615 , \13614 );
and \U$12754 ( \13616 , \13539 , \13615 );
and \U$12755 ( \13617 , \13521 , \13538 );
or \U$12756 ( \13618 , \13616 , \13617 );
not \U$12757 ( \13619 , \13618 );
nand \U$12758 ( \13620 , \13607_nR28bb , \12288 );
and \U$12759 ( \13621 , \13322_nR2a51 , \12426 );
and \U$12760 ( \13622 , \12388 , \13388_nR2979 );
nand \U$12761 ( \13623 , \13322_nR2a51 , \12381 );
or \U$12762 ( \13624 , \12387 , \13388_nR2979 );
nand \U$12763 ( \13625 , \13624 , \12422 );
and \U$12764 ( \13626 , \13623 , \13625 );
nor \U$12765 ( \13627 , \13621 , \13622 , \13626 );
xor \U$12766 ( \13628 , \13620 , \13627 );
not \U$12767 ( \13629 , \13628 );
not \U$12768 ( \13630 , \13629 );
and \U$12769 ( \13631 , \13619 , \13630 );
and \U$12770 ( \13632 , \13618 , \13629 );
xor \U$12771 ( \13633 , \13273 , \13280 );
xor \U$12772 ( \13634 , \13633 , \13288 );
xor \U$12773 ( \13635 , \13405 , \13409 );
xor \U$12774 ( \13636 , \13634 , \13635 );
nor \U$12775 ( \13637 , \13632 , \13636 );
nor \U$12776 ( \13638 , \13631 , \13637 );
not \U$12777 ( \13639 , \13414 );
not \U$12778 ( \13640 , \13463 );
and \U$12779 ( \13641 , \13639 , \13640 );
and \U$12780 ( \13642 , \13414 , \13463 );
nor \U$12781 ( \13643 , \13641 , \13642 );
xor \U$12782 ( \13644 , \13638 , \13643 );
not \U$12783 ( \13645 , \13358 );
not \U$12784 ( \13646 , \13399 );
and \U$12785 ( \13647 , \13645 , \13646 );
and \U$12786 ( \13648 , \13358 , \13399 );
nor \U$12787 ( \13649 , \13647 , \13648 );
and \U$12788 ( \13650 , \13644 , \13649 );
and \U$12789 ( \13651 , \13638 , \13643 );
or \U$12790 ( \13652 , \13650 , \13651 );
not \U$12791 ( \13653 , \13336 );
not \U$12792 ( \13654 , \13292 );
and \U$12793 ( \13655 , \13653 , \13654 );
and \U$12794 ( \13656 , \13336 , \13292 );
nor \U$12795 ( \13657 , \13655 , \13656 );
xor \U$12796 ( \13658 , \13652 , \13657 );
xor \U$12797 ( \13659 , \13400 , \13464 );
xor \U$12798 ( \13660 , \13659 , \13471 );
and \U$12799 ( \13661 , \13658 , \13660 );
and \U$12800 ( \13662 , \13652 , \13657 );
or \U$12801 ( \13663 , \13661 , \13662 );
xor \U$12802 ( \13664 , \13496 , \13663 );
and \U$12803 ( \13665 , \12952_nR2c3a , \12712 );
or \U$12804 ( \13666 , \12562 , \13175_nR2b34 );
nand \U$12805 ( \13667 , \13666 , \12658 );
nand \U$12806 ( \13668 , \12952_nR2c3a , \12651 );
and \U$12807 ( \13669 , \13667 , \13668 );
and \U$12808 ( \13670 , \13175_nR2b34 , \12654 );
nor \U$12809 ( \13671 , \13665 , \13669 , \13670 );
and \U$12810 ( \13672 , \12843_nR2d1d , \12803 );
or \U$12811 ( \13673 , \12733 , \12762_nR2e29 );
nand \U$12812 ( \13674 , \13673 , \12891 );
nand \U$12813 ( \13675 , \12843_nR2d1d , \12801 );
and \U$12814 ( \13676 , \13674 , \13675 );
and \U$12815 ( \13677 , \12762_nR2e29 , \12895 );
nor \U$12816 ( \13678 , \13672 , \13676 , \13677 );
xor \U$12817 ( \13679 , \13671 , \13678 );
and \U$12818 ( \13680 , \13388_nR2979 , \12485 );
and \U$12819 ( \13681 , \12512 , \13322_nR2a51 );
nand \U$12820 ( \13682 , \13388_nR2979 , \12482 );
or \U$12821 ( \13683 , \12440 , \13322_nR2a51 );
nand \U$12822 ( \13684 , \13683 , \12516 );
and \U$12823 ( \13685 , \13682 , \13684 );
nor \U$12824 ( \13686 , \13680 , \13681 , \13685 );
and \U$12825 ( \13687 , \13679 , \13686 );
and \U$12826 ( \13688 , \13671 , \13678 );
or \U$12827 ( \13689 , \13687 , \13688 );
nand \U$12828 ( \13690 , \12549_nR3150 , \13248 );
or \U$12829 ( \13691 , \13213 , \12470_nR3271 );
nand \U$12830 ( \13692 , \13691 , \13445 );
and \U$12831 ( \13693 , \13690 , \13692 );
and \U$12832 ( \13694 , \13448 , \12470_nR3271 );
and \U$12833 ( \13695 , \12549_nR3150 , \13251 );
nor \U$12834 ( \13696 , \13693 , \13694 , \13695 );
not \U$12835 ( \13697 , \13696 );
not \U$12836 ( \13698 , \13536 );
and \U$12837 ( \13699 , \12419 , \13698 );
and \U$12838 ( \13700 , \13534 , \12371 );
nand \U$12839 ( \13701 , \13533 , \13530 );
not \U$12840 ( \13702 , \13701 );
and \U$12841 ( \13703 , \12418_nR349f , \13702 );
nor \U$12842 ( \13704 , \13699 , \13700 , \13703 );
not \U$12843 ( \13705 , \13704 );
and \U$12844 ( \13706 , \13697 , \13705 );
and \U$12845 ( \13707 , \13696 , \13704 );
nand \U$12846 ( \13708 , \12690_nR2f21 , \13018 );
or \U$12847 ( \13709 , \12913 , \12631_nR3038 );
nand \U$12848 ( \13710 , \13709 , \13187 );
and \U$12849 ( \13711 , \13708 , \13710 );
and \U$12850 ( \13712 , \13190 , \12631_nR3038 );
and \U$12851 ( \13713 , \12690_nR2f21 , \13021 );
nor \U$12852 ( \13714 , \13711 , \13712 , \13713 );
nor \U$12853 ( \13715 , \13707 , \13714 );
nor \U$12854 ( \13716 , \13706 , \13715 );
nor \U$12855 ( \13717 , \13689 , \13716 );
not \U$12856 ( \13718 , \13441 );
nand \U$12857 ( \13719 , \13718 , \13439 );
not \U$12858 ( \13720 , \13719 );
not \U$12859 ( \13721 , \13424 );
or \U$12860 ( \13722 , \13720 , \13721 );
or \U$12861 ( \13723 , \13424 , \13719 );
nand \U$12862 ( \13724 , \13722 , \13723 );
xor \U$12863 ( \13725 , \13717 , \13724 );
not \U$12864 ( \13726 , \13576 );
not \U$12865 ( \13727 , \13613 );
not \U$12866 ( \13728 , \13546 );
and \U$12867 ( \13729 , \13727 , \13728 );
and \U$12868 ( \13730 , \13613 , \13546 );
nor \U$12869 ( \13731 , \13729 , \13730 );
not \U$12870 ( \13732 , \13731 );
or \U$12871 ( \13733 , \13726 , \13732 );
or \U$12872 ( \13734 , \13731 , \13576 );
nand \U$12873 ( \13735 , \13733 , \13734 );
not \U$12874 ( \13736 , \13735 );
xor \U$12875 ( \13737 , \13503 , \13510 );
xor \U$12876 ( \13738 , \13737 , \13518 );
nor \U$12877 ( \13739 , \13736 , \13738 );
and \U$12878 ( \13740 , \13725 , \13739 );
and \U$12879 ( \13741 , \13717 , \13724 );
or \U$12880 ( \13742 , \13740 , \13741 );
not \U$12881 ( \13743 , \13742 );
xor \U$12882 ( \13744 , \13451 , \13208 );
xor \U$12883 ( \13745 , \13744 , \13459 );
xor \U$12884 ( \13746 , \13628 , \13745 );
xor \U$12885 ( \13747 , \13521 , \13538 );
xor \U$12886 ( \13748 , \13747 , \13615 );
and \U$12887 ( \13749 , \13746 , \13748 );
and \U$12888 ( \13750 , \13628 , \13745 );
or \U$12889 ( \13751 , \13749 , \13750 );
nand \U$12890 ( \13752 , \13743 , \13751 );
not \U$12891 ( \13753 , \13462 );
or \U$12892 ( \13754 , \13442 , \13753 );
or \U$12893 ( \13755 , \13620 , \13627 );
not \U$12894 ( \13756 , \13442 );
or \U$12895 ( \13757 , \13462 , \13756 );
nand \U$12896 ( \13758 , \13754 , \13755 , \13757 );
not \U$12897 ( \13759 , \13618 );
and \U$12898 ( \13760 , \13636 , \13629 );
not \U$12899 ( \13761 , \13636 );
and \U$12900 ( \13762 , \13761 , \13628 );
nor \U$12901 ( \13763 , \13760 , \13762 );
not \U$12902 ( \13764 , \13763 );
or \U$12903 ( \13765 , \13759 , \13764 );
or \U$12904 ( \13766 , \13763 , \13618 );
nand \U$12905 ( \13767 , \13765 , \13766 );
and \U$12906 ( \13768 , \13758 , \13767 );
xnor \U$12907 ( \13769 , \13752 , \13768 );
not \U$12908 ( \13770 , \13769 );
xor \U$12909 ( \13771 , \13638 , \13643 );
xor \U$12910 ( \13772 , \13771 , \13649 );
not \U$12911 ( \13773 , \13772 );
and \U$12912 ( \13774 , \13770 , \13773 );
and \U$12913 ( \13775 , \13769 , \13772 );
nor \U$12914 ( \13776 , \13774 , \13775 );
xor \U$12915 ( \13777 , \13758 , \13767 );
not \U$12916 ( \13778 , \13751 );
not \U$12917 ( \13779 , \13742 );
and \U$12918 ( \13780 , \13778 , \13779 );
and \U$12919 ( \13781 , \13751 , \13742 );
nor \U$12920 ( \13782 , \13780 , \13781 );
xor \U$12921 ( \13783 , \13777 , \13782 );
xor \U$12922 ( \13784 , \13628 , \13745 );
xor \U$12923 ( \13785 , \13784 , \13748 );
not \U$12924 ( \13786 , \13528 );
not \U$12925 ( \13787 , \13537 );
and \U$12926 ( \13788 , \13786 , \13787 );
and \U$12927 ( \13789 , \13528 , \13537 );
nor \U$12928 ( \13790 , \13788 , \13789 );
and \U$12929 ( \13791 , \13607_nR28bb , \12485 );
and \U$12930 ( \13792 , \12512 , \13388_nR2979 );
nand \U$12931 ( \13793 , \13607_nR28bb , \12482 );
or \U$12932 ( \13794 , \12440 , \13388_nR2979 );
nand \U$12933 ( \13795 , \13794 , \12516 );
and \U$12934 ( \13796 , \13793 , \13795 );
nor \U$12935 ( \13797 , \13791 , \13792 , \13796 );
and \U$12936 ( \13798 , RIb558a00_491, \12333 );
and \U$12937 ( \13799 , RIb558eb0_501, \12317 );
and \U$12938 ( \13800 , \12356 , RIb558c58_496);
and \U$12939 ( \13801 , RIb558be0_495, \12358 );
nor \U$12940 ( \13802 , \13800 , \13801 );
and \U$12941 ( \13803 , \12360 , RIb558898_488);
and \U$12942 ( \13804 , RIb558820_487, \12363 );
nor \U$12943 ( \13805 , \13803 , \13804 );
and \U$12944 ( \13806 , \12313 , RIb5587a8_486);
and \U$12945 ( \13807 , RIb558cd0_497, \12351 );
nor \U$12946 ( \13808 , \13806 , \13807 );
and \U$12947 ( \13809 , \12338 , RIb558988_490);
and \U$12948 ( \13810 , RIb558910_489, \12341 );
nor \U$12949 ( \13811 , \13809 , \13810 );
nand \U$12950 ( \13812 , \13802 , \13805 , \13808 , \13811 );
nor \U$12951 ( \13813 , \13798 , \13799 , \13812 );
and \U$12952 ( \13814 , \12309 , RIb558e38_500);
and \U$12953 ( \13815 , RIb558dc0_499, \12320 );
nor \U$12954 ( \13816 , \13814 , \13815 );
nand \U$12955 ( \13817 , RIb558f28_502, \8856 );
and \U$12956 ( \13818 , RIb558af0_493, \12327 );
and \U$12957 ( \13819 , RIb558a78_492, \12330 );
and \U$12958 ( \13820 , \12324 , RIb558b68_494);
and \U$12959 ( \13821 , RIb558d48_498, \12349 );
nor \U$12960 ( \13822 , \13820 , \13821 );
not \U$12961 ( \13823 , \13822 );
nor \U$12962 ( \13824 , \13818 , \13819 , \13823 );
nand \U$12963 ( \13825 , \13813 , \13816 , \13817 , \13824 );
_DC r26a6 ( \13826_nR26a6 , \13825 , \12369 );
nand \U$12964 ( \13827 , \13826_nR26a6 , \12288 );
and \U$12965 ( \13828 , \13797 , \13827 );
and \U$12966 ( \13829 , \13575_nR27ee , \12426 );
and \U$12967 ( \13830 , RIb559180_507, \12338 );
and \U$12968 ( \13831 , RIb5596a8_518, \12317 );
and \U$12969 ( \13832 , \12351 , RIb5594c8_514);
and \U$12970 ( \13833 , RIb559450_513, \12356 );
nor \U$12971 ( \13834 , \13832 , \13833 );
and \U$12972 ( \13835 , \12320 , RIb5595b8_516);
and \U$12973 ( \13836 , RIb559108_506, \12341 );
nor \U$12974 ( \13837 , \13835 , \13836 );
and \U$12975 ( \13838 , \12313 , RIb558fa0_503);
and \U$12976 ( \13839 , RIb559018_504, \12363 );
nor \U$12977 ( \13840 , \13838 , \13839 );
and \U$12978 ( \13841 , \12358 , RIb5593d8_512);
and \U$12979 ( \13842 , RIb559090_505, \12360 );
nor \U$12980 ( \13843 , \13841 , \13842 );
nand \U$12981 ( \13844 , \13834 , \13837 , \13840 , \13843 );
nor \U$12982 ( \13845 , \13830 , \13831 , \13844 );
and \U$12983 ( \13846 , \12309 , RIb559630_517);
and \U$12984 ( \13847 , RIb559540_515, \12349 );
nor \U$12985 ( \13848 , \13846 , \13847 );
nand \U$12986 ( \13849 , RIb559720_519, \8856 );
and \U$12987 ( \13850 , RIb559270_509, \12330 );
and \U$12988 ( \13851 , RIb5591f8_508, \12333 );
and \U$12989 ( \13852 , \12324 , RIb559360_511);
and \U$12990 ( \13853 , RIb5592e8_510, \12327 );
nor \U$12991 ( \13854 , \13852 , \13853 );
not \U$12992 ( \13855 , \13854 );
nor \U$12993 ( \13856 , \13850 , \13851 , \13855 );
nand \U$12994 ( \13857 , \13845 , \13848 , \13849 , \13856 );
_DC r274c ( \13858_nR274c , \13857 , \12369 );
and \U$12995 ( \13859 , \12388 , \13858_nR274c );
nand \U$12996 ( \13860 , \13575_nR27ee , \12381 );
or \U$12997 ( \13861 , \12387 , \13858_nR274c );
nand \U$12998 ( \13862 , \13861 , \12422 );
and \U$12999 ( \13863 , \13860 , \13862 );
nor \U$13000 ( \13864 , \13829 , \13859 , \13863 );
nor \U$13001 ( \13865 , \13828 , \13864 );
not \U$13002 ( \13866 , \13865 );
and \U$13003 ( \13867 , \12952_nR2c3a , \12803 );
or \U$13004 ( \13868 , \12733 , \12843_nR2d1d );
nand \U$13005 ( \13869 , \13868 , \12891 );
nand \U$13006 ( \13870 , \12952_nR2c3a , \12801 );
and \U$13007 ( \13871 , \13869 , \13870 );
and \U$13008 ( \13872 , \12843_nR2d1d , \12895 );
nor \U$13009 ( \13873 , \13867 , \13871 , \13872 );
nand \U$13010 ( \13874 , \12762_nR2e29 , \13018 );
or \U$13011 ( \13875 , \12913 , \12690_nR2f21 );
nand \U$13012 ( \13876 , \13875 , \13187 );
and \U$13013 ( \13877 , \13874 , \13876 );
and \U$13014 ( \13878 , \13190 , \12690_nR2f21 );
and \U$13015 ( \13879 , \12762_nR2e29 , \13021 );
nor \U$13016 ( \13880 , \13877 , \13878 , \13879 );
xor \U$13017 ( \13881 , \13873 , \13880 );
and \U$13018 ( \13882 , \13175_nR2b34 , \12712 );
or \U$13019 ( \13883 , \12562 , \13322_nR2a51 );
nand \U$13020 ( \13884 , \13883 , \12658 );
nand \U$13021 ( \13885 , \13175_nR2b34 , \12651 );
and \U$13022 ( \13886 , \13884 , \13885 );
and \U$13023 ( \13887 , \13322_nR2a51 , \12654 );
nor \U$13024 ( \13888 , \13882 , \13886 , \13887 );
and \U$13025 ( \13889 , \13881 , \13888 );
and \U$13026 ( \13890 , \13873 , \13880 );
or \U$13027 ( \13891 , \13889 , \13890 );
nand \U$13028 ( \13892 , \13866 , \13891 );
or \U$13029 ( \13893 , \13701 , \12371 );
or \U$13030 ( \13894 , \12370_nR3379 , \13536 );
or \U$13031 ( \13895 , \12470_nR3271 , \13535 );
nand \U$13032 ( \13896 , \13893 , \13894 , \13895 );
or \U$13033 ( \13897 , \13252 , \12632 );
or \U$13034 ( \13898 , \13213 , \12549_nR3150 );
nand \U$13035 ( \13899 , \13898 , \13445 );
nand \U$13036 ( \13900 , \12631_nR3038 , \13248 );
and \U$13037 ( \13901 , \13899 , \13900 );
and \U$13038 ( \13902 , \12549_nR3150 , \13448 );
nor \U$13039 ( \13903 , \13901 , \13902 );
nand \U$13040 ( \13904 , \13897 , \13903 );
and \U$13041 ( \13905 , \13896 , \13904 );
and \U$13042 ( \13906 , \13892 , \13905 );
not \U$13043 ( \13907 , \13865 );
nor \U$13044 ( \13908 , \13907 , \13891 );
nor \U$13045 ( \13909 , \13906 , \13908 );
nand \U$13046 ( \13910 , \13790 , \13909 );
xor \U$13047 ( \13911 , \13671 , \13678 );
xor \U$13048 ( \13912 , \13911 , \13686 );
not \U$13049 ( \13913 , \13912 );
nand \U$13050 ( \13914 , \13858_nR274c , \12288 );
and \U$13051 ( \13915 , \13607_nR28bb , \12426 );
and \U$13052 ( \13916 , \12388 , \13575_nR27ee );
nand \U$13053 ( \13917 , \13607_nR28bb , \12381 );
or \U$13054 ( \13918 , \12387 , \13575_nR27ee );
nand \U$13055 ( \13919 , \13918 , \12422 );
and \U$13056 ( \13920 , \13917 , \13919 );
nor \U$13057 ( \13921 , \13915 , \13916 , \13920 );
xor \U$13058 ( \13922 , \13914 , \13921 );
and \U$13059 ( \13923 , \13913 , \13922 );
and \U$13060 ( \13924 , \13910 , \13923 );
nor \U$13061 ( \13925 , \13909 , \13790 );
nor \U$13062 ( \13926 , \13924 , \13925 );
and \U$13063 ( \13927 , \13785 , \13926 );
not \U$13064 ( \13928 , \13927 );
not \U$13065 ( \13929 , \13735 );
not \U$13066 ( \13930 , \13738 );
and \U$13067 ( \13931 , \13929 , \13930 );
and \U$13068 ( \13932 , \13735 , \13738 );
nor \U$13069 ( \13933 , \13931 , \13932 );
not \U$13070 ( \13934 , \13933 );
or \U$13071 ( \13935 , \13921 , \13914 );
not \U$13072 ( \13936 , \13716 );
or \U$13073 ( \13937 , \13936 , \13689 );
not \U$13074 ( \13938 , \13689 );
or \U$13075 ( \13939 , \13716 , \13938 );
nand \U$13076 ( \13940 , \13935 , \13937 , \13939 );
nand \U$13077 ( \13941 , \13934 , \13940 );
not \U$13078 ( \13942 , \13941 );
and \U$13079 ( \13943 , \13928 , \13942 );
nor \U$13080 ( \13944 , \13785 , \13926 );
nor \U$13081 ( \13945 , \13943 , \13944 );
not \U$13082 ( \13946 , \13945 );
and \U$13083 ( \13947 , \13783 , \13946 );
and \U$13084 ( \13948 , \13777 , \13782 );
or \U$13085 ( \13949 , \13947 , \13948 );
xor \U$13086 ( \13950 , \13776 , \13949 );
not \U$13087 ( \13951 , \13940 );
not \U$13088 ( \13952 , \13933 );
or \U$13089 ( \13953 , \13951 , \13952 );
or \U$13090 ( \13954 , \13933 , \13940 );
nand \U$13091 ( \13955 , \13953 , \13954 );
not \U$13092 ( \13956 , \13696 );
xor \U$13093 ( \13957 , \13704 , \13714 );
not \U$13094 ( \13958 , \13957 );
or \U$13095 ( \13959 , \13956 , \13958 );
or \U$13096 ( \13960 , \13957 , \13696 );
nand \U$13097 ( \13961 , \13959 , \13960 );
and \U$13098 ( \13962 , \13322_nR2a51 , \12712 );
or \U$13099 ( \13963 , \12562 , \13388_nR2979 );
nand \U$13100 ( \13964 , \13963 , \12658 );
nand \U$13101 ( \13965 , \13322_nR2a51 , \12651 );
and \U$13102 ( \13966 , \13964 , \13965 );
and \U$13103 ( \13967 , \13388_nR2979 , \12654 );
nor \U$13104 ( \13968 , \13962 , \13966 , \13967 );
and \U$13105 ( \13969 , \13175_nR2b34 , \12803 );
or \U$13106 ( \13970 , \12733 , \12952_nR2c3a );
nand \U$13107 ( \13971 , \13970 , \12891 );
nand \U$13108 ( \13972 , \13175_nR2b34 , \12801 );
and \U$13109 ( \13973 , \13971 , \13972 );
and \U$13110 ( \13974 , \12952_nR2c3a , \12895 );
nor \U$13111 ( \13975 , \13969 , \13973 , \13974 );
xor \U$13112 ( \13976 , \13968 , \13975 );
and \U$13113 ( \13977 , \13575_nR27ee , \12485 );
and \U$13114 ( \13978 , \12512 , \13607_nR28bb );
nand \U$13115 ( \13979 , \13575_nR27ee , \12482 );
or \U$13116 ( \13980 , \12440 , \13607_nR28bb );
nand \U$13117 ( \13981 , \13980 , \12516 );
and \U$13118 ( \13982 , \13979 , \13981 );
nor \U$13119 ( \13983 , \13977 , \13978 , \13982 );
and \U$13120 ( \13984 , \13976 , \13983 );
and \U$13121 ( \13985 , \13968 , \13975 );
or \U$13122 ( \13986 , \13984 , \13985 );
nand \U$13123 ( \13987 , \12690_nR2f21 , \13248 );
or \U$13124 ( \13988 , \13213 , \12631_nR3038 );
nand \U$13125 ( \13989 , \13988 , \13445 );
and \U$13126 ( \13990 , \13987 , \13989 );
and \U$13127 ( \13991 , \13448 , \12631_nR3038 );
and \U$13128 ( \13992 , \12690_nR2f21 , \13251 );
nor \U$13129 ( \13993 , \13990 , \13991 , \13992 );
and \U$13130 ( \13994 , \12492 , \13698 );
not \U$13131 ( \13995 , \12549_nR3150 );
and \U$13132 ( \13996 , \13534 , \13995 );
and \U$13133 ( \13997 , \12470_nR3271 , \13702 );
nor \U$13134 ( \13998 , \13994 , \13996 , \13997 );
xor \U$13135 ( \13999 , \13993 , \13998 );
nand \U$13136 ( \14000 , \12843_nR2d1d , \13018 );
or \U$13137 ( \14001 , \12913 , \12762_nR2e29 );
nand \U$13138 ( \14002 , \14001 , \13187 );
and \U$13139 ( \14003 , \14000 , \14002 );
and \U$13140 ( \14004 , \13190 , \12762_nR2e29 );
and \U$13141 ( \14005 , \12843_nR2d1d , \13021 );
nor \U$13142 ( \14006 , \14003 , \14004 , \14005 );
and \U$13143 ( \14007 , \13999 , \14006 );
and \U$13144 ( \14008 , \13993 , \13998 );
or \U$13145 ( \14009 , \14007 , \14008 );
nor \U$13146 ( \14010 , \13986 , \14009 );
and \U$13147 ( \14011 , \13961 , \14010 );
xor \U$13148 ( \14012 , \13955 , \14011 );
not \U$13149 ( \14013 , \13923 );
not \U$13150 ( \14014 , \13925 );
nand \U$13151 ( \14015 , \14014 , \13910 );
not \U$13152 ( \14016 , \14015 );
or \U$13153 ( \14017 , \14013 , \14016 );
or \U$13154 ( \14018 , \14015 , \13923 );
nand \U$13155 ( \14019 , \14017 , \14018 );
and \U$13156 ( \14020 , \14012 , \14019 );
and \U$13157 ( \14021 , \13955 , \14011 );
or \U$13158 ( \14022 , \14020 , \14021 );
xor \U$13159 ( \14023 , \13717 , \13724 );
xor \U$13160 ( \14024 , \14023 , \13739 );
xor \U$13161 ( \14025 , \14022 , \14024 );
not \U$13162 ( \14026 , \13941 );
nor \U$13163 ( \14027 , \13944 , \13927 );
not \U$13164 ( \14028 , \14027 );
or \U$13165 ( \14029 , \14026 , \14028 );
or \U$13166 ( \14030 , \14027 , \13941 );
nand \U$13167 ( \14031 , \14029 , \14030 );
and \U$13168 ( \14032 , \14025 , \14031 );
and \U$13169 ( \14033 , \14022 , \14024 );
or \U$13170 ( \14034 , \14032 , \14033 );
xor \U$13171 ( \14035 , \13777 , \13782 );
xor \U$13172 ( \14036 , \14035 , \13946 );
xor \U$13173 ( \14037 , \14034 , \14036 );
xor \U$13174 ( \14038 , \14022 , \14024 );
xor \U$13175 ( \14039 , \14038 , \14031 );
not \U$13176 ( \14040 , \14009 );
or \U$13177 ( \14041 , \13986 , \14040 );
and \U$13178 ( \14042 , RIb55a698_552, \12317 );
and \U$13179 ( \14043 , RIb559f90_537, \12313 );
and \U$13180 ( \14044 , \12351 , RIb55a4b8_548);
and \U$13181 ( \14045 , RIb55a440_547, \12356 );
nor \U$13182 ( \14046 , \14044 , \14045 );
and \U$13183 ( \14047 , \12324 , RIb55a350_545);
and \U$13184 ( \14048 , RIb55a2d8_544, \12327 );
nor \U$13185 ( \14049 , \14047 , \14048 );
and \U$13186 ( \14050 , \12330 , RIb55a260_543);
and \U$13187 ( \14051 , RIb55a1e8_542, \12333 );
nor \U$13188 ( \14052 , \14050 , \14051 );
and \U$13189 ( \14053 , \12309 , RIb55a620_551);
and \U$13190 ( \14054 , RIb55a530_549, \12349 );
nor \U$13191 ( \14055 , \14053 , \14054 );
nand \U$13192 ( \14056 , \14046 , \14049 , \14052 , \14055 );
nor \U$13193 ( \14057 , \14042 , \14043 , \14056 );
and \U$13194 ( \14058 , \12320 , RIb55a5a8_550);
and \U$13195 ( \14059 , RIb55a3c8_546, \12358 );
nor \U$13196 ( \14060 , \14058 , \14059 );
and \U$13197 ( \14061 , RIb55a170_541, \12338 );
and \U$13198 ( \14062 , RIb55a0f8_540, \12341 );
and \U$13199 ( \14063 , \12360 , RIb55a080_539);
and \U$13200 ( \14064 , RIb55a008_538, \12363 );
nor \U$13201 ( \14065 , \14063 , \14064 );
not \U$13202 ( \14066 , \14065 );
nor \U$13203 ( \14067 , \14061 , \14062 , \14066 );
nand \U$13204 ( \14068 , \14057 , \14060 , \10540 , \14067 );
_DC r2626 ( \14069_nR2626 , \14068 , \12369 );
nand \U$13205 ( \14070 , \14069_nR2626 , \12288 );
and \U$13206 ( \14071 , \13858_nR274c , \12426 );
and \U$13207 ( \14072 , \12388 , \13826_nR26a6 );
nand \U$13208 ( \14073 , \13858_nR274c , \12381 );
or \U$13209 ( \14074 , \12387 , \13826_nR26a6 );
nand \U$13210 ( \14075 , \14074 , \12422 );
and \U$13211 ( \14076 , \14073 , \14075 );
nor \U$13212 ( \14077 , \14071 , \14072 , \14076 );
or \U$13213 ( \14078 , \14070 , \14077 );
not \U$13214 ( \14079 , \13986 );
or \U$13215 ( \14080 , \14009 , \14079 );
nand \U$13216 ( \14081 , \14041 , \14078 , \14080 );
xor \U$13217 ( \14082 , \13896 , \13904 );
xor \U$13218 ( \14083 , \14081 , \14082 );
not \U$13219 ( \14084 , \13827 );
not \U$13220 ( \14085 , \13864 );
not \U$13221 ( \14086 , \13797 );
and \U$13222 ( \14087 , \14085 , \14086 );
and \U$13223 ( \14088 , \13864 , \13797 );
nor \U$13224 ( \14089 , \14087 , \14088 );
not \U$13225 ( \14090 , \14089 );
or \U$13226 ( \14091 , \14084 , \14090 );
or \U$13227 ( \14092 , \14089 , \13827 );
nand \U$13228 ( \14093 , \14091 , \14092 );
and \U$13229 ( \14094 , \14083 , \14093 );
and \U$13230 ( \14095 , \14081 , \14082 );
or \U$13231 ( \14096 , \14094 , \14095 );
xor \U$13232 ( \14097 , \13913 , \13922 );
xor \U$13233 ( \14098 , \14096 , \14097 );
and \U$13234 ( \14099 , \13322_nR2a51 , \12803 );
or \U$13235 ( \14100 , \12733 , \13175_nR2b34 );
nand \U$13236 ( \14101 , \14100 , \12891 );
nand \U$13237 ( \14102 , \13322_nR2a51 , \12801 );
and \U$13238 ( \14103 , \14101 , \14102 );
and \U$13239 ( \14104 , \13175_nR2b34 , \12895 );
nor \U$13240 ( \14105 , \14099 , \14103 , \14104 );
nand \U$13241 ( \14106 , \12952_nR2c3a , \13018 );
or \U$13242 ( \14107 , \12913 , \12843_nR2d1d );
nand \U$13243 ( \14108 , \14107 , \13187 );
and \U$13244 ( \14109 , \14106 , \14108 );
and \U$13245 ( \14110 , \13190 , \12843_nR2d1d );
and \U$13246 ( \14111 , \12952_nR2c3a , \13021 );
nor \U$13247 ( \14112 , \14109 , \14110 , \14111 );
xor \U$13248 ( \14113 , \14105 , \14112 );
and \U$13249 ( \14114 , \13388_nR2979 , \12712 );
or \U$13250 ( \14115 , \12562 , \13607_nR28bb );
nand \U$13251 ( \14116 , \14115 , \12658 );
nand \U$13252 ( \14117 , \13388_nR2979 , \12651 );
and \U$13253 ( \14118 , \14116 , \14117 );
and \U$13254 ( \14119 , \13607_nR28bb , \12654 );
nor \U$13255 ( \14120 , \14114 , \14118 , \14119 );
and \U$13256 ( \14121 , \14113 , \14120 );
and \U$13257 ( \14122 , \14105 , \14112 );
or \U$13258 ( \14123 , \14121 , \14122 );
nand \U$13259 ( \14124 , \12762_nR2e29 , \13248 );
or \U$13260 ( \14125 , \13213 , \12690_nR2f21 );
nand \U$13261 ( \14126 , \14125 , \13445 );
and \U$13262 ( \14127 , \14124 , \14126 );
and \U$13263 ( \14128 , \13448 , \12690_nR2f21 );
and \U$13264 ( \14129 , \12762_nR2e29 , \13251 );
nor \U$13265 ( \14130 , \14127 , \14128 , \14129 );
not \U$13266 ( \14131 , \14130 );
or \U$13267 ( \14132 , \13701 , \13995 );
or \U$13268 ( \14133 , \12549_nR3150 , \13536 );
or \U$13269 ( \14134 , \12631_nR3038 , \13535 );
nand \U$13270 ( \14135 , \14132 , \14133 , \14134 );
nand \U$13271 ( \14136 , \14131 , \14135 );
xor \U$13272 ( \14137 , \14123 , \14136 );
and \U$13273 ( \14138 , \13858_nR274c , \12485 );
and \U$13274 ( \14139 , \12512 , \13575_nR27ee );
nand \U$13275 ( \14140 , \13858_nR274c , \12482 );
or \U$13276 ( \14141 , \12440 , \13575_nR27ee );
nand \U$13277 ( \14142 , \14141 , \12516 );
and \U$13278 ( \14143 , \14140 , \14142 );
nor \U$13279 ( \14144 , \14138 , \14139 , \14143 );
and \U$13280 ( \14145 , RIb559900_523, \12341 );
and \U$13281 ( \14146 , RIb559ea0_535, \12317 );
and \U$13282 ( \14147 , \12356 , RIb559c48_530);
and \U$13283 ( \14148 , RIb559bd0_529, \12358 );
nor \U$13284 ( \14149 , \14147 , \14148 );
and \U$13285 ( \14150 , \12360 , RIb559888_522);
and \U$13286 ( \14151 , RIb559810_521, \12363 );
nor \U$13287 ( \14152 , \14150 , \14151 );
and \U$13288 ( \14153 , \12309 , RIb559e28_534);
and \U$13289 ( \14154 , RIb559798_520, \12313 );
nor \U$13290 ( \14155 , \14153 , \14154 );
and \U$13291 ( \14156 , \12320 , RIb559db0_533);
and \U$13292 ( \14157 , RIb559cc0_531, \12351 );
nor \U$13293 ( \14158 , \14156 , \14157 );
nand \U$13294 ( \14159 , \14149 , \14152 , \14155 , \14158 );
nor \U$13295 ( \14160 , \14145 , \14146 , \14159 );
and \U$13296 ( \14161 , \12324 , RIb559b58_528);
and \U$13297 ( \14162 , RIb559d38_532, \12349 );
nor \U$13298 ( \14163 , \14161 , \14162 );
and \U$13299 ( \14164 , RIb559978_524, \12338 );
and \U$13300 ( \14165 , RIb5599f0_525, \12333 );
and \U$13301 ( \14166 , \12327 , RIb559ae0_527);
and \U$13302 ( \14167 , RIb559a68_526, \12330 );
nor \U$13303 ( \14168 , \14166 , \14167 );
not \U$13304 ( \14169 , \14168 );
nor \U$13305 ( \14170 , \14164 , \14165 , \14169 );
nand \U$13306 ( \14171 , \14160 , \14163 , \10658 , \14170 );
_DC r25a7 ( \14172_nR25a7 , \14171 , \12369 );
nand \U$13307 ( \14173 , \14172_nR25a7 , \12288 );
and \U$13308 ( \14174 , \14144 , \14173 );
and \U$13309 ( \14175 , \13826_nR26a6 , \12426 );
and \U$13310 ( \14176 , \12388 , \14069_nR2626 );
nand \U$13311 ( \14177 , \13826_nR26a6 , \12381 );
or \U$13312 ( \14178 , \12387 , \14069_nR2626 );
nand \U$13313 ( \14179 , \14178 , \12422 );
and \U$13314 ( \14180 , \14177 , \14179 );
nor \U$13315 ( \14181 , \14175 , \14176 , \14180 );
nor \U$13316 ( \14182 , \14174 , \14181 );
not \U$13317 ( \14183 , \14182 );
and \U$13318 ( \14184 , \14137 , \14183 );
and \U$13319 ( \14185 , \14123 , \14136 );
or \U$13320 ( \14186 , \14184 , \14185 );
xor \U$13321 ( \14187 , \13873 , \13880 );
xor \U$13322 ( \14188 , \14187 , \13888 );
xor \U$13323 ( \14189 , \14186 , \14188 );
xnor \U$13324 ( \14190 , \14070 , \14077 );
xor \U$13325 ( \14191 , \13968 , \13975 );
xor \U$13326 ( \14192 , \14191 , \13983 );
and \U$13327 ( \14193 , \14190 , \14192 );
not \U$13328 ( \14194 , \14193 );
xor \U$13329 ( \14195 , \13993 , \13998 );
xor \U$13330 ( \14196 , \14195 , \14006 );
not \U$13331 ( \14197 , \14196 );
and \U$13332 ( \14198 , \14194 , \14197 );
nor \U$13333 ( \14199 , \14190 , \14192 );
nor \U$13334 ( \14200 , \14198 , \14199 );
and \U$13335 ( \14201 , \14189 , \14200 );
and \U$13336 ( \14202 , \14186 , \14188 );
or \U$13337 ( \14203 , \14201 , \14202 );
not \U$13338 ( \14204 , \14203 );
and \U$13339 ( \14205 , \14098 , \14204 );
and \U$13340 ( \14206 , \14096 , \14097 );
or \U$13341 ( \14207 , \14205 , \14206 );
xor \U$13342 ( \14208 , \13961 , \14010 );
not \U$13343 ( \14209 , \13905 );
not \U$13344 ( \14210 , \13908 );
nand \U$13345 ( \14211 , \14210 , \13892 );
not \U$13346 ( \14212 , \14211 );
or \U$13347 ( \14213 , \14209 , \14212 );
or \U$13348 ( \14214 , \14211 , \13905 );
nand \U$13349 ( \14215 , \14213 , \14214 );
and \U$13350 ( \14216 , \14208 , \14215 );
xor \U$13351 ( \14217 , \14207 , \14216 );
xor \U$13352 ( \14218 , \13955 , \14011 );
xor \U$13353 ( \14219 , \14218 , \14019 );
and \U$13354 ( \14220 , \14217 , \14219 );
and \U$13355 ( \14221 , \14207 , \14216 );
or \U$13356 ( \14222 , \14220 , \14221 );
xor \U$13357 ( \14223 , \14039 , \14222 );
xor \U$13358 ( \14224 , \14186 , \14188 );
xor \U$13359 ( \14225 , \14224 , \14200 );
xor \U$13360 ( \14226 , \14081 , \14082 );
xor \U$13361 ( \14227 , \14226 , \14093 );
not \U$13362 ( \14228 , \14227 );
or \U$13363 ( \14229 , \14225 , \14228 );
not \U$13364 ( \14230 , \14228 );
not \U$13365 ( \14231 , \14225 );
or \U$13366 ( \14232 , \14230 , \14231 );
not \U$13367 ( \14233 , \14173 );
not \U$13368 ( \14234 , \14181 );
not \U$13369 ( \14235 , \14144 );
and \U$13370 ( \14236 , \14234 , \14235 );
and \U$13371 ( \14237 , \14181 , \14144 );
nor \U$13372 ( \14238 , \14236 , \14237 );
not \U$13373 ( \14239 , \14238 );
or \U$13374 ( \14240 , \14233 , \14239 );
or \U$13375 ( \14241 , \14238 , \14173 );
nand \U$13376 ( \14242 , \14240 , \14241 );
not \U$13377 ( \14243 , \14242 );
xor \U$13378 ( \14244 , \14105 , \14112 );
xor \U$13379 ( \14245 , \14244 , \14120 );
nor \U$13380 ( \14246 , \14243 , \14245 );
and \U$13381 ( \14247 , \13607_nR28bb , \12712 );
or \U$13382 ( \14248 , \12562 , \13575_nR27ee );
nand \U$13383 ( \14249 , \14248 , \12658 );
nand \U$13384 ( \14250 , \13607_nR28bb , \12651 );
and \U$13385 ( \14251 , \14249 , \14250 );
and \U$13386 ( \14252 , \13575_nR27ee , \12654 );
nor \U$13387 ( \14253 , \14247 , \14251 , \14252 );
and \U$13388 ( \14254 , \13388_nR2979 , \12803 );
or \U$13389 ( \14255 , \12733 , \13322_nR2a51 );
nand \U$13390 ( \14256 , \14255 , \12891 );
nand \U$13391 ( \14257 , \13388_nR2979 , \12801 );
and \U$13392 ( \14258 , \14256 , \14257 );
and \U$13393 ( \14259 , \13322_nR2a51 , \12895 );
nor \U$13394 ( \14260 , \14254 , \14258 , \14259 );
xor \U$13395 ( \14261 , \14253 , \14260 );
and \U$13396 ( \14262 , \13826_nR26a6 , \12485 );
and \U$13397 ( \14263 , \12512 , \13858_nR274c );
nand \U$13398 ( \14264 , \13826_nR26a6 , \12482 );
or \U$13399 ( \14265 , \12440 , \13858_nR274c );
nand \U$13400 ( \14266 , \14265 , \12516 );
and \U$13401 ( \14267 , \14264 , \14266 );
nor \U$13402 ( \14268 , \14262 , \14263 , \14267 );
and \U$13403 ( \14269 , \14261 , \14268 );
and \U$13404 ( \14270 , \14253 , \14260 );
or \U$13405 ( \14271 , \14269 , \14270 );
nand \U$13406 ( \14272 , \12843_nR2d1d , \13248 );
or \U$13407 ( \14273 , \13213 , \12762_nR2e29 );
nand \U$13408 ( \14274 , \14273 , \13445 );
and \U$13409 ( \14275 , \14272 , \14274 );
and \U$13410 ( \14276 , \13448 , \12762_nR2e29 );
and \U$13411 ( \14277 , \12843_nR2d1d , \13251 );
nor \U$13412 ( \14278 , \14275 , \14276 , \14277 );
and \U$13413 ( \14279 , \12632 , \13698 );
not \U$13414 ( \14280 , \12690_nR2f21 );
and \U$13415 ( \14281 , \13534 , \14280 );
and \U$13416 ( \14282 , \12631_nR3038 , \13702 );
nor \U$13417 ( \14283 , \14279 , \14281 , \14282 );
xor \U$13418 ( \14284 , \14278 , \14283 );
nand \U$13419 ( \14285 , \13175_nR2b34 , \13018 );
or \U$13420 ( \14286 , \12913 , \12952_nR2c3a );
nand \U$13421 ( \14287 , \14286 , \13187 );
and \U$13422 ( \14288 , \14285 , \14287 );
and \U$13423 ( \14289 , \13190 , \12952_nR2c3a );
and \U$13424 ( \14290 , \13175_nR2b34 , \13021 );
nor \U$13425 ( \14291 , \14288 , \14289 , \14290 );
and \U$13426 ( \14292 , \14284 , \14291 );
and \U$13427 ( \14293 , \14278 , \14283 );
or \U$13428 ( \14294 , \14292 , \14293 );
nor \U$13429 ( \14295 , \14271 , \14294 );
xor \U$13430 ( \14296 , \14246 , \14295 );
not \U$13431 ( \14297 , \14196 );
nor \U$13432 ( \14298 , \14199 , \14193 );
not \U$13433 ( \14299 , \14298 );
or \U$13434 ( \14300 , \14297 , \14299 );
or \U$13435 ( \14301 , \14298 , \14196 );
nand \U$13436 ( \14302 , \14300 , \14301 );
and \U$13437 ( \14303 , \14296 , \14302 );
and \U$13438 ( \14304 , \14246 , \14295 );
or \U$13439 ( \14305 , \14303 , \14304 );
nand \U$13440 ( \14306 , \14232 , \14305 );
nand \U$13441 ( \14307 , \14229 , \14306 );
xor \U$13442 ( \14308 , \14208 , \14215 );
xor \U$13443 ( \14309 , \14307 , \14308 );
xor \U$13444 ( \14310 , \14096 , \14097 );
xor \U$13445 ( \14311 , \14310 , \14204 );
and \U$13446 ( \14312 , \14309 , \14311 );
and \U$13447 ( \14313 , \14307 , \14308 );
or \U$13448 ( \14314 , \14312 , \14313 );
xor \U$13449 ( \14315 , \14207 , \14216 );
xor \U$13450 ( \14316 , \14315 , \14219 );
xor \U$13451 ( \14317 , \14314 , \14316 );
xor \U$13452 ( \14318 , \14307 , \14308 );
xor \U$13453 ( \14319 , \14318 , \14311 );
not \U$13454 ( \14320 , \14225 );
not \U$13455 ( \14321 , \14305 );
and \U$13456 ( \14322 , \14320 , \14321 );
and \U$13457 ( \14323 , \14225 , \14305 );
nor \U$13458 ( \14324 , \14322 , \14323 );
not \U$13459 ( \14325 , \14324 );
not \U$13460 ( \14326 , \14227 );
and \U$13461 ( \14327 , \14325 , \14326 );
and \U$13462 ( \14328 , \14324 , \14227 );
nor \U$13463 ( \14329 , \14327 , \14328 );
and \U$13464 ( \14330 , RIb55aa58_560, \12330 );
and \U$13465 ( \14331 , RIb55ae90_569, \12317 );
and \U$13466 ( \14332 , \12356 , RIb55ac38_564);
and \U$13467 ( \14333 , RIb55abc0_563, \12358 );
nor \U$13468 ( \14334 , \14332 , \14333 );
and \U$13469 ( \14335 , \12360 , RIb55a878_556);
and \U$13470 ( \14336 , RIb55a800_555, \12363 );
nor \U$13471 ( \14337 , \14335 , \14336 );
and \U$13472 ( \14338 , \12313 , RIb55a788_554);
and \U$13473 ( \14339 , RIb55a8f0_557, \12341 );
nor \U$13474 ( \14340 , \14338 , \14339 );
and \U$13475 ( \14341 , \12338 , RIb55a968_558);
and \U$13476 ( \14342 , RIb55a9e0_559, \12333 );
nor \U$13477 ( \14343 , \14341 , \14342 );
nand \U$13478 ( \14344 , \14334 , \14337 , \14340 , \14343 );
nor \U$13479 ( \14345 , \14330 , \14331 , \14344 );
and \U$13480 ( \14346 , \12309 , RIb55ae18_568);
and \U$13481 ( \14347 , RIb55ada0_567, \12320 );
nor \U$13482 ( \14348 , \14346 , \14347 );
nand \U$13483 ( \14349 , RIb55af08_570, \8856 );
and \U$13484 ( \14350 , RIb55ab48_562, \12324 );
and \U$13485 ( \14351 , RIb55aad0_561, \12327 );
and \U$13486 ( \14352 , \12349 , RIb55ad28_566);
and \U$13487 ( \14353 , RIb55acb0_565, \12351 );
nor \U$13488 ( \14354 , \14352 , \14353 );
not \U$13489 ( \14355 , \14354 );
nor \U$13490 ( \14356 , \14350 , \14351 , \14355 );
nand \U$13491 ( \14357 , \14345 , \14348 , \14349 , \14356 );
_DC r2538 ( \14358_nR2538 , \14357 , \12369 );
nand \U$13492 ( \14359 , \14358_nR2538 , \12288 );
and \U$13493 ( \14360 , \14069_nR2626 , \12426 );
and \U$13494 ( \14361 , \12388 , \14172_nR25a7 );
nand \U$13495 ( \14362 , \14069_nR2626 , \12381 );
or \U$13496 ( \14363 , \12387 , \14172_nR25a7 );
nand \U$13497 ( \14364 , \14363 , \12422 );
and \U$13498 ( \14365 , \14362 , \14364 );
nor \U$13499 ( \14366 , \14360 , \14361 , \14365 );
xnor \U$13500 ( \14367 , \14359 , \14366 );
xor \U$13501 ( \14368 , \14253 , \14260 );
xor \U$13502 ( \14369 , \14368 , \14268 );
and \U$13503 ( \14370 , \14367 , \14369 );
not \U$13504 ( \14371 , \14370 );
xor \U$13505 ( \14372 , \14278 , \14283 );
xor \U$13506 ( \14373 , \14372 , \14291 );
not \U$13507 ( \14374 , \14373 );
and \U$13508 ( \14375 , \14371 , \14374 );
nor \U$13509 ( \14376 , \14367 , \14369 );
nor \U$13510 ( \14377 , \14375 , \14376 );
and \U$13511 ( \14378 , \14069_nR2626 , \12485 );
and \U$13512 ( \14379 , \12512 , \13826_nR26a6 );
nand \U$13513 ( \14380 , \14069_nR2626 , \12482 );
or \U$13514 ( \14381 , \12440 , \13826_nR26a6 );
nand \U$13515 ( \14382 , \14381 , \12516 );
and \U$13516 ( \14383 , \14380 , \14382 );
nor \U$13517 ( \14384 , \14378 , \14379 , \14383 );
and \U$13518 ( \14385 , RIb55b4a8_582, \12351 );
and \U$13519 ( \14386 , RIb55af80_571, \12313 );
and \U$13520 ( \14387 , \12349 , RIb55b520_583);
and \U$13521 ( \14388 , RIb55b598_584, \12320 );
nor \U$13522 ( \14389 , \14387 , \14388 );
and \U$13523 ( \14390 , \12324 , RIb55b340_579);
and \U$13524 ( \14391 , RIb55b2c8_578, \12327 );
nor \U$13525 ( \14392 , \14390 , \14391 );
and \U$13526 ( \14393 , \12330 , RIb55b250_577);
and \U$13527 ( \14394 , RIb55b1d8_576, \12333 );
nor \U$13528 ( \14395 , \14393 , \14394 );
and \U$13529 ( \14396 , \12317 , RIb55b688_586);
and \U$13530 ( \14397 , RIb55b610_585, \12309 );
nor \U$13531 ( \14398 , \14396 , \14397 );
nand \U$13532 ( \14399 , \14389 , \14392 , \14395 , \14398 );
nor \U$13533 ( \14400 , \14385 , \14386 , \14399 );
and \U$13534 ( \14401 , \12356 , RIb55b430_581);
and \U$13535 ( \14402 , RIb55b3b8_580, \12358 );
nor \U$13536 ( \14403 , \14401 , \14402 );
nand \U$13537 ( \14404 , RIb55b700_587, \8856 );
and \U$13538 ( \14405 , RIb55b160_575, \12338 );
and \U$13539 ( \14406 , RIb55b0e8_574, \12341 );
and \U$13540 ( \14407 , \12360 , RIb55b070_573);
and \U$13541 ( \14408 , RIb55aff8_572, \12363 );
nor \U$13542 ( \14409 , \14407 , \14408 );
not \U$13543 ( \14410 , \14409 );
nor \U$13544 ( \14411 , \14405 , \14406 , \14410 );
nand \U$13545 ( \14412 , \14400 , \14403 , \14404 , \14411 );
_DC r2430 ( \14413_nR2430 , \14412 , \12369 );
nand \U$13546 ( \14414 , \14413_nR2430 , \12288 );
and \U$13547 ( \14415 , \14384 , \14414 );
and \U$13548 ( \14416 , \14172_nR25a7 , \12426 );
and \U$13549 ( \14417 , \12388 , \14358_nR2538 );
nand \U$13550 ( \14418 , \14172_nR25a7 , \12381 );
or \U$13551 ( \14419 , \12387 , \14358_nR2538 );
nand \U$13552 ( \14420 , \14419 , \12422 );
and \U$13553 ( \14421 , \14418 , \14420 );
nor \U$13554 ( \14422 , \14416 , \14417 , \14421 );
nor \U$13555 ( \14423 , \14415 , \14422 );
not \U$13556 ( \14424 , \14423 );
and \U$13557 ( \14425 , \13607_nR28bb , \12803 );
or \U$13558 ( \14426 , \12733 , \13388_nR2979 );
nand \U$13559 ( \14427 , \14426 , \12891 );
nand \U$13560 ( \14428 , \13607_nR28bb , \12801 );
and \U$13561 ( \14429 , \14427 , \14428 );
and \U$13562 ( \14430 , \13388_nR2979 , \12895 );
nor \U$13563 ( \14431 , \14425 , \14429 , \14430 );
nand \U$13564 ( \14432 , \13322_nR2a51 , \13018 );
or \U$13565 ( \14433 , \12913 , \13175_nR2b34 );
nand \U$13566 ( \14434 , \14433 , \13187 );
and \U$13567 ( \14435 , \14432 , \14434 );
and \U$13568 ( \14436 , \13190 , \13175_nR2b34 );
and \U$13569 ( \14437 , \13322_nR2a51 , \13021 );
nor \U$13570 ( \14438 , \14435 , \14436 , \14437 );
xor \U$13571 ( \14439 , \14431 , \14438 );
and \U$13572 ( \14440 , \13575_nR27ee , \12712 );
or \U$13573 ( \14441 , \12562 , \13858_nR274c );
nand \U$13574 ( \14442 , \14441 , \12658 );
nand \U$13575 ( \14443 , \13575_nR27ee , \12651 );
and \U$13576 ( \14444 , \14442 , \14443 );
and \U$13577 ( \14445 , \13858_nR274c , \12654 );
nor \U$13578 ( \14446 , \14440 , \14444 , \14445 );
and \U$13579 ( \14447 , \14439 , \14446 );
and \U$13580 ( \14448 , \14431 , \14438 );
or \U$13581 ( \14449 , \14447 , \14448 );
nand \U$13582 ( \14450 , \14424 , \14449 );
or \U$13583 ( \14451 , \13701 , \14280 );
or \U$13584 ( \14452 , \12690_nR2f21 , \13536 );
or \U$13585 ( \14453 , \12762_nR2e29 , \13535 );
nand \U$13586 ( \14454 , \14451 , \14452 , \14453 );
not \U$13587 ( \14455 , \12952_nR2c3a );
or \U$13588 ( \14456 , \13252 , \14455 );
or \U$13589 ( \14457 , \13213 , \12843_nR2d1d );
nand \U$13590 ( \14458 , \14457 , \13445 );
nand \U$13591 ( \14459 , \12952_nR2c3a , \13248 );
and \U$13592 ( \14460 , \14458 , \14459 );
and \U$13593 ( \14461 , \12843_nR2d1d , \13448 );
nor \U$13594 ( \14462 , \14460 , \14461 );
nand \U$13595 ( \14463 , \14456 , \14462 );
and \U$13596 ( \14464 , \14454 , \14463 );
and \U$13597 ( \14465 , \14450 , \14464 );
not \U$13598 ( \14466 , \14423 );
nor \U$13599 ( \14467 , \14466 , \14449 );
nor \U$13600 ( \14468 , \14465 , \14467 );
and \U$13601 ( \14469 , \14377 , \14468 );
not \U$13602 ( \14470 , \14469 );
not \U$13603 ( \14471 , \14130 );
not \U$13604 ( \14472 , \14135 );
and \U$13605 ( \14473 , \14471 , \14472 );
and \U$13606 ( \14474 , \14130 , \14135 );
nor \U$13607 ( \14475 , \14473 , \14474 );
not \U$13608 ( \14476 , \14475 );
and \U$13609 ( \14477 , \14470 , \14476 );
nor \U$13610 ( \14478 , \14377 , \14468 );
nor \U$13611 ( \14479 , \14477 , \14478 );
xor \U$13612 ( \14480 , \14123 , \14136 );
xor \U$13613 ( \14481 , \14480 , \14183 );
and \U$13614 ( \14482 , \14479 , \14481 );
not \U$13615 ( \14483 , \14482 );
not \U$13616 ( \14484 , \14242 );
not \U$13617 ( \14485 , \14245 );
and \U$13618 ( \14486 , \14484 , \14485 );
and \U$13619 ( \14487 , \14242 , \14245 );
nor \U$13620 ( \14488 , \14486 , \14487 );
not \U$13621 ( \14489 , \14488 );
or \U$13622 ( \14490 , \14366 , \14359 );
not \U$13623 ( \14491 , \14294 );
or \U$13624 ( \14492 , \14491 , \14271 );
not \U$13625 ( \14493 , \14271 );
or \U$13626 ( \14494 , \14294 , \14493 );
nand \U$13627 ( \14495 , \14490 , \14492 , \14494 );
nand \U$13628 ( \14496 , \14489 , \14495 );
not \U$13629 ( \14497 , \14496 );
and \U$13630 ( \14498 , \14483 , \14497 );
nor \U$13631 ( \14499 , \14479 , \14481 );
nor \U$13632 ( \14500 , \14498 , \14499 );
nor \U$13633 ( \14501 , \14329 , \14500 );
xor \U$13634 ( \14502 , \14319 , \14501 );
and \U$13635 ( \14503 , \14329 , \14500 );
nor \U$13636 ( \14504 , \14503 , \14501 );
xor \U$13637 ( \14505 , \14246 , \14295 );
xor \U$13638 ( \14506 , \14505 , \14302 );
not \U$13639 ( \14507 , \14496 );
nor \U$13640 ( \14508 , \14499 , \14482 );
not \U$13641 ( \14509 , \14508 );
or \U$13642 ( \14510 , \14507 , \14509 );
or \U$13643 ( \14511 , \14508 , \14496 );
nand \U$13644 ( \14512 , \14510 , \14511 );
and \U$13645 ( \14513 , \14506 , \14512 );
xor \U$13646 ( \14514 , \14504 , \14513 );
xor \U$13647 ( \14515 , \14506 , \14512 );
and \U$13648 ( \14516 , \13858_nR274c , \12712 );
or \U$13649 ( \14517 , \12562 , \13826_nR26a6 );
nand \U$13650 ( \14518 , \14517 , \12658 );
nand \U$13651 ( \14519 , \13858_nR274c , \12651 );
and \U$13652 ( \14520 , \14518 , \14519 );
and \U$13653 ( \14521 , \13826_nR26a6 , \12654 );
nor \U$13654 ( \14522 , \14516 , \14520 , \14521 );
and \U$13655 ( \14523 , \13575_nR27ee , \12803 );
or \U$13656 ( \14524 , \12733 , \13607_nR28bb );
nand \U$13657 ( \14525 , \14524 , \12891 );
nand \U$13658 ( \14526 , \13575_nR27ee , \12801 );
and \U$13659 ( \14527 , \14525 , \14526 );
and \U$13660 ( \14528 , \13607_nR28bb , \12895 );
nor \U$13661 ( \14529 , \14523 , \14527 , \14528 );
xor \U$13662 ( \14530 , \14522 , \14529 );
and \U$13663 ( \14531 , \14172_nR25a7 , \12485 );
and \U$13664 ( \14532 , \12512 , \14069_nR2626 );
nand \U$13665 ( \14533 , \14172_nR25a7 , \12482 );
or \U$13666 ( \14534 , \12440 , \14069_nR2626 );
nand \U$13667 ( \14535 , \14534 , \12516 );
and \U$13668 ( \14536 , \14533 , \14535 );
nor \U$13669 ( \14537 , \14531 , \14532 , \14536 );
and \U$13670 ( \14538 , \14530 , \14537 );
and \U$13671 ( \14539 , \14522 , \14529 );
or \U$13672 ( \14540 , \14538 , \14539 );
nand \U$13673 ( \14541 , \13175_nR2b34 , \13248 );
or \U$13674 ( \14542 , \13213 , \12952_nR2c3a );
nand \U$13675 ( \14543 , \14542 , \13445 );
and \U$13676 ( \14544 , \14541 , \14543 );
and \U$13677 ( \14545 , \13448 , \12952_nR2c3a );
and \U$13678 ( \14546 , \13175_nR2b34 , \13251 );
nor \U$13679 ( \14547 , \14544 , \14545 , \14546 );
and \U$13680 ( \14548 , \12763 , \13698 );
not \U$13681 ( \14549 , \12843_nR2d1d );
and \U$13682 ( \14550 , \13534 , \14549 );
and \U$13683 ( \14551 , \12762_nR2e29 , \13702 );
nor \U$13684 ( \14552 , \14548 , \14550 , \14551 );
xor \U$13685 ( \14553 , \14547 , \14552 );
nand \U$13686 ( \14554 , \13388_nR2979 , \13018 );
or \U$13687 ( \14555 , \12913 , \13322_nR2a51 );
nand \U$13688 ( \14556 , \14555 , \13187 );
and \U$13689 ( \14557 , \14554 , \14556 );
and \U$13690 ( \14558 , \13190 , \13322_nR2a51 );
and \U$13691 ( \14559 , \13388_nR2979 , \13021 );
nor \U$13692 ( \14560 , \14557 , \14558 , \14559 );
and \U$13693 ( \14561 , \14553 , \14560 );
and \U$13694 ( \14562 , \14547 , \14552 );
or \U$13695 ( \14563 , \14561 , \14562 );
xor \U$13696 ( \14564 , \14540 , \14563 );
not \U$13697 ( \14565 , \14422 );
not \U$13698 ( \14566 , \14384 );
and \U$13699 ( \14567 , \14565 , \14566 );
and \U$13700 ( \14568 , \14422 , \14384 );
nor \U$13701 ( \14569 , \14567 , \14568 );
not \U$13702 ( \14570 , \14569 );
not \U$13703 ( \14571 , \14414 );
and \U$13704 ( \14572 , \14570 , \14571 );
and \U$13705 ( \14573 , \14569 , \14414 );
nor \U$13706 ( \14574 , \14572 , \14573 );
and \U$13707 ( \14575 , \14564 , \14574 );
and \U$13708 ( \14576 , \14540 , \14563 );
or \U$13709 ( \14577 , \14575 , \14576 );
not \U$13710 ( \14578 , \14577 );
xor \U$13711 ( \14579 , \14454 , \14463 );
not \U$13712 ( \14580 , \14579 );
xor \U$13713 ( \14581 , \14431 , \14438 );
xor \U$13714 ( \14582 , \14581 , \14446 );
nor \U$13715 ( \14583 , \14580 , \14582 );
xor \U$13716 ( \14584 , \14578 , \14583 );
not \U$13717 ( \14585 , \14373 );
nor \U$13718 ( \14586 , \14376 , \14370 );
not \U$13719 ( \14587 , \14586 );
or \U$13720 ( \14588 , \14585 , \14587 );
or \U$13721 ( \14589 , \14586 , \14373 );
nand \U$13722 ( \14590 , \14588 , \14589 );
and \U$13723 ( \14591 , \14584 , \14590 );
and \U$13724 ( \14592 , \14578 , \14583 );
or \U$13725 ( \14593 , \14591 , \14592 );
not \U$13726 ( \14594 , \14495 );
not \U$13727 ( \14595 , \14488 );
or \U$13728 ( \14596 , \14594 , \14595 );
or \U$13729 ( \14597 , \14488 , \14495 );
nand \U$13730 ( \14598 , \14596 , \14597 );
xor \U$13731 ( \14599 , \14593 , \14598 );
not \U$13732 ( \14600 , \14475 );
nor \U$13733 ( \14601 , \14478 , \14469 );
not \U$13734 ( \14602 , \14601 );
or \U$13735 ( \14603 , \14600 , \14602 );
or \U$13736 ( \14604 , \14601 , \14475 );
nand \U$13737 ( \14605 , \14603 , \14604 );
and \U$13738 ( \14606 , \14599 , \14605 );
and \U$13739 ( \14607 , \14593 , \14598 );
or \U$13740 ( \14608 , \14606 , \14607 );
xor \U$13741 ( \14609 , \14515 , \14608 );
xor \U$13742 ( \14610 , \14578 , \14583 );
xor \U$13743 ( \14611 , \14610 , \14590 );
not \U$13744 ( \14612 , \14464 );
not \U$13745 ( \14613 , \14467 );
nand \U$13746 ( \14614 , \14613 , \14450 );
not \U$13747 ( \14615 , \14614 );
or \U$13748 ( \14616 , \14612 , \14615 );
or \U$13749 ( \14617 , \14614 , \14464 );
nand \U$13750 ( \14618 , \14616 , \14617 );
nor \U$13751 ( \14619 , \14611 , \14618 );
nand \U$13752 ( \14620 , \13322_nR2a51 , \13248 );
or \U$13753 ( \14621 , \13213 , \13175_nR2b34 );
nand \U$13754 ( \14622 , \14621 , \13445 );
and \U$13755 ( \14623 , \14620 , \14622 );
and \U$13756 ( \14624 , \13448 , \13175_nR2b34 );
and \U$13757 ( \14625 , \13322_nR2a51 , \13251 );
nor \U$13758 ( \14626 , \14623 , \14624 , \14625 );
and \U$13759 ( \14627 , \14549 , \13698 );
and \U$13760 ( \14628 , \13534 , \14455 );
and \U$13761 ( \14629 , \12843_nR2d1d , \13702 );
nor \U$13762 ( \14630 , \14627 , \14628 , \14629 );
xor \U$13763 ( \14631 , \14626 , \14630 );
and \U$13764 ( \14632 , \14631 , \12387 );
and \U$13765 ( \14633 , \14626 , \14630 );
or \U$13766 ( \14634 , \14632 , \14633 );
and \U$13767 ( \14635 , \13858_nR274c , \12803 );
or \U$13768 ( \14636 , \12733 , \13575_nR27ee );
nand \U$13769 ( \14637 , \14636 , \12891 );
nand \U$13770 ( \14638 , \13858_nR274c , \12801 );
and \U$13771 ( \14639 , \14637 , \14638 );
and \U$13772 ( \14640 , \13575_nR27ee , \12895 );
nor \U$13773 ( \14641 , \14635 , \14639 , \14640 );
nand \U$13774 ( \14642 , \13607_nR28bb , \13018 );
or \U$13775 ( \14643 , \12913 , \13388_nR2979 );
nand \U$13776 ( \14644 , \14643 , \13187 );
and \U$13777 ( \14645 , \14642 , \14644 );
and \U$13778 ( \14646 , \13190 , \13388_nR2979 );
and \U$13779 ( \14647 , \13607_nR28bb , \13021 );
nor \U$13780 ( \14648 , \14645 , \14646 , \14647 );
xor \U$13781 ( \14649 , \14641 , \14648 );
and \U$13782 ( \14650 , \13826_nR26a6 , \12712 );
or \U$13783 ( \14651 , \12562 , \14069_nR2626 );
nand \U$13784 ( \14652 , \14651 , \12658 );
nand \U$13785 ( \14653 , \13826_nR26a6 , \12651 );
and \U$13786 ( \14654 , \14652 , \14653 );
and \U$13787 ( \14655 , \14069_nR2626 , \12654 );
nor \U$13788 ( \14656 , \14650 , \14654 , \14655 );
and \U$13789 ( \14657 , \14649 , \14656 );
and \U$13790 ( \14658 , \14641 , \14648 );
or \U$13791 ( \14659 , \14657 , \14658 );
xor \U$13792 ( \14660 , \14634 , \14659 );
and \U$13793 ( \14661 , \14358_nR2538 , \12426 );
and \U$13794 ( \14662 , \12388 , \14413_nR2430 );
nand \U$13795 ( \14663 , \14358_nR2538 , \12381 );
or \U$13796 ( \14664 , \12387 , \14413_nR2430 );
nand \U$13797 ( \14665 , \14664 , \12422 );
and \U$13798 ( \14666 , \14663 , \14665 );
nor \U$13799 ( \14667 , \14661 , \14662 , \14666 );
and \U$13800 ( \14668 , \14660 , \14667 );
and \U$13801 ( \14669 , \14634 , \14659 );
or \U$13802 ( \14670 , \14668 , \14669 );
not \U$13803 ( \14671 , \14582 );
not \U$13804 ( \14672 , \14579 );
and \U$13805 ( \14673 , \14671 , \14672 );
and \U$13806 ( \14674 , \14582 , \14579 );
nor \U$13807 ( \14675 , \14673 , \14674 );
xor \U$13808 ( \14676 , \14670 , \14675 );
xor \U$13809 ( \14677 , \14540 , \14563 );
xor \U$13810 ( \14678 , \14677 , \14574 );
and \U$13811 ( \14679 , \14676 , \14678 );
and \U$13812 ( \14680 , \14670 , \14675 );
or \U$13813 ( \14681 , \14679 , \14680 );
or \U$13814 ( \14682 , \14619 , \14681 );
nand \U$13815 ( \14683 , \14618 , \14611 );
nand \U$13816 ( \14684 , \14682 , \14683 );
xor \U$13817 ( \14685 , \14593 , \14598 );
xor \U$13818 ( \14686 , \14685 , \14605 );
xor \U$13819 ( \14687 , \14684 , \14686 );
not \U$13820 ( \14688 , \14681 );
not \U$13821 ( \14689 , \14619 );
nand \U$13822 ( \14690 , \14689 , \14683 );
not \U$13823 ( \14691 , \14690 );
or \U$13824 ( \14692 , \14688 , \14691 );
or \U$13825 ( \14693 , \14690 , \14681 );
nand \U$13826 ( \14694 , \14692 , \14693 );
xor \U$13827 ( \14695 , \14634 , \14659 );
xor \U$13828 ( \14696 , \14695 , \14667 );
xor \U$13829 ( \14697 , \14547 , \14552 );
xor \U$13830 ( \14698 , \14697 , \14560 );
or \U$13831 ( \14699 , \14696 , \14698 );
and \U$13832 ( \14700 , \14358_nR2538 , \12485 );
and \U$13833 ( \14701 , \12512 , \14172_nR25a7 );
nand \U$13834 ( \14702 , \14358_nR2538 , \12482 );
or \U$13835 ( \14703 , \12440 , \14172_nR25a7 );
nand \U$13836 ( \14704 , \14703 , \12516 );
and \U$13837 ( \14705 , \14702 , \14704 );
nor \U$13838 ( \14706 , \14700 , \14701 , \14705 );
nand \U$13839 ( \14707 , \13388_nR2979 , \13248 );
or \U$13840 ( \14708 , \13213 , \13322_nR2a51 );
nand \U$13841 ( \14709 , \14708 , \13445 );
and \U$13842 ( \14710 , \14707 , \14709 );
and \U$13843 ( \14711 , \13448 , \13322_nR2a51 );
and \U$13844 ( \14712 , \13388_nR2979 , \13251 );
nor \U$13845 ( \14713 , \14710 , \14711 , \14712 );
and \U$13846 ( \14714 , \14455 , \13698 );
and \U$13847 ( \14715 , \13534 , \13416 );
and \U$13848 ( \14716 , \12952_nR2c3a , \13702 );
nor \U$13849 ( \14717 , \14714 , \14715 , \14716 );
xor \U$13850 ( \14718 , \14713 , \14717 );
nand \U$13851 ( \14719 , \13575_nR27ee , \13018 );
or \U$13852 ( \14720 , \12913 , \13607_nR28bb );
nand \U$13853 ( \14721 , \14720 , \13187 );
and \U$13854 ( \14722 , \14719 , \14721 );
and \U$13855 ( \14723 , \13190 , \13607_nR28bb );
and \U$13856 ( \14724 , \13575_nR27ee , \13021 );
nor \U$13857 ( \14725 , \14722 , \14723 , \14724 );
and \U$13858 ( \14726 , \14718 , \14725 );
and \U$13859 ( \14727 , \14713 , \14717 );
or \U$13860 ( \14728 , \14726 , \14727 );
xor \U$13861 ( \14729 , \14706 , \14728 );
and \U$13862 ( \14730 , \14069_nR2626 , \12712 );
or \U$13863 ( \14731 , \12562 , \14172_nR25a7 );
nand \U$13864 ( \14732 , \14731 , \12658 );
nand \U$13865 ( \14733 , \14069_nR2626 , \12651 );
and \U$13866 ( \14734 , \14732 , \14733 );
and \U$13867 ( \14735 , \14172_nR25a7 , \12654 );
nor \U$13868 ( \14736 , \14730 , \14734 , \14735 );
and \U$13869 ( \14737 , \13826_nR26a6 , \12803 );
or \U$13870 ( \14738 , \12733 , \13858_nR274c );
nand \U$13871 ( \14739 , \14738 , \12891 );
nand \U$13872 ( \14740 , \13826_nR26a6 , \12801 );
and \U$13873 ( \14741 , \14739 , \14740 );
and \U$13874 ( \14742 , \13858_nR274c , \12895 );
nor \U$13875 ( \14743 , \14737 , \14741 , \14742 );
xor \U$13876 ( \14744 , \14736 , \14743 );
and \U$13877 ( \14745 , \14413_nR2430 , \12485 );
and \U$13878 ( \14746 , \12512 , \14358_nR2538 );
nand \U$13879 ( \14747 , \14413_nR2430 , \12482 );
or \U$13880 ( \14748 , \12440 , \14358_nR2538 );
nand \U$13881 ( \14749 , \14748 , \12516 );
and \U$13882 ( \14750 , \14747 , \14749 );
nor \U$13883 ( \14751 , \14745 , \14746 , \14750 );
and \U$13884 ( \14752 , \14744 , \14751 );
and \U$13885 ( \14753 , \14736 , \14743 );
or \U$13886 ( \14754 , \14752 , \14753 );
and \U$13887 ( \14755 , \14729 , \14754 );
and \U$13888 ( \14756 , \14706 , \14728 );
or \U$13889 ( \14757 , \14755 , \14756 );
xor \U$13890 ( \14758 , \14522 , \14529 );
xor \U$13891 ( \14759 , \14758 , \14537 );
xor \U$13892 ( \14760 , \14757 , \14759 );
xor \U$13893 ( \14761 , \14641 , \14648 );
xor \U$13894 ( \14762 , \14761 , \14656 );
xor \U$13895 ( \14763 , \14626 , \14630 );
xor \U$13896 ( \14764 , \14763 , \12387 );
and \U$13897 ( \14765 , \14762 , \14764 );
and \U$13898 ( \14766 , \12426 , \14413_nR2430 );
nand \U$13899 ( \14767 , \14413_nR2430 , \12381 );
and \U$13900 ( \14768 , \14767 , \12386 );
nor \U$13901 ( \14769 , \14766 , \14768 );
xor \U$13902 ( \14770 , \14626 , \14630 );
xor \U$13903 ( \14771 , \14770 , \12387 );
and \U$13904 ( \14772 , \14769 , \14771 );
and \U$13905 ( \14773 , \14762 , \14769 );
or \U$13906 ( \14774 , \14765 , \14772 , \14773 );
and \U$13907 ( \14775 , \14760 , \14774 );
and \U$13908 ( \14776 , \14757 , \14759 );
or \U$13909 ( \14777 , \14775 , \14776 );
xor \U$13910 ( \14778 , \14699 , \14777 );
xor \U$13911 ( \14779 , \14670 , \14675 );
xor \U$13912 ( \14780 , \14779 , \14678 );
and \U$13913 ( \14781 , \14778 , \14780 );
and \U$13914 ( \14782 , \14699 , \14777 );
or \U$13915 ( \14783 , \14781 , \14782 );
xor \U$13916 ( \14784 , \14694 , \14783 );
nand \U$13917 ( \14785 , \13607_nR28bb , \13248 );
or \U$13918 ( \14786 , \13213 , \13388_nR2979 );
nand \U$13919 ( \14787 , \14786 , \13445 );
and \U$13920 ( \14788 , \14785 , \14787 );
and \U$13921 ( \14789 , \13448 , \13388_nR2979 );
and \U$13922 ( \14790 , \13607_nR28bb , \13251 );
nor \U$13923 ( \14791 , \14788 , \14789 , \14790 );
and \U$13924 ( \14792 , \13416 , \13698 );
not \U$13925 ( \14793 , \13322_nR2a51 );
and \U$13926 ( \14794 , \13534 , \14793 );
and \U$13927 ( \14795 , \13175_nR2b34 , \13702 );
nor \U$13928 ( \14796 , \14792 , \14794 , \14795 );
xor \U$13929 ( \14797 , \14791 , \14796 );
and \U$13930 ( \14798 , \14797 , \12440 );
and \U$13931 ( \14799 , \14791 , \14796 );
or \U$13932 ( \14800 , \14798 , \14799 );
and \U$13933 ( \14801 , \14069_nR2626 , \12803 );
or \U$13934 ( \14802 , \12733 , \13826_nR26a6 );
nand \U$13935 ( \14803 , \14802 , \12891 );
nand \U$13936 ( \14804 , \14069_nR2626 , \12801 );
and \U$13937 ( \14805 , \14803 , \14804 );
and \U$13938 ( \14806 , \13826_nR26a6 , \12895 );
nor \U$13939 ( \14807 , \14801 , \14805 , \14806 );
nand \U$13940 ( \14808 , \13858_nR274c , \13018 );
or \U$13941 ( \14809 , \12913 , \13575_nR27ee );
nand \U$13942 ( \14810 , \14809 , \13187 );
and \U$13943 ( \14811 , \14808 , \14810 );
and \U$13944 ( \14812 , \13190 , \13575_nR27ee );
and \U$13945 ( \14813 , \13858_nR274c , \13021 );
nor \U$13946 ( \14814 , \14811 , \14812 , \14813 );
xor \U$13947 ( \14815 , \14807 , \14814 );
and \U$13948 ( \14816 , \14172_nR25a7 , \12712 );
or \U$13949 ( \14817 , \12562 , \14358_nR2538 );
nand \U$13950 ( \14818 , \14817 , \12658 );
nand \U$13951 ( \14819 , \14172_nR25a7 , \12651 );
and \U$13952 ( \14820 , \14818 , \14819 );
and \U$13953 ( \14821 , \14358_nR2538 , \12654 );
nor \U$13954 ( \14822 , \14816 , \14820 , \14821 );
and \U$13955 ( \14823 , \14815 , \14822 );
and \U$13956 ( \14824 , \14807 , \14814 );
or \U$13957 ( \14825 , \14823 , \14824 );
xor \U$13958 ( \14826 , \14800 , \14825 );
xor \U$13959 ( \14827 , \14736 , \14743 );
xor \U$13960 ( \14828 , \14827 , \14751 );
and \U$13961 ( \14829 , \14826 , \14828 );
and \U$13962 ( \14830 , \14800 , \14825 );
or \U$13963 ( \14831 , \14829 , \14830 );
xor \U$13964 ( \14832 , \14706 , \14728 );
xor \U$13965 ( \14833 , \14832 , \14754 );
xor \U$13966 ( \14834 , \14831 , \14833 );
xor \U$13967 ( \14835 , \14626 , \14630 );
xor \U$13968 ( \14836 , \14835 , \12387 );
xor \U$13969 ( \14837 , \14762 , \14769 );
xor \U$13970 ( \14838 , \14836 , \14837 );
and \U$13971 ( \14839 , \14834 , \14838 );
and \U$13972 ( \14840 , \14831 , \14833 );
or \U$13973 ( \14841 , \14839 , \14840 );
xor \U$13974 ( \14842 , \14757 , \14759 );
xor \U$13975 ( \14843 , \14842 , \14774 );
xor \U$13976 ( \14844 , \14841 , \14843 );
xnor \U$13977 ( \14845 , \14698 , \14696 );
xor \U$13978 ( \14846 , \14844 , \14845 );
not \U$13979 ( \14847 , \14846 );
xor \U$13980 ( \14848 , \14831 , \14833 );
xor \U$13981 ( \14849 , \14848 , \14838 );
nand \U$13982 ( \14850 , \13575_nR27ee , \13248 );
or \U$13983 ( \14851 , \13213 , \13607_nR28bb );
nand \U$13984 ( \14852 , \14851 , \13445 );
and \U$13985 ( \14853 , \14850 , \14852 );
and \U$13986 ( \14854 , \13448 , \13607_nR28bb );
and \U$13987 ( \14855 , \13575_nR27ee , \13251 );
nor \U$13988 ( \14856 , \14853 , \14854 , \14855 );
not \U$13989 ( \14857 , \14856 );
and \U$13990 ( \14858 , \14793 , \13698 );
not \U$13991 ( \14859 , \13388_nR2979 );
and \U$13992 ( \14860 , \13534 , \14859 );
and \U$13993 ( \14861 , \13322_nR2a51 , \13702 );
nor \U$13994 ( \14862 , \14858 , \14860 , \14861 );
not \U$13995 ( \14863 , \14862 );
and \U$13996 ( \14864 , \14857 , \14863 );
and \U$13997 ( \14865 , \14856 , \14862 );
nand \U$13998 ( \14866 , \13826_nR26a6 , \13018 );
or \U$13999 ( \14867 , \12913 , \13858_nR274c );
nand \U$14000 ( \14868 , \14867 , \13187 );
and \U$14001 ( \14869 , \14866 , \14868 );
and \U$14002 ( \14870 , \13190 , \13858_nR274c );
and \U$14003 ( \14871 , \13826_nR26a6 , \13021 );
nor \U$14004 ( \14872 , \14869 , \14870 , \14871 );
nor \U$14005 ( \14873 , \14865 , \14872 );
nor \U$14006 ( \14874 , \14864 , \14873 );
xor \U$14007 ( \14875 , \14807 , \14814 );
xor \U$14008 ( \14876 , \14875 , \14822 );
and \U$14009 ( \14877 , \14874 , \14876 );
and \U$14010 ( \14878 , \14413_nR2430 , \12512 );
not \U$14011 ( \14879 , \14413_nR2430 );
and \U$14012 ( \14880 , \14879 , \12484 );
not \U$14013 ( \14881 , \12516 );
nor \U$14014 ( \14882 , \14878 , \14880 , \14881 );
xor \U$14015 ( \14883 , \14807 , \14814 );
xor \U$14016 ( \14884 , \14883 , \14822 );
and \U$14017 ( \14885 , \14882 , \14884 );
and \U$14018 ( \14886 , \14874 , \14882 );
or \U$14019 ( \14887 , \14877 , \14885 , \14886 );
xor \U$14020 ( \14888 , \14713 , \14717 );
xor \U$14021 ( \14889 , \14888 , \14725 );
xor \U$14022 ( \14890 , \14887 , \14889 );
xor \U$14023 ( \14891 , \14800 , \14825 );
xor \U$14024 ( \14892 , \14891 , \14828 );
and \U$14025 ( \14893 , \14890 , \14892 );
and \U$14026 ( \14894 , \14887 , \14889 );
or \U$14027 ( \14895 , \14893 , \14894 );
nor \U$14028 ( \14896 , \14849 , \14895 );
xor \U$14029 ( \14897 , \14847 , \14896 );
and \U$14030 ( \14898 , \14849 , \14895 );
nor \U$14031 ( \14899 , \14898 , \14896 );
xor \U$14032 ( \14900 , \14887 , \14889 );
xor \U$14033 ( \14901 , \14900 , \14892 );
and \U$14034 ( \14902 , \14172_nR25a7 , \12803 );
or \U$14035 ( \14903 , \12733 , \14069_nR2626 );
nand \U$14036 ( \14904 , \14903 , \12891 );
nand \U$14037 ( \14905 , \14172_nR25a7 , \12801 );
and \U$14038 ( \14906 , \14904 , \14905 );
and \U$14039 ( \14907 , \14069_nR2626 , \12895 );
nor \U$14040 ( \14908 , \14902 , \14906 , \14907 );
nand \U$14041 ( \14909 , \13858_nR274c , \13248 );
or \U$14042 ( \14910 , \13213 , \13575_nR27ee );
nand \U$14043 ( \14911 , \14910 , \13445 );
and \U$14044 ( \14912 , \14909 , \14911 );
and \U$14045 ( \14913 , \13448 , \13575_nR27ee );
and \U$14046 ( \14914 , \13858_nR274c , \13251 );
nor \U$14047 ( \14915 , \14912 , \14913 , \14914 );
and \U$14048 ( \14916 , \14859 , \13698 );
not \U$14049 ( \14917 , \13607_nR28bb );
and \U$14050 ( \14918 , \13534 , \14917 );
and \U$14051 ( \14919 , \13388_nR2979 , \13702 );
nor \U$14052 ( \14920 , \14916 , \14918 , \14919 );
xor \U$14053 ( \14921 , \14915 , \14920 );
and \U$14054 ( \14922 , \14921 , \12562 );
and \U$14055 ( \14923 , \14915 , \14920 );
or \U$14056 ( \14924 , \14922 , \14923 );
xor \U$14057 ( \14925 , \14908 , \14924 );
and \U$14058 ( \14926 , \14358_nR2538 , \12803 );
or \U$14059 ( \14927 , \12733 , \14172_nR25a7 );
nand \U$14060 ( \14928 , \14927 , \12891 );
nand \U$14061 ( \14929 , \14358_nR2538 , \12801 );
and \U$14062 ( \14930 , \14928 , \14929 );
and \U$14063 ( \14931 , \14172_nR25a7 , \12895 );
nor \U$14064 ( \14932 , \14926 , \14930 , \14931 );
nand \U$14065 ( \14933 , \14069_nR2626 , \13018 );
or \U$14066 ( \14934 , \12913 , \13826_nR26a6 );
nand \U$14067 ( \14935 , \14934 , \13187 );
and \U$14068 ( \14936 , \14933 , \14935 );
and \U$14069 ( \14937 , \13190 , \13826_nR26a6 );
and \U$14070 ( \14938 , \14069_nR2626 , \13021 );
nor \U$14071 ( \14939 , \14936 , \14937 , \14938 );
xor \U$14072 ( \14940 , \14932 , \14939 );
and \U$14073 ( \14941 , \12712 , \14413_nR2430 );
nand \U$14074 ( \14942 , \14413_nR2430 , \12651 );
and \U$14075 ( \14943 , \12656 , \14942 );
nor \U$14076 ( \14944 , \14941 , \14943 );
and \U$14077 ( \14945 , \14940 , \14944 );
and \U$14078 ( \14946 , \14932 , \14939 );
or \U$14079 ( \14947 , \14945 , \14946 );
and \U$14080 ( \14948 , \14925 , \14947 );
and \U$14081 ( \14949 , \14908 , \14924 );
or \U$14082 ( \14950 , \14948 , \14949 );
xor \U$14083 ( \14951 , \14791 , \14796 );
xor \U$14084 ( \14952 , \14951 , \12440 );
nand \U$14085 ( \14953 , \14950 , \14952 );
not \U$14086 ( \14954 , \14856 );
xor \U$14087 ( \14955 , \14862 , \14872 );
not \U$14088 ( \14956 , \14955 );
or \U$14089 ( \14957 , \14954 , \14956 );
or \U$14090 ( \14958 , \14955 , \14856 );
nand \U$14091 ( \14959 , \14957 , \14958 );
not \U$14092 ( \14960 , \14358_nR2538 );
or \U$14093 ( \14961 , \12784 , \14960 );
or \U$14094 ( \14962 , \14879 , \12786 );
or \U$14095 ( \14963 , \12711 , \14960 );
or \U$14096 ( \14964 , \12562 , \14413_nR2430 );
nand \U$14097 ( \14965 , \14964 , \12658 );
nand \U$14098 ( \14966 , \14963 , \14965 );
nand \U$14099 ( \14967 , \14961 , \14962 , \14966 );
and \U$14100 ( \14968 , \14959 , \14967 );
and \U$14101 ( \14969 , \14953 , \14968 );
nor \U$14102 ( \14970 , \14952 , \14950 );
nor \U$14103 ( \14971 , \14969 , \14970 );
nor \U$14104 ( \14972 , \14901 , \14971 );
xor \U$14105 ( \14973 , \14899 , \14972 );
not \U$14106 ( \14974 , \14968 );
not \U$14107 ( \14975 , \14970 );
nand \U$14108 ( \14976 , \14975 , \14953 );
not \U$14109 ( \14977 , \14976 );
or \U$14110 ( \14978 , \14974 , \14977 );
or \U$14111 ( \14979 , \14976 , \14968 );
nand \U$14112 ( \14980 , \14978 , \14979 );
xor \U$14113 ( \14981 , \14807 , \14814 );
xor \U$14114 ( \14982 , \14981 , \14822 );
xor \U$14115 ( \14983 , \14874 , \14882 );
xor \U$14116 ( \14984 , \14982 , \14983 );
not \U$14117 ( \14985 , \14984 );
xor \U$14118 ( \14986 , \14980 , \14985 );
xor \U$14119 ( \14987 , \14908 , \14924 );
xor \U$14120 ( \14988 , \14987 , \14947 );
nand \U$14121 ( \14989 , \13826_nR26a6 , \13248 );
or \U$14122 ( \14990 , \13213 , \13858_nR274c );
nand \U$14123 ( \14991 , \14990 , \13445 );
and \U$14124 ( \14992 , \14989 , \14991 );
and \U$14125 ( \14993 , \13448 , \13858_nR274c );
and \U$14126 ( \14994 , \13826_nR26a6 , \13251 );
nor \U$14127 ( \14995 , \14992 , \14993 , \14994 );
not \U$14128 ( \14996 , \14995 );
and \U$14129 ( \14997 , \14917 , \13698 );
not \U$14130 ( \14998 , \13575_nR27ee );
and \U$14131 ( \14999 , \13534 , \14998 );
and \U$14132 ( \15000 , \13607_nR28bb , \13702 );
nor \U$14133 ( \15001 , \14997 , \14999 , \15000 );
not \U$14134 ( \15002 , \15001 );
and \U$14135 ( \15003 , \14996 , \15002 );
and \U$14136 ( \15004 , \14995 , \15001 );
nand \U$14137 ( \15005 , \14172_nR25a7 , \13018 );
or \U$14138 ( \15006 , \12913 , \14069_nR2626 );
nand \U$14139 ( \15007 , \15006 , \13187 );
and \U$14140 ( \15008 , \15005 , \15007 );
and \U$14141 ( \15009 , \13190 , \14069_nR2626 );
and \U$14142 ( \15010 , \14172_nR25a7 , \13021 );
nor \U$14143 ( \15011 , \15008 , \15009 , \15010 );
nor \U$14144 ( \15012 , \15004 , \15011 );
nor \U$14145 ( \15013 , \15003 , \15012 );
xor \U$14146 ( \15014 , \14915 , \14920 );
xor \U$14147 ( \15015 , \15014 , \12562 );
and \U$14148 ( \15016 , \15013 , \15015 );
xor \U$14149 ( \15017 , \14932 , \14939 );
xor \U$14150 ( \15018 , \15017 , \14944 );
xor \U$14151 ( \15019 , \14915 , \14920 );
xor \U$14152 ( \15020 , \15019 , \12562 );
and \U$14153 ( \15021 , \15018 , \15020 );
and \U$14154 ( \15022 , \15013 , \15018 );
or \U$14155 ( \15023 , \15016 , \15021 , \15022 );
nand \U$14156 ( \15024 , \14988 , \15023 );
xor \U$14157 ( \15025 , \14959 , \14967 );
and \U$14158 ( \15026 , \15024 , \15025 );
nor \U$14159 ( \15027 , \15023 , \14988 );
nor \U$14160 ( \15028 , \15026 , \15027 );
not \U$14161 ( \15029 , \15028 );
xor \U$14162 ( \15030 , \14986 , \15029 );
not \U$14163 ( \15031 , \15024 );
nor \U$14164 ( \15032 , \15031 , \15027 );
not \U$14165 ( \15033 , \15032 );
not \U$14166 ( \15034 , \15025 );
and \U$14167 ( \15035 , \15033 , \15034 );
and \U$14168 ( \15036 , \15032 , \15025 );
nor \U$14169 ( \15037 , \15035 , \15036 );
xor \U$14170 ( \15038 , \14915 , \14920 );
xor \U$14171 ( \15039 , \15038 , \12562 );
xor \U$14172 ( \15040 , \15013 , \15018 );
xor \U$14173 ( \15041 , \15039 , \15040 );
nand \U$14174 ( \15042 , \14069_nR2626 , \13248 );
or \U$14175 ( \15043 , \13213 , \13826_nR26a6 );
nand \U$14176 ( \15044 , \15043 , \13445 );
and \U$14177 ( \15045 , \15042 , \15044 );
and \U$14178 ( \15046 , \13448 , \13826_nR26a6 );
and \U$14179 ( \15047 , \14069_nR2626 , \13251 );
nor \U$14180 ( \15048 , \15045 , \15046 , \15047 );
and \U$14181 ( \15049 , \14998 , \13698 );
not \U$14182 ( \15050 , \13858_nR274c );
and \U$14183 ( \15051 , \13534 , \15050 );
and \U$14184 ( \15052 , \13575_nR27ee , \13702 );
nor \U$14185 ( \15053 , \15049 , \15051 , \15052 );
xor \U$14186 ( \15054 , \15048 , \15053 );
and \U$14187 ( \15055 , \15054 , \12733 );
and \U$14188 ( \15056 , \15048 , \15053 );
or \U$14189 ( \15057 , \15055 , \15056 );
and \U$14190 ( \15058 , \14413_nR2430 , \12803 );
or \U$14191 ( \15059 , \12733 , \14358_nR2538 );
nand \U$14192 ( \15060 , \15059 , \12891 );
nand \U$14193 ( \15061 , \14413_nR2430 , \12801 );
and \U$14194 ( \15062 , \15060 , \15061 );
and \U$14195 ( \15063 , \14358_nR2538 , \12895 );
nor \U$14196 ( \15064 , \15058 , \15062 , \15063 );
nand \U$14197 ( \15065 , \15057 , \15064 );
or \U$14198 ( \15066 , \13022 , \14960 );
or \U$14199 ( \15067 , \12913 , \14172_nR25a7 );
nand \U$14200 ( \15068 , \15067 , \13187 );
nand \U$14201 ( \15069 , \14358_nR2538 , \13018 );
and \U$14202 ( \15070 , \15068 , \15069 );
and \U$14203 ( \15071 , \14172_nR25a7 , \13190 );
nor \U$14204 ( \15072 , \15070 , \15071 );
nand \U$14205 ( \15073 , \15066 , \15072 );
or \U$14206 ( \15074 , \13029 , \14879 );
or \U$14207 ( \15075 , \14413_nR2430 , \12733 );
nand \U$14208 ( \15076 , \15074 , \15075 , \12891 );
and \U$14209 ( \15077 , \15073 , \15076 );
and \U$14210 ( \15078 , \15065 , \15077 );
nor \U$14211 ( \15079 , \15064 , \15057 );
nor \U$14212 ( \15080 , \15078 , \15079 );
nor \U$14213 ( \15081 , \15041 , \15080 );
xor \U$14214 ( \15082 , \15037 , \15081 );
xor \U$14215 ( \15083 , \15073 , \15076 );
not \U$14216 ( \15084 , \15083 );
xor \U$14217 ( \15085 , \15048 , \15053 );
xor \U$14218 ( \15086 , \15085 , \12733 );
nand \U$14219 ( \15087 , \14172_nR25a7 , \13248 );
or \U$14220 ( \15088 , \13213 , \14069_nR2626 );
nand \U$14221 ( \15089 , \15088 , \13445 );
and \U$14222 ( \15090 , \15087 , \15089 );
and \U$14223 ( \15091 , \13448 , \14069_nR2626 );
and \U$14224 ( \15092 , \14172_nR25a7 , \13251 );
nor \U$14225 ( \15093 , \15090 , \15091 , \15092 );
and \U$14226 ( \15094 , \15050 , \13698 );
not \U$14227 ( \15095 , \13826_nR26a6 );
and \U$14228 ( \15096 , \13534 , \15095 );
and \U$14229 ( \15097 , \13858_nR274c , \13702 );
nor \U$14230 ( \15098 , \15094 , \15096 , \15097 );
xor \U$14231 ( \15099 , \15093 , \15098 );
nand \U$14232 ( \15100 , \14413_nR2430 , \13018 );
or \U$14233 ( \15101 , \12913 , \14358_nR2538 );
nand \U$14234 ( \15102 , \15101 , \13187 );
and \U$14235 ( \15103 , \15100 , \15102 );
and \U$14236 ( \15104 , \13190 , \14358_nR2538 );
and \U$14237 ( \15105 , \14413_nR2430 , \13021 );
nor \U$14238 ( \15106 , \15103 , \15104 , \15105 );
and \U$14239 ( \15107 , \15099 , \15106 );
and \U$14240 ( \15108 , \15093 , \15098 );
or \U$14241 ( \15109 , \15107 , \15108 );
nand \U$14242 ( \15110 , \15086 , \15109 );
not \U$14243 ( \15111 , \15110 );
nor \U$14244 ( \15112 , \15109 , \15086 );
nor \U$14245 ( \15113 , \15111 , \15112 );
not \U$14246 ( \15114 , \15113 );
and \U$14247 ( \15115 , \15084 , \15114 );
and \U$14248 ( \15116 , \15083 , \15113 );
nor \U$14249 ( \15117 , \15115 , \15116 );
xor \U$14250 ( \15118 , \15093 , \15098 );
xor \U$14251 ( \15119 , \15118 , \15106 );
nand \U$14252 ( \15120 , \14358_nR2538 , \13248 );
or \U$14253 ( \15121 , \13213 , \14172_nR25a7 );
nand \U$14254 ( \15122 , \15121 , \13445 );
and \U$14255 ( \15123 , \15120 , \15122 );
and \U$14256 ( \15124 , \13448 , \14172_nR25a7 );
and \U$14257 ( \15125 , \14358_nR2538 , \13251 );
nor \U$14258 ( \15126 , \15123 , \15124 , \15125 );
and \U$14259 ( \15127 , \15095 , \13698 );
not \U$14260 ( \15128 , \14069_nR2626 );
and \U$14261 ( \15129 , \13534 , \15128 );
and \U$14262 ( \15130 , \13826_nR26a6 , \13702 );
nor \U$14263 ( \15131 , \15127 , \15129 , \15130 );
xor \U$14264 ( \15132 , \15126 , \15131 );
and \U$14265 ( \15133 , \15132 , \12913 );
and \U$14266 ( \15134 , \15126 , \15131 );
or \U$14267 ( \15135 , \15133 , \15134 );
nor \U$14268 ( \15136 , \15119 , \15135 );
xor \U$14269 ( \15137 , \15117 , \15136 );
not \U$14270 ( \15138 , \14172_nR25a7 );
or \U$14271 ( \15139 , \13701 , \15138 );
or \U$14272 ( \15140 , \14172_nR25a7 , \13536 );
or \U$14273 ( \15141 , \14358_nR2538 , \13535 );
nand \U$14274 ( \15142 , \15139 , \15140 , \15141 );
xor \U$14275 ( \15143 , \15142 , \13250 );
or \U$14276 ( \15144 , \13701 , \14960 );
or \U$14277 ( \15145 , \14358_nR2538 , \13536 );
or \U$14278 ( \15146 , \14413_nR2430 , \13535 );
nand \U$14279 ( \15147 , \15144 , \15145 , \15146 );
nand \U$14280 ( \15148 , \14413_nR2430 , \13533 );
and \U$14281 ( \15149 , \15147 , \13208 , \15148 );
xor \U$14282 ( \15150 , \15143 , \15149 );
not \U$14283 ( \15151 , \13448 );
or \U$14284 ( \15152 , \15151 , \14879 );
or \U$14285 ( \15153 , \14413_nR2430 , \13213 );
nand \U$14286 ( \15154 , \15152 , \15153 , \13445 );
and \U$14287 ( \15155 , \15150 , \15154 );
and \U$14288 ( \15156 , \15143 , \15149 );
or \U$14289 ( \15157 , \15155 , \15156 );
and \U$14290 ( \15158 , \15142 , \13250 );
xor \U$14291 ( \15159 , \15157 , \15158 );
nand \U$14292 ( \15160 , \14413_nR2430 , \13248 );
or \U$14293 ( \15161 , \13213 , \14358_nR2538 );
nand \U$14294 ( \15162 , \15161 , \13445 );
and \U$14295 ( \15163 , \15160 , \15162 );
and \U$14296 ( \15164 , \13448 , \14358_nR2538 );
and \U$14297 ( \15165 , \14413_nR2430 , \13251 );
nor \U$14298 ( \15166 , \15163 , \15164 , \15165 );
and \U$14299 ( \15167 , \15128 , \13698 );
and \U$14300 ( \15168 , \13534 , \15138 );
and \U$14301 ( \15169 , \14069_nR2626 , \13702 );
nor \U$14302 ( \15170 , \15167 , \15168 , \15169 );
and \U$14303 ( \15171 , \15166 , \15170 );
nor \U$14304 ( \15172 , \15166 , \15170 );
nor \U$14305 ( \15173 , \15171 , \15172 );
and \U$14306 ( \15174 , \15159 , \15173 );
and \U$14307 ( \15175 , \15157 , \15158 );
or \U$14308 ( \15176 , \15174 , \15175 );
xor \U$14309 ( \15177 , \15176 , \15172 );
and \U$14310 ( \15178 , \14413_nR2430 , \13190 );
and \U$14311 ( \15179 , \14879 , \13020 );
not \U$14312 ( \15180 , \13187 );
nor \U$14313 ( \15181 , \15178 , \15179 , \15180 );
xor \U$14314 ( \15182 , \15126 , \15131 );
xor \U$14315 ( \15183 , \15182 , \12913 );
and \U$14316 ( \15184 , \15181 , \15183 );
nor \U$14317 ( \15185 , \15181 , \15183 );
nor \U$14318 ( \15186 , \15184 , \15185 );
and \U$14319 ( \15187 , \15177 , \15186 );
and \U$14320 ( \15188 , \15176 , \15172 );
or \U$14321 ( \15189 , \15187 , \15188 );
xor \U$14322 ( \15190 , \15189 , \15185 );
and \U$14323 ( \15191 , \15119 , \15135 );
nor \U$14324 ( \15192 , \15191 , \15136 );
and \U$14325 ( \15193 , \15190 , \15192 );
and \U$14326 ( \15194 , \15189 , \15185 );
or \U$14327 ( \15195 , \15193 , \15194 );
and \U$14328 ( \15196 , \15137 , \15195 );
and \U$14329 ( \15197 , \15117 , \15136 );
or \U$14330 ( \15198 , \15196 , \15197 );
and \U$14331 ( \15199 , \15083 , \15110 );
nor \U$14332 ( \15200 , \15199 , \15112 );
not \U$14333 ( \15201 , \15200 );
xor \U$14334 ( \15202 , \15198 , \15201 );
not \U$14335 ( \15203 , \14995 );
xor \U$14336 ( \15204 , \15001 , \15011 );
not \U$14337 ( \15205 , \15204 );
or \U$14338 ( \15206 , \15203 , \15205 );
or \U$14339 ( \15207 , \15204 , \14995 );
nand \U$14340 ( \15208 , \15206 , \15207 );
not \U$14341 ( \15209 , \15077 );
not \U$14342 ( \15210 , \15079 );
nand \U$14343 ( \15211 , \15210 , \15065 );
not \U$14344 ( \15212 , \15211 );
or \U$14345 ( \15213 , \15209 , \15212 );
or \U$14346 ( \15214 , \15211 , \15077 );
nand \U$14347 ( \15215 , \15213 , \15214 );
xor \U$14348 ( \15216 , \15208 , \15215 );
and \U$14349 ( \15217 , \15202 , \15216 );
and \U$14350 ( \15218 , \15198 , \15201 );
or \U$14351 ( \15219 , \15217 , \15218 );
and \U$14352 ( \15220 , \15208 , \15215 );
xor \U$14353 ( \15221 , \15219 , \15220 );
and \U$14354 ( \15222 , \15041 , \15080 );
nor \U$14355 ( \15223 , \15222 , \15081 );
and \U$14356 ( \15224 , \15221 , \15223 );
and \U$14357 ( \15225 , \15219 , \15220 );
or \U$14358 ( \15226 , \15224 , \15225 );
and \U$14359 ( \15227 , \15082 , \15226 );
and \U$14360 ( \15228 , \15037 , \15081 );
or \U$14361 ( \15229 , \15227 , \15228 );
and \U$14362 ( \15230 , \15030 , \15229 );
and \U$14363 ( \15231 , \14986 , \15029 );
or \U$14364 ( \15232 , \15230 , \15231 );
and \U$14365 ( \15233 , \14980 , \14985 );
xor \U$14366 ( \15234 , \15232 , \15233 );
and \U$14367 ( \15235 , \14901 , \14971 );
nor \U$14368 ( \15236 , \15235 , \14972 );
and \U$14369 ( \15237 , \15234 , \15236 );
and \U$14370 ( \15238 , \15232 , \15233 );
or \U$14371 ( \15239 , \15237 , \15238 );
and \U$14372 ( \15240 , \14973 , \15239 );
and \U$14373 ( \15241 , \14899 , \14972 );
or \U$14374 ( \15242 , \15240 , \15241 );
and \U$14375 ( \15243 , \14897 , \15242 );
and \U$14376 ( \15244 , \14847 , \14896 );
or \U$14377 ( \15245 , \15243 , \15244 );
xor \U$14378 ( \15246 , \14841 , \14843 );
and \U$14379 ( \15247 , \15246 , \14845 );
and \U$14380 ( \15248 , \14841 , \14843 );
or \U$14381 ( \15249 , \15247 , \15248 );
xor \U$14382 ( \15250 , \14699 , \14777 );
xor \U$14383 ( \15251 , \15250 , \14780 );
nand \U$14384 ( \15252 , \15249 , \15251 );
and \U$14385 ( \15253 , \15245 , \15252 );
nor \U$14386 ( \15254 , \15251 , \15249 );
nor \U$14387 ( \15255 , \15253 , \15254 );
and \U$14388 ( \15256 , \14784 , \15255 );
and \U$14389 ( \15257 , \14694 , \14783 );
or \U$14390 ( \15258 , \15256 , \15257 );
not \U$14391 ( \15259 , \15258 );
and \U$14392 ( \15260 , \14687 , \15259 );
and \U$14393 ( \15261 , \14684 , \14686 );
or \U$14394 ( \15262 , \15260 , \15261 );
and \U$14395 ( \15263 , \14609 , \15262 );
and \U$14396 ( \15264 , \14515 , \14608 );
or \U$14397 ( \15265 , \15263 , \15264 );
and \U$14398 ( \15266 , \14514 , \15265 );
and \U$14399 ( \15267 , \14504 , \14513 );
or \U$14400 ( \15268 , \15266 , \15267 );
and \U$14401 ( \15269 , \14502 , \15268 );
and \U$14402 ( \15270 , \14319 , \14501 );
or \U$14403 ( \15271 , \15269 , \15270 );
and \U$14404 ( \15272 , \14317 , \15271 );
and \U$14405 ( \15273 , \14314 , \14316 );
or \U$14406 ( \15274 , \15272 , \15273 );
and \U$14407 ( \15275 , \14223 , \15274 );
and \U$14408 ( \15276 , \14039 , \14222 );
or \U$14409 ( \15277 , \15275 , \15276 );
and \U$14410 ( \15278 , \14037 , \15277 );
and \U$14411 ( \15279 , \14034 , \14036 );
or \U$14412 ( \15280 , \15278 , \15279 );
and \U$14413 ( \15281 , \13950 , \15280 );
and \U$14414 ( \15282 , \13776 , \13949 );
or \U$14415 ( \15283 , \15281 , \15282 );
and \U$14416 ( \15284 , \13768 , \13752 );
not \U$14417 ( \15285 , \13768 );
not \U$14418 ( \15286 , \13752 );
and \U$14419 ( \15287 , \15285 , \15286 );
nor \U$14420 ( \15288 , \15287 , \13772 );
nor \U$14421 ( \15289 , \15284 , \15288 );
xor \U$14422 ( \15290 , \13652 , \13657 );
xor \U$14423 ( \15291 , \15290 , \13660 );
nand \U$14424 ( \15292 , \15289 , \15291 );
and \U$14425 ( \15293 , \15283 , \15292 );
nor \U$14426 ( \15294 , \15291 , \15289 );
nor \U$14427 ( \15295 , \15293 , \15294 );
and \U$14428 ( \15296 , \13664 , \15295 );
and \U$14429 ( \15297 , \13496 , \13663 );
or \U$14430 ( \15298 , \15296 , \15297 );
not \U$14431 ( \15299 , \15298 );
and \U$14432 ( \15300 , \13490 , \15299 );
and \U$14433 ( \15301 , \13352 , \13489 );
or \U$14434 ( \15302 , \15300 , \15301 );
and \U$14435 ( \15303 , \13350 , \15302 );
and \U$14436 ( \15304 , \13236 , \13349 );
or \U$14437 ( \15305 , \15303 , \15304 );
and \U$14438 ( \15306 , \13232 , \15305 );
and \U$14439 ( \15307 , \13229 , \13231 );
or \U$14440 ( \15308 , \15306 , \15307 );
and \U$14441 ( \15309 , \13115 , \15308 );
and \U$14442 ( \15310 , \13112 , \13114 );
or \U$14443 ( \15311 , \15309 , \15310 );
and \U$14444 ( \15312 , \13006 , \15311 );
and \U$14445 ( \15313 , \12888 , \13005 );
or \U$14446 ( \15314 , \15312 , \15313 );
and \U$14447 ( \15315 , \12886 , \15314 );
and \U$14448 ( \15316 , \12709 , \12885 );
or \U$14449 ( \15317 , \15315 , \15316 );
and \U$14450 ( \15318 , \12707 , \15317 );
and \U$14451 ( \15319 , \12705 , \12706 );
or \U$14452 ( \15320 , \15318 , \15319 );
not \U$14453 ( \15321 , \15320 );
or \U$14454 ( \15322 , \12596 , \15321 );
or \U$14455 ( \15323 , \15320 , \12595 );
nand \U$14456 ( \15324 , \15322 , \15323 );
buf \U$14457 ( \15325 , \8726 );
buf \U$14458 ( \15326 , \8307 );
_DC r9a1 ( \15327_nR9a1 , \15325 , \15326 );
not \U$14459 ( \15328 , \15327_nR9a1 );
not \U$14460 ( \15329 , \15328 );
buf \U$14461 ( \15330 , \12248 );
buf \U$14462 ( \15331 , \8307 );
_DC r9a3 ( \15332_nR9a3 , \15330 , \15331 );
not \U$14463 ( \15333 , \15332_nR9a3 );
and \U$14464 ( \15334 , \15329 , \15333 );
buf \U$14465 ( \15335 , \8694 );
_DC r9c0 ( \15336_nR9c0 , \15335 , \15326 );
nor \U$14466 ( \15337 , \15334 , \15336_nR9c0 );
buf \U$14467 ( \15338 , \12218 );
_DC r9c2 ( \15339_nR9c2 , \15338 , \15331 );
and \U$14468 ( \15340 , \15337 , \15339_nR9c2 );
and \U$14469 ( \15341 , \15332_nR9a3 , \15328 );
nor \U$14470 ( \15342 , \15340 , \15341 );
buf \U$14471 ( \15343 , \12188 );
_DC r984 ( \15344_nR984 , \15343 , \15331 );
not \U$14472 ( \15345 , \15344_nR984 );
and \U$14473 ( \15346 , \15342 , \15345 );
buf \U$14474 ( \15347 , \8663 );
_DC r982 ( \15348_nR982 , \15347 , \15326 );
or \U$14475 ( \15349 , \15346 , \15348_nR982 );
or \U$14476 ( \15350 , \15345 , \15342 );
nand \U$14477 ( \15351 , \15349 , \15350 );
buf \U$14478 ( \15352 , \12158 );
_DC r965 ( \15353_nR965 , \15352 , \15331 );
and \U$14479 ( \15354 , \15351 , \15353_nR965 );
not \U$14480 ( \15355 , \15351 );
not \U$14481 ( \15356 , \15353_nR965 );
and \U$14482 ( \15357 , \15355 , \15356 );
buf \U$14483 ( \15358 , \8631 );
_DC r963 ( \15359_nR963 , \15358 , \15326 );
nor \U$14484 ( \15360 , \15357 , \15359_nR963 );
nor \U$14485 ( \15361 , \15354 , \15360 );
buf \U$14486 ( \15362 , \12128 );
_DC r946 ( \15363_nR946 , \15362 , \15331 );
not \U$14487 ( \15364 , \15363_nR946 );
buf \U$14488 ( \15365 , \8595 );
_DC r944 ( \15366_nR944 , \15365 , \15326 );
and \U$14489 ( \15367 , \15364 , \15366_nR944 );
or \U$14490 ( \15368 , \15361 , \15367 );
or \U$14491 ( \15369 , \15366_nR944 , \15364 );
nand \U$14492 ( \15370 , \15368 , \15369 );
buf \U$14493 ( \15371 , \12098 );
_DC r927 ( \15372_nR927 , \15371 , \15331 );
and \U$14494 ( \15373 , \15370 , \15372_nR927 );
not \U$14495 ( \15374 , \15370 );
not \U$14496 ( \15375 , \15372_nR927 );
and \U$14497 ( \15376 , \15374 , \15375 );
buf \U$14498 ( \15377 , \8559 );
_DC r925 ( \15378_nR925 , \15377 , \15326 );
nor \U$14499 ( \15379 , \15376 , \15378_nR925 );
nor \U$14500 ( \15380 , \15373 , \15379 );
buf \U$14501 ( \15381 , \8523 );
_DC r906 ( \15382_nR906 , \15381 , \15326 );
or \U$14502 ( \15383 , \15380 , \15382_nR906 );
not \U$14503 ( \15384 , \15382_nR906 );
not \U$14504 ( \15385 , \15380 );
or \U$14505 ( \15386 , \15384 , \15385 );
buf \U$14506 ( \15387 , \12068 );
_DC r908 ( \15388_nR908 , \15387 , \15331 );
nand \U$14507 ( \15389 , \15386 , \15388_nR908 );
nand \U$14508 ( \15390 , \15383 , \15389 );
buf \U$14509 ( \15391 , \12038 );
_DC r8e9 ( \15392_nR8e9 , \15391 , \15331 );
and \U$14510 ( \15393 , \15390 , \15392_nR8e9 );
not \U$14511 ( \15394 , \15390 );
not \U$14512 ( \15395 , \15392_nR8e9 );
and \U$14513 ( \15396 , \15394 , \15395 );
buf \U$14514 ( \15397 , \8487 );
_DC r8e7 ( \15398_nR8e7 , \15397 , \15326 );
nor \U$14515 ( \15399 , \15396 , \15398_nR8e7 );
nor \U$14516 ( \15400 , \15393 , \15399 );
buf \U$14517 ( \15401 , \12008 );
_DC r8ca ( \15402_nR8ca , \15401 , \15331 );
not \U$14518 ( \15403 , \15402_nR8ca );
buf \U$14519 ( \15404 , \8451 );
_DC r8c8 ( \15405_nR8c8 , \15404 , \15326 );
and \U$14520 ( \15406 , \15403 , \15405_nR8c8 );
or \U$14521 ( \15407 , \15400 , \15406 );
or \U$14522 ( \15408 , \15405_nR8c8 , \15403 );
nand \U$14523 ( \15409 , \15407 , \15408 );
buf \U$14524 ( \15410 , \11978 );
_DC r8ab ( \15411_nR8ab , \15410 , \15331 );
and \U$14525 ( \15412 , \15409 , \15411_nR8ab );
not \U$14526 ( \15413 , \15409 );
not \U$14527 ( \15414 , \15411_nR8ab );
and \U$14528 ( \15415 , \15413 , \15414 );
buf \U$14529 ( \15416 , \8415 );
_DC r8a9 ( \15417_nR8a9 , \15416 , \15326 );
nor \U$14530 ( \15418 , \15415 , \15417_nR8a9 );
nor \U$14531 ( \15419 , \15412 , \15418 );
buf \U$14532 ( \15420 , \11948 );
_DC r88c ( \15421_nR88c , \15420 , \15331 );
not \U$14533 ( \15422 , \15421_nR88c );
buf \U$14534 ( \15423 , \8379 );
_DC r88a ( \15424_nR88a , \15423 , \15326 );
and \U$14535 ( \15425 , \15422 , \15424_nR88a );
or \U$14536 ( \15426 , \15419 , \15425 );
or \U$14537 ( \15427 , \15424_nR88a , \15422 );
nand \U$14538 ( \15428 , \15426 , \15427 );
buf \U$14539 ( \15429 , \11918 );
_DC r86d ( \15430_nR86d , \15429 , \15331 );
and \U$14540 ( \15431 , \15428 , \15430_nR86d );
not \U$14541 ( \15432 , \15428 );
not \U$14542 ( \15433 , \15430_nR86d );
and \U$14543 ( \15434 , \15432 , \15433 );
buf \U$14544 ( \15435 , \8343 );
_DC r86b ( \15436_nR86b , \15435 , \15326 );
nor \U$14545 ( \15437 , \15434 , \15436_nR86b );
nor \U$14546 ( \15438 , \15431 , \15437 );
buf \U$14547 ( \15439 , \11887 );
_DC r84e ( \15440_nR84e , \15439 , \15331 );
not \U$14548 ( \15441 , \15440_nR84e );
buf \U$14549 ( \15442 , \8305 );
_DC r84b ( \15443_nR84b , \15442 , \15326 );
and \U$14550 ( \15444 , \15441 , \15443_nR84b );
or \U$14551 ( \15445 , \15438 , \15444 );
or \U$14552 ( \15446 , \15443_nR84b , \15441 );
nand \U$14553 ( \15447 , \15445 , \15446 );
nor \U$14554 ( \15448 , \8215 , RIb55b778_588);
nand \U$14555 ( \15449 , RIb55bb38_596, \15448 );
not \U$14556 ( \15450 , \15449 );
nand \U$14557 ( \15451 , RIb55bac0_595, \15450 );
not \U$14558 ( \15452 , \15451 );
nand \U$14559 ( \15453 , RIb55ba48_594, \15452 );
not \U$14560 ( \15454 , \15453 );
nand \U$14561 ( \15455 , RIb55b9d0_593, \15454 );
nor \U$14562 ( \15456 , \15455 , \8421 );
nand \U$14563 ( \15457 , RIb55b8e0_591, \15456 );
not \U$14564 ( \15458 , \15457 );
nand \U$14565 ( \15459 , RIb55b868_590, \15458 );
not \U$14566 ( \15460 , \15459 );
nand \U$14567 ( \15461 , \15460 , RIb55b7f0_589);
not \U$14568 ( \15462 , \15461 );
not \U$14569 ( \15463 , RIb55c3a8_614);
and \U$14570 ( \15464 , \15462 , \15463 );
and \U$14571 ( \15465 , \15461 , RIb55c3a8_614);
nor \U$14572 ( \15466 , \15464 , \15465 );
buf \U$14573 ( \15467 , \11887 );
buf \U$14574 ( \15468 , \8307 );
_DC r6ad ( \15469_nR6ad , \15467 , \15468 );
or \U$14575 ( \15470 , \15466 , \15469_nR6ad );
buf \U$14576 ( \15471 , \11918 );
_DC r6cb ( \15472_nR6cb , \15471 , \15468 );
not \U$14577 ( \15473 , \15459 );
not \U$14578 ( \15474 , RIb55b7f0_589);
and \U$14579 ( \15475 , \15473 , \15474 );
and \U$14580 ( \15476 , \15459 , RIb55b7f0_589);
nor \U$14581 ( \15477 , \15475 , \15476 );
or \U$14582 ( \15478 , \15472_nR6cb , \15477 );
not \U$14583 ( \15479 , \15472_nR6cb );
not \U$14584 ( \15480 , \15477 );
or \U$14585 ( \15481 , \15479 , \15480 );
buf \U$14586 ( \15482 , \11978 );
_DC r707 ( \15483_nR707 , \15482 , \15468 );
not \U$14587 ( \15484 , \15483_nR707 );
or \U$14588 ( \15485 , \15456 , RIb55b8e0_591);
nand \U$14589 ( \15486 , \15485 , \15457 );
not \U$14590 ( \15487 , \15486 );
or \U$14591 ( \15488 , \15484 , \15487 );
or \U$14592 ( \15489 , \15486 , \15483_nR707 );
buf \U$14593 ( \15490 , \12008 );
_DC r725 ( \15491_nR725 , \15490 , \15468 );
not \U$14594 ( \15492 , \15491_nR725 );
not \U$14595 ( \15493 , \15455 );
not \U$14596 ( \15494 , RIb55b958_592);
and \U$14597 ( \15495 , \15493 , \15494 );
and \U$14598 ( \15496 , \15455 , RIb55b958_592);
nor \U$14599 ( \15497 , \15495 , \15496 );
not \U$14600 ( \15498 , \15497 );
or \U$14601 ( \15499 , \15492 , \15498 );
or \U$14602 ( \15500 , \15497 , \15491_nR725 );
buf \U$14603 ( \15501 , \12038 );
_DC r743 ( \15502_nR743 , \15501 , \15468 );
not \U$14604 ( \15503 , \15502_nR743 );
or \U$14605 ( \15504 , \15454 , RIb55b9d0_593);
nand \U$14606 ( \15505 , \15504 , \15455 );
not \U$14607 ( \15506 , \15505 );
or \U$14608 ( \15507 , \15503 , \15506 );
or \U$14609 ( \15508 , \15505 , \15502_nR743 );
buf \U$14610 ( \15509 , \12068 );
_DC r761 ( \15510_nR761 , \15509 , \15468 );
not \U$14611 ( \15511 , \15510_nR761 );
or \U$14612 ( \15512 , \15452 , RIb55ba48_594);
nand \U$14613 ( \15513 , \15512 , \15453 );
not \U$14614 ( \15514 , \15513 );
or \U$14615 ( \15515 , \15511 , \15514 );
or \U$14616 ( \15516 , \15513 , \15510_nR761 );
buf \U$14617 ( \15517 , \12098 );
_DC r77f ( \15518_nR77f , \15517 , \15468 );
not \U$14618 ( \15519 , \15518_nR77f );
or \U$14619 ( \15520 , \15450 , RIb55bac0_595);
nand \U$14620 ( \15521 , \15520 , \15451 );
not \U$14621 ( \15522 , \15521 );
or \U$14622 ( \15523 , \15519 , \15522 );
or \U$14623 ( \15524 , \15521 , \15518_nR77f );
buf \U$14624 ( \15525 , \12128 );
_DC r79d ( \15526_nR79d , \15525 , \15468 );
not \U$14625 ( \15527 , \15526_nR79d );
buf \U$14626 ( \15528 , \12248 );
_DC r7f7 ( \15529_nR7f7 , \15528 , \15468 );
not \U$14627 ( \15530 , \15529_nR7f7 );
buf \U$14628 ( \15531 , \12218 );
_DC r815 ( \15532_nR815 , \15531 , \15468 );
and \U$14629 ( \15533 , \8697 , \15532_nR815 );
not \U$14630 ( \15534 , \15533 );
or \U$14631 ( \15535 , \15530 , \15534 );
or \U$14632 ( \15536 , \15533 , \15529_nR7f7 );
or \U$14633 ( \15537 , \7913 , RIb55bca0_599);
nand \U$14634 ( \15538 , RIb55bca0_599, \7913 );
nand \U$14635 ( \15539 , \15537 , \15538 );
nand \U$14636 ( \15540 , \15536 , \15539 );
nand \U$14637 ( \15541 , \15535 , \15540 );
buf \U$14638 ( \15542 , \12188 );
_DC r7d9 ( \15543_nR7d9 , \15542 , \15468 );
and \U$14639 ( \15544 , \15541 , \15543_nR7d9 );
and \U$14640 ( \15545 , \15538 , RIb55bc28_598);
nor \U$14641 ( \15546 , \15541 , \15543_nR7d9 );
nor \U$14642 ( \15547 , \15538 , RIb55bc28_598);
nor \U$14643 ( \15548 , \15545 , \15546 , \15547 );
nor \U$14644 ( \15549 , \15544 , \15548 );
not \U$14645 ( \15550 , \8213 );
not \U$14646 ( \15551 , RIb55b778_588);
and \U$14647 ( \15552 , \15550 , \15551 );
nor \U$14648 ( \15553 , \15552 , RIb55bbb0_597);
buf \U$14649 ( \15554 , \12158 );
_DC r7bb ( \15555_nR7bb , \15554 , \15468 );
nor \U$14650 ( \15556 , \15448 , \15553 , \15555_nR7bb );
or \U$14651 ( \15557 , \15549 , \15556 );
or \U$14652 ( \15558 , \15448 , \15553 );
nand \U$14653 ( \15559 , \15558 , \15555_nR7bb );
nand \U$14654 ( \15560 , \15557 , \15559 );
not \U$14655 ( \15561 , \15560 );
or \U$14656 ( \15562 , \15527 , \15561 );
or \U$14657 ( \15563 , \15560 , \15526_nR79d );
or \U$14658 ( \15564 , \15448 , RIb55bb38_596);
nand \U$14659 ( \15565 , \15564 , \15449 );
nand \U$14660 ( \15566 , \15563 , \15565 );
nand \U$14661 ( \15567 , \15562 , \15566 );
nand \U$14662 ( \15568 , \15524 , \15567 );
nand \U$14663 ( \15569 , \15523 , \15568 );
nand \U$14664 ( \15570 , \15516 , \15569 );
nand \U$14665 ( \15571 , \15515 , \15570 );
nand \U$14666 ( \15572 , \15508 , \15571 );
nand \U$14667 ( \15573 , \15507 , \15572 );
nand \U$14668 ( \15574 , \15500 , \15573 );
nand \U$14669 ( \15575 , \15499 , \15574 );
nand \U$14670 ( \15576 , \15489 , \15575 );
nand \U$14671 ( \15577 , \15488 , \15576 );
or \U$14672 ( \15578 , \15458 , RIb55b868_590);
nand \U$14673 ( \15579 , \15578 , \15459 );
buf \U$14674 ( \15580 , \11948 );
_DC r6e9 ( \15581_nR6e9 , \15580 , \15468 );
or \U$14675 ( \15582 , \15579 , \15581_nR6e9 );
and \U$14676 ( \15583 , \15577 , \15582 );
and \U$14677 ( \15584 , \15581_nR6e9 , \15579 );
nor \U$14678 ( \15585 , \15583 , \15584 );
nand \U$14679 ( \15586 , \15481 , \15585 );
nand \U$14680 ( \15587 , \15470 , \15478 , \15586 );
nand \U$14681 ( \15588 , \15469_nR6ad , \15466 );
and \U$14682 ( \15589 , \15447 , \15587 , \8783 , \15588 );
_HMUX r3dc1 ( \15590_nR3dc1 , \11849 , \15324 , \15589 );
buf \U$14683 ( \15591 , \15590_nR3dc1 );
xor \U$14684 ( \15592 , \9200 , \9199 );
not \U$14685 ( \15593 , \15592 );
not \U$14686 ( \15594 , \11843 );
or \U$14687 ( \15595 , \15593 , \15594 );
or \U$14688 ( \15596 , \11843 , \15592 );
nand \U$14689 ( \15597 , \15595 , \15596 );
xor \U$14690 ( \15598 , \12705 , \12706 );
xor \U$14691 ( \15599 , \15598 , \15317 );
_HMUX r3d84 ( \15600_nR3d84 , \15597 , \15599 , \15589 );
buf \U$14692 ( \15601 , \15600_nR3d84 );
not \U$14693 ( \15602 , \11842 );
nand \U$14694 ( \15603 , \15602 , \11840 );
not \U$14695 ( \15604 , \15603 );
not \U$14696 ( \15605 , \11830 );
or \U$14697 ( \15606 , \15604 , \15605 );
or \U$14698 ( \15607 , \11830 , \15603 );
nand \U$14699 ( \15608 , \15606 , \15607 );
xor \U$14700 ( \15609 , \12709 , \12885 );
xor \U$14701 ( \15610 , \15609 , \15314 );
_HMUX r3d54 ( \15611_nR3d54 , \15608 , \15610 , \15589 );
buf \U$14702 ( \15612 , \15611_nR3d54 );
xor \U$14703 ( \15613 , \9393 , \9515 );
xor \U$14704 ( \15614 , \15613 , \11827 );
xor \U$14705 ( \15615 , \12888 , \13005 );
xor \U$14706 ( \15616 , \15615 , \15311 );
_HMUX r3d07 ( \15617_nR3d07 , \15614 , \15616 , \15589 );
buf \U$14707 ( \15618 , \15617_nR3d07 );
xor \U$14708 ( \15619 , \9518 , \9624 );
xor \U$14709 ( \15620 , \15619 , \11824 );
xor \U$14710 ( \15621 , \13112 , \13114 );
xor \U$14711 ( \15622 , \15621 , \15308 );
_HMUX r3c96 ( \15623_nR3c96 , \15620 , \15622 , \15589 );
buf \U$14712 ( \15624 , \15623_nR3c96 );
xor \U$14713 ( \15625 , \9742 , \9744 );
xor \U$14714 ( \15626 , \15625 , \11821 );
xor \U$14715 ( \15627 , \13229 , \13231 );
xor \U$14716 ( \15628 , \15627 , \15305 );
_HMUX r3c30 ( \15629_nR3c30 , \15626 , \15628 , \15589 );
buf \U$14717 ( \15630 , \15629_nR3c30 );
xor \U$14718 ( \15631 , \9749 , \9858 );
xor \U$14719 ( \15632 , \15631 , \11818 );
xor \U$14720 ( \15633 , \13236 , \13349 );
xor \U$14721 ( \15634 , \15633 , \15302 );
_HMUX r3b9b ( \15635_nR3b9b , \15632 , \15634 , \15589 );
buf \U$14722 ( \15636 , \15635_nR3b9b );
xor \U$14723 ( \15637 , \9995 , \9997 );
xor \U$14724 ( \15638 , \15637 , \11815 );
xor \U$14725 ( \15639 , \13352 , \13489 );
xor \U$14726 ( \15640 , \15639 , \15299 );
_HMUX r3afb ( \15641_nR3afb , \15638 , \15640 , \15589 );
buf \U$14727 ( \15642 , \15641_nR3afb );
xor \U$14728 ( \15643 , \10002 , \10159 );
xor \U$14729 ( \15644 , \15643 , \11812 );
xor \U$14730 ( \15645 , \13496 , \13663 );
xor \U$14731 ( \15646 , \15645 , \15295 );
not \U$14732 ( \15647 , \15646 );
_HMUX r3a4f ( \15648_nR3a4f , \15644 , \15647 , \15589 );
buf \U$14733 ( \15649 , \15648_nR3a4f );
xor \U$14734 ( \15650 , \10162 , \10269 );
xor \U$14735 ( \15651 , \15650 , \11809 );
not \U$14736 ( \15652 , \15294 );
nand \U$14737 ( \15653 , \15652 , \15292 );
not \U$14738 ( \15654 , \15653 );
not \U$14739 ( \15655 , \15283 );
or \U$14740 ( \15656 , \15654 , \15655 );
or \U$14741 ( \15657 , \15283 , \15653 );
nand \U$14742 ( \15658 , \15656 , \15657 );
_HMUX r3999 ( \15659_nR3999 , \15651 , \15658 , \15589 );
buf \U$14743 ( \15660 , \15659_nR3999 );
xor \U$14744 ( \15661 , \10272 , \10443 );
xor \U$14745 ( \15662 , \15661 , \11806 );
xor \U$14746 ( \15663 , \13776 , \13949 );
xor \U$14747 ( \15664 , \15663 , \15280 );
_HMUX r38e8 ( \15665_nR38e8 , \15662 , \15664 , \15589 );
buf \U$14748 ( \15666 , \15665_nR38e8 );
xor \U$14749 ( \15667 , \11798 , \11802 );
xnor \U$14750 ( \15668 , \11796 , \15667 );
xor \U$14751 ( \15669 , \14034 , \14036 );
xor \U$14752 ( \15670 , \15669 , \15277 );
_HMUX r381f ( \15671_nR381f , \15668 , \15670 , \15589 );
buf \U$14753 ( \15672 , \15671_nR381f );
not \U$14754 ( \15673 , \11795 );
nand \U$14755 ( \15674 , \15673 , \11793 );
not \U$14756 ( \15675 , \15674 );
not \U$14757 ( \15676 , \11774 );
or \U$14758 ( \15677 , \15675 , \15676 );
or \U$14759 ( \15678 , \11774 , \15674 );
nand \U$14760 ( \15679 , \15677 , \15678 );
xor \U$14761 ( \15680 , \14039 , \14222 );
xor \U$14762 ( \15681 , \15680 , \15274 );
_HMUX r374a ( \15682_nR374a , \15679 , \15681 , \15589 );
buf \U$14763 ( \15683 , \15682_nR374a );
xor \U$14764 ( \15684 , \10713 , \10809 );
xor \U$14765 ( \15685 , \15684 , \11771 );
xor \U$14766 ( \15686 , \14314 , \14316 );
xor \U$14767 ( \15687 , \15686 , \15271 );
_HMUX r3678 ( \15688_nR3678 , \15685 , \15687 , \15589 );
buf \U$14768 ( \15689 , \15688_nR3678 );
xor \U$14769 ( \15690 , \10812 , \10988 );
xor \U$14770 ( \15691 , \15690 , \11768 );
xor \U$14771 ( \15692 , \14319 , \14501 );
xor \U$14772 ( \15693 , \15692 , \15268 );
_HMUX r3576 ( \15694_nR3576 , \15691 , \15693 , \15589 );
buf \U$14773 ( \15695 , \15694_nR3576 );
xor \U$14774 ( \15696 , \10991 , \11000 );
xor \U$14775 ( \15697 , \15696 , \11765 );
xor \U$14776 ( \15698 , \14504 , \14513 );
xor \U$14777 ( \15699 , \15698 , \15265 );
_HMUX r3464 ( \15700_nR3464 , \15697 , \15699 , \15589 );
buf \U$14778 ( \15701 , \15700_nR3464 );
xor \U$14779 ( \15702 , \11003 , \11090 );
xor \U$14780 ( \15703 , \15702 , \11762 );
xor \U$14781 ( \15704 , \14515 , \14608 );
xor \U$14782 ( \15705 , \15704 , \15262 );
_HMUX r333e ( \15706_nR333e , \15703 , \15705 , \15589 );
buf \U$14783 ( \15707 , \15706_nR333e );
xor \U$14784 ( \15708 , \11171 , \11176 );
xor \U$14785 ( \15709 , \15708 , \11759 );
xor \U$14786 ( \15710 , \14684 , \14686 );
xor \U$14787 ( \15711 , \15710 , \15259 );
_HMUX r3236 ( \15712_nR3236 , \15709 , \15711 , \15589 );
buf \U$14788 ( \15713 , \15712_nR3236 );
xor \U$14789 ( \15714 , \11184 , \11271 );
xor \U$14790 ( \15715 , \15714 , \11755 );
not \U$14791 ( \15716 , \15715 );
xor \U$14792 ( \15717 , \14694 , \14783 );
xor \U$14793 ( \15718 , \15717 , \15255 );
not \U$14794 ( \15719 , \15718 );
_HMUX r3115 ( \15720_nR3115 , \15716 , \15719 , \15589 );
buf \U$14795 ( \15721 , \15720_nR3115 );
not \U$14796 ( \15722 , \11754 );
nand \U$14797 ( \15723 , \15722 , \11752 );
not \U$14798 ( \15724 , \15723 );
not \U$14799 ( \15725 , \11741 );
or \U$14800 ( \15726 , \15724 , \15725 );
or \U$14801 ( \15727 , \11741 , \15723 );
nand \U$14802 ( \15728 , \15726 , \15727 );
not \U$14803 ( \15729 , \15254 );
nand \U$14804 ( \15730 , \15729 , \15252 );
not \U$14805 ( \15731 , \15730 );
not \U$14806 ( \15732 , \15245 );
or \U$14807 ( \15733 , \15731 , \15732 );
or \U$14808 ( \15734 , \15245 , \15730 );
nand \U$14809 ( \15735 , \15733 , \15734 );
_HMUX r2ffe ( \15736_nR2ffe , \15728 , \15735 , \15589 );
buf \U$14810 ( \15737 , \15736_nR2ffe );
xor \U$14811 ( \15738 , \11335 , \11386 );
xor \U$14812 ( \15739 , \15738 , \11738 );
xor \U$14813 ( \15740 , \14847 , \14896 );
xor \U$14814 ( \15741 , \15740 , \15242 );
_HMUX r2ee6 ( \15742_nR2ee6 , \15739 , \15741 , \15589 );
buf \U$14815 ( \15743 , \15742_nR2ee6 );
xor \U$14816 ( \15744 , \11389 , \11462 );
xor \U$14817 ( \15745 , \15744 , \11735 );
xor \U$14818 ( \15746 , \14899 , \14972 );
xor \U$14819 ( \15747 , \15746 , \15239 );
_HMUX r2def ( \15748_nR2def , \15745 , \15747 , \15589 );
buf \U$14820 ( \15749 , \15748_nR2def );
xor \U$14821 ( \15750 , \11728 , \11729 );
xor \U$14822 ( \15751 , \15750 , \11732 );
xor \U$14823 ( \15752 , \15232 , \15233 );
xor \U$14824 ( \15753 , \15752 , \15236 );
_HMUX r2cdf ( \15754_nR2cdf , \15751 , \15753 , \15589 );
buf \U$14825 ( \15755 , \15754_nR2cdf );
xor \U$14826 ( \15756 , \11477 , \11518 );
xor \U$14827 ( \15757 , \15756 , \11725 );
xor \U$14828 ( \15758 , \14986 , \15029 );
xor \U$14829 ( \15759 , \15758 , \15229 );
_HMUX r2c00 ( \15760_nR2c00 , \15757 , \15759 , \15589 );
buf \U$14830 ( \15761 , \15760_nR2c00 );
xor \U$14831 ( \15762 , \11526 , \11572 );
xor \U$14832 ( \15763 , \15762 , \11722 );
xor \U$14833 ( \15764 , \15037 , \15081 );
xor \U$14834 ( \15765 , \15764 , \15226 );
_HMUX r2af2 ( \15766_nR2af2 , \15763 , \15765 , \15589 );
buf \U$14835 ( \15767 , \15766_nR2af2 );
xor \U$14836 ( \15768 , \11716 , \11579 );
xor \U$14837 ( \15769 , \15768 , \11719 );
xor \U$14838 ( \15770 , \15219 , \15220 );
xor \U$14839 ( \15771 , \15770 , \15223 );
_HMUX r2a16 ( \15772_nR2a16 , \15769 , \15771 , \15589 );
buf \U$14840 ( \15773 , \15772_nR2a16 );
xor \U$14841 ( \15774 , \11580 , \11621 );
xor \U$14842 ( \15775 , \15774 , \11713 );
xor \U$14843 ( \15776 , \15198 , \15201 );
xor \U$14844 ( \15777 , \15776 , \15216 );
_HMUX r2937 ( \15778_nR2937 , \15775 , \15777 , \15589 );
buf \U$14845 ( \15779 , \15778_nR2937 );
endmodule

